module tt_um_urish_spell (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire clknet_leaf_0_clk;
 wire \delay_counter[0] ;
 wire \delay_counter[1] ;
 wire \delay_counter[2] ;
 wire \delay_counter[3] ;
 wire \delay_counter[4] ;
 wire \delay_counter[5] ;
 wire \delay_counter[6] ;
 wire \delay_counter[7] ;
 wire \delay_cycles[0] ;
 wire \delay_cycles[10] ;
 wire \delay_cycles[11] ;
 wire \delay_cycles[12] ;
 wire \delay_cycles[13] ;
 wire \delay_cycles[14] ;
 wire \delay_cycles[15] ;
 wire \delay_cycles[16] ;
 wire \delay_cycles[17] ;
 wire \delay_cycles[18] ;
 wire \delay_cycles[19] ;
 wire \delay_cycles[1] ;
 wire \delay_cycles[20] ;
 wire \delay_cycles[21] ;
 wire \delay_cycles[22] ;
 wire \delay_cycles[23] ;
 wire \delay_cycles[2] ;
 wire \delay_cycles[3] ;
 wire \delay_cycles[4] ;
 wire \delay_cycles[5] ;
 wire \delay_cycles[6] ;
 wire \delay_cycles[7] ;
 wire \delay_cycles[8] ;
 wire \delay_cycles[9] ;
 wire \exec.memory_input[0] ;
 wire \exec.memory_input[1] ;
 wire \exec.memory_input[2] ;
 wire \exec.memory_input[3] ;
 wire \exec.memory_input[4] ;
 wire \exec.memory_input[5] ;
 wire \exec.memory_input[6] ;
 wire \exec.memory_input[7] ;
 wire \exec.opcode[0] ;
 wire \exec.opcode[1] ;
 wire \exec.opcode[2] ;
 wire \exec.opcode[3] ;
 wire \exec.opcode[4] ;
 wire \exec.opcode[5] ;
 wire \exec.opcode[6] ;
 wire \exec.opcode[7] ;
 wire \exec.out_of_order_exec ;
 wire \exec.pc[0] ;
 wire \exec.pc[1] ;
 wire \exec.pc[2] ;
 wire \exec.pc[3] ;
 wire \exec.pc[4] ;
 wire \exec.pc[5] ;
 wire \exec.pc[6] ;
 wire \exec.pc[7] ;
 wire \exec.sp[0] ;
 wire \exec.sp[1] ;
 wire \exec.sp[2] ;
 wire \exec.sp[3] ;
 wire \exec.sp[4] ;
 wire \mem.addr[0] ;
 wire \mem.addr[1] ;
 wire \mem.addr[2] ;
 wire \mem.addr[3] ;
 wire \mem.addr[4] ;
 wire \mem.addr[5] ;
 wire \mem.addr[6] ;
 wire \mem.addr[7] ;
 wire \mem.data_in[0] ;
 wire \mem.data_in[1] ;
 wire \mem.data_in[2] ;
 wire \mem.data_in[3] ;
 wire \mem.data_in[4] ;
 wire \mem.data_in[5] ;
 wire \mem.data_in[6] ;
 wire \mem.data_in[7] ;
 wire \mem.internal_data_out[0] ;
 wire \mem.internal_data_out[1] ;
 wire \mem.internal_data_out[2] ;
 wire \mem.internal_data_out[3] ;
 wire \mem.internal_data_out[4] ;
 wire \mem.internal_data_out[5] ;
 wire \mem.internal_data_out[6] ;
 wire \mem.internal_data_out[7] ;
 wire \mem.internal_data_ready ;
 wire \mem.io_data_out[0] ;
 wire \mem.io_data_out[1] ;
 wire \mem.io_data_out[2] ;
 wire \mem.io_data_out[3] ;
 wire \mem.io_data_out[4] ;
 wire \mem.io_data_out[5] ;
 wire \mem.io_data_out[6] ;
 wire \mem.io_data_out[7] ;
 wire \mem.io_data_ready ;
 wire \mem.mem_internal.code_mem[0][0] ;
 wire \mem.mem_internal.code_mem[0][1] ;
 wire \mem.mem_internal.code_mem[0][2] ;
 wire \mem.mem_internal.code_mem[0][3] ;
 wire \mem.mem_internal.code_mem[0][4] ;
 wire \mem.mem_internal.code_mem[0][5] ;
 wire \mem.mem_internal.code_mem[0][6] ;
 wire \mem.mem_internal.code_mem[0][7] ;
 wire \mem.mem_internal.code_mem[100][0] ;
 wire \mem.mem_internal.code_mem[100][1] ;
 wire \mem.mem_internal.code_mem[100][2] ;
 wire \mem.mem_internal.code_mem[100][3] ;
 wire \mem.mem_internal.code_mem[100][4] ;
 wire \mem.mem_internal.code_mem[100][5] ;
 wire \mem.mem_internal.code_mem[100][6] ;
 wire \mem.mem_internal.code_mem[100][7] ;
 wire \mem.mem_internal.code_mem[101][0] ;
 wire \mem.mem_internal.code_mem[101][1] ;
 wire \mem.mem_internal.code_mem[101][2] ;
 wire \mem.mem_internal.code_mem[101][3] ;
 wire \mem.mem_internal.code_mem[101][4] ;
 wire \mem.mem_internal.code_mem[101][5] ;
 wire \mem.mem_internal.code_mem[101][6] ;
 wire \mem.mem_internal.code_mem[101][7] ;
 wire \mem.mem_internal.code_mem[102][0] ;
 wire \mem.mem_internal.code_mem[102][1] ;
 wire \mem.mem_internal.code_mem[102][2] ;
 wire \mem.mem_internal.code_mem[102][3] ;
 wire \mem.mem_internal.code_mem[102][4] ;
 wire \mem.mem_internal.code_mem[102][5] ;
 wire \mem.mem_internal.code_mem[102][6] ;
 wire \mem.mem_internal.code_mem[102][7] ;
 wire \mem.mem_internal.code_mem[103][0] ;
 wire \mem.mem_internal.code_mem[103][1] ;
 wire \mem.mem_internal.code_mem[103][2] ;
 wire \mem.mem_internal.code_mem[103][3] ;
 wire \mem.mem_internal.code_mem[103][4] ;
 wire \mem.mem_internal.code_mem[103][5] ;
 wire \mem.mem_internal.code_mem[103][6] ;
 wire \mem.mem_internal.code_mem[103][7] ;
 wire \mem.mem_internal.code_mem[104][0] ;
 wire \mem.mem_internal.code_mem[104][1] ;
 wire \mem.mem_internal.code_mem[104][2] ;
 wire \mem.mem_internal.code_mem[104][3] ;
 wire \mem.mem_internal.code_mem[104][4] ;
 wire \mem.mem_internal.code_mem[104][5] ;
 wire \mem.mem_internal.code_mem[104][6] ;
 wire \mem.mem_internal.code_mem[104][7] ;
 wire \mem.mem_internal.code_mem[105][0] ;
 wire \mem.mem_internal.code_mem[105][1] ;
 wire \mem.mem_internal.code_mem[105][2] ;
 wire \mem.mem_internal.code_mem[105][3] ;
 wire \mem.mem_internal.code_mem[105][4] ;
 wire \mem.mem_internal.code_mem[105][5] ;
 wire \mem.mem_internal.code_mem[105][6] ;
 wire \mem.mem_internal.code_mem[105][7] ;
 wire \mem.mem_internal.code_mem[106][0] ;
 wire \mem.mem_internal.code_mem[106][1] ;
 wire \mem.mem_internal.code_mem[106][2] ;
 wire \mem.mem_internal.code_mem[106][3] ;
 wire \mem.mem_internal.code_mem[106][4] ;
 wire \mem.mem_internal.code_mem[106][5] ;
 wire \mem.mem_internal.code_mem[106][6] ;
 wire \mem.mem_internal.code_mem[106][7] ;
 wire \mem.mem_internal.code_mem[107][0] ;
 wire \mem.mem_internal.code_mem[107][1] ;
 wire \mem.mem_internal.code_mem[107][2] ;
 wire \mem.mem_internal.code_mem[107][3] ;
 wire \mem.mem_internal.code_mem[107][4] ;
 wire \mem.mem_internal.code_mem[107][5] ;
 wire \mem.mem_internal.code_mem[107][6] ;
 wire \mem.mem_internal.code_mem[107][7] ;
 wire \mem.mem_internal.code_mem[108][0] ;
 wire \mem.mem_internal.code_mem[108][1] ;
 wire \mem.mem_internal.code_mem[108][2] ;
 wire \mem.mem_internal.code_mem[108][3] ;
 wire \mem.mem_internal.code_mem[108][4] ;
 wire \mem.mem_internal.code_mem[108][5] ;
 wire \mem.mem_internal.code_mem[108][6] ;
 wire \mem.mem_internal.code_mem[108][7] ;
 wire \mem.mem_internal.code_mem[109][0] ;
 wire \mem.mem_internal.code_mem[109][1] ;
 wire \mem.mem_internal.code_mem[109][2] ;
 wire \mem.mem_internal.code_mem[109][3] ;
 wire \mem.mem_internal.code_mem[109][4] ;
 wire \mem.mem_internal.code_mem[109][5] ;
 wire \mem.mem_internal.code_mem[109][6] ;
 wire \mem.mem_internal.code_mem[109][7] ;
 wire \mem.mem_internal.code_mem[10][0] ;
 wire \mem.mem_internal.code_mem[10][1] ;
 wire \mem.mem_internal.code_mem[10][2] ;
 wire \mem.mem_internal.code_mem[10][3] ;
 wire \mem.mem_internal.code_mem[10][4] ;
 wire \mem.mem_internal.code_mem[10][5] ;
 wire \mem.mem_internal.code_mem[10][6] ;
 wire \mem.mem_internal.code_mem[10][7] ;
 wire \mem.mem_internal.code_mem[110][0] ;
 wire \mem.mem_internal.code_mem[110][1] ;
 wire \mem.mem_internal.code_mem[110][2] ;
 wire \mem.mem_internal.code_mem[110][3] ;
 wire \mem.mem_internal.code_mem[110][4] ;
 wire \mem.mem_internal.code_mem[110][5] ;
 wire \mem.mem_internal.code_mem[110][6] ;
 wire \mem.mem_internal.code_mem[110][7] ;
 wire \mem.mem_internal.code_mem[111][0] ;
 wire \mem.mem_internal.code_mem[111][1] ;
 wire \mem.mem_internal.code_mem[111][2] ;
 wire \mem.mem_internal.code_mem[111][3] ;
 wire \mem.mem_internal.code_mem[111][4] ;
 wire \mem.mem_internal.code_mem[111][5] ;
 wire \mem.mem_internal.code_mem[111][6] ;
 wire \mem.mem_internal.code_mem[111][7] ;
 wire \mem.mem_internal.code_mem[112][0] ;
 wire \mem.mem_internal.code_mem[112][1] ;
 wire \mem.mem_internal.code_mem[112][2] ;
 wire \mem.mem_internal.code_mem[112][3] ;
 wire \mem.mem_internal.code_mem[112][4] ;
 wire \mem.mem_internal.code_mem[112][5] ;
 wire \mem.mem_internal.code_mem[112][6] ;
 wire \mem.mem_internal.code_mem[112][7] ;
 wire \mem.mem_internal.code_mem[113][0] ;
 wire \mem.mem_internal.code_mem[113][1] ;
 wire \mem.mem_internal.code_mem[113][2] ;
 wire \mem.mem_internal.code_mem[113][3] ;
 wire \mem.mem_internal.code_mem[113][4] ;
 wire \mem.mem_internal.code_mem[113][5] ;
 wire \mem.mem_internal.code_mem[113][6] ;
 wire \mem.mem_internal.code_mem[113][7] ;
 wire \mem.mem_internal.code_mem[114][0] ;
 wire \mem.mem_internal.code_mem[114][1] ;
 wire \mem.mem_internal.code_mem[114][2] ;
 wire \mem.mem_internal.code_mem[114][3] ;
 wire \mem.mem_internal.code_mem[114][4] ;
 wire \mem.mem_internal.code_mem[114][5] ;
 wire \mem.mem_internal.code_mem[114][6] ;
 wire \mem.mem_internal.code_mem[114][7] ;
 wire \mem.mem_internal.code_mem[115][0] ;
 wire \mem.mem_internal.code_mem[115][1] ;
 wire \mem.mem_internal.code_mem[115][2] ;
 wire \mem.mem_internal.code_mem[115][3] ;
 wire \mem.mem_internal.code_mem[115][4] ;
 wire \mem.mem_internal.code_mem[115][5] ;
 wire \mem.mem_internal.code_mem[115][6] ;
 wire \mem.mem_internal.code_mem[115][7] ;
 wire \mem.mem_internal.code_mem[116][0] ;
 wire \mem.mem_internal.code_mem[116][1] ;
 wire \mem.mem_internal.code_mem[116][2] ;
 wire \mem.mem_internal.code_mem[116][3] ;
 wire \mem.mem_internal.code_mem[116][4] ;
 wire \mem.mem_internal.code_mem[116][5] ;
 wire \mem.mem_internal.code_mem[116][6] ;
 wire \mem.mem_internal.code_mem[116][7] ;
 wire \mem.mem_internal.code_mem[117][0] ;
 wire \mem.mem_internal.code_mem[117][1] ;
 wire \mem.mem_internal.code_mem[117][2] ;
 wire \mem.mem_internal.code_mem[117][3] ;
 wire \mem.mem_internal.code_mem[117][4] ;
 wire \mem.mem_internal.code_mem[117][5] ;
 wire \mem.mem_internal.code_mem[117][6] ;
 wire \mem.mem_internal.code_mem[117][7] ;
 wire \mem.mem_internal.code_mem[118][0] ;
 wire \mem.mem_internal.code_mem[118][1] ;
 wire \mem.mem_internal.code_mem[118][2] ;
 wire \mem.mem_internal.code_mem[118][3] ;
 wire \mem.mem_internal.code_mem[118][4] ;
 wire \mem.mem_internal.code_mem[118][5] ;
 wire \mem.mem_internal.code_mem[118][6] ;
 wire \mem.mem_internal.code_mem[118][7] ;
 wire \mem.mem_internal.code_mem[119][0] ;
 wire \mem.mem_internal.code_mem[119][1] ;
 wire \mem.mem_internal.code_mem[119][2] ;
 wire \mem.mem_internal.code_mem[119][3] ;
 wire \mem.mem_internal.code_mem[119][4] ;
 wire \mem.mem_internal.code_mem[119][5] ;
 wire \mem.mem_internal.code_mem[119][6] ;
 wire \mem.mem_internal.code_mem[119][7] ;
 wire \mem.mem_internal.code_mem[11][0] ;
 wire \mem.mem_internal.code_mem[11][1] ;
 wire \mem.mem_internal.code_mem[11][2] ;
 wire \mem.mem_internal.code_mem[11][3] ;
 wire \mem.mem_internal.code_mem[11][4] ;
 wire \mem.mem_internal.code_mem[11][5] ;
 wire \mem.mem_internal.code_mem[11][6] ;
 wire \mem.mem_internal.code_mem[11][7] ;
 wire \mem.mem_internal.code_mem[120][0] ;
 wire \mem.mem_internal.code_mem[120][1] ;
 wire \mem.mem_internal.code_mem[120][2] ;
 wire \mem.mem_internal.code_mem[120][3] ;
 wire \mem.mem_internal.code_mem[120][4] ;
 wire \mem.mem_internal.code_mem[120][5] ;
 wire \mem.mem_internal.code_mem[120][6] ;
 wire \mem.mem_internal.code_mem[120][7] ;
 wire \mem.mem_internal.code_mem[121][0] ;
 wire \mem.mem_internal.code_mem[121][1] ;
 wire \mem.mem_internal.code_mem[121][2] ;
 wire \mem.mem_internal.code_mem[121][3] ;
 wire \mem.mem_internal.code_mem[121][4] ;
 wire \mem.mem_internal.code_mem[121][5] ;
 wire \mem.mem_internal.code_mem[121][6] ;
 wire \mem.mem_internal.code_mem[121][7] ;
 wire \mem.mem_internal.code_mem[122][0] ;
 wire \mem.mem_internal.code_mem[122][1] ;
 wire \mem.mem_internal.code_mem[122][2] ;
 wire \mem.mem_internal.code_mem[122][3] ;
 wire \mem.mem_internal.code_mem[122][4] ;
 wire \mem.mem_internal.code_mem[122][5] ;
 wire \mem.mem_internal.code_mem[122][6] ;
 wire \mem.mem_internal.code_mem[122][7] ;
 wire \mem.mem_internal.code_mem[123][0] ;
 wire \mem.mem_internal.code_mem[123][1] ;
 wire \mem.mem_internal.code_mem[123][2] ;
 wire \mem.mem_internal.code_mem[123][3] ;
 wire \mem.mem_internal.code_mem[123][4] ;
 wire \mem.mem_internal.code_mem[123][5] ;
 wire \mem.mem_internal.code_mem[123][6] ;
 wire \mem.mem_internal.code_mem[123][7] ;
 wire \mem.mem_internal.code_mem[124][0] ;
 wire \mem.mem_internal.code_mem[124][1] ;
 wire \mem.mem_internal.code_mem[124][2] ;
 wire \mem.mem_internal.code_mem[124][3] ;
 wire \mem.mem_internal.code_mem[124][4] ;
 wire \mem.mem_internal.code_mem[124][5] ;
 wire \mem.mem_internal.code_mem[124][6] ;
 wire \mem.mem_internal.code_mem[124][7] ;
 wire \mem.mem_internal.code_mem[125][0] ;
 wire \mem.mem_internal.code_mem[125][1] ;
 wire \mem.mem_internal.code_mem[125][2] ;
 wire \mem.mem_internal.code_mem[125][3] ;
 wire \mem.mem_internal.code_mem[125][4] ;
 wire \mem.mem_internal.code_mem[125][5] ;
 wire \mem.mem_internal.code_mem[125][6] ;
 wire \mem.mem_internal.code_mem[125][7] ;
 wire \mem.mem_internal.code_mem[126][0] ;
 wire \mem.mem_internal.code_mem[126][1] ;
 wire \mem.mem_internal.code_mem[126][2] ;
 wire \mem.mem_internal.code_mem[126][3] ;
 wire \mem.mem_internal.code_mem[126][4] ;
 wire \mem.mem_internal.code_mem[126][5] ;
 wire \mem.mem_internal.code_mem[126][6] ;
 wire \mem.mem_internal.code_mem[126][7] ;
 wire \mem.mem_internal.code_mem[127][0] ;
 wire \mem.mem_internal.code_mem[127][1] ;
 wire \mem.mem_internal.code_mem[127][2] ;
 wire \mem.mem_internal.code_mem[127][3] ;
 wire \mem.mem_internal.code_mem[127][4] ;
 wire \mem.mem_internal.code_mem[127][5] ;
 wire \mem.mem_internal.code_mem[127][6] ;
 wire \mem.mem_internal.code_mem[127][7] ;
 wire \mem.mem_internal.code_mem[128][0] ;
 wire \mem.mem_internal.code_mem[128][1] ;
 wire \mem.mem_internal.code_mem[128][2] ;
 wire \mem.mem_internal.code_mem[128][3] ;
 wire \mem.mem_internal.code_mem[128][4] ;
 wire \mem.mem_internal.code_mem[128][5] ;
 wire \mem.mem_internal.code_mem[128][6] ;
 wire \mem.mem_internal.code_mem[128][7] ;
 wire \mem.mem_internal.code_mem[129][0] ;
 wire \mem.mem_internal.code_mem[129][1] ;
 wire \mem.mem_internal.code_mem[129][2] ;
 wire \mem.mem_internal.code_mem[129][3] ;
 wire \mem.mem_internal.code_mem[129][4] ;
 wire \mem.mem_internal.code_mem[129][5] ;
 wire \mem.mem_internal.code_mem[129][6] ;
 wire \mem.mem_internal.code_mem[129][7] ;
 wire \mem.mem_internal.code_mem[12][0] ;
 wire \mem.mem_internal.code_mem[12][1] ;
 wire \mem.mem_internal.code_mem[12][2] ;
 wire \mem.mem_internal.code_mem[12][3] ;
 wire \mem.mem_internal.code_mem[12][4] ;
 wire \mem.mem_internal.code_mem[12][5] ;
 wire \mem.mem_internal.code_mem[12][6] ;
 wire \mem.mem_internal.code_mem[12][7] ;
 wire \mem.mem_internal.code_mem[130][0] ;
 wire \mem.mem_internal.code_mem[130][1] ;
 wire \mem.mem_internal.code_mem[130][2] ;
 wire \mem.mem_internal.code_mem[130][3] ;
 wire \mem.mem_internal.code_mem[130][4] ;
 wire \mem.mem_internal.code_mem[130][5] ;
 wire \mem.mem_internal.code_mem[130][6] ;
 wire \mem.mem_internal.code_mem[130][7] ;
 wire \mem.mem_internal.code_mem[131][0] ;
 wire \mem.mem_internal.code_mem[131][1] ;
 wire \mem.mem_internal.code_mem[131][2] ;
 wire \mem.mem_internal.code_mem[131][3] ;
 wire \mem.mem_internal.code_mem[131][4] ;
 wire \mem.mem_internal.code_mem[131][5] ;
 wire \mem.mem_internal.code_mem[131][6] ;
 wire \mem.mem_internal.code_mem[131][7] ;
 wire \mem.mem_internal.code_mem[132][0] ;
 wire \mem.mem_internal.code_mem[132][1] ;
 wire \mem.mem_internal.code_mem[132][2] ;
 wire \mem.mem_internal.code_mem[132][3] ;
 wire \mem.mem_internal.code_mem[132][4] ;
 wire \mem.mem_internal.code_mem[132][5] ;
 wire \mem.mem_internal.code_mem[132][6] ;
 wire \mem.mem_internal.code_mem[132][7] ;
 wire \mem.mem_internal.code_mem[133][0] ;
 wire \mem.mem_internal.code_mem[133][1] ;
 wire \mem.mem_internal.code_mem[133][2] ;
 wire \mem.mem_internal.code_mem[133][3] ;
 wire \mem.mem_internal.code_mem[133][4] ;
 wire \mem.mem_internal.code_mem[133][5] ;
 wire \mem.mem_internal.code_mem[133][6] ;
 wire \mem.mem_internal.code_mem[133][7] ;
 wire \mem.mem_internal.code_mem[134][0] ;
 wire \mem.mem_internal.code_mem[134][1] ;
 wire \mem.mem_internal.code_mem[134][2] ;
 wire \mem.mem_internal.code_mem[134][3] ;
 wire \mem.mem_internal.code_mem[134][4] ;
 wire \mem.mem_internal.code_mem[134][5] ;
 wire \mem.mem_internal.code_mem[134][6] ;
 wire \mem.mem_internal.code_mem[134][7] ;
 wire \mem.mem_internal.code_mem[135][0] ;
 wire \mem.mem_internal.code_mem[135][1] ;
 wire \mem.mem_internal.code_mem[135][2] ;
 wire \mem.mem_internal.code_mem[135][3] ;
 wire \mem.mem_internal.code_mem[135][4] ;
 wire \mem.mem_internal.code_mem[135][5] ;
 wire \mem.mem_internal.code_mem[135][6] ;
 wire \mem.mem_internal.code_mem[135][7] ;
 wire \mem.mem_internal.code_mem[136][0] ;
 wire \mem.mem_internal.code_mem[136][1] ;
 wire \mem.mem_internal.code_mem[136][2] ;
 wire \mem.mem_internal.code_mem[136][3] ;
 wire \mem.mem_internal.code_mem[136][4] ;
 wire \mem.mem_internal.code_mem[136][5] ;
 wire \mem.mem_internal.code_mem[136][6] ;
 wire \mem.mem_internal.code_mem[136][7] ;
 wire \mem.mem_internal.code_mem[137][0] ;
 wire \mem.mem_internal.code_mem[137][1] ;
 wire \mem.mem_internal.code_mem[137][2] ;
 wire \mem.mem_internal.code_mem[137][3] ;
 wire \mem.mem_internal.code_mem[137][4] ;
 wire \mem.mem_internal.code_mem[137][5] ;
 wire \mem.mem_internal.code_mem[137][6] ;
 wire \mem.mem_internal.code_mem[137][7] ;
 wire \mem.mem_internal.code_mem[138][0] ;
 wire \mem.mem_internal.code_mem[138][1] ;
 wire \mem.mem_internal.code_mem[138][2] ;
 wire \mem.mem_internal.code_mem[138][3] ;
 wire \mem.mem_internal.code_mem[138][4] ;
 wire \mem.mem_internal.code_mem[138][5] ;
 wire \mem.mem_internal.code_mem[138][6] ;
 wire \mem.mem_internal.code_mem[138][7] ;
 wire \mem.mem_internal.code_mem[139][0] ;
 wire \mem.mem_internal.code_mem[139][1] ;
 wire \mem.mem_internal.code_mem[139][2] ;
 wire \mem.mem_internal.code_mem[139][3] ;
 wire \mem.mem_internal.code_mem[139][4] ;
 wire \mem.mem_internal.code_mem[139][5] ;
 wire \mem.mem_internal.code_mem[139][6] ;
 wire \mem.mem_internal.code_mem[139][7] ;
 wire \mem.mem_internal.code_mem[13][0] ;
 wire \mem.mem_internal.code_mem[13][1] ;
 wire \mem.mem_internal.code_mem[13][2] ;
 wire \mem.mem_internal.code_mem[13][3] ;
 wire \mem.mem_internal.code_mem[13][4] ;
 wire \mem.mem_internal.code_mem[13][5] ;
 wire \mem.mem_internal.code_mem[13][6] ;
 wire \mem.mem_internal.code_mem[13][7] ;
 wire \mem.mem_internal.code_mem[140][0] ;
 wire \mem.mem_internal.code_mem[140][1] ;
 wire \mem.mem_internal.code_mem[140][2] ;
 wire \mem.mem_internal.code_mem[140][3] ;
 wire \mem.mem_internal.code_mem[140][4] ;
 wire \mem.mem_internal.code_mem[140][5] ;
 wire \mem.mem_internal.code_mem[140][6] ;
 wire \mem.mem_internal.code_mem[140][7] ;
 wire \mem.mem_internal.code_mem[141][0] ;
 wire \mem.mem_internal.code_mem[141][1] ;
 wire \mem.mem_internal.code_mem[141][2] ;
 wire \mem.mem_internal.code_mem[141][3] ;
 wire \mem.mem_internal.code_mem[141][4] ;
 wire \mem.mem_internal.code_mem[141][5] ;
 wire \mem.mem_internal.code_mem[141][6] ;
 wire \mem.mem_internal.code_mem[141][7] ;
 wire \mem.mem_internal.code_mem[142][0] ;
 wire \mem.mem_internal.code_mem[142][1] ;
 wire \mem.mem_internal.code_mem[142][2] ;
 wire \mem.mem_internal.code_mem[142][3] ;
 wire \mem.mem_internal.code_mem[142][4] ;
 wire \mem.mem_internal.code_mem[142][5] ;
 wire \mem.mem_internal.code_mem[142][6] ;
 wire \mem.mem_internal.code_mem[142][7] ;
 wire \mem.mem_internal.code_mem[143][0] ;
 wire \mem.mem_internal.code_mem[143][1] ;
 wire \mem.mem_internal.code_mem[143][2] ;
 wire \mem.mem_internal.code_mem[143][3] ;
 wire \mem.mem_internal.code_mem[143][4] ;
 wire \mem.mem_internal.code_mem[143][5] ;
 wire \mem.mem_internal.code_mem[143][6] ;
 wire \mem.mem_internal.code_mem[143][7] ;
 wire \mem.mem_internal.code_mem[144][0] ;
 wire \mem.mem_internal.code_mem[144][1] ;
 wire \mem.mem_internal.code_mem[144][2] ;
 wire \mem.mem_internal.code_mem[144][3] ;
 wire \mem.mem_internal.code_mem[144][4] ;
 wire \mem.mem_internal.code_mem[144][5] ;
 wire \mem.mem_internal.code_mem[144][6] ;
 wire \mem.mem_internal.code_mem[144][7] ;
 wire \mem.mem_internal.code_mem[145][0] ;
 wire \mem.mem_internal.code_mem[145][1] ;
 wire \mem.mem_internal.code_mem[145][2] ;
 wire \mem.mem_internal.code_mem[145][3] ;
 wire \mem.mem_internal.code_mem[145][4] ;
 wire \mem.mem_internal.code_mem[145][5] ;
 wire \mem.mem_internal.code_mem[145][6] ;
 wire \mem.mem_internal.code_mem[145][7] ;
 wire \mem.mem_internal.code_mem[146][0] ;
 wire \mem.mem_internal.code_mem[146][1] ;
 wire \mem.mem_internal.code_mem[146][2] ;
 wire \mem.mem_internal.code_mem[146][3] ;
 wire \mem.mem_internal.code_mem[146][4] ;
 wire \mem.mem_internal.code_mem[146][5] ;
 wire \mem.mem_internal.code_mem[146][6] ;
 wire \mem.mem_internal.code_mem[146][7] ;
 wire \mem.mem_internal.code_mem[147][0] ;
 wire \mem.mem_internal.code_mem[147][1] ;
 wire \mem.mem_internal.code_mem[147][2] ;
 wire \mem.mem_internal.code_mem[147][3] ;
 wire \mem.mem_internal.code_mem[147][4] ;
 wire \mem.mem_internal.code_mem[147][5] ;
 wire \mem.mem_internal.code_mem[147][6] ;
 wire \mem.mem_internal.code_mem[147][7] ;
 wire \mem.mem_internal.code_mem[148][0] ;
 wire \mem.mem_internal.code_mem[148][1] ;
 wire \mem.mem_internal.code_mem[148][2] ;
 wire \mem.mem_internal.code_mem[148][3] ;
 wire \mem.mem_internal.code_mem[148][4] ;
 wire \mem.mem_internal.code_mem[148][5] ;
 wire \mem.mem_internal.code_mem[148][6] ;
 wire \mem.mem_internal.code_mem[148][7] ;
 wire \mem.mem_internal.code_mem[149][0] ;
 wire \mem.mem_internal.code_mem[149][1] ;
 wire \mem.mem_internal.code_mem[149][2] ;
 wire \mem.mem_internal.code_mem[149][3] ;
 wire \mem.mem_internal.code_mem[149][4] ;
 wire \mem.mem_internal.code_mem[149][5] ;
 wire \mem.mem_internal.code_mem[149][6] ;
 wire \mem.mem_internal.code_mem[149][7] ;
 wire \mem.mem_internal.code_mem[14][0] ;
 wire \mem.mem_internal.code_mem[14][1] ;
 wire \mem.mem_internal.code_mem[14][2] ;
 wire \mem.mem_internal.code_mem[14][3] ;
 wire \mem.mem_internal.code_mem[14][4] ;
 wire \mem.mem_internal.code_mem[14][5] ;
 wire \mem.mem_internal.code_mem[14][6] ;
 wire \mem.mem_internal.code_mem[14][7] ;
 wire \mem.mem_internal.code_mem[150][0] ;
 wire \mem.mem_internal.code_mem[150][1] ;
 wire \mem.mem_internal.code_mem[150][2] ;
 wire \mem.mem_internal.code_mem[150][3] ;
 wire \mem.mem_internal.code_mem[150][4] ;
 wire \mem.mem_internal.code_mem[150][5] ;
 wire \mem.mem_internal.code_mem[150][6] ;
 wire \mem.mem_internal.code_mem[150][7] ;
 wire \mem.mem_internal.code_mem[151][0] ;
 wire \mem.mem_internal.code_mem[151][1] ;
 wire \mem.mem_internal.code_mem[151][2] ;
 wire \mem.mem_internal.code_mem[151][3] ;
 wire \mem.mem_internal.code_mem[151][4] ;
 wire \mem.mem_internal.code_mem[151][5] ;
 wire \mem.mem_internal.code_mem[151][6] ;
 wire \mem.mem_internal.code_mem[151][7] ;
 wire \mem.mem_internal.code_mem[152][0] ;
 wire \mem.mem_internal.code_mem[152][1] ;
 wire \mem.mem_internal.code_mem[152][2] ;
 wire \mem.mem_internal.code_mem[152][3] ;
 wire \mem.mem_internal.code_mem[152][4] ;
 wire \mem.mem_internal.code_mem[152][5] ;
 wire \mem.mem_internal.code_mem[152][6] ;
 wire \mem.mem_internal.code_mem[152][7] ;
 wire \mem.mem_internal.code_mem[153][0] ;
 wire \mem.mem_internal.code_mem[153][1] ;
 wire \mem.mem_internal.code_mem[153][2] ;
 wire \mem.mem_internal.code_mem[153][3] ;
 wire \mem.mem_internal.code_mem[153][4] ;
 wire \mem.mem_internal.code_mem[153][5] ;
 wire \mem.mem_internal.code_mem[153][6] ;
 wire \mem.mem_internal.code_mem[153][7] ;
 wire \mem.mem_internal.code_mem[154][0] ;
 wire \mem.mem_internal.code_mem[154][1] ;
 wire \mem.mem_internal.code_mem[154][2] ;
 wire \mem.mem_internal.code_mem[154][3] ;
 wire \mem.mem_internal.code_mem[154][4] ;
 wire \mem.mem_internal.code_mem[154][5] ;
 wire \mem.mem_internal.code_mem[154][6] ;
 wire \mem.mem_internal.code_mem[154][7] ;
 wire \mem.mem_internal.code_mem[155][0] ;
 wire \mem.mem_internal.code_mem[155][1] ;
 wire \mem.mem_internal.code_mem[155][2] ;
 wire \mem.mem_internal.code_mem[155][3] ;
 wire \mem.mem_internal.code_mem[155][4] ;
 wire \mem.mem_internal.code_mem[155][5] ;
 wire \mem.mem_internal.code_mem[155][6] ;
 wire \mem.mem_internal.code_mem[155][7] ;
 wire \mem.mem_internal.code_mem[156][0] ;
 wire \mem.mem_internal.code_mem[156][1] ;
 wire \mem.mem_internal.code_mem[156][2] ;
 wire \mem.mem_internal.code_mem[156][3] ;
 wire \mem.mem_internal.code_mem[156][4] ;
 wire \mem.mem_internal.code_mem[156][5] ;
 wire \mem.mem_internal.code_mem[156][6] ;
 wire \mem.mem_internal.code_mem[156][7] ;
 wire \mem.mem_internal.code_mem[157][0] ;
 wire \mem.mem_internal.code_mem[157][1] ;
 wire \mem.mem_internal.code_mem[157][2] ;
 wire \mem.mem_internal.code_mem[157][3] ;
 wire \mem.mem_internal.code_mem[157][4] ;
 wire \mem.mem_internal.code_mem[157][5] ;
 wire \mem.mem_internal.code_mem[157][6] ;
 wire \mem.mem_internal.code_mem[157][7] ;
 wire \mem.mem_internal.code_mem[158][0] ;
 wire \mem.mem_internal.code_mem[158][1] ;
 wire \mem.mem_internal.code_mem[158][2] ;
 wire \mem.mem_internal.code_mem[158][3] ;
 wire \mem.mem_internal.code_mem[158][4] ;
 wire \mem.mem_internal.code_mem[158][5] ;
 wire \mem.mem_internal.code_mem[158][6] ;
 wire \mem.mem_internal.code_mem[158][7] ;
 wire \mem.mem_internal.code_mem[159][0] ;
 wire \mem.mem_internal.code_mem[159][1] ;
 wire \mem.mem_internal.code_mem[159][2] ;
 wire \mem.mem_internal.code_mem[159][3] ;
 wire \mem.mem_internal.code_mem[159][4] ;
 wire \mem.mem_internal.code_mem[159][5] ;
 wire \mem.mem_internal.code_mem[159][6] ;
 wire \mem.mem_internal.code_mem[159][7] ;
 wire \mem.mem_internal.code_mem[15][0] ;
 wire \mem.mem_internal.code_mem[15][1] ;
 wire \mem.mem_internal.code_mem[15][2] ;
 wire \mem.mem_internal.code_mem[15][3] ;
 wire \mem.mem_internal.code_mem[15][4] ;
 wire \mem.mem_internal.code_mem[15][5] ;
 wire \mem.mem_internal.code_mem[15][6] ;
 wire \mem.mem_internal.code_mem[15][7] ;
 wire \mem.mem_internal.code_mem[160][0] ;
 wire \mem.mem_internal.code_mem[160][1] ;
 wire \mem.mem_internal.code_mem[160][2] ;
 wire \mem.mem_internal.code_mem[160][3] ;
 wire \mem.mem_internal.code_mem[160][4] ;
 wire \mem.mem_internal.code_mem[160][5] ;
 wire \mem.mem_internal.code_mem[160][6] ;
 wire \mem.mem_internal.code_mem[160][7] ;
 wire \mem.mem_internal.code_mem[161][0] ;
 wire \mem.mem_internal.code_mem[161][1] ;
 wire \mem.mem_internal.code_mem[161][2] ;
 wire \mem.mem_internal.code_mem[161][3] ;
 wire \mem.mem_internal.code_mem[161][4] ;
 wire \mem.mem_internal.code_mem[161][5] ;
 wire \mem.mem_internal.code_mem[161][6] ;
 wire \mem.mem_internal.code_mem[161][7] ;
 wire \mem.mem_internal.code_mem[162][0] ;
 wire \mem.mem_internal.code_mem[162][1] ;
 wire \mem.mem_internal.code_mem[162][2] ;
 wire \mem.mem_internal.code_mem[162][3] ;
 wire \mem.mem_internal.code_mem[162][4] ;
 wire \mem.mem_internal.code_mem[162][5] ;
 wire \mem.mem_internal.code_mem[162][6] ;
 wire \mem.mem_internal.code_mem[162][7] ;
 wire \mem.mem_internal.code_mem[163][0] ;
 wire \mem.mem_internal.code_mem[163][1] ;
 wire \mem.mem_internal.code_mem[163][2] ;
 wire \mem.mem_internal.code_mem[163][3] ;
 wire \mem.mem_internal.code_mem[163][4] ;
 wire \mem.mem_internal.code_mem[163][5] ;
 wire \mem.mem_internal.code_mem[163][6] ;
 wire \mem.mem_internal.code_mem[163][7] ;
 wire \mem.mem_internal.code_mem[164][0] ;
 wire \mem.mem_internal.code_mem[164][1] ;
 wire \mem.mem_internal.code_mem[164][2] ;
 wire \mem.mem_internal.code_mem[164][3] ;
 wire \mem.mem_internal.code_mem[164][4] ;
 wire \mem.mem_internal.code_mem[164][5] ;
 wire \mem.mem_internal.code_mem[164][6] ;
 wire \mem.mem_internal.code_mem[164][7] ;
 wire \mem.mem_internal.code_mem[165][0] ;
 wire \mem.mem_internal.code_mem[165][1] ;
 wire \mem.mem_internal.code_mem[165][2] ;
 wire \mem.mem_internal.code_mem[165][3] ;
 wire \mem.mem_internal.code_mem[165][4] ;
 wire \mem.mem_internal.code_mem[165][5] ;
 wire \mem.mem_internal.code_mem[165][6] ;
 wire \mem.mem_internal.code_mem[165][7] ;
 wire \mem.mem_internal.code_mem[166][0] ;
 wire \mem.mem_internal.code_mem[166][1] ;
 wire \mem.mem_internal.code_mem[166][2] ;
 wire \mem.mem_internal.code_mem[166][3] ;
 wire \mem.mem_internal.code_mem[166][4] ;
 wire \mem.mem_internal.code_mem[166][5] ;
 wire \mem.mem_internal.code_mem[166][6] ;
 wire \mem.mem_internal.code_mem[166][7] ;
 wire \mem.mem_internal.code_mem[167][0] ;
 wire \mem.mem_internal.code_mem[167][1] ;
 wire \mem.mem_internal.code_mem[167][2] ;
 wire \mem.mem_internal.code_mem[167][3] ;
 wire \mem.mem_internal.code_mem[167][4] ;
 wire \mem.mem_internal.code_mem[167][5] ;
 wire \mem.mem_internal.code_mem[167][6] ;
 wire \mem.mem_internal.code_mem[167][7] ;
 wire \mem.mem_internal.code_mem[168][0] ;
 wire \mem.mem_internal.code_mem[168][1] ;
 wire \mem.mem_internal.code_mem[168][2] ;
 wire \mem.mem_internal.code_mem[168][3] ;
 wire \mem.mem_internal.code_mem[168][4] ;
 wire \mem.mem_internal.code_mem[168][5] ;
 wire \mem.mem_internal.code_mem[168][6] ;
 wire \mem.mem_internal.code_mem[168][7] ;
 wire \mem.mem_internal.code_mem[169][0] ;
 wire \mem.mem_internal.code_mem[169][1] ;
 wire \mem.mem_internal.code_mem[169][2] ;
 wire \mem.mem_internal.code_mem[169][3] ;
 wire \mem.mem_internal.code_mem[169][4] ;
 wire \mem.mem_internal.code_mem[169][5] ;
 wire \mem.mem_internal.code_mem[169][6] ;
 wire \mem.mem_internal.code_mem[169][7] ;
 wire \mem.mem_internal.code_mem[16][0] ;
 wire \mem.mem_internal.code_mem[16][1] ;
 wire \mem.mem_internal.code_mem[16][2] ;
 wire \mem.mem_internal.code_mem[16][3] ;
 wire \mem.mem_internal.code_mem[16][4] ;
 wire \mem.mem_internal.code_mem[16][5] ;
 wire \mem.mem_internal.code_mem[16][6] ;
 wire \mem.mem_internal.code_mem[16][7] ;
 wire \mem.mem_internal.code_mem[170][0] ;
 wire \mem.mem_internal.code_mem[170][1] ;
 wire \mem.mem_internal.code_mem[170][2] ;
 wire \mem.mem_internal.code_mem[170][3] ;
 wire \mem.mem_internal.code_mem[170][4] ;
 wire \mem.mem_internal.code_mem[170][5] ;
 wire \mem.mem_internal.code_mem[170][6] ;
 wire \mem.mem_internal.code_mem[170][7] ;
 wire \mem.mem_internal.code_mem[171][0] ;
 wire \mem.mem_internal.code_mem[171][1] ;
 wire \mem.mem_internal.code_mem[171][2] ;
 wire \mem.mem_internal.code_mem[171][3] ;
 wire \mem.mem_internal.code_mem[171][4] ;
 wire \mem.mem_internal.code_mem[171][5] ;
 wire \mem.mem_internal.code_mem[171][6] ;
 wire \mem.mem_internal.code_mem[171][7] ;
 wire \mem.mem_internal.code_mem[172][0] ;
 wire \mem.mem_internal.code_mem[172][1] ;
 wire \mem.mem_internal.code_mem[172][2] ;
 wire \mem.mem_internal.code_mem[172][3] ;
 wire \mem.mem_internal.code_mem[172][4] ;
 wire \mem.mem_internal.code_mem[172][5] ;
 wire \mem.mem_internal.code_mem[172][6] ;
 wire \mem.mem_internal.code_mem[172][7] ;
 wire \mem.mem_internal.code_mem[173][0] ;
 wire \mem.mem_internal.code_mem[173][1] ;
 wire \mem.mem_internal.code_mem[173][2] ;
 wire \mem.mem_internal.code_mem[173][3] ;
 wire \mem.mem_internal.code_mem[173][4] ;
 wire \mem.mem_internal.code_mem[173][5] ;
 wire \mem.mem_internal.code_mem[173][6] ;
 wire \mem.mem_internal.code_mem[173][7] ;
 wire \mem.mem_internal.code_mem[174][0] ;
 wire \mem.mem_internal.code_mem[174][1] ;
 wire \mem.mem_internal.code_mem[174][2] ;
 wire \mem.mem_internal.code_mem[174][3] ;
 wire \mem.mem_internal.code_mem[174][4] ;
 wire \mem.mem_internal.code_mem[174][5] ;
 wire \mem.mem_internal.code_mem[174][6] ;
 wire \mem.mem_internal.code_mem[174][7] ;
 wire \mem.mem_internal.code_mem[175][0] ;
 wire \mem.mem_internal.code_mem[175][1] ;
 wire \mem.mem_internal.code_mem[175][2] ;
 wire \mem.mem_internal.code_mem[175][3] ;
 wire \mem.mem_internal.code_mem[175][4] ;
 wire \mem.mem_internal.code_mem[175][5] ;
 wire \mem.mem_internal.code_mem[175][6] ;
 wire \mem.mem_internal.code_mem[175][7] ;
 wire \mem.mem_internal.code_mem[176][0] ;
 wire \mem.mem_internal.code_mem[176][1] ;
 wire \mem.mem_internal.code_mem[176][2] ;
 wire \mem.mem_internal.code_mem[176][3] ;
 wire \mem.mem_internal.code_mem[176][4] ;
 wire \mem.mem_internal.code_mem[176][5] ;
 wire \mem.mem_internal.code_mem[176][6] ;
 wire \mem.mem_internal.code_mem[176][7] ;
 wire \mem.mem_internal.code_mem[177][0] ;
 wire \mem.mem_internal.code_mem[177][1] ;
 wire \mem.mem_internal.code_mem[177][2] ;
 wire \mem.mem_internal.code_mem[177][3] ;
 wire \mem.mem_internal.code_mem[177][4] ;
 wire \mem.mem_internal.code_mem[177][5] ;
 wire \mem.mem_internal.code_mem[177][6] ;
 wire \mem.mem_internal.code_mem[177][7] ;
 wire \mem.mem_internal.code_mem[178][0] ;
 wire \mem.mem_internal.code_mem[178][1] ;
 wire \mem.mem_internal.code_mem[178][2] ;
 wire \mem.mem_internal.code_mem[178][3] ;
 wire \mem.mem_internal.code_mem[178][4] ;
 wire \mem.mem_internal.code_mem[178][5] ;
 wire \mem.mem_internal.code_mem[178][6] ;
 wire \mem.mem_internal.code_mem[178][7] ;
 wire \mem.mem_internal.code_mem[179][0] ;
 wire \mem.mem_internal.code_mem[179][1] ;
 wire \mem.mem_internal.code_mem[179][2] ;
 wire \mem.mem_internal.code_mem[179][3] ;
 wire \mem.mem_internal.code_mem[179][4] ;
 wire \mem.mem_internal.code_mem[179][5] ;
 wire \mem.mem_internal.code_mem[179][6] ;
 wire \mem.mem_internal.code_mem[179][7] ;
 wire \mem.mem_internal.code_mem[17][0] ;
 wire \mem.mem_internal.code_mem[17][1] ;
 wire \mem.mem_internal.code_mem[17][2] ;
 wire \mem.mem_internal.code_mem[17][3] ;
 wire \mem.mem_internal.code_mem[17][4] ;
 wire \mem.mem_internal.code_mem[17][5] ;
 wire \mem.mem_internal.code_mem[17][6] ;
 wire \mem.mem_internal.code_mem[17][7] ;
 wire \mem.mem_internal.code_mem[180][0] ;
 wire \mem.mem_internal.code_mem[180][1] ;
 wire \mem.mem_internal.code_mem[180][2] ;
 wire \mem.mem_internal.code_mem[180][3] ;
 wire \mem.mem_internal.code_mem[180][4] ;
 wire \mem.mem_internal.code_mem[180][5] ;
 wire \mem.mem_internal.code_mem[180][6] ;
 wire \mem.mem_internal.code_mem[180][7] ;
 wire \mem.mem_internal.code_mem[181][0] ;
 wire \mem.mem_internal.code_mem[181][1] ;
 wire \mem.mem_internal.code_mem[181][2] ;
 wire \mem.mem_internal.code_mem[181][3] ;
 wire \mem.mem_internal.code_mem[181][4] ;
 wire \mem.mem_internal.code_mem[181][5] ;
 wire \mem.mem_internal.code_mem[181][6] ;
 wire \mem.mem_internal.code_mem[181][7] ;
 wire \mem.mem_internal.code_mem[182][0] ;
 wire \mem.mem_internal.code_mem[182][1] ;
 wire \mem.mem_internal.code_mem[182][2] ;
 wire \mem.mem_internal.code_mem[182][3] ;
 wire \mem.mem_internal.code_mem[182][4] ;
 wire \mem.mem_internal.code_mem[182][5] ;
 wire \mem.mem_internal.code_mem[182][6] ;
 wire \mem.mem_internal.code_mem[182][7] ;
 wire \mem.mem_internal.code_mem[183][0] ;
 wire \mem.mem_internal.code_mem[183][1] ;
 wire \mem.mem_internal.code_mem[183][2] ;
 wire \mem.mem_internal.code_mem[183][3] ;
 wire \mem.mem_internal.code_mem[183][4] ;
 wire \mem.mem_internal.code_mem[183][5] ;
 wire \mem.mem_internal.code_mem[183][6] ;
 wire \mem.mem_internal.code_mem[183][7] ;
 wire \mem.mem_internal.code_mem[184][0] ;
 wire \mem.mem_internal.code_mem[184][1] ;
 wire \mem.mem_internal.code_mem[184][2] ;
 wire \mem.mem_internal.code_mem[184][3] ;
 wire \mem.mem_internal.code_mem[184][4] ;
 wire \mem.mem_internal.code_mem[184][5] ;
 wire \mem.mem_internal.code_mem[184][6] ;
 wire \mem.mem_internal.code_mem[184][7] ;
 wire \mem.mem_internal.code_mem[185][0] ;
 wire \mem.mem_internal.code_mem[185][1] ;
 wire \mem.mem_internal.code_mem[185][2] ;
 wire \mem.mem_internal.code_mem[185][3] ;
 wire \mem.mem_internal.code_mem[185][4] ;
 wire \mem.mem_internal.code_mem[185][5] ;
 wire \mem.mem_internal.code_mem[185][6] ;
 wire \mem.mem_internal.code_mem[185][7] ;
 wire \mem.mem_internal.code_mem[186][0] ;
 wire \mem.mem_internal.code_mem[186][1] ;
 wire \mem.mem_internal.code_mem[186][2] ;
 wire \mem.mem_internal.code_mem[186][3] ;
 wire \mem.mem_internal.code_mem[186][4] ;
 wire \mem.mem_internal.code_mem[186][5] ;
 wire \mem.mem_internal.code_mem[186][6] ;
 wire \mem.mem_internal.code_mem[186][7] ;
 wire \mem.mem_internal.code_mem[187][0] ;
 wire \mem.mem_internal.code_mem[187][1] ;
 wire \mem.mem_internal.code_mem[187][2] ;
 wire \mem.mem_internal.code_mem[187][3] ;
 wire \mem.mem_internal.code_mem[187][4] ;
 wire \mem.mem_internal.code_mem[187][5] ;
 wire \mem.mem_internal.code_mem[187][6] ;
 wire \mem.mem_internal.code_mem[187][7] ;
 wire \mem.mem_internal.code_mem[188][0] ;
 wire \mem.mem_internal.code_mem[188][1] ;
 wire \mem.mem_internal.code_mem[188][2] ;
 wire \mem.mem_internal.code_mem[188][3] ;
 wire \mem.mem_internal.code_mem[188][4] ;
 wire \mem.mem_internal.code_mem[188][5] ;
 wire \mem.mem_internal.code_mem[188][6] ;
 wire \mem.mem_internal.code_mem[188][7] ;
 wire \mem.mem_internal.code_mem[189][0] ;
 wire \mem.mem_internal.code_mem[189][1] ;
 wire \mem.mem_internal.code_mem[189][2] ;
 wire \mem.mem_internal.code_mem[189][3] ;
 wire \mem.mem_internal.code_mem[189][4] ;
 wire \mem.mem_internal.code_mem[189][5] ;
 wire \mem.mem_internal.code_mem[189][6] ;
 wire \mem.mem_internal.code_mem[189][7] ;
 wire \mem.mem_internal.code_mem[18][0] ;
 wire \mem.mem_internal.code_mem[18][1] ;
 wire \mem.mem_internal.code_mem[18][2] ;
 wire \mem.mem_internal.code_mem[18][3] ;
 wire \mem.mem_internal.code_mem[18][4] ;
 wire \mem.mem_internal.code_mem[18][5] ;
 wire \mem.mem_internal.code_mem[18][6] ;
 wire \mem.mem_internal.code_mem[18][7] ;
 wire \mem.mem_internal.code_mem[190][0] ;
 wire \mem.mem_internal.code_mem[190][1] ;
 wire \mem.mem_internal.code_mem[190][2] ;
 wire \mem.mem_internal.code_mem[190][3] ;
 wire \mem.mem_internal.code_mem[190][4] ;
 wire \mem.mem_internal.code_mem[190][5] ;
 wire \mem.mem_internal.code_mem[190][6] ;
 wire \mem.mem_internal.code_mem[190][7] ;
 wire \mem.mem_internal.code_mem[191][0] ;
 wire \mem.mem_internal.code_mem[191][1] ;
 wire \mem.mem_internal.code_mem[191][2] ;
 wire \mem.mem_internal.code_mem[191][3] ;
 wire \mem.mem_internal.code_mem[191][4] ;
 wire \mem.mem_internal.code_mem[191][5] ;
 wire \mem.mem_internal.code_mem[191][6] ;
 wire \mem.mem_internal.code_mem[191][7] ;
 wire \mem.mem_internal.code_mem[192][0] ;
 wire \mem.mem_internal.code_mem[192][1] ;
 wire \mem.mem_internal.code_mem[192][2] ;
 wire \mem.mem_internal.code_mem[192][3] ;
 wire \mem.mem_internal.code_mem[192][4] ;
 wire \mem.mem_internal.code_mem[192][5] ;
 wire \mem.mem_internal.code_mem[192][6] ;
 wire \mem.mem_internal.code_mem[192][7] ;
 wire \mem.mem_internal.code_mem[193][0] ;
 wire \mem.mem_internal.code_mem[193][1] ;
 wire \mem.mem_internal.code_mem[193][2] ;
 wire \mem.mem_internal.code_mem[193][3] ;
 wire \mem.mem_internal.code_mem[193][4] ;
 wire \mem.mem_internal.code_mem[193][5] ;
 wire \mem.mem_internal.code_mem[193][6] ;
 wire \mem.mem_internal.code_mem[193][7] ;
 wire \mem.mem_internal.code_mem[194][0] ;
 wire \mem.mem_internal.code_mem[194][1] ;
 wire \mem.mem_internal.code_mem[194][2] ;
 wire \mem.mem_internal.code_mem[194][3] ;
 wire \mem.mem_internal.code_mem[194][4] ;
 wire \mem.mem_internal.code_mem[194][5] ;
 wire \mem.mem_internal.code_mem[194][6] ;
 wire \mem.mem_internal.code_mem[194][7] ;
 wire \mem.mem_internal.code_mem[195][0] ;
 wire \mem.mem_internal.code_mem[195][1] ;
 wire \mem.mem_internal.code_mem[195][2] ;
 wire \mem.mem_internal.code_mem[195][3] ;
 wire \mem.mem_internal.code_mem[195][4] ;
 wire \mem.mem_internal.code_mem[195][5] ;
 wire \mem.mem_internal.code_mem[195][6] ;
 wire \mem.mem_internal.code_mem[195][7] ;
 wire \mem.mem_internal.code_mem[196][0] ;
 wire \mem.mem_internal.code_mem[196][1] ;
 wire \mem.mem_internal.code_mem[196][2] ;
 wire \mem.mem_internal.code_mem[196][3] ;
 wire \mem.mem_internal.code_mem[196][4] ;
 wire \mem.mem_internal.code_mem[196][5] ;
 wire \mem.mem_internal.code_mem[196][6] ;
 wire \mem.mem_internal.code_mem[196][7] ;
 wire \mem.mem_internal.code_mem[197][0] ;
 wire \mem.mem_internal.code_mem[197][1] ;
 wire \mem.mem_internal.code_mem[197][2] ;
 wire \mem.mem_internal.code_mem[197][3] ;
 wire \mem.mem_internal.code_mem[197][4] ;
 wire \mem.mem_internal.code_mem[197][5] ;
 wire \mem.mem_internal.code_mem[197][6] ;
 wire \mem.mem_internal.code_mem[197][7] ;
 wire \mem.mem_internal.code_mem[198][0] ;
 wire \mem.mem_internal.code_mem[198][1] ;
 wire \mem.mem_internal.code_mem[198][2] ;
 wire \mem.mem_internal.code_mem[198][3] ;
 wire \mem.mem_internal.code_mem[198][4] ;
 wire \mem.mem_internal.code_mem[198][5] ;
 wire \mem.mem_internal.code_mem[198][6] ;
 wire \mem.mem_internal.code_mem[198][7] ;
 wire \mem.mem_internal.code_mem[199][0] ;
 wire \mem.mem_internal.code_mem[199][1] ;
 wire \mem.mem_internal.code_mem[199][2] ;
 wire \mem.mem_internal.code_mem[199][3] ;
 wire \mem.mem_internal.code_mem[199][4] ;
 wire \mem.mem_internal.code_mem[199][5] ;
 wire \mem.mem_internal.code_mem[199][6] ;
 wire \mem.mem_internal.code_mem[199][7] ;
 wire \mem.mem_internal.code_mem[19][0] ;
 wire \mem.mem_internal.code_mem[19][1] ;
 wire \mem.mem_internal.code_mem[19][2] ;
 wire \mem.mem_internal.code_mem[19][3] ;
 wire \mem.mem_internal.code_mem[19][4] ;
 wire \mem.mem_internal.code_mem[19][5] ;
 wire \mem.mem_internal.code_mem[19][6] ;
 wire \mem.mem_internal.code_mem[19][7] ;
 wire \mem.mem_internal.code_mem[1][0] ;
 wire \mem.mem_internal.code_mem[1][1] ;
 wire \mem.mem_internal.code_mem[1][2] ;
 wire \mem.mem_internal.code_mem[1][3] ;
 wire \mem.mem_internal.code_mem[1][4] ;
 wire \mem.mem_internal.code_mem[1][5] ;
 wire \mem.mem_internal.code_mem[1][6] ;
 wire \mem.mem_internal.code_mem[1][7] ;
 wire \mem.mem_internal.code_mem[200][0] ;
 wire \mem.mem_internal.code_mem[200][1] ;
 wire \mem.mem_internal.code_mem[200][2] ;
 wire \mem.mem_internal.code_mem[200][3] ;
 wire \mem.mem_internal.code_mem[200][4] ;
 wire \mem.mem_internal.code_mem[200][5] ;
 wire \mem.mem_internal.code_mem[200][6] ;
 wire \mem.mem_internal.code_mem[200][7] ;
 wire \mem.mem_internal.code_mem[201][0] ;
 wire \mem.mem_internal.code_mem[201][1] ;
 wire \mem.mem_internal.code_mem[201][2] ;
 wire \mem.mem_internal.code_mem[201][3] ;
 wire \mem.mem_internal.code_mem[201][4] ;
 wire \mem.mem_internal.code_mem[201][5] ;
 wire \mem.mem_internal.code_mem[201][6] ;
 wire \mem.mem_internal.code_mem[201][7] ;
 wire \mem.mem_internal.code_mem[202][0] ;
 wire \mem.mem_internal.code_mem[202][1] ;
 wire \mem.mem_internal.code_mem[202][2] ;
 wire \mem.mem_internal.code_mem[202][3] ;
 wire \mem.mem_internal.code_mem[202][4] ;
 wire \mem.mem_internal.code_mem[202][5] ;
 wire \mem.mem_internal.code_mem[202][6] ;
 wire \mem.mem_internal.code_mem[202][7] ;
 wire \mem.mem_internal.code_mem[203][0] ;
 wire \mem.mem_internal.code_mem[203][1] ;
 wire \mem.mem_internal.code_mem[203][2] ;
 wire \mem.mem_internal.code_mem[203][3] ;
 wire \mem.mem_internal.code_mem[203][4] ;
 wire \mem.mem_internal.code_mem[203][5] ;
 wire \mem.mem_internal.code_mem[203][6] ;
 wire \mem.mem_internal.code_mem[203][7] ;
 wire \mem.mem_internal.code_mem[204][0] ;
 wire \mem.mem_internal.code_mem[204][1] ;
 wire \mem.mem_internal.code_mem[204][2] ;
 wire \mem.mem_internal.code_mem[204][3] ;
 wire \mem.mem_internal.code_mem[204][4] ;
 wire \mem.mem_internal.code_mem[204][5] ;
 wire \mem.mem_internal.code_mem[204][6] ;
 wire \mem.mem_internal.code_mem[204][7] ;
 wire \mem.mem_internal.code_mem[205][0] ;
 wire \mem.mem_internal.code_mem[205][1] ;
 wire \mem.mem_internal.code_mem[205][2] ;
 wire \mem.mem_internal.code_mem[205][3] ;
 wire \mem.mem_internal.code_mem[205][4] ;
 wire \mem.mem_internal.code_mem[205][5] ;
 wire \mem.mem_internal.code_mem[205][6] ;
 wire \mem.mem_internal.code_mem[205][7] ;
 wire \mem.mem_internal.code_mem[206][0] ;
 wire \mem.mem_internal.code_mem[206][1] ;
 wire \mem.mem_internal.code_mem[206][2] ;
 wire \mem.mem_internal.code_mem[206][3] ;
 wire \mem.mem_internal.code_mem[206][4] ;
 wire \mem.mem_internal.code_mem[206][5] ;
 wire \mem.mem_internal.code_mem[206][6] ;
 wire \mem.mem_internal.code_mem[206][7] ;
 wire \mem.mem_internal.code_mem[207][0] ;
 wire \mem.mem_internal.code_mem[207][1] ;
 wire \mem.mem_internal.code_mem[207][2] ;
 wire \mem.mem_internal.code_mem[207][3] ;
 wire \mem.mem_internal.code_mem[207][4] ;
 wire \mem.mem_internal.code_mem[207][5] ;
 wire \mem.mem_internal.code_mem[207][6] ;
 wire \mem.mem_internal.code_mem[207][7] ;
 wire \mem.mem_internal.code_mem[208][0] ;
 wire \mem.mem_internal.code_mem[208][1] ;
 wire \mem.mem_internal.code_mem[208][2] ;
 wire \mem.mem_internal.code_mem[208][3] ;
 wire \mem.mem_internal.code_mem[208][4] ;
 wire \mem.mem_internal.code_mem[208][5] ;
 wire \mem.mem_internal.code_mem[208][6] ;
 wire \mem.mem_internal.code_mem[208][7] ;
 wire \mem.mem_internal.code_mem[209][0] ;
 wire \mem.mem_internal.code_mem[209][1] ;
 wire \mem.mem_internal.code_mem[209][2] ;
 wire \mem.mem_internal.code_mem[209][3] ;
 wire \mem.mem_internal.code_mem[209][4] ;
 wire \mem.mem_internal.code_mem[209][5] ;
 wire \mem.mem_internal.code_mem[209][6] ;
 wire \mem.mem_internal.code_mem[209][7] ;
 wire \mem.mem_internal.code_mem[20][0] ;
 wire \mem.mem_internal.code_mem[20][1] ;
 wire \mem.mem_internal.code_mem[20][2] ;
 wire \mem.mem_internal.code_mem[20][3] ;
 wire \mem.mem_internal.code_mem[20][4] ;
 wire \mem.mem_internal.code_mem[20][5] ;
 wire \mem.mem_internal.code_mem[20][6] ;
 wire \mem.mem_internal.code_mem[20][7] ;
 wire \mem.mem_internal.code_mem[210][0] ;
 wire \mem.mem_internal.code_mem[210][1] ;
 wire \mem.mem_internal.code_mem[210][2] ;
 wire \mem.mem_internal.code_mem[210][3] ;
 wire \mem.mem_internal.code_mem[210][4] ;
 wire \mem.mem_internal.code_mem[210][5] ;
 wire \mem.mem_internal.code_mem[210][6] ;
 wire \mem.mem_internal.code_mem[210][7] ;
 wire \mem.mem_internal.code_mem[211][0] ;
 wire \mem.mem_internal.code_mem[211][1] ;
 wire \mem.mem_internal.code_mem[211][2] ;
 wire \mem.mem_internal.code_mem[211][3] ;
 wire \mem.mem_internal.code_mem[211][4] ;
 wire \mem.mem_internal.code_mem[211][5] ;
 wire \mem.mem_internal.code_mem[211][6] ;
 wire \mem.mem_internal.code_mem[211][7] ;
 wire \mem.mem_internal.code_mem[212][0] ;
 wire \mem.mem_internal.code_mem[212][1] ;
 wire \mem.mem_internal.code_mem[212][2] ;
 wire \mem.mem_internal.code_mem[212][3] ;
 wire \mem.mem_internal.code_mem[212][4] ;
 wire \mem.mem_internal.code_mem[212][5] ;
 wire \mem.mem_internal.code_mem[212][6] ;
 wire \mem.mem_internal.code_mem[212][7] ;
 wire \mem.mem_internal.code_mem[213][0] ;
 wire \mem.mem_internal.code_mem[213][1] ;
 wire \mem.mem_internal.code_mem[213][2] ;
 wire \mem.mem_internal.code_mem[213][3] ;
 wire \mem.mem_internal.code_mem[213][4] ;
 wire \mem.mem_internal.code_mem[213][5] ;
 wire \mem.mem_internal.code_mem[213][6] ;
 wire \mem.mem_internal.code_mem[213][7] ;
 wire \mem.mem_internal.code_mem[214][0] ;
 wire \mem.mem_internal.code_mem[214][1] ;
 wire \mem.mem_internal.code_mem[214][2] ;
 wire \mem.mem_internal.code_mem[214][3] ;
 wire \mem.mem_internal.code_mem[214][4] ;
 wire \mem.mem_internal.code_mem[214][5] ;
 wire \mem.mem_internal.code_mem[214][6] ;
 wire \mem.mem_internal.code_mem[214][7] ;
 wire \mem.mem_internal.code_mem[215][0] ;
 wire \mem.mem_internal.code_mem[215][1] ;
 wire \mem.mem_internal.code_mem[215][2] ;
 wire \mem.mem_internal.code_mem[215][3] ;
 wire \mem.mem_internal.code_mem[215][4] ;
 wire \mem.mem_internal.code_mem[215][5] ;
 wire \mem.mem_internal.code_mem[215][6] ;
 wire \mem.mem_internal.code_mem[215][7] ;
 wire \mem.mem_internal.code_mem[216][0] ;
 wire \mem.mem_internal.code_mem[216][1] ;
 wire \mem.mem_internal.code_mem[216][2] ;
 wire \mem.mem_internal.code_mem[216][3] ;
 wire \mem.mem_internal.code_mem[216][4] ;
 wire \mem.mem_internal.code_mem[216][5] ;
 wire \mem.mem_internal.code_mem[216][6] ;
 wire \mem.mem_internal.code_mem[216][7] ;
 wire \mem.mem_internal.code_mem[217][0] ;
 wire \mem.mem_internal.code_mem[217][1] ;
 wire \mem.mem_internal.code_mem[217][2] ;
 wire \mem.mem_internal.code_mem[217][3] ;
 wire \mem.mem_internal.code_mem[217][4] ;
 wire \mem.mem_internal.code_mem[217][5] ;
 wire \mem.mem_internal.code_mem[217][6] ;
 wire \mem.mem_internal.code_mem[217][7] ;
 wire \mem.mem_internal.code_mem[218][0] ;
 wire \mem.mem_internal.code_mem[218][1] ;
 wire \mem.mem_internal.code_mem[218][2] ;
 wire \mem.mem_internal.code_mem[218][3] ;
 wire \mem.mem_internal.code_mem[218][4] ;
 wire \mem.mem_internal.code_mem[218][5] ;
 wire \mem.mem_internal.code_mem[218][6] ;
 wire \mem.mem_internal.code_mem[218][7] ;
 wire \mem.mem_internal.code_mem[219][0] ;
 wire \mem.mem_internal.code_mem[219][1] ;
 wire \mem.mem_internal.code_mem[219][2] ;
 wire \mem.mem_internal.code_mem[219][3] ;
 wire \mem.mem_internal.code_mem[219][4] ;
 wire \mem.mem_internal.code_mem[219][5] ;
 wire \mem.mem_internal.code_mem[219][6] ;
 wire \mem.mem_internal.code_mem[219][7] ;
 wire \mem.mem_internal.code_mem[21][0] ;
 wire \mem.mem_internal.code_mem[21][1] ;
 wire \mem.mem_internal.code_mem[21][2] ;
 wire \mem.mem_internal.code_mem[21][3] ;
 wire \mem.mem_internal.code_mem[21][4] ;
 wire \mem.mem_internal.code_mem[21][5] ;
 wire \mem.mem_internal.code_mem[21][6] ;
 wire \mem.mem_internal.code_mem[21][7] ;
 wire \mem.mem_internal.code_mem[220][0] ;
 wire \mem.mem_internal.code_mem[220][1] ;
 wire \mem.mem_internal.code_mem[220][2] ;
 wire \mem.mem_internal.code_mem[220][3] ;
 wire \mem.mem_internal.code_mem[220][4] ;
 wire \mem.mem_internal.code_mem[220][5] ;
 wire \mem.mem_internal.code_mem[220][6] ;
 wire \mem.mem_internal.code_mem[220][7] ;
 wire \mem.mem_internal.code_mem[221][0] ;
 wire \mem.mem_internal.code_mem[221][1] ;
 wire \mem.mem_internal.code_mem[221][2] ;
 wire \mem.mem_internal.code_mem[221][3] ;
 wire \mem.mem_internal.code_mem[221][4] ;
 wire \mem.mem_internal.code_mem[221][5] ;
 wire \mem.mem_internal.code_mem[221][6] ;
 wire \mem.mem_internal.code_mem[221][7] ;
 wire \mem.mem_internal.code_mem[222][0] ;
 wire \mem.mem_internal.code_mem[222][1] ;
 wire \mem.mem_internal.code_mem[222][2] ;
 wire \mem.mem_internal.code_mem[222][3] ;
 wire \mem.mem_internal.code_mem[222][4] ;
 wire \mem.mem_internal.code_mem[222][5] ;
 wire \mem.mem_internal.code_mem[222][6] ;
 wire \mem.mem_internal.code_mem[222][7] ;
 wire \mem.mem_internal.code_mem[223][0] ;
 wire \mem.mem_internal.code_mem[223][1] ;
 wire \mem.mem_internal.code_mem[223][2] ;
 wire \mem.mem_internal.code_mem[223][3] ;
 wire \mem.mem_internal.code_mem[223][4] ;
 wire \mem.mem_internal.code_mem[223][5] ;
 wire \mem.mem_internal.code_mem[223][6] ;
 wire \mem.mem_internal.code_mem[223][7] ;
 wire \mem.mem_internal.code_mem[224][0] ;
 wire \mem.mem_internal.code_mem[224][1] ;
 wire \mem.mem_internal.code_mem[224][2] ;
 wire \mem.mem_internal.code_mem[224][3] ;
 wire \mem.mem_internal.code_mem[224][4] ;
 wire \mem.mem_internal.code_mem[224][5] ;
 wire \mem.mem_internal.code_mem[224][6] ;
 wire \mem.mem_internal.code_mem[224][7] ;
 wire \mem.mem_internal.code_mem[225][0] ;
 wire \mem.mem_internal.code_mem[225][1] ;
 wire \mem.mem_internal.code_mem[225][2] ;
 wire \mem.mem_internal.code_mem[225][3] ;
 wire \mem.mem_internal.code_mem[225][4] ;
 wire \mem.mem_internal.code_mem[225][5] ;
 wire \mem.mem_internal.code_mem[225][6] ;
 wire \mem.mem_internal.code_mem[225][7] ;
 wire \mem.mem_internal.code_mem[226][0] ;
 wire \mem.mem_internal.code_mem[226][1] ;
 wire \mem.mem_internal.code_mem[226][2] ;
 wire \mem.mem_internal.code_mem[226][3] ;
 wire \mem.mem_internal.code_mem[226][4] ;
 wire \mem.mem_internal.code_mem[226][5] ;
 wire \mem.mem_internal.code_mem[226][6] ;
 wire \mem.mem_internal.code_mem[226][7] ;
 wire \mem.mem_internal.code_mem[227][0] ;
 wire \mem.mem_internal.code_mem[227][1] ;
 wire \mem.mem_internal.code_mem[227][2] ;
 wire \mem.mem_internal.code_mem[227][3] ;
 wire \mem.mem_internal.code_mem[227][4] ;
 wire \mem.mem_internal.code_mem[227][5] ;
 wire \mem.mem_internal.code_mem[227][6] ;
 wire \mem.mem_internal.code_mem[227][7] ;
 wire \mem.mem_internal.code_mem[228][0] ;
 wire \mem.mem_internal.code_mem[228][1] ;
 wire \mem.mem_internal.code_mem[228][2] ;
 wire \mem.mem_internal.code_mem[228][3] ;
 wire \mem.mem_internal.code_mem[228][4] ;
 wire \mem.mem_internal.code_mem[228][5] ;
 wire \mem.mem_internal.code_mem[228][6] ;
 wire \mem.mem_internal.code_mem[228][7] ;
 wire \mem.mem_internal.code_mem[229][0] ;
 wire \mem.mem_internal.code_mem[229][1] ;
 wire \mem.mem_internal.code_mem[229][2] ;
 wire \mem.mem_internal.code_mem[229][3] ;
 wire \mem.mem_internal.code_mem[229][4] ;
 wire \mem.mem_internal.code_mem[229][5] ;
 wire \mem.mem_internal.code_mem[229][6] ;
 wire \mem.mem_internal.code_mem[229][7] ;
 wire \mem.mem_internal.code_mem[22][0] ;
 wire \mem.mem_internal.code_mem[22][1] ;
 wire \mem.mem_internal.code_mem[22][2] ;
 wire \mem.mem_internal.code_mem[22][3] ;
 wire \mem.mem_internal.code_mem[22][4] ;
 wire \mem.mem_internal.code_mem[22][5] ;
 wire \mem.mem_internal.code_mem[22][6] ;
 wire \mem.mem_internal.code_mem[22][7] ;
 wire \mem.mem_internal.code_mem[230][0] ;
 wire \mem.mem_internal.code_mem[230][1] ;
 wire \mem.mem_internal.code_mem[230][2] ;
 wire \mem.mem_internal.code_mem[230][3] ;
 wire \mem.mem_internal.code_mem[230][4] ;
 wire \mem.mem_internal.code_mem[230][5] ;
 wire \mem.mem_internal.code_mem[230][6] ;
 wire \mem.mem_internal.code_mem[230][7] ;
 wire \mem.mem_internal.code_mem[231][0] ;
 wire \mem.mem_internal.code_mem[231][1] ;
 wire \mem.mem_internal.code_mem[231][2] ;
 wire \mem.mem_internal.code_mem[231][3] ;
 wire \mem.mem_internal.code_mem[231][4] ;
 wire \mem.mem_internal.code_mem[231][5] ;
 wire \mem.mem_internal.code_mem[231][6] ;
 wire \mem.mem_internal.code_mem[231][7] ;
 wire \mem.mem_internal.code_mem[232][0] ;
 wire \mem.mem_internal.code_mem[232][1] ;
 wire \mem.mem_internal.code_mem[232][2] ;
 wire \mem.mem_internal.code_mem[232][3] ;
 wire \mem.mem_internal.code_mem[232][4] ;
 wire \mem.mem_internal.code_mem[232][5] ;
 wire \mem.mem_internal.code_mem[232][6] ;
 wire \mem.mem_internal.code_mem[232][7] ;
 wire \mem.mem_internal.code_mem[233][0] ;
 wire \mem.mem_internal.code_mem[233][1] ;
 wire \mem.mem_internal.code_mem[233][2] ;
 wire \mem.mem_internal.code_mem[233][3] ;
 wire \mem.mem_internal.code_mem[233][4] ;
 wire \mem.mem_internal.code_mem[233][5] ;
 wire \mem.mem_internal.code_mem[233][6] ;
 wire \mem.mem_internal.code_mem[233][7] ;
 wire \mem.mem_internal.code_mem[234][0] ;
 wire \mem.mem_internal.code_mem[234][1] ;
 wire \mem.mem_internal.code_mem[234][2] ;
 wire \mem.mem_internal.code_mem[234][3] ;
 wire \mem.mem_internal.code_mem[234][4] ;
 wire \mem.mem_internal.code_mem[234][5] ;
 wire \mem.mem_internal.code_mem[234][6] ;
 wire \mem.mem_internal.code_mem[234][7] ;
 wire \mem.mem_internal.code_mem[235][0] ;
 wire \mem.mem_internal.code_mem[235][1] ;
 wire \mem.mem_internal.code_mem[235][2] ;
 wire \mem.mem_internal.code_mem[235][3] ;
 wire \mem.mem_internal.code_mem[235][4] ;
 wire \mem.mem_internal.code_mem[235][5] ;
 wire \mem.mem_internal.code_mem[235][6] ;
 wire \mem.mem_internal.code_mem[235][7] ;
 wire \mem.mem_internal.code_mem[236][0] ;
 wire \mem.mem_internal.code_mem[236][1] ;
 wire \mem.mem_internal.code_mem[236][2] ;
 wire \mem.mem_internal.code_mem[236][3] ;
 wire \mem.mem_internal.code_mem[236][4] ;
 wire \mem.mem_internal.code_mem[236][5] ;
 wire \mem.mem_internal.code_mem[236][6] ;
 wire \mem.mem_internal.code_mem[236][7] ;
 wire \mem.mem_internal.code_mem[237][0] ;
 wire \mem.mem_internal.code_mem[237][1] ;
 wire \mem.mem_internal.code_mem[237][2] ;
 wire \mem.mem_internal.code_mem[237][3] ;
 wire \mem.mem_internal.code_mem[237][4] ;
 wire \mem.mem_internal.code_mem[237][5] ;
 wire \mem.mem_internal.code_mem[237][6] ;
 wire \mem.mem_internal.code_mem[237][7] ;
 wire \mem.mem_internal.code_mem[238][0] ;
 wire \mem.mem_internal.code_mem[238][1] ;
 wire \mem.mem_internal.code_mem[238][2] ;
 wire \mem.mem_internal.code_mem[238][3] ;
 wire \mem.mem_internal.code_mem[238][4] ;
 wire \mem.mem_internal.code_mem[238][5] ;
 wire \mem.mem_internal.code_mem[238][6] ;
 wire \mem.mem_internal.code_mem[238][7] ;
 wire \mem.mem_internal.code_mem[239][0] ;
 wire \mem.mem_internal.code_mem[239][1] ;
 wire \mem.mem_internal.code_mem[239][2] ;
 wire \mem.mem_internal.code_mem[239][3] ;
 wire \mem.mem_internal.code_mem[239][4] ;
 wire \mem.mem_internal.code_mem[239][5] ;
 wire \mem.mem_internal.code_mem[239][6] ;
 wire \mem.mem_internal.code_mem[239][7] ;
 wire \mem.mem_internal.code_mem[23][0] ;
 wire \mem.mem_internal.code_mem[23][1] ;
 wire \mem.mem_internal.code_mem[23][2] ;
 wire \mem.mem_internal.code_mem[23][3] ;
 wire \mem.mem_internal.code_mem[23][4] ;
 wire \mem.mem_internal.code_mem[23][5] ;
 wire \mem.mem_internal.code_mem[23][6] ;
 wire \mem.mem_internal.code_mem[23][7] ;
 wire \mem.mem_internal.code_mem[240][0] ;
 wire \mem.mem_internal.code_mem[240][1] ;
 wire \mem.mem_internal.code_mem[240][2] ;
 wire \mem.mem_internal.code_mem[240][3] ;
 wire \mem.mem_internal.code_mem[240][4] ;
 wire \mem.mem_internal.code_mem[240][5] ;
 wire \mem.mem_internal.code_mem[240][6] ;
 wire \mem.mem_internal.code_mem[240][7] ;
 wire \mem.mem_internal.code_mem[241][0] ;
 wire \mem.mem_internal.code_mem[241][1] ;
 wire \mem.mem_internal.code_mem[241][2] ;
 wire \mem.mem_internal.code_mem[241][3] ;
 wire \mem.mem_internal.code_mem[241][4] ;
 wire \mem.mem_internal.code_mem[241][5] ;
 wire \mem.mem_internal.code_mem[241][6] ;
 wire \mem.mem_internal.code_mem[241][7] ;
 wire \mem.mem_internal.code_mem[242][0] ;
 wire \mem.mem_internal.code_mem[242][1] ;
 wire \mem.mem_internal.code_mem[242][2] ;
 wire \mem.mem_internal.code_mem[242][3] ;
 wire \mem.mem_internal.code_mem[242][4] ;
 wire \mem.mem_internal.code_mem[242][5] ;
 wire \mem.mem_internal.code_mem[242][6] ;
 wire \mem.mem_internal.code_mem[242][7] ;
 wire \mem.mem_internal.code_mem[243][0] ;
 wire \mem.mem_internal.code_mem[243][1] ;
 wire \mem.mem_internal.code_mem[243][2] ;
 wire \mem.mem_internal.code_mem[243][3] ;
 wire \mem.mem_internal.code_mem[243][4] ;
 wire \mem.mem_internal.code_mem[243][5] ;
 wire \mem.mem_internal.code_mem[243][6] ;
 wire \mem.mem_internal.code_mem[243][7] ;
 wire \mem.mem_internal.code_mem[244][0] ;
 wire \mem.mem_internal.code_mem[244][1] ;
 wire \mem.mem_internal.code_mem[244][2] ;
 wire \mem.mem_internal.code_mem[244][3] ;
 wire \mem.mem_internal.code_mem[244][4] ;
 wire \mem.mem_internal.code_mem[244][5] ;
 wire \mem.mem_internal.code_mem[244][6] ;
 wire \mem.mem_internal.code_mem[244][7] ;
 wire \mem.mem_internal.code_mem[245][0] ;
 wire \mem.mem_internal.code_mem[245][1] ;
 wire \mem.mem_internal.code_mem[245][2] ;
 wire \mem.mem_internal.code_mem[245][3] ;
 wire \mem.mem_internal.code_mem[245][4] ;
 wire \mem.mem_internal.code_mem[245][5] ;
 wire \mem.mem_internal.code_mem[245][6] ;
 wire \mem.mem_internal.code_mem[245][7] ;
 wire \mem.mem_internal.code_mem[246][0] ;
 wire \mem.mem_internal.code_mem[246][1] ;
 wire \mem.mem_internal.code_mem[246][2] ;
 wire \mem.mem_internal.code_mem[246][3] ;
 wire \mem.mem_internal.code_mem[246][4] ;
 wire \mem.mem_internal.code_mem[246][5] ;
 wire \mem.mem_internal.code_mem[246][6] ;
 wire \mem.mem_internal.code_mem[246][7] ;
 wire \mem.mem_internal.code_mem[247][0] ;
 wire \mem.mem_internal.code_mem[247][1] ;
 wire \mem.mem_internal.code_mem[247][2] ;
 wire \mem.mem_internal.code_mem[247][3] ;
 wire \mem.mem_internal.code_mem[247][4] ;
 wire \mem.mem_internal.code_mem[247][5] ;
 wire \mem.mem_internal.code_mem[247][6] ;
 wire \mem.mem_internal.code_mem[247][7] ;
 wire \mem.mem_internal.code_mem[248][0] ;
 wire \mem.mem_internal.code_mem[248][1] ;
 wire \mem.mem_internal.code_mem[248][2] ;
 wire \mem.mem_internal.code_mem[248][3] ;
 wire \mem.mem_internal.code_mem[248][4] ;
 wire \mem.mem_internal.code_mem[248][5] ;
 wire \mem.mem_internal.code_mem[248][6] ;
 wire \mem.mem_internal.code_mem[248][7] ;
 wire \mem.mem_internal.code_mem[249][0] ;
 wire \mem.mem_internal.code_mem[249][1] ;
 wire \mem.mem_internal.code_mem[249][2] ;
 wire \mem.mem_internal.code_mem[249][3] ;
 wire \mem.mem_internal.code_mem[249][4] ;
 wire \mem.mem_internal.code_mem[249][5] ;
 wire \mem.mem_internal.code_mem[249][6] ;
 wire \mem.mem_internal.code_mem[249][7] ;
 wire \mem.mem_internal.code_mem[24][0] ;
 wire \mem.mem_internal.code_mem[24][1] ;
 wire \mem.mem_internal.code_mem[24][2] ;
 wire \mem.mem_internal.code_mem[24][3] ;
 wire \mem.mem_internal.code_mem[24][4] ;
 wire \mem.mem_internal.code_mem[24][5] ;
 wire \mem.mem_internal.code_mem[24][6] ;
 wire \mem.mem_internal.code_mem[24][7] ;
 wire \mem.mem_internal.code_mem[250][0] ;
 wire \mem.mem_internal.code_mem[250][1] ;
 wire \mem.mem_internal.code_mem[250][2] ;
 wire \mem.mem_internal.code_mem[250][3] ;
 wire \mem.mem_internal.code_mem[250][4] ;
 wire \mem.mem_internal.code_mem[250][5] ;
 wire \mem.mem_internal.code_mem[250][6] ;
 wire \mem.mem_internal.code_mem[250][7] ;
 wire \mem.mem_internal.code_mem[251][0] ;
 wire \mem.mem_internal.code_mem[251][1] ;
 wire \mem.mem_internal.code_mem[251][2] ;
 wire \mem.mem_internal.code_mem[251][3] ;
 wire \mem.mem_internal.code_mem[251][4] ;
 wire \mem.mem_internal.code_mem[251][5] ;
 wire \mem.mem_internal.code_mem[251][6] ;
 wire \mem.mem_internal.code_mem[251][7] ;
 wire \mem.mem_internal.code_mem[252][0] ;
 wire \mem.mem_internal.code_mem[252][1] ;
 wire \mem.mem_internal.code_mem[252][2] ;
 wire \mem.mem_internal.code_mem[252][3] ;
 wire \mem.mem_internal.code_mem[252][4] ;
 wire \mem.mem_internal.code_mem[252][5] ;
 wire \mem.mem_internal.code_mem[252][6] ;
 wire \mem.mem_internal.code_mem[252][7] ;
 wire \mem.mem_internal.code_mem[253][0] ;
 wire \mem.mem_internal.code_mem[253][1] ;
 wire \mem.mem_internal.code_mem[253][2] ;
 wire \mem.mem_internal.code_mem[253][3] ;
 wire \mem.mem_internal.code_mem[253][4] ;
 wire \mem.mem_internal.code_mem[253][5] ;
 wire \mem.mem_internal.code_mem[253][6] ;
 wire \mem.mem_internal.code_mem[253][7] ;
 wire \mem.mem_internal.code_mem[254][0] ;
 wire \mem.mem_internal.code_mem[254][1] ;
 wire \mem.mem_internal.code_mem[254][2] ;
 wire \mem.mem_internal.code_mem[254][3] ;
 wire \mem.mem_internal.code_mem[254][4] ;
 wire \mem.mem_internal.code_mem[254][5] ;
 wire \mem.mem_internal.code_mem[254][6] ;
 wire \mem.mem_internal.code_mem[254][7] ;
 wire \mem.mem_internal.code_mem[255][0] ;
 wire \mem.mem_internal.code_mem[255][1] ;
 wire \mem.mem_internal.code_mem[255][2] ;
 wire \mem.mem_internal.code_mem[255][3] ;
 wire \mem.mem_internal.code_mem[255][4] ;
 wire \mem.mem_internal.code_mem[255][5] ;
 wire \mem.mem_internal.code_mem[255][6] ;
 wire \mem.mem_internal.code_mem[255][7] ;
 wire \mem.mem_internal.code_mem[25][0] ;
 wire \mem.mem_internal.code_mem[25][1] ;
 wire \mem.mem_internal.code_mem[25][2] ;
 wire \mem.mem_internal.code_mem[25][3] ;
 wire \mem.mem_internal.code_mem[25][4] ;
 wire \mem.mem_internal.code_mem[25][5] ;
 wire \mem.mem_internal.code_mem[25][6] ;
 wire \mem.mem_internal.code_mem[25][7] ;
 wire \mem.mem_internal.code_mem[26][0] ;
 wire \mem.mem_internal.code_mem[26][1] ;
 wire \mem.mem_internal.code_mem[26][2] ;
 wire \mem.mem_internal.code_mem[26][3] ;
 wire \mem.mem_internal.code_mem[26][4] ;
 wire \mem.mem_internal.code_mem[26][5] ;
 wire \mem.mem_internal.code_mem[26][6] ;
 wire \mem.mem_internal.code_mem[26][7] ;
 wire \mem.mem_internal.code_mem[27][0] ;
 wire \mem.mem_internal.code_mem[27][1] ;
 wire \mem.mem_internal.code_mem[27][2] ;
 wire \mem.mem_internal.code_mem[27][3] ;
 wire \mem.mem_internal.code_mem[27][4] ;
 wire \mem.mem_internal.code_mem[27][5] ;
 wire \mem.mem_internal.code_mem[27][6] ;
 wire \mem.mem_internal.code_mem[27][7] ;
 wire \mem.mem_internal.code_mem[28][0] ;
 wire \mem.mem_internal.code_mem[28][1] ;
 wire \mem.mem_internal.code_mem[28][2] ;
 wire \mem.mem_internal.code_mem[28][3] ;
 wire \mem.mem_internal.code_mem[28][4] ;
 wire \mem.mem_internal.code_mem[28][5] ;
 wire \mem.mem_internal.code_mem[28][6] ;
 wire \mem.mem_internal.code_mem[28][7] ;
 wire \mem.mem_internal.code_mem[29][0] ;
 wire \mem.mem_internal.code_mem[29][1] ;
 wire \mem.mem_internal.code_mem[29][2] ;
 wire \mem.mem_internal.code_mem[29][3] ;
 wire \mem.mem_internal.code_mem[29][4] ;
 wire \mem.mem_internal.code_mem[29][5] ;
 wire \mem.mem_internal.code_mem[29][6] ;
 wire \mem.mem_internal.code_mem[29][7] ;
 wire \mem.mem_internal.code_mem[2][0] ;
 wire \mem.mem_internal.code_mem[2][1] ;
 wire \mem.mem_internal.code_mem[2][2] ;
 wire \mem.mem_internal.code_mem[2][3] ;
 wire \mem.mem_internal.code_mem[2][4] ;
 wire \mem.mem_internal.code_mem[2][5] ;
 wire \mem.mem_internal.code_mem[2][6] ;
 wire \mem.mem_internal.code_mem[2][7] ;
 wire \mem.mem_internal.code_mem[30][0] ;
 wire \mem.mem_internal.code_mem[30][1] ;
 wire \mem.mem_internal.code_mem[30][2] ;
 wire \mem.mem_internal.code_mem[30][3] ;
 wire \mem.mem_internal.code_mem[30][4] ;
 wire \mem.mem_internal.code_mem[30][5] ;
 wire \mem.mem_internal.code_mem[30][6] ;
 wire \mem.mem_internal.code_mem[30][7] ;
 wire \mem.mem_internal.code_mem[31][0] ;
 wire \mem.mem_internal.code_mem[31][1] ;
 wire \mem.mem_internal.code_mem[31][2] ;
 wire \mem.mem_internal.code_mem[31][3] ;
 wire \mem.mem_internal.code_mem[31][4] ;
 wire \mem.mem_internal.code_mem[31][5] ;
 wire \mem.mem_internal.code_mem[31][6] ;
 wire \mem.mem_internal.code_mem[31][7] ;
 wire \mem.mem_internal.code_mem[32][0] ;
 wire \mem.mem_internal.code_mem[32][1] ;
 wire \mem.mem_internal.code_mem[32][2] ;
 wire \mem.mem_internal.code_mem[32][3] ;
 wire \mem.mem_internal.code_mem[32][4] ;
 wire \mem.mem_internal.code_mem[32][5] ;
 wire \mem.mem_internal.code_mem[32][6] ;
 wire \mem.mem_internal.code_mem[32][7] ;
 wire \mem.mem_internal.code_mem[33][0] ;
 wire \mem.mem_internal.code_mem[33][1] ;
 wire \mem.mem_internal.code_mem[33][2] ;
 wire \mem.mem_internal.code_mem[33][3] ;
 wire \mem.mem_internal.code_mem[33][4] ;
 wire \mem.mem_internal.code_mem[33][5] ;
 wire \mem.mem_internal.code_mem[33][6] ;
 wire \mem.mem_internal.code_mem[33][7] ;
 wire \mem.mem_internal.code_mem[34][0] ;
 wire \mem.mem_internal.code_mem[34][1] ;
 wire \mem.mem_internal.code_mem[34][2] ;
 wire \mem.mem_internal.code_mem[34][3] ;
 wire \mem.mem_internal.code_mem[34][4] ;
 wire \mem.mem_internal.code_mem[34][5] ;
 wire \mem.mem_internal.code_mem[34][6] ;
 wire \mem.mem_internal.code_mem[34][7] ;
 wire \mem.mem_internal.code_mem[35][0] ;
 wire \mem.mem_internal.code_mem[35][1] ;
 wire \mem.mem_internal.code_mem[35][2] ;
 wire \mem.mem_internal.code_mem[35][3] ;
 wire \mem.mem_internal.code_mem[35][4] ;
 wire \mem.mem_internal.code_mem[35][5] ;
 wire \mem.mem_internal.code_mem[35][6] ;
 wire \mem.mem_internal.code_mem[35][7] ;
 wire \mem.mem_internal.code_mem[36][0] ;
 wire \mem.mem_internal.code_mem[36][1] ;
 wire \mem.mem_internal.code_mem[36][2] ;
 wire \mem.mem_internal.code_mem[36][3] ;
 wire \mem.mem_internal.code_mem[36][4] ;
 wire \mem.mem_internal.code_mem[36][5] ;
 wire \mem.mem_internal.code_mem[36][6] ;
 wire \mem.mem_internal.code_mem[36][7] ;
 wire \mem.mem_internal.code_mem[37][0] ;
 wire \mem.mem_internal.code_mem[37][1] ;
 wire \mem.mem_internal.code_mem[37][2] ;
 wire \mem.mem_internal.code_mem[37][3] ;
 wire \mem.mem_internal.code_mem[37][4] ;
 wire \mem.mem_internal.code_mem[37][5] ;
 wire \mem.mem_internal.code_mem[37][6] ;
 wire \mem.mem_internal.code_mem[37][7] ;
 wire \mem.mem_internal.code_mem[38][0] ;
 wire \mem.mem_internal.code_mem[38][1] ;
 wire \mem.mem_internal.code_mem[38][2] ;
 wire \mem.mem_internal.code_mem[38][3] ;
 wire \mem.mem_internal.code_mem[38][4] ;
 wire \mem.mem_internal.code_mem[38][5] ;
 wire \mem.mem_internal.code_mem[38][6] ;
 wire \mem.mem_internal.code_mem[38][7] ;
 wire \mem.mem_internal.code_mem[39][0] ;
 wire \mem.mem_internal.code_mem[39][1] ;
 wire \mem.mem_internal.code_mem[39][2] ;
 wire \mem.mem_internal.code_mem[39][3] ;
 wire \mem.mem_internal.code_mem[39][4] ;
 wire \mem.mem_internal.code_mem[39][5] ;
 wire \mem.mem_internal.code_mem[39][6] ;
 wire \mem.mem_internal.code_mem[39][7] ;
 wire \mem.mem_internal.code_mem[3][0] ;
 wire \mem.mem_internal.code_mem[3][1] ;
 wire \mem.mem_internal.code_mem[3][2] ;
 wire \mem.mem_internal.code_mem[3][3] ;
 wire \mem.mem_internal.code_mem[3][4] ;
 wire \mem.mem_internal.code_mem[3][5] ;
 wire \mem.mem_internal.code_mem[3][6] ;
 wire \mem.mem_internal.code_mem[3][7] ;
 wire \mem.mem_internal.code_mem[40][0] ;
 wire \mem.mem_internal.code_mem[40][1] ;
 wire \mem.mem_internal.code_mem[40][2] ;
 wire \mem.mem_internal.code_mem[40][3] ;
 wire \mem.mem_internal.code_mem[40][4] ;
 wire \mem.mem_internal.code_mem[40][5] ;
 wire \mem.mem_internal.code_mem[40][6] ;
 wire \mem.mem_internal.code_mem[40][7] ;
 wire \mem.mem_internal.code_mem[41][0] ;
 wire \mem.mem_internal.code_mem[41][1] ;
 wire \mem.mem_internal.code_mem[41][2] ;
 wire \mem.mem_internal.code_mem[41][3] ;
 wire \mem.mem_internal.code_mem[41][4] ;
 wire \mem.mem_internal.code_mem[41][5] ;
 wire \mem.mem_internal.code_mem[41][6] ;
 wire \mem.mem_internal.code_mem[41][7] ;
 wire \mem.mem_internal.code_mem[42][0] ;
 wire \mem.mem_internal.code_mem[42][1] ;
 wire \mem.mem_internal.code_mem[42][2] ;
 wire \mem.mem_internal.code_mem[42][3] ;
 wire \mem.mem_internal.code_mem[42][4] ;
 wire \mem.mem_internal.code_mem[42][5] ;
 wire \mem.mem_internal.code_mem[42][6] ;
 wire \mem.mem_internal.code_mem[42][7] ;
 wire \mem.mem_internal.code_mem[43][0] ;
 wire \mem.mem_internal.code_mem[43][1] ;
 wire \mem.mem_internal.code_mem[43][2] ;
 wire \mem.mem_internal.code_mem[43][3] ;
 wire \mem.mem_internal.code_mem[43][4] ;
 wire \mem.mem_internal.code_mem[43][5] ;
 wire \mem.mem_internal.code_mem[43][6] ;
 wire \mem.mem_internal.code_mem[43][7] ;
 wire \mem.mem_internal.code_mem[44][0] ;
 wire \mem.mem_internal.code_mem[44][1] ;
 wire \mem.mem_internal.code_mem[44][2] ;
 wire \mem.mem_internal.code_mem[44][3] ;
 wire \mem.mem_internal.code_mem[44][4] ;
 wire \mem.mem_internal.code_mem[44][5] ;
 wire \mem.mem_internal.code_mem[44][6] ;
 wire \mem.mem_internal.code_mem[44][7] ;
 wire \mem.mem_internal.code_mem[45][0] ;
 wire \mem.mem_internal.code_mem[45][1] ;
 wire \mem.mem_internal.code_mem[45][2] ;
 wire \mem.mem_internal.code_mem[45][3] ;
 wire \mem.mem_internal.code_mem[45][4] ;
 wire \mem.mem_internal.code_mem[45][5] ;
 wire \mem.mem_internal.code_mem[45][6] ;
 wire \mem.mem_internal.code_mem[45][7] ;
 wire \mem.mem_internal.code_mem[46][0] ;
 wire \mem.mem_internal.code_mem[46][1] ;
 wire \mem.mem_internal.code_mem[46][2] ;
 wire \mem.mem_internal.code_mem[46][3] ;
 wire \mem.mem_internal.code_mem[46][4] ;
 wire \mem.mem_internal.code_mem[46][5] ;
 wire \mem.mem_internal.code_mem[46][6] ;
 wire \mem.mem_internal.code_mem[46][7] ;
 wire \mem.mem_internal.code_mem[47][0] ;
 wire \mem.mem_internal.code_mem[47][1] ;
 wire \mem.mem_internal.code_mem[47][2] ;
 wire \mem.mem_internal.code_mem[47][3] ;
 wire \mem.mem_internal.code_mem[47][4] ;
 wire \mem.mem_internal.code_mem[47][5] ;
 wire \mem.mem_internal.code_mem[47][6] ;
 wire \mem.mem_internal.code_mem[47][7] ;
 wire \mem.mem_internal.code_mem[48][0] ;
 wire \mem.mem_internal.code_mem[48][1] ;
 wire \mem.mem_internal.code_mem[48][2] ;
 wire \mem.mem_internal.code_mem[48][3] ;
 wire \mem.mem_internal.code_mem[48][4] ;
 wire \mem.mem_internal.code_mem[48][5] ;
 wire \mem.mem_internal.code_mem[48][6] ;
 wire \mem.mem_internal.code_mem[48][7] ;
 wire \mem.mem_internal.code_mem[49][0] ;
 wire \mem.mem_internal.code_mem[49][1] ;
 wire \mem.mem_internal.code_mem[49][2] ;
 wire \mem.mem_internal.code_mem[49][3] ;
 wire \mem.mem_internal.code_mem[49][4] ;
 wire \mem.mem_internal.code_mem[49][5] ;
 wire \mem.mem_internal.code_mem[49][6] ;
 wire \mem.mem_internal.code_mem[49][7] ;
 wire \mem.mem_internal.code_mem[4][0] ;
 wire \mem.mem_internal.code_mem[4][1] ;
 wire \mem.mem_internal.code_mem[4][2] ;
 wire \mem.mem_internal.code_mem[4][3] ;
 wire \mem.mem_internal.code_mem[4][4] ;
 wire \mem.mem_internal.code_mem[4][5] ;
 wire \mem.mem_internal.code_mem[4][6] ;
 wire \mem.mem_internal.code_mem[4][7] ;
 wire \mem.mem_internal.code_mem[50][0] ;
 wire \mem.mem_internal.code_mem[50][1] ;
 wire \mem.mem_internal.code_mem[50][2] ;
 wire \mem.mem_internal.code_mem[50][3] ;
 wire \mem.mem_internal.code_mem[50][4] ;
 wire \mem.mem_internal.code_mem[50][5] ;
 wire \mem.mem_internal.code_mem[50][6] ;
 wire \mem.mem_internal.code_mem[50][7] ;
 wire \mem.mem_internal.code_mem[51][0] ;
 wire \mem.mem_internal.code_mem[51][1] ;
 wire \mem.mem_internal.code_mem[51][2] ;
 wire \mem.mem_internal.code_mem[51][3] ;
 wire \mem.mem_internal.code_mem[51][4] ;
 wire \mem.mem_internal.code_mem[51][5] ;
 wire \mem.mem_internal.code_mem[51][6] ;
 wire \mem.mem_internal.code_mem[51][7] ;
 wire \mem.mem_internal.code_mem[52][0] ;
 wire \mem.mem_internal.code_mem[52][1] ;
 wire \mem.mem_internal.code_mem[52][2] ;
 wire \mem.mem_internal.code_mem[52][3] ;
 wire \mem.mem_internal.code_mem[52][4] ;
 wire \mem.mem_internal.code_mem[52][5] ;
 wire \mem.mem_internal.code_mem[52][6] ;
 wire \mem.mem_internal.code_mem[52][7] ;
 wire \mem.mem_internal.code_mem[53][0] ;
 wire \mem.mem_internal.code_mem[53][1] ;
 wire \mem.mem_internal.code_mem[53][2] ;
 wire \mem.mem_internal.code_mem[53][3] ;
 wire \mem.mem_internal.code_mem[53][4] ;
 wire \mem.mem_internal.code_mem[53][5] ;
 wire \mem.mem_internal.code_mem[53][6] ;
 wire \mem.mem_internal.code_mem[53][7] ;
 wire \mem.mem_internal.code_mem[54][0] ;
 wire \mem.mem_internal.code_mem[54][1] ;
 wire \mem.mem_internal.code_mem[54][2] ;
 wire \mem.mem_internal.code_mem[54][3] ;
 wire \mem.mem_internal.code_mem[54][4] ;
 wire \mem.mem_internal.code_mem[54][5] ;
 wire \mem.mem_internal.code_mem[54][6] ;
 wire \mem.mem_internal.code_mem[54][7] ;
 wire \mem.mem_internal.code_mem[55][0] ;
 wire \mem.mem_internal.code_mem[55][1] ;
 wire \mem.mem_internal.code_mem[55][2] ;
 wire \mem.mem_internal.code_mem[55][3] ;
 wire \mem.mem_internal.code_mem[55][4] ;
 wire \mem.mem_internal.code_mem[55][5] ;
 wire \mem.mem_internal.code_mem[55][6] ;
 wire \mem.mem_internal.code_mem[55][7] ;
 wire \mem.mem_internal.code_mem[56][0] ;
 wire \mem.mem_internal.code_mem[56][1] ;
 wire \mem.mem_internal.code_mem[56][2] ;
 wire \mem.mem_internal.code_mem[56][3] ;
 wire \mem.mem_internal.code_mem[56][4] ;
 wire \mem.mem_internal.code_mem[56][5] ;
 wire \mem.mem_internal.code_mem[56][6] ;
 wire \mem.mem_internal.code_mem[56][7] ;
 wire \mem.mem_internal.code_mem[57][0] ;
 wire \mem.mem_internal.code_mem[57][1] ;
 wire \mem.mem_internal.code_mem[57][2] ;
 wire \mem.mem_internal.code_mem[57][3] ;
 wire \mem.mem_internal.code_mem[57][4] ;
 wire \mem.mem_internal.code_mem[57][5] ;
 wire \mem.mem_internal.code_mem[57][6] ;
 wire \mem.mem_internal.code_mem[57][7] ;
 wire \mem.mem_internal.code_mem[58][0] ;
 wire \mem.mem_internal.code_mem[58][1] ;
 wire \mem.mem_internal.code_mem[58][2] ;
 wire \mem.mem_internal.code_mem[58][3] ;
 wire \mem.mem_internal.code_mem[58][4] ;
 wire \mem.mem_internal.code_mem[58][5] ;
 wire \mem.mem_internal.code_mem[58][6] ;
 wire \mem.mem_internal.code_mem[58][7] ;
 wire \mem.mem_internal.code_mem[59][0] ;
 wire \mem.mem_internal.code_mem[59][1] ;
 wire \mem.mem_internal.code_mem[59][2] ;
 wire \mem.mem_internal.code_mem[59][3] ;
 wire \mem.mem_internal.code_mem[59][4] ;
 wire \mem.mem_internal.code_mem[59][5] ;
 wire \mem.mem_internal.code_mem[59][6] ;
 wire \mem.mem_internal.code_mem[59][7] ;
 wire \mem.mem_internal.code_mem[5][0] ;
 wire \mem.mem_internal.code_mem[5][1] ;
 wire \mem.mem_internal.code_mem[5][2] ;
 wire \mem.mem_internal.code_mem[5][3] ;
 wire \mem.mem_internal.code_mem[5][4] ;
 wire \mem.mem_internal.code_mem[5][5] ;
 wire \mem.mem_internal.code_mem[5][6] ;
 wire \mem.mem_internal.code_mem[5][7] ;
 wire \mem.mem_internal.code_mem[60][0] ;
 wire \mem.mem_internal.code_mem[60][1] ;
 wire \mem.mem_internal.code_mem[60][2] ;
 wire \mem.mem_internal.code_mem[60][3] ;
 wire \mem.mem_internal.code_mem[60][4] ;
 wire \mem.mem_internal.code_mem[60][5] ;
 wire \mem.mem_internal.code_mem[60][6] ;
 wire \mem.mem_internal.code_mem[60][7] ;
 wire \mem.mem_internal.code_mem[61][0] ;
 wire \mem.mem_internal.code_mem[61][1] ;
 wire \mem.mem_internal.code_mem[61][2] ;
 wire \mem.mem_internal.code_mem[61][3] ;
 wire \mem.mem_internal.code_mem[61][4] ;
 wire \mem.mem_internal.code_mem[61][5] ;
 wire \mem.mem_internal.code_mem[61][6] ;
 wire \mem.mem_internal.code_mem[61][7] ;
 wire \mem.mem_internal.code_mem[62][0] ;
 wire \mem.mem_internal.code_mem[62][1] ;
 wire \mem.mem_internal.code_mem[62][2] ;
 wire \mem.mem_internal.code_mem[62][3] ;
 wire \mem.mem_internal.code_mem[62][4] ;
 wire \mem.mem_internal.code_mem[62][5] ;
 wire \mem.mem_internal.code_mem[62][6] ;
 wire \mem.mem_internal.code_mem[62][7] ;
 wire \mem.mem_internal.code_mem[63][0] ;
 wire \mem.mem_internal.code_mem[63][1] ;
 wire \mem.mem_internal.code_mem[63][2] ;
 wire \mem.mem_internal.code_mem[63][3] ;
 wire \mem.mem_internal.code_mem[63][4] ;
 wire \mem.mem_internal.code_mem[63][5] ;
 wire \mem.mem_internal.code_mem[63][6] ;
 wire \mem.mem_internal.code_mem[63][7] ;
 wire \mem.mem_internal.code_mem[64][0] ;
 wire \mem.mem_internal.code_mem[64][1] ;
 wire \mem.mem_internal.code_mem[64][2] ;
 wire \mem.mem_internal.code_mem[64][3] ;
 wire \mem.mem_internal.code_mem[64][4] ;
 wire \mem.mem_internal.code_mem[64][5] ;
 wire \mem.mem_internal.code_mem[64][6] ;
 wire \mem.mem_internal.code_mem[64][7] ;
 wire \mem.mem_internal.code_mem[65][0] ;
 wire \mem.mem_internal.code_mem[65][1] ;
 wire \mem.mem_internal.code_mem[65][2] ;
 wire \mem.mem_internal.code_mem[65][3] ;
 wire \mem.mem_internal.code_mem[65][4] ;
 wire \mem.mem_internal.code_mem[65][5] ;
 wire \mem.mem_internal.code_mem[65][6] ;
 wire \mem.mem_internal.code_mem[65][7] ;
 wire \mem.mem_internal.code_mem[66][0] ;
 wire \mem.mem_internal.code_mem[66][1] ;
 wire \mem.mem_internal.code_mem[66][2] ;
 wire \mem.mem_internal.code_mem[66][3] ;
 wire \mem.mem_internal.code_mem[66][4] ;
 wire \mem.mem_internal.code_mem[66][5] ;
 wire \mem.mem_internal.code_mem[66][6] ;
 wire \mem.mem_internal.code_mem[66][7] ;
 wire \mem.mem_internal.code_mem[67][0] ;
 wire \mem.mem_internal.code_mem[67][1] ;
 wire \mem.mem_internal.code_mem[67][2] ;
 wire \mem.mem_internal.code_mem[67][3] ;
 wire \mem.mem_internal.code_mem[67][4] ;
 wire \mem.mem_internal.code_mem[67][5] ;
 wire \mem.mem_internal.code_mem[67][6] ;
 wire \mem.mem_internal.code_mem[67][7] ;
 wire \mem.mem_internal.code_mem[68][0] ;
 wire \mem.mem_internal.code_mem[68][1] ;
 wire \mem.mem_internal.code_mem[68][2] ;
 wire \mem.mem_internal.code_mem[68][3] ;
 wire \mem.mem_internal.code_mem[68][4] ;
 wire \mem.mem_internal.code_mem[68][5] ;
 wire \mem.mem_internal.code_mem[68][6] ;
 wire \mem.mem_internal.code_mem[68][7] ;
 wire \mem.mem_internal.code_mem[69][0] ;
 wire \mem.mem_internal.code_mem[69][1] ;
 wire \mem.mem_internal.code_mem[69][2] ;
 wire \mem.mem_internal.code_mem[69][3] ;
 wire \mem.mem_internal.code_mem[69][4] ;
 wire \mem.mem_internal.code_mem[69][5] ;
 wire \mem.mem_internal.code_mem[69][6] ;
 wire \mem.mem_internal.code_mem[69][7] ;
 wire \mem.mem_internal.code_mem[6][0] ;
 wire \mem.mem_internal.code_mem[6][1] ;
 wire \mem.mem_internal.code_mem[6][2] ;
 wire \mem.mem_internal.code_mem[6][3] ;
 wire \mem.mem_internal.code_mem[6][4] ;
 wire \mem.mem_internal.code_mem[6][5] ;
 wire \mem.mem_internal.code_mem[6][6] ;
 wire \mem.mem_internal.code_mem[6][7] ;
 wire \mem.mem_internal.code_mem[70][0] ;
 wire \mem.mem_internal.code_mem[70][1] ;
 wire \mem.mem_internal.code_mem[70][2] ;
 wire \mem.mem_internal.code_mem[70][3] ;
 wire \mem.mem_internal.code_mem[70][4] ;
 wire \mem.mem_internal.code_mem[70][5] ;
 wire \mem.mem_internal.code_mem[70][6] ;
 wire \mem.mem_internal.code_mem[70][7] ;
 wire \mem.mem_internal.code_mem[71][0] ;
 wire \mem.mem_internal.code_mem[71][1] ;
 wire \mem.mem_internal.code_mem[71][2] ;
 wire \mem.mem_internal.code_mem[71][3] ;
 wire \mem.mem_internal.code_mem[71][4] ;
 wire \mem.mem_internal.code_mem[71][5] ;
 wire \mem.mem_internal.code_mem[71][6] ;
 wire \mem.mem_internal.code_mem[71][7] ;
 wire \mem.mem_internal.code_mem[72][0] ;
 wire \mem.mem_internal.code_mem[72][1] ;
 wire \mem.mem_internal.code_mem[72][2] ;
 wire \mem.mem_internal.code_mem[72][3] ;
 wire \mem.mem_internal.code_mem[72][4] ;
 wire \mem.mem_internal.code_mem[72][5] ;
 wire \mem.mem_internal.code_mem[72][6] ;
 wire \mem.mem_internal.code_mem[72][7] ;
 wire \mem.mem_internal.code_mem[73][0] ;
 wire \mem.mem_internal.code_mem[73][1] ;
 wire \mem.mem_internal.code_mem[73][2] ;
 wire \mem.mem_internal.code_mem[73][3] ;
 wire \mem.mem_internal.code_mem[73][4] ;
 wire \mem.mem_internal.code_mem[73][5] ;
 wire \mem.mem_internal.code_mem[73][6] ;
 wire \mem.mem_internal.code_mem[73][7] ;
 wire \mem.mem_internal.code_mem[74][0] ;
 wire \mem.mem_internal.code_mem[74][1] ;
 wire \mem.mem_internal.code_mem[74][2] ;
 wire \mem.mem_internal.code_mem[74][3] ;
 wire \mem.mem_internal.code_mem[74][4] ;
 wire \mem.mem_internal.code_mem[74][5] ;
 wire \mem.mem_internal.code_mem[74][6] ;
 wire \mem.mem_internal.code_mem[74][7] ;
 wire \mem.mem_internal.code_mem[75][0] ;
 wire \mem.mem_internal.code_mem[75][1] ;
 wire \mem.mem_internal.code_mem[75][2] ;
 wire \mem.mem_internal.code_mem[75][3] ;
 wire \mem.mem_internal.code_mem[75][4] ;
 wire \mem.mem_internal.code_mem[75][5] ;
 wire \mem.mem_internal.code_mem[75][6] ;
 wire \mem.mem_internal.code_mem[75][7] ;
 wire \mem.mem_internal.code_mem[76][0] ;
 wire \mem.mem_internal.code_mem[76][1] ;
 wire \mem.mem_internal.code_mem[76][2] ;
 wire \mem.mem_internal.code_mem[76][3] ;
 wire \mem.mem_internal.code_mem[76][4] ;
 wire \mem.mem_internal.code_mem[76][5] ;
 wire \mem.mem_internal.code_mem[76][6] ;
 wire \mem.mem_internal.code_mem[76][7] ;
 wire \mem.mem_internal.code_mem[77][0] ;
 wire \mem.mem_internal.code_mem[77][1] ;
 wire \mem.mem_internal.code_mem[77][2] ;
 wire \mem.mem_internal.code_mem[77][3] ;
 wire \mem.mem_internal.code_mem[77][4] ;
 wire \mem.mem_internal.code_mem[77][5] ;
 wire \mem.mem_internal.code_mem[77][6] ;
 wire \mem.mem_internal.code_mem[77][7] ;
 wire \mem.mem_internal.code_mem[78][0] ;
 wire \mem.mem_internal.code_mem[78][1] ;
 wire \mem.mem_internal.code_mem[78][2] ;
 wire \mem.mem_internal.code_mem[78][3] ;
 wire \mem.mem_internal.code_mem[78][4] ;
 wire \mem.mem_internal.code_mem[78][5] ;
 wire \mem.mem_internal.code_mem[78][6] ;
 wire \mem.mem_internal.code_mem[78][7] ;
 wire \mem.mem_internal.code_mem[79][0] ;
 wire \mem.mem_internal.code_mem[79][1] ;
 wire \mem.mem_internal.code_mem[79][2] ;
 wire \mem.mem_internal.code_mem[79][3] ;
 wire \mem.mem_internal.code_mem[79][4] ;
 wire \mem.mem_internal.code_mem[79][5] ;
 wire \mem.mem_internal.code_mem[79][6] ;
 wire \mem.mem_internal.code_mem[79][7] ;
 wire \mem.mem_internal.code_mem[7][0] ;
 wire \mem.mem_internal.code_mem[7][1] ;
 wire \mem.mem_internal.code_mem[7][2] ;
 wire \mem.mem_internal.code_mem[7][3] ;
 wire \mem.mem_internal.code_mem[7][4] ;
 wire \mem.mem_internal.code_mem[7][5] ;
 wire \mem.mem_internal.code_mem[7][6] ;
 wire \mem.mem_internal.code_mem[7][7] ;
 wire \mem.mem_internal.code_mem[80][0] ;
 wire \mem.mem_internal.code_mem[80][1] ;
 wire \mem.mem_internal.code_mem[80][2] ;
 wire \mem.mem_internal.code_mem[80][3] ;
 wire \mem.mem_internal.code_mem[80][4] ;
 wire \mem.mem_internal.code_mem[80][5] ;
 wire \mem.mem_internal.code_mem[80][6] ;
 wire \mem.mem_internal.code_mem[80][7] ;
 wire \mem.mem_internal.code_mem[81][0] ;
 wire \mem.mem_internal.code_mem[81][1] ;
 wire \mem.mem_internal.code_mem[81][2] ;
 wire \mem.mem_internal.code_mem[81][3] ;
 wire \mem.mem_internal.code_mem[81][4] ;
 wire \mem.mem_internal.code_mem[81][5] ;
 wire \mem.mem_internal.code_mem[81][6] ;
 wire \mem.mem_internal.code_mem[81][7] ;
 wire \mem.mem_internal.code_mem[82][0] ;
 wire \mem.mem_internal.code_mem[82][1] ;
 wire \mem.mem_internal.code_mem[82][2] ;
 wire \mem.mem_internal.code_mem[82][3] ;
 wire \mem.mem_internal.code_mem[82][4] ;
 wire \mem.mem_internal.code_mem[82][5] ;
 wire \mem.mem_internal.code_mem[82][6] ;
 wire \mem.mem_internal.code_mem[82][7] ;
 wire \mem.mem_internal.code_mem[83][0] ;
 wire \mem.mem_internal.code_mem[83][1] ;
 wire \mem.mem_internal.code_mem[83][2] ;
 wire \mem.mem_internal.code_mem[83][3] ;
 wire \mem.mem_internal.code_mem[83][4] ;
 wire \mem.mem_internal.code_mem[83][5] ;
 wire \mem.mem_internal.code_mem[83][6] ;
 wire \mem.mem_internal.code_mem[83][7] ;
 wire \mem.mem_internal.code_mem[84][0] ;
 wire \mem.mem_internal.code_mem[84][1] ;
 wire \mem.mem_internal.code_mem[84][2] ;
 wire \mem.mem_internal.code_mem[84][3] ;
 wire \mem.mem_internal.code_mem[84][4] ;
 wire \mem.mem_internal.code_mem[84][5] ;
 wire \mem.mem_internal.code_mem[84][6] ;
 wire \mem.mem_internal.code_mem[84][7] ;
 wire \mem.mem_internal.code_mem[85][0] ;
 wire \mem.mem_internal.code_mem[85][1] ;
 wire \mem.mem_internal.code_mem[85][2] ;
 wire \mem.mem_internal.code_mem[85][3] ;
 wire \mem.mem_internal.code_mem[85][4] ;
 wire \mem.mem_internal.code_mem[85][5] ;
 wire \mem.mem_internal.code_mem[85][6] ;
 wire \mem.mem_internal.code_mem[85][7] ;
 wire \mem.mem_internal.code_mem[86][0] ;
 wire \mem.mem_internal.code_mem[86][1] ;
 wire \mem.mem_internal.code_mem[86][2] ;
 wire \mem.mem_internal.code_mem[86][3] ;
 wire \mem.mem_internal.code_mem[86][4] ;
 wire \mem.mem_internal.code_mem[86][5] ;
 wire \mem.mem_internal.code_mem[86][6] ;
 wire \mem.mem_internal.code_mem[86][7] ;
 wire \mem.mem_internal.code_mem[87][0] ;
 wire \mem.mem_internal.code_mem[87][1] ;
 wire \mem.mem_internal.code_mem[87][2] ;
 wire \mem.mem_internal.code_mem[87][3] ;
 wire \mem.mem_internal.code_mem[87][4] ;
 wire \mem.mem_internal.code_mem[87][5] ;
 wire \mem.mem_internal.code_mem[87][6] ;
 wire \mem.mem_internal.code_mem[87][7] ;
 wire \mem.mem_internal.code_mem[88][0] ;
 wire \mem.mem_internal.code_mem[88][1] ;
 wire \mem.mem_internal.code_mem[88][2] ;
 wire \mem.mem_internal.code_mem[88][3] ;
 wire \mem.mem_internal.code_mem[88][4] ;
 wire \mem.mem_internal.code_mem[88][5] ;
 wire \mem.mem_internal.code_mem[88][6] ;
 wire \mem.mem_internal.code_mem[88][7] ;
 wire \mem.mem_internal.code_mem[89][0] ;
 wire \mem.mem_internal.code_mem[89][1] ;
 wire \mem.mem_internal.code_mem[89][2] ;
 wire \mem.mem_internal.code_mem[89][3] ;
 wire \mem.mem_internal.code_mem[89][4] ;
 wire \mem.mem_internal.code_mem[89][5] ;
 wire \mem.mem_internal.code_mem[89][6] ;
 wire \mem.mem_internal.code_mem[89][7] ;
 wire \mem.mem_internal.code_mem[8][0] ;
 wire \mem.mem_internal.code_mem[8][1] ;
 wire \mem.mem_internal.code_mem[8][2] ;
 wire \mem.mem_internal.code_mem[8][3] ;
 wire \mem.mem_internal.code_mem[8][4] ;
 wire \mem.mem_internal.code_mem[8][5] ;
 wire \mem.mem_internal.code_mem[8][6] ;
 wire \mem.mem_internal.code_mem[8][7] ;
 wire \mem.mem_internal.code_mem[90][0] ;
 wire \mem.mem_internal.code_mem[90][1] ;
 wire \mem.mem_internal.code_mem[90][2] ;
 wire \mem.mem_internal.code_mem[90][3] ;
 wire \mem.mem_internal.code_mem[90][4] ;
 wire \mem.mem_internal.code_mem[90][5] ;
 wire \mem.mem_internal.code_mem[90][6] ;
 wire \mem.mem_internal.code_mem[90][7] ;
 wire \mem.mem_internal.code_mem[91][0] ;
 wire \mem.mem_internal.code_mem[91][1] ;
 wire \mem.mem_internal.code_mem[91][2] ;
 wire \mem.mem_internal.code_mem[91][3] ;
 wire \mem.mem_internal.code_mem[91][4] ;
 wire \mem.mem_internal.code_mem[91][5] ;
 wire \mem.mem_internal.code_mem[91][6] ;
 wire \mem.mem_internal.code_mem[91][7] ;
 wire \mem.mem_internal.code_mem[92][0] ;
 wire \mem.mem_internal.code_mem[92][1] ;
 wire \mem.mem_internal.code_mem[92][2] ;
 wire \mem.mem_internal.code_mem[92][3] ;
 wire \mem.mem_internal.code_mem[92][4] ;
 wire \mem.mem_internal.code_mem[92][5] ;
 wire \mem.mem_internal.code_mem[92][6] ;
 wire \mem.mem_internal.code_mem[92][7] ;
 wire \mem.mem_internal.code_mem[93][0] ;
 wire \mem.mem_internal.code_mem[93][1] ;
 wire \mem.mem_internal.code_mem[93][2] ;
 wire \mem.mem_internal.code_mem[93][3] ;
 wire \mem.mem_internal.code_mem[93][4] ;
 wire \mem.mem_internal.code_mem[93][5] ;
 wire \mem.mem_internal.code_mem[93][6] ;
 wire \mem.mem_internal.code_mem[93][7] ;
 wire \mem.mem_internal.code_mem[94][0] ;
 wire \mem.mem_internal.code_mem[94][1] ;
 wire \mem.mem_internal.code_mem[94][2] ;
 wire \mem.mem_internal.code_mem[94][3] ;
 wire \mem.mem_internal.code_mem[94][4] ;
 wire \mem.mem_internal.code_mem[94][5] ;
 wire \mem.mem_internal.code_mem[94][6] ;
 wire \mem.mem_internal.code_mem[94][7] ;
 wire \mem.mem_internal.code_mem[95][0] ;
 wire \mem.mem_internal.code_mem[95][1] ;
 wire \mem.mem_internal.code_mem[95][2] ;
 wire \mem.mem_internal.code_mem[95][3] ;
 wire \mem.mem_internal.code_mem[95][4] ;
 wire \mem.mem_internal.code_mem[95][5] ;
 wire \mem.mem_internal.code_mem[95][6] ;
 wire \mem.mem_internal.code_mem[95][7] ;
 wire \mem.mem_internal.code_mem[96][0] ;
 wire \mem.mem_internal.code_mem[96][1] ;
 wire \mem.mem_internal.code_mem[96][2] ;
 wire \mem.mem_internal.code_mem[96][3] ;
 wire \mem.mem_internal.code_mem[96][4] ;
 wire \mem.mem_internal.code_mem[96][5] ;
 wire \mem.mem_internal.code_mem[96][6] ;
 wire \mem.mem_internal.code_mem[96][7] ;
 wire \mem.mem_internal.code_mem[97][0] ;
 wire \mem.mem_internal.code_mem[97][1] ;
 wire \mem.mem_internal.code_mem[97][2] ;
 wire \mem.mem_internal.code_mem[97][3] ;
 wire \mem.mem_internal.code_mem[97][4] ;
 wire \mem.mem_internal.code_mem[97][5] ;
 wire \mem.mem_internal.code_mem[97][6] ;
 wire \mem.mem_internal.code_mem[97][7] ;
 wire \mem.mem_internal.code_mem[98][0] ;
 wire \mem.mem_internal.code_mem[98][1] ;
 wire \mem.mem_internal.code_mem[98][2] ;
 wire \mem.mem_internal.code_mem[98][3] ;
 wire \mem.mem_internal.code_mem[98][4] ;
 wire \mem.mem_internal.code_mem[98][5] ;
 wire \mem.mem_internal.code_mem[98][6] ;
 wire \mem.mem_internal.code_mem[98][7] ;
 wire \mem.mem_internal.code_mem[99][0] ;
 wire \mem.mem_internal.code_mem[99][1] ;
 wire \mem.mem_internal.code_mem[99][2] ;
 wire \mem.mem_internal.code_mem[99][3] ;
 wire \mem.mem_internal.code_mem[99][4] ;
 wire \mem.mem_internal.code_mem[99][5] ;
 wire \mem.mem_internal.code_mem[99][6] ;
 wire \mem.mem_internal.code_mem[99][7] ;
 wire \mem.mem_internal.code_mem[9][0] ;
 wire \mem.mem_internal.code_mem[9][1] ;
 wire \mem.mem_internal.code_mem[9][2] ;
 wire \mem.mem_internal.code_mem[9][3] ;
 wire \mem.mem_internal.code_mem[9][4] ;
 wire \mem.mem_internal.code_mem[9][5] ;
 wire \mem.mem_internal.code_mem[9][6] ;
 wire \mem.mem_internal.code_mem[9][7] ;
 wire \mem.mem_internal.cycles[0] ;
 wire \mem.mem_internal.cycles[1] ;
 wire \mem.mem_internal.data_mem[0][0] ;
 wire \mem.mem_internal.data_mem[0][1] ;
 wire \mem.mem_internal.data_mem[0][2] ;
 wire \mem.mem_internal.data_mem[0][3] ;
 wire \mem.mem_internal.data_mem[0][4] ;
 wire \mem.mem_internal.data_mem[0][5] ;
 wire \mem.mem_internal.data_mem[0][6] ;
 wire \mem.mem_internal.data_mem[0][7] ;
 wire \mem.mem_internal.data_mem[10][0] ;
 wire \mem.mem_internal.data_mem[10][1] ;
 wire \mem.mem_internal.data_mem[10][2] ;
 wire \mem.mem_internal.data_mem[10][3] ;
 wire \mem.mem_internal.data_mem[10][4] ;
 wire \mem.mem_internal.data_mem[10][5] ;
 wire \mem.mem_internal.data_mem[10][6] ;
 wire \mem.mem_internal.data_mem[10][7] ;
 wire \mem.mem_internal.data_mem[11][0] ;
 wire \mem.mem_internal.data_mem[11][1] ;
 wire \mem.mem_internal.data_mem[11][2] ;
 wire \mem.mem_internal.data_mem[11][3] ;
 wire \mem.mem_internal.data_mem[11][4] ;
 wire \mem.mem_internal.data_mem[11][5] ;
 wire \mem.mem_internal.data_mem[11][6] ;
 wire \mem.mem_internal.data_mem[11][7] ;
 wire \mem.mem_internal.data_mem[12][0] ;
 wire \mem.mem_internal.data_mem[12][1] ;
 wire \mem.mem_internal.data_mem[12][2] ;
 wire \mem.mem_internal.data_mem[12][3] ;
 wire \mem.mem_internal.data_mem[12][4] ;
 wire \mem.mem_internal.data_mem[12][5] ;
 wire \mem.mem_internal.data_mem[12][6] ;
 wire \mem.mem_internal.data_mem[12][7] ;
 wire \mem.mem_internal.data_mem[13][0] ;
 wire \mem.mem_internal.data_mem[13][1] ;
 wire \mem.mem_internal.data_mem[13][2] ;
 wire \mem.mem_internal.data_mem[13][3] ;
 wire \mem.mem_internal.data_mem[13][4] ;
 wire \mem.mem_internal.data_mem[13][5] ;
 wire \mem.mem_internal.data_mem[13][6] ;
 wire \mem.mem_internal.data_mem[13][7] ;
 wire \mem.mem_internal.data_mem[14][0] ;
 wire \mem.mem_internal.data_mem[14][1] ;
 wire \mem.mem_internal.data_mem[14][2] ;
 wire \mem.mem_internal.data_mem[14][3] ;
 wire \mem.mem_internal.data_mem[14][4] ;
 wire \mem.mem_internal.data_mem[14][5] ;
 wire \mem.mem_internal.data_mem[14][6] ;
 wire \mem.mem_internal.data_mem[14][7] ;
 wire \mem.mem_internal.data_mem[15][0] ;
 wire \mem.mem_internal.data_mem[15][1] ;
 wire \mem.mem_internal.data_mem[15][2] ;
 wire \mem.mem_internal.data_mem[15][3] ;
 wire \mem.mem_internal.data_mem[15][4] ;
 wire \mem.mem_internal.data_mem[15][5] ;
 wire \mem.mem_internal.data_mem[15][6] ;
 wire \mem.mem_internal.data_mem[15][7] ;
 wire \mem.mem_internal.data_mem[16][0] ;
 wire \mem.mem_internal.data_mem[16][1] ;
 wire \mem.mem_internal.data_mem[16][2] ;
 wire \mem.mem_internal.data_mem[16][3] ;
 wire \mem.mem_internal.data_mem[16][4] ;
 wire \mem.mem_internal.data_mem[16][5] ;
 wire \mem.mem_internal.data_mem[16][6] ;
 wire \mem.mem_internal.data_mem[16][7] ;
 wire \mem.mem_internal.data_mem[17][0] ;
 wire \mem.mem_internal.data_mem[17][1] ;
 wire \mem.mem_internal.data_mem[17][2] ;
 wire \mem.mem_internal.data_mem[17][3] ;
 wire \mem.mem_internal.data_mem[17][4] ;
 wire \mem.mem_internal.data_mem[17][5] ;
 wire \mem.mem_internal.data_mem[17][6] ;
 wire \mem.mem_internal.data_mem[17][7] ;
 wire \mem.mem_internal.data_mem[18][0] ;
 wire \mem.mem_internal.data_mem[18][1] ;
 wire \mem.mem_internal.data_mem[18][2] ;
 wire \mem.mem_internal.data_mem[18][3] ;
 wire \mem.mem_internal.data_mem[18][4] ;
 wire \mem.mem_internal.data_mem[18][5] ;
 wire \mem.mem_internal.data_mem[18][6] ;
 wire \mem.mem_internal.data_mem[18][7] ;
 wire \mem.mem_internal.data_mem[19][0] ;
 wire \mem.mem_internal.data_mem[19][1] ;
 wire \mem.mem_internal.data_mem[19][2] ;
 wire \mem.mem_internal.data_mem[19][3] ;
 wire \mem.mem_internal.data_mem[19][4] ;
 wire \mem.mem_internal.data_mem[19][5] ;
 wire \mem.mem_internal.data_mem[19][6] ;
 wire \mem.mem_internal.data_mem[19][7] ;
 wire \mem.mem_internal.data_mem[1][0] ;
 wire \mem.mem_internal.data_mem[1][1] ;
 wire \mem.mem_internal.data_mem[1][2] ;
 wire \mem.mem_internal.data_mem[1][3] ;
 wire \mem.mem_internal.data_mem[1][4] ;
 wire \mem.mem_internal.data_mem[1][5] ;
 wire \mem.mem_internal.data_mem[1][6] ;
 wire \mem.mem_internal.data_mem[1][7] ;
 wire \mem.mem_internal.data_mem[20][0] ;
 wire \mem.mem_internal.data_mem[20][1] ;
 wire \mem.mem_internal.data_mem[20][2] ;
 wire \mem.mem_internal.data_mem[20][3] ;
 wire \mem.mem_internal.data_mem[20][4] ;
 wire \mem.mem_internal.data_mem[20][5] ;
 wire \mem.mem_internal.data_mem[20][6] ;
 wire \mem.mem_internal.data_mem[20][7] ;
 wire \mem.mem_internal.data_mem[21][0] ;
 wire \mem.mem_internal.data_mem[21][1] ;
 wire \mem.mem_internal.data_mem[21][2] ;
 wire \mem.mem_internal.data_mem[21][3] ;
 wire \mem.mem_internal.data_mem[21][4] ;
 wire \mem.mem_internal.data_mem[21][5] ;
 wire \mem.mem_internal.data_mem[21][6] ;
 wire \mem.mem_internal.data_mem[21][7] ;
 wire \mem.mem_internal.data_mem[22][0] ;
 wire \mem.mem_internal.data_mem[22][1] ;
 wire \mem.mem_internal.data_mem[22][2] ;
 wire \mem.mem_internal.data_mem[22][3] ;
 wire \mem.mem_internal.data_mem[22][4] ;
 wire \mem.mem_internal.data_mem[22][5] ;
 wire \mem.mem_internal.data_mem[22][6] ;
 wire \mem.mem_internal.data_mem[22][7] ;
 wire \mem.mem_internal.data_mem[23][0] ;
 wire \mem.mem_internal.data_mem[23][1] ;
 wire \mem.mem_internal.data_mem[23][2] ;
 wire \mem.mem_internal.data_mem[23][3] ;
 wire \mem.mem_internal.data_mem[23][4] ;
 wire \mem.mem_internal.data_mem[23][5] ;
 wire \mem.mem_internal.data_mem[23][6] ;
 wire \mem.mem_internal.data_mem[23][7] ;
 wire \mem.mem_internal.data_mem[24][0] ;
 wire \mem.mem_internal.data_mem[24][1] ;
 wire \mem.mem_internal.data_mem[24][2] ;
 wire \mem.mem_internal.data_mem[24][3] ;
 wire \mem.mem_internal.data_mem[24][4] ;
 wire \mem.mem_internal.data_mem[24][5] ;
 wire \mem.mem_internal.data_mem[24][6] ;
 wire \mem.mem_internal.data_mem[24][7] ;
 wire \mem.mem_internal.data_mem[25][0] ;
 wire \mem.mem_internal.data_mem[25][1] ;
 wire \mem.mem_internal.data_mem[25][2] ;
 wire \mem.mem_internal.data_mem[25][3] ;
 wire \mem.mem_internal.data_mem[25][4] ;
 wire \mem.mem_internal.data_mem[25][5] ;
 wire \mem.mem_internal.data_mem[25][6] ;
 wire \mem.mem_internal.data_mem[25][7] ;
 wire \mem.mem_internal.data_mem[26][0] ;
 wire \mem.mem_internal.data_mem[26][1] ;
 wire \mem.mem_internal.data_mem[26][2] ;
 wire \mem.mem_internal.data_mem[26][3] ;
 wire \mem.mem_internal.data_mem[26][4] ;
 wire \mem.mem_internal.data_mem[26][5] ;
 wire \mem.mem_internal.data_mem[26][6] ;
 wire \mem.mem_internal.data_mem[26][7] ;
 wire \mem.mem_internal.data_mem[27][0] ;
 wire \mem.mem_internal.data_mem[27][1] ;
 wire \mem.mem_internal.data_mem[27][2] ;
 wire \mem.mem_internal.data_mem[27][3] ;
 wire \mem.mem_internal.data_mem[27][4] ;
 wire \mem.mem_internal.data_mem[27][5] ;
 wire \mem.mem_internal.data_mem[27][6] ;
 wire \mem.mem_internal.data_mem[27][7] ;
 wire \mem.mem_internal.data_mem[28][0] ;
 wire \mem.mem_internal.data_mem[28][1] ;
 wire \mem.mem_internal.data_mem[28][2] ;
 wire \mem.mem_internal.data_mem[28][3] ;
 wire \mem.mem_internal.data_mem[28][4] ;
 wire \mem.mem_internal.data_mem[28][5] ;
 wire \mem.mem_internal.data_mem[28][6] ;
 wire \mem.mem_internal.data_mem[28][7] ;
 wire \mem.mem_internal.data_mem[29][0] ;
 wire \mem.mem_internal.data_mem[29][1] ;
 wire \mem.mem_internal.data_mem[29][2] ;
 wire \mem.mem_internal.data_mem[29][3] ;
 wire \mem.mem_internal.data_mem[29][4] ;
 wire \mem.mem_internal.data_mem[29][5] ;
 wire \mem.mem_internal.data_mem[29][6] ;
 wire \mem.mem_internal.data_mem[29][7] ;
 wire \mem.mem_internal.data_mem[2][0] ;
 wire \mem.mem_internal.data_mem[2][1] ;
 wire \mem.mem_internal.data_mem[2][2] ;
 wire \mem.mem_internal.data_mem[2][3] ;
 wire \mem.mem_internal.data_mem[2][4] ;
 wire \mem.mem_internal.data_mem[2][5] ;
 wire \mem.mem_internal.data_mem[2][6] ;
 wire \mem.mem_internal.data_mem[2][7] ;
 wire \mem.mem_internal.data_mem[30][0] ;
 wire \mem.mem_internal.data_mem[30][1] ;
 wire \mem.mem_internal.data_mem[30][2] ;
 wire \mem.mem_internal.data_mem[30][3] ;
 wire \mem.mem_internal.data_mem[30][4] ;
 wire \mem.mem_internal.data_mem[30][5] ;
 wire \mem.mem_internal.data_mem[30][6] ;
 wire \mem.mem_internal.data_mem[30][7] ;
 wire \mem.mem_internal.data_mem[31][0] ;
 wire \mem.mem_internal.data_mem[31][1] ;
 wire \mem.mem_internal.data_mem[31][2] ;
 wire \mem.mem_internal.data_mem[31][3] ;
 wire \mem.mem_internal.data_mem[31][4] ;
 wire \mem.mem_internal.data_mem[31][5] ;
 wire \mem.mem_internal.data_mem[31][6] ;
 wire \mem.mem_internal.data_mem[31][7] ;
 wire \mem.mem_internal.data_mem[3][0] ;
 wire \mem.mem_internal.data_mem[3][1] ;
 wire \mem.mem_internal.data_mem[3][2] ;
 wire \mem.mem_internal.data_mem[3][3] ;
 wire \mem.mem_internal.data_mem[3][4] ;
 wire \mem.mem_internal.data_mem[3][5] ;
 wire \mem.mem_internal.data_mem[3][6] ;
 wire \mem.mem_internal.data_mem[3][7] ;
 wire \mem.mem_internal.data_mem[4][0] ;
 wire \mem.mem_internal.data_mem[4][1] ;
 wire \mem.mem_internal.data_mem[4][2] ;
 wire \mem.mem_internal.data_mem[4][3] ;
 wire \mem.mem_internal.data_mem[4][4] ;
 wire \mem.mem_internal.data_mem[4][5] ;
 wire \mem.mem_internal.data_mem[4][6] ;
 wire \mem.mem_internal.data_mem[4][7] ;
 wire \mem.mem_internal.data_mem[5][0] ;
 wire \mem.mem_internal.data_mem[5][1] ;
 wire \mem.mem_internal.data_mem[5][2] ;
 wire \mem.mem_internal.data_mem[5][3] ;
 wire \mem.mem_internal.data_mem[5][4] ;
 wire \mem.mem_internal.data_mem[5][5] ;
 wire \mem.mem_internal.data_mem[5][6] ;
 wire \mem.mem_internal.data_mem[5][7] ;
 wire \mem.mem_internal.data_mem[6][0] ;
 wire \mem.mem_internal.data_mem[6][1] ;
 wire \mem.mem_internal.data_mem[6][2] ;
 wire \mem.mem_internal.data_mem[6][3] ;
 wire \mem.mem_internal.data_mem[6][4] ;
 wire \mem.mem_internal.data_mem[6][5] ;
 wire \mem.mem_internal.data_mem[6][6] ;
 wire \mem.mem_internal.data_mem[6][7] ;
 wire \mem.mem_internal.data_mem[7][0] ;
 wire \mem.mem_internal.data_mem[7][1] ;
 wire \mem.mem_internal.data_mem[7][2] ;
 wire \mem.mem_internal.data_mem[7][3] ;
 wire \mem.mem_internal.data_mem[7][4] ;
 wire \mem.mem_internal.data_mem[7][5] ;
 wire \mem.mem_internal.data_mem[7][6] ;
 wire \mem.mem_internal.data_mem[7][7] ;
 wire \mem.mem_internal.data_mem[8][0] ;
 wire \mem.mem_internal.data_mem[8][1] ;
 wire \mem.mem_internal.data_mem[8][2] ;
 wire \mem.mem_internal.data_mem[8][3] ;
 wire \mem.mem_internal.data_mem[8][4] ;
 wire \mem.mem_internal.data_mem[8][5] ;
 wire \mem.mem_internal.data_mem[8][6] ;
 wire \mem.mem_internal.data_mem[8][7] ;
 wire \mem.mem_internal.data_mem[9][0] ;
 wire \mem.mem_internal.data_mem[9][1] ;
 wire \mem.mem_internal.data_mem[9][2] ;
 wire \mem.mem_internal.data_mem[9][3] ;
 wire \mem.mem_internal.data_mem[9][4] ;
 wire \mem.mem_internal.data_mem[9][5] ;
 wire \mem.mem_internal.data_mem[9][6] ;
 wire \mem.mem_internal.data_mem[9][7] ;
 wire \mem.mem_internal.memory_type_data ;
 wire \mem.mem_internal.write ;
 wire \mem.mem_io.past_write ;
 wire \mem.mem_io.porta_oe[0] ;
 wire \mem.mem_io.porta_oe[1] ;
 wire \mem.mem_io.porta_oe[2] ;
 wire \mem.mem_io.porta_oe[3] ;
 wire \mem.mem_io.porta_oe[4] ;
 wire \mem.mem_io.porta_oe[5] ;
 wire \mem.mem_io.porta_oe[6] ;
 wire \mem.mem_io.porta_oe[7] ;
 wire \mem.mem_io.porta_out[0] ;
 wire \mem.mem_io.porta_out[1] ;
 wire \mem.mem_io.porta_out[2] ;
 wire \mem.mem_io.porta_out[3] ;
 wire \mem.mem_io.porta_out[4] ;
 wire \mem.mem_io.porta_out[5] ;
 wire \mem.mem_io.porta_out[6] ;
 wire \mem.mem_io.porta_out[7] ;
 wire \mem.select ;
 wire o_shift_out;
 wire o_sleep;
 wire o_wait_delay;
 wire past_i_run;
 wire \shift_reg[0] ;
 wire \shift_reg[1] ;
 wire \shift_reg[2] ;
 wire \shift_reg[3] ;
 wire \shift_reg[4] ;
 wire \shift_reg[5] ;
 wire \shift_reg[6] ;
 wire \shift_reg[7] ;
 wire single_step;
 wire \stack[0][0] ;
 wire \stack[0][1] ;
 wire \stack[0][2] ;
 wire \stack[0][3] ;
 wire \stack[0][4] ;
 wire \stack[0][5] ;
 wire \stack[0][6] ;
 wire \stack[0][7] ;
 wire \stack[10][0] ;
 wire \stack[10][1] ;
 wire \stack[10][2] ;
 wire \stack[10][3] ;
 wire \stack[10][4] ;
 wire \stack[10][5] ;
 wire \stack[10][6] ;
 wire \stack[10][7] ;
 wire \stack[11][0] ;
 wire \stack[11][1] ;
 wire \stack[11][2] ;
 wire \stack[11][3] ;
 wire \stack[11][4] ;
 wire \stack[11][5] ;
 wire \stack[11][6] ;
 wire \stack[11][7] ;
 wire \stack[12][0] ;
 wire \stack[12][1] ;
 wire \stack[12][2] ;
 wire \stack[12][3] ;
 wire \stack[12][4] ;
 wire \stack[12][5] ;
 wire \stack[12][6] ;
 wire \stack[12][7] ;
 wire \stack[13][0] ;
 wire \stack[13][1] ;
 wire \stack[13][2] ;
 wire \stack[13][3] ;
 wire \stack[13][4] ;
 wire \stack[13][5] ;
 wire \stack[13][6] ;
 wire \stack[13][7] ;
 wire \stack[14][0] ;
 wire \stack[14][1] ;
 wire \stack[14][2] ;
 wire \stack[14][3] ;
 wire \stack[14][4] ;
 wire \stack[14][5] ;
 wire \stack[14][6] ;
 wire \stack[14][7] ;
 wire \stack[15][0] ;
 wire \stack[15][1] ;
 wire \stack[15][2] ;
 wire \stack[15][3] ;
 wire \stack[15][4] ;
 wire \stack[15][5] ;
 wire \stack[15][6] ;
 wire \stack[15][7] ;
 wire \stack[16][0] ;
 wire \stack[16][1] ;
 wire \stack[16][2] ;
 wire \stack[16][3] ;
 wire \stack[16][4] ;
 wire \stack[16][5] ;
 wire \stack[16][6] ;
 wire \stack[16][7] ;
 wire \stack[17][0] ;
 wire \stack[17][1] ;
 wire \stack[17][2] ;
 wire \stack[17][3] ;
 wire \stack[17][4] ;
 wire \stack[17][5] ;
 wire \stack[17][6] ;
 wire \stack[17][7] ;
 wire \stack[18][0] ;
 wire \stack[18][1] ;
 wire \stack[18][2] ;
 wire \stack[18][3] ;
 wire \stack[18][4] ;
 wire \stack[18][5] ;
 wire \stack[18][6] ;
 wire \stack[18][7] ;
 wire \stack[19][0] ;
 wire \stack[19][1] ;
 wire \stack[19][2] ;
 wire \stack[19][3] ;
 wire \stack[19][4] ;
 wire \stack[19][5] ;
 wire \stack[19][6] ;
 wire \stack[19][7] ;
 wire \stack[1][0] ;
 wire \stack[1][1] ;
 wire \stack[1][2] ;
 wire \stack[1][3] ;
 wire \stack[1][4] ;
 wire \stack[1][5] ;
 wire \stack[1][6] ;
 wire \stack[1][7] ;
 wire \stack[20][0] ;
 wire \stack[20][1] ;
 wire \stack[20][2] ;
 wire \stack[20][3] ;
 wire \stack[20][4] ;
 wire \stack[20][5] ;
 wire \stack[20][6] ;
 wire \stack[20][7] ;
 wire \stack[21][0] ;
 wire \stack[21][1] ;
 wire \stack[21][2] ;
 wire \stack[21][3] ;
 wire \stack[21][4] ;
 wire \stack[21][5] ;
 wire \stack[21][6] ;
 wire \stack[21][7] ;
 wire \stack[22][0] ;
 wire \stack[22][1] ;
 wire \stack[22][2] ;
 wire \stack[22][3] ;
 wire \stack[22][4] ;
 wire \stack[22][5] ;
 wire \stack[22][6] ;
 wire \stack[22][7] ;
 wire \stack[23][0] ;
 wire \stack[23][1] ;
 wire \stack[23][2] ;
 wire \stack[23][3] ;
 wire \stack[23][4] ;
 wire \stack[23][5] ;
 wire \stack[23][6] ;
 wire \stack[23][7] ;
 wire \stack[24][0] ;
 wire \stack[24][1] ;
 wire \stack[24][2] ;
 wire \stack[24][3] ;
 wire \stack[24][4] ;
 wire \stack[24][5] ;
 wire \stack[24][6] ;
 wire \stack[24][7] ;
 wire \stack[25][0] ;
 wire \stack[25][1] ;
 wire \stack[25][2] ;
 wire \stack[25][3] ;
 wire \stack[25][4] ;
 wire \stack[25][5] ;
 wire \stack[25][6] ;
 wire \stack[25][7] ;
 wire \stack[26][0] ;
 wire \stack[26][1] ;
 wire \stack[26][2] ;
 wire \stack[26][3] ;
 wire \stack[26][4] ;
 wire \stack[26][5] ;
 wire \stack[26][6] ;
 wire \stack[26][7] ;
 wire \stack[27][0] ;
 wire \stack[27][1] ;
 wire \stack[27][2] ;
 wire \stack[27][3] ;
 wire \stack[27][4] ;
 wire \stack[27][5] ;
 wire \stack[27][6] ;
 wire \stack[27][7] ;
 wire \stack[28][0] ;
 wire \stack[28][1] ;
 wire \stack[28][2] ;
 wire \stack[28][3] ;
 wire \stack[28][4] ;
 wire \stack[28][5] ;
 wire \stack[28][6] ;
 wire \stack[28][7] ;
 wire \stack[29][0] ;
 wire \stack[29][1] ;
 wire \stack[29][2] ;
 wire \stack[29][3] ;
 wire \stack[29][4] ;
 wire \stack[29][5] ;
 wire \stack[29][6] ;
 wire \stack[29][7] ;
 wire \stack[2][0] ;
 wire \stack[2][1] ;
 wire \stack[2][2] ;
 wire \stack[2][3] ;
 wire \stack[2][4] ;
 wire \stack[2][5] ;
 wire \stack[2][6] ;
 wire \stack[2][7] ;
 wire \stack[30][0] ;
 wire \stack[30][1] ;
 wire \stack[30][2] ;
 wire \stack[30][3] ;
 wire \stack[30][4] ;
 wire \stack[30][5] ;
 wire \stack[30][6] ;
 wire \stack[30][7] ;
 wire \stack[31][0] ;
 wire \stack[31][1] ;
 wire \stack[31][2] ;
 wire \stack[31][3] ;
 wire \stack[31][4] ;
 wire \stack[31][5] ;
 wire \stack[31][6] ;
 wire \stack[31][7] ;
 wire \stack[3][0] ;
 wire \stack[3][1] ;
 wire \stack[3][2] ;
 wire \stack[3][3] ;
 wire \stack[3][4] ;
 wire \stack[3][5] ;
 wire \stack[3][6] ;
 wire \stack[3][7] ;
 wire \stack[4][0] ;
 wire \stack[4][1] ;
 wire \stack[4][2] ;
 wire \stack[4][3] ;
 wire \stack[4][4] ;
 wire \stack[4][5] ;
 wire \stack[4][6] ;
 wire \stack[4][7] ;
 wire \stack[5][0] ;
 wire \stack[5][1] ;
 wire \stack[5][2] ;
 wire \stack[5][3] ;
 wire \stack[5][4] ;
 wire \stack[5][5] ;
 wire \stack[5][6] ;
 wire \stack[5][7] ;
 wire \stack[6][0] ;
 wire \stack[6][1] ;
 wire \stack[6][2] ;
 wire \stack[6][3] ;
 wire \stack[6][4] ;
 wire \stack[6][5] ;
 wire \stack[6][6] ;
 wire \stack[6][7] ;
 wire \stack[7][0] ;
 wire \stack[7][1] ;
 wire \stack[7][2] ;
 wire \stack[7][3] ;
 wire \stack[7][4] ;
 wire \stack[7][5] ;
 wire \stack[7][6] ;
 wire \stack[7][7] ;
 wire \stack[8][0] ;
 wire \stack[8][1] ;
 wire \stack[8][2] ;
 wire \stack[8][3] ;
 wire \stack[8][4] ;
 wire \stack[8][5] ;
 wire \stack[8][6] ;
 wire \stack[8][7] ;
 wire \stack[9][0] ;
 wire \stack[9][1] ;
 wire \stack[9][2] ;
 wire \stack[9][3] ;
 wire \stack[9][4] ;
 wire \stack[9][5] ;
 wire \stack[9][6] ;
 wire \stack[9][7] ;
 wire \state[1] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_leaf_326_clk;
 wire clknet_leaf_327_clk;
 wire clknet_leaf_328_clk;
 wire clknet_leaf_329_clk;
 wire clknet_leaf_330_clk;
 wire clknet_leaf_331_clk;
 wire clknet_leaf_332_clk;
 wire clknet_leaf_333_clk;
 wire clknet_leaf_334_clk;
 wire clknet_leaf_335_clk;
 wire clknet_leaf_336_clk;
 wire clknet_leaf_337_clk;
 wire clknet_leaf_338_clk;
 wire clknet_leaf_339_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_8 _15705_ (.A(\exec.sp[0] ),
    .X(_09614_));
 sg13g2_buf_8 _15706_ (.A(_09614_),
    .X(_09615_));
 sg13g2_buf_8 _15707_ (.A(_09615_),
    .X(_09616_));
 sg13g2_buf_8 _15708_ (.A(net1206),
    .X(_09617_));
 sg13g2_buf_8 _15709_ (.A(net874),
    .X(_09618_));
 sg13g2_buf_8 _15710_ (.A(net788),
    .X(_09619_));
 sg13g2_buf_2 _15711_ (.A(net565),
    .X(_09620_));
 sg13g2_buf_8 _15712_ (.A(\exec.sp[1] ),
    .X(_09621_));
 sg13g2_buf_8 _15713_ (.A(net1311),
    .X(_09622_));
 sg13g2_buf_8 _15714_ (.A(net1281),
    .X(_09623_));
 sg13g2_buf_1 _15715_ (.A(net1205),
    .X(_09624_));
 sg13g2_buf_8 _15716_ (.A(net873),
    .X(_09625_));
 sg13g2_buf_1 _15717_ (.A(net787),
    .X(_09626_));
 sg13g2_buf_1 _15718_ (.A(net564),
    .X(_09627_));
 sg13g2_mux4_1 _15719_ (.S0(_09620_),
    .A0(\stack[27][7] ),
    .A1(\stack[24][7] ),
    .A2(\stack[25][7] ),
    .A3(\stack[26][7] ),
    .S1(net530),
    .X(_09628_));
 sg13g2_mux4_1 _15720_ (.S0(_09620_),
    .A0(\stack[19][7] ),
    .A1(\stack[16][7] ),
    .A2(\stack[17][7] ),
    .A3(\stack[18][7] ),
    .S1(net530),
    .X(_09629_));
 sg13g2_mux4_1 _15721_ (.S0(_09619_),
    .A0(\stack[31][7] ),
    .A1(\stack[28][7] ),
    .A2(\stack[29][7] ),
    .A3(\stack[30][7] ),
    .S1(_09627_),
    .X(_09630_));
 sg13g2_mux4_1 _15722_ (.S0(net565),
    .A0(\stack[23][7] ),
    .A1(\stack[20][7] ),
    .A2(\stack[21][7] ),
    .A3(\stack[22][7] ),
    .S1(_09627_),
    .X(_09631_));
 sg13g2_buf_2 _15723_ (.A(_00039_),
    .X(_09632_));
 sg13g2_inv_2 _15724_ (.Y(_09633_),
    .A(_09632_));
 sg13g2_buf_1 _15725_ (.A(\exec.sp[2] ),
    .X(_09634_));
 sg13g2_nor3_2 _15726_ (.A(net1282),
    .B(net1311),
    .C(net1310),
    .Y(_09635_));
 sg13g2_xnor2_1 _15727_ (.Y(_09636_),
    .A(_09633_),
    .B(_09635_));
 sg13g2_buf_1 _15728_ (.A(_09636_),
    .X(_09637_));
 sg13g2_buf_2 _15729_ (.A(_09637_),
    .X(_09638_));
 sg13g2_or3_1 _15730_ (.A(_09614_),
    .B(\exec.sp[1] ),
    .C(net1310),
    .X(_09639_));
 sg13g2_buf_1 _15731_ (.A(_09639_),
    .X(_09640_));
 sg13g2_o21ai_1 _15732_ (.B1(net1310),
    .Y(_09641_),
    .A1(_09614_),
    .A2(net1311));
 sg13g2_buf_2 _15733_ (.A(_09641_),
    .X(_09642_));
 sg13g2_nand2_1 _15734_ (.Y(_09643_),
    .A(_09640_),
    .B(_09642_));
 sg13g2_buf_2 _15735_ (.A(_09643_),
    .X(_09644_));
 sg13g2_buf_8 _15736_ (.A(_09644_),
    .X(_09645_));
 sg13g2_mux4_1 _15737_ (.S0(_09638_),
    .A0(_09628_),
    .A1(_09629_),
    .A2(_09630_),
    .A3(_09631_),
    .S1(_09645_),
    .X(_09646_));
 sg13g2_mux4_1 _15738_ (.S0(net565),
    .A0(\stack[11][7] ),
    .A1(\stack[8][7] ),
    .A2(\stack[9][7] ),
    .A3(\stack[10][7] ),
    .S1(net530),
    .X(_09647_));
 sg13g2_mux4_1 _15739_ (.S0(net531),
    .A0(\stack[3][7] ),
    .A1(\stack[0][7] ),
    .A2(\stack[1][7] ),
    .A3(\stack[2][7] ),
    .S1(net530),
    .X(_09648_));
 sg13g2_mux4_1 _15740_ (.S0(net565),
    .A0(\stack[15][7] ),
    .A1(\stack[12][7] ),
    .A2(\stack[13][7] ),
    .A3(\stack[14][7] ),
    .S1(net530),
    .X(_09649_));
 sg13g2_mux4_1 _15741_ (.S0(net565),
    .A0(\stack[7][7] ),
    .A1(\stack[4][7] ),
    .A2(\stack[5][7] ),
    .A3(\stack[6][7] ),
    .S1(net530),
    .X(_09650_));
 sg13g2_mux4_1 _15742_ (.S0(net563),
    .A0(_09647_),
    .A1(_09648_),
    .A2(_09649_),
    .A3(_09650_),
    .S1(net562),
    .X(_09651_));
 sg13g2_buf_8 _15743_ (.A(_00048_),
    .X(_09652_));
 sg13g2_inv_1 _15744_ (.Y(_09653_),
    .A(_09652_));
 sg13g2_buf_2 _15745_ (.A(\exec.sp[3] ),
    .X(_09654_));
 sg13g2_nor4_2 _15746_ (.A(_09614_),
    .B(net1311),
    .C(net1310),
    .Y(_09655_),
    .D(_09654_));
 sg13g2_xnor2_1 _15747_ (.Y(_09656_),
    .A(_09653_),
    .B(_09655_));
 sg13g2_buf_8 _15748_ (.A(_09656_),
    .X(_09657_));
 sg13g2_mux2_1 _15749_ (.A0(_09646_),
    .A1(_09651_),
    .S(net872),
    .X(_09658_));
 sg13g2_buf_1 _15750_ (.A(_09658_),
    .X(_09659_));
 sg13g2_buf_1 _15751_ (.A(_09659_),
    .X(_09660_));
 sg13g2_buf_1 _15752_ (.A(net1281),
    .X(_09661_));
 sg13g2_mux4_1 _15753_ (.S0(_09616_),
    .A0(\stack[19][1] ),
    .A1(\stack[16][1] ),
    .A2(\stack[17][1] ),
    .A3(\stack[18][1] ),
    .S1(net1204),
    .X(_09662_));
 sg13g2_mux4_1 _15754_ (.S0(_09616_),
    .A0(\stack[3][1] ),
    .A1(\stack[0][1] ),
    .A2(\stack[1][1] ),
    .A3(\stack[2][1] ),
    .S1(_09623_),
    .X(_09663_));
 sg13g2_buf_8 _15755_ (.A(net1282),
    .X(_09664_));
 sg13g2_mux4_1 _15756_ (.S0(net1203),
    .A0(\stack[23][1] ),
    .A1(\stack[20][1] ),
    .A2(\stack[21][1] ),
    .A3(\stack[22][1] ),
    .S1(net1204),
    .X(_09665_));
 sg13g2_mux4_1 _15757_ (.S0(net1206),
    .A0(\stack[7][1] ),
    .A1(\stack[4][1] ),
    .A2(\stack[5][1] ),
    .A3(\stack[6][1] ),
    .S1(net1204),
    .X(_09666_));
 sg13g2_mux4_1 _15758_ (.S0(net872),
    .A0(_09662_),
    .A1(_09663_),
    .A2(_09665_),
    .A3(_09666_),
    .S1(net562),
    .X(_09667_));
 sg13g2_nand2_1 _15759_ (.Y(_09668_),
    .A(_09637_),
    .B(_09667_));
 sg13g2_buf_8 _15760_ (.A(_09640_),
    .X(_09669_));
 sg13g2_xor2_1 _15761_ (.B(_09652_),
    .A(_09654_),
    .X(_09670_));
 sg13g2_or3_1 _15762_ (.A(_09633_),
    .B(net871),
    .C(_09670_),
    .X(_09671_));
 sg13g2_nand3_1 _15763_ (.B(_09652_),
    .C(net871),
    .A(_09633_),
    .Y(_09672_));
 sg13g2_nand2_1 _15764_ (.Y(_09673_),
    .A(_09671_),
    .B(_09672_));
 sg13g2_buf_8 _15765_ (.A(_09673_),
    .X(_09674_));
 sg13g2_buf_8 _15766_ (.A(_09621_),
    .X(_09675_));
 sg13g2_buf_2 _15767_ (.A(net1280),
    .X(_09676_));
 sg13g2_buf_8 _15768_ (.A(net1310),
    .X(_09677_));
 sg13g2_buf_8 _15769_ (.A(net1279),
    .X(_09678_));
 sg13g2_mux2_1 _15770_ (.A0(\stack[15][1] ),
    .A1(\stack[11][1] ),
    .S(net1201),
    .X(_09679_));
 sg13g2_nor2_1 _15771_ (.A(net1202),
    .B(_09679_),
    .Y(_09680_));
 sg13g2_nand2_1 _15772_ (.Y(_09681_),
    .A(net1281),
    .B(net1279));
 sg13g2_inv_1 _15773_ (.Y(_09682_),
    .A(net1282));
 sg13g2_buf_1 _15774_ (.A(_09682_),
    .X(_09683_));
 sg13g2_o21ai_1 _15775_ (.B1(net870),
    .Y(_09684_),
    .A1(\stack[13][1] ),
    .A2(_09681_));
 sg13g2_and2_1 _15776_ (.A(net1282),
    .B(net1281),
    .X(_09685_));
 sg13g2_buf_1 _15777_ (.A(_09685_),
    .X(_09686_));
 sg13g2_buf_1 _15778_ (.A(\stack[10][1] ),
    .X(_09687_));
 sg13g2_mux2_1 _15779_ (.A0(_09687_),
    .A1(\stack[14][1] ),
    .S(net1201),
    .X(_09688_));
 sg13g2_nor2b_1 _15780_ (.A(net1280),
    .B_N(net1282),
    .Y(_09689_));
 sg13g2_mux2_1 _15781_ (.A0(\stack[8][1] ),
    .A1(\stack[12][1] ),
    .S(net1201),
    .X(_09690_));
 sg13g2_a22oi_1 _15782_ (.Y(_09691_),
    .B1(_09689_),
    .B2(_09690_),
    .A2(_09688_),
    .A1(_09686_));
 sg13g2_o21ai_1 _15783_ (.B1(_09691_),
    .Y(_09692_),
    .A1(_09680_),
    .A2(_09684_));
 sg13g2_nor2b_1 _15784_ (.A(net1279),
    .B_N(net1281),
    .Y(_09693_));
 sg13g2_buf_2 _15785_ (.A(_09693_),
    .X(_09694_));
 sg13g2_buf_8 _15786_ (.A(_09615_),
    .X(_09695_));
 sg13g2_buf_8 _15787_ (.A(net1200),
    .X(_09696_));
 sg13g2_nand2_1 _15788_ (.Y(_09697_),
    .A(net869),
    .B(_09687_));
 sg13g2_nand2_1 _15789_ (.Y(_09698_),
    .A(net870),
    .B(\stack[9][1] ));
 sg13g2_nand3_1 _15790_ (.B(_09697_),
    .C(_09698_),
    .A(_09694_),
    .Y(_09699_));
 sg13g2_nand3_1 _15791_ (.B(_09692_),
    .C(_09699_),
    .A(_09674_),
    .Y(_09700_));
 sg13g2_nor2_1 _15792_ (.A(_09637_),
    .B(net872),
    .Y(_09701_));
 sg13g2_buf_8 _15793_ (.A(net1280),
    .X(_09702_));
 sg13g2_mux4_1 _15794_ (.S0(net1200),
    .A0(\stack[27][1] ),
    .A1(\stack[24][1] ),
    .A2(\stack[25][1] ),
    .A3(\stack[26][1] ),
    .S1(net1199),
    .X(_09703_));
 sg13g2_mux4_1 _15795_ (.S0(net1200),
    .A0(\stack[31][1] ),
    .A1(\stack[28][1] ),
    .A2(\stack[29][1] ),
    .A3(\stack[30][1] ),
    .S1(net1199),
    .X(_09704_));
 sg13g2_mux2_1 _15796_ (.A0(_09703_),
    .A1(_09704_),
    .S(_09644_),
    .X(_09705_));
 sg13g2_nand2_1 _15797_ (.Y(_09706_),
    .A(_09701_),
    .B(_09705_));
 sg13g2_and3_1 _15798_ (.X(_09707_),
    .A(_09668_),
    .B(_09700_),
    .C(_09706_));
 sg13g2_buf_2 _15799_ (.A(_09707_),
    .X(_09708_));
 sg13g2_xnor2_1 _15800_ (.Y(_09709_),
    .A(_09632_),
    .B(_09635_));
 sg13g2_buf_2 _15801_ (.A(_09709_),
    .X(_09710_));
 sg13g2_buf_1 _15802_ (.A(net1279),
    .X(_09711_));
 sg13g2_buf_1 _15803_ (.A(net1198),
    .X(_09712_));
 sg13g2_buf_8 _15804_ (.A(net1203),
    .X(_09713_));
 sg13g2_buf_8 _15805_ (.A(net867),
    .X(_09714_));
 sg13g2_mux2_1 _15806_ (.A0(_00044_),
    .A1(_00046_),
    .S(net1204),
    .X(_09715_));
 sg13g2_nor2b_1 _15807_ (.A(_09614_),
    .B_N(net1311),
    .Y(_09716_));
 sg13g2_buf_1 _15808_ (.A(_09716_),
    .X(_09717_));
 sg13g2_a22oi_1 _15809_ (.Y(_09718_),
    .B1(net1197),
    .B2(_00045_),
    .A2(_09715_),
    .A1(net786));
 sg13g2_nor2_2 _15810_ (.A(net1282),
    .B(net1281),
    .Y(_09719_));
 sg13g2_mux2_1 _15811_ (.A0(_00040_),
    .A1(_00042_),
    .S(net1204),
    .X(_09720_));
 sg13g2_a221oi_1 _15812_ (.B2(net786),
    .C1(net868),
    .B1(_09720_),
    .A1(_00047_),
    .Y(_09721_),
    .A2(_09719_));
 sg13g2_a21o_1 _15813_ (.A2(_09718_),
    .A1(net868),
    .B1(_09721_),
    .X(_09722_));
 sg13g2_buf_1 _15814_ (.A(net870),
    .X(_09723_));
 sg13g2_inv_1 _15815_ (.Y(_09724_),
    .A(_00043_));
 sg13g2_nand2b_1 _15816_ (.Y(_09725_),
    .B(net1310),
    .A_N(net1311));
 sg13g2_buf_2 _15817_ (.A(_09725_),
    .X(_09726_));
 sg13g2_buf_8 _15818_ (.A(_09726_),
    .X(_09727_));
 sg13g2_nand3b_1 _15819_ (.B(_00041_),
    .C(net1202),
    .Y(_09728_),
    .A_N(net1198));
 sg13g2_o21ai_1 _15820_ (.B1(_09728_),
    .Y(_09729_),
    .A1(_09724_),
    .A2(net866));
 sg13g2_xnor2_1 _15821_ (.Y(_09730_),
    .A(_09652_),
    .B(_09655_));
 sg13g2_a21oi_1 _15822_ (.A1(net785),
    .A2(_09729_),
    .Y(_09731_),
    .B1(_09730_));
 sg13g2_buf_8 _15823_ (.A(_09719_),
    .X(_09732_));
 sg13g2_mux2_1 _15824_ (.A0(_00061_),
    .A1(_00063_),
    .S(net1205),
    .X(_09733_));
 sg13g2_buf_8 _15825_ (.A(net1206),
    .X(_09734_));
 sg13g2_buf_8 _15826_ (.A(net864),
    .X(_09735_));
 sg13g2_a22oi_1 _15827_ (.Y(_09736_),
    .B1(_09733_),
    .B2(net784),
    .A2(net865),
    .A1(_00060_));
 sg13g2_mux2_1 _15828_ (.A0(_00057_),
    .A1(_00059_),
    .S(net1205),
    .X(_09737_));
 sg13g2_a221oi_1 _15829_ (.B2(net786),
    .C1(net868),
    .B1(_09737_),
    .A1(_00058_),
    .Y(_09738_),
    .A2(net1197));
 sg13g2_a21o_1 _15830_ (.A2(_09736_),
    .A1(net868),
    .B1(_09738_),
    .X(_09739_));
 sg13g2_inv_1 _15831_ (.Y(_09740_),
    .A(_00064_));
 sg13g2_or2_1 _15832_ (.X(_09741_),
    .B(net1310),
    .A(_09621_));
 sg13g2_buf_2 _15833_ (.A(_09741_),
    .X(_09742_));
 sg13g2_buf_1 _15834_ (.A(_09742_),
    .X(_09743_));
 sg13g2_buf_8 _15835_ (.A(net1281),
    .X(_09744_));
 sg13g2_buf_1 _15836_ (.A(net1196),
    .X(_09745_));
 sg13g2_buf_1 _15837_ (.A(net1201),
    .X(_09746_));
 sg13g2_nand3_1 _15838_ (.B(net861),
    .C(_00062_),
    .A(net862),
    .Y(_09747_));
 sg13g2_o21ai_1 _15839_ (.B1(_09747_),
    .Y(_09748_),
    .A1(_09740_),
    .A2(net863));
 sg13g2_a21oi_1 _15840_ (.A1(net785),
    .A2(_09748_),
    .Y(_09749_),
    .B1(net872));
 sg13g2_a22oi_1 _15841_ (.Y(_09750_),
    .B1(_09739_),
    .B2(_09749_),
    .A2(_09731_),
    .A1(_09722_));
 sg13g2_mux2_1 _15842_ (.A0(_00035_),
    .A1(_00037_),
    .S(net1196),
    .X(_09751_));
 sg13g2_a22oi_1 _15843_ (.Y(_09752_),
    .B1(_09751_),
    .B2(net786),
    .A2(net1197),
    .A1(_00036_));
 sg13g2_mux2_1 _15844_ (.A0(_00031_),
    .A1(_00033_),
    .S(net1196),
    .X(_09753_));
 sg13g2_a221oi_1 _15845_ (.B2(net869),
    .C1(net861),
    .B1(_09753_),
    .A1(_00038_),
    .Y(_09754_),
    .A2(_09719_));
 sg13g2_a21o_1 _15846_ (.A2(_09752_),
    .A1(net868),
    .B1(_09754_),
    .X(_09755_));
 sg13g2_inv_1 _15847_ (.Y(_09756_),
    .A(_00034_));
 sg13g2_nand3b_1 _15848_ (.B(net1199),
    .C(_00032_),
    .Y(_09757_),
    .A_N(_09711_));
 sg13g2_o21ai_1 _15849_ (.B1(_09757_),
    .Y(_09758_),
    .A1(_09756_),
    .A2(_09727_));
 sg13g2_a21oi_1 _15850_ (.A1(net870),
    .A2(_09758_),
    .Y(_09759_),
    .B1(_09730_));
 sg13g2_mux2_1 _15851_ (.A0(_00053_),
    .A1(_00055_),
    .S(net1204),
    .X(_09760_));
 sg13g2_a22oi_1 _15852_ (.Y(_09761_),
    .B1(_09760_),
    .B2(net786),
    .A2(net865),
    .A1(_00052_));
 sg13g2_mux2_1 _15853_ (.A0(_00049_),
    .A1(_00051_),
    .S(net1196),
    .X(_09762_));
 sg13g2_a221oi_1 _15854_ (.B2(net869),
    .C1(net861),
    .B1(_09762_),
    .A1(_00050_),
    .Y(_09763_),
    .A2(net1197));
 sg13g2_a21o_1 _15855_ (.A2(_09761_),
    .A1(net868),
    .B1(_09763_),
    .X(_09764_));
 sg13g2_inv_1 _15856_ (.Y(_09765_),
    .A(_00056_));
 sg13g2_nand3_1 _15857_ (.B(net1198),
    .C(_00054_),
    .A(net1202),
    .Y(_09766_));
 sg13g2_o21ai_1 _15858_ (.B1(_09766_),
    .Y(_09767_),
    .A1(_09765_),
    .A2(_09742_));
 sg13g2_a21oi_1 _15859_ (.A1(net785),
    .A2(_09767_),
    .Y(_09768_),
    .B1(_09657_));
 sg13g2_a221oi_1 _15860_ (.B2(_09768_),
    .C1(_09710_),
    .B1(_09764_),
    .A1(_09755_),
    .Y(_09769_),
    .A2(_09759_));
 sg13g2_a21o_1 _15861_ (.A2(_09750_),
    .A1(_09710_),
    .B1(_09769_),
    .X(_09770_));
 sg13g2_buf_2 _15862_ (.A(_09770_),
    .X(_09771_));
 sg13g2_buf_8 _15863_ (.A(_09771_),
    .X(_09772_));
 sg13g2_mux4_1 _15864_ (.S0(net1203),
    .A0(\stack[19][3] ),
    .A1(\stack[16][3] ),
    .A2(\stack[17][3] ),
    .A3(\stack[18][3] ),
    .S1(net1196),
    .X(_09773_));
 sg13g2_mux4_1 _15865_ (.S0(net1203),
    .A0(\stack[3][3] ),
    .A1(\stack[0][3] ),
    .A2(\stack[1][3] ),
    .A3(\stack[2][3] ),
    .S1(net1196),
    .X(_09774_));
 sg13g2_mux4_1 _15866_ (.S0(_09664_),
    .A0(\stack[23][3] ),
    .A1(\stack[20][3] ),
    .A2(\stack[21][3] ),
    .A3(\stack[22][3] ),
    .S1(_09744_),
    .X(_09775_));
 sg13g2_mux4_1 _15867_ (.S0(net1203),
    .A0(\stack[7][3] ),
    .A1(\stack[4][3] ),
    .A2(\stack[5][3] ),
    .A3(\stack[6][3] ),
    .S1(net1196),
    .X(_09776_));
 sg13g2_mux4_1 _15868_ (.S0(net872),
    .A0(_09773_),
    .A1(_09774_),
    .A2(_09775_),
    .A3(_09776_),
    .S1(_09644_),
    .X(_09777_));
 sg13g2_mux4_1 _15869_ (.S0(net1200),
    .A0(\stack[27][3] ),
    .A1(\stack[24][3] ),
    .A2(\stack[25][3] ),
    .A3(\stack[26][3] ),
    .S1(net1199),
    .X(_09778_));
 sg13g2_mux4_1 _15870_ (.S0(net1206),
    .A0(\stack[31][3] ),
    .A1(\stack[28][3] ),
    .A2(\stack[29][3] ),
    .A3(\stack[30][3] ),
    .S1(net1205),
    .X(_09779_));
 sg13g2_mux2_1 _15871_ (.A0(_09778_),
    .A1(_09779_),
    .S(_09644_),
    .X(_09780_));
 sg13g2_mux4_1 _15872_ (.S0(net1206),
    .A0(\stack[11][3] ),
    .A1(\stack[12][3] ),
    .A2(\stack[13][3] ),
    .A3(\stack[14][3] ),
    .S1(net1205),
    .X(_09781_));
 sg13g2_nand2_1 _15873_ (.Y(_09782_),
    .A(net861),
    .B(_09781_));
 sg13g2_buf_2 _15874_ (.A(net1282),
    .X(_09783_));
 sg13g2_mux4_1 _15875_ (.S0(net1280),
    .A0(\stack[15][3] ),
    .A1(\stack[9][3] ),
    .A2(\stack[8][3] ),
    .A3(\stack[10][3] ),
    .S1(net1195),
    .X(_09784_));
 sg13g2_nand2b_1 _15876_ (.Y(_09785_),
    .B(_09784_),
    .A_N(net861));
 sg13g2_a22oi_1 _15877_ (.Y(_09786_),
    .B1(_09782_),
    .B2(_09785_),
    .A2(_09672_),
    .A1(_09671_));
 sg13g2_a221oi_1 _15878_ (.B2(_09701_),
    .C1(_09786_),
    .B1(_09780_),
    .A1(_09637_),
    .Y(_09787_),
    .A2(_09777_));
 sg13g2_buf_2 _15879_ (.A(_09787_),
    .X(_09788_));
 sg13g2_mux4_1 _15880_ (.S0(net1206),
    .A0(\stack[11][2] ),
    .A1(\stack[8][2] ),
    .A2(\stack[9][2] ),
    .A3(\stack[10][2] ),
    .S1(net1205),
    .X(_09789_));
 sg13g2_mux4_1 _15881_ (.S0(net1206),
    .A0(\stack[15][2] ),
    .A1(\stack[12][2] ),
    .A2(\stack[13][2] ),
    .A3(\stack[14][2] ),
    .S1(net1205),
    .X(_09790_));
 sg13g2_mux2_1 _15882_ (.A0(_09789_),
    .A1(_09790_),
    .S(_09644_),
    .X(_09791_));
 sg13g2_mux4_1 _15883_ (.S0(net1203),
    .A0(\stack[19][2] ),
    .A1(\stack[16][2] ),
    .A2(\stack[17][2] ),
    .A3(\stack[18][2] ),
    .S1(net1204),
    .X(_09792_));
 sg13g2_mux4_1 _15884_ (.S0(net1203),
    .A0(\stack[3][2] ),
    .A1(\stack[0][2] ),
    .A2(\stack[1][2] ),
    .A3(\stack[2][2] ),
    .S1(_09661_),
    .X(_09793_));
 sg13g2_mux4_1 _15885_ (.S0(_09664_),
    .A0(\stack[23][2] ),
    .A1(\stack[20][2] ),
    .A2(\stack[21][2] ),
    .A3(\stack[22][2] ),
    .S1(_09744_),
    .X(_09794_));
 sg13g2_mux4_1 _15886_ (.S0(net1203),
    .A0(\stack[7][2] ),
    .A1(\stack[4][2] ),
    .A2(\stack[5][2] ),
    .A3(\stack[6][2] ),
    .S1(net1196),
    .X(_09795_));
 sg13g2_mux4_1 _15887_ (.S0(_09657_),
    .A0(_09792_),
    .A1(_09793_),
    .A2(_09794_),
    .A3(_09795_),
    .S1(_09645_),
    .X(_09796_));
 sg13g2_nand3_1 _15888_ (.B(_09635_),
    .C(_09670_),
    .A(_09632_),
    .Y(_09797_));
 sg13g2_buf_1 _15889_ (.A(_09797_),
    .X(_09798_));
 sg13g2_nand3_1 _15890_ (.B(_09653_),
    .C(net871),
    .A(_09633_),
    .Y(_09799_));
 sg13g2_buf_1 _15891_ (.A(_09799_),
    .X(_09800_));
 sg13g2_mux4_1 _15892_ (.S0(net1201),
    .A0(\stack[24][2] ),
    .A1(\stack[28][2] ),
    .A2(\stack[26][2] ),
    .A3(\stack[30][2] ),
    .S1(net1205),
    .X(_09801_));
 sg13g2_nand2_1 _15893_ (.Y(_09802_),
    .A(net786),
    .B(_09801_));
 sg13g2_mux4_1 _15894_ (.S0(net1280),
    .A0(\stack[31][2] ),
    .A1(\stack[25][2] ),
    .A2(\stack[27][2] ),
    .A3(\stack[29][2] ),
    .S1(net1198),
    .X(_09803_));
 sg13g2_nand2_1 _15895_ (.Y(_09804_),
    .A(net870),
    .B(_09803_));
 sg13g2_a22oi_1 _15896_ (.Y(_09805_),
    .B1(_09802_),
    .B2(_09804_),
    .A2(_09800_),
    .A1(_09798_));
 sg13g2_a221oi_1 _15897_ (.B2(_09637_),
    .C1(_09805_),
    .B1(_09796_),
    .A1(_09674_),
    .Y(_09806_),
    .A2(_09791_));
 sg13g2_buf_2 _15898_ (.A(_09806_),
    .X(_09807_));
 sg13g2_and2_1 _15899_ (.A(_09788_),
    .B(_09807_),
    .X(_09808_));
 sg13g2_buf_8 _15900_ (.A(_09808_),
    .X(_09809_));
 sg13g2_mux4_1 _15901_ (.S0(_09619_),
    .A0(\stack[27][6] ),
    .A1(\stack[24][6] ),
    .A2(\stack[25][6] ),
    .A3(\stack[26][6] ),
    .S1(net564),
    .X(_09810_));
 sg13g2_mux4_1 _15902_ (.S0(net565),
    .A0(\stack[19][6] ),
    .A1(\stack[16][6] ),
    .A2(\stack[17][6] ),
    .A3(\stack[18][6] ),
    .S1(_09626_),
    .X(_09811_));
 sg13g2_buf_8 _15903_ (.A(net784),
    .X(_09812_));
 sg13g2_mux4_1 _15904_ (.S0(net561),
    .A0(\stack[31][6] ),
    .A1(\stack[28][6] ),
    .A2(\stack[29][6] ),
    .A3(\stack[30][6] ),
    .S1(_09626_),
    .X(_09813_));
 sg13g2_mux4_1 _15905_ (.S0(net561),
    .A0(\stack[23][6] ),
    .A1(\stack[20][6] ),
    .A2(\stack[21][6] ),
    .A3(\stack[22][6] ),
    .S1(net564),
    .X(_09814_));
 sg13g2_mux4_1 _15906_ (.S0(_09638_),
    .A0(_09810_),
    .A1(_09811_),
    .A2(_09813_),
    .A3(_09814_),
    .S1(net562),
    .X(_09815_));
 sg13g2_mux4_1 _15907_ (.S0(net561),
    .A0(\stack[11][6] ),
    .A1(\stack[8][6] ),
    .A2(\stack[9][6] ),
    .A3(\stack[10][6] ),
    .S1(net564),
    .X(_09816_));
 sg13g2_mux4_1 _15908_ (.S0(net561),
    .A0(\stack[3][6] ),
    .A1(\stack[0][6] ),
    .A2(\stack[1][6] ),
    .A3(\stack[2][6] ),
    .S1(net564),
    .X(_09817_));
 sg13g2_mux4_1 _15909_ (.S0(net561),
    .A0(\stack[15][6] ),
    .A1(\stack[12][6] ),
    .A2(\stack[13][6] ),
    .A3(\stack[14][6] ),
    .S1(net787),
    .X(_09818_));
 sg13g2_mux4_1 _15910_ (.S0(_09812_),
    .A0(\stack[7][6] ),
    .A1(\stack[4][6] ),
    .A2(\stack[5][6] ),
    .A3(\stack[6][6] ),
    .S1(net787),
    .X(_09819_));
 sg13g2_mux4_1 _15911_ (.S0(net563),
    .A0(_09816_),
    .A1(_09817_),
    .A2(_09818_),
    .A3(_09819_),
    .S1(net562),
    .X(_09820_));
 sg13g2_mux2_1 _15912_ (.A0(_09815_),
    .A1(_09820_),
    .S(net872),
    .X(_09821_));
 sg13g2_buf_1 _15913_ (.A(_09821_),
    .X(_09822_));
 sg13g2_buf_8 _15914_ (.A(net786),
    .X(_09823_));
 sg13g2_mux4_1 _15915_ (.S0(net560),
    .A0(\stack[23][5] ),
    .A1(\stack[20][5] ),
    .A2(\stack[21][5] ),
    .A3(\stack[22][5] ),
    .S1(net787),
    .X(_09824_));
 sg13g2_inv_1 _15916_ (.Y(_09825_),
    .A(_09824_));
 sg13g2_mux4_1 _15917_ (.S0(net560),
    .A0(\stack[7][5] ),
    .A1(\stack[4][5] ),
    .A2(\stack[5][5] ),
    .A3(\stack[6][5] ),
    .S1(_09625_),
    .X(_09826_));
 sg13g2_inv_1 _15918_ (.Y(_09827_),
    .A(_09826_));
 sg13g2_mux4_1 _15919_ (.S0(net788),
    .A0(\stack[19][5] ),
    .A1(\stack[16][5] ),
    .A2(\stack[17][5] ),
    .A3(\stack[18][5] ),
    .S1(net787),
    .X(_09828_));
 sg13g2_inv_1 _15920_ (.Y(_09829_),
    .A(_09828_));
 sg13g2_mux4_1 _15921_ (.S0(net788),
    .A0(\stack[3][5] ),
    .A1(\stack[0][5] ),
    .A2(\stack[1][5] ),
    .A3(\stack[2][5] ),
    .S1(_09625_),
    .X(_09830_));
 sg13g2_inv_1 _15922_ (.Y(_09831_),
    .A(_09830_));
 sg13g2_and2_1 _15923_ (.A(_09669_),
    .B(_09642_),
    .X(_09832_));
 sg13g2_mux4_1 _15924_ (.S0(net872),
    .A0(_09825_),
    .A1(_09827_),
    .A2(_09829_),
    .A3(_09831_),
    .S1(_09832_),
    .X(_09833_));
 sg13g2_mux4_1 _15925_ (.S0(net565),
    .A0(\stack[11][5] ),
    .A1(\stack[8][5] ),
    .A2(\stack[9][5] ),
    .A3(\stack[10][5] ),
    .S1(net564),
    .X(_09834_));
 sg13g2_mux4_1 _15926_ (.S0(net560),
    .A0(\stack[15][5] ),
    .A1(\stack[12][5] ),
    .A2(\stack[13][5] ),
    .A3(\stack[14][5] ),
    .S1(net787),
    .X(_09835_));
 sg13g2_a21o_1 _15927_ (.A2(_09642_),
    .A1(net871),
    .B1(_09835_),
    .X(_09836_));
 sg13g2_o21ai_1 _15928_ (.B1(_09836_),
    .Y(_09837_),
    .A1(net562),
    .A2(_09834_));
 sg13g2_mux4_1 _15929_ (.S0(net565),
    .A0(\stack[31][5] ),
    .A1(\stack[28][5] ),
    .A2(\stack[29][5] ),
    .A3(\stack[30][5] ),
    .S1(net564),
    .X(_09838_));
 sg13g2_mux4_1 _15930_ (.S0(net560),
    .A0(\stack[27][5] ),
    .A1(\stack[24][5] ),
    .A2(\stack[25][5] ),
    .A3(\stack[26][5] ),
    .S1(net787),
    .X(_09839_));
 sg13g2_and3_1 _15931_ (.X(_09840_),
    .A(net871),
    .B(_09642_),
    .C(_09839_));
 sg13g2_a221oi_1 _15932_ (.B2(net562),
    .C1(_09840_),
    .B1(_09838_),
    .A1(_09798_),
    .Y(_09841_),
    .A2(_09800_));
 sg13g2_a221oi_1 _15933_ (.B2(_09837_),
    .C1(_09841_),
    .B1(_09674_),
    .A1(net563),
    .Y(_09842_),
    .A2(_09833_));
 sg13g2_buf_1 _15934_ (.A(_09842_),
    .X(_09843_));
 sg13g2_mux4_1 _15935_ (.S0(net874),
    .A0(\stack[23][4] ),
    .A1(\stack[20][4] ),
    .A2(\stack[21][4] ),
    .A3(\stack[22][4] ),
    .S1(net873),
    .X(_09844_));
 sg13g2_inv_1 _15936_ (.Y(_09845_),
    .A(_09844_));
 sg13g2_mux4_1 _15937_ (.S0(net874),
    .A0(\stack[7][4] ),
    .A1(\stack[4][4] ),
    .A2(\stack[5][4] ),
    .A3(\stack[6][4] ),
    .S1(net873),
    .X(_09846_));
 sg13g2_inv_1 _15938_ (.Y(_09847_),
    .A(_09846_));
 sg13g2_mux4_1 _15939_ (.S0(net864),
    .A0(\stack[19][4] ),
    .A1(\stack[16][4] ),
    .A2(\stack[17][4] ),
    .A3(\stack[18][4] ),
    .S1(_09624_),
    .X(_09848_));
 sg13g2_inv_1 _15940_ (.Y(_09849_),
    .A(_09848_));
 sg13g2_mux4_1 _15941_ (.S0(net874),
    .A0(\stack[3][4] ),
    .A1(\stack[0][4] ),
    .A2(\stack[1][4] ),
    .A3(\stack[2][4] ),
    .S1(net873),
    .X(_09850_));
 sg13g2_inv_1 _15942_ (.Y(_09851_),
    .A(_09850_));
 sg13g2_mux4_1 _15943_ (.S0(net872),
    .A0(_09845_),
    .A1(_09847_),
    .A2(_09849_),
    .A3(_09851_),
    .S1(_09832_),
    .X(_09852_));
 sg13g2_buf_2 _15944_ (.A(net1199),
    .X(_09853_));
 sg13g2_mux4_1 _15945_ (.S0(net784),
    .A0(\stack[11][4] ),
    .A1(\stack[8][4] ),
    .A2(\stack[9][4] ),
    .A3(\stack[10][4] ),
    .S1(net860),
    .X(_09854_));
 sg13g2_mux4_1 _15946_ (.S0(net869),
    .A0(\stack[15][4] ),
    .A1(\stack[12][4] ),
    .A2(\stack[13][4] ),
    .A3(\stack[14][4] ),
    .S1(net860),
    .X(_09855_));
 sg13g2_a21o_1 _15947_ (.A2(_09642_),
    .A1(net871),
    .B1(_09855_),
    .X(_09856_));
 sg13g2_o21ai_1 _15948_ (.B1(_09856_),
    .Y(_09857_),
    .A1(net562),
    .A2(_09854_));
 sg13g2_buf_1 _15949_ (.A(\stack[31][4] ),
    .X(_09858_));
 sg13g2_mux4_1 _15950_ (.S0(net784),
    .A0(_09858_),
    .A1(\stack[28][4] ),
    .A2(\stack[29][4] ),
    .A3(\stack[30][4] ),
    .S1(net860),
    .X(_09859_));
 sg13g2_mux4_1 _15951_ (.S0(_09696_),
    .A0(\stack[27][4] ),
    .A1(\stack[24][4] ),
    .A2(\stack[25][4] ),
    .A3(\stack[26][4] ),
    .S1(net860),
    .X(_09860_));
 sg13g2_and3_1 _15952_ (.X(_09861_),
    .A(net871),
    .B(_09642_),
    .C(_09860_));
 sg13g2_a221oi_1 _15953_ (.B2(net562),
    .C1(_09861_),
    .B1(_09859_),
    .A1(_09798_),
    .Y(_09862_),
    .A2(_09800_));
 sg13g2_a221oi_1 _15954_ (.B2(_09674_),
    .C1(_09862_),
    .B1(_09857_),
    .A1(net563),
    .Y(_09863_),
    .A2(_09852_));
 sg13g2_buf_2 _15955_ (.A(_09863_),
    .X(_09864_));
 sg13g2_nor3_1 _15956_ (.A(net497),
    .B(_09843_),
    .C(_09864_),
    .Y(_09865_));
 sg13g2_nand4_1 _15957_ (.B(net487),
    .C(_09809_),
    .A(_09708_),
    .Y(_09866_),
    .D(_09865_));
 sg13g2_buf_1 _15958_ (.A(_09866_),
    .X(_09867_));
 sg13g2_buf_1 _15959_ (.A(\exec.opcode[7] ),
    .X(_09868_));
 sg13g2_buf_1 _15960_ (.A(\exec.opcode[5] ),
    .X(_09869_));
 sg13g2_nand2b_1 _15961_ (.Y(_09870_),
    .B(net1308),
    .A_N(net1309));
 sg13g2_buf_8 _15962_ (.A(\exec.opcode[6] ),
    .X(_09871_));
 sg13g2_or2_1 _15963_ (.X(_09872_),
    .B(net1307),
    .A(\exec.opcode[4] ));
 sg13g2_buf_1 _15964_ (.A(_09872_),
    .X(_09873_));
 sg13g2_nor2_1 _15965_ (.A(_09870_),
    .B(_09873_),
    .Y(_09874_));
 sg13g2_buf_2 _15966_ (.A(_09874_),
    .X(_09875_));
 sg13g2_buf_2 _15967_ (.A(\exec.opcode[1] ),
    .X(_09876_));
 sg13g2_buf_1 _15968_ (.A(_09876_),
    .X(_09877_));
 sg13g2_buf_1 _15969_ (.A(\exec.opcode[0] ),
    .X(_09878_));
 sg13g2_nor2_1 _15970_ (.A(net1278),
    .B(net1306),
    .Y(_09879_));
 sg13g2_buf_1 _15971_ (.A(\exec.opcode[3] ),
    .X(_09880_));
 sg13g2_buf_2 _15972_ (.A(\exec.opcode[2] ),
    .X(_09881_));
 sg13g2_and2_1 _15973_ (.A(_09880_),
    .B(_09881_),
    .X(_09882_));
 sg13g2_buf_1 _15974_ (.A(_09882_),
    .X(_09883_));
 sg13g2_and2_1 _15975_ (.A(_09879_),
    .B(_09883_),
    .X(_09884_));
 sg13g2_buf_1 _15976_ (.A(_09884_),
    .X(_09885_));
 sg13g2_and2_1 _15977_ (.A(_09875_),
    .B(_09885_),
    .X(_09886_));
 sg13g2_buf_1 _15978_ (.A(_09886_),
    .X(_09887_));
 sg13g2_o21ai_1 _15979_ (.B1(_09887_),
    .Y(_09888_),
    .A1(net474),
    .A2(_09867_));
 sg13g2_buf_1 _15980_ (.A(_09880_),
    .X(_09889_));
 sg13g2_inv_2 _15981_ (.Y(_09890_),
    .A(net1277));
 sg13g2_nor2b_1 _15982_ (.A(net1309),
    .B_N(net1308),
    .Y(_09891_));
 sg13g2_or2_1 _15983_ (.X(_09892_),
    .B(_09881_),
    .A(_09876_));
 sg13g2_buf_1 _15984_ (.A(\exec.opcode[4] ),
    .X(_09893_));
 sg13g2_nand4_1 _15985_ (.B(_09881_),
    .C(net1305),
    .A(_09876_),
    .Y(_09894_),
    .D(net1307));
 sg13g2_o21ai_1 _15986_ (.B1(_09894_),
    .Y(_09895_),
    .A1(_09873_),
    .A2(_09892_));
 sg13g2_nand4_1 _15987_ (.B(_09890_),
    .C(_09891_),
    .A(net1306),
    .Y(_09896_),
    .D(_09895_));
 sg13g2_buf_1 _15988_ (.A(_09896_),
    .X(_09897_));
 sg13g2_nand2_1 _15989_ (.Y(_09898_),
    .A(net1278),
    .B(_09871_));
 sg13g2_nand2_1 _15990_ (.Y(_09899_),
    .A(net1306),
    .B(_09868_));
 sg13g2_nand2_1 _15991_ (.Y(_09900_),
    .A(net1305),
    .B(net1308));
 sg13g2_buf_2 _15992_ (.A(_09900_),
    .X(_09901_));
 sg13g2_nor3_1 _15993_ (.A(_09898_),
    .B(_09899_),
    .C(_09901_),
    .Y(_09902_));
 sg13g2_buf_1 _15994_ (.A(single_step),
    .X(_09903_));
 sg13g2_a21oi_1 _15995_ (.A1(_09883_),
    .A2(_09902_),
    .Y(_09904_),
    .B1(_09903_));
 sg13g2_nand2_1 _15996_ (.Y(_09905_),
    .A(net559),
    .B(_09904_));
 sg13g2_buf_2 _15997_ (.A(rst_n),
    .X(_09906_));
 sg13g2_buf_1 _15998_ (.A(_09906_),
    .X(_09907_));
 sg13g2_buf_1 _15999_ (.A(net1304),
    .X(_09908_));
 sg13g2_buf_1 _16000_ (.A(\state[3] ),
    .X(_09909_));
 sg13g2_nand2_1 _16001_ (.Y(_09910_),
    .A(net1276),
    .B(_09909_));
 sg13g2_buf_1 _16002_ (.A(_09910_),
    .X(_09911_));
 sg13g2_inv_1 _16003_ (.Y(_09912_),
    .A(_09881_));
 sg13g2_inv_1 _16004_ (.Y(_09913_),
    .A(net1278));
 sg13g2_buf_1 _16005_ (.A(net1306),
    .X(_09914_));
 sg13g2_nor2_1 _16006_ (.A(_09913_),
    .B(_09914_),
    .Y(_09915_));
 sg13g2_buf_1 _16007_ (.A(_09915_),
    .X(_09916_));
 sg13g2_nand2b_1 _16008_ (.Y(_09917_),
    .B(net1307),
    .A_N(net1309));
 sg13g2_buf_2 _16009_ (.A(_09917_),
    .X(_09918_));
 sg13g2_nor2_1 _16010_ (.A(_09901_),
    .B(_09918_),
    .Y(_09919_));
 sg13g2_and4_1 _16011_ (.A(net1277),
    .B(_09912_),
    .C(_09916_),
    .D(_09919_),
    .X(_09920_));
 sg13g2_or3_1 _16012_ (.A(_09905_),
    .B(net859),
    .C(_09920_),
    .X(_09921_));
 sg13g2_buf_1 _16013_ (.A(ui_in[6]),
    .X(_09922_));
 sg13g2_buf_1 _16014_ (.A(_09922_),
    .X(_09923_));
 sg13g2_buf_1 _16015_ (.A(ui_in[5]),
    .X(_09924_));
 sg13g2_nor2b_1 _16016_ (.A(_09924_),
    .B_N(net3),
    .Y(_09925_));
 sg13g2_nand2_1 _16017_ (.Y(_09926_),
    .A(net1303),
    .B(_09925_));
 sg13g2_buf_1 _16018_ (.A(_09926_),
    .X(_09927_));
 sg13g2_buf_2 _16019_ (.A(o_sleep),
    .X(_09928_));
 sg13g2_or2_2 _16020_ (.X(_09929_),
    .B(_09928_),
    .A(\state[4] ));
 sg13g2_nand3b_1 _16021_ (.B(_09929_),
    .C(net1),
    .Y(_09930_),
    .A_N(past_i_run));
 sg13g2_buf_1 _16022_ (.A(_09930_),
    .X(_09931_));
 sg13g2_nand2_1 _16023_ (.Y(_09932_),
    .A(_09906_),
    .B(_09931_));
 sg13g2_buf_1 _16024_ (.A(_09932_),
    .X(_09933_));
 sg13g2_buf_1 _16025_ (.A(o_wait_delay),
    .X(_09934_));
 sg13g2_inv_2 _16026_ (.Y(_09935_),
    .A(_09934_));
 sg13g2_nor2_1 _16027_ (.A(\delay_cycles[14] ),
    .B(\delay_cycles[19] ),
    .Y(_09936_));
 sg13g2_nor4_1 _16028_ (.A(\delay_cycles[20] ),
    .B(\delay_cycles[21] ),
    .C(\delay_cycles[22] ),
    .D(\delay_cycles[23] ),
    .Y(_09937_));
 sg13g2_nor4_1 _16029_ (.A(\delay_cycles[15] ),
    .B(\delay_cycles[16] ),
    .C(\delay_cycles[17] ),
    .D(\delay_cycles[18] ),
    .Y(_09938_));
 sg13g2_buf_1 _16030_ (.A(\delay_cycles[11] ),
    .X(_09939_));
 sg13g2_buf_1 _16031_ (.A(\delay_cycles[12] ),
    .X(_09940_));
 sg13g2_or2_1 _16032_ (.X(_09941_),
    .B(_09940_),
    .A(_09939_));
 sg13g2_inv_1 _16033_ (.Y(_09942_),
    .A(\delay_cycles[3] ));
 sg13g2_buf_1 _16034_ (.A(\delay_cycles[1] ),
    .X(_09943_));
 sg13g2_buf_1 _16035_ (.A(\delay_cycles[0] ),
    .X(_09944_));
 sg13g2_buf_1 _16036_ (.A(\delay_cycles[2] ),
    .X(_09945_));
 sg13g2_nand3_1 _16037_ (.B(_09944_),
    .C(_09945_),
    .A(_09943_),
    .Y(_09946_));
 sg13g2_buf_1 _16038_ (.A(_09946_),
    .X(_09947_));
 sg13g2_or2_1 _16039_ (.X(_09948_),
    .B(_09947_),
    .A(_09942_));
 sg13g2_buf_1 _16040_ (.A(_09948_),
    .X(_09949_));
 sg13g2_buf_1 _16041_ (.A(\delay_cycles[4] ),
    .X(_09950_));
 sg13g2_buf_1 _16042_ (.A(\delay_cycles[5] ),
    .X(_09951_));
 sg13g2_buf_1 _16043_ (.A(\delay_cycles[6] ),
    .X(_09952_));
 sg13g2_buf_1 _16044_ (.A(\delay_cycles[7] ),
    .X(_09953_));
 sg13g2_nor4_1 _16045_ (.A(_09950_),
    .B(_09951_),
    .C(_09952_),
    .D(_09953_),
    .Y(_09954_));
 sg13g2_buf_1 _16046_ (.A(\delay_cycles[8] ),
    .X(_09955_));
 sg13g2_buf_1 _16047_ (.A(\delay_cycles[9] ),
    .X(_09956_));
 sg13g2_buf_1 _16048_ (.A(\delay_cycles[10] ),
    .X(_09957_));
 sg13g2_nand3_1 _16049_ (.B(_09956_),
    .C(_09957_),
    .A(_09955_),
    .Y(_09958_));
 sg13g2_a21oi_1 _16050_ (.A1(_09949_),
    .A2(_09954_),
    .Y(_09959_),
    .B1(_09958_));
 sg13g2_o21ai_1 _16051_ (.B1(\delay_cycles[13] ),
    .Y(_09960_),
    .A1(_09941_),
    .A2(_09959_));
 sg13g2_nand4_1 _16052_ (.B(_09937_),
    .C(_09938_),
    .A(_09936_),
    .Y(_09961_),
    .D(_09960_));
 sg13g2_buf_1 _16053_ (.A(_09961_),
    .X(_09962_));
 sg13g2_or2_1 _16054_ (.X(_09963_),
    .B(_09962_),
    .A(_09935_));
 sg13g2_buf_1 _16055_ (.A(_09963_),
    .X(_09964_));
 sg13g2_buf_1 _16056_ (.A(_09934_),
    .X(_09965_));
 sg13g2_buf_1 _16057_ (.A(\delay_counter[7] ),
    .X(_09966_));
 sg13g2_buf_1 _16058_ (.A(\delay_counter[6] ),
    .X(_09967_));
 sg13g2_buf_1 _16059_ (.A(\delay_counter[4] ),
    .X(_09968_));
 sg13g2_buf_1 _16060_ (.A(\delay_counter[3] ),
    .X(_09969_));
 sg13g2_buf_1 _16061_ (.A(\delay_counter[0] ),
    .X(_09970_));
 sg13g2_buf_1 _16062_ (.A(\delay_counter[1] ),
    .X(_09971_));
 sg13g2_buf_1 _16063_ (.A(\delay_counter[2] ),
    .X(_09972_));
 sg13g2_nor3_1 _16064_ (.A(_09970_),
    .B(_09971_),
    .C(_09972_),
    .Y(_09973_));
 sg13g2_nor2b_1 _16065_ (.A(_09969_),
    .B_N(_09973_),
    .Y(_09974_));
 sg13g2_nand2b_1 _16066_ (.Y(_09975_),
    .B(_09974_),
    .A_N(_09968_));
 sg13g2_or2_1 _16067_ (.X(_09976_),
    .B(_09975_),
    .A(\delay_counter[5] ));
 sg13g2_buf_1 _16068_ (.A(_09976_),
    .X(_09977_));
 sg13g2_nor3_1 _16069_ (.A(_09966_),
    .B(_09967_),
    .C(_09977_),
    .Y(_09978_));
 sg13g2_nor2_1 _16070_ (.A(_09933_),
    .B(_09978_),
    .Y(_09979_));
 sg13g2_nand3_1 _16071_ (.B(_09962_),
    .C(_09979_),
    .A(net1274),
    .Y(_09980_));
 sg13g2_o21ai_1 _16072_ (.B1(_09980_),
    .Y(_09981_),
    .A1(_09933_),
    .A2(_09964_));
 sg13g2_nand2_1 _16073_ (.Y(_09982_),
    .A(net1194),
    .B(_09981_));
 sg13g2_o21ai_1 _16074_ (.B1(_09982_),
    .Y(_00010_),
    .A1(_09888_),
    .A2(_09921_));
 sg13g2_inv_1 _16075_ (.Y(_09983_),
    .A(_09888_));
 sg13g2_buf_1 _16076_ (.A(net1304),
    .X(_09984_));
 sg13g2_buf_1 _16077_ (.A(net1273),
    .X(_09985_));
 sg13g2_buf_2 _16078_ (.A(\mem.internal_data_ready ),
    .X(_09986_));
 sg13g2_buf_2 _16079_ (.A(\state[6] ),
    .X(_09987_));
 sg13g2_o21ai_1 _16080_ (.B1(_09987_),
    .Y(_09988_),
    .A1(_09986_),
    .A2(\mem.io_data_ready ));
 sg13g2_o21ai_1 _16081_ (.B1(_09931_),
    .Y(_09989_),
    .A1(_09903_),
    .A2(_09988_));
 sg13g2_buf_1 _16082_ (.A(\state[1] ),
    .X(_09990_));
 sg13g2_buf_2 _16083_ (.A(\mem.select ),
    .X(_09991_));
 sg13g2_o21ai_1 _16084_ (.B1(_09991_),
    .Y(_09992_),
    .A1(_09986_),
    .A2(\mem.io_data_ready ));
 sg13g2_nand3_1 _16085_ (.B(_09926_),
    .C(_09992_),
    .A(_09990_),
    .Y(_09993_));
 sg13g2_nand2b_1 _16086_ (.Y(_09994_),
    .B(_09993_),
    .A_N(_09989_));
 sg13g2_buf_1 _16087_ (.A(net1273),
    .X(_09995_));
 sg13g2_and4_1 _16088_ (.A(net1274),
    .B(net1192),
    .C(_09962_),
    .D(_09978_),
    .X(_09996_));
 sg13g2_a22oi_1 _16089_ (.Y(_09997_),
    .B1(_09996_),
    .B2(_00069_),
    .A2(_09994_),
    .A1(_09985_));
 sg13g2_o21ai_1 _16090_ (.B1(_09997_),
    .Y(_00009_),
    .A1(_09983_),
    .A2(_09921_));
 sg13g2_and2_1 _16091_ (.A(net1303),
    .B(_09925_),
    .X(_09998_));
 sg13g2_buf_1 _16092_ (.A(_09998_),
    .X(_09999_));
 sg13g2_nor2_1 _16093_ (.A(_09999_),
    .B(_09933_),
    .Y(_10000_));
 sg13g2_and4_1 _16094_ (.A(net1275),
    .B(_09890_),
    .C(_09891_),
    .D(_09895_),
    .X(_10001_));
 sg13g2_buf_1 _16095_ (.A(_10001_),
    .X(_10002_));
 sg13g2_nor3_1 _16096_ (.A(_10002_),
    .B(_09904_),
    .C(net859),
    .Y(_10003_));
 sg13g2_a21o_1 _16097_ (.A2(_10000_),
    .A1(\state[4] ),
    .B1(_10003_),
    .X(_00012_));
 sg13g2_nor2_2 _16098_ (.A(_09986_),
    .B(\mem.io_data_ready ),
    .Y(_10004_));
 sg13g2_nor2b_1 _16099_ (.A(_10004_),
    .B_N(_09991_),
    .Y(_10005_));
 sg13g2_buf_1 _16100_ (.A(\state[5] ),
    .X(_10006_));
 sg13g2_or2_1 _16101_ (.X(_10007_),
    .B(_10006_),
    .A(_09990_));
 sg13g2_buf_1 _16102_ (.A(_10007_),
    .X(_10008_));
 sg13g2_a21oi_1 _16103_ (.A1(_09987_),
    .A2(_10004_),
    .Y(_10009_),
    .B1(_10008_));
 sg13g2_nor2_1 _16104_ (.A(\state[4] ),
    .B(_09928_),
    .Y(_10010_));
 sg13g2_o21ai_1 _16105_ (.B1(_10010_),
    .Y(_10011_),
    .A1(_10005_),
    .A2(_10009_));
 sg13g2_a21oi_1 _16106_ (.A1(_09962_),
    .A2(_09978_),
    .Y(_10012_),
    .B1(_09935_));
 sg13g2_nor2_1 _16107_ (.A(_10011_),
    .B(_10012_),
    .Y(_10013_));
 sg13g2_buf_1 _16108_ (.A(\shift_reg[0] ),
    .X(_10014_));
 sg13g2_buf_1 _16109_ (.A(\shift_reg[2] ),
    .X(_10015_));
 sg13g2_buf_1 _16110_ (.A(\shift_reg[3] ),
    .X(_10016_));
 sg13g2_buf_1 _16111_ (.A(\shift_reg[6] ),
    .X(_10017_));
 sg13g2_inv_2 _16112_ (.Y(_10018_),
    .A(_10017_));
 sg13g2_nand4_1 _16113_ (.B(net1301),
    .C(_10016_),
    .A(_10014_),
    .Y(_10019_),
    .D(_10018_));
 sg13g2_or4_1 _16114_ (.A(\shift_reg[0] ),
    .B(\shift_reg[2] ),
    .C(\shift_reg[3] ),
    .D(_10018_),
    .X(_10020_));
 sg13g2_buf_1 _16115_ (.A(\shift_reg[1] ),
    .X(_10021_));
 sg13g2_buf_1 _16116_ (.A(\shift_reg[4] ),
    .X(_10022_));
 sg13g2_buf_1 _16117_ (.A(\shift_reg[5] ),
    .X(_10023_));
 sg13g2_buf_1 _16118_ (.A(\shift_reg[7] ),
    .X(_10024_));
 sg13g2_inv_2 _16119_ (.Y(_10025_),
    .A(_10024_));
 sg13g2_nand4_1 _16120_ (.B(_10022_),
    .C(net1298),
    .A(net1299),
    .Y(_10026_),
    .D(_10025_));
 sg13g2_a21oi_1 _16121_ (.A1(_10019_),
    .A2(_10020_),
    .Y(_10027_),
    .B1(_10026_));
 sg13g2_nor4_1 _16122_ (.A(_09927_),
    .B(_09933_),
    .C(_10013_),
    .D(_10027_),
    .Y(_10028_));
 sg13g2_and3_1 _16123_ (.X(_10029_),
    .A(net1273),
    .B(_10006_),
    .C(_10005_));
 sg13g2_buf_1 _16124_ (.A(_10029_),
    .X(_10030_));
 sg13g2_buf_1 _16125_ (.A(\mem.addr[7] ),
    .X(_10031_));
 sg13g2_nand2b_1 _16126_ (.Y(_10032_),
    .B(\mem.mem_internal.memory_type_data ),
    .A_N(net1297));
 sg13g2_buf_1 _16127_ (.A(\mem.addr[6] ),
    .X(_10033_));
 sg13g2_buf_2 _16128_ (.A(\mem.addr[5] ),
    .X(_10034_));
 sg13g2_xnor2_1 _16129_ (.Y(_10035_),
    .A(net1296),
    .B(_10034_));
 sg13g2_nor2_1 _16130_ (.A(_10032_),
    .B(_10035_),
    .Y(_10036_));
 sg13g2_and2_1 _16131_ (.A(_09991_),
    .B(_10036_),
    .X(_10037_));
 sg13g2_buf_1 _16132_ (.A(_10037_),
    .X(_10038_));
 sg13g2_buf_1 _16133_ (.A(_10038_),
    .X(_10039_));
 sg13g2_mux2_2 _16134_ (.A0(\mem.internal_data_out[4] ),
    .A1(\mem.io_data_out[4] ),
    .S(net558),
    .X(_10040_));
 sg13g2_mux2_2 _16135_ (.A0(\mem.internal_data_out[1] ),
    .A1(\mem.io_data_out[1] ),
    .S(net558),
    .X(_10041_));
 sg13g2_mux2_1 _16136_ (.A0(\mem.internal_data_out[7] ),
    .A1(\mem.io_data_out[7] ),
    .S(net558),
    .X(_10042_));
 sg13g2_inv_1 _16137_ (.Y(_10043_),
    .A(_10042_));
 sg13g2_mux2_2 _16138_ (.A0(\mem.internal_data_out[5] ),
    .A1(\mem.io_data_out[5] ),
    .S(net558),
    .X(_10044_));
 sg13g2_nand4_1 _16139_ (.B(_10041_),
    .C(_10043_),
    .A(_10040_),
    .Y(_10045_),
    .D(_10044_));
 sg13g2_mux2_1 _16140_ (.A0(\mem.internal_data_out[0] ),
    .A1(\mem.io_data_out[0] ),
    .S(_10039_),
    .X(_10046_));
 sg13g2_buf_1 _16141_ (.A(_10046_),
    .X(_10047_));
 sg13g2_mux2_1 _16142_ (.A0(\mem.internal_data_out[3] ),
    .A1(\mem.io_data_out[3] ),
    .S(net558),
    .X(_10048_));
 sg13g2_buf_1 _16143_ (.A(_10048_),
    .X(_10049_));
 sg13g2_nor2_1 _16144_ (.A(_10047_),
    .B(_10049_),
    .Y(_10050_));
 sg13g2_mux2_1 _16145_ (.A0(\mem.internal_data_out[2] ),
    .A1(\mem.io_data_out[2] ),
    .S(_10039_),
    .X(_10051_));
 sg13g2_buf_1 _16146_ (.A(_10051_),
    .X(_10052_));
 sg13g2_mux2_1 _16147_ (.A0(\mem.internal_data_out[6] ),
    .A1(\mem.io_data_out[6] ),
    .S(_10038_),
    .X(_10053_));
 sg13g2_buf_1 _16148_ (.A(_10053_),
    .X(_10054_));
 sg13g2_nor2b_1 _16149_ (.A(_10052_),
    .B_N(_10054_),
    .Y(_10055_));
 sg13g2_and2_1 _16150_ (.A(_10047_),
    .B(_10049_),
    .X(_10056_));
 sg13g2_nor2b_1 _16151_ (.A(_10054_),
    .B_N(_10052_),
    .Y(_10057_));
 sg13g2_a22oi_1 _16152_ (.Y(_10058_),
    .B1(_10056_),
    .B2(_10057_),
    .A2(_10055_),
    .A1(_10050_));
 sg13g2_nor2_1 _16153_ (.A(_10045_),
    .B(_10058_),
    .Y(_10059_));
 sg13g2_and2_1 _16154_ (.A(_09990_),
    .B(_10005_),
    .X(_10060_));
 sg13g2_buf_1 _16155_ (.A(_10060_),
    .X(_10061_));
 sg13g2_nand2_1 _16156_ (.Y(_10062_),
    .A(_09985_),
    .B(_10061_));
 sg13g2_nor2_1 _16157_ (.A(_10059_),
    .B(_10062_),
    .Y(_10063_));
 sg13g2_or3_1 _16158_ (.A(_10028_),
    .B(_10030_),
    .C(_10063_),
    .X(_00011_));
 sg13g2_buf_1 _16159_ (.A(_09999_),
    .X(_10064_));
 sg13g2_nor2_1 _16160_ (.A(_09935_),
    .B(_09962_),
    .Y(_10065_));
 sg13g2_buf_1 _16161_ (.A(_10065_),
    .X(_10066_));
 sg13g2_nor2_1 _16162_ (.A(_10066_),
    .B(_10011_),
    .Y(_10067_));
 sg13g2_o21ai_1 _16163_ (.B1(_09980_),
    .Y(_10068_),
    .A1(_09933_),
    .A2(_10067_));
 sg13g2_nand3_1 _16164_ (.B(_10027_),
    .C(_10068_),
    .A(net858),
    .Y(_10069_));
 sg13g2_buf_2 _16165_ (.A(net1273),
    .X(_10070_));
 sg13g2_buf_2 _16166_ (.A(_10070_),
    .X(_10071_));
 sg13g2_buf_1 _16167_ (.A(net782),
    .X(_10072_));
 sg13g2_nand3_1 _16168_ (.B(_10059_),
    .C(_10072_),
    .A(_10071_),
    .Y(_10073_));
 sg13g2_nand3_1 _16169_ (.B(_09992_),
    .C(_10000_),
    .A(_10006_),
    .Y(_10074_));
 sg13g2_nand3_1 _16170_ (.B(_10073_),
    .C(_10074_),
    .A(_10069_),
    .Y(_00013_));
 sg13g2_buf_1 _16171_ (.A(_09909_),
    .X(_10075_));
 sg13g2_nand2_1 _16172_ (.Y(_10076_),
    .A(net1272),
    .B(_09920_));
 sg13g2_o21ai_1 _16173_ (.B1(net1192),
    .Y(_10077_),
    .A1(_00069_),
    .A2(_09988_));
 sg13g2_a21oi_1 _16174_ (.A1(_09928_),
    .A2(_10000_),
    .Y(_10078_),
    .B1(_10077_));
 sg13g2_o21ai_1 _16175_ (.B1(_10078_),
    .Y(_10079_),
    .A1(_09905_),
    .A2(_10076_));
 sg13g2_a21o_1 _16176_ (.A2(_09996_),
    .A1(_09903_),
    .B1(_10079_),
    .X(_00008_));
 sg13g2_buf_1 _16177_ (.A(net859),
    .X(_10080_));
 sg13g2_nand3_1 _16178_ (.B(_10004_),
    .C(_10000_),
    .A(_09987_),
    .Y(_10081_));
 sg13g2_o21ai_1 _16179_ (.B1(_10081_),
    .Y(_00014_),
    .A1(net559),
    .A2(_10080_));
 sg13g2_nand2b_1 _16180_ (.Y(_10082_),
    .B(_00072_),
    .A_N(_09990_));
 sg13g2_o21ai_1 _16181_ (.B1(net1276),
    .Y(_10083_),
    .A1(_09909_),
    .A2(_10082_));
 sg13g2_buf_1 _16182_ (.A(_10083_),
    .X(_10084_));
 sg13g2_buf_1 _16183_ (.A(_10084_),
    .X(_10085_));
 sg13g2_buf_2 _16184_ (.A(\exec.pc[0] ),
    .X(_10086_));
 sg13g2_nor2_1 _16185_ (.A(_09909_),
    .B(_10006_),
    .Y(_10087_));
 sg13g2_buf_2 _16186_ (.A(_10087_),
    .X(_10088_));
 sg13g2_buf_1 _16187_ (.A(_10088_),
    .X(_10089_));
 sg13g2_nor2_1 _16188_ (.A(net487),
    .B(net856),
    .Y(_10090_));
 sg13g2_a21oi_1 _16189_ (.A1(_10086_),
    .A2(_10089_),
    .Y(_10091_),
    .B1(_10090_));
 sg13g2_buf_1 _16190_ (.A(\mem.addr[0] ),
    .X(_10092_));
 sg13g2_nand2_1 _16191_ (.Y(_10093_),
    .A(_10092_),
    .B(_10085_));
 sg13g2_o21ai_1 _16192_ (.B1(_10093_),
    .Y(_00015_),
    .A1(net780),
    .A2(_10091_));
 sg13g2_nand3_1 _16193_ (.B(_09700_),
    .C(_09706_),
    .A(_09668_),
    .Y(_10094_));
 sg13g2_buf_1 _16194_ (.A(_10094_),
    .X(_10095_));
 sg13g2_buf_8 _16195_ (.A(_10095_),
    .X(_10096_));
 sg13g2_buf_1 _16196_ (.A(net486),
    .X(_10097_));
 sg13g2_buf_2 _16197_ (.A(net473),
    .X(_10098_));
 sg13g2_buf_1 _16198_ (.A(\exec.pc[1] ),
    .X(_10099_));
 sg13g2_nand2b_1 _16199_ (.Y(_10100_),
    .B(_10088_),
    .A_N(_10099_));
 sg13g2_o21ai_1 _16200_ (.B1(_10100_),
    .Y(_10101_),
    .A1(net447),
    .A2(_10089_));
 sg13g2_buf_1 _16201_ (.A(\mem.addr[1] ),
    .X(_10102_));
 sg13g2_nand2_1 _16202_ (.Y(_10103_),
    .A(_10102_),
    .B(_10084_));
 sg13g2_o21ai_1 _16203_ (.B1(_10103_),
    .Y(_00016_),
    .A1(net780),
    .A2(_10101_));
 sg13g2_buf_1 _16204_ (.A(\exec.pc[2] ),
    .X(_10104_));
 sg13g2_nand2_1 _16205_ (.Y(_10105_),
    .A(_10104_),
    .B(_10088_));
 sg13g2_o21ai_1 _16206_ (.B1(_10105_),
    .Y(_10106_),
    .A1(_09807_),
    .A2(net856));
 sg13g2_buf_1 _16207_ (.A(\mem.addr[2] ),
    .X(_10107_));
 sg13g2_mux2_1 _16208_ (.A0(_10106_),
    .A1(net1293),
    .S(net780),
    .X(_00017_));
 sg13g2_buf_1 _16209_ (.A(\exec.pc[3] ),
    .X(_10108_));
 sg13g2_nand2_1 _16210_ (.Y(_10109_),
    .A(_10108_),
    .B(_10088_));
 sg13g2_o21ai_1 _16211_ (.B1(_10109_),
    .Y(_10110_),
    .A1(_09788_),
    .A2(net856));
 sg13g2_buf_1 _16212_ (.A(\mem.addr[3] ),
    .X(_10111_));
 sg13g2_buf_1 _16213_ (.A(_10111_),
    .X(_10112_));
 sg13g2_mux2_1 _16214_ (.A0(_10110_),
    .A1(net1271),
    .S(net780),
    .X(_00018_));
 sg13g2_buf_1 _16215_ (.A(\mem.addr[4] ),
    .X(_10113_));
 sg13g2_inv_2 _16216_ (.Y(_10114_),
    .A(_10113_));
 sg13g2_nand2_1 _16217_ (.Y(_10115_),
    .A(net563),
    .B(_09852_));
 sg13g2_a21oi_1 _16218_ (.A1(_09674_),
    .A2(_09857_),
    .Y(_10116_),
    .B1(_09862_));
 sg13g2_nand2_1 _16219_ (.Y(_10117_),
    .A(_10115_),
    .B(_10116_));
 sg13g2_buf_1 _16220_ (.A(_10117_),
    .X(_10118_));
 sg13g2_buf_1 _16221_ (.A(\exec.pc[4] ),
    .X(_10119_));
 sg13g2_nand2_1 _16222_ (.Y(_10120_),
    .A(_10119_),
    .B(_10088_));
 sg13g2_o21ai_1 _16223_ (.B1(_10120_),
    .Y(_10121_),
    .A1(_10118_),
    .A2(net856));
 sg13g2_nor2_1 _16224_ (.A(_10084_),
    .B(_10121_),
    .Y(_10122_));
 sg13g2_a21oi_1 _16225_ (.A1(_10114_),
    .A2(net780),
    .Y(_00019_),
    .B1(_10122_));
 sg13g2_inv_1 _16226_ (.Y(_10123_),
    .A(_10034_));
 sg13g2_nand2_1 _16227_ (.Y(_10124_),
    .A(net563),
    .B(_09833_));
 sg13g2_a21oi_1 _16228_ (.A1(_09674_),
    .A2(_09837_),
    .Y(_10125_),
    .B1(_09841_));
 sg13g2_nand2_1 _16229_ (.Y(_10126_),
    .A(_10124_),
    .B(_10125_));
 sg13g2_buf_1 _16230_ (.A(_10126_),
    .X(_10127_));
 sg13g2_buf_1 _16231_ (.A(net472),
    .X(_10128_));
 sg13g2_buf_1 _16232_ (.A(\exec.pc[5] ),
    .X(_10129_));
 sg13g2_nand2_1 _16233_ (.Y(_10130_),
    .A(_10129_),
    .B(_10088_));
 sg13g2_o21ai_1 _16234_ (.B1(_10130_),
    .Y(_10131_),
    .A1(_10128_),
    .A2(net856));
 sg13g2_nor2_1 _16235_ (.A(_10084_),
    .B(_10131_),
    .Y(_10132_));
 sg13g2_a21oi_1 _16236_ (.A1(_10123_),
    .A2(net780),
    .Y(_00020_),
    .B1(_10132_));
 sg13g2_buf_1 _16237_ (.A(\exec.pc[6] ),
    .X(_10133_));
 sg13g2_inv_1 _16238_ (.Y(_10134_),
    .A(net497));
 sg13g2_nor2_1 _16239_ (.A(_10134_),
    .B(net856),
    .Y(_10135_));
 sg13g2_a21oi_1 _16240_ (.A1(_10133_),
    .A2(net856),
    .Y(_10136_),
    .B1(_10135_));
 sg13g2_nand2_1 _16241_ (.Y(_10137_),
    .A(net1296),
    .B(_10084_));
 sg13g2_o21ai_1 _16242_ (.B1(_10137_),
    .Y(_00021_),
    .A1(_10085_),
    .A2(_10136_));
 sg13g2_inv_2 _16243_ (.Y(_10138_),
    .A(net474));
 sg13g2_nor2_1 _16244_ (.A(_10138_),
    .B(_10088_),
    .Y(_10139_));
 sg13g2_a21oi_1 _16245_ (.A1(\exec.pc[7] ),
    .A2(net856),
    .Y(_10140_),
    .B1(_10139_));
 sg13g2_nand2_1 _16246_ (.Y(_10141_),
    .A(net1297),
    .B(_10084_));
 sg13g2_o21ai_1 _16247_ (.B1(_10141_),
    .Y(_00022_),
    .A1(net780),
    .A2(_10140_));
 sg13g2_inv_1 _16248_ (.Y(_10142_),
    .A(_09906_));
 sg13g2_buf_1 _16249_ (.A(_10142_),
    .X(_10143_));
 sg13g2_buf_1 _16250_ (.A(net1270),
    .X(_10144_));
 sg13g2_nand2b_1 _16251_ (.Y(_10145_),
    .B(_09888_),
    .A_N(_00068_));
 sg13g2_nor2_1 _16252_ (.A(_09934_),
    .B(_09909_),
    .Y(_10146_));
 sg13g2_a21oi_1 _16253_ (.A1(_09909_),
    .A2(_09905_),
    .Y(_10147_),
    .B1(_10146_));
 sg13g2_o21ai_1 _16254_ (.B1(_10147_),
    .Y(_10148_),
    .A1(_09905_),
    .A2(_10145_));
 sg13g2_buf_1 _16255_ (.A(_10148_),
    .X(_10149_));
 sg13g2_or3_1 _16256_ (.A(net1191),
    .B(_10066_),
    .C(_10149_),
    .X(_10150_));
 sg13g2_buf_1 _16257_ (.A(_10150_),
    .X(_10151_));
 sg13g2_nand2_1 _16258_ (.Y(_10152_),
    .A(_09875_),
    .B(_09885_));
 sg13g2_o21ai_1 _16259_ (.B1(_09935_),
    .Y(_10153_),
    .A1(_10152_),
    .A2(net487));
 sg13g2_nor3_1 _16260_ (.A(_09970_),
    .B(_09935_),
    .C(net106),
    .Y(_10154_));
 sg13g2_a21oi_1 _16261_ (.A1(_09970_),
    .A2(_10151_),
    .Y(_10155_),
    .B1(_10154_));
 sg13g2_o21ai_1 _16262_ (.B1(_10155_),
    .Y(_00082_),
    .A1(net106),
    .A2(_10153_));
 sg13g2_nor2_1 _16263_ (.A(_09970_),
    .B(_09971_),
    .Y(_10156_));
 sg13g2_buf_1 _16264_ (.A(_10149_),
    .X(_10157_));
 sg13g2_nor3_1 _16265_ (.A(net1191),
    .B(_10066_),
    .C(net120),
    .Y(_10158_));
 sg13g2_buf_1 _16266_ (.A(_10158_),
    .X(_10159_));
 sg13g2_and2_1 _16267_ (.A(_09970_),
    .B(_09971_),
    .X(_10160_));
 sg13g2_a21oi_1 _16268_ (.A1(_10156_),
    .A2(net92),
    .Y(_10161_),
    .B1(_10160_));
 sg13g2_nor2_2 _16269_ (.A(net1274),
    .B(net106),
    .Y(_10162_));
 sg13g2_nand2_1 _16270_ (.Y(_10163_),
    .A(_09708_),
    .B(net487));
 sg13g2_a21oi_1 _16271_ (.A1(_09710_),
    .A2(_09750_),
    .Y(_10164_),
    .B1(_09769_));
 sg13g2_buf_1 _16272_ (.A(_10164_),
    .X(_10165_));
 sg13g2_nand2_1 _16273_ (.Y(_10166_),
    .A(net473),
    .B(net495));
 sg13g2_nand3_1 _16274_ (.B(_10163_),
    .C(_10166_),
    .A(_09887_),
    .Y(_10167_));
 sg13g2_a22oi_1 _16275_ (.Y(_10168_),
    .B1(_10162_),
    .B2(_10167_),
    .A2(_10151_),
    .A1(_09971_));
 sg13g2_o21ai_1 _16276_ (.B1(_10168_),
    .Y(_00083_),
    .A1(_09935_),
    .A2(_10161_));
 sg13g2_nor3_1 _16277_ (.A(net1274),
    .B(_10152_),
    .C(net106),
    .Y(_10169_));
 sg13g2_xnor2_1 _16278_ (.Y(_10170_),
    .A(_10163_),
    .B(_09807_));
 sg13g2_nand3_1 _16279_ (.B(_10156_),
    .C(_10159_),
    .A(_09972_),
    .Y(_10171_));
 sg13g2_o21ai_1 _16280_ (.B1(_10171_),
    .Y(_10172_),
    .A1(_09972_),
    .A2(_10156_));
 sg13g2_nor2_1 _16281_ (.A(_09972_),
    .B(net92),
    .Y(_10173_));
 sg13g2_a221oi_1 _16282_ (.B2(net1274),
    .C1(_10173_),
    .B1(_10172_),
    .A1(_10169_),
    .Y(_00084_),
    .A2(_10170_));
 sg13g2_nand2_1 _16283_ (.Y(_10174_),
    .A(net563),
    .B(_09777_));
 sg13g2_a21oi_1 _16284_ (.A1(_09701_),
    .A2(_09780_),
    .Y(_10175_),
    .B1(_09786_));
 sg13g2_nand2_1 _16285_ (.Y(_10176_),
    .A(_10174_),
    .B(_10175_));
 sg13g2_buf_1 _16286_ (.A(_10176_),
    .X(_10177_));
 sg13g2_buf_1 _16287_ (.A(net510),
    .X(_10178_));
 sg13g2_inv_1 _16288_ (.Y(_10179_),
    .A(_09796_));
 sg13g2_a21oi_1 _16289_ (.A1(_09674_),
    .A2(_09791_),
    .Y(_10180_),
    .B1(_09805_));
 sg13g2_o21ai_1 _16290_ (.B1(_10180_),
    .Y(_10181_),
    .A1(_09710_),
    .A2(_10179_));
 sg13g2_buf_2 _16291_ (.A(_10181_),
    .X(_10182_));
 sg13g2_buf_1 _16292_ (.A(_10182_),
    .X(_10183_));
 sg13g2_nor2_1 _16293_ (.A(_10163_),
    .B(net485),
    .Y(_10184_));
 sg13g2_xnor2_1 _16294_ (.Y(_10185_),
    .A(net494),
    .B(_10184_));
 sg13g2_nand3_1 _16295_ (.B(_09973_),
    .C(net92),
    .A(_09969_),
    .Y(_10186_));
 sg13g2_o21ai_1 _16296_ (.B1(_10186_),
    .Y(_10187_),
    .A1(_09969_),
    .A2(_09973_));
 sg13g2_nor2_1 _16297_ (.A(_09969_),
    .B(net92),
    .Y(_10188_));
 sg13g2_a221oi_1 _16298_ (.B2(net1274),
    .C1(_10188_),
    .B1(_10187_),
    .A1(_10169_),
    .Y(_00085_),
    .A2(_10185_));
 sg13g2_nor4_2 _16299_ (.A(_10176_),
    .B(_10095_),
    .C(_10164_),
    .Y(_10189_),
    .D(_10182_));
 sg13g2_buf_1 _16300_ (.A(_09864_),
    .X(_10190_));
 sg13g2_buf_1 _16301_ (.A(net493),
    .X(_10191_));
 sg13g2_xnor2_1 _16302_ (.Y(_10192_),
    .A(_10189_),
    .B(net484));
 sg13g2_nand3_1 _16303_ (.B(_09974_),
    .C(net92),
    .A(_09968_),
    .Y(_10193_));
 sg13g2_o21ai_1 _16304_ (.B1(_10193_),
    .Y(_10194_),
    .A1(_09968_),
    .A2(_09974_));
 sg13g2_nor2_1 _16305_ (.A(_09968_),
    .B(net92),
    .Y(_10195_));
 sg13g2_a221oi_1 _16306_ (.B2(_09965_),
    .C1(_10195_),
    .B1(_10194_),
    .A1(_10169_),
    .Y(_00086_),
    .A2(_10192_));
 sg13g2_and4_1 _16307_ (.A(_09708_),
    .B(_09771_),
    .C(_09809_),
    .D(_10117_),
    .X(_10196_));
 sg13g2_buf_1 _16308_ (.A(_10196_),
    .X(_10197_));
 sg13g2_nand2_1 _16309_ (.Y(_10198_),
    .A(net472),
    .B(_10197_));
 sg13g2_buf_1 _16310_ (.A(_09843_),
    .X(_10199_));
 sg13g2_nand4_1 _16311_ (.B(_09771_),
    .C(_09809_),
    .A(_09708_),
    .Y(_10200_),
    .D(_10117_));
 sg13g2_buf_1 _16312_ (.A(_10200_),
    .X(_10201_));
 sg13g2_nand2_1 _16313_ (.Y(_10202_),
    .A(net471),
    .B(_10201_));
 sg13g2_nand3_1 _16314_ (.B(_10198_),
    .C(_10202_),
    .A(_09887_),
    .Y(_10203_));
 sg13g2_nand2_1 _16315_ (.Y(_10204_),
    .A(\delay_counter[5] ),
    .B(_09975_));
 sg13g2_o21ai_1 _16316_ (.B1(_10204_),
    .Y(_10205_),
    .A1(_09977_),
    .A2(net106));
 sg13g2_and2_1 _16317_ (.A(\delay_counter[5] ),
    .B(net106),
    .X(_10206_));
 sg13g2_a221oi_1 _16318_ (.B2(_09965_),
    .C1(_10206_),
    .B1(_10205_),
    .A1(_10162_),
    .Y(_10207_),
    .A2(_10203_));
 sg13g2_inv_1 _16319_ (.Y(_00087_),
    .A(_10207_));
 sg13g2_nor2_1 _16320_ (.A(_09934_),
    .B(_10152_),
    .Y(_10208_));
 sg13g2_a22oi_1 _16321_ (.Y(_10209_),
    .B1(_10208_),
    .B2(_10198_),
    .A2(_09977_),
    .A1(_09934_));
 sg13g2_buf_1 _16322_ (.A(_10209_),
    .X(_10210_));
 sg13g2_buf_1 _16323_ (.A(net497),
    .X(_10211_));
 sg13g2_nand2_1 _16324_ (.Y(_10212_),
    .A(_09887_),
    .B(net483));
 sg13g2_xor2_1 _16325_ (.B(_10212_),
    .A(_10210_),
    .X(_10213_));
 sg13g2_nand3_1 _16326_ (.B(net92),
    .C(_10210_),
    .A(_09967_),
    .Y(_10214_));
 sg13g2_o21ai_1 _16327_ (.B1(_10214_),
    .Y(_10215_),
    .A1(_09967_),
    .A2(_10210_));
 sg13g2_nor2_1 _16328_ (.A(_09967_),
    .B(net92),
    .Y(_10216_));
 sg13g2_a221oi_1 _16329_ (.B2(net1274),
    .C1(_10216_),
    .B1(_10215_),
    .A1(_10162_),
    .Y(_00088_),
    .A2(_10213_));
 sg13g2_nor2_1 _16330_ (.A(_09934_),
    .B(_10212_),
    .Y(_10217_));
 sg13g2_a21oi_1 _16331_ (.A1(net1274),
    .A2(_09967_),
    .Y(_10218_),
    .B1(_10217_));
 sg13g2_nand2_1 _16332_ (.Y(_10219_),
    .A(_10210_),
    .B(_10218_));
 sg13g2_nor3_1 _16333_ (.A(_09966_),
    .B(net106),
    .C(_10219_),
    .Y(_10220_));
 sg13g2_a21oi_1 _16334_ (.A1(_09966_),
    .A2(_10219_),
    .Y(_10221_),
    .B1(_10220_));
 sg13g2_buf_1 _16335_ (.A(net474),
    .X(_10222_));
 sg13g2_nand2_1 _16336_ (.Y(_10223_),
    .A(_09887_),
    .B(net445));
 sg13g2_xor2_1 _16337_ (.B(_10223_),
    .A(_10219_),
    .X(_10224_));
 sg13g2_a22oi_1 _16338_ (.Y(_10225_),
    .B1(_10162_),
    .B2(_10224_),
    .A2(net106),
    .A1(_09966_));
 sg13g2_o21ai_1 _16339_ (.B1(_10225_),
    .Y(_00089_),
    .A1(_09935_),
    .A2(_10221_));
 sg13g2_buf_1 _16340_ (.A(_10070_),
    .X(_10226_));
 sg13g2_nand2_1 _16341_ (.Y(_10227_),
    .A(net855),
    .B(\mem.mem_internal.code_mem[0][0] ));
 sg13g2_nor2_1 _16342_ (.A(net1293),
    .B(net1271),
    .Y(_10228_));
 sg13g2_buf_2 _16343_ (.A(_10228_),
    .X(_10229_));
 sg13g2_nor2_2 _16344_ (.A(net1295),
    .B(net1294),
    .Y(_10230_));
 sg13g2_nand2_1 _16345_ (.Y(_10231_),
    .A(_10229_),
    .B(_10230_));
 sg13g2_buf_2 _16346_ (.A(_10231_),
    .X(_10232_));
 sg13g2_buf_2 _16347_ (.A(_10232_),
    .X(_10233_));
 sg13g2_nor2_1 _16348_ (.A(net1297),
    .B(net1296),
    .Y(_10234_));
 sg13g2_buf_1 _16349_ (.A(_10113_),
    .X(_10235_));
 sg13g2_buf_2 _16350_ (.A(\mem.mem_internal.write ),
    .X(_10236_));
 sg13g2_buf_1 _16351_ (.A(\mem.mem_internal.cycles[1] ),
    .X(_10237_));
 sg13g2_buf_1 _16352_ (.A(\mem.mem_internal.cycles[0] ),
    .X(_10238_));
 sg13g2_nor2b_1 _16353_ (.A(_10036_),
    .B_N(_09991_),
    .Y(_10239_));
 sg13g2_nand2_1 _16354_ (.Y(_10240_),
    .A(_09906_),
    .B(_10239_));
 sg13g2_nor3_1 _16355_ (.A(_10237_),
    .B(_10238_),
    .C(_10240_),
    .Y(_10241_));
 sg13g2_nand3b_1 _16356_ (.B(_10236_),
    .C(_10241_),
    .Y(_10242_),
    .A_N(\mem.mem_internal.memory_type_data ));
 sg13g2_buf_2 _16357_ (.A(_10242_),
    .X(_10243_));
 sg13g2_nor3_2 _16358_ (.A(_10235_),
    .B(_10034_),
    .C(_10243_),
    .Y(_10244_));
 sg13g2_nand2_1 _16359_ (.Y(_10245_),
    .A(_10234_),
    .B(_10244_));
 sg13g2_buf_2 _16360_ (.A(_10245_),
    .X(_10246_));
 sg13g2_buf_1 _16361_ (.A(_10246_),
    .X(_10247_));
 sg13g2_nor2_1 _16362_ (.A(net529),
    .B(net470),
    .Y(_10248_));
 sg13g2_buf_2 _16363_ (.A(_10248_),
    .X(_10249_));
 sg13g2_buf_1 _16364_ (.A(_10249_),
    .X(_10250_));
 sg13g2_buf_1 _16365_ (.A(_00023_),
    .X(_10251_));
 sg13g2_buf_1 _16366_ (.A(_10251_),
    .X(_10252_));
 sg13g2_buf_1 _16367_ (.A(net1268),
    .X(_10253_));
 sg13g2_nand2_1 _16368_ (.Y(_10254_),
    .A(_10253_),
    .B(net293));
 sg13g2_o21ai_1 _16369_ (.B1(_10254_),
    .Y(_00114_),
    .A1(_10227_),
    .A2(net293));
 sg13g2_nand2_1 _16370_ (.Y(_10255_),
    .A(_10071_),
    .B(\mem.mem_internal.code_mem[0][1] ));
 sg13g2_buf_1 _16371_ (.A(_00024_),
    .X(_10256_));
 sg13g2_buf_1 _16372_ (.A(_10256_),
    .X(_10257_));
 sg13g2_buf_1 _16373_ (.A(net1267),
    .X(_10258_));
 sg13g2_nand2_1 _16374_ (.Y(_10259_),
    .A(_10258_),
    .B(net293));
 sg13g2_o21ai_1 _16375_ (.B1(_10259_),
    .Y(_00115_),
    .A1(net293),
    .A2(_10255_));
 sg13g2_buf_1 _16376_ (.A(net1193),
    .X(_10260_));
 sg13g2_nand2_1 _16377_ (.Y(_10261_),
    .A(net854),
    .B(\mem.mem_internal.code_mem[0][2] ));
 sg13g2_buf_1 _16378_ (.A(_00025_),
    .X(_10262_));
 sg13g2_buf_1 _16379_ (.A(_10262_),
    .X(_10263_));
 sg13g2_buf_1 _16380_ (.A(net1266),
    .X(_10264_));
 sg13g2_nand2_1 _16381_ (.Y(_10265_),
    .A(_10264_),
    .B(_10249_));
 sg13g2_o21ai_1 _16382_ (.B1(_10265_),
    .Y(_00116_),
    .A1(net293),
    .A2(_10261_));
 sg13g2_nand2_1 _16383_ (.Y(_10266_),
    .A(net854),
    .B(\mem.mem_internal.code_mem[0][3] ));
 sg13g2_buf_1 _16384_ (.A(_00026_),
    .X(_10267_));
 sg13g2_buf_1 _16385_ (.A(_10267_),
    .X(_10268_));
 sg13g2_buf_1 _16386_ (.A(net1265),
    .X(_10269_));
 sg13g2_nand2_1 _16387_ (.Y(_10270_),
    .A(_10269_),
    .B(_10249_));
 sg13g2_o21ai_1 _16388_ (.B1(_10270_),
    .Y(_00117_),
    .A1(net293),
    .A2(_10266_));
 sg13g2_nand2_1 _16389_ (.Y(_10271_),
    .A(net854),
    .B(\mem.mem_internal.code_mem[0][4] ));
 sg13g2_buf_1 _16390_ (.A(_00027_),
    .X(_10272_));
 sg13g2_buf_1 _16391_ (.A(_10272_),
    .X(_10273_));
 sg13g2_buf_1 _16392_ (.A(net1264),
    .X(_10274_));
 sg13g2_nand2_1 _16393_ (.Y(_10275_),
    .A(_10274_),
    .B(_10249_));
 sg13g2_o21ai_1 _16394_ (.B1(_10275_),
    .Y(_00118_),
    .A1(_10250_),
    .A2(_10271_));
 sg13g2_nand2_1 _16395_ (.Y(_10276_),
    .A(net854),
    .B(\mem.mem_internal.code_mem[0][5] ));
 sg13g2_buf_1 _16396_ (.A(_00028_),
    .X(_10277_));
 sg13g2_buf_1 _16397_ (.A(_10277_),
    .X(_10278_));
 sg13g2_buf_1 _16398_ (.A(net1263),
    .X(_10279_));
 sg13g2_nand2_1 _16399_ (.Y(_10280_),
    .A(_10279_),
    .B(_10249_));
 sg13g2_o21ai_1 _16400_ (.B1(_10280_),
    .Y(_00119_),
    .A1(_10250_),
    .A2(_10276_));
 sg13g2_nand2_1 _16401_ (.Y(_10281_),
    .A(net854),
    .B(\mem.mem_internal.code_mem[0][6] ));
 sg13g2_buf_1 _16402_ (.A(_00029_),
    .X(_10282_));
 sg13g2_buf_1 _16403_ (.A(_10282_),
    .X(_10283_));
 sg13g2_buf_1 _16404_ (.A(net1262),
    .X(_10284_));
 sg13g2_nand2_1 _16405_ (.Y(_10285_),
    .A(_10284_),
    .B(_10249_));
 sg13g2_o21ai_1 _16406_ (.B1(_10285_),
    .Y(_00120_),
    .A1(net293),
    .A2(_10281_));
 sg13g2_nand2_1 _16407_ (.Y(_10286_),
    .A(net854),
    .B(\mem.mem_internal.code_mem[0][7] ));
 sg13g2_buf_1 _16408_ (.A(_00030_),
    .X(_10287_));
 sg13g2_buf_1 _16409_ (.A(_10287_),
    .X(_10288_));
 sg13g2_buf_1 _16410_ (.A(net1261),
    .X(_10289_));
 sg13g2_nand2_1 _16411_ (.Y(_10290_),
    .A(_10289_),
    .B(_10249_));
 sg13g2_o21ai_1 _16412_ (.B1(_10290_),
    .Y(_00121_),
    .A1(net293),
    .A2(_10286_));
 sg13g2_nand2_1 _16413_ (.Y(_10291_),
    .A(net855),
    .B(\mem.mem_internal.code_mem[100][0] ));
 sg13g2_nor2b_1 _16414_ (.A(_10111_),
    .B_N(net1293),
    .Y(_10292_));
 sg13g2_buf_1 _16415_ (.A(_10292_),
    .X(_10293_));
 sg13g2_nand2_1 _16416_ (.Y(_10294_),
    .A(_10230_),
    .B(_10293_));
 sg13g2_buf_2 _16417_ (.A(_10294_),
    .X(_10295_));
 sg13g2_buf_2 _16418_ (.A(_10295_),
    .X(_10296_));
 sg13g2_nor2b_1 _16419_ (.A(_10031_),
    .B_N(_10033_),
    .Y(_10297_));
 sg13g2_nor3_2 _16420_ (.A(_10235_),
    .B(_10123_),
    .C(_10243_),
    .Y(_10298_));
 sg13g2_nand2_1 _16421_ (.Y(_10299_),
    .A(_10297_),
    .B(_10298_));
 sg13g2_buf_2 _16422_ (.A(_10299_),
    .X(_10300_));
 sg13g2_buf_1 _16423_ (.A(_10300_),
    .X(_10301_));
 sg13g2_nor2_1 _16424_ (.A(net556),
    .B(net469),
    .Y(_10302_));
 sg13g2_buf_2 _16425_ (.A(_10302_),
    .X(_10303_));
 sg13g2_buf_1 _16426_ (.A(_10303_),
    .X(_10304_));
 sg13g2_nand2_1 _16427_ (.Y(_10305_),
    .A(net1190),
    .B(net292));
 sg13g2_o21ai_1 _16428_ (.B1(_10305_),
    .Y(_00122_),
    .A1(_10291_),
    .A2(net292));
 sg13g2_nand2_1 _16429_ (.Y(_10306_),
    .A(net854),
    .B(\mem.mem_internal.code_mem[100][1] ));
 sg13g2_nand2_1 _16430_ (.Y(_10307_),
    .A(net1189),
    .B(net292));
 sg13g2_o21ai_1 _16431_ (.B1(_10307_),
    .Y(_00123_),
    .A1(net292),
    .A2(_10306_));
 sg13g2_nand2_1 _16432_ (.Y(_10308_),
    .A(net854),
    .B(\mem.mem_internal.code_mem[100][2] ));
 sg13g2_nand2_1 _16433_ (.Y(_10309_),
    .A(net1188),
    .B(_10303_));
 sg13g2_o21ai_1 _16434_ (.B1(_10309_),
    .Y(_00124_),
    .A1(net292),
    .A2(_10308_));
 sg13g2_nand2_1 _16435_ (.Y(_10310_),
    .A(_10260_),
    .B(\mem.mem_internal.code_mem[100][3] ));
 sg13g2_nand2_1 _16436_ (.Y(_10311_),
    .A(net1187),
    .B(_10303_));
 sg13g2_o21ai_1 _16437_ (.B1(_10311_),
    .Y(_00125_),
    .A1(net292),
    .A2(_10310_));
 sg13g2_nand2_1 _16438_ (.Y(_10312_),
    .A(_10260_),
    .B(\mem.mem_internal.code_mem[100][4] ));
 sg13g2_nand2_1 _16439_ (.Y(_10313_),
    .A(net1186),
    .B(_10303_));
 sg13g2_o21ai_1 _16440_ (.B1(_10313_),
    .Y(_00126_),
    .A1(net292),
    .A2(_10312_));
 sg13g2_buf_1 _16441_ (.A(net1193),
    .X(_10314_));
 sg13g2_nand2_1 _16442_ (.Y(_10315_),
    .A(net853),
    .B(\mem.mem_internal.code_mem[100][5] ));
 sg13g2_nand2_1 _16443_ (.Y(_10316_),
    .A(net1185),
    .B(_10303_));
 sg13g2_o21ai_1 _16444_ (.B1(_10316_),
    .Y(_00127_),
    .A1(_10304_),
    .A2(_10315_));
 sg13g2_nand2_1 _16445_ (.Y(_10317_),
    .A(net853),
    .B(\mem.mem_internal.code_mem[100][6] ));
 sg13g2_nand2_1 _16446_ (.Y(_10318_),
    .A(net1184),
    .B(_10303_));
 sg13g2_o21ai_1 _16447_ (.B1(_10318_),
    .Y(_00128_),
    .A1(_10304_),
    .A2(_10317_));
 sg13g2_nand2_1 _16448_ (.Y(_10319_),
    .A(net853),
    .B(\mem.mem_internal.code_mem[100][7] ));
 sg13g2_nand2_1 _16449_ (.Y(_10320_),
    .A(net1183),
    .B(_10303_));
 sg13g2_o21ai_1 _16450_ (.B1(_10320_),
    .Y(_00129_),
    .A1(net292),
    .A2(_10319_));
 sg13g2_nand2_1 _16451_ (.Y(_10321_),
    .A(net855),
    .B(\mem.mem_internal.code_mem[101][0] ));
 sg13g2_nor2b_1 _16452_ (.A(net1294),
    .B_N(net1295),
    .Y(_10322_));
 sg13g2_buf_1 _16453_ (.A(_10322_),
    .X(_10323_));
 sg13g2_nand2_1 _16454_ (.Y(_10324_),
    .A(_10293_),
    .B(_10323_));
 sg13g2_buf_2 _16455_ (.A(_10324_),
    .X(_10325_));
 sg13g2_buf_2 _16456_ (.A(_10325_),
    .X(_10326_));
 sg13g2_nor2_1 _16457_ (.A(_10301_),
    .B(net555),
    .Y(_10327_));
 sg13g2_buf_2 _16458_ (.A(_10327_),
    .X(_10328_));
 sg13g2_buf_1 _16459_ (.A(_10328_),
    .X(_10329_));
 sg13g2_nand2_1 _16460_ (.Y(_10330_),
    .A(net1190),
    .B(net291));
 sg13g2_o21ai_1 _16461_ (.B1(_10330_),
    .Y(_00130_),
    .A1(_10321_),
    .A2(net291));
 sg13g2_nand2_1 _16462_ (.Y(_10331_),
    .A(net853),
    .B(\mem.mem_internal.code_mem[101][1] ));
 sg13g2_nand2_1 _16463_ (.Y(_10332_),
    .A(net1189),
    .B(net291));
 sg13g2_o21ai_1 _16464_ (.B1(_10332_),
    .Y(_00131_),
    .A1(net291),
    .A2(_10331_));
 sg13g2_nand2_1 _16465_ (.Y(_10333_),
    .A(net853),
    .B(\mem.mem_internal.code_mem[101][2] ));
 sg13g2_nand2_1 _16466_ (.Y(_10334_),
    .A(net1188),
    .B(_10328_));
 sg13g2_o21ai_1 _16467_ (.B1(_10334_),
    .Y(_00132_),
    .A1(net291),
    .A2(_10333_));
 sg13g2_nand2_1 _16468_ (.Y(_10335_),
    .A(_10314_),
    .B(\mem.mem_internal.code_mem[101][3] ));
 sg13g2_nand2_1 _16469_ (.Y(_10336_),
    .A(net1187),
    .B(_10328_));
 sg13g2_o21ai_1 _16470_ (.B1(_10336_),
    .Y(_00133_),
    .A1(net291),
    .A2(_10335_));
 sg13g2_nand2_1 _16471_ (.Y(_10337_),
    .A(_10314_),
    .B(\mem.mem_internal.code_mem[101][4] ));
 sg13g2_nand2_1 _16472_ (.Y(_10338_),
    .A(net1186),
    .B(_10328_));
 sg13g2_o21ai_1 _16473_ (.B1(_10338_),
    .Y(_00134_),
    .A1(net291),
    .A2(_10337_));
 sg13g2_nand2_1 _16474_ (.Y(_10339_),
    .A(net853),
    .B(\mem.mem_internal.code_mem[101][5] ));
 sg13g2_nand2_1 _16475_ (.Y(_10340_),
    .A(net1185),
    .B(_10328_));
 sg13g2_o21ai_1 _16476_ (.B1(_10340_),
    .Y(_00135_),
    .A1(_10329_),
    .A2(_10339_));
 sg13g2_nand2_1 _16477_ (.Y(_10341_),
    .A(net853),
    .B(\mem.mem_internal.code_mem[101][6] ));
 sg13g2_nand2_1 _16478_ (.Y(_10342_),
    .A(net1184),
    .B(_10328_));
 sg13g2_o21ai_1 _16479_ (.B1(_10342_),
    .Y(_00136_),
    .A1(_10329_),
    .A2(_10341_));
 sg13g2_nand2_1 _16480_ (.Y(_10343_),
    .A(net853),
    .B(\mem.mem_internal.code_mem[101][7] ));
 sg13g2_nand2_1 _16481_ (.Y(_10344_),
    .A(net1183),
    .B(_10328_));
 sg13g2_o21ai_1 _16482_ (.B1(_10344_),
    .Y(_00137_),
    .A1(net291),
    .A2(_10343_));
 sg13g2_nand2_1 _16483_ (.Y(_10345_),
    .A(net855),
    .B(\mem.mem_internal.code_mem[102][0] ));
 sg13g2_nor2b_1 _16484_ (.A(net1295),
    .B_N(net1294),
    .Y(_10346_));
 sg13g2_buf_1 _16485_ (.A(_10346_),
    .X(_10347_));
 sg13g2_nand2_1 _16486_ (.Y(_10348_),
    .A(_10293_),
    .B(_10347_));
 sg13g2_buf_1 _16487_ (.A(_10348_),
    .X(_10349_));
 sg13g2_buf_2 _16488_ (.A(net779),
    .X(_10350_));
 sg13g2_nor2_1 _16489_ (.A(net469),
    .B(net554),
    .Y(_10351_));
 sg13g2_buf_2 _16490_ (.A(_10351_),
    .X(_10352_));
 sg13g2_buf_1 _16491_ (.A(_10352_),
    .X(_10353_));
 sg13g2_nand2_1 _16492_ (.Y(_10354_),
    .A(net1190),
    .B(net290));
 sg13g2_o21ai_1 _16493_ (.B1(_10354_),
    .Y(_00138_),
    .A1(_10345_),
    .A2(net290));
 sg13g2_buf_1 _16494_ (.A(net1193),
    .X(_10355_));
 sg13g2_nand2_1 _16495_ (.Y(_10356_),
    .A(net852),
    .B(\mem.mem_internal.code_mem[102][1] ));
 sg13g2_nand2_1 _16496_ (.Y(_10357_),
    .A(net1189),
    .B(net290));
 sg13g2_o21ai_1 _16497_ (.B1(_10357_),
    .Y(_00139_),
    .A1(net290),
    .A2(_10356_));
 sg13g2_nand2_1 _16498_ (.Y(_10358_),
    .A(net852),
    .B(\mem.mem_internal.code_mem[102][2] ));
 sg13g2_nand2_1 _16499_ (.Y(_10359_),
    .A(net1188),
    .B(_10352_));
 sg13g2_o21ai_1 _16500_ (.B1(_10359_),
    .Y(_00140_),
    .A1(net290),
    .A2(_10358_));
 sg13g2_nand2_1 _16501_ (.Y(_10360_),
    .A(net852),
    .B(\mem.mem_internal.code_mem[102][3] ));
 sg13g2_nand2_1 _16502_ (.Y(_10361_),
    .A(net1187),
    .B(_10352_));
 sg13g2_o21ai_1 _16503_ (.B1(_10361_),
    .Y(_00141_),
    .A1(net290),
    .A2(_10360_));
 sg13g2_nand2_1 _16504_ (.Y(_10362_),
    .A(net852),
    .B(\mem.mem_internal.code_mem[102][4] ));
 sg13g2_nand2_1 _16505_ (.Y(_10363_),
    .A(net1186),
    .B(_10352_));
 sg13g2_o21ai_1 _16506_ (.B1(_10363_),
    .Y(_00142_),
    .A1(net290),
    .A2(_10362_));
 sg13g2_nand2_1 _16507_ (.Y(_10364_),
    .A(net852),
    .B(\mem.mem_internal.code_mem[102][5] ));
 sg13g2_nand2_1 _16508_ (.Y(_10365_),
    .A(net1185),
    .B(_10352_));
 sg13g2_o21ai_1 _16509_ (.B1(_10365_),
    .Y(_00143_),
    .A1(_10353_),
    .A2(_10364_));
 sg13g2_nand2_1 _16510_ (.Y(_10366_),
    .A(_10355_),
    .B(\mem.mem_internal.code_mem[102][6] ));
 sg13g2_nand2_1 _16511_ (.Y(_10367_),
    .A(net1184),
    .B(_10352_));
 sg13g2_o21ai_1 _16512_ (.B1(_10367_),
    .Y(_00144_),
    .A1(_10353_),
    .A2(_10366_));
 sg13g2_nand2_1 _16513_ (.Y(_10368_),
    .A(net852),
    .B(\mem.mem_internal.code_mem[102][7] ));
 sg13g2_nand2_1 _16514_ (.Y(_10369_),
    .A(net1183),
    .B(_10352_));
 sg13g2_o21ai_1 _16515_ (.B1(_10369_),
    .Y(_00145_),
    .A1(net290),
    .A2(_10368_));
 sg13g2_nand2_1 _16516_ (.Y(_10370_),
    .A(net855),
    .B(\mem.mem_internal.code_mem[103][0] ));
 sg13g2_nand3_1 _16517_ (.B(_10102_),
    .C(_10293_),
    .A(net1295),
    .Y(_10371_));
 sg13g2_buf_4 _16518_ (.X(_10372_),
    .A(_10371_));
 sg13g2_buf_2 _16519_ (.A(_10372_),
    .X(_10373_));
 sg13g2_nor2_1 _16520_ (.A(net469),
    .B(net553),
    .Y(_10374_));
 sg13g2_buf_2 _16521_ (.A(_10374_),
    .X(_10375_));
 sg13g2_buf_1 _16522_ (.A(_10375_),
    .X(_10376_));
 sg13g2_nand2_1 _16523_ (.Y(_10377_),
    .A(_10253_),
    .B(net289));
 sg13g2_o21ai_1 _16524_ (.B1(_10377_),
    .Y(_00146_),
    .A1(_10370_),
    .A2(net289));
 sg13g2_nand2_1 _16525_ (.Y(_10378_),
    .A(net852),
    .B(\mem.mem_internal.code_mem[103][1] ));
 sg13g2_nand2_1 _16526_ (.Y(_10379_),
    .A(_10258_),
    .B(net289));
 sg13g2_o21ai_1 _16527_ (.B1(_10379_),
    .Y(_00147_),
    .A1(net289),
    .A2(_10378_));
 sg13g2_nand2_1 _16528_ (.Y(_10380_),
    .A(net852),
    .B(\mem.mem_internal.code_mem[103][2] ));
 sg13g2_nand2_1 _16529_ (.Y(_10381_),
    .A(_10264_),
    .B(_10375_));
 sg13g2_o21ai_1 _16530_ (.B1(_10381_),
    .Y(_00148_),
    .A1(net289),
    .A2(_10380_));
 sg13g2_nand2_1 _16531_ (.Y(_10382_),
    .A(_10355_),
    .B(\mem.mem_internal.code_mem[103][3] ));
 sg13g2_nand2_1 _16532_ (.Y(_10383_),
    .A(_10269_),
    .B(_10375_));
 sg13g2_o21ai_1 _16533_ (.B1(_10383_),
    .Y(_00149_),
    .A1(net289),
    .A2(_10382_));
 sg13g2_buf_1 _16534_ (.A(net1193),
    .X(_10384_));
 sg13g2_nand2_1 _16535_ (.Y(_10385_),
    .A(_10384_),
    .B(\mem.mem_internal.code_mem[103][4] ));
 sg13g2_nand2_1 _16536_ (.Y(_10386_),
    .A(_10274_),
    .B(_10375_));
 sg13g2_o21ai_1 _16537_ (.B1(_10386_),
    .Y(_00150_),
    .A1(net289),
    .A2(_10385_));
 sg13g2_nand2_1 _16538_ (.Y(_10387_),
    .A(net851),
    .B(\mem.mem_internal.code_mem[103][5] ));
 sg13g2_nand2_1 _16539_ (.Y(_10388_),
    .A(_10279_),
    .B(_10375_));
 sg13g2_o21ai_1 _16540_ (.B1(_10388_),
    .Y(_00151_),
    .A1(_10376_),
    .A2(_10387_));
 sg13g2_nand2_1 _16541_ (.Y(_10389_),
    .A(_10384_),
    .B(\mem.mem_internal.code_mem[103][6] ));
 sg13g2_nand2_1 _16542_ (.Y(_10390_),
    .A(_10284_),
    .B(_10375_));
 sg13g2_o21ai_1 _16543_ (.B1(_10390_),
    .Y(_00152_),
    .A1(_10376_),
    .A2(_10389_));
 sg13g2_nand2_1 _16544_ (.Y(_10391_),
    .A(net851),
    .B(\mem.mem_internal.code_mem[103][7] ));
 sg13g2_nand2_1 _16545_ (.Y(_10392_),
    .A(_10289_),
    .B(_10375_));
 sg13g2_o21ai_1 _16546_ (.B1(_10392_),
    .Y(_00153_),
    .A1(net289),
    .A2(_10391_));
 sg13g2_nand2_1 _16547_ (.Y(_10393_),
    .A(net855),
    .B(\mem.mem_internal.code_mem[104][0] ));
 sg13g2_nor2b_1 _16548_ (.A(net1293),
    .B_N(_10111_),
    .Y(_10394_));
 sg13g2_buf_2 _16549_ (.A(_10394_),
    .X(_10395_));
 sg13g2_nand2_1 _16550_ (.Y(_10396_),
    .A(_10230_),
    .B(_10395_));
 sg13g2_buf_2 _16551_ (.A(_10396_),
    .X(_10397_));
 sg13g2_buf_1 _16552_ (.A(net778),
    .X(_10398_));
 sg13g2_nor2_1 _16553_ (.A(net469),
    .B(net552),
    .Y(_10399_));
 sg13g2_buf_2 _16554_ (.A(_10399_),
    .X(_10400_));
 sg13g2_buf_1 _16555_ (.A(_10400_),
    .X(_10401_));
 sg13g2_nand2_1 _16556_ (.Y(_10402_),
    .A(net1190),
    .B(net288));
 sg13g2_o21ai_1 _16557_ (.B1(_10402_),
    .Y(_00154_),
    .A1(_10393_),
    .A2(net288));
 sg13g2_nand2_1 _16558_ (.Y(_10403_),
    .A(net851),
    .B(\mem.mem_internal.code_mem[104][1] ));
 sg13g2_nand2_1 _16559_ (.Y(_10404_),
    .A(net1189),
    .B(net288));
 sg13g2_o21ai_1 _16560_ (.B1(_10404_),
    .Y(_00155_),
    .A1(net288),
    .A2(_10403_));
 sg13g2_nand2_1 _16561_ (.Y(_10405_),
    .A(net851),
    .B(\mem.mem_internal.code_mem[104][2] ));
 sg13g2_nand2_1 _16562_ (.Y(_10406_),
    .A(net1188),
    .B(_10400_));
 sg13g2_o21ai_1 _16563_ (.B1(_10406_),
    .Y(_00156_),
    .A1(net288),
    .A2(_10405_));
 sg13g2_nand2_1 _16564_ (.Y(_10407_),
    .A(net851),
    .B(\mem.mem_internal.code_mem[104][3] ));
 sg13g2_nand2_1 _16565_ (.Y(_10408_),
    .A(net1187),
    .B(_10400_));
 sg13g2_o21ai_1 _16566_ (.B1(_10408_),
    .Y(_00157_),
    .A1(net288),
    .A2(_10407_));
 sg13g2_nand2_1 _16567_ (.Y(_10409_),
    .A(net851),
    .B(\mem.mem_internal.code_mem[104][4] ));
 sg13g2_nand2_1 _16568_ (.Y(_10410_),
    .A(net1186),
    .B(_10400_));
 sg13g2_o21ai_1 _16569_ (.B1(_10410_),
    .Y(_00158_),
    .A1(_10401_),
    .A2(_10409_));
 sg13g2_nand2_1 _16570_ (.Y(_10411_),
    .A(net851),
    .B(\mem.mem_internal.code_mem[104][5] ));
 sg13g2_nand2_1 _16571_ (.Y(_10412_),
    .A(net1185),
    .B(_10400_));
 sg13g2_o21ai_1 _16572_ (.B1(_10412_),
    .Y(_00159_),
    .A1(_10401_),
    .A2(_10411_));
 sg13g2_nand2_1 _16573_ (.Y(_10413_),
    .A(net851),
    .B(\mem.mem_internal.code_mem[104][6] ));
 sg13g2_nand2_1 _16574_ (.Y(_10414_),
    .A(net1184),
    .B(_10400_));
 sg13g2_o21ai_1 _16575_ (.B1(_10414_),
    .Y(_00160_),
    .A1(net288),
    .A2(_10413_));
 sg13g2_buf_2 _16576_ (.A(net1276),
    .X(_10415_));
 sg13g2_buf_1 _16577_ (.A(_10415_),
    .X(_10416_));
 sg13g2_buf_1 _16578_ (.A(_10416_),
    .X(_10417_));
 sg13g2_nand2_1 _16579_ (.Y(_10418_),
    .A(_10417_),
    .B(\mem.mem_internal.code_mem[104][7] ));
 sg13g2_nand2_1 _16580_ (.Y(_10419_),
    .A(net1183),
    .B(_10400_));
 sg13g2_o21ai_1 _16581_ (.B1(_10419_),
    .Y(_00161_),
    .A1(net288),
    .A2(_10418_));
 sg13g2_nand2_1 _16582_ (.Y(_10420_),
    .A(net855),
    .B(\mem.mem_internal.code_mem[105][0] ));
 sg13g2_nand2_1 _16583_ (.Y(_10421_),
    .A(_10323_),
    .B(_10395_));
 sg13g2_buf_4 _16584_ (.X(_10422_),
    .A(_10421_));
 sg13g2_buf_2 _16585_ (.A(_10422_),
    .X(_10423_));
 sg13g2_nor2_1 _16586_ (.A(net469),
    .B(net551),
    .Y(_10424_));
 sg13g2_buf_2 _16587_ (.A(_10424_),
    .X(_10425_));
 sg13g2_buf_1 _16588_ (.A(_10425_),
    .X(_10426_));
 sg13g2_nand2_1 _16589_ (.Y(_10427_),
    .A(net1190),
    .B(net287));
 sg13g2_o21ai_1 _16590_ (.B1(_10427_),
    .Y(_00162_),
    .A1(_10420_),
    .A2(net287));
 sg13g2_nand2_1 _16591_ (.Y(_10428_),
    .A(net777),
    .B(\mem.mem_internal.code_mem[105][1] ));
 sg13g2_nand2_1 _16592_ (.Y(_10429_),
    .A(net1189),
    .B(net287));
 sg13g2_o21ai_1 _16593_ (.B1(_10429_),
    .Y(_00163_),
    .A1(net287),
    .A2(_10428_));
 sg13g2_nand2_1 _16594_ (.Y(_10430_),
    .A(net777),
    .B(\mem.mem_internal.code_mem[105][2] ));
 sg13g2_nand2_1 _16595_ (.Y(_10431_),
    .A(net1188),
    .B(_10425_));
 sg13g2_o21ai_1 _16596_ (.B1(_10431_),
    .Y(_00164_),
    .A1(net287),
    .A2(_10430_));
 sg13g2_nand2_1 _16597_ (.Y(_10432_),
    .A(net777),
    .B(\mem.mem_internal.code_mem[105][3] ));
 sg13g2_nand2_1 _16598_ (.Y(_10433_),
    .A(net1187),
    .B(_10425_));
 sg13g2_o21ai_1 _16599_ (.B1(_10433_),
    .Y(_00165_),
    .A1(net287),
    .A2(_10432_));
 sg13g2_nand2_1 _16600_ (.Y(_10434_),
    .A(net777),
    .B(\mem.mem_internal.code_mem[105][4] ));
 sg13g2_nand2_1 _16601_ (.Y(_10435_),
    .A(net1186),
    .B(_10425_));
 sg13g2_o21ai_1 _16602_ (.B1(_10435_),
    .Y(_00166_),
    .A1(net287),
    .A2(_10434_));
 sg13g2_nand2_1 _16603_ (.Y(_10436_),
    .A(net777),
    .B(\mem.mem_internal.code_mem[105][5] ));
 sg13g2_nand2_1 _16604_ (.Y(_10437_),
    .A(net1185),
    .B(_10425_));
 sg13g2_o21ai_1 _16605_ (.B1(_10437_),
    .Y(_00167_),
    .A1(net287),
    .A2(_10436_));
 sg13g2_nand2_1 _16606_ (.Y(_10438_),
    .A(net777),
    .B(\mem.mem_internal.code_mem[105][6] ));
 sg13g2_nand2_1 _16607_ (.Y(_10439_),
    .A(net1184),
    .B(_10425_));
 sg13g2_o21ai_1 _16608_ (.B1(_10439_),
    .Y(_00168_),
    .A1(_10426_),
    .A2(_10438_));
 sg13g2_nand2_1 _16609_ (.Y(_10440_),
    .A(_10417_),
    .B(\mem.mem_internal.code_mem[105][7] ));
 sg13g2_nand2_1 _16610_ (.Y(_10441_),
    .A(net1183),
    .B(_10425_));
 sg13g2_o21ai_1 _16611_ (.B1(_10441_),
    .Y(_00169_),
    .A1(_10426_),
    .A2(_10440_));
 sg13g2_nand2_1 _16612_ (.Y(_10442_),
    .A(net855),
    .B(\mem.mem_internal.code_mem[106][0] ));
 sg13g2_nand2_1 _16613_ (.Y(_10443_),
    .A(_10347_),
    .B(_10395_));
 sg13g2_buf_4 _16614_ (.X(_10444_),
    .A(_10443_));
 sg13g2_buf_1 _16615_ (.A(_10444_),
    .X(_10445_));
 sg13g2_nor2_1 _16616_ (.A(net469),
    .B(net550),
    .Y(_10446_));
 sg13g2_buf_2 _16617_ (.A(_10446_),
    .X(_10447_));
 sg13g2_buf_1 _16618_ (.A(_10447_),
    .X(_10448_));
 sg13g2_nand2_1 _16619_ (.Y(_10449_),
    .A(net1190),
    .B(net286));
 sg13g2_o21ai_1 _16620_ (.B1(_10449_),
    .Y(_00170_),
    .A1(_10442_),
    .A2(net286));
 sg13g2_nand2_1 _16621_ (.Y(_10450_),
    .A(net777),
    .B(\mem.mem_internal.code_mem[106][1] ));
 sg13g2_nand2_1 _16622_ (.Y(_10451_),
    .A(net1189),
    .B(net286));
 sg13g2_o21ai_1 _16623_ (.B1(_10451_),
    .Y(_00171_),
    .A1(net286),
    .A2(_10450_));
 sg13g2_nand2_1 _16624_ (.Y(_10452_),
    .A(net777),
    .B(\mem.mem_internal.code_mem[106][2] ));
 sg13g2_nand2_1 _16625_ (.Y(_10453_),
    .A(net1188),
    .B(_10447_));
 sg13g2_o21ai_1 _16626_ (.B1(_10453_),
    .Y(_00172_),
    .A1(net286),
    .A2(_10452_));
 sg13g2_buf_1 _16627_ (.A(_10416_),
    .X(_10454_));
 sg13g2_nand2_1 _16628_ (.Y(_10455_),
    .A(_10454_),
    .B(\mem.mem_internal.code_mem[106][3] ));
 sg13g2_nand2_1 _16629_ (.Y(_10456_),
    .A(net1187),
    .B(_10447_));
 sg13g2_o21ai_1 _16630_ (.B1(_10456_),
    .Y(_00173_),
    .A1(net286),
    .A2(_10455_));
 sg13g2_nand2_1 _16631_ (.Y(_10457_),
    .A(net776),
    .B(\mem.mem_internal.code_mem[106][4] ));
 sg13g2_nand2_1 _16632_ (.Y(_10458_),
    .A(net1186),
    .B(_10447_));
 sg13g2_o21ai_1 _16633_ (.B1(_10458_),
    .Y(_00174_),
    .A1(net286),
    .A2(_10457_));
 sg13g2_nand2_1 _16634_ (.Y(_10459_),
    .A(net776),
    .B(\mem.mem_internal.code_mem[106][5] ));
 sg13g2_nand2_1 _16635_ (.Y(_10460_),
    .A(net1185),
    .B(_10447_));
 sg13g2_o21ai_1 _16636_ (.B1(_10460_),
    .Y(_00175_),
    .A1(net286),
    .A2(_10459_));
 sg13g2_nand2_1 _16637_ (.Y(_10461_),
    .A(net776),
    .B(\mem.mem_internal.code_mem[106][6] ));
 sg13g2_nand2_1 _16638_ (.Y(_10462_),
    .A(net1184),
    .B(_10447_));
 sg13g2_o21ai_1 _16639_ (.B1(_10462_),
    .Y(_00176_),
    .A1(_10448_),
    .A2(_10461_));
 sg13g2_nand2_1 _16640_ (.Y(_10463_),
    .A(net776),
    .B(\mem.mem_internal.code_mem[106][7] ));
 sg13g2_nand2_1 _16641_ (.Y(_10464_),
    .A(net1183),
    .B(_10447_));
 sg13g2_o21ai_1 _16642_ (.B1(_10464_),
    .Y(_00177_),
    .A1(_10448_),
    .A2(_10463_));
 sg13g2_nand2_1 _16643_ (.Y(_10465_),
    .A(_10226_),
    .B(\mem.mem_internal.code_mem[107][0] ));
 sg13g2_nand3_1 _16644_ (.B(net1294),
    .C(_10395_),
    .A(net1295),
    .Y(_10466_));
 sg13g2_buf_1 _16645_ (.A(_10466_),
    .X(_10467_));
 sg13g2_buf_2 _16646_ (.A(net775),
    .X(_10468_));
 sg13g2_nor2_1 _16647_ (.A(net469),
    .B(net549),
    .Y(_10469_));
 sg13g2_buf_2 _16648_ (.A(_10469_),
    .X(_10470_));
 sg13g2_buf_1 _16649_ (.A(_10470_),
    .X(_10471_));
 sg13g2_nand2_1 _16650_ (.Y(_10472_),
    .A(net1190),
    .B(net285));
 sg13g2_o21ai_1 _16651_ (.B1(_10472_),
    .Y(_00178_),
    .A1(_10465_),
    .A2(net285));
 sg13g2_nand2_1 _16652_ (.Y(_10473_),
    .A(net776),
    .B(\mem.mem_internal.code_mem[107][1] ));
 sg13g2_nand2_1 _16653_ (.Y(_10474_),
    .A(net1189),
    .B(net285));
 sg13g2_o21ai_1 _16654_ (.B1(_10474_),
    .Y(_00179_),
    .A1(net285),
    .A2(_10473_));
 sg13g2_nand2_1 _16655_ (.Y(_10475_),
    .A(net776),
    .B(\mem.mem_internal.code_mem[107][2] ));
 sg13g2_nand2_1 _16656_ (.Y(_10476_),
    .A(net1188),
    .B(_10470_));
 sg13g2_o21ai_1 _16657_ (.B1(_10476_),
    .Y(_00180_),
    .A1(net285),
    .A2(_10475_));
 sg13g2_nand2_1 _16658_ (.Y(_10477_),
    .A(_10454_),
    .B(\mem.mem_internal.code_mem[107][3] ));
 sg13g2_nand2_1 _16659_ (.Y(_10478_),
    .A(net1187),
    .B(_10470_));
 sg13g2_o21ai_1 _16660_ (.B1(_10478_),
    .Y(_00181_),
    .A1(net285),
    .A2(_10477_));
 sg13g2_nand2_1 _16661_ (.Y(_10479_),
    .A(net776),
    .B(\mem.mem_internal.code_mem[107][4] ));
 sg13g2_nand2_1 _16662_ (.Y(_10480_),
    .A(net1186),
    .B(_10470_));
 sg13g2_o21ai_1 _16663_ (.B1(_10480_),
    .Y(_00182_),
    .A1(net285),
    .A2(_10479_));
 sg13g2_nand2_1 _16664_ (.Y(_10481_),
    .A(net776),
    .B(\mem.mem_internal.code_mem[107][5] ));
 sg13g2_nand2_1 _16665_ (.Y(_10482_),
    .A(net1185),
    .B(_10470_));
 sg13g2_o21ai_1 _16666_ (.B1(_10482_),
    .Y(_00183_),
    .A1(net285),
    .A2(_10481_));
 sg13g2_buf_1 _16667_ (.A(_10416_),
    .X(_10483_));
 sg13g2_nand2_1 _16668_ (.Y(_10484_),
    .A(net774),
    .B(\mem.mem_internal.code_mem[107][6] ));
 sg13g2_nand2_1 _16669_ (.Y(_10485_),
    .A(net1184),
    .B(_10470_));
 sg13g2_o21ai_1 _16670_ (.B1(_10485_),
    .Y(_00184_),
    .A1(_10471_),
    .A2(_10484_));
 sg13g2_nand2_1 _16671_ (.Y(_10486_),
    .A(net774),
    .B(\mem.mem_internal.code_mem[107][7] ));
 sg13g2_nand2_1 _16672_ (.Y(_10487_),
    .A(net1183),
    .B(_10470_));
 sg13g2_o21ai_1 _16673_ (.B1(_10487_),
    .Y(_00185_),
    .A1(_10471_),
    .A2(_10486_));
 sg13g2_buf_1 _16674_ (.A(_10070_),
    .X(_10488_));
 sg13g2_nand2_1 _16675_ (.Y(_10489_),
    .A(net850),
    .B(\mem.mem_internal.code_mem[108][0] ));
 sg13g2_nand3_1 _16676_ (.B(net1271),
    .C(_10230_),
    .A(net1293),
    .Y(_10490_));
 sg13g2_buf_2 _16677_ (.A(_10490_),
    .X(_10491_));
 sg13g2_buf_1 _16678_ (.A(_10491_),
    .X(_10492_));
 sg13g2_nor2_1 _16679_ (.A(net469),
    .B(net773),
    .Y(_10493_));
 sg13g2_buf_2 _16680_ (.A(_10493_),
    .X(_10494_));
 sg13g2_buf_1 _16681_ (.A(_10494_),
    .X(_10495_));
 sg13g2_nand2_1 _16682_ (.Y(_10496_),
    .A(net1190),
    .B(net284));
 sg13g2_o21ai_1 _16683_ (.B1(_10496_),
    .Y(_00186_),
    .A1(_10489_),
    .A2(net284));
 sg13g2_nand2_1 _16684_ (.Y(_10497_),
    .A(net774),
    .B(\mem.mem_internal.code_mem[108][1] ));
 sg13g2_nand2_1 _16685_ (.Y(_10498_),
    .A(net1189),
    .B(net284));
 sg13g2_o21ai_1 _16686_ (.B1(_10498_),
    .Y(_00187_),
    .A1(net284),
    .A2(_10497_));
 sg13g2_nand2_1 _16687_ (.Y(_10499_),
    .A(_10483_),
    .B(\mem.mem_internal.code_mem[108][2] ));
 sg13g2_nand2_1 _16688_ (.Y(_10500_),
    .A(net1188),
    .B(_10494_));
 sg13g2_o21ai_1 _16689_ (.B1(_10500_),
    .Y(_00188_),
    .A1(net284),
    .A2(_10499_));
 sg13g2_nand2_1 _16690_ (.Y(_10501_),
    .A(_10483_),
    .B(\mem.mem_internal.code_mem[108][3] ));
 sg13g2_nand2_1 _16691_ (.Y(_10502_),
    .A(net1187),
    .B(_10494_));
 sg13g2_o21ai_1 _16692_ (.B1(_10502_),
    .Y(_00189_),
    .A1(net284),
    .A2(_10501_));
 sg13g2_nand2_1 _16693_ (.Y(_10503_),
    .A(net774),
    .B(\mem.mem_internal.code_mem[108][4] ));
 sg13g2_nand2_1 _16694_ (.Y(_10504_),
    .A(net1186),
    .B(_10494_));
 sg13g2_o21ai_1 _16695_ (.B1(_10504_),
    .Y(_00190_),
    .A1(net284),
    .A2(_10503_));
 sg13g2_nand2_1 _16696_ (.Y(_10505_),
    .A(net774),
    .B(\mem.mem_internal.code_mem[108][5] ));
 sg13g2_nand2_1 _16697_ (.Y(_10506_),
    .A(net1185),
    .B(_10494_));
 sg13g2_o21ai_1 _16698_ (.B1(_10506_),
    .Y(_00191_),
    .A1(net284),
    .A2(_10505_));
 sg13g2_nand2_1 _16699_ (.Y(_10507_),
    .A(net774),
    .B(\mem.mem_internal.code_mem[108][6] ));
 sg13g2_nand2_1 _16700_ (.Y(_10508_),
    .A(net1184),
    .B(_10494_));
 sg13g2_o21ai_1 _16701_ (.B1(_10508_),
    .Y(_00192_),
    .A1(_10495_),
    .A2(_10507_));
 sg13g2_nand2_1 _16702_ (.Y(_10509_),
    .A(net774),
    .B(\mem.mem_internal.code_mem[108][7] ));
 sg13g2_nand2_1 _16703_ (.Y(_10510_),
    .A(net1183),
    .B(_10494_));
 sg13g2_o21ai_1 _16704_ (.B1(_10510_),
    .Y(_00193_),
    .A1(_10495_),
    .A2(_10509_));
 sg13g2_nand2_1 _16705_ (.Y(_10511_),
    .A(net850),
    .B(\mem.mem_internal.code_mem[109][0] ));
 sg13g2_nand3_1 _16706_ (.B(_10112_),
    .C(_10323_),
    .A(net1293),
    .Y(_10512_));
 sg13g2_buf_2 _16707_ (.A(_10512_),
    .X(_10513_));
 sg13g2_buf_1 _16708_ (.A(_10513_),
    .X(_10514_));
 sg13g2_nor2_1 _16709_ (.A(_10300_),
    .B(net548),
    .Y(_10515_));
 sg13g2_buf_2 _16710_ (.A(_10515_),
    .X(_10516_));
 sg13g2_buf_1 _16711_ (.A(_10516_),
    .X(_10517_));
 sg13g2_buf_1 _16712_ (.A(net1268),
    .X(_10518_));
 sg13g2_nand2_1 _16713_ (.Y(_10519_),
    .A(net1182),
    .B(net399));
 sg13g2_o21ai_1 _16714_ (.B1(_10519_),
    .Y(_00194_),
    .A1(_10511_),
    .A2(net399));
 sg13g2_nand2_1 _16715_ (.Y(_10520_),
    .A(net774),
    .B(\mem.mem_internal.code_mem[109][1] ));
 sg13g2_buf_1 _16716_ (.A(net1267),
    .X(_10521_));
 sg13g2_nand2_1 _16717_ (.Y(_10522_),
    .A(net1181),
    .B(net399));
 sg13g2_o21ai_1 _16718_ (.B1(_10522_),
    .Y(_00195_),
    .A1(_10517_),
    .A2(_10520_));
 sg13g2_buf_1 _16719_ (.A(_10416_),
    .X(_10523_));
 sg13g2_nand2_1 _16720_ (.Y(_10524_),
    .A(net772),
    .B(\mem.mem_internal.code_mem[109][2] ));
 sg13g2_buf_1 _16721_ (.A(net1266),
    .X(_10525_));
 sg13g2_nand2_1 _16722_ (.Y(_10526_),
    .A(net1180),
    .B(_10516_));
 sg13g2_o21ai_1 _16723_ (.B1(_10526_),
    .Y(_00196_),
    .A1(net399),
    .A2(_10524_));
 sg13g2_nand2_1 _16724_ (.Y(_10527_),
    .A(net772),
    .B(\mem.mem_internal.code_mem[109][3] ));
 sg13g2_buf_1 _16725_ (.A(net1265),
    .X(_10528_));
 sg13g2_nand2_1 _16726_ (.Y(_10529_),
    .A(net1179),
    .B(_10516_));
 sg13g2_o21ai_1 _16727_ (.B1(_10529_),
    .Y(_00197_),
    .A1(_10517_),
    .A2(_10527_));
 sg13g2_nand2_1 _16728_ (.Y(_10530_),
    .A(net772),
    .B(\mem.mem_internal.code_mem[109][4] ));
 sg13g2_buf_1 _16729_ (.A(net1264),
    .X(_10531_));
 sg13g2_nand2_1 _16730_ (.Y(_10532_),
    .A(net1178),
    .B(_10516_));
 sg13g2_o21ai_1 _16731_ (.B1(_10532_),
    .Y(_00198_),
    .A1(net399),
    .A2(_10530_));
 sg13g2_nand2_1 _16732_ (.Y(_10533_),
    .A(net772),
    .B(\mem.mem_internal.code_mem[109][5] ));
 sg13g2_buf_1 _16733_ (.A(net1263),
    .X(_10534_));
 sg13g2_nand2_1 _16734_ (.Y(_10535_),
    .A(net1177),
    .B(_10516_));
 sg13g2_o21ai_1 _16735_ (.B1(_10535_),
    .Y(_00199_),
    .A1(net399),
    .A2(_10533_));
 sg13g2_nand2_1 _16736_ (.Y(_10536_),
    .A(net772),
    .B(\mem.mem_internal.code_mem[109][6] ));
 sg13g2_buf_1 _16737_ (.A(net1262),
    .X(_10537_));
 sg13g2_nand2_1 _16738_ (.Y(_10538_),
    .A(net1176),
    .B(_10516_));
 sg13g2_o21ai_1 _16739_ (.B1(_10538_),
    .Y(_00200_),
    .A1(net399),
    .A2(_10536_));
 sg13g2_nand2_1 _16740_ (.Y(_10539_),
    .A(net772),
    .B(\mem.mem_internal.code_mem[109][7] ));
 sg13g2_buf_1 _16741_ (.A(net1261),
    .X(_10540_));
 sg13g2_nand2_1 _16742_ (.Y(_10541_),
    .A(net1175),
    .B(_10516_));
 sg13g2_o21ai_1 _16743_ (.B1(_10541_),
    .Y(_00201_),
    .A1(net399),
    .A2(_10539_));
 sg13g2_nand2_1 _16744_ (.Y(_10542_),
    .A(net850),
    .B(\mem.mem_internal.code_mem[10][0] ));
 sg13g2_nor2_1 _16745_ (.A(net470),
    .B(net550),
    .Y(_10543_));
 sg13g2_buf_2 _16746_ (.A(_10543_),
    .X(_10544_));
 sg13g2_buf_1 _16747_ (.A(_10544_),
    .X(_10545_));
 sg13g2_nand2_1 _16748_ (.Y(_10546_),
    .A(net1182),
    .B(net283));
 sg13g2_o21ai_1 _16749_ (.B1(_10546_),
    .Y(_00202_),
    .A1(_10542_),
    .A2(net283));
 sg13g2_nand2_1 _16750_ (.Y(_10547_),
    .A(net772),
    .B(\mem.mem_internal.code_mem[10][1] ));
 sg13g2_nand2_1 _16751_ (.Y(_10548_),
    .A(net1181),
    .B(net283));
 sg13g2_o21ai_1 _16752_ (.B1(_10548_),
    .Y(_00203_),
    .A1(net283),
    .A2(_10547_));
 sg13g2_nand2_1 _16753_ (.Y(_10549_),
    .A(net772),
    .B(\mem.mem_internal.code_mem[10][2] ));
 sg13g2_nand2_1 _16754_ (.Y(_10550_),
    .A(net1180),
    .B(_10544_));
 sg13g2_o21ai_1 _16755_ (.B1(_10550_),
    .Y(_00204_),
    .A1(net283),
    .A2(_10549_));
 sg13g2_nand2_1 _16756_ (.Y(_10551_),
    .A(_10523_),
    .B(\mem.mem_internal.code_mem[10][3] ));
 sg13g2_nand2_1 _16757_ (.Y(_10552_),
    .A(net1179),
    .B(_10544_));
 sg13g2_o21ai_1 _16758_ (.B1(_10552_),
    .Y(_00205_),
    .A1(net283),
    .A2(_10551_));
 sg13g2_nand2_1 _16759_ (.Y(_10553_),
    .A(_10523_),
    .B(\mem.mem_internal.code_mem[10][4] ));
 sg13g2_nand2_1 _16760_ (.Y(_10554_),
    .A(net1178),
    .B(_10544_));
 sg13g2_o21ai_1 _16761_ (.B1(_10554_),
    .Y(_00206_),
    .A1(net283),
    .A2(_10553_));
 sg13g2_buf_1 _16762_ (.A(_10416_),
    .X(_10555_));
 sg13g2_nand2_1 _16763_ (.Y(_10556_),
    .A(_10555_),
    .B(\mem.mem_internal.code_mem[10][5] ));
 sg13g2_nand2_1 _16764_ (.Y(_10557_),
    .A(net1177),
    .B(_10544_));
 sg13g2_o21ai_1 _16765_ (.B1(_10557_),
    .Y(_00207_),
    .A1(net283),
    .A2(_10556_));
 sg13g2_nand2_1 _16766_ (.Y(_10558_),
    .A(_10555_),
    .B(\mem.mem_internal.code_mem[10][6] ));
 sg13g2_nand2_1 _16767_ (.Y(_10559_),
    .A(net1176),
    .B(_10544_));
 sg13g2_o21ai_1 _16768_ (.B1(_10559_),
    .Y(_00208_),
    .A1(_10545_),
    .A2(_10558_));
 sg13g2_nand2_1 _16769_ (.Y(_10560_),
    .A(net771),
    .B(\mem.mem_internal.code_mem[10][7] ));
 sg13g2_nand2_1 _16770_ (.Y(_10561_),
    .A(net1175),
    .B(_10544_));
 sg13g2_o21ai_1 _16771_ (.B1(_10561_),
    .Y(_00209_),
    .A1(_10545_),
    .A2(_10560_));
 sg13g2_nand2_1 _16772_ (.Y(_10562_),
    .A(net850),
    .B(\mem.mem_internal.code_mem[110][0] ));
 sg13g2_nand3_1 _16773_ (.B(_10112_),
    .C(_10347_),
    .A(_10107_),
    .Y(_10563_));
 sg13g2_buf_2 _16774_ (.A(_10563_),
    .X(_10564_));
 sg13g2_buf_1 _16775_ (.A(_10564_),
    .X(_10565_));
 sg13g2_nor2_1 _16776_ (.A(_10300_),
    .B(net547),
    .Y(_10566_));
 sg13g2_buf_2 _16777_ (.A(_10566_),
    .X(_10567_));
 sg13g2_buf_1 _16778_ (.A(_10567_),
    .X(_10568_));
 sg13g2_nand2_1 _16779_ (.Y(_10569_),
    .A(net1182),
    .B(net398));
 sg13g2_o21ai_1 _16780_ (.B1(_10569_),
    .Y(_00210_),
    .A1(_10562_),
    .A2(net398));
 sg13g2_nand2_1 _16781_ (.Y(_10570_),
    .A(net771),
    .B(\mem.mem_internal.code_mem[110][1] ));
 sg13g2_nand2_1 _16782_ (.Y(_10571_),
    .A(net1181),
    .B(net398));
 sg13g2_o21ai_1 _16783_ (.B1(_10571_),
    .Y(_00211_),
    .A1(net398),
    .A2(_10570_));
 sg13g2_nand2_1 _16784_ (.Y(_10572_),
    .A(net771),
    .B(\mem.mem_internal.code_mem[110][2] ));
 sg13g2_nand2_1 _16785_ (.Y(_10573_),
    .A(net1180),
    .B(_10567_));
 sg13g2_o21ai_1 _16786_ (.B1(_10573_),
    .Y(_00212_),
    .A1(net398),
    .A2(_10572_));
 sg13g2_nand2_1 _16787_ (.Y(_10574_),
    .A(net771),
    .B(\mem.mem_internal.code_mem[110][3] ));
 sg13g2_nand2_1 _16788_ (.Y(_10575_),
    .A(net1179),
    .B(_10567_));
 sg13g2_o21ai_1 _16789_ (.B1(_10575_),
    .Y(_00213_),
    .A1(net398),
    .A2(_10574_));
 sg13g2_nand2_1 _16790_ (.Y(_10576_),
    .A(net771),
    .B(\mem.mem_internal.code_mem[110][4] ));
 sg13g2_nand2_1 _16791_ (.Y(_10577_),
    .A(net1178),
    .B(_10567_));
 sg13g2_o21ai_1 _16792_ (.B1(_10577_),
    .Y(_00214_),
    .A1(net398),
    .A2(_10576_));
 sg13g2_nand2_1 _16793_ (.Y(_10578_),
    .A(net771),
    .B(\mem.mem_internal.code_mem[110][5] ));
 sg13g2_nand2_1 _16794_ (.Y(_10579_),
    .A(net1177),
    .B(_10567_));
 sg13g2_o21ai_1 _16795_ (.B1(_10579_),
    .Y(_00215_),
    .A1(net398),
    .A2(_10578_));
 sg13g2_nand2_1 _16796_ (.Y(_10580_),
    .A(net771),
    .B(\mem.mem_internal.code_mem[110][6] ));
 sg13g2_nand2_1 _16797_ (.Y(_10581_),
    .A(net1176),
    .B(_10567_));
 sg13g2_o21ai_1 _16798_ (.B1(_10581_),
    .Y(_00216_),
    .A1(_10568_),
    .A2(_10580_));
 sg13g2_nand2_1 _16799_ (.Y(_10582_),
    .A(net771),
    .B(\mem.mem_internal.code_mem[110][7] ));
 sg13g2_nand2_1 _16800_ (.Y(_10583_),
    .A(net1175),
    .B(_10567_));
 sg13g2_o21ai_1 _16801_ (.B1(_10583_),
    .Y(_00217_),
    .A1(_10568_),
    .A2(_10582_));
 sg13g2_nand2_1 _16802_ (.Y(_10584_),
    .A(net850),
    .B(\mem.mem_internal.code_mem[111][0] ));
 sg13g2_nand4_1 _16803_ (.B(net1271),
    .C(net1295),
    .A(net1293),
    .Y(_10585_),
    .D(net1294));
 sg13g2_buf_2 _16804_ (.A(_10585_),
    .X(_10586_));
 sg13g2_buf_1 _16805_ (.A(_10586_),
    .X(_10587_));
 sg13g2_nor2_1 _16806_ (.A(_10300_),
    .B(net770),
    .Y(_10588_));
 sg13g2_buf_2 _16807_ (.A(_10588_),
    .X(_10589_));
 sg13g2_buf_1 _16808_ (.A(_10589_),
    .X(_10590_));
 sg13g2_nand2_1 _16809_ (.Y(_10591_),
    .A(net1182),
    .B(net397));
 sg13g2_o21ai_1 _16810_ (.B1(_10591_),
    .Y(_00218_),
    .A1(_10584_),
    .A2(net397));
 sg13g2_buf_1 _16811_ (.A(_10416_),
    .X(_10592_));
 sg13g2_nand2_1 _16812_ (.Y(_10593_),
    .A(net769),
    .B(\mem.mem_internal.code_mem[111][1] ));
 sg13g2_nand2_1 _16813_ (.Y(_10594_),
    .A(net1181),
    .B(net397));
 sg13g2_o21ai_1 _16814_ (.B1(_10594_),
    .Y(_00219_),
    .A1(net397),
    .A2(_10593_));
 sg13g2_nand2_1 _16815_ (.Y(_10595_),
    .A(net769),
    .B(\mem.mem_internal.code_mem[111][2] ));
 sg13g2_nand2_1 _16816_ (.Y(_10596_),
    .A(net1180),
    .B(_10589_));
 sg13g2_o21ai_1 _16817_ (.B1(_10596_),
    .Y(_00220_),
    .A1(net397),
    .A2(_10595_));
 sg13g2_nand2_1 _16818_ (.Y(_10597_),
    .A(net769),
    .B(\mem.mem_internal.code_mem[111][3] ));
 sg13g2_nand2_1 _16819_ (.Y(_10598_),
    .A(net1179),
    .B(_10589_));
 sg13g2_o21ai_1 _16820_ (.B1(_10598_),
    .Y(_00221_),
    .A1(net397),
    .A2(_10597_));
 sg13g2_nand2_1 _16821_ (.Y(_10599_),
    .A(net769),
    .B(\mem.mem_internal.code_mem[111][4] ));
 sg13g2_nand2_1 _16822_ (.Y(_10600_),
    .A(net1178),
    .B(_10589_));
 sg13g2_o21ai_1 _16823_ (.B1(_10600_),
    .Y(_00222_),
    .A1(net397),
    .A2(_10599_));
 sg13g2_nand2_1 _16824_ (.Y(_10601_),
    .A(net769),
    .B(\mem.mem_internal.code_mem[111][5] ));
 sg13g2_nand2_1 _16825_ (.Y(_10602_),
    .A(net1177),
    .B(_10589_));
 sg13g2_o21ai_1 _16826_ (.B1(_10602_),
    .Y(_00223_),
    .A1(_10590_),
    .A2(_10601_));
 sg13g2_nand2_1 _16827_ (.Y(_10603_),
    .A(net769),
    .B(\mem.mem_internal.code_mem[111][6] ));
 sg13g2_nand2_1 _16828_ (.Y(_10604_),
    .A(net1176),
    .B(_10589_));
 sg13g2_o21ai_1 _16829_ (.B1(_10604_),
    .Y(_00224_),
    .A1(_10590_),
    .A2(_10603_));
 sg13g2_nand2_1 _16830_ (.Y(_10605_),
    .A(net769),
    .B(\mem.mem_internal.code_mem[111][7] ));
 sg13g2_nand2_1 _16831_ (.Y(_10606_),
    .A(net1175),
    .B(_10589_));
 sg13g2_o21ai_1 _16832_ (.B1(_10606_),
    .Y(_00225_),
    .A1(net397),
    .A2(_10605_));
 sg13g2_nor3_1 _16833_ (.A(_10114_),
    .B(_10123_),
    .C(_10243_),
    .Y(_10607_));
 sg13g2_nand2_1 _16834_ (.Y(_10608_),
    .A(_10297_),
    .B(_10607_));
 sg13g2_buf_2 _16835_ (.A(_10608_),
    .X(_10609_));
 sg13g2_buf_1 _16836_ (.A(_10609_),
    .X(_10610_));
 sg13g2_nor2_1 _16837_ (.A(net529),
    .B(_10610_),
    .Y(_10611_));
 sg13g2_buf_2 _16838_ (.A(_10611_),
    .X(_10612_));
 sg13g2_buf_1 _16839_ (.A(_10612_),
    .X(_10613_));
 sg13g2_nand2_1 _16840_ (.Y(_10614_),
    .A(net769),
    .B(\mem.mem_internal.code_mem[112][0] ));
 sg13g2_nand2_1 _16841_ (.Y(_10615_),
    .A(net1182),
    .B(net282));
 sg13g2_o21ai_1 _16842_ (.B1(_10615_),
    .Y(_00226_),
    .A1(net282),
    .A2(_10614_));
 sg13g2_nand2_1 _16843_ (.Y(_10616_),
    .A(_10592_),
    .B(\mem.mem_internal.code_mem[112][1] ));
 sg13g2_nand2_1 _16844_ (.Y(_10617_),
    .A(net1181),
    .B(net282));
 sg13g2_o21ai_1 _16845_ (.B1(_10617_),
    .Y(_00227_),
    .A1(net282),
    .A2(_10616_));
 sg13g2_nand2_1 _16846_ (.Y(_10618_),
    .A(_10592_),
    .B(\mem.mem_internal.code_mem[112][2] ));
 sg13g2_nand2_1 _16847_ (.Y(_10619_),
    .A(net1180),
    .B(_10612_));
 sg13g2_o21ai_1 _16848_ (.B1(_10619_),
    .Y(_00228_),
    .A1(net282),
    .A2(_10618_));
 sg13g2_buf_1 _16849_ (.A(_10416_),
    .X(_10620_));
 sg13g2_nand2_1 _16850_ (.Y(_10621_),
    .A(net768),
    .B(\mem.mem_internal.code_mem[112][3] ));
 sg13g2_nand2_1 _16851_ (.Y(_10622_),
    .A(net1179),
    .B(_10612_));
 sg13g2_o21ai_1 _16852_ (.B1(_10622_),
    .Y(_00229_),
    .A1(_10613_),
    .A2(_10621_));
 sg13g2_nand2_1 _16853_ (.Y(_10623_),
    .A(net768),
    .B(\mem.mem_internal.code_mem[112][4] ));
 sg13g2_nand2_1 _16854_ (.Y(_10624_),
    .A(net1178),
    .B(_10612_));
 sg13g2_o21ai_1 _16855_ (.B1(_10624_),
    .Y(_00230_),
    .A1(net282),
    .A2(_10623_));
 sg13g2_nand2_1 _16856_ (.Y(_10625_),
    .A(net768),
    .B(\mem.mem_internal.code_mem[112][5] ));
 sg13g2_nand2_1 _16857_ (.Y(_10626_),
    .A(net1177),
    .B(_10612_));
 sg13g2_o21ai_1 _16858_ (.B1(_10626_),
    .Y(_00231_),
    .A1(net282),
    .A2(_10625_));
 sg13g2_nand2_1 _16859_ (.Y(_10627_),
    .A(_10620_),
    .B(\mem.mem_internal.code_mem[112][6] ));
 sg13g2_nand2_1 _16860_ (.Y(_10628_),
    .A(net1176),
    .B(_10612_));
 sg13g2_o21ai_1 _16861_ (.B1(_10628_),
    .Y(_00232_),
    .A1(net282),
    .A2(_10627_));
 sg13g2_nand2_1 _16862_ (.Y(_10629_),
    .A(net768),
    .B(\mem.mem_internal.code_mem[112][7] ));
 sg13g2_nand2_1 _16863_ (.Y(_10630_),
    .A(net1175),
    .B(_10612_));
 sg13g2_o21ai_1 _16864_ (.B1(_10630_),
    .Y(_00233_),
    .A1(_10613_),
    .A2(_10629_));
 sg13g2_nand2_1 _16865_ (.Y(_10631_),
    .A(_10229_),
    .B(_10323_));
 sg13g2_buf_2 _16866_ (.A(_10631_),
    .X(_10632_));
 sg13g2_buf_1 _16867_ (.A(_10632_),
    .X(_10633_));
 sg13g2_nor2_1 _16868_ (.A(_10609_),
    .B(net528),
    .Y(_10634_));
 sg13g2_buf_2 _16869_ (.A(_10634_),
    .X(_10635_));
 sg13g2_buf_1 _16870_ (.A(_10635_),
    .X(_10636_));
 sg13g2_nand2_1 _16871_ (.Y(_10637_),
    .A(net768),
    .B(\mem.mem_internal.code_mem[113][0] ));
 sg13g2_nand2_1 _16872_ (.Y(_10638_),
    .A(net1182),
    .B(net396));
 sg13g2_o21ai_1 _16873_ (.B1(_10638_),
    .Y(_00234_),
    .A1(net396),
    .A2(_10637_));
 sg13g2_nand2_1 _16874_ (.Y(_10639_),
    .A(net768),
    .B(\mem.mem_internal.code_mem[113][1] ));
 sg13g2_nand2_1 _16875_ (.Y(_10640_),
    .A(net1181),
    .B(net396));
 sg13g2_o21ai_1 _16876_ (.B1(_10640_),
    .Y(_00235_),
    .A1(net396),
    .A2(_10639_));
 sg13g2_nand2_1 _16877_ (.Y(_10641_),
    .A(net768),
    .B(\mem.mem_internal.code_mem[113][2] ));
 sg13g2_nand2_1 _16878_ (.Y(_10642_),
    .A(net1180),
    .B(_10635_));
 sg13g2_o21ai_1 _16879_ (.B1(_10642_),
    .Y(_00236_),
    .A1(net396),
    .A2(_10641_));
 sg13g2_nand2_1 _16880_ (.Y(_10643_),
    .A(_10620_),
    .B(\mem.mem_internal.code_mem[113][3] ));
 sg13g2_nand2_1 _16881_ (.Y(_10644_),
    .A(net1179),
    .B(_10635_));
 sg13g2_o21ai_1 _16882_ (.B1(_10644_),
    .Y(_00237_),
    .A1(_10636_),
    .A2(_10643_));
 sg13g2_nand2_1 _16883_ (.Y(_10645_),
    .A(net768),
    .B(\mem.mem_internal.code_mem[113][4] ));
 sg13g2_nand2_1 _16884_ (.Y(_10646_),
    .A(net1178),
    .B(_10635_));
 sg13g2_o21ai_1 _16885_ (.B1(_10646_),
    .Y(_00238_),
    .A1(net396),
    .A2(_10645_));
 sg13g2_buf_1 _16886_ (.A(_10415_),
    .X(_10647_));
 sg13g2_buf_1 _16887_ (.A(_10647_),
    .X(_10648_));
 sg13g2_nand2_1 _16888_ (.Y(_10649_),
    .A(net767),
    .B(\mem.mem_internal.code_mem[113][5] ));
 sg13g2_nand2_1 _16889_ (.Y(_10650_),
    .A(net1177),
    .B(_10635_));
 sg13g2_o21ai_1 _16890_ (.B1(_10650_),
    .Y(_00239_),
    .A1(net396),
    .A2(_10649_));
 sg13g2_nand2_1 _16891_ (.Y(_10651_),
    .A(net767),
    .B(\mem.mem_internal.code_mem[113][6] ));
 sg13g2_nand2_1 _16892_ (.Y(_10652_),
    .A(net1176),
    .B(_10635_));
 sg13g2_o21ai_1 _16893_ (.B1(_10652_),
    .Y(_00240_),
    .A1(net396),
    .A2(_10651_));
 sg13g2_nand2_1 _16894_ (.Y(_10653_),
    .A(_10648_),
    .B(\mem.mem_internal.code_mem[113][7] ));
 sg13g2_nand2_1 _16895_ (.Y(_10654_),
    .A(net1175),
    .B(_10635_));
 sg13g2_o21ai_1 _16896_ (.B1(_10654_),
    .Y(_00241_),
    .A1(_10636_),
    .A2(_10653_));
 sg13g2_nand2_1 _16897_ (.Y(_10655_),
    .A(_10229_),
    .B(_10347_));
 sg13g2_buf_2 _16898_ (.A(_10655_),
    .X(_10656_));
 sg13g2_buf_1 _16899_ (.A(_10656_),
    .X(_10657_));
 sg13g2_nor2_1 _16900_ (.A(_10609_),
    .B(net527),
    .Y(_10658_));
 sg13g2_buf_2 _16901_ (.A(_10658_),
    .X(_10659_));
 sg13g2_buf_1 _16902_ (.A(_10659_),
    .X(_10660_));
 sg13g2_nand2_1 _16903_ (.Y(_10661_),
    .A(net767),
    .B(\mem.mem_internal.code_mem[114][0] ));
 sg13g2_nand2_1 _16904_ (.Y(_10662_),
    .A(net1182),
    .B(net395));
 sg13g2_o21ai_1 _16905_ (.B1(_10662_),
    .Y(_00242_),
    .A1(net395),
    .A2(_10661_));
 sg13g2_nand2_1 _16906_ (.Y(_10663_),
    .A(net767),
    .B(\mem.mem_internal.code_mem[114][1] ));
 sg13g2_nand2_1 _16907_ (.Y(_10664_),
    .A(net1181),
    .B(net395));
 sg13g2_o21ai_1 _16908_ (.B1(_10664_),
    .Y(_00243_),
    .A1(net395),
    .A2(_10663_));
 sg13g2_nand2_1 _16909_ (.Y(_10665_),
    .A(net767),
    .B(\mem.mem_internal.code_mem[114][2] ));
 sg13g2_nand2_1 _16910_ (.Y(_10666_),
    .A(net1180),
    .B(_10659_));
 sg13g2_o21ai_1 _16911_ (.B1(_10666_),
    .Y(_00244_),
    .A1(net395),
    .A2(_10665_));
 sg13g2_nand2_1 _16912_ (.Y(_10667_),
    .A(_10648_),
    .B(\mem.mem_internal.code_mem[114][3] ));
 sg13g2_nand2_1 _16913_ (.Y(_10668_),
    .A(net1179),
    .B(_10659_));
 sg13g2_o21ai_1 _16914_ (.B1(_10668_),
    .Y(_00245_),
    .A1(_10660_),
    .A2(_10667_));
 sg13g2_nand2_1 _16915_ (.Y(_10669_),
    .A(net767),
    .B(\mem.mem_internal.code_mem[114][4] ));
 sg13g2_nand2_1 _16916_ (.Y(_10670_),
    .A(net1178),
    .B(_10659_));
 sg13g2_o21ai_1 _16917_ (.B1(_10670_),
    .Y(_00246_),
    .A1(net395),
    .A2(_10669_));
 sg13g2_nand2_1 _16918_ (.Y(_10671_),
    .A(net767),
    .B(\mem.mem_internal.code_mem[114][5] ));
 sg13g2_nand2_1 _16919_ (.Y(_10672_),
    .A(net1177),
    .B(_10659_));
 sg13g2_o21ai_1 _16920_ (.B1(_10672_),
    .Y(_00247_),
    .A1(net395),
    .A2(_10671_));
 sg13g2_nand2_1 _16921_ (.Y(_10673_),
    .A(net767),
    .B(\mem.mem_internal.code_mem[114][6] ));
 sg13g2_nand2_1 _16922_ (.Y(_10674_),
    .A(net1176),
    .B(_10659_));
 sg13g2_o21ai_1 _16923_ (.B1(_10674_),
    .Y(_00248_),
    .A1(net395),
    .A2(_10673_));
 sg13g2_buf_1 _16924_ (.A(_10647_),
    .X(_10675_));
 sg13g2_nand2_1 _16925_ (.Y(_10676_),
    .A(net766),
    .B(\mem.mem_internal.code_mem[114][7] ));
 sg13g2_nand2_1 _16926_ (.Y(_10677_),
    .A(net1175),
    .B(_10659_));
 sg13g2_o21ai_1 _16927_ (.B1(_10677_),
    .Y(_00249_),
    .A1(_10660_),
    .A2(_10676_));
 sg13g2_nand3_1 _16928_ (.B(net1294),
    .C(_10229_),
    .A(net1295),
    .Y(_10678_));
 sg13g2_buf_2 _16929_ (.A(_10678_),
    .X(_10679_));
 sg13g2_buf_1 _16930_ (.A(_10679_),
    .X(_10680_));
 sg13g2_nor2_1 _16931_ (.A(_10609_),
    .B(net526),
    .Y(_10681_));
 sg13g2_buf_2 _16932_ (.A(_10681_),
    .X(_10682_));
 sg13g2_buf_1 _16933_ (.A(_10682_),
    .X(_10683_));
 sg13g2_nand2_1 _16934_ (.Y(_10684_),
    .A(net766),
    .B(\mem.mem_internal.code_mem[115][0] ));
 sg13g2_nand2_1 _16935_ (.Y(_10685_),
    .A(net1182),
    .B(net394));
 sg13g2_o21ai_1 _16936_ (.B1(_10685_),
    .Y(_00250_),
    .A1(net394),
    .A2(_10684_));
 sg13g2_nand2_1 _16937_ (.Y(_10686_),
    .A(net766),
    .B(\mem.mem_internal.code_mem[115][1] ));
 sg13g2_nand2_1 _16938_ (.Y(_10687_),
    .A(net1181),
    .B(net394));
 sg13g2_o21ai_1 _16939_ (.B1(_10687_),
    .Y(_00251_),
    .A1(net394),
    .A2(_10686_));
 sg13g2_nand2_1 _16940_ (.Y(_10688_),
    .A(net766),
    .B(\mem.mem_internal.code_mem[115][2] ));
 sg13g2_nand2_1 _16941_ (.Y(_10689_),
    .A(net1180),
    .B(_10682_));
 sg13g2_o21ai_1 _16942_ (.B1(_10689_),
    .Y(_00252_),
    .A1(net394),
    .A2(_10688_));
 sg13g2_nand2_1 _16943_ (.Y(_10690_),
    .A(net766),
    .B(\mem.mem_internal.code_mem[115][3] ));
 sg13g2_nand2_1 _16944_ (.Y(_10691_),
    .A(net1179),
    .B(_10682_));
 sg13g2_o21ai_1 _16945_ (.B1(_10691_),
    .Y(_00253_),
    .A1(_10683_),
    .A2(_10690_));
 sg13g2_nand2_1 _16946_ (.Y(_10692_),
    .A(net766),
    .B(\mem.mem_internal.code_mem[115][4] ));
 sg13g2_nand2_1 _16947_ (.Y(_10693_),
    .A(net1178),
    .B(_10682_));
 sg13g2_o21ai_1 _16948_ (.B1(_10693_),
    .Y(_00254_),
    .A1(net394),
    .A2(_10692_));
 sg13g2_nand2_1 _16949_ (.Y(_10694_),
    .A(net766),
    .B(\mem.mem_internal.code_mem[115][5] ));
 sg13g2_nand2_1 _16950_ (.Y(_10695_),
    .A(net1177),
    .B(_10682_));
 sg13g2_o21ai_1 _16951_ (.B1(_10695_),
    .Y(_00255_),
    .A1(net394),
    .A2(_10694_));
 sg13g2_nand2_1 _16952_ (.Y(_10696_),
    .A(_10675_),
    .B(\mem.mem_internal.code_mem[115][6] ));
 sg13g2_nand2_1 _16953_ (.Y(_10697_),
    .A(net1176),
    .B(_10682_));
 sg13g2_o21ai_1 _16954_ (.B1(_10697_),
    .Y(_00256_),
    .A1(net394),
    .A2(_10696_));
 sg13g2_nand2_1 _16955_ (.Y(_10698_),
    .A(_10675_),
    .B(\mem.mem_internal.code_mem[115][7] ));
 sg13g2_nand2_1 _16956_ (.Y(_10699_),
    .A(net1175),
    .B(_10682_));
 sg13g2_o21ai_1 _16957_ (.B1(_10699_),
    .Y(_00257_),
    .A1(_10683_),
    .A2(_10698_));
 sg13g2_nor2_1 _16958_ (.A(net556),
    .B(net468),
    .Y(_10700_));
 sg13g2_buf_2 _16959_ (.A(_10700_),
    .X(_10701_));
 sg13g2_buf_1 _16960_ (.A(_10701_),
    .X(_10702_));
 sg13g2_nand2_1 _16961_ (.Y(_10703_),
    .A(net766),
    .B(\mem.mem_internal.code_mem[116][0] ));
 sg13g2_nand2_1 _16962_ (.Y(_10704_),
    .A(_10518_),
    .B(net281));
 sg13g2_o21ai_1 _16963_ (.B1(_10704_),
    .Y(_00258_),
    .A1(net281),
    .A2(_10703_));
 sg13g2_buf_1 _16964_ (.A(_10647_),
    .X(_10705_));
 sg13g2_nand2_1 _16965_ (.Y(_10706_),
    .A(net765),
    .B(\mem.mem_internal.code_mem[116][1] ));
 sg13g2_nand2_1 _16966_ (.Y(_10707_),
    .A(_10521_),
    .B(net281));
 sg13g2_o21ai_1 _16967_ (.B1(_10707_),
    .Y(_00259_),
    .A1(net281),
    .A2(_10706_));
 sg13g2_nand2_1 _16968_ (.Y(_10708_),
    .A(net765),
    .B(\mem.mem_internal.code_mem[116][2] ));
 sg13g2_nand2_1 _16969_ (.Y(_10709_),
    .A(_10525_),
    .B(_10701_));
 sg13g2_o21ai_1 _16970_ (.B1(_10709_),
    .Y(_00260_),
    .A1(net281),
    .A2(_10708_));
 sg13g2_nand2_1 _16971_ (.Y(_10710_),
    .A(net765),
    .B(\mem.mem_internal.code_mem[116][3] ));
 sg13g2_nand2_1 _16972_ (.Y(_10711_),
    .A(_10528_),
    .B(_10701_));
 sg13g2_o21ai_1 _16973_ (.B1(_10711_),
    .Y(_00261_),
    .A1(net281),
    .A2(_10710_));
 sg13g2_nand2_1 _16974_ (.Y(_10712_),
    .A(net765),
    .B(\mem.mem_internal.code_mem[116][4] ));
 sg13g2_nand2_1 _16975_ (.Y(_10713_),
    .A(_10531_),
    .B(_10701_));
 sg13g2_o21ai_1 _16976_ (.B1(_10713_),
    .Y(_00262_),
    .A1(net281),
    .A2(_10712_));
 sg13g2_nand2_1 _16977_ (.Y(_10714_),
    .A(_10705_),
    .B(\mem.mem_internal.code_mem[116][5] ));
 sg13g2_nand2_1 _16978_ (.Y(_10715_),
    .A(_10534_),
    .B(_10701_));
 sg13g2_o21ai_1 _16979_ (.B1(_10715_),
    .Y(_00263_),
    .A1(_10702_),
    .A2(_10714_));
 sg13g2_nand2_1 _16980_ (.Y(_10716_),
    .A(_10705_),
    .B(\mem.mem_internal.code_mem[116][6] ));
 sg13g2_nand2_1 _16981_ (.Y(_10717_),
    .A(_10537_),
    .B(_10701_));
 sg13g2_o21ai_1 _16982_ (.B1(_10717_),
    .Y(_00264_),
    .A1(_10702_),
    .A2(_10716_));
 sg13g2_nand2_1 _16983_ (.Y(_10718_),
    .A(net765),
    .B(\mem.mem_internal.code_mem[116][7] ));
 sg13g2_nand2_1 _16984_ (.Y(_10719_),
    .A(_10540_),
    .B(_10701_));
 sg13g2_o21ai_1 _16985_ (.B1(_10719_),
    .Y(_00265_),
    .A1(net281),
    .A2(_10718_));
 sg13g2_nor2_1 _16986_ (.A(net555),
    .B(_10610_),
    .Y(_10720_));
 sg13g2_buf_2 _16987_ (.A(_10720_),
    .X(_10721_));
 sg13g2_buf_1 _16988_ (.A(_10721_),
    .X(_10722_));
 sg13g2_nand2_1 _16989_ (.Y(_10723_),
    .A(net765),
    .B(\mem.mem_internal.code_mem[117][0] ));
 sg13g2_nand2_1 _16990_ (.Y(_10724_),
    .A(_10518_),
    .B(net280));
 sg13g2_o21ai_1 _16991_ (.B1(_10724_),
    .Y(_00266_),
    .A1(net280),
    .A2(_10723_));
 sg13g2_nand2_1 _16992_ (.Y(_10725_),
    .A(net765),
    .B(\mem.mem_internal.code_mem[117][1] ));
 sg13g2_nand2_1 _16993_ (.Y(_10726_),
    .A(_10521_),
    .B(net280));
 sg13g2_o21ai_1 _16994_ (.B1(_10726_),
    .Y(_00267_),
    .A1(net280),
    .A2(_10725_));
 sg13g2_nand2_1 _16995_ (.Y(_10727_),
    .A(net765),
    .B(\mem.mem_internal.code_mem[117][2] ));
 sg13g2_nand2_1 _16996_ (.Y(_10728_),
    .A(_10525_),
    .B(_10721_));
 sg13g2_o21ai_1 _16997_ (.B1(_10728_),
    .Y(_00268_),
    .A1(net280),
    .A2(_10727_));
 sg13g2_buf_1 _16998_ (.A(_10647_),
    .X(_10729_));
 sg13g2_nand2_1 _16999_ (.Y(_10730_),
    .A(net764),
    .B(\mem.mem_internal.code_mem[117][3] ));
 sg13g2_nand2_1 _17000_ (.Y(_10731_),
    .A(_10528_),
    .B(_10721_));
 sg13g2_o21ai_1 _17001_ (.B1(_10731_),
    .Y(_00269_),
    .A1(net280),
    .A2(_10730_));
 sg13g2_nand2_1 _17002_ (.Y(_10732_),
    .A(net764),
    .B(\mem.mem_internal.code_mem[117][4] ));
 sg13g2_nand2_1 _17003_ (.Y(_10733_),
    .A(_10531_),
    .B(_10721_));
 sg13g2_o21ai_1 _17004_ (.B1(_10733_),
    .Y(_00270_),
    .A1(net280),
    .A2(_10732_));
 sg13g2_nand2_1 _17005_ (.Y(_10734_),
    .A(net764),
    .B(\mem.mem_internal.code_mem[117][5] ));
 sg13g2_nand2_1 _17006_ (.Y(_10735_),
    .A(_10534_),
    .B(_10721_));
 sg13g2_o21ai_1 _17007_ (.B1(_10735_),
    .Y(_00271_),
    .A1(_10722_),
    .A2(_10734_));
 sg13g2_nand2_1 _17008_ (.Y(_10736_),
    .A(net764),
    .B(\mem.mem_internal.code_mem[117][6] ));
 sg13g2_nand2_1 _17009_ (.Y(_10737_),
    .A(_10537_),
    .B(_10721_));
 sg13g2_o21ai_1 _17010_ (.B1(_10737_),
    .Y(_00272_),
    .A1(_10722_),
    .A2(_10736_));
 sg13g2_nand2_1 _17011_ (.Y(_10738_),
    .A(net764),
    .B(\mem.mem_internal.code_mem[117][7] ));
 sg13g2_nand2_1 _17012_ (.Y(_10739_),
    .A(_10540_),
    .B(_10721_));
 sg13g2_o21ai_1 _17013_ (.B1(_10739_),
    .Y(_00273_),
    .A1(net280),
    .A2(_10738_));
 sg13g2_nor2_1 _17014_ (.A(net554),
    .B(net468),
    .Y(_10740_));
 sg13g2_buf_2 _17015_ (.A(_10740_),
    .X(_10741_));
 sg13g2_buf_1 _17016_ (.A(_10741_),
    .X(_10742_));
 sg13g2_nand2_1 _17017_ (.Y(_10743_),
    .A(net764),
    .B(\mem.mem_internal.code_mem[118][0] ));
 sg13g2_buf_1 _17018_ (.A(net1268),
    .X(_10744_));
 sg13g2_nand2_1 _17019_ (.Y(_10745_),
    .A(net1174),
    .B(net279));
 sg13g2_o21ai_1 _17020_ (.B1(_10745_),
    .Y(_00274_),
    .A1(net279),
    .A2(_10743_));
 sg13g2_nand2_1 _17021_ (.Y(_10746_),
    .A(net764),
    .B(\mem.mem_internal.code_mem[118][1] ));
 sg13g2_buf_1 _17022_ (.A(net1267),
    .X(_10747_));
 sg13g2_nand2_1 _17023_ (.Y(_10748_),
    .A(_10747_),
    .B(net279));
 sg13g2_o21ai_1 _17024_ (.B1(_10748_),
    .Y(_00275_),
    .A1(net279),
    .A2(_10746_));
 sg13g2_nand2_1 _17025_ (.Y(_10749_),
    .A(net764),
    .B(\mem.mem_internal.code_mem[118][2] ));
 sg13g2_buf_1 _17026_ (.A(net1266),
    .X(_10750_));
 sg13g2_nand2_1 _17027_ (.Y(_10751_),
    .A(_10750_),
    .B(_10741_));
 sg13g2_o21ai_1 _17028_ (.B1(_10751_),
    .Y(_00276_),
    .A1(net279),
    .A2(_10749_));
 sg13g2_nand2_1 _17029_ (.Y(_10752_),
    .A(_10729_),
    .B(\mem.mem_internal.code_mem[118][3] ));
 sg13g2_buf_1 _17030_ (.A(net1265),
    .X(_10753_));
 sg13g2_nand2_1 _17031_ (.Y(_10754_),
    .A(_10753_),
    .B(_10741_));
 sg13g2_o21ai_1 _17032_ (.B1(_10754_),
    .Y(_00277_),
    .A1(net279),
    .A2(_10752_));
 sg13g2_nand2_1 _17033_ (.Y(_10755_),
    .A(_10729_),
    .B(\mem.mem_internal.code_mem[118][4] ));
 sg13g2_buf_1 _17034_ (.A(net1264),
    .X(_10756_));
 sg13g2_nand2_1 _17035_ (.Y(_10757_),
    .A(_10756_),
    .B(_10741_));
 sg13g2_o21ai_1 _17036_ (.B1(_10757_),
    .Y(_00278_),
    .A1(net279),
    .A2(_10755_));
 sg13g2_buf_1 _17037_ (.A(_10647_),
    .X(_10758_));
 sg13g2_nand2_1 _17038_ (.Y(_10759_),
    .A(net763),
    .B(\mem.mem_internal.code_mem[118][5] ));
 sg13g2_buf_1 _17039_ (.A(net1263),
    .X(_10760_));
 sg13g2_nand2_1 _17040_ (.Y(_10761_),
    .A(_10760_),
    .B(_10741_));
 sg13g2_o21ai_1 _17041_ (.B1(_10761_),
    .Y(_00279_),
    .A1(_10742_),
    .A2(_10759_));
 sg13g2_nand2_1 _17042_ (.Y(_10762_),
    .A(net763),
    .B(\mem.mem_internal.code_mem[118][6] ));
 sg13g2_buf_1 _17043_ (.A(net1262),
    .X(_10763_));
 sg13g2_nand2_1 _17044_ (.Y(_10764_),
    .A(_10763_),
    .B(_10741_));
 sg13g2_o21ai_1 _17045_ (.B1(_10764_),
    .Y(_00280_),
    .A1(_10742_),
    .A2(_10762_));
 sg13g2_nand2_1 _17046_ (.Y(_10765_),
    .A(net763),
    .B(\mem.mem_internal.code_mem[118][7] ));
 sg13g2_buf_1 _17047_ (.A(net1261),
    .X(_10766_));
 sg13g2_nand2_1 _17048_ (.Y(_10767_),
    .A(net1167),
    .B(_10741_));
 sg13g2_o21ai_1 _17049_ (.B1(_10767_),
    .Y(_00281_),
    .A1(net279),
    .A2(_10765_));
 sg13g2_nor2_1 _17050_ (.A(net553),
    .B(net468),
    .Y(_10768_));
 sg13g2_buf_2 _17051_ (.A(_10768_),
    .X(_10769_));
 sg13g2_buf_1 _17052_ (.A(_10769_),
    .X(_10770_));
 sg13g2_nand2_1 _17053_ (.Y(_10771_),
    .A(_10758_),
    .B(\mem.mem_internal.code_mem[119][0] ));
 sg13g2_nand2_1 _17054_ (.Y(_10772_),
    .A(_10744_),
    .B(net278));
 sg13g2_o21ai_1 _17055_ (.B1(_10772_),
    .Y(_00282_),
    .A1(net278),
    .A2(_10771_));
 sg13g2_nand2_1 _17056_ (.Y(_10773_),
    .A(net763),
    .B(\mem.mem_internal.code_mem[119][1] ));
 sg13g2_nand2_1 _17057_ (.Y(_10774_),
    .A(_10747_),
    .B(net278));
 sg13g2_o21ai_1 _17058_ (.B1(_10774_),
    .Y(_00283_),
    .A1(net278),
    .A2(_10773_));
 sg13g2_nand2_1 _17059_ (.Y(_10775_),
    .A(net763),
    .B(\mem.mem_internal.code_mem[119][2] ));
 sg13g2_nand2_1 _17060_ (.Y(_10776_),
    .A(_10750_),
    .B(_10769_));
 sg13g2_o21ai_1 _17061_ (.B1(_10776_),
    .Y(_00284_),
    .A1(net278),
    .A2(_10775_));
 sg13g2_nand2_1 _17062_ (.Y(_10777_),
    .A(net763),
    .B(\mem.mem_internal.code_mem[119][3] ));
 sg13g2_nand2_1 _17063_ (.Y(_10778_),
    .A(net1171),
    .B(_10769_));
 sg13g2_o21ai_1 _17064_ (.B1(_10778_),
    .Y(_00285_),
    .A1(net278),
    .A2(_10777_));
 sg13g2_nand2_1 _17065_ (.Y(_10779_),
    .A(net763),
    .B(\mem.mem_internal.code_mem[119][4] ));
 sg13g2_nand2_1 _17066_ (.Y(_10780_),
    .A(net1170),
    .B(_10769_));
 sg13g2_o21ai_1 _17067_ (.B1(_10780_),
    .Y(_00286_),
    .A1(net278),
    .A2(_10779_));
 sg13g2_nand2_1 _17068_ (.Y(_10781_),
    .A(net763),
    .B(\mem.mem_internal.code_mem[119][5] ));
 sg13g2_nand2_1 _17069_ (.Y(_10782_),
    .A(net1169),
    .B(_10769_));
 sg13g2_o21ai_1 _17070_ (.B1(_10782_),
    .Y(_00287_),
    .A1(_10770_),
    .A2(_10781_));
 sg13g2_nand2_1 _17071_ (.Y(_10783_),
    .A(_10758_),
    .B(\mem.mem_internal.code_mem[119][6] ));
 sg13g2_nand2_1 _17072_ (.Y(_10784_),
    .A(net1168),
    .B(_10769_));
 sg13g2_o21ai_1 _17073_ (.B1(_10784_),
    .Y(_00288_),
    .A1(_10770_),
    .A2(_10783_));
 sg13g2_buf_1 _17074_ (.A(_10647_),
    .X(_10785_));
 sg13g2_nand2_1 _17075_ (.Y(_10786_),
    .A(net762),
    .B(\mem.mem_internal.code_mem[119][7] ));
 sg13g2_nand2_1 _17076_ (.Y(_10787_),
    .A(net1167),
    .B(_10769_));
 sg13g2_o21ai_1 _17077_ (.B1(_10787_),
    .Y(_00289_),
    .A1(net278),
    .A2(_10786_));
 sg13g2_nand2_1 _17078_ (.Y(_10788_),
    .A(_10488_),
    .B(\mem.mem_internal.code_mem[11][0] ));
 sg13g2_nor2_1 _17079_ (.A(net470),
    .B(net549),
    .Y(_10789_));
 sg13g2_buf_2 _17080_ (.A(_10789_),
    .X(_10790_));
 sg13g2_buf_1 _17081_ (.A(_10790_),
    .X(_10791_));
 sg13g2_nand2_1 _17082_ (.Y(_10792_),
    .A(net1174),
    .B(_10791_));
 sg13g2_o21ai_1 _17083_ (.B1(_10792_),
    .Y(_00290_),
    .A1(_10788_),
    .A2(_10791_));
 sg13g2_nand2_1 _17084_ (.Y(_10793_),
    .A(net762),
    .B(\mem.mem_internal.code_mem[11][1] ));
 sg13g2_nand2_1 _17085_ (.Y(_10794_),
    .A(net1173),
    .B(net277));
 sg13g2_o21ai_1 _17086_ (.B1(_10794_),
    .Y(_00291_),
    .A1(net277),
    .A2(_10793_));
 sg13g2_nand2_1 _17087_ (.Y(_10795_),
    .A(net762),
    .B(\mem.mem_internal.code_mem[11][2] ));
 sg13g2_nand2_1 _17088_ (.Y(_10796_),
    .A(net1172),
    .B(_10790_));
 sg13g2_o21ai_1 _17089_ (.B1(_10796_),
    .Y(_00292_),
    .A1(net277),
    .A2(_10795_));
 sg13g2_nand2_1 _17090_ (.Y(_10797_),
    .A(net762),
    .B(\mem.mem_internal.code_mem[11][3] ));
 sg13g2_nand2_1 _17091_ (.Y(_10798_),
    .A(net1171),
    .B(_10790_));
 sg13g2_o21ai_1 _17092_ (.B1(_10798_),
    .Y(_00293_),
    .A1(net277),
    .A2(_10797_));
 sg13g2_nand2_1 _17093_ (.Y(_10799_),
    .A(net762),
    .B(\mem.mem_internal.code_mem[11][4] ));
 sg13g2_nand2_1 _17094_ (.Y(_10800_),
    .A(net1170),
    .B(_10790_));
 sg13g2_o21ai_1 _17095_ (.B1(_10800_),
    .Y(_00294_),
    .A1(net277),
    .A2(_10799_));
 sg13g2_nand2_1 _17096_ (.Y(_10801_),
    .A(net762),
    .B(\mem.mem_internal.code_mem[11][5] ));
 sg13g2_nand2_1 _17097_ (.Y(_10802_),
    .A(net1169),
    .B(_10790_));
 sg13g2_o21ai_1 _17098_ (.B1(_10802_),
    .Y(_00295_),
    .A1(net277),
    .A2(_10801_));
 sg13g2_nand2_1 _17099_ (.Y(_10803_),
    .A(net762),
    .B(\mem.mem_internal.code_mem[11][6] ));
 sg13g2_nand2_1 _17100_ (.Y(_10804_),
    .A(net1168),
    .B(_10790_));
 sg13g2_o21ai_1 _17101_ (.B1(_10804_),
    .Y(_00296_),
    .A1(net277),
    .A2(_10803_));
 sg13g2_nand2_1 _17102_ (.Y(_10805_),
    .A(net762),
    .B(\mem.mem_internal.code_mem[11][7] ));
 sg13g2_nand2_1 _17103_ (.Y(_10806_),
    .A(net1167),
    .B(_10790_));
 sg13g2_o21ai_1 _17104_ (.B1(_10806_),
    .Y(_00297_),
    .A1(net277),
    .A2(_10805_));
 sg13g2_nor2_1 _17105_ (.A(net552),
    .B(net468),
    .Y(_10807_));
 sg13g2_buf_2 _17106_ (.A(_10807_),
    .X(_10808_));
 sg13g2_buf_1 _17107_ (.A(_10808_),
    .X(_10809_));
 sg13g2_nand2_1 _17108_ (.Y(_10810_),
    .A(_10785_),
    .B(\mem.mem_internal.code_mem[120][0] ));
 sg13g2_nand2_1 _17109_ (.Y(_10811_),
    .A(net1174),
    .B(net276));
 sg13g2_o21ai_1 _17110_ (.B1(_10811_),
    .Y(_00298_),
    .A1(net276),
    .A2(_10810_));
 sg13g2_nand2_1 _17111_ (.Y(_10812_),
    .A(_10785_),
    .B(\mem.mem_internal.code_mem[120][1] ));
 sg13g2_nand2_1 _17112_ (.Y(_10813_),
    .A(net1173),
    .B(net276));
 sg13g2_o21ai_1 _17113_ (.B1(_10813_),
    .Y(_00299_),
    .A1(net276),
    .A2(_10812_));
 sg13g2_buf_1 _17114_ (.A(_10647_),
    .X(_10814_));
 sg13g2_nand2_1 _17115_ (.Y(_10815_),
    .A(net761),
    .B(\mem.mem_internal.code_mem[120][2] ));
 sg13g2_nand2_1 _17116_ (.Y(_10816_),
    .A(net1172),
    .B(_10808_));
 sg13g2_o21ai_1 _17117_ (.B1(_10816_),
    .Y(_00300_),
    .A1(net276),
    .A2(_10815_));
 sg13g2_nand2_1 _17118_ (.Y(_10817_),
    .A(net761),
    .B(\mem.mem_internal.code_mem[120][3] ));
 sg13g2_nand2_1 _17119_ (.Y(_10818_),
    .A(_10753_),
    .B(_10808_));
 sg13g2_o21ai_1 _17120_ (.B1(_10818_),
    .Y(_00301_),
    .A1(net276),
    .A2(_10817_));
 sg13g2_nand2_1 _17121_ (.Y(_10819_),
    .A(net761),
    .B(\mem.mem_internal.code_mem[120][4] ));
 sg13g2_nand2_1 _17122_ (.Y(_10820_),
    .A(_10756_),
    .B(_10808_));
 sg13g2_o21ai_1 _17123_ (.B1(_10820_),
    .Y(_00302_),
    .A1(net276),
    .A2(_10819_));
 sg13g2_nand2_1 _17124_ (.Y(_10821_),
    .A(net761),
    .B(\mem.mem_internal.code_mem[120][5] ));
 sg13g2_nand2_1 _17125_ (.Y(_10822_),
    .A(_10760_),
    .B(_10808_));
 sg13g2_o21ai_1 _17126_ (.B1(_10822_),
    .Y(_00303_),
    .A1(net276),
    .A2(_10821_));
 sg13g2_nand2_1 _17127_ (.Y(_10823_),
    .A(_10814_),
    .B(\mem.mem_internal.code_mem[120][6] ));
 sg13g2_nand2_1 _17128_ (.Y(_10824_),
    .A(_10763_),
    .B(_10808_));
 sg13g2_o21ai_1 _17129_ (.B1(_10824_),
    .Y(_00304_),
    .A1(_10809_),
    .A2(_10823_));
 sg13g2_nand2_1 _17130_ (.Y(_10825_),
    .A(_10814_),
    .B(\mem.mem_internal.code_mem[120][7] ));
 sg13g2_nand2_1 _17131_ (.Y(_10826_),
    .A(net1167),
    .B(_10808_));
 sg13g2_o21ai_1 _17132_ (.B1(_10826_),
    .Y(_00305_),
    .A1(_10809_),
    .A2(_10825_));
 sg13g2_nor2_1 _17133_ (.A(net551),
    .B(net468),
    .Y(_10827_));
 sg13g2_buf_2 _17134_ (.A(_10827_),
    .X(_10828_));
 sg13g2_buf_1 _17135_ (.A(_10828_),
    .X(_10829_));
 sg13g2_nand2_1 _17136_ (.Y(_10830_),
    .A(net761),
    .B(\mem.mem_internal.code_mem[121][0] ));
 sg13g2_nand2_1 _17137_ (.Y(_10831_),
    .A(net1174),
    .B(net275));
 sg13g2_o21ai_1 _17138_ (.B1(_10831_),
    .Y(_00306_),
    .A1(net275),
    .A2(_10830_));
 sg13g2_nand2_1 _17139_ (.Y(_10832_),
    .A(net761),
    .B(\mem.mem_internal.code_mem[121][1] ));
 sg13g2_nand2_1 _17140_ (.Y(_10833_),
    .A(net1173),
    .B(net275));
 sg13g2_o21ai_1 _17141_ (.B1(_10833_),
    .Y(_00307_),
    .A1(_10829_),
    .A2(_10832_));
 sg13g2_nand2_1 _17142_ (.Y(_10834_),
    .A(net761),
    .B(\mem.mem_internal.code_mem[121][2] ));
 sg13g2_nand2_1 _17143_ (.Y(_10835_),
    .A(net1172),
    .B(_10828_));
 sg13g2_o21ai_1 _17144_ (.B1(_10835_),
    .Y(_00308_),
    .A1(net275),
    .A2(_10834_));
 sg13g2_nand2_1 _17145_ (.Y(_10836_),
    .A(net761),
    .B(\mem.mem_internal.code_mem[121][3] ));
 sg13g2_nand2_1 _17146_ (.Y(_10837_),
    .A(net1171),
    .B(_10828_));
 sg13g2_o21ai_1 _17147_ (.B1(_10837_),
    .Y(_00309_),
    .A1(net275),
    .A2(_10836_));
 sg13g2_buf_1 _17148_ (.A(_10415_),
    .X(_10838_));
 sg13g2_buf_1 _17149_ (.A(_10838_),
    .X(_10839_));
 sg13g2_nand2_1 _17150_ (.Y(_10840_),
    .A(net760),
    .B(\mem.mem_internal.code_mem[121][4] ));
 sg13g2_nand2_1 _17151_ (.Y(_10841_),
    .A(net1170),
    .B(_10828_));
 sg13g2_o21ai_1 _17152_ (.B1(_10841_),
    .Y(_00310_),
    .A1(net275),
    .A2(_10840_));
 sg13g2_nand2_1 _17153_ (.Y(_10842_),
    .A(net760),
    .B(\mem.mem_internal.code_mem[121][5] ));
 sg13g2_nand2_1 _17154_ (.Y(_10843_),
    .A(net1169),
    .B(_10828_));
 sg13g2_o21ai_1 _17155_ (.B1(_10843_),
    .Y(_00311_),
    .A1(net275),
    .A2(_10842_));
 sg13g2_nand2_1 _17156_ (.Y(_10844_),
    .A(_10839_),
    .B(\mem.mem_internal.code_mem[121][6] ));
 sg13g2_nand2_1 _17157_ (.Y(_10845_),
    .A(net1168),
    .B(_10828_));
 sg13g2_o21ai_1 _17158_ (.B1(_10845_),
    .Y(_00312_),
    .A1(_10829_),
    .A2(_10844_));
 sg13g2_nand2_1 _17159_ (.Y(_10846_),
    .A(_10839_),
    .B(\mem.mem_internal.code_mem[121][7] ));
 sg13g2_nand2_1 _17160_ (.Y(_10847_),
    .A(net1167),
    .B(_10828_));
 sg13g2_o21ai_1 _17161_ (.B1(_10847_),
    .Y(_00313_),
    .A1(net275),
    .A2(_10846_));
 sg13g2_nor2_1 _17162_ (.A(net550),
    .B(net468),
    .Y(_10848_));
 sg13g2_buf_2 _17163_ (.A(_10848_),
    .X(_10849_));
 sg13g2_buf_1 _17164_ (.A(_10849_),
    .X(_10850_));
 sg13g2_nand2_1 _17165_ (.Y(_10851_),
    .A(net760),
    .B(\mem.mem_internal.code_mem[122][0] ));
 sg13g2_nand2_1 _17166_ (.Y(_10852_),
    .A(net1174),
    .B(_10850_));
 sg13g2_o21ai_1 _17167_ (.B1(_10852_),
    .Y(_00314_),
    .A1(_10850_),
    .A2(_10851_));
 sg13g2_nand2_1 _17168_ (.Y(_10853_),
    .A(net760),
    .B(\mem.mem_internal.code_mem[122][1] ));
 sg13g2_nand2_1 _17169_ (.Y(_10854_),
    .A(net1173),
    .B(net274));
 sg13g2_o21ai_1 _17170_ (.B1(_10854_),
    .Y(_00315_),
    .A1(net274),
    .A2(_10853_));
 sg13g2_nand2_1 _17171_ (.Y(_10855_),
    .A(net760),
    .B(\mem.mem_internal.code_mem[122][2] ));
 sg13g2_nand2_1 _17172_ (.Y(_10856_),
    .A(net1172),
    .B(_10849_));
 sg13g2_o21ai_1 _17173_ (.B1(_10856_),
    .Y(_00316_),
    .A1(net274),
    .A2(_10855_));
 sg13g2_nand2_1 _17174_ (.Y(_10857_),
    .A(net760),
    .B(\mem.mem_internal.code_mem[122][3] ));
 sg13g2_nand2_1 _17175_ (.Y(_10858_),
    .A(net1171),
    .B(_10849_));
 sg13g2_o21ai_1 _17176_ (.B1(_10858_),
    .Y(_00317_),
    .A1(net274),
    .A2(_10857_));
 sg13g2_nand2_1 _17177_ (.Y(_10859_),
    .A(net760),
    .B(\mem.mem_internal.code_mem[122][4] ));
 sg13g2_nand2_1 _17178_ (.Y(_10860_),
    .A(net1170),
    .B(_10849_));
 sg13g2_o21ai_1 _17179_ (.B1(_10860_),
    .Y(_00318_),
    .A1(net274),
    .A2(_10859_));
 sg13g2_nand2_1 _17180_ (.Y(_10861_),
    .A(net760),
    .B(\mem.mem_internal.code_mem[122][5] ));
 sg13g2_nand2_1 _17181_ (.Y(_10862_),
    .A(net1169),
    .B(_10849_));
 sg13g2_o21ai_1 _17182_ (.B1(_10862_),
    .Y(_00319_),
    .A1(net274),
    .A2(_10861_));
 sg13g2_buf_1 _17183_ (.A(_10838_),
    .X(_10863_));
 sg13g2_nand2_1 _17184_ (.Y(_10864_),
    .A(net759),
    .B(\mem.mem_internal.code_mem[122][6] ));
 sg13g2_nand2_1 _17185_ (.Y(_10865_),
    .A(net1168),
    .B(_10849_));
 sg13g2_o21ai_1 _17186_ (.B1(_10865_),
    .Y(_00320_),
    .A1(net274),
    .A2(_10864_));
 sg13g2_nand2_1 _17187_ (.Y(_10866_),
    .A(net759),
    .B(\mem.mem_internal.code_mem[122][7] ));
 sg13g2_nand2_1 _17188_ (.Y(_10867_),
    .A(_10766_),
    .B(_10849_));
 sg13g2_o21ai_1 _17189_ (.B1(_10867_),
    .Y(_00321_),
    .A1(net274),
    .A2(_10866_));
 sg13g2_nor2_1 _17190_ (.A(net549),
    .B(net468),
    .Y(_10868_));
 sg13g2_buf_2 _17191_ (.A(_10868_),
    .X(_10869_));
 sg13g2_buf_1 _17192_ (.A(_10869_),
    .X(_10870_));
 sg13g2_nand2_1 _17193_ (.Y(_10871_),
    .A(net759),
    .B(\mem.mem_internal.code_mem[123][0] ));
 sg13g2_nand2_1 _17194_ (.Y(_10872_),
    .A(_10744_),
    .B(_10870_));
 sg13g2_o21ai_1 _17195_ (.B1(_10872_),
    .Y(_00322_),
    .A1(net273),
    .A2(_10871_));
 sg13g2_nand2_1 _17196_ (.Y(_10873_),
    .A(net759),
    .B(\mem.mem_internal.code_mem[123][1] ));
 sg13g2_nand2_1 _17197_ (.Y(_10874_),
    .A(net1173),
    .B(net273));
 sg13g2_o21ai_1 _17198_ (.B1(_10874_),
    .Y(_00323_),
    .A1(net273),
    .A2(_10873_));
 sg13g2_nand2_1 _17199_ (.Y(_10875_),
    .A(net759),
    .B(\mem.mem_internal.code_mem[123][2] ));
 sg13g2_nand2_1 _17200_ (.Y(_10876_),
    .A(net1172),
    .B(_10869_));
 sg13g2_o21ai_1 _17201_ (.B1(_10876_),
    .Y(_00324_),
    .A1(net273),
    .A2(_10875_));
 sg13g2_nand2_1 _17202_ (.Y(_10877_),
    .A(net759),
    .B(\mem.mem_internal.code_mem[123][3] ));
 sg13g2_nand2_1 _17203_ (.Y(_10878_),
    .A(net1171),
    .B(_10869_));
 sg13g2_o21ai_1 _17204_ (.B1(_10878_),
    .Y(_00325_),
    .A1(_10870_),
    .A2(_10877_));
 sg13g2_nand2_1 _17205_ (.Y(_10879_),
    .A(_10863_),
    .B(\mem.mem_internal.code_mem[123][4] ));
 sg13g2_nand2_1 _17206_ (.Y(_10880_),
    .A(net1170),
    .B(_10869_));
 sg13g2_o21ai_1 _17207_ (.B1(_10880_),
    .Y(_00326_),
    .A1(net273),
    .A2(_10879_));
 sg13g2_nand2_1 _17208_ (.Y(_10881_),
    .A(_10863_),
    .B(\mem.mem_internal.code_mem[123][5] ));
 sg13g2_nand2_1 _17209_ (.Y(_10882_),
    .A(net1169),
    .B(_10869_));
 sg13g2_o21ai_1 _17210_ (.B1(_10882_),
    .Y(_00327_),
    .A1(net273),
    .A2(_10881_));
 sg13g2_nand2_1 _17211_ (.Y(_10883_),
    .A(net759),
    .B(\mem.mem_internal.code_mem[123][6] ));
 sg13g2_nand2_1 _17212_ (.Y(_10884_),
    .A(net1168),
    .B(_10869_));
 sg13g2_o21ai_1 _17213_ (.B1(_10884_),
    .Y(_00328_),
    .A1(net273),
    .A2(_10883_));
 sg13g2_nand2_1 _17214_ (.Y(_10885_),
    .A(net759),
    .B(\mem.mem_internal.code_mem[123][7] ));
 sg13g2_nand2_1 _17215_ (.Y(_10886_),
    .A(_10766_),
    .B(_10869_));
 sg13g2_o21ai_1 _17216_ (.B1(_10886_),
    .Y(_00329_),
    .A1(net273),
    .A2(_10885_));
 sg13g2_nor2_1 _17217_ (.A(net773),
    .B(net468),
    .Y(_10887_));
 sg13g2_buf_2 _17218_ (.A(_10887_),
    .X(_10888_));
 sg13g2_buf_1 _17219_ (.A(_10888_),
    .X(_10889_));
 sg13g2_buf_1 _17220_ (.A(_10838_),
    .X(_10890_));
 sg13g2_nand2_1 _17221_ (.Y(_10891_),
    .A(net758),
    .B(\mem.mem_internal.code_mem[124][0] ));
 sg13g2_nand2_1 _17222_ (.Y(_10892_),
    .A(net1174),
    .B(net272));
 sg13g2_o21ai_1 _17223_ (.B1(_10892_),
    .Y(_00330_),
    .A1(net272),
    .A2(_10891_));
 sg13g2_nand2_1 _17224_ (.Y(_10893_),
    .A(net758),
    .B(\mem.mem_internal.code_mem[124][1] ));
 sg13g2_nand2_1 _17225_ (.Y(_10894_),
    .A(net1173),
    .B(net272));
 sg13g2_o21ai_1 _17226_ (.B1(_10894_),
    .Y(_00331_),
    .A1(net272),
    .A2(_10893_));
 sg13g2_nand2_1 _17227_ (.Y(_10895_),
    .A(net758),
    .B(\mem.mem_internal.code_mem[124][2] ));
 sg13g2_nand2_1 _17228_ (.Y(_10896_),
    .A(net1172),
    .B(_10888_));
 sg13g2_o21ai_1 _17229_ (.B1(_10896_),
    .Y(_00332_),
    .A1(net272),
    .A2(_10895_));
 sg13g2_nand2_1 _17230_ (.Y(_10897_),
    .A(net758),
    .B(\mem.mem_internal.code_mem[124][3] ));
 sg13g2_nand2_1 _17231_ (.Y(_10898_),
    .A(net1171),
    .B(_10888_));
 sg13g2_o21ai_1 _17232_ (.B1(_10898_),
    .Y(_00333_),
    .A1(_10889_),
    .A2(_10897_));
 sg13g2_nand2_1 _17233_ (.Y(_10899_),
    .A(net758),
    .B(\mem.mem_internal.code_mem[124][4] ));
 sg13g2_nand2_1 _17234_ (.Y(_10900_),
    .A(net1170),
    .B(_10888_));
 sg13g2_o21ai_1 _17235_ (.B1(_10900_),
    .Y(_00334_),
    .A1(net272),
    .A2(_10899_));
 sg13g2_nand2_1 _17236_ (.Y(_10901_),
    .A(_10890_),
    .B(\mem.mem_internal.code_mem[124][5] ));
 sg13g2_nand2_1 _17237_ (.Y(_10902_),
    .A(net1169),
    .B(_10888_));
 sg13g2_o21ai_1 _17238_ (.B1(_10902_),
    .Y(_00335_),
    .A1(net272),
    .A2(_10901_));
 sg13g2_nand2_1 _17239_ (.Y(_10903_),
    .A(net758),
    .B(\mem.mem_internal.code_mem[124][6] ));
 sg13g2_nand2_1 _17240_ (.Y(_10904_),
    .A(net1168),
    .B(_10888_));
 sg13g2_o21ai_1 _17241_ (.B1(_10904_),
    .Y(_00336_),
    .A1(net272),
    .A2(_10903_));
 sg13g2_nand2_1 _17242_ (.Y(_10905_),
    .A(_10890_),
    .B(\mem.mem_internal.code_mem[124][7] ));
 sg13g2_nand2_1 _17243_ (.Y(_10906_),
    .A(net1167),
    .B(_10888_));
 sg13g2_o21ai_1 _17244_ (.B1(_10906_),
    .Y(_00337_),
    .A1(_10889_),
    .A2(_10905_));
 sg13g2_nor2_1 _17245_ (.A(net548),
    .B(_10609_),
    .Y(_10907_));
 sg13g2_buf_2 _17246_ (.A(_10907_),
    .X(_10908_));
 sg13g2_buf_1 _17247_ (.A(_10908_),
    .X(_10909_));
 sg13g2_nand2_1 _17248_ (.Y(_10910_),
    .A(net758),
    .B(\mem.mem_internal.code_mem[125][0] ));
 sg13g2_nand2_1 _17249_ (.Y(_10911_),
    .A(net1174),
    .B(_10909_));
 sg13g2_o21ai_1 _17250_ (.B1(_10911_),
    .Y(_00338_),
    .A1(_10909_),
    .A2(_10910_));
 sg13g2_nand2_1 _17251_ (.Y(_10912_),
    .A(net758),
    .B(\mem.mem_internal.code_mem[125][1] ));
 sg13g2_nand2_1 _17252_ (.Y(_10913_),
    .A(net1173),
    .B(net393));
 sg13g2_o21ai_1 _17253_ (.B1(_10913_),
    .Y(_00339_),
    .A1(net393),
    .A2(_10912_));
 sg13g2_buf_1 _17254_ (.A(_10838_),
    .X(_10914_));
 sg13g2_nand2_1 _17255_ (.Y(_10915_),
    .A(net757),
    .B(\mem.mem_internal.code_mem[125][2] ));
 sg13g2_nand2_1 _17256_ (.Y(_10916_),
    .A(net1172),
    .B(_10908_));
 sg13g2_o21ai_1 _17257_ (.B1(_10916_),
    .Y(_00340_),
    .A1(net393),
    .A2(_10915_));
 sg13g2_nand2_1 _17258_ (.Y(_10917_),
    .A(net757),
    .B(\mem.mem_internal.code_mem[125][3] ));
 sg13g2_nand2_1 _17259_ (.Y(_10918_),
    .A(net1171),
    .B(_10908_));
 sg13g2_o21ai_1 _17260_ (.B1(_10918_),
    .Y(_00341_),
    .A1(net393),
    .A2(_10917_));
 sg13g2_nand2_1 _17261_ (.Y(_10919_),
    .A(net757),
    .B(\mem.mem_internal.code_mem[125][4] ));
 sg13g2_nand2_1 _17262_ (.Y(_10920_),
    .A(net1170),
    .B(_10908_));
 sg13g2_o21ai_1 _17263_ (.B1(_10920_),
    .Y(_00342_),
    .A1(net393),
    .A2(_10919_));
 sg13g2_nand2_1 _17264_ (.Y(_10921_),
    .A(net757),
    .B(\mem.mem_internal.code_mem[125][5] ));
 sg13g2_nand2_1 _17265_ (.Y(_10922_),
    .A(net1169),
    .B(_10908_));
 sg13g2_o21ai_1 _17266_ (.B1(_10922_),
    .Y(_00343_),
    .A1(net393),
    .A2(_10921_));
 sg13g2_nand2_1 _17267_ (.Y(_10923_),
    .A(net757),
    .B(\mem.mem_internal.code_mem[125][6] ));
 sg13g2_nand2_1 _17268_ (.Y(_10924_),
    .A(net1168),
    .B(_10908_));
 sg13g2_o21ai_1 _17269_ (.B1(_10924_),
    .Y(_00344_),
    .A1(net393),
    .A2(_10923_));
 sg13g2_nand2_1 _17270_ (.Y(_10925_),
    .A(_10914_),
    .B(\mem.mem_internal.code_mem[125][7] ));
 sg13g2_nand2_1 _17271_ (.Y(_10926_),
    .A(net1167),
    .B(_10908_));
 sg13g2_o21ai_1 _17272_ (.B1(_10926_),
    .Y(_00345_),
    .A1(net393),
    .A2(_10925_));
 sg13g2_nor2_1 _17273_ (.A(net547),
    .B(_10609_),
    .Y(_10927_));
 sg13g2_buf_2 _17274_ (.A(_10927_),
    .X(_10928_));
 sg13g2_buf_1 _17275_ (.A(_10928_),
    .X(_10929_));
 sg13g2_nand2_1 _17276_ (.Y(_10930_),
    .A(net757),
    .B(\mem.mem_internal.code_mem[126][0] ));
 sg13g2_nand2_1 _17277_ (.Y(_10931_),
    .A(net1174),
    .B(net392));
 sg13g2_o21ai_1 _17278_ (.B1(_10931_),
    .Y(_00346_),
    .A1(net392),
    .A2(_10930_));
 sg13g2_nand2_1 _17279_ (.Y(_10932_),
    .A(net757),
    .B(\mem.mem_internal.code_mem[126][1] ));
 sg13g2_nand2_1 _17280_ (.Y(_10933_),
    .A(net1173),
    .B(net392));
 sg13g2_o21ai_1 _17281_ (.B1(_10933_),
    .Y(_00347_),
    .A1(net392),
    .A2(_10932_));
 sg13g2_nand2_1 _17282_ (.Y(_10934_),
    .A(net757),
    .B(\mem.mem_internal.code_mem[126][2] ));
 sg13g2_nand2_1 _17283_ (.Y(_10935_),
    .A(net1172),
    .B(_10928_));
 sg13g2_o21ai_1 _17284_ (.B1(_10935_),
    .Y(_00348_),
    .A1(net392),
    .A2(_10934_));
 sg13g2_nand2_1 _17285_ (.Y(_10936_),
    .A(_10914_),
    .B(\mem.mem_internal.code_mem[126][3] ));
 sg13g2_nand2_1 _17286_ (.Y(_10937_),
    .A(net1171),
    .B(_10928_));
 sg13g2_o21ai_1 _17287_ (.B1(_10937_),
    .Y(_00349_),
    .A1(_10929_),
    .A2(_10936_));
 sg13g2_buf_1 _17288_ (.A(_10838_),
    .X(_10938_));
 sg13g2_nand2_1 _17289_ (.Y(_10939_),
    .A(net756),
    .B(\mem.mem_internal.code_mem[126][4] ));
 sg13g2_nand2_1 _17290_ (.Y(_10940_),
    .A(net1170),
    .B(_10928_));
 sg13g2_o21ai_1 _17291_ (.B1(_10940_),
    .Y(_00350_),
    .A1(net392),
    .A2(_10939_));
 sg13g2_nand2_1 _17292_ (.Y(_10941_),
    .A(net756),
    .B(\mem.mem_internal.code_mem[126][5] ));
 sg13g2_nand2_1 _17293_ (.Y(_10942_),
    .A(net1169),
    .B(_10928_));
 sg13g2_o21ai_1 _17294_ (.B1(_10942_),
    .Y(_00351_),
    .A1(net392),
    .A2(_10941_));
 sg13g2_nand2_1 _17295_ (.Y(_10943_),
    .A(net756),
    .B(\mem.mem_internal.code_mem[126][6] ));
 sg13g2_nand2_1 _17296_ (.Y(_10944_),
    .A(net1168),
    .B(_10928_));
 sg13g2_o21ai_1 _17297_ (.B1(_10944_),
    .Y(_00352_),
    .A1(net392),
    .A2(_10943_));
 sg13g2_nand2_1 _17298_ (.Y(_10945_),
    .A(net756),
    .B(\mem.mem_internal.code_mem[126][7] ));
 sg13g2_nand2_1 _17299_ (.Y(_10946_),
    .A(net1167),
    .B(_10928_));
 sg13g2_o21ai_1 _17300_ (.B1(_10946_),
    .Y(_00353_),
    .A1(_10929_),
    .A2(_10945_));
 sg13g2_nor2_1 _17301_ (.A(net770),
    .B(_10609_),
    .Y(_10947_));
 sg13g2_buf_2 _17302_ (.A(_10947_),
    .X(_10948_));
 sg13g2_buf_1 _17303_ (.A(_10948_),
    .X(_10949_));
 sg13g2_nand2_1 _17304_ (.Y(_10950_),
    .A(_10938_),
    .B(\mem.mem_internal.code_mem[127][0] ));
 sg13g2_buf_1 _17305_ (.A(net1268),
    .X(_10951_));
 sg13g2_nand2_1 _17306_ (.Y(_10952_),
    .A(_10951_),
    .B(_10949_));
 sg13g2_o21ai_1 _17307_ (.B1(_10952_),
    .Y(_00354_),
    .A1(net391),
    .A2(_10950_));
 sg13g2_nand2_1 _17308_ (.Y(_10953_),
    .A(net756),
    .B(\mem.mem_internal.code_mem[127][1] ));
 sg13g2_buf_1 _17309_ (.A(net1267),
    .X(_10954_));
 sg13g2_nand2_1 _17310_ (.Y(_10955_),
    .A(net1165),
    .B(net391));
 sg13g2_o21ai_1 _17311_ (.B1(_10955_),
    .Y(_00355_),
    .A1(net391),
    .A2(_10953_));
 sg13g2_nand2_1 _17312_ (.Y(_10956_),
    .A(net756),
    .B(\mem.mem_internal.code_mem[127][2] ));
 sg13g2_buf_1 _17313_ (.A(net1266),
    .X(_10957_));
 sg13g2_nand2_1 _17314_ (.Y(_10958_),
    .A(_10957_),
    .B(_10948_));
 sg13g2_o21ai_1 _17315_ (.B1(_10958_),
    .Y(_00356_),
    .A1(net391),
    .A2(_10956_));
 sg13g2_nand2_1 _17316_ (.Y(_10959_),
    .A(_10938_),
    .B(\mem.mem_internal.code_mem[127][3] ));
 sg13g2_buf_1 _17317_ (.A(net1265),
    .X(_10960_));
 sg13g2_nand2_1 _17318_ (.Y(_10961_),
    .A(_10960_),
    .B(_10948_));
 sg13g2_o21ai_1 _17319_ (.B1(_10961_),
    .Y(_00357_),
    .A1(net391),
    .A2(_10959_));
 sg13g2_nand2_1 _17320_ (.Y(_10962_),
    .A(net756),
    .B(\mem.mem_internal.code_mem[127][4] ));
 sg13g2_buf_1 _17321_ (.A(net1264),
    .X(_10963_));
 sg13g2_nand2_1 _17322_ (.Y(_10964_),
    .A(_10963_),
    .B(_10948_));
 sg13g2_o21ai_1 _17323_ (.B1(_10964_),
    .Y(_00358_),
    .A1(net391),
    .A2(_10962_));
 sg13g2_nand2_1 _17324_ (.Y(_10965_),
    .A(net756),
    .B(\mem.mem_internal.code_mem[127][5] ));
 sg13g2_buf_1 _17325_ (.A(net1263),
    .X(_10966_));
 sg13g2_nand2_1 _17326_ (.Y(_10967_),
    .A(_10966_),
    .B(_10948_));
 sg13g2_o21ai_1 _17327_ (.B1(_10967_),
    .Y(_00359_),
    .A1(net391),
    .A2(_10965_));
 sg13g2_buf_1 _17328_ (.A(_10838_),
    .X(_10968_));
 sg13g2_nand2_1 _17329_ (.Y(_10969_),
    .A(net755),
    .B(\mem.mem_internal.code_mem[127][6] ));
 sg13g2_buf_1 _17330_ (.A(net1262),
    .X(_10970_));
 sg13g2_nand2_1 _17331_ (.Y(_10971_),
    .A(_10970_),
    .B(_10948_));
 sg13g2_o21ai_1 _17332_ (.B1(_10971_),
    .Y(_00360_),
    .A1(net391),
    .A2(_10969_));
 sg13g2_nand2_1 _17333_ (.Y(_10972_),
    .A(net755),
    .B(\mem.mem_internal.code_mem[127][7] ));
 sg13g2_buf_1 _17334_ (.A(net1261),
    .X(_10973_));
 sg13g2_nand2_1 _17335_ (.Y(_10974_),
    .A(_10973_),
    .B(_10948_));
 sg13g2_o21ai_1 _17336_ (.B1(_10974_),
    .Y(_00361_),
    .A1(_10949_),
    .A2(_10972_));
 sg13g2_nand2_1 _17337_ (.Y(_10975_),
    .A(net850),
    .B(\mem.mem_internal.code_mem[128][0] ));
 sg13g2_nor2b_1 _17338_ (.A(net1296),
    .B_N(net1297),
    .Y(_10976_));
 sg13g2_nand2_1 _17339_ (.Y(_10977_),
    .A(_10244_),
    .B(_10976_));
 sg13g2_buf_2 _17340_ (.A(_10977_),
    .X(_10978_));
 sg13g2_buf_1 _17341_ (.A(_10978_),
    .X(_10979_));
 sg13g2_nor2_1 _17342_ (.A(_10233_),
    .B(net467),
    .Y(_10980_));
 sg13g2_buf_2 _17343_ (.A(_10980_),
    .X(_10981_));
 sg13g2_buf_1 _17344_ (.A(_10981_),
    .X(_10982_));
 sg13g2_nand2_1 _17345_ (.Y(_10983_),
    .A(net1166),
    .B(_10982_));
 sg13g2_o21ai_1 _17346_ (.B1(_10983_),
    .Y(_00362_),
    .A1(_10975_),
    .A2(_10982_));
 sg13g2_nand2_1 _17347_ (.Y(_10984_),
    .A(net755),
    .B(\mem.mem_internal.code_mem[128][1] ));
 sg13g2_nand2_1 _17348_ (.Y(_10985_),
    .A(net1165),
    .B(net271));
 sg13g2_o21ai_1 _17349_ (.B1(_10985_),
    .Y(_00363_),
    .A1(net271),
    .A2(_10984_));
 sg13g2_nand2_1 _17350_ (.Y(_10986_),
    .A(_10968_),
    .B(\mem.mem_internal.code_mem[128][2] ));
 sg13g2_nand2_1 _17351_ (.Y(_10987_),
    .A(_10957_),
    .B(_10981_));
 sg13g2_o21ai_1 _17352_ (.B1(_10987_),
    .Y(_00364_),
    .A1(net271),
    .A2(_10986_));
 sg13g2_nand2_1 _17353_ (.Y(_10988_),
    .A(_10968_),
    .B(\mem.mem_internal.code_mem[128][3] ));
 sg13g2_nand2_1 _17354_ (.Y(_10989_),
    .A(_10960_),
    .B(_10981_));
 sg13g2_o21ai_1 _17355_ (.B1(_10989_),
    .Y(_00365_),
    .A1(net271),
    .A2(_10988_));
 sg13g2_nand2_1 _17356_ (.Y(_10990_),
    .A(net755),
    .B(\mem.mem_internal.code_mem[128][4] ));
 sg13g2_nand2_1 _17357_ (.Y(_10991_),
    .A(_10963_),
    .B(_10981_));
 sg13g2_o21ai_1 _17358_ (.B1(_10991_),
    .Y(_00366_),
    .A1(net271),
    .A2(_10990_));
 sg13g2_nand2_1 _17359_ (.Y(_10992_),
    .A(net755),
    .B(\mem.mem_internal.code_mem[128][5] ));
 sg13g2_nand2_1 _17360_ (.Y(_10993_),
    .A(_10966_),
    .B(_10981_));
 sg13g2_o21ai_1 _17361_ (.B1(_10993_),
    .Y(_00367_),
    .A1(net271),
    .A2(_10992_));
 sg13g2_nand2_1 _17362_ (.Y(_10994_),
    .A(net755),
    .B(\mem.mem_internal.code_mem[128][6] ));
 sg13g2_nand2_1 _17363_ (.Y(_10995_),
    .A(net1160),
    .B(_10981_));
 sg13g2_o21ai_1 _17364_ (.B1(_10995_),
    .Y(_00368_),
    .A1(net271),
    .A2(_10994_));
 sg13g2_nand2_1 _17365_ (.Y(_10996_),
    .A(net755),
    .B(\mem.mem_internal.code_mem[128][7] ));
 sg13g2_nand2_1 _17366_ (.Y(_10997_),
    .A(_10973_),
    .B(_10981_));
 sg13g2_o21ai_1 _17367_ (.B1(_10997_),
    .Y(_00369_),
    .A1(net271),
    .A2(_10996_));
 sg13g2_nand2_1 _17368_ (.Y(_10998_),
    .A(net850),
    .B(\mem.mem_internal.code_mem[129][0] ));
 sg13g2_nor2_1 _17369_ (.A(_10633_),
    .B(net467),
    .Y(_10999_));
 sg13g2_buf_2 _17370_ (.A(_10999_),
    .X(_11000_));
 sg13g2_buf_1 _17371_ (.A(_11000_),
    .X(_11001_));
 sg13g2_nand2_1 _17372_ (.Y(_11002_),
    .A(net1166),
    .B(net270));
 sg13g2_o21ai_1 _17373_ (.B1(_11002_),
    .Y(_00370_),
    .A1(_10998_),
    .A2(net270));
 sg13g2_nand2_1 _17374_ (.Y(_11003_),
    .A(net755),
    .B(\mem.mem_internal.code_mem[129][1] ));
 sg13g2_nand2_1 _17375_ (.Y(_11004_),
    .A(net1165),
    .B(net270));
 sg13g2_o21ai_1 _17376_ (.B1(_11004_),
    .Y(_00371_),
    .A1(net270),
    .A2(_11003_));
 sg13g2_buf_1 _17377_ (.A(_10838_),
    .X(_11005_));
 sg13g2_nand2_1 _17378_ (.Y(_11006_),
    .A(net754),
    .B(\mem.mem_internal.code_mem[129][2] ));
 sg13g2_nand2_1 _17379_ (.Y(_11007_),
    .A(net1164),
    .B(_11000_));
 sg13g2_o21ai_1 _17380_ (.B1(_11007_),
    .Y(_00372_),
    .A1(net270),
    .A2(_11006_));
 sg13g2_nand2_1 _17381_ (.Y(_11008_),
    .A(net754),
    .B(\mem.mem_internal.code_mem[129][3] ));
 sg13g2_nand2_1 _17382_ (.Y(_11009_),
    .A(net1163),
    .B(_11000_));
 sg13g2_o21ai_1 _17383_ (.B1(_11009_),
    .Y(_00373_),
    .A1(_11001_),
    .A2(_11008_));
 sg13g2_nand2_1 _17384_ (.Y(_11010_),
    .A(net754),
    .B(\mem.mem_internal.code_mem[129][4] ));
 sg13g2_nand2_1 _17385_ (.Y(_11011_),
    .A(net1162),
    .B(_11000_));
 sg13g2_o21ai_1 _17386_ (.B1(_11011_),
    .Y(_00374_),
    .A1(_11001_),
    .A2(_11010_));
 sg13g2_nand2_1 _17387_ (.Y(_11012_),
    .A(net754),
    .B(\mem.mem_internal.code_mem[129][5] ));
 sg13g2_nand2_1 _17388_ (.Y(_11013_),
    .A(net1161),
    .B(_11000_));
 sg13g2_o21ai_1 _17389_ (.B1(_11013_),
    .Y(_00375_),
    .A1(net270),
    .A2(_11012_));
 sg13g2_nand2_1 _17390_ (.Y(_11014_),
    .A(_11005_),
    .B(\mem.mem_internal.code_mem[129][6] ));
 sg13g2_nand2_1 _17391_ (.Y(_11015_),
    .A(net1160),
    .B(_11000_));
 sg13g2_o21ai_1 _17392_ (.B1(_11015_),
    .Y(_00376_),
    .A1(net270),
    .A2(_11014_));
 sg13g2_nand2_1 _17393_ (.Y(_11016_),
    .A(_11005_),
    .B(\mem.mem_internal.code_mem[129][7] ));
 sg13g2_nand2_1 _17394_ (.Y(_11017_),
    .A(net1159),
    .B(_11000_));
 sg13g2_o21ai_1 _17395_ (.B1(_11017_),
    .Y(_00377_),
    .A1(net270),
    .A2(_11016_));
 sg13g2_nand2_1 _17396_ (.Y(_11018_),
    .A(net850),
    .B(\mem.mem_internal.code_mem[12][0] ));
 sg13g2_nor2_1 _17397_ (.A(_10247_),
    .B(_10492_),
    .Y(_11019_));
 sg13g2_buf_2 _17398_ (.A(_11019_),
    .X(_11020_));
 sg13g2_buf_1 _17399_ (.A(_11020_),
    .X(_11021_));
 sg13g2_nand2_1 _17400_ (.Y(_11022_),
    .A(net1166),
    .B(net269));
 sg13g2_o21ai_1 _17401_ (.B1(_11022_),
    .Y(_00378_),
    .A1(_11018_),
    .A2(net269));
 sg13g2_nand2_1 _17402_ (.Y(_11023_),
    .A(net754),
    .B(\mem.mem_internal.code_mem[12][1] ));
 sg13g2_nand2_1 _17403_ (.Y(_11024_),
    .A(_10954_),
    .B(net269));
 sg13g2_o21ai_1 _17404_ (.B1(_11024_),
    .Y(_00379_),
    .A1(net269),
    .A2(_11023_));
 sg13g2_nand2_1 _17405_ (.Y(_11025_),
    .A(net754),
    .B(\mem.mem_internal.code_mem[12][2] ));
 sg13g2_nand2_1 _17406_ (.Y(_11026_),
    .A(net1164),
    .B(_11020_));
 sg13g2_o21ai_1 _17407_ (.B1(_11026_),
    .Y(_00380_),
    .A1(net269),
    .A2(_11025_));
 sg13g2_nand2_1 _17408_ (.Y(_11027_),
    .A(net754),
    .B(\mem.mem_internal.code_mem[12][3] ));
 sg13g2_nand2_1 _17409_ (.Y(_11028_),
    .A(net1163),
    .B(_11020_));
 sg13g2_o21ai_1 _17410_ (.B1(_11028_),
    .Y(_00381_),
    .A1(_11021_),
    .A2(_11027_));
 sg13g2_nand2_1 _17411_ (.Y(_11029_),
    .A(net754),
    .B(\mem.mem_internal.code_mem[12][4] ));
 sg13g2_nand2_1 _17412_ (.Y(_11030_),
    .A(net1162),
    .B(_11020_));
 sg13g2_o21ai_1 _17413_ (.B1(_11030_),
    .Y(_00382_),
    .A1(_11021_),
    .A2(_11029_));
 sg13g2_buf_1 _17414_ (.A(_10415_),
    .X(_11031_));
 sg13g2_buf_1 _17415_ (.A(_11031_),
    .X(_11032_));
 sg13g2_nand2_1 _17416_ (.Y(_11033_),
    .A(net753),
    .B(\mem.mem_internal.code_mem[12][5] ));
 sg13g2_nand2_1 _17417_ (.Y(_11034_),
    .A(net1161),
    .B(_11020_));
 sg13g2_o21ai_1 _17418_ (.B1(_11034_),
    .Y(_00383_),
    .A1(net269),
    .A2(_11033_));
 sg13g2_nand2_1 _17419_ (.Y(_11035_),
    .A(net753),
    .B(\mem.mem_internal.code_mem[12][6] ));
 sg13g2_nand2_1 _17420_ (.Y(_11036_),
    .A(net1160),
    .B(_11020_));
 sg13g2_o21ai_1 _17421_ (.B1(_11036_),
    .Y(_00384_),
    .A1(net269),
    .A2(_11035_));
 sg13g2_nand2_1 _17422_ (.Y(_11037_),
    .A(net753),
    .B(\mem.mem_internal.code_mem[12][7] ));
 sg13g2_nand2_1 _17423_ (.Y(_11038_),
    .A(net1159),
    .B(_11020_));
 sg13g2_o21ai_1 _17424_ (.B1(_11038_),
    .Y(_00385_),
    .A1(net269),
    .A2(_11037_));
 sg13g2_nand2_1 _17425_ (.Y(_11039_),
    .A(_10488_),
    .B(\mem.mem_internal.code_mem[130][0] ));
 sg13g2_nor2_1 _17426_ (.A(_10657_),
    .B(net467),
    .Y(_11040_));
 sg13g2_buf_2 _17427_ (.A(_11040_),
    .X(_11041_));
 sg13g2_buf_1 _17428_ (.A(_11041_),
    .X(_11042_));
 sg13g2_nand2_1 _17429_ (.Y(_11043_),
    .A(_10951_),
    .B(net268));
 sg13g2_o21ai_1 _17430_ (.B1(_11043_),
    .Y(_00386_),
    .A1(_11039_),
    .A2(net268));
 sg13g2_nand2_1 _17431_ (.Y(_11044_),
    .A(net753),
    .B(\mem.mem_internal.code_mem[130][1] ));
 sg13g2_nand2_1 _17432_ (.Y(_11045_),
    .A(_10954_),
    .B(net268));
 sg13g2_o21ai_1 _17433_ (.B1(_11045_),
    .Y(_00387_),
    .A1(net268),
    .A2(_11044_));
 sg13g2_nand2_1 _17434_ (.Y(_11046_),
    .A(net753),
    .B(\mem.mem_internal.code_mem[130][2] ));
 sg13g2_nand2_1 _17435_ (.Y(_11047_),
    .A(net1164),
    .B(_11041_));
 sg13g2_o21ai_1 _17436_ (.B1(_11047_),
    .Y(_00388_),
    .A1(_11042_),
    .A2(_11046_));
 sg13g2_nand2_1 _17437_ (.Y(_11048_),
    .A(net753),
    .B(\mem.mem_internal.code_mem[130][3] ));
 sg13g2_nand2_1 _17438_ (.Y(_11049_),
    .A(net1163),
    .B(_11041_));
 sg13g2_o21ai_1 _17439_ (.B1(_11049_),
    .Y(_00389_),
    .A1(_11042_),
    .A2(_11048_));
 sg13g2_nand2_1 _17440_ (.Y(_11050_),
    .A(net753),
    .B(\mem.mem_internal.code_mem[130][4] ));
 sg13g2_nand2_1 _17441_ (.Y(_11051_),
    .A(net1162),
    .B(_11041_));
 sg13g2_o21ai_1 _17442_ (.B1(_11051_),
    .Y(_00390_),
    .A1(net268),
    .A2(_11050_));
 sg13g2_nand2_1 _17443_ (.Y(_11052_),
    .A(net753),
    .B(\mem.mem_internal.code_mem[130][5] ));
 sg13g2_nand2_1 _17444_ (.Y(_11053_),
    .A(net1161),
    .B(_11041_));
 sg13g2_o21ai_1 _17445_ (.B1(_11053_),
    .Y(_00391_),
    .A1(net268),
    .A2(_11052_));
 sg13g2_nand2_1 _17446_ (.Y(_11054_),
    .A(_11032_),
    .B(\mem.mem_internal.code_mem[130][6] ));
 sg13g2_nand2_1 _17447_ (.Y(_11055_),
    .A(_10970_),
    .B(_11041_));
 sg13g2_o21ai_1 _17448_ (.B1(_11055_),
    .Y(_00392_),
    .A1(net268),
    .A2(_11054_));
 sg13g2_nand2_1 _17449_ (.Y(_11056_),
    .A(_11032_),
    .B(\mem.mem_internal.code_mem[130][7] ));
 sg13g2_nand2_1 _17450_ (.Y(_11057_),
    .A(net1159),
    .B(_11041_));
 sg13g2_o21ai_1 _17451_ (.B1(_11057_),
    .Y(_00393_),
    .A1(net268),
    .A2(_11056_));
 sg13g2_buf_1 _17452_ (.A(net1273),
    .X(_11058_));
 sg13g2_buf_1 _17453_ (.A(_11058_),
    .X(_11059_));
 sg13g2_nand2_1 _17454_ (.Y(_11060_),
    .A(net849),
    .B(\mem.mem_internal.code_mem[131][0] ));
 sg13g2_nor2_1 _17455_ (.A(_10680_),
    .B(net467),
    .Y(_11061_));
 sg13g2_buf_2 _17456_ (.A(_11061_),
    .X(_11062_));
 sg13g2_buf_1 _17457_ (.A(_11062_),
    .X(_11063_));
 sg13g2_nand2_1 _17458_ (.Y(_11064_),
    .A(net1166),
    .B(_11063_));
 sg13g2_o21ai_1 _17459_ (.B1(_11064_),
    .Y(_00394_),
    .A1(_11060_),
    .A2(_11063_));
 sg13g2_buf_1 _17460_ (.A(_11031_),
    .X(_11065_));
 sg13g2_nand2_1 _17461_ (.Y(_11066_),
    .A(net752),
    .B(\mem.mem_internal.code_mem[131][1] ));
 sg13g2_nand2_1 _17462_ (.Y(_11067_),
    .A(net1165),
    .B(net267));
 sg13g2_o21ai_1 _17463_ (.B1(_11067_),
    .Y(_00395_),
    .A1(net267),
    .A2(_11066_));
 sg13g2_nand2_1 _17464_ (.Y(_11068_),
    .A(net752),
    .B(\mem.mem_internal.code_mem[131][2] ));
 sg13g2_nand2_1 _17465_ (.Y(_11069_),
    .A(net1164),
    .B(_11062_));
 sg13g2_o21ai_1 _17466_ (.B1(_11069_),
    .Y(_00396_),
    .A1(net267),
    .A2(_11068_));
 sg13g2_nand2_1 _17467_ (.Y(_11070_),
    .A(net752),
    .B(\mem.mem_internal.code_mem[131][3] ));
 sg13g2_nand2_1 _17468_ (.Y(_11071_),
    .A(net1163),
    .B(_11062_));
 sg13g2_o21ai_1 _17469_ (.B1(_11071_),
    .Y(_00397_),
    .A1(net267),
    .A2(_11070_));
 sg13g2_nand2_1 _17470_ (.Y(_11072_),
    .A(net752),
    .B(\mem.mem_internal.code_mem[131][4] ));
 sg13g2_nand2_1 _17471_ (.Y(_11073_),
    .A(net1162),
    .B(_11062_));
 sg13g2_o21ai_1 _17472_ (.B1(_11073_),
    .Y(_00398_),
    .A1(net267),
    .A2(_11072_));
 sg13g2_nand2_1 _17473_ (.Y(_11074_),
    .A(net752),
    .B(\mem.mem_internal.code_mem[131][5] ));
 sg13g2_nand2_1 _17474_ (.Y(_11075_),
    .A(net1161),
    .B(_11062_));
 sg13g2_o21ai_1 _17475_ (.B1(_11075_),
    .Y(_00399_),
    .A1(net267),
    .A2(_11074_));
 sg13g2_nand2_1 _17476_ (.Y(_11076_),
    .A(_11065_),
    .B(\mem.mem_internal.code_mem[131][6] ));
 sg13g2_nand2_1 _17477_ (.Y(_11077_),
    .A(net1160),
    .B(_11062_));
 sg13g2_o21ai_1 _17478_ (.B1(_11077_),
    .Y(_00400_),
    .A1(net267),
    .A2(_11076_));
 sg13g2_nand2_1 _17479_ (.Y(_11078_),
    .A(_11065_),
    .B(\mem.mem_internal.code_mem[131][7] ));
 sg13g2_nand2_1 _17480_ (.Y(_11079_),
    .A(net1159),
    .B(_11062_));
 sg13g2_o21ai_1 _17481_ (.B1(_11079_),
    .Y(_00401_),
    .A1(net267),
    .A2(_11078_));
 sg13g2_nand2_1 _17482_ (.Y(_11080_),
    .A(net849),
    .B(\mem.mem_internal.code_mem[132][0] ));
 sg13g2_nor2_1 _17483_ (.A(_10296_),
    .B(net467),
    .Y(_11081_));
 sg13g2_buf_2 _17484_ (.A(_11081_),
    .X(_11082_));
 sg13g2_buf_1 _17485_ (.A(_11082_),
    .X(_11083_));
 sg13g2_nand2_1 _17486_ (.Y(_11084_),
    .A(net1166),
    .B(net266));
 sg13g2_o21ai_1 _17487_ (.B1(_11084_),
    .Y(_00402_),
    .A1(_11080_),
    .A2(net266));
 sg13g2_nand2_1 _17488_ (.Y(_11085_),
    .A(net752),
    .B(\mem.mem_internal.code_mem[132][1] ));
 sg13g2_nand2_1 _17489_ (.Y(_11086_),
    .A(net1165),
    .B(net266));
 sg13g2_o21ai_1 _17490_ (.B1(_11086_),
    .Y(_00403_),
    .A1(net266),
    .A2(_11085_));
 sg13g2_nand2_1 _17491_ (.Y(_11087_),
    .A(net752),
    .B(\mem.mem_internal.code_mem[132][2] ));
 sg13g2_nand2_1 _17492_ (.Y(_11088_),
    .A(net1164),
    .B(_11082_));
 sg13g2_o21ai_1 _17493_ (.B1(_11088_),
    .Y(_00404_),
    .A1(net266),
    .A2(_11087_));
 sg13g2_nand2_1 _17494_ (.Y(_11089_),
    .A(net752),
    .B(\mem.mem_internal.code_mem[132][3] ));
 sg13g2_nand2_1 _17495_ (.Y(_11090_),
    .A(net1163),
    .B(_11082_));
 sg13g2_o21ai_1 _17496_ (.B1(_11090_),
    .Y(_00405_),
    .A1(net266),
    .A2(_11089_));
 sg13g2_buf_1 _17497_ (.A(_11031_),
    .X(_11091_));
 sg13g2_nand2_1 _17498_ (.Y(_11092_),
    .A(net751),
    .B(\mem.mem_internal.code_mem[132][4] ));
 sg13g2_nand2_1 _17499_ (.Y(_11093_),
    .A(net1162),
    .B(_11082_));
 sg13g2_o21ai_1 _17500_ (.B1(_11093_),
    .Y(_00406_),
    .A1(net266),
    .A2(_11092_));
 sg13g2_nand2_1 _17501_ (.Y(_11094_),
    .A(net751),
    .B(\mem.mem_internal.code_mem[132][5] ));
 sg13g2_nand2_1 _17502_ (.Y(_11095_),
    .A(net1161),
    .B(_11082_));
 sg13g2_o21ai_1 _17503_ (.B1(_11095_),
    .Y(_00407_),
    .A1(_11083_),
    .A2(_11094_));
 sg13g2_nand2_1 _17504_ (.Y(_11096_),
    .A(net751),
    .B(\mem.mem_internal.code_mem[132][6] ));
 sg13g2_nand2_1 _17505_ (.Y(_11097_),
    .A(net1160),
    .B(_11082_));
 sg13g2_o21ai_1 _17506_ (.B1(_11097_),
    .Y(_00408_),
    .A1(_11083_),
    .A2(_11096_));
 sg13g2_nand2_1 _17507_ (.Y(_11098_),
    .A(net751),
    .B(\mem.mem_internal.code_mem[132][7] ));
 sg13g2_nand2_1 _17508_ (.Y(_11099_),
    .A(net1159),
    .B(_11082_));
 sg13g2_o21ai_1 _17509_ (.B1(_11099_),
    .Y(_00409_),
    .A1(net266),
    .A2(_11098_));
 sg13g2_nand2_1 _17510_ (.Y(_11100_),
    .A(net849),
    .B(\mem.mem_internal.code_mem[133][0] ));
 sg13g2_nor2_1 _17511_ (.A(_10326_),
    .B(_10979_),
    .Y(_11101_));
 sg13g2_buf_2 _17512_ (.A(_11101_),
    .X(_11102_));
 sg13g2_buf_1 _17513_ (.A(_11102_),
    .X(_11103_));
 sg13g2_nand2_1 _17514_ (.Y(_11104_),
    .A(net1166),
    .B(net265));
 sg13g2_o21ai_1 _17515_ (.B1(_11104_),
    .Y(_00410_),
    .A1(_11100_),
    .A2(net265));
 sg13g2_nand2_1 _17516_ (.Y(_11105_),
    .A(net751),
    .B(\mem.mem_internal.code_mem[133][1] ));
 sg13g2_nand2_1 _17517_ (.Y(_11106_),
    .A(net1165),
    .B(net265));
 sg13g2_o21ai_1 _17518_ (.B1(_11106_),
    .Y(_00411_),
    .A1(net265),
    .A2(_11105_));
 sg13g2_nand2_1 _17519_ (.Y(_11107_),
    .A(net751),
    .B(\mem.mem_internal.code_mem[133][2] ));
 sg13g2_nand2_1 _17520_ (.Y(_11108_),
    .A(net1164),
    .B(_11102_));
 sg13g2_o21ai_1 _17521_ (.B1(_11108_),
    .Y(_00412_),
    .A1(net265),
    .A2(_11107_));
 sg13g2_nand2_1 _17522_ (.Y(_11109_),
    .A(_11091_),
    .B(\mem.mem_internal.code_mem[133][3] ));
 sg13g2_nand2_1 _17523_ (.Y(_11110_),
    .A(net1163),
    .B(_11102_));
 sg13g2_o21ai_1 _17524_ (.B1(_11110_),
    .Y(_00413_),
    .A1(net265),
    .A2(_11109_));
 sg13g2_nand2_1 _17525_ (.Y(_11111_),
    .A(net751),
    .B(\mem.mem_internal.code_mem[133][4] ));
 sg13g2_nand2_1 _17526_ (.Y(_11112_),
    .A(net1162),
    .B(_11102_));
 sg13g2_o21ai_1 _17527_ (.B1(_11112_),
    .Y(_00414_),
    .A1(net265),
    .A2(_11111_));
 sg13g2_nand2_1 _17528_ (.Y(_11113_),
    .A(_11091_),
    .B(\mem.mem_internal.code_mem[133][5] ));
 sg13g2_nand2_1 _17529_ (.Y(_11114_),
    .A(net1161),
    .B(_11102_));
 sg13g2_o21ai_1 _17530_ (.B1(_11114_),
    .Y(_00415_),
    .A1(net265),
    .A2(_11113_));
 sg13g2_nand2_1 _17531_ (.Y(_11115_),
    .A(net751),
    .B(\mem.mem_internal.code_mem[133][6] ));
 sg13g2_nand2_1 _17532_ (.Y(_11116_),
    .A(net1160),
    .B(_11102_));
 sg13g2_o21ai_1 _17533_ (.B1(_11116_),
    .Y(_00416_),
    .A1(_11103_),
    .A2(_11115_));
 sg13g2_buf_1 _17534_ (.A(_11031_),
    .X(_11117_));
 sg13g2_nand2_1 _17535_ (.Y(_11118_),
    .A(net750),
    .B(\mem.mem_internal.code_mem[133][7] ));
 sg13g2_nand2_1 _17536_ (.Y(_11119_),
    .A(net1159),
    .B(_11102_));
 sg13g2_o21ai_1 _17537_ (.B1(_11119_),
    .Y(_00417_),
    .A1(_11103_),
    .A2(_11118_));
 sg13g2_nand2_1 _17538_ (.Y(_11120_),
    .A(_11059_),
    .B(\mem.mem_internal.code_mem[134][0] ));
 sg13g2_nor2_1 _17539_ (.A(_10350_),
    .B(net467),
    .Y(_11121_));
 sg13g2_buf_2 _17540_ (.A(_11121_),
    .X(_11122_));
 sg13g2_buf_1 _17541_ (.A(_11122_),
    .X(_11123_));
 sg13g2_nand2_1 _17542_ (.Y(_11124_),
    .A(net1166),
    .B(net264));
 sg13g2_o21ai_1 _17543_ (.B1(_11124_),
    .Y(_00418_),
    .A1(_11120_),
    .A2(net264));
 sg13g2_nand2_1 _17544_ (.Y(_11125_),
    .A(net750),
    .B(\mem.mem_internal.code_mem[134][1] ));
 sg13g2_nand2_1 _17545_ (.Y(_11126_),
    .A(net1165),
    .B(net264));
 sg13g2_o21ai_1 _17546_ (.B1(_11126_),
    .Y(_00419_),
    .A1(net264),
    .A2(_11125_));
 sg13g2_nand2_1 _17547_ (.Y(_11127_),
    .A(net750),
    .B(\mem.mem_internal.code_mem[134][2] ));
 sg13g2_nand2_1 _17548_ (.Y(_11128_),
    .A(net1164),
    .B(_11122_));
 sg13g2_o21ai_1 _17549_ (.B1(_11128_),
    .Y(_00420_),
    .A1(net264),
    .A2(_11127_));
 sg13g2_nand2_1 _17550_ (.Y(_11129_),
    .A(_11117_),
    .B(\mem.mem_internal.code_mem[134][3] ));
 sg13g2_nand2_1 _17551_ (.Y(_11130_),
    .A(net1163),
    .B(_11122_));
 sg13g2_o21ai_1 _17552_ (.B1(_11130_),
    .Y(_00421_),
    .A1(net264),
    .A2(_11129_));
 sg13g2_nand2_1 _17553_ (.Y(_11131_),
    .A(net750),
    .B(\mem.mem_internal.code_mem[134][4] ));
 sg13g2_nand2_1 _17554_ (.Y(_11132_),
    .A(net1162),
    .B(_11122_));
 sg13g2_o21ai_1 _17555_ (.B1(_11132_),
    .Y(_00422_),
    .A1(net264),
    .A2(_11131_));
 sg13g2_nand2_1 _17556_ (.Y(_11133_),
    .A(net750),
    .B(\mem.mem_internal.code_mem[134][5] ));
 sg13g2_nand2_1 _17557_ (.Y(_11134_),
    .A(net1161),
    .B(_11122_));
 sg13g2_o21ai_1 _17558_ (.B1(_11134_),
    .Y(_00423_),
    .A1(_11123_),
    .A2(_11133_));
 sg13g2_nand2_1 _17559_ (.Y(_11135_),
    .A(_11117_),
    .B(\mem.mem_internal.code_mem[134][6] ));
 sg13g2_nand2_1 _17560_ (.Y(_11136_),
    .A(net1160),
    .B(_11122_));
 sg13g2_o21ai_1 _17561_ (.B1(_11136_),
    .Y(_00424_),
    .A1(_11123_),
    .A2(_11135_));
 sg13g2_nand2_1 _17562_ (.Y(_11137_),
    .A(net750),
    .B(\mem.mem_internal.code_mem[134][7] ));
 sg13g2_nand2_1 _17563_ (.Y(_11138_),
    .A(net1159),
    .B(_11122_));
 sg13g2_o21ai_1 _17564_ (.B1(_11138_),
    .Y(_00425_),
    .A1(net264),
    .A2(_11137_));
 sg13g2_nand2_1 _17565_ (.Y(_11139_),
    .A(_11059_),
    .B(\mem.mem_internal.code_mem[135][0] ));
 sg13g2_nor2_1 _17566_ (.A(_10373_),
    .B(_10979_),
    .Y(_11140_));
 sg13g2_buf_2 _17567_ (.A(_11140_),
    .X(_11141_));
 sg13g2_buf_1 _17568_ (.A(_11141_),
    .X(_11142_));
 sg13g2_nand2_1 _17569_ (.Y(_11143_),
    .A(net1166),
    .B(net263));
 sg13g2_o21ai_1 _17570_ (.B1(_11143_),
    .Y(_00426_),
    .A1(_11139_),
    .A2(net263));
 sg13g2_nand2_1 _17571_ (.Y(_11144_),
    .A(net750),
    .B(\mem.mem_internal.code_mem[135][1] ));
 sg13g2_nand2_1 _17572_ (.Y(_11145_),
    .A(net1165),
    .B(net263));
 sg13g2_o21ai_1 _17573_ (.B1(_11145_),
    .Y(_00427_),
    .A1(net263),
    .A2(_11144_));
 sg13g2_nand2_1 _17574_ (.Y(_11146_),
    .A(net750),
    .B(\mem.mem_internal.code_mem[135][2] ));
 sg13g2_nand2_1 _17575_ (.Y(_11147_),
    .A(net1164),
    .B(_11141_));
 sg13g2_o21ai_1 _17576_ (.B1(_11147_),
    .Y(_00428_),
    .A1(net263),
    .A2(_11146_));
 sg13g2_buf_1 _17577_ (.A(_11031_),
    .X(_11148_));
 sg13g2_nand2_1 _17578_ (.Y(_11149_),
    .A(net749),
    .B(\mem.mem_internal.code_mem[135][3] ));
 sg13g2_nand2_1 _17579_ (.Y(_11150_),
    .A(net1163),
    .B(_11141_));
 sg13g2_o21ai_1 _17580_ (.B1(_11150_),
    .Y(_00429_),
    .A1(net263),
    .A2(_11149_));
 sg13g2_nand2_1 _17581_ (.Y(_11151_),
    .A(net749),
    .B(\mem.mem_internal.code_mem[135][4] ));
 sg13g2_nand2_1 _17582_ (.Y(_11152_),
    .A(net1162),
    .B(_11141_));
 sg13g2_o21ai_1 _17583_ (.B1(_11152_),
    .Y(_00430_),
    .A1(net263),
    .A2(_11151_));
 sg13g2_nand2_1 _17584_ (.Y(_11153_),
    .A(net749),
    .B(\mem.mem_internal.code_mem[135][5] ));
 sg13g2_nand2_1 _17585_ (.Y(_11154_),
    .A(net1161),
    .B(_11141_));
 sg13g2_o21ai_1 _17586_ (.B1(_11154_),
    .Y(_00431_),
    .A1(_11142_),
    .A2(_11153_));
 sg13g2_nand2_1 _17587_ (.Y(_11155_),
    .A(_11148_),
    .B(\mem.mem_internal.code_mem[135][6] ));
 sg13g2_nand2_1 _17588_ (.Y(_11156_),
    .A(net1160),
    .B(_11141_));
 sg13g2_o21ai_1 _17589_ (.B1(_11156_),
    .Y(_00432_),
    .A1(_11142_),
    .A2(_11155_));
 sg13g2_nand2_1 _17590_ (.Y(_11157_),
    .A(_11148_),
    .B(\mem.mem_internal.code_mem[135][7] ));
 sg13g2_nand2_1 _17591_ (.Y(_11158_),
    .A(net1159),
    .B(_11141_));
 sg13g2_o21ai_1 _17592_ (.B1(_11158_),
    .Y(_00433_),
    .A1(net263),
    .A2(_11157_));
 sg13g2_nand2_1 _17593_ (.Y(_11159_),
    .A(net849),
    .B(\mem.mem_internal.code_mem[136][0] ));
 sg13g2_nor2_1 _17594_ (.A(net552),
    .B(net467),
    .Y(_11160_));
 sg13g2_buf_2 _17595_ (.A(_11160_),
    .X(_11161_));
 sg13g2_buf_1 _17596_ (.A(_11161_),
    .X(_11162_));
 sg13g2_buf_2 _17597_ (.A(_10251_),
    .X(_11163_));
 sg13g2_buf_1 _17598_ (.A(_11163_),
    .X(_11164_));
 sg13g2_nand2_1 _17599_ (.Y(_11165_),
    .A(_11164_),
    .B(net262));
 sg13g2_o21ai_1 _17600_ (.B1(_11165_),
    .Y(_00434_),
    .A1(_11159_),
    .A2(net262));
 sg13g2_nand2_1 _17601_ (.Y(_11166_),
    .A(net749),
    .B(\mem.mem_internal.code_mem[136][1] ));
 sg13g2_buf_1 _17602_ (.A(_10256_),
    .X(_11167_));
 sg13g2_buf_1 _17603_ (.A(_11167_),
    .X(_11168_));
 sg13g2_nand2_1 _17604_ (.Y(_11169_),
    .A(net1157),
    .B(net262));
 sg13g2_o21ai_1 _17605_ (.B1(_11169_),
    .Y(_00435_),
    .A1(net262),
    .A2(_11166_));
 sg13g2_nand2_1 _17606_ (.Y(_11170_),
    .A(net749),
    .B(\mem.mem_internal.code_mem[136][2] ));
 sg13g2_buf_2 _17607_ (.A(_10262_),
    .X(_11171_));
 sg13g2_buf_1 _17608_ (.A(_11171_),
    .X(_11172_));
 sg13g2_nand2_1 _17609_ (.Y(_11173_),
    .A(_11172_),
    .B(_11161_));
 sg13g2_o21ai_1 _17610_ (.B1(_11173_),
    .Y(_00436_),
    .A1(_11162_),
    .A2(_11170_));
 sg13g2_nand2_1 _17611_ (.Y(_11174_),
    .A(net749),
    .B(\mem.mem_internal.code_mem[136][3] ));
 sg13g2_buf_2 _17612_ (.A(_10267_),
    .X(_11175_));
 sg13g2_buf_1 _17613_ (.A(_11175_),
    .X(_11176_));
 sg13g2_nand2_1 _17614_ (.Y(_11177_),
    .A(net1155),
    .B(_11161_));
 sg13g2_o21ai_1 _17615_ (.B1(_11177_),
    .Y(_00437_),
    .A1(_11162_),
    .A2(_11174_));
 sg13g2_nand2_1 _17616_ (.Y(_11178_),
    .A(net749),
    .B(\mem.mem_internal.code_mem[136][4] ));
 sg13g2_buf_2 _17617_ (.A(_10272_),
    .X(_11179_));
 sg13g2_buf_1 _17618_ (.A(_11179_),
    .X(_11180_));
 sg13g2_nand2_1 _17619_ (.Y(_11181_),
    .A(net1154),
    .B(_11161_));
 sg13g2_o21ai_1 _17620_ (.B1(_11181_),
    .Y(_00438_),
    .A1(net262),
    .A2(_11178_));
 sg13g2_nand2_1 _17621_ (.Y(_11182_),
    .A(net749),
    .B(\mem.mem_internal.code_mem[136][5] ));
 sg13g2_buf_2 _17622_ (.A(_10277_),
    .X(_11183_));
 sg13g2_buf_1 _17623_ (.A(_11183_),
    .X(_11184_));
 sg13g2_nand2_1 _17624_ (.Y(_11185_),
    .A(_11184_),
    .B(_11161_));
 sg13g2_o21ai_1 _17625_ (.B1(_11185_),
    .Y(_00439_),
    .A1(net262),
    .A2(_11182_));
 sg13g2_buf_1 _17626_ (.A(_11031_),
    .X(_11186_));
 sg13g2_nand2_1 _17627_ (.Y(_11187_),
    .A(net748),
    .B(\mem.mem_internal.code_mem[136][6] ));
 sg13g2_buf_2 _17628_ (.A(_10282_),
    .X(_11188_));
 sg13g2_buf_1 _17629_ (.A(_11188_),
    .X(_11189_));
 sg13g2_nand2_1 _17630_ (.Y(_11190_),
    .A(net1152),
    .B(_11161_));
 sg13g2_o21ai_1 _17631_ (.B1(_11190_),
    .Y(_00440_),
    .A1(net262),
    .A2(_11187_));
 sg13g2_nand2_1 _17632_ (.Y(_11191_),
    .A(net748),
    .B(\mem.mem_internal.code_mem[136][7] ));
 sg13g2_buf_2 _17633_ (.A(_10287_),
    .X(_11192_));
 sg13g2_buf_1 _17634_ (.A(_11192_),
    .X(_11193_));
 sg13g2_nand2_1 _17635_ (.Y(_11194_),
    .A(net1151),
    .B(_11161_));
 sg13g2_o21ai_1 _17636_ (.B1(_11194_),
    .Y(_00441_),
    .A1(net262),
    .A2(_11191_));
 sg13g2_nand2_1 _17637_ (.Y(_11195_),
    .A(net849),
    .B(\mem.mem_internal.code_mem[137][0] ));
 sg13g2_nor2_1 _17638_ (.A(net551),
    .B(net467),
    .Y(_11196_));
 sg13g2_buf_2 _17639_ (.A(_11196_),
    .X(_11197_));
 sg13g2_buf_1 _17640_ (.A(_11197_),
    .X(_11198_));
 sg13g2_nand2_1 _17641_ (.Y(_11199_),
    .A(net1158),
    .B(net261));
 sg13g2_o21ai_1 _17642_ (.B1(_11199_),
    .Y(_00442_),
    .A1(_11195_),
    .A2(net261));
 sg13g2_nand2_1 _17643_ (.Y(_11200_),
    .A(net748),
    .B(\mem.mem_internal.code_mem[137][1] ));
 sg13g2_nand2_1 _17644_ (.Y(_11201_),
    .A(net1157),
    .B(net261));
 sg13g2_o21ai_1 _17645_ (.B1(_11201_),
    .Y(_00443_),
    .A1(net261),
    .A2(_11200_));
 sg13g2_nand2_1 _17646_ (.Y(_11202_),
    .A(net748),
    .B(\mem.mem_internal.code_mem[137][2] ));
 sg13g2_nand2_1 _17647_ (.Y(_11203_),
    .A(net1156),
    .B(_11197_));
 sg13g2_o21ai_1 _17648_ (.B1(_11203_),
    .Y(_00444_),
    .A1(_11198_),
    .A2(_11202_));
 sg13g2_nand2_1 _17649_ (.Y(_11204_),
    .A(net748),
    .B(\mem.mem_internal.code_mem[137][3] ));
 sg13g2_nand2_1 _17650_ (.Y(_11205_),
    .A(net1155),
    .B(_11197_));
 sg13g2_o21ai_1 _17651_ (.B1(_11205_),
    .Y(_00445_),
    .A1(_11198_),
    .A2(_11204_));
 sg13g2_nand2_1 _17652_ (.Y(_11206_),
    .A(net748),
    .B(\mem.mem_internal.code_mem[137][4] ));
 sg13g2_nand2_1 _17653_ (.Y(_11207_),
    .A(net1154),
    .B(_11197_));
 sg13g2_o21ai_1 _17654_ (.B1(_11207_),
    .Y(_00446_),
    .A1(net261),
    .A2(_11206_));
 sg13g2_nand2_1 _17655_ (.Y(_11208_),
    .A(_11186_),
    .B(\mem.mem_internal.code_mem[137][5] ));
 sg13g2_nand2_1 _17656_ (.Y(_11209_),
    .A(_11184_),
    .B(_11197_));
 sg13g2_o21ai_1 _17657_ (.B1(_11209_),
    .Y(_00447_),
    .A1(net261),
    .A2(_11208_));
 sg13g2_nand2_1 _17658_ (.Y(_11210_),
    .A(_11186_),
    .B(\mem.mem_internal.code_mem[137][6] ));
 sg13g2_nand2_1 _17659_ (.Y(_11211_),
    .A(net1152),
    .B(_11197_));
 sg13g2_o21ai_1 _17660_ (.B1(_11211_),
    .Y(_00448_),
    .A1(net261),
    .A2(_11210_));
 sg13g2_nand2_1 _17661_ (.Y(_11212_),
    .A(net748),
    .B(\mem.mem_internal.code_mem[137][7] ));
 sg13g2_nand2_1 _17662_ (.Y(_11213_),
    .A(net1151),
    .B(_11197_));
 sg13g2_o21ai_1 _17663_ (.B1(_11213_),
    .Y(_00449_),
    .A1(net261),
    .A2(_11212_));
 sg13g2_nand2_1 _17664_ (.Y(_11214_),
    .A(net849),
    .B(\mem.mem_internal.code_mem[138][0] ));
 sg13g2_nor2_1 _17665_ (.A(net550),
    .B(_10978_),
    .Y(_11215_));
 sg13g2_buf_2 _17666_ (.A(_11215_),
    .X(_11216_));
 sg13g2_buf_1 _17667_ (.A(_11216_),
    .X(_11217_));
 sg13g2_nand2_1 _17668_ (.Y(_11218_),
    .A(net1158),
    .B(_11217_));
 sg13g2_o21ai_1 _17669_ (.B1(_11218_),
    .Y(_00450_),
    .A1(_11214_),
    .A2(_11217_));
 sg13g2_nand2_1 _17670_ (.Y(_11219_),
    .A(net748),
    .B(\mem.mem_internal.code_mem[138][1] ));
 sg13g2_nand2_1 _17671_ (.Y(_11220_),
    .A(net1157),
    .B(net390));
 sg13g2_o21ai_1 _17672_ (.B1(_11220_),
    .Y(_00451_),
    .A1(net390),
    .A2(_11219_));
 sg13g2_buf_1 _17673_ (.A(_11031_),
    .X(_11221_));
 sg13g2_nand2_1 _17674_ (.Y(_11222_),
    .A(net747),
    .B(\mem.mem_internal.code_mem[138][2] ));
 sg13g2_nand2_1 _17675_ (.Y(_11223_),
    .A(net1156),
    .B(_11216_));
 sg13g2_o21ai_1 _17676_ (.B1(_11223_),
    .Y(_00452_),
    .A1(net390),
    .A2(_11222_));
 sg13g2_nand2_1 _17677_ (.Y(_11224_),
    .A(net747),
    .B(\mem.mem_internal.code_mem[138][3] ));
 sg13g2_nand2_1 _17678_ (.Y(_11225_),
    .A(net1155),
    .B(_11216_));
 sg13g2_o21ai_1 _17679_ (.B1(_11225_),
    .Y(_00453_),
    .A1(net390),
    .A2(_11224_));
 sg13g2_nand2_1 _17680_ (.Y(_11226_),
    .A(net747),
    .B(\mem.mem_internal.code_mem[138][4] ));
 sg13g2_nand2_1 _17681_ (.Y(_11227_),
    .A(_11180_),
    .B(_11216_));
 sg13g2_o21ai_1 _17682_ (.B1(_11227_),
    .Y(_00454_),
    .A1(net390),
    .A2(_11226_));
 sg13g2_nand2_1 _17683_ (.Y(_11228_),
    .A(_11221_),
    .B(\mem.mem_internal.code_mem[138][5] ));
 sg13g2_nand2_1 _17684_ (.Y(_11229_),
    .A(net1153),
    .B(_11216_));
 sg13g2_o21ai_1 _17685_ (.B1(_11229_),
    .Y(_00455_),
    .A1(net390),
    .A2(_11228_));
 sg13g2_nand2_1 _17686_ (.Y(_11230_),
    .A(net747),
    .B(\mem.mem_internal.code_mem[138][6] ));
 sg13g2_nand2_1 _17687_ (.Y(_11231_),
    .A(net1152),
    .B(_11216_));
 sg13g2_o21ai_1 _17688_ (.B1(_11231_),
    .Y(_00456_),
    .A1(net390),
    .A2(_11230_));
 sg13g2_nand2_1 _17689_ (.Y(_11232_),
    .A(net747),
    .B(\mem.mem_internal.code_mem[138][7] ));
 sg13g2_nand2_1 _17690_ (.Y(_11233_),
    .A(net1151),
    .B(_11216_));
 sg13g2_o21ai_1 _17691_ (.B1(_11233_),
    .Y(_00457_),
    .A1(net390),
    .A2(_11232_));
 sg13g2_nand2_1 _17692_ (.Y(_11234_),
    .A(net849),
    .B(\mem.mem_internal.code_mem[139][0] ));
 sg13g2_nor2_1 _17693_ (.A(net549),
    .B(_10978_),
    .Y(_11235_));
 sg13g2_buf_2 _17694_ (.A(_11235_),
    .X(_11236_));
 sg13g2_buf_1 _17695_ (.A(_11236_),
    .X(_11237_));
 sg13g2_nand2_1 _17696_ (.Y(_11238_),
    .A(_11164_),
    .B(net389));
 sg13g2_o21ai_1 _17697_ (.B1(_11238_),
    .Y(_00458_),
    .A1(_11234_),
    .A2(net389));
 sg13g2_nand2_1 _17698_ (.Y(_11239_),
    .A(net747),
    .B(\mem.mem_internal.code_mem[139][1] ));
 sg13g2_nand2_1 _17699_ (.Y(_11240_),
    .A(net1157),
    .B(net389));
 sg13g2_o21ai_1 _17700_ (.B1(_11240_),
    .Y(_00459_),
    .A1(net389),
    .A2(_11239_));
 sg13g2_nand2_1 _17701_ (.Y(_11241_),
    .A(net747),
    .B(\mem.mem_internal.code_mem[139][2] ));
 sg13g2_nand2_1 _17702_ (.Y(_11242_),
    .A(_11172_),
    .B(_11236_));
 sg13g2_o21ai_1 _17703_ (.B1(_11242_),
    .Y(_00460_),
    .A1(net389),
    .A2(_11241_));
 sg13g2_nand2_1 _17704_ (.Y(_11243_),
    .A(net747),
    .B(\mem.mem_internal.code_mem[139][3] ));
 sg13g2_nand2_1 _17705_ (.Y(_11244_),
    .A(net1155),
    .B(_11236_));
 sg13g2_o21ai_1 _17706_ (.B1(_11244_),
    .Y(_00461_),
    .A1(net389),
    .A2(_11243_));
 sg13g2_nand2_1 _17707_ (.Y(_11245_),
    .A(_11221_),
    .B(\mem.mem_internal.code_mem[139][4] ));
 sg13g2_nand2_1 _17708_ (.Y(_11246_),
    .A(_11180_),
    .B(_11236_));
 sg13g2_o21ai_1 _17709_ (.B1(_11246_),
    .Y(_00462_),
    .A1(_11237_),
    .A2(_11245_));
 sg13g2_buf_1 _17710_ (.A(_10415_),
    .X(_11247_));
 sg13g2_buf_1 _17711_ (.A(_11247_),
    .X(_11248_));
 sg13g2_nand2_1 _17712_ (.Y(_11249_),
    .A(_11248_),
    .B(\mem.mem_internal.code_mem[139][5] ));
 sg13g2_nand2_1 _17713_ (.Y(_11250_),
    .A(net1153),
    .B(_11236_));
 sg13g2_o21ai_1 _17714_ (.B1(_11250_),
    .Y(_00463_),
    .A1(net389),
    .A2(_11249_));
 sg13g2_nand2_1 _17715_ (.Y(_11251_),
    .A(_11248_),
    .B(\mem.mem_internal.code_mem[139][6] ));
 sg13g2_nand2_1 _17716_ (.Y(_11252_),
    .A(_11189_),
    .B(_11236_));
 sg13g2_o21ai_1 _17717_ (.B1(_11252_),
    .Y(_00464_),
    .A1(_11237_),
    .A2(_11251_));
 sg13g2_nand2_1 _17718_ (.Y(_11253_),
    .A(net746),
    .B(\mem.mem_internal.code_mem[139][7] ));
 sg13g2_nand2_1 _17719_ (.Y(_11254_),
    .A(net1151),
    .B(_11236_));
 sg13g2_o21ai_1 _17720_ (.B1(_11254_),
    .Y(_00465_),
    .A1(net389),
    .A2(_11253_));
 sg13g2_nand2_1 _17721_ (.Y(_11255_),
    .A(net849),
    .B(\mem.mem_internal.code_mem[13][0] ));
 sg13g2_nor2_1 _17722_ (.A(net470),
    .B(net548),
    .Y(_11256_));
 sg13g2_buf_2 _17723_ (.A(_11256_),
    .X(_11257_));
 sg13g2_buf_1 _17724_ (.A(_11257_),
    .X(_11258_));
 sg13g2_nand2_1 _17725_ (.Y(_11259_),
    .A(net1158),
    .B(net260));
 sg13g2_o21ai_1 _17726_ (.B1(_11259_),
    .Y(_00466_),
    .A1(_11255_),
    .A2(net260));
 sg13g2_nand2_1 _17727_ (.Y(_11260_),
    .A(net746),
    .B(\mem.mem_internal.code_mem[13][1] ));
 sg13g2_nand2_1 _17728_ (.Y(_11261_),
    .A(_11168_),
    .B(_11258_));
 sg13g2_o21ai_1 _17729_ (.B1(_11261_),
    .Y(_00467_),
    .A1(net260),
    .A2(_11260_));
 sg13g2_nand2_1 _17730_ (.Y(_11262_),
    .A(net746),
    .B(\mem.mem_internal.code_mem[13][2] ));
 sg13g2_nand2_1 _17731_ (.Y(_11263_),
    .A(net1156),
    .B(_11257_));
 sg13g2_o21ai_1 _17732_ (.B1(_11263_),
    .Y(_00468_),
    .A1(net260),
    .A2(_11262_));
 sg13g2_nand2_1 _17733_ (.Y(_11264_),
    .A(net746),
    .B(\mem.mem_internal.code_mem[13][3] ));
 sg13g2_nand2_1 _17734_ (.Y(_11265_),
    .A(_11176_),
    .B(_11257_));
 sg13g2_o21ai_1 _17735_ (.B1(_11265_),
    .Y(_00469_),
    .A1(net260),
    .A2(_11264_));
 sg13g2_nand2_1 _17736_ (.Y(_11266_),
    .A(net746),
    .B(\mem.mem_internal.code_mem[13][4] ));
 sg13g2_nand2_1 _17737_ (.Y(_11267_),
    .A(net1154),
    .B(_11257_));
 sg13g2_o21ai_1 _17738_ (.B1(_11267_),
    .Y(_00470_),
    .A1(_11258_),
    .A2(_11266_));
 sg13g2_nand2_1 _17739_ (.Y(_11268_),
    .A(net746),
    .B(\mem.mem_internal.code_mem[13][5] ));
 sg13g2_nand2_1 _17740_ (.Y(_11269_),
    .A(net1153),
    .B(_11257_));
 sg13g2_o21ai_1 _17741_ (.B1(_11269_),
    .Y(_00471_),
    .A1(net260),
    .A2(_11268_));
 sg13g2_nand2_1 _17742_ (.Y(_11270_),
    .A(net746),
    .B(\mem.mem_internal.code_mem[13][6] ));
 sg13g2_nand2_1 _17743_ (.Y(_11271_),
    .A(_11189_),
    .B(_11257_));
 sg13g2_o21ai_1 _17744_ (.B1(_11271_),
    .Y(_00472_),
    .A1(net260),
    .A2(_11270_));
 sg13g2_nand2_1 _17745_ (.Y(_11272_),
    .A(net746),
    .B(\mem.mem_internal.code_mem[13][7] ));
 sg13g2_nand2_1 _17746_ (.Y(_11273_),
    .A(_11193_),
    .B(_11257_));
 sg13g2_o21ai_1 _17747_ (.B1(_11273_),
    .Y(_00473_),
    .A1(net260),
    .A2(_11272_));
 sg13g2_buf_1 _17748_ (.A(_11058_),
    .X(_11274_));
 sg13g2_nand2_1 _17749_ (.Y(_11275_),
    .A(net848),
    .B(\mem.mem_internal.code_mem[140][0] ));
 sg13g2_nor2_1 _17750_ (.A(net773),
    .B(_10978_),
    .Y(_11276_));
 sg13g2_buf_2 _17751_ (.A(_11276_),
    .X(_11277_));
 sg13g2_buf_1 _17752_ (.A(_11277_),
    .X(_11278_));
 sg13g2_nand2_1 _17753_ (.Y(_11279_),
    .A(net1158),
    .B(net388));
 sg13g2_o21ai_1 _17754_ (.B1(_11279_),
    .Y(_00474_),
    .A1(_11275_),
    .A2(_11278_));
 sg13g2_buf_1 _17755_ (.A(_11247_),
    .X(_11280_));
 sg13g2_nand2_1 _17756_ (.Y(_11281_),
    .A(net745),
    .B(\mem.mem_internal.code_mem[140][1] ));
 sg13g2_nand2_1 _17757_ (.Y(_11282_),
    .A(net1157),
    .B(net388));
 sg13g2_o21ai_1 _17758_ (.B1(_11282_),
    .Y(_00475_),
    .A1(net388),
    .A2(_11281_));
 sg13g2_nand2_1 _17759_ (.Y(_11283_),
    .A(net745),
    .B(\mem.mem_internal.code_mem[140][2] ));
 sg13g2_nand2_1 _17760_ (.Y(_11284_),
    .A(net1156),
    .B(_11277_));
 sg13g2_o21ai_1 _17761_ (.B1(_11284_),
    .Y(_00476_),
    .A1(net388),
    .A2(_11283_));
 sg13g2_nand2_1 _17762_ (.Y(_11285_),
    .A(net745),
    .B(\mem.mem_internal.code_mem[140][3] ));
 sg13g2_nand2_1 _17763_ (.Y(_11286_),
    .A(net1155),
    .B(_11277_));
 sg13g2_o21ai_1 _17764_ (.B1(_11286_),
    .Y(_00477_),
    .A1(net388),
    .A2(_11285_));
 sg13g2_nand2_1 _17765_ (.Y(_11287_),
    .A(_11280_),
    .B(\mem.mem_internal.code_mem[140][4] ));
 sg13g2_nand2_1 _17766_ (.Y(_11288_),
    .A(net1154),
    .B(_11277_));
 sg13g2_o21ai_1 _17767_ (.B1(_11288_),
    .Y(_00478_),
    .A1(net388),
    .A2(_11287_));
 sg13g2_nand2_1 _17768_ (.Y(_11289_),
    .A(_11280_),
    .B(\mem.mem_internal.code_mem[140][5] ));
 sg13g2_nand2_1 _17769_ (.Y(_11290_),
    .A(net1153),
    .B(_11277_));
 sg13g2_o21ai_1 _17770_ (.B1(_11290_),
    .Y(_00479_),
    .A1(_11278_),
    .A2(_11289_));
 sg13g2_nand2_1 _17771_ (.Y(_11291_),
    .A(net745),
    .B(\mem.mem_internal.code_mem[140][6] ));
 sg13g2_nand2_1 _17772_ (.Y(_11292_),
    .A(net1152),
    .B(_11277_));
 sg13g2_o21ai_1 _17773_ (.B1(_11292_),
    .Y(_00480_),
    .A1(net388),
    .A2(_11291_));
 sg13g2_nand2_1 _17774_ (.Y(_11293_),
    .A(net745),
    .B(\mem.mem_internal.code_mem[140][7] ));
 sg13g2_nand2_1 _17775_ (.Y(_11294_),
    .A(net1151),
    .B(_11277_));
 sg13g2_o21ai_1 _17776_ (.B1(_11294_),
    .Y(_00481_),
    .A1(net388),
    .A2(_11293_));
 sg13g2_nand2_1 _17777_ (.Y(_11295_),
    .A(net848),
    .B(\mem.mem_internal.code_mem[141][0] ));
 sg13g2_nor2_1 _17778_ (.A(net548),
    .B(_10978_),
    .Y(_11296_));
 sg13g2_buf_2 _17779_ (.A(_11296_),
    .X(_11297_));
 sg13g2_buf_1 _17780_ (.A(_11297_),
    .X(_11298_));
 sg13g2_nand2_1 _17781_ (.Y(_11299_),
    .A(net1158),
    .B(_11298_));
 sg13g2_o21ai_1 _17782_ (.B1(_11299_),
    .Y(_00482_),
    .A1(_11295_),
    .A2(net387));
 sg13g2_nand2_1 _17783_ (.Y(_11300_),
    .A(net745),
    .B(\mem.mem_internal.code_mem[141][1] ));
 sg13g2_nand2_1 _17784_ (.Y(_11301_),
    .A(net1157),
    .B(net387));
 sg13g2_o21ai_1 _17785_ (.B1(_11301_),
    .Y(_00483_),
    .A1(net387),
    .A2(_11300_));
 sg13g2_nand2_1 _17786_ (.Y(_11302_),
    .A(net745),
    .B(\mem.mem_internal.code_mem[141][2] ));
 sg13g2_nand2_1 _17787_ (.Y(_11303_),
    .A(net1156),
    .B(_11297_));
 sg13g2_o21ai_1 _17788_ (.B1(_11303_),
    .Y(_00484_),
    .A1(net387),
    .A2(_11302_));
 sg13g2_nand2_1 _17789_ (.Y(_11304_),
    .A(net745),
    .B(\mem.mem_internal.code_mem[141][3] ));
 sg13g2_nand2_1 _17790_ (.Y(_11305_),
    .A(net1155),
    .B(_11297_));
 sg13g2_o21ai_1 _17791_ (.B1(_11305_),
    .Y(_00485_),
    .A1(net387),
    .A2(_11304_));
 sg13g2_buf_1 _17792_ (.A(_11247_),
    .X(_11306_));
 sg13g2_nand2_1 _17793_ (.Y(_11307_),
    .A(net744),
    .B(\mem.mem_internal.code_mem[141][4] ));
 sg13g2_nand2_1 _17794_ (.Y(_11308_),
    .A(net1154),
    .B(_11297_));
 sg13g2_o21ai_1 _17795_ (.B1(_11308_),
    .Y(_00486_),
    .A1(net387),
    .A2(_11307_));
 sg13g2_nand2_1 _17796_ (.Y(_11309_),
    .A(net744),
    .B(\mem.mem_internal.code_mem[141][5] ));
 sg13g2_nand2_1 _17797_ (.Y(_11310_),
    .A(net1153),
    .B(_11297_));
 sg13g2_o21ai_1 _17798_ (.B1(_11310_),
    .Y(_00487_),
    .A1(_11298_),
    .A2(_11309_));
 sg13g2_nand2_1 _17799_ (.Y(_11311_),
    .A(net744),
    .B(\mem.mem_internal.code_mem[141][6] ));
 sg13g2_nand2_1 _17800_ (.Y(_11312_),
    .A(net1152),
    .B(_11297_));
 sg13g2_o21ai_1 _17801_ (.B1(_11312_),
    .Y(_00488_),
    .A1(net387),
    .A2(_11311_));
 sg13g2_nand2_1 _17802_ (.Y(_11313_),
    .A(net744),
    .B(\mem.mem_internal.code_mem[141][7] ));
 sg13g2_nand2_1 _17803_ (.Y(_11314_),
    .A(net1151),
    .B(_11297_));
 sg13g2_o21ai_1 _17804_ (.B1(_11314_),
    .Y(_00489_),
    .A1(net387),
    .A2(_11313_));
 sg13g2_nand2_1 _17805_ (.Y(_11315_),
    .A(net848),
    .B(\mem.mem_internal.code_mem[142][0] ));
 sg13g2_nor2_1 _17806_ (.A(net547),
    .B(_10978_),
    .Y(_11316_));
 sg13g2_buf_2 _17807_ (.A(_11316_),
    .X(_11317_));
 sg13g2_buf_1 _17808_ (.A(_11317_),
    .X(_11318_));
 sg13g2_nand2_1 _17809_ (.Y(_11319_),
    .A(net1158),
    .B(net386));
 sg13g2_o21ai_1 _17810_ (.B1(_11319_),
    .Y(_00490_),
    .A1(_11315_),
    .A2(_11318_));
 sg13g2_nand2_1 _17811_ (.Y(_11320_),
    .A(net744),
    .B(\mem.mem_internal.code_mem[142][1] ));
 sg13g2_nand2_1 _17812_ (.Y(_11321_),
    .A(net1157),
    .B(net386));
 sg13g2_o21ai_1 _17813_ (.B1(_11321_),
    .Y(_00491_),
    .A1(net386),
    .A2(_11320_));
 sg13g2_nand2_1 _17814_ (.Y(_11322_),
    .A(net744),
    .B(\mem.mem_internal.code_mem[142][2] ));
 sg13g2_nand2_1 _17815_ (.Y(_11323_),
    .A(net1156),
    .B(_11317_));
 sg13g2_o21ai_1 _17816_ (.B1(_11323_),
    .Y(_00492_),
    .A1(net386),
    .A2(_11322_));
 sg13g2_nand2_1 _17817_ (.Y(_11324_),
    .A(net744),
    .B(\mem.mem_internal.code_mem[142][3] ));
 sg13g2_nand2_1 _17818_ (.Y(_11325_),
    .A(net1155),
    .B(_11317_));
 sg13g2_o21ai_1 _17819_ (.B1(_11325_),
    .Y(_00493_),
    .A1(net386),
    .A2(_11324_));
 sg13g2_nand2_1 _17820_ (.Y(_11326_),
    .A(_11306_),
    .B(\mem.mem_internal.code_mem[142][4] ));
 sg13g2_nand2_1 _17821_ (.Y(_11327_),
    .A(net1154),
    .B(_11317_));
 sg13g2_o21ai_1 _17822_ (.B1(_11327_),
    .Y(_00494_),
    .A1(net386),
    .A2(_11326_));
 sg13g2_nand2_1 _17823_ (.Y(_11328_),
    .A(_11306_),
    .B(\mem.mem_internal.code_mem[142][5] ));
 sg13g2_nand2_1 _17824_ (.Y(_11329_),
    .A(net1153),
    .B(_11317_));
 sg13g2_o21ai_1 _17825_ (.B1(_11329_),
    .Y(_00495_),
    .A1(_11318_),
    .A2(_11328_));
 sg13g2_nand2_1 _17826_ (.Y(_11330_),
    .A(net744),
    .B(\mem.mem_internal.code_mem[142][6] ));
 sg13g2_nand2_1 _17827_ (.Y(_11331_),
    .A(net1152),
    .B(_11317_));
 sg13g2_o21ai_1 _17828_ (.B1(_11331_),
    .Y(_00496_),
    .A1(net386),
    .A2(_11330_));
 sg13g2_buf_1 _17829_ (.A(_11247_),
    .X(_11332_));
 sg13g2_nand2_1 _17830_ (.Y(_11333_),
    .A(net743),
    .B(\mem.mem_internal.code_mem[142][7] ));
 sg13g2_nand2_1 _17831_ (.Y(_11334_),
    .A(net1151),
    .B(_11317_));
 sg13g2_o21ai_1 _17832_ (.B1(_11334_),
    .Y(_00497_),
    .A1(net386),
    .A2(_11333_));
 sg13g2_nand2_1 _17833_ (.Y(_11335_),
    .A(net848),
    .B(\mem.mem_internal.code_mem[143][0] ));
 sg13g2_nor2_1 _17834_ (.A(net770),
    .B(_10978_),
    .Y(_11336_));
 sg13g2_buf_2 _17835_ (.A(_11336_),
    .X(_11337_));
 sg13g2_buf_1 _17836_ (.A(_11337_),
    .X(_11338_));
 sg13g2_nand2_1 _17837_ (.Y(_11339_),
    .A(net1158),
    .B(net385));
 sg13g2_o21ai_1 _17838_ (.B1(_11339_),
    .Y(_00498_),
    .A1(_11335_),
    .A2(_11338_));
 sg13g2_nand2_1 _17839_ (.Y(_11340_),
    .A(net743),
    .B(\mem.mem_internal.code_mem[143][1] ));
 sg13g2_nand2_1 _17840_ (.Y(_11341_),
    .A(net1157),
    .B(net385));
 sg13g2_o21ai_1 _17841_ (.B1(_11341_),
    .Y(_00499_),
    .A1(net385),
    .A2(_11340_));
 sg13g2_nand2_1 _17842_ (.Y(_11342_),
    .A(net743),
    .B(\mem.mem_internal.code_mem[143][2] ));
 sg13g2_nand2_1 _17843_ (.Y(_11343_),
    .A(net1156),
    .B(_11337_));
 sg13g2_o21ai_1 _17844_ (.B1(_11343_),
    .Y(_00500_),
    .A1(net385),
    .A2(_11342_));
 sg13g2_nand2_1 _17845_ (.Y(_11344_),
    .A(net743),
    .B(\mem.mem_internal.code_mem[143][3] ));
 sg13g2_nand2_1 _17846_ (.Y(_11345_),
    .A(net1155),
    .B(_11337_));
 sg13g2_o21ai_1 _17847_ (.B1(_11345_),
    .Y(_00501_),
    .A1(net385),
    .A2(_11344_));
 sg13g2_nand2_1 _17848_ (.Y(_11346_),
    .A(net743),
    .B(\mem.mem_internal.code_mem[143][4] ));
 sg13g2_nand2_1 _17849_ (.Y(_11347_),
    .A(net1154),
    .B(_11337_));
 sg13g2_o21ai_1 _17850_ (.B1(_11347_),
    .Y(_00502_),
    .A1(_11338_),
    .A2(_11346_));
 sg13g2_nand2_1 _17851_ (.Y(_11348_),
    .A(_11332_),
    .B(\mem.mem_internal.code_mem[143][5] ));
 sg13g2_nand2_1 _17852_ (.Y(_11349_),
    .A(net1153),
    .B(_11337_));
 sg13g2_o21ai_1 _17853_ (.B1(_11349_),
    .Y(_00503_),
    .A1(net385),
    .A2(_11348_));
 sg13g2_nand2_1 _17854_ (.Y(_11350_),
    .A(net743),
    .B(\mem.mem_internal.code_mem[143][6] ));
 sg13g2_nand2_1 _17855_ (.Y(_11351_),
    .A(net1152),
    .B(_11337_));
 sg13g2_o21ai_1 _17856_ (.B1(_11351_),
    .Y(_00504_),
    .A1(net385),
    .A2(_11350_));
 sg13g2_nand2_1 _17857_ (.Y(_11352_),
    .A(net743),
    .B(\mem.mem_internal.code_mem[143][7] ));
 sg13g2_nand2_1 _17858_ (.Y(_11353_),
    .A(net1151),
    .B(_11337_));
 sg13g2_o21ai_1 _17859_ (.B1(_11353_),
    .Y(_00505_),
    .A1(net385),
    .A2(_11352_));
 sg13g2_nand2_1 _17860_ (.Y(_11354_),
    .A(_11274_),
    .B(\mem.mem_internal.code_mem[144][0] ));
 sg13g2_nor3_2 _17861_ (.A(_10114_),
    .B(_10034_),
    .C(_10243_),
    .Y(_11355_));
 sg13g2_nand2_1 _17862_ (.Y(_11356_),
    .A(_10976_),
    .B(_11355_));
 sg13g2_buf_2 _17863_ (.A(_11356_),
    .X(_11357_));
 sg13g2_buf_1 _17864_ (.A(_11357_),
    .X(_11358_));
 sg13g2_nor2_1 _17865_ (.A(net529),
    .B(net466),
    .Y(_11359_));
 sg13g2_buf_2 _17866_ (.A(_11359_),
    .X(_11360_));
 sg13g2_buf_1 _17867_ (.A(_11360_),
    .X(_11361_));
 sg13g2_nand2_1 _17868_ (.Y(_11362_),
    .A(net1158),
    .B(net259));
 sg13g2_o21ai_1 _17869_ (.B1(_11362_),
    .Y(_00506_),
    .A1(_11354_),
    .A2(net259));
 sg13g2_nand2_1 _17870_ (.Y(_11363_),
    .A(_11332_),
    .B(\mem.mem_internal.code_mem[144][1] ));
 sg13g2_nand2_1 _17871_ (.Y(_11364_),
    .A(_11168_),
    .B(net259));
 sg13g2_o21ai_1 _17872_ (.B1(_11364_),
    .Y(_00507_),
    .A1(net259),
    .A2(_11363_));
 sg13g2_nand2_1 _17873_ (.Y(_11365_),
    .A(net743),
    .B(\mem.mem_internal.code_mem[144][2] ));
 sg13g2_nand2_1 _17874_ (.Y(_11366_),
    .A(net1156),
    .B(_11360_));
 sg13g2_o21ai_1 _17875_ (.B1(_11366_),
    .Y(_00508_),
    .A1(net259),
    .A2(_11365_));
 sg13g2_buf_1 _17876_ (.A(_11247_),
    .X(_11367_));
 sg13g2_nand2_1 _17877_ (.Y(_11368_),
    .A(net742),
    .B(\mem.mem_internal.code_mem[144][3] ));
 sg13g2_nand2_1 _17878_ (.Y(_11369_),
    .A(_11176_),
    .B(_11360_));
 sg13g2_o21ai_1 _17879_ (.B1(_11369_),
    .Y(_00509_),
    .A1(net259),
    .A2(_11368_));
 sg13g2_nand2_1 _17880_ (.Y(_11370_),
    .A(net742),
    .B(\mem.mem_internal.code_mem[144][4] ));
 sg13g2_nand2_1 _17881_ (.Y(_11371_),
    .A(net1154),
    .B(_11360_));
 sg13g2_o21ai_1 _17882_ (.B1(_11371_),
    .Y(_00510_),
    .A1(net259),
    .A2(_11370_));
 sg13g2_nand2_1 _17883_ (.Y(_11372_),
    .A(net742),
    .B(\mem.mem_internal.code_mem[144][5] ));
 sg13g2_nand2_1 _17884_ (.Y(_11373_),
    .A(net1153),
    .B(_11360_));
 sg13g2_o21ai_1 _17885_ (.B1(_11373_),
    .Y(_00511_),
    .A1(net259),
    .A2(_11372_));
 sg13g2_nand2_1 _17886_ (.Y(_11374_),
    .A(net742),
    .B(\mem.mem_internal.code_mem[144][6] ));
 sg13g2_nand2_1 _17887_ (.Y(_11375_),
    .A(net1152),
    .B(_11360_));
 sg13g2_o21ai_1 _17888_ (.B1(_11375_),
    .Y(_00512_),
    .A1(_11361_),
    .A2(_11374_));
 sg13g2_nand2_1 _17889_ (.Y(_11376_),
    .A(net742),
    .B(\mem.mem_internal.code_mem[144][7] ));
 sg13g2_nand2_1 _17890_ (.Y(_11377_),
    .A(_11193_),
    .B(_11360_));
 sg13g2_o21ai_1 _17891_ (.B1(_11377_),
    .Y(_00513_),
    .A1(_11361_),
    .A2(_11376_));
 sg13g2_nand2_1 _17892_ (.Y(_11378_),
    .A(_11274_),
    .B(\mem.mem_internal.code_mem[145][0] ));
 sg13g2_nor2_1 _17893_ (.A(net528),
    .B(_11358_),
    .Y(_11379_));
 sg13g2_buf_2 _17894_ (.A(_11379_),
    .X(_11380_));
 sg13g2_buf_1 _17895_ (.A(_11380_),
    .X(_11381_));
 sg13g2_buf_1 _17896_ (.A(_11163_),
    .X(_11382_));
 sg13g2_nand2_1 _17897_ (.Y(_11383_),
    .A(_11382_),
    .B(net258));
 sg13g2_o21ai_1 _17898_ (.B1(_11383_),
    .Y(_00514_),
    .A1(_11378_),
    .A2(net258));
 sg13g2_nand2_1 _17899_ (.Y(_11384_),
    .A(net742),
    .B(\mem.mem_internal.code_mem[145][1] ));
 sg13g2_buf_1 _17900_ (.A(_11167_),
    .X(_11385_));
 sg13g2_nand2_1 _17901_ (.Y(_11386_),
    .A(net1149),
    .B(net258));
 sg13g2_o21ai_1 _17902_ (.B1(_11386_),
    .Y(_00515_),
    .A1(net258),
    .A2(_11384_));
 sg13g2_nand2_1 _17903_ (.Y(_11387_),
    .A(net742),
    .B(\mem.mem_internal.code_mem[145][2] ));
 sg13g2_buf_1 _17904_ (.A(_11171_),
    .X(_11388_));
 sg13g2_nand2_1 _17905_ (.Y(_11389_),
    .A(net1148),
    .B(_11380_));
 sg13g2_o21ai_1 _17906_ (.B1(_11389_),
    .Y(_00516_),
    .A1(net258),
    .A2(_11387_));
 sg13g2_nand2_1 _17907_ (.Y(_11390_),
    .A(_11367_),
    .B(\mem.mem_internal.code_mem[145][3] ));
 sg13g2_buf_1 _17908_ (.A(_11175_),
    .X(_11391_));
 sg13g2_nand2_1 _17909_ (.Y(_11392_),
    .A(net1147),
    .B(_11380_));
 sg13g2_o21ai_1 _17910_ (.B1(_11392_),
    .Y(_00517_),
    .A1(net258),
    .A2(_11390_));
 sg13g2_nand2_1 _17911_ (.Y(_11393_),
    .A(_11367_),
    .B(\mem.mem_internal.code_mem[145][4] ));
 sg13g2_buf_1 _17912_ (.A(_11179_),
    .X(_11394_));
 sg13g2_nand2_1 _17913_ (.Y(_11395_),
    .A(net1146),
    .B(_11380_));
 sg13g2_o21ai_1 _17914_ (.B1(_11395_),
    .Y(_00518_),
    .A1(_11381_),
    .A2(_11393_));
 sg13g2_nand2_1 _17915_ (.Y(_11396_),
    .A(net742),
    .B(\mem.mem_internal.code_mem[145][5] ));
 sg13g2_buf_1 _17916_ (.A(_11183_),
    .X(_11397_));
 sg13g2_nand2_1 _17917_ (.Y(_11398_),
    .A(net1145),
    .B(_11380_));
 sg13g2_o21ai_1 _17918_ (.B1(_11398_),
    .Y(_00519_),
    .A1(_11381_),
    .A2(_11396_));
 sg13g2_buf_1 _17919_ (.A(_11247_),
    .X(_11399_));
 sg13g2_nand2_1 _17920_ (.Y(_11400_),
    .A(net741),
    .B(\mem.mem_internal.code_mem[145][6] ));
 sg13g2_buf_1 _17921_ (.A(_11188_),
    .X(_11401_));
 sg13g2_nand2_1 _17922_ (.Y(_11402_),
    .A(net1144),
    .B(_11380_));
 sg13g2_o21ai_1 _17923_ (.B1(_11402_),
    .Y(_00520_),
    .A1(net258),
    .A2(_11400_));
 sg13g2_nand2_1 _17924_ (.Y(_11403_),
    .A(net741),
    .B(\mem.mem_internal.code_mem[145][7] ));
 sg13g2_buf_1 _17925_ (.A(_11192_),
    .X(_11404_));
 sg13g2_nand2_1 _17926_ (.Y(_11405_),
    .A(net1143),
    .B(_11380_));
 sg13g2_o21ai_1 _17927_ (.B1(_11405_),
    .Y(_00521_),
    .A1(net258),
    .A2(_11403_));
 sg13g2_nand2_1 _17928_ (.Y(_11406_),
    .A(net848),
    .B(\mem.mem_internal.code_mem[146][0] ));
 sg13g2_nor2_1 _17929_ (.A(net527),
    .B(_11358_),
    .Y(_11407_));
 sg13g2_buf_2 _17930_ (.A(_11407_),
    .X(_11408_));
 sg13g2_buf_1 _17931_ (.A(_11408_),
    .X(_11409_));
 sg13g2_nand2_1 _17932_ (.Y(_11410_),
    .A(_11382_),
    .B(net257));
 sg13g2_o21ai_1 _17933_ (.B1(_11410_),
    .Y(_00522_),
    .A1(_11406_),
    .A2(net257));
 sg13g2_nand2_1 _17934_ (.Y(_11411_),
    .A(net741),
    .B(\mem.mem_internal.code_mem[146][1] ));
 sg13g2_nand2_1 _17935_ (.Y(_11412_),
    .A(net1149),
    .B(net257));
 sg13g2_o21ai_1 _17936_ (.B1(_11412_),
    .Y(_00523_),
    .A1(net257),
    .A2(_11411_));
 sg13g2_nand2_1 _17937_ (.Y(_11413_),
    .A(net741),
    .B(\mem.mem_internal.code_mem[146][2] ));
 sg13g2_nand2_1 _17938_ (.Y(_11414_),
    .A(net1148),
    .B(_11408_));
 sg13g2_o21ai_1 _17939_ (.B1(_11414_),
    .Y(_00524_),
    .A1(_11409_),
    .A2(_11413_));
 sg13g2_nand2_1 _17940_ (.Y(_11415_),
    .A(_11399_),
    .B(\mem.mem_internal.code_mem[146][3] ));
 sg13g2_nand2_1 _17941_ (.Y(_11416_),
    .A(net1147),
    .B(_11408_));
 sg13g2_o21ai_1 _17942_ (.B1(_11416_),
    .Y(_00525_),
    .A1(net257),
    .A2(_11415_));
 sg13g2_nand2_1 _17943_ (.Y(_11417_),
    .A(net741),
    .B(\mem.mem_internal.code_mem[146][4] ));
 sg13g2_nand2_1 _17944_ (.Y(_11418_),
    .A(net1146),
    .B(_11408_));
 sg13g2_o21ai_1 _17945_ (.B1(_11418_),
    .Y(_00526_),
    .A1(_11409_),
    .A2(_11417_));
 sg13g2_nand2_1 _17946_ (.Y(_11419_),
    .A(net741),
    .B(\mem.mem_internal.code_mem[146][5] ));
 sg13g2_nand2_1 _17947_ (.Y(_11420_),
    .A(net1145),
    .B(_11408_));
 sg13g2_o21ai_1 _17948_ (.B1(_11420_),
    .Y(_00527_),
    .A1(net257),
    .A2(_11419_));
 sg13g2_nand2_1 _17949_ (.Y(_11421_),
    .A(net741),
    .B(\mem.mem_internal.code_mem[146][6] ));
 sg13g2_nand2_1 _17950_ (.Y(_11422_),
    .A(net1144),
    .B(_11408_));
 sg13g2_o21ai_1 _17951_ (.B1(_11422_),
    .Y(_00528_),
    .A1(net257),
    .A2(_11421_));
 sg13g2_nand2_1 _17952_ (.Y(_11423_),
    .A(net741),
    .B(\mem.mem_internal.code_mem[146][7] ));
 sg13g2_nand2_1 _17953_ (.Y(_11424_),
    .A(_11404_),
    .B(_11408_));
 sg13g2_o21ai_1 _17954_ (.B1(_11424_),
    .Y(_00529_),
    .A1(net257),
    .A2(_11423_));
 sg13g2_nand2_1 _17955_ (.Y(_11425_),
    .A(net848),
    .B(\mem.mem_internal.code_mem[147][0] ));
 sg13g2_nor2_1 _17956_ (.A(net526),
    .B(net466),
    .Y(_11426_));
 sg13g2_buf_2 _17957_ (.A(_11426_),
    .X(_11427_));
 sg13g2_buf_1 _17958_ (.A(_11427_),
    .X(_11428_));
 sg13g2_nand2_1 _17959_ (.Y(_11429_),
    .A(net1150),
    .B(net256));
 sg13g2_o21ai_1 _17960_ (.B1(_11429_),
    .Y(_00530_),
    .A1(_11425_),
    .A2(net256));
 sg13g2_nand2_1 _17961_ (.Y(_11430_),
    .A(_11399_),
    .B(\mem.mem_internal.code_mem[147][1] ));
 sg13g2_nand2_1 _17962_ (.Y(_11431_),
    .A(net1149),
    .B(_11428_));
 sg13g2_o21ai_1 _17963_ (.B1(_11431_),
    .Y(_00531_),
    .A1(net256),
    .A2(_11430_));
 sg13g2_buf_1 _17964_ (.A(_11247_),
    .X(_11432_));
 sg13g2_nand2_1 _17965_ (.Y(_11433_),
    .A(net740),
    .B(\mem.mem_internal.code_mem[147][2] ));
 sg13g2_nand2_1 _17966_ (.Y(_11434_),
    .A(net1148),
    .B(_11427_));
 sg13g2_o21ai_1 _17967_ (.B1(_11434_),
    .Y(_00532_),
    .A1(_11428_),
    .A2(_11433_));
 sg13g2_nand2_1 _17968_ (.Y(_11435_),
    .A(net740),
    .B(\mem.mem_internal.code_mem[147][3] ));
 sg13g2_nand2_1 _17969_ (.Y(_11436_),
    .A(net1147),
    .B(_11427_));
 sg13g2_o21ai_1 _17970_ (.B1(_11436_),
    .Y(_00533_),
    .A1(net256),
    .A2(_11435_));
 sg13g2_nand2_1 _17971_ (.Y(_11437_),
    .A(net740),
    .B(\mem.mem_internal.code_mem[147][4] ));
 sg13g2_nand2_1 _17972_ (.Y(_11438_),
    .A(net1146),
    .B(_11427_));
 sg13g2_o21ai_1 _17973_ (.B1(_11438_),
    .Y(_00534_),
    .A1(net256),
    .A2(_11437_));
 sg13g2_nand2_1 _17974_ (.Y(_11439_),
    .A(_11432_),
    .B(\mem.mem_internal.code_mem[147][5] ));
 sg13g2_nand2_1 _17975_ (.Y(_11440_),
    .A(_11397_),
    .B(_11427_));
 sg13g2_o21ai_1 _17976_ (.B1(_11440_),
    .Y(_00535_),
    .A1(net256),
    .A2(_11439_));
 sg13g2_nand2_1 _17977_ (.Y(_11441_),
    .A(net740),
    .B(\mem.mem_internal.code_mem[147][6] ));
 sg13g2_nand2_1 _17978_ (.Y(_11442_),
    .A(_11401_),
    .B(_11427_));
 sg13g2_o21ai_1 _17979_ (.B1(_11442_),
    .Y(_00536_),
    .A1(net256),
    .A2(_11441_));
 sg13g2_nand2_1 _17980_ (.Y(_11443_),
    .A(net740),
    .B(\mem.mem_internal.code_mem[147][7] ));
 sg13g2_nand2_1 _17981_ (.Y(_11444_),
    .A(net1143),
    .B(_11427_));
 sg13g2_o21ai_1 _17982_ (.B1(_11444_),
    .Y(_00537_),
    .A1(net256),
    .A2(_11443_));
 sg13g2_nand2_1 _17983_ (.Y(_11445_),
    .A(net848),
    .B(\mem.mem_internal.code_mem[148][0] ));
 sg13g2_nor2_1 _17984_ (.A(net556),
    .B(net466),
    .Y(_11446_));
 sg13g2_buf_2 _17985_ (.A(_11446_),
    .X(_11447_));
 sg13g2_buf_1 _17986_ (.A(_11447_),
    .X(_11448_));
 sg13g2_nand2_1 _17987_ (.Y(_11449_),
    .A(net1150),
    .B(net255));
 sg13g2_o21ai_1 _17988_ (.B1(_11449_),
    .Y(_00538_),
    .A1(_11445_),
    .A2(net255));
 sg13g2_nand2_1 _17989_ (.Y(_11450_),
    .A(_11432_),
    .B(\mem.mem_internal.code_mem[148][1] ));
 sg13g2_nand2_1 _17990_ (.Y(_11451_),
    .A(net1149),
    .B(net255));
 sg13g2_o21ai_1 _17991_ (.B1(_11451_),
    .Y(_00539_),
    .A1(net255),
    .A2(_11450_));
 sg13g2_nand2_1 _17992_ (.Y(_11452_),
    .A(net740),
    .B(\mem.mem_internal.code_mem[148][2] ));
 sg13g2_nand2_1 _17993_ (.Y(_11453_),
    .A(net1148),
    .B(_11447_));
 sg13g2_o21ai_1 _17994_ (.B1(_11453_),
    .Y(_00540_),
    .A1(net255),
    .A2(_11452_));
 sg13g2_nand2_1 _17995_ (.Y(_11454_),
    .A(net740),
    .B(\mem.mem_internal.code_mem[148][3] ));
 sg13g2_nand2_1 _17996_ (.Y(_11455_),
    .A(net1147),
    .B(_11447_));
 sg13g2_o21ai_1 _17997_ (.B1(_11455_),
    .Y(_00541_),
    .A1(net255),
    .A2(_11454_));
 sg13g2_nand2_1 _17998_ (.Y(_11456_),
    .A(net740),
    .B(\mem.mem_internal.code_mem[148][4] ));
 sg13g2_nand2_1 _17999_ (.Y(_11457_),
    .A(net1146),
    .B(_11447_));
 sg13g2_o21ai_1 _18000_ (.B1(_11457_),
    .Y(_00542_),
    .A1(_11448_),
    .A2(_11456_));
 sg13g2_buf_1 _18001_ (.A(_10415_),
    .X(_11458_));
 sg13g2_buf_1 _18002_ (.A(_11458_),
    .X(_11459_));
 sg13g2_nand2_1 _18003_ (.Y(_11460_),
    .A(net739),
    .B(\mem.mem_internal.code_mem[148][5] ));
 sg13g2_nand2_1 _18004_ (.Y(_11461_),
    .A(net1145),
    .B(_11447_));
 sg13g2_o21ai_1 _18005_ (.B1(_11461_),
    .Y(_00543_),
    .A1(_11448_),
    .A2(_11460_));
 sg13g2_nand2_1 _18006_ (.Y(_11462_),
    .A(net739),
    .B(\mem.mem_internal.code_mem[148][6] ));
 sg13g2_nand2_1 _18007_ (.Y(_11463_),
    .A(net1144),
    .B(_11447_));
 sg13g2_o21ai_1 _18008_ (.B1(_11463_),
    .Y(_00544_),
    .A1(net255),
    .A2(_11462_));
 sg13g2_nand2_1 _18009_ (.Y(_11464_),
    .A(net739),
    .B(\mem.mem_internal.code_mem[148][7] ));
 sg13g2_nand2_1 _18010_ (.Y(_11465_),
    .A(net1143),
    .B(_11447_));
 sg13g2_o21ai_1 _18011_ (.B1(_11465_),
    .Y(_00545_),
    .A1(net255),
    .A2(_11464_));
 sg13g2_nand2_1 _18012_ (.Y(_11466_),
    .A(net848),
    .B(\mem.mem_internal.code_mem[149][0] ));
 sg13g2_nor2_1 _18013_ (.A(net555),
    .B(net466),
    .Y(_11467_));
 sg13g2_buf_2 _18014_ (.A(_11467_),
    .X(_11468_));
 sg13g2_buf_1 _18015_ (.A(_11468_),
    .X(_11469_));
 sg13g2_nand2_1 _18016_ (.Y(_11470_),
    .A(net1150),
    .B(net254));
 sg13g2_o21ai_1 _18017_ (.B1(_11470_),
    .Y(_00546_),
    .A1(_11466_),
    .A2(net254));
 sg13g2_nand2_1 _18018_ (.Y(_11471_),
    .A(net739),
    .B(\mem.mem_internal.code_mem[149][1] ));
 sg13g2_nand2_1 _18019_ (.Y(_11472_),
    .A(net1149),
    .B(net254));
 sg13g2_o21ai_1 _18020_ (.B1(_11472_),
    .Y(_00547_),
    .A1(net254),
    .A2(_11471_));
 sg13g2_nand2_1 _18021_ (.Y(_11473_),
    .A(net739),
    .B(\mem.mem_internal.code_mem[149][2] ));
 sg13g2_nand2_1 _18022_ (.Y(_11474_),
    .A(net1148),
    .B(_11468_));
 sg13g2_o21ai_1 _18023_ (.B1(_11474_),
    .Y(_00548_),
    .A1(net254),
    .A2(_11473_));
 sg13g2_nand2_1 _18024_ (.Y(_11475_),
    .A(net739),
    .B(\mem.mem_internal.code_mem[149][3] ));
 sg13g2_nand2_1 _18025_ (.Y(_11476_),
    .A(net1147),
    .B(_11468_));
 sg13g2_o21ai_1 _18026_ (.B1(_11476_),
    .Y(_00549_),
    .A1(net254),
    .A2(_11475_));
 sg13g2_nand2_1 _18027_ (.Y(_11477_),
    .A(_11459_),
    .B(\mem.mem_internal.code_mem[149][4] ));
 sg13g2_nand2_1 _18028_ (.Y(_11478_),
    .A(net1146),
    .B(_11468_));
 sg13g2_o21ai_1 _18029_ (.B1(_11478_),
    .Y(_00550_),
    .A1(_11469_),
    .A2(_11477_));
 sg13g2_nand2_1 _18030_ (.Y(_11479_),
    .A(_11459_),
    .B(\mem.mem_internal.code_mem[149][5] ));
 sg13g2_nand2_1 _18031_ (.Y(_11480_),
    .A(net1145),
    .B(_11468_));
 sg13g2_o21ai_1 _18032_ (.B1(_11480_),
    .Y(_00551_),
    .A1(_11469_),
    .A2(_11479_));
 sg13g2_nand2_1 _18033_ (.Y(_11481_),
    .A(net739),
    .B(\mem.mem_internal.code_mem[149][6] ));
 sg13g2_nand2_1 _18034_ (.Y(_11482_),
    .A(net1144),
    .B(_11468_));
 sg13g2_o21ai_1 _18035_ (.B1(_11482_),
    .Y(_00552_),
    .A1(net254),
    .A2(_11481_));
 sg13g2_nand2_1 _18036_ (.Y(_11483_),
    .A(net739),
    .B(\mem.mem_internal.code_mem[149][7] ));
 sg13g2_nand2_1 _18037_ (.Y(_11484_),
    .A(net1143),
    .B(_11468_));
 sg13g2_o21ai_1 _18038_ (.B1(_11484_),
    .Y(_00553_),
    .A1(net254),
    .A2(_11483_));
 sg13g2_buf_1 _18039_ (.A(_11058_),
    .X(_11485_));
 sg13g2_nand2_1 _18040_ (.Y(_11486_),
    .A(net847),
    .B(\mem.mem_internal.code_mem[14][0] ));
 sg13g2_nor2_1 _18041_ (.A(net470),
    .B(net547),
    .Y(_11487_));
 sg13g2_buf_2 _18042_ (.A(_11487_),
    .X(_11488_));
 sg13g2_buf_1 _18043_ (.A(_11488_),
    .X(_11489_));
 sg13g2_nand2_1 _18044_ (.Y(_11490_),
    .A(net1150),
    .B(net253));
 sg13g2_o21ai_1 _18045_ (.B1(_11490_),
    .Y(_00554_),
    .A1(_11486_),
    .A2(net253));
 sg13g2_buf_1 _18046_ (.A(_11458_),
    .X(_11491_));
 sg13g2_nand2_1 _18047_ (.Y(_11492_),
    .A(net738),
    .B(\mem.mem_internal.code_mem[14][1] ));
 sg13g2_nand2_1 _18048_ (.Y(_11493_),
    .A(_11385_),
    .B(net253));
 sg13g2_o21ai_1 _18049_ (.B1(_11493_),
    .Y(_00555_),
    .A1(_11489_),
    .A2(_11492_));
 sg13g2_nand2_1 _18050_ (.Y(_11494_),
    .A(net738),
    .B(\mem.mem_internal.code_mem[14][2] ));
 sg13g2_nand2_1 _18051_ (.Y(_11495_),
    .A(_11388_),
    .B(_11488_));
 sg13g2_o21ai_1 _18052_ (.B1(_11495_),
    .Y(_00556_),
    .A1(net253),
    .A2(_11494_));
 sg13g2_nand2_1 _18053_ (.Y(_11496_),
    .A(net738),
    .B(\mem.mem_internal.code_mem[14][3] ));
 sg13g2_nand2_1 _18054_ (.Y(_11497_),
    .A(_11391_),
    .B(_11488_));
 sg13g2_o21ai_1 _18055_ (.B1(_11497_),
    .Y(_00557_),
    .A1(net253),
    .A2(_11496_));
 sg13g2_nand2_1 _18056_ (.Y(_11498_),
    .A(net738),
    .B(\mem.mem_internal.code_mem[14][4] ));
 sg13g2_nand2_1 _18057_ (.Y(_11499_),
    .A(net1146),
    .B(_11488_));
 sg13g2_o21ai_1 _18058_ (.B1(_11499_),
    .Y(_00558_),
    .A1(net253),
    .A2(_11498_));
 sg13g2_nand2_1 _18059_ (.Y(_11500_),
    .A(net738),
    .B(\mem.mem_internal.code_mem[14][5] ));
 sg13g2_nand2_1 _18060_ (.Y(_11501_),
    .A(_11397_),
    .B(_11488_));
 sg13g2_o21ai_1 _18061_ (.B1(_11501_),
    .Y(_00559_),
    .A1(_11489_),
    .A2(_11500_));
 sg13g2_nand2_1 _18062_ (.Y(_11502_),
    .A(_11491_),
    .B(\mem.mem_internal.code_mem[14][6] ));
 sg13g2_nand2_1 _18063_ (.Y(_11503_),
    .A(_11401_),
    .B(_11488_));
 sg13g2_o21ai_1 _18064_ (.B1(_11503_),
    .Y(_00560_),
    .A1(net253),
    .A2(_11502_));
 sg13g2_nand2_1 _18065_ (.Y(_11504_),
    .A(_11491_),
    .B(\mem.mem_internal.code_mem[14][7] ));
 sg13g2_nand2_1 _18066_ (.Y(_11505_),
    .A(_11404_),
    .B(_11488_));
 sg13g2_o21ai_1 _18067_ (.B1(_11505_),
    .Y(_00561_),
    .A1(net253),
    .A2(_11504_));
 sg13g2_nand2_1 _18068_ (.Y(_11506_),
    .A(net847),
    .B(\mem.mem_internal.code_mem[150][0] ));
 sg13g2_nor2_1 _18069_ (.A(net554),
    .B(net466),
    .Y(_11507_));
 sg13g2_buf_2 _18070_ (.A(_11507_),
    .X(_11508_));
 sg13g2_buf_1 _18071_ (.A(_11508_),
    .X(_11509_));
 sg13g2_nand2_1 _18072_ (.Y(_11510_),
    .A(net1150),
    .B(net252));
 sg13g2_o21ai_1 _18073_ (.B1(_11510_),
    .Y(_00562_),
    .A1(_11506_),
    .A2(net252));
 sg13g2_nand2_1 _18074_ (.Y(_11511_),
    .A(net738),
    .B(\mem.mem_internal.code_mem[150][1] ));
 sg13g2_nand2_1 _18075_ (.Y(_11512_),
    .A(_11385_),
    .B(_11509_));
 sg13g2_o21ai_1 _18076_ (.B1(_11512_),
    .Y(_00563_),
    .A1(net252),
    .A2(_11511_));
 sg13g2_nand2_1 _18077_ (.Y(_11513_),
    .A(net738),
    .B(\mem.mem_internal.code_mem[150][2] ));
 sg13g2_nand2_1 _18078_ (.Y(_11514_),
    .A(_11388_),
    .B(_11508_));
 sg13g2_o21ai_1 _18079_ (.B1(_11514_),
    .Y(_00564_),
    .A1(_11509_),
    .A2(_11513_));
 sg13g2_nand2_1 _18080_ (.Y(_11515_),
    .A(net738),
    .B(\mem.mem_internal.code_mem[150][3] ));
 sg13g2_nand2_1 _18081_ (.Y(_11516_),
    .A(_11391_),
    .B(_11508_));
 sg13g2_o21ai_1 _18082_ (.B1(_11516_),
    .Y(_00565_),
    .A1(net252),
    .A2(_11515_));
 sg13g2_buf_1 _18083_ (.A(_11458_),
    .X(_11517_));
 sg13g2_nand2_1 _18084_ (.Y(_11518_),
    .A(net737),
    .B(\mem.mem_internal.code_mem[150][4] ));
 sg13g2_nand2_1 _18085_ (.Y(_11519_),
    .A(_11394_),
    .B(_11508_));
 sg13g2_o21ai_1 _18086_ (.B1(_11519_),
    .Y(_00566_),
    .A1(net252),
    .A2(_11518_));
 sg13g2_nand2_1 _18087_ (.Y(_11520_),
    .A(net737),
    .B(\mem.mem_internal.code_mem[150][5] ));
 sg13g2_nand2_1 _18088_ (.Y(_11521_),
    .A(net1145),
    .B(_11508_));
 sg13g2_o21ai_1 _18089_ (.B1(_11521_),
    .Y(_00567_),
    .A1(net252),
    .A2(_11520_));
 sg13g2_nand2_1 _18090_ (.Y(_11522_),
    .A(net737),
    .B(\mem.mem_internal.code_mem[150][6] ));
 sg13g2_nand2_1 _18091_ (.Y(_11523_),
    .A(net1144),
    .B(_11508_));
 sg13g2_o21ai_1 _18092_ (.B1(_11523_),
    .Y(_00568_),
    .A1(net252),
    .A2(_11522_));
 sg13g2_nand2_1 _18093_ (.Y(_11524_),
    .A(net737),
    .B(\mem.mem_internal.code_mem[150][7] ));
 sg13g2_nand2_1 _18094_ (.Y(_11525_),
    .A(net1143),
    .B(_11508_));
 sg13g2_o21ai_1 _18095_ (.B1(_11525_),
    .Y(_00569_),
    .A1(net252),
    .A2(_11524_));
 sg13g2_nand2_1 _18096_ (.Y(_11526_),
    .A(_11485_),
    .B(\mem.mem_internal.code_mem[151][0] ));
 sg13g2_nor2_1 _18097_ (.A(net553),
    .B(net466),
    .Y(_11527_));
 sg13g2_buf_2 _18098_ (.A(_11527_),
    .X(_11528_));
 sg13g2_buf_1 _18099_ (.A(_11528_),
    .X(_11529_));
 sg13g2_nand2_1 _18100_ (.Y(_11530_),
    .A(net1150),
    .B(net251));
 sg13g2_o21ai_1 _18101_ (.B1(_11530_),
    .Y(_00570_),
    .A1(_11526_),
    .A2(net251));
 sg13g2_nand2_1 _18102_ (.Y(_11531_),
    .A(net737),
    .B(\mem.mem_internal.code_mem[151][1] ));
 sg13g2_nand2_1 _18103_ (.Y(_11532_),
    .A(net1149),
    .B(net251));
 sg13g2_o21ai_1 _18104_ (.B1(_11532_),
    .Y(_00571_),
    .A1(net251),
    .A2(_11531_));
 sg13g2_nand2_1 _18105_ (.Y(_11533_),
    .A(net737),
    .B(\mem.mem_internal.code_mem[151][2] ));
 sg13g2_nand2_1 _18106_ (.Y(_11534_),
    .A(net1148),
    .B(_11528_));
 sg13g2_o21ai_1 _18107_ (.B1(_11534_),
    .Y(_00572_),
    .A1(net251),
    .A2(_11533_));
 sg13g2_nand2_1 _18108_ (.Y(_11535_),
    .A(_11517_),
    .B(\mem.mem_internal.code_mem[151][3] ));
 sg13g2_nand2_1 _18109_ (.Y(_11536_),
    .A(net1147),
    .B(_11528_));
 sg13g2_o21ai_1 _18110_ (.B1(_11536_),
    .Y(_00573_),
    .A1(net251),
    .A2(_11535_));
 sg13g2_nand2_1 _18111_ (.Y(_11537_),
    .A(_11517_),
    .B(\mem.mem_internal.code_mem[151][4] ));
 sg13g2_nand2_1 _18112_ (.Y(_11538_),
    .A(_11394_),
    .B(_11528_));
 sg13g2_o21ai_1 _18113_ (.B1(_11538_),
    .Y(_00574_),
    .A1(_11529_),
    .A2(_11537_));
 sg13g2_nand2_1 _18114_ (.Y(_11539_),
    .A(net737),
    .B(\mem.mem_internal.code_mem[151][5] ));
 sg13g2_nand2_1 _18115_ (.Y(_11540_),
    .A(net1145),
    .B(_11528_));
 sg13g2_o21ai_1 _18116_ (.B1(_11540_),
    .Y(_00575_),
    .A1(_11529_),
    .A2(_11539_));
 sg13g2_nand2_1 _18117_ (.Y(_11541_),
    .A(net737),
    .B(\mem.mem_internal.code_mem[151][6] ));
 sg13g2_nand2_1 _18118_ (.Y(_11542_),
    .A(net1144),
    .B(_11528_));
 sg13g2_o21ai_1 _18119_ (.B1(_11542_),
    .Y(_00576_),
    .A1(net251),
    .A2(_11541_));
 sg13g2_buf_1 _18120_ (.A(_11458_),
    .X(_11543_));
 sg13g2_nand2_1 _18121_ (.Y(_11544_),
    .A(_11543_),
    .B(\mem.mem_internal.code_mem[151][7] ));
 sg13g2_nand2_1 _18122_ (.Y(_11545_),
    .A(net1143),
    .B(_11528_));
 sg13g2_o21ai_1 _18123_ (.B1(_11545_),
    .Y(_00577_),
    .A1(net251),
    .A2(_11544_));
 sg13g2_nand2_1 _18124_ (.Y(_11546_),
    .A(net847),
    .B(\mem.mem_internal.code_mem[152][0] ));
 sg13g2_nor2_1 _18125_ (.A(net552),
    .B(net466),
    .Y(_11547_));
 sg13g2_buf_2 _18126_ (.A(_11547_),
    .X(_11548_));
 sg13g2_buf_1 _18127_ (.A(_11548_),
    .X(_11549_));
 sg13g2_nand2_1 _18128_ (.Y(_11550_),
    .A(net1150),
    .B(_11549_));
 sg13g2_o21ai_1 _18129_ (.B1(_11550_),
    .Y(_00578_),
    .A1(_11546_),
    .A2(net250));
 sg13g2_nand2_1 _18130_ (.Y(_11551_),
    .A(net736),
    .B(\mem.mem_internal.code_mem[152][1] ));
 sg13g2_nand2_1 _18131_ (.Y(_11552_),
    .A(net1149),
    .B(net250));
 sg13g2_o21ai_1 _18132_ (.B1(_11552_),
    .Y(_00579_),
    .A1(net250),
    .A2(_11551_));
 sg13g2_nand2_1 _18133_ (.Y(_11553_),
    .A(net736),
    .B(\mem.mem_internal.code_mem[152][2] ));
 sg13g2_nand2_1 _18134_ (.Y(_11554_),
    .A(net1148),
    .B(_11548_));
 sg13g2_o21ai_1 _18135_ (.B1(_11554_),
    .Y(_00580_),
    .A1(net250),
    .A2(_11553_));
 sg13g2_nand2_1 _18136_ (.Y(_11555_),
    .A(net736),
    .B(\mem.mem_internal.code_mem[152][3] ));
 sg13g2_nand2_1 _18137_ (.Y(_11556_),
    .A(net1147),
    .B(_11548_));
 sg13g2_o21ai_1 _18138_ (.B1(_11556_),
    .Y(_00581_),
    .A1(_11549_),
    .A2(_11555_));
 sg13g2_nand2_1 _18139_ (.Y(_11557_),
    .A(net736),
    .B(\mem.mem_internal.code_mem[152][4] ));
 sg13g2_nand2_1 _18140_ (.Y(_11558_),
    .A(net1146),
    .B(_11548_));
 sg13g2_o21ai_1 _18141_ (.B1(_11558_),
    .Y(_00582_),
    .A1(net250),
    .A2(_11557_));
 sg13g2_nand2_1 _18142_ (.Y(_11559_),
    .A(net736),
    .B(\mem.mem_internal.code_mem[152][5] ));
 sg13g2_nand2_1 _18143_ (.Y(_11560_),
    .A(net1145),
    .B(_11548_));
 sg13g2_o21ai_1 _18144_ (.B1(_11560_),
    .Y(_00583_),
    .A1(net250),
    .A2(_11559_));
 sg13g2_nand2_1 _18145_ (.Y(_11561_),
    .A(net736),
    .B(\mem.mem_internal.code_mem[152][6] ));
 sg13g2_nand2_1 _18146_ (.Y(_11562_),
    .A(net1144),
    .B(_11548_));
 sg13g2_o21ai_1 _18147_ (.B1(_11562_),
    .Y(_00584_),
    .A1(net250),
    .A2(_11561_));
 sg13g2_nand2_1 _18148_ (.Y(_11563_),
    .A(net736),
    .B(\mem.mem_internal.code_mem[152][7] ));
 sg13g2_nand2_1 _18149_ (.Y(_11564_),
    .A(net1143),
    .B(_11548_));
 sg13g2_o21ai_1 _18150_ (.B1(_11564_),
    .Y(_00585_),
    .A1(net250),
    .A2(_11563_));
 sg13g2_nand2_1 _18151_ (.Y(_11565_),
    .A(_11485_),
    .B(\mem.mem_internal.code_mem[153][0] ));
 sg13g2_nor2_1 _18152_ (.A(net551),
    .B(net466),
    .Y(_11566_));
 sg13g2_buf_2 _18153_ (.A(_11566_),
    .X(_11567_));
 sg13g2_buf_1 _18154_ (.A(_11567_),
    .X(_11568_));
 sg13g2_nand2_1 _18155_ (.Y(_11569_),
    .A(net1150),
    .B(_11568_));
 sg13g2_o21ai_1 _18156_ (.B1(_11569_),
    .Y(_00586_),
    .A1(_11565_),
    .A2(net249));
 sg13g2_nand2_1 _18157_ (.Y(_11570_),
    .A(net736),
    .B(\mem.mem_internal.code_mem[153][1] ));
 sg13g2_nand2_1 _18158_ (.Y(_11571_),
    .A(net1149),
    .B(net249));
 sg13g2_o21ai_1 _18159_ (.B1(_11571_),
    .Y(_00587_),
    .A1(net249),
    .A2(_11570_));
 sg13g2_nand2_1 _18160_ (.Y(_11572_),
    .A(_11543_),
    .B(\mem.mem_internal.code_mem[153][2] ));
 sg13g2_nand2_1 _18161_ (.Y(_11573_),
    .A(net1148),
    .B(_11567_));
 sg13g2_o21ai_1 _18162_ (.B1(_11573_),
    .Y(_00588_),
    .A1(net249),
    .A2(_11572_));
 sg13g2_buf_1 _18163_ (.A(_11458_),
    .X(_11574_));
 sg13g2_nand2_1 _18164_ (.Y(_11575_),
    .A(net735),
    .B(\mem.mem_internal.code_mem[153][3] ));
 sg13g2_nand2_1 _18165_ (.Y(_11576_),
    .A(net1147),
    .B(_11567_));
 sg13g2_o21ai_1 _18166_ (.B1(_11576_),
    .Y(_00589_),
    .A1(_11568_),
    .A2(_11575_));
 sg13g2_nand2_1 _18167_ (.Y(_11577_),
    .A(net735),
    .B(\mem.mem_internal.code_mem[153][4] ));
 sg13g2_nand2_1 _18168_ (.Y(_11578_),
    .A(net1146),
    .B(_11567_));
 sg13g2_o21ai_1 _18169_ (.B1(_11578_),
    .Y(_00590_),
    .A1(net249),
    .A2(_11577_));
 sg13g2_nand2_1 _18170_ (.Y(_11579_),
    .A(net735),
    .B(\mem.mem_internal.code_mem[153][5] ));
 sg13g2_nand2_1 _18171_ (.Y(_11580_),
    .A(net1145),
    .B(_11567_));
 sg13g2_o21ai_1 _18172_ (.B1(_11580_),
    .Y(_00591_),
    .A1(net249),
    .A2(_11579_));
 sg13g2_nand2_1 _18173_ (.Y(_11581_),
    .A(net735),
    .B(\mem.mem_internal.code_mem[153][6] ));
 sg13g2_nand2_1 _18174_ (.Y(_11582_),
    .A(net1144),
    .B(_11567_));
 sg13g2_o21ai_1 _18175_ (.B1(_11582_),
    .Y(_00592_),
    .A1(net249),
    .A2(_11581_));
 sg13g2_nand2_1 _18176_ (.Y(_11583_),
    .A(net735),
    .B(\mem.mem_internal.code_mem[153][7] ));
 sg13g2_nand2_1 _18177_ (.Y(_11584_),
    .A(net1143),
    .B(_11567_));
 sg13g2_o21ai_1 _18178_ (.B1(_11584_),
    .Y(_00593_),
    .A1(net249),
    .A2(_11583_));
 sg13g2_nand2_1 _18179_ (.Y(_11585_),
    .A(net847),
    .B(\mem.mem_internal.code_mem[154][0] ));
 sg13g2_nor2_1 _18180_ (.A(net550),
    .B(_11357_),
    .Y(_11586_));
 sg13g2_buf_1 _18181_ (.A(_11586_),
    .X(_11587_));
 sg13g2_buf_1 _18182_ (.A(_11587_),
    .X(_11588_));
 sg13g2_buf_1 _18183_ (.A(_11163_),
    .X(_11589_));
 sg13g2_nand2_1 _18184_ (.Y(_11590_),
    .A(net1142),
    .B(_11588_));
 sg13g2_o21ai_1 _18185_ (.B1(_11590_),
    .Y(_00594_),
    .A1(_11585_),
    .A2(_11588_));
 sg13g2_nand2_1 _18186_ (.Y(_11591_),
    .A(net735),
    .B(\mem.mem_internal.code_mem[154][1] ));
 sg13g2_buf_1 _18187_ (.A(_11167_),
    .X(_11592_));
 sg13g2_nand2_1 _18188_ (.Y(_11593_),
    .A(_11592_),
    .B(net384));
 sg13g2_o21ai_1 _18189_ (.B1(_11593_),
    .Y(_00595_),
    .A1(net384),
    .A2(_11591_));
 sg13g2_nand2_1 _18190_ (.Y(_11594_),
    .A(_11574_),
    .B(\mem.mem_internal.code_mem[154][2] ));
 sg13g2_buf_1 _18191_ (.A(_11171_),
    .X(_11595_));
 sg13g2_nand2_1 _18192_ (.Y(_11596_),
    .A(_11595_),
    .B(_11587_));
 sg13g2_o21ai_1 _18193_ (.B1(_11596_),
    .Y(_00596_),
    .A1(net384),
    .A2(_11594_));
 sg13g2_nand2_1 _18194_ (.Y(_11597_),
    .A(_11574_),
    .B(\mem.mem_internal.code_mem[154][3] ));
 sg13g2_buf_1 _18195_ (.A(_11175_),
    .X(_11598_));
 sg13g2_nand2_1 _18196_ (.Y(_11599_),
    .A(_11598_),
    .B(_11587_));
 sg13g2_o21ai_1 _18197_ (.B1(_11599_),
    .Y(_00597_),
    .A1(net384),
    .A2(_11597_));
 sg13g2_nand2_1 _18198_ (.Y(_11600_),
    .A(net735),
    .B(\mem.mem_internal.code_mem[154][4] ));
 sg13g2_buf_1 _18199_ (.A(_11179_),
    .X(_11601_));
 sg13g2_nand2_1 _18200_ (.Y(_11602_),
    .A(net1138),
    .B(_11587_));
 sg13g2_o21ai_1 _18201_ (.B1(_11602_),
    .Y(_00598_),
    .A1(net384),
    .A2(_11600_));
 sg13g2_nand2_1 _18202_ (.Y(_11603_),
    .A(net735),
    .B(\mem.mem_internal.code_mem[154][5] ));
 sg13g2_buf_1 _18203_ (.A(_11183_),
    .X(_11604_));
 sg13g2_nand2_1 _18204_ (.Y(_11605_),
    .A(net1137),
    .B(_11587_));
 sg13g2_o21ai_1 _18205_ (.B1(_11605_),
    .Y(_00599_),
    .A1(net384),
    .A2(_11603_));
 sg13g2_buf_1 _18206_ (.A(_11458_),
    .X(_11606_));
 sg13g2_nand2_1 _18207_ (.Y(_11607_),
    .A(net734),
    .B(\mem.mem_internal.code_mem[154][6] ));
 sg13g2_buf_1 _18208_ (.A(_11188_),
    .X(_11608_));
 sg13g2_nand2_1 _18209_ (.Y(_11609_),
    .A(net1136),
    .B(_11587_));
 sg13g2_o21ai_1 _18210_ (.B1(_11609_),
    .Y(_00600_),
    .A1(net384),
    .A2(_11607_));
 sg13g2_nand2_1 _18211_ (.Y(_11610_),
    .A(net734),
    .B(\mem.mem_internal.code_mem[154][7] ));
 sg13g2_buf_1 _18212_ (.A(_11192_),
    .X(_11611_));
 sg13g2_nand2_1 _18213_ (.Y(_11612_),
    .A(net1135),
    .B(_11587_));
 sg13g2_o21ai_1 _18214_ (.B1(_11612_),
    .Y(_00601_),
    .A1(net384),
    .A2(_11610_));
 sg13g2_nand2_1 _18215_ (.Y(_11613_),
    .A(net847),
    .B(\mem.mem_internal.code_mem[155][0] ));
 sg13g2_nor2_1 _18216_ (.A(net549),
    .B(_11357_),
    .Y(_11614_));
 sg13g2_buf_2 _18217_ (.A(_11614_),
    .X(_11615_));
 sg13g2_buf_1 _18218_ (.A(_11615_),
    .X(_11616_));
 sg13g2_nand2_1 _18219_ (.Y(_11617_),
    .A(_11589_),
    .B(_11616_));
 sg13g2_o21ai_1 _18220_ (.B1(_11617_),
    .Y(_00602_),
    .A1(_11613_),
    .A2(net383));
 sg13g2_nand2_1 _18221_ (.Y(_11618_),
    .A(_11606_),
    .B(\mem.mem_internal.code_mem[155][1] ));
 sg13g2_nand2_1 _18222_ (.Y(_11619_),
    .A(net1141),
    .B(net383));
 sg13g2_o21ai_1 _18223_ (.B1(_11619_),
    .Y(_00603_),
    .A1(net383),
    .A2(_11618_));
 sg13g2_nand2_1 _18224_ (.Y(_11620_),
    .A(_11606_),
    .B(\mem.mem_internal.code_mem[155][2] ));
 sg13g2_nand2_1 _18225_ (.Y(_11621_),
    .A(_11595_),
    .B(_11615_));
 sg13g2_o21ai_1 _18226_ (.B1(_11621_),
    .Y(_00604_),
    .A1(_11616_),
    .A2(_11620_));
 sg13g2_nand2_1 _18227_ (.Y(_11622_),
    .A(net734),
    .B(\mem.mem_internal.code_mem[155][3] ));
 sg13g2_nand2_1 _18228_ (.Y(_11623_),
    .A(_11598_),
    .B(_11615_));
 sg13g2_o21ai_1 _18229_ (.B1(_11623_),
    .Y(_00605_),
    .A1(net383),
    .A2(_11622_));
 sg13g2_nand2_1 _18230_ (.Y(_11624_),
    .A(net734),
    .B(\mem.mem_internal.code_mem[155][4] ));
 sg13g2_nand2_1 _18231_ (.Y(_11625_),
    .A(net1138),
    .B(_11615_));
 sg13g2_o21ai_1 _18232_ (.B1(_11625_),
    .Y(_00606_),
    .A1(net383),
    .A2(_11624_));
 sg13g2_nand2_1 _18233_ (.Y(_11626_),
    .A(net734),
    .B(\mem.mem_internal.code_mem[155][5] ));
 sg13g2_nand2_1 _18234_ (.Y(_11627_),
    .A(net1137),
    .B(_11615_));
 sg13g2_o21ai_1 _18235_ (.B1(_11627_),
    .Y(_00607_),
    .A1(net383),
    .A2(_11626_));
 sg13g2_nand2_1 _18236_ (.Y(_11628_),
    .A(net734),
    .B(\mem.mem_internal.code_mem[155][6] ));
 sg13g2_nand2_1 _18237_ (.Y(_11629_),
    .A(net1136),
    .B(_11615_));
 sg13g2_o21ai_1 _18238_ (.B1(_11629_),
    .Y(_00608_),
    .A1(net383),
    .A2(_11628_));
 sg13g2_nand2_1 _18239_ (.Y(_11630_),
    .A(net734),
    .B(\mem.mem_internal.code_mem[155][7] ));
 sg13g2_nand2_1 _18240_ (.Y(_11631_),
    .A(net1135),
    .B(_11615_));
 sg13g2_o21ai_1 _18241_ (.B1(_11631_),
    .Y(_00609_),
    .A1(net383),
    .A2(_11630_));
 sg13g2_nand2_1 _18242_ (.Y(_11632_),
    .A(net847),
    .B(\mem.mem_internal.code_mem[156][0] ));
 sg13g2_nor2_1 _18243_ (.A(net773),
    .B(_11357_),
    .Y(_11633_));
 sg13g2_buf_2 _18244_ (.A(_11633_),
    .X(_11634_));
 sg13g2_buf_1 _18245_ (.A(_11634_),
    .X(_11635_));
 sg13g2_nand2_1 _18246_ (.Y(_11636_),
    .A(net1142),
    .B(net382));
 sg13g2_o21ai_1 _18247_ (.B1(_11636_),
    .Y(_00610_),
    .A1(_11632_),
    .A2(net382));
 sg13g2_nand2_1 _18248_ (.Y(_11637_),
    .A(net734),
    .B(\mem.mem_internal.code_mem[156][1] ));
 sg13g2_nand2_1 _18249_ (.Y(_11638_),
    .A(net1141),
    .B(net382));
 sg13g2_o21ai_1 _18250_ (.B1(_11638_),
    .Y(_00611_),
    .A1(net382),
    .A2(_11637_));
 sg13g2_buf_1 _18251_ (.A(_11458_),
    .X(_11639_));
 sg13g2_nand2_1 _18252_ (.Y(_11640_),
    .A(net733),
    .B(\mem.mem_internal.code_mem[156][2] ));
 sg13g2_nand2_1 _18253_ (.Y(_11641_),
    .A(net1140),
    .B(_11634_));
 sg13g2_o21ai_1 _18254_ (.B1(_11641_),
    .Y(_00612_),
    .A1(net382),
    .A2(_11640_));
 sg13g2_nand2_1 _18255_ (.Y(_11642_),
    .A(net733),
    .B(\mem.mem_internal.code_mem[156][3] ));
 sg13g2_nand2_1 _18256_ (.Y(_11643_),
    .A(net1139),
    .B(_11634_));
 sg13g2_o21ai_1 _18257_ (.B1(_11643_),
    .Y(_00613_),
    .A1(_11635_),
    .A2(_11642_));
 sg13g2_nand2_1 _18258_ (.Y(_11644_),
    .A(net733),
    .B(\mem.mem_internal.code_mem[156][4] ));
 sg13g2_nand2_1 _18259_ (.Y(_11645_),
    .A(net1138),
    .B(_11634_));
 sg13g2_o21ai_1 _18260_ (.B1(_11645_),
    .Y(_00614_),
    .A1(net382),
    .A2(_11644_));
 sg13g2_nand2_1 _18261_ (.Y(_11646_),
    .A(net733),
    .B(\mem.mem_internal.code_mem[156][5] ));
 sg13g2_nand2_1 _18262_ (.Y(_11647_),
    .A(net1137),
    .B(_11634_));
 sg13g2_o21ai_1 _18263_ (.B1(_11647_),
    .Y(_00615_),
    .A1(net382),
    .A2(_11646_));
 sg13g2_nand2_1 _18264_ (.Y(_11648_),
    .A(_11639_),
    .B(\mem.mem_internal.code_mem[156][6] ));
 sg13g2_nand2_1 _18265_ (.Y(_11649_),
    .A(net1136),
    .B(_11634_));
 sg13g2_o21ai_1 _18266_ (.B1(_11649_),
    .Y(_00616_),
    .A1(net382),
    .A2(_11648_));
 sg13g2_nand2_1 _18267_ (.Y(_11650_),
    .A(net733),
    .B(\mem.mem_internal.code_mem[156][7] ));
 sg13g2_nand2_1 _18268_ (.Y(_11651_),
    .A(net1135),
    .B(_11634_));
 sg13g2_o21ai_1 _18269_ (.B1(_11651_),
    .Y(_00617_),
    .A1(_11635_),
    .A2(_11650_));
 sg13g2_nand2_1 _18270_ (.Y(_11652_),
    .A(net847),
    .B(\mem.mem_internal.code_mem[157][0] ));
 sg13g2_nor2_1 _18271_ (.A(net548),
    .B(_11357_),
    .Y(_11653_));
 sg13g2_buf_2 _18272_ (.A(_11653_),
    .X(_11654_));
 sg13g2_buf_1 _18273_ (.A(_11654_),
    .X(_11655_));
 sg13g2_nand2_1 _18274_ (.Y(_11656_),
    .A(net1142),
    .B(net381));
 sg13g2_o21ai_1 _18275_ (.B1(_11656_),
    .Y(_00618_),
    .A1(_11652_),
    .A2(net381));
 sg13g2_nand2_1 _18276_ (.Y(_11657_),
    .A(net733),
    .B(\mem.mem_internal.code_mem[157][1] ));
 sg13g2_nand2_1 _18277_ (.Y(_11658_),
    .A(net1141),
    .B(net381));
 sg13g2_o21ai_1 _18278_ (.B1(_11658_),
    .Y(_00619_),
    .A1(net381),
    .A2(_11657_));
 sg13g2_nand2_1 _18279_ (.Y(_11659_),
    .A(net733),
    .B(\mem.mem_internal.code_mem[157][2] ));
 sg13g2_nand2_1 _18280_ (.Y(_11660_),
    .A(net1140),
    .B(_11654_));
 sg13g2_o21ai_1 _18281_ (.B1(_11660_),
    .Y(_00620_),
    .A1(net381),
    .A2(_11659_));
 sg13g2_nand2_1 _18282_ (.Y(_11661_),
    .A(_11639_),
    .B(\mem.mem_internal.code_mem[157][3] ));
 sg13g2_nand2_1 _18283_ (.Y(_11662_),
    .A(net1139),
    .B(_11654_));
 sg13g2_o21ai_1 _18284_ (.B1(_11662_),
    .Y(_00621_),
    .A1(_11655_),
    .A2(_11661_));
 sg13g2_nand2_1 _18285_ (.Y(_11663_),
    .A(net733),
    .B(\mem.mem_internal.code_mem[157][4] ));
 sg13g2_nand2_1 _18286_ (.Y(_11664_),
    .A(net1138),
    .B(_11654_));
 sg13g2_o21ai_1 _18287_ (.B1(_11664_),
    .Y(_00622_),
    .A1(net381),
    .A2(_11663_));
 sg13g2_buf_1 _18288_ (.A(_10415_),
    .X(_11665_));
 sg13g2_buf_1 _18289_ (.A(_11665_),
    .X(_11666_));
 sg13g2_nand2_1 _18290_ (.Y(_11667_),
    .A(net732),
    .B(\mem.mem_internal.code_mem[157][5] ));
 sg13g2_nand2_1 _18291_ (.Y(_11668_),
    .A(net1137),
    .B(_11654_));
 sg13g2_o21ai_1 _18292_ (.B1(_11668_),
    .Y(_00623_),
    .A1(net381),
    .A2(_11667_));
 sg13g2_nand2_1 _18293_ (.Y(_11669_),
    .A(net732),
    .B(\mem.mem_internal.code_mem[157][6] ));
 sg13g2_nand2_1 _18294_ (.Y(_11670_),
    .A(net1136),
    .B(_11654_));
 sg13g2_o21ai_1 _18295_ (.B1(_11670_),
    .Y(_00624_),
    .A1(_11655_),
    .A2(_11669_));
 sg13g2_nand2_1 _18296_ (.Y(_11671_),
    .A(_11666_),
    .B(\mem.mem_internal.code_mem[157][7] ));
 sg13g2_nand2_1 _18297_ (.Y(_11672_),
    .A(net1135),
    .B(_11654_));
 sg13g2_o21ai_1 _18298_ (.B1(_11672_),
    .Y(_00625_),
    .A1(net381),
    .A2(_11671_));
 sg13g2_nand2_1 _18299_ (.Y(_11673_),
    .A(net847),
    .B(\mem.mem_internal.code_mem[158][0] ));
 sg13g2_nor2_1 _18300_ (.A(net547),
    .B(_11357_),
    .Y(_11674_));
 sg13g2_buf_2 _18301_ (.A(_11674_),
    .X(_11675_));
 sg13g2_buf_1 _18302_ (.A(_11675_),
    .X(_11676_));
 sg13g2_nand2_1 _18303_ (.Y(_11677_),
    .A(net1142),
    .B(net380));
 sg13g2_o21ai_1 _18304_ (.B1(_11677_),
    .Y(_00626_),
    .A1(_11673_),
    .A2(net380));
 sg13g2_nand2_1 _18305_ (.Y(_11678_),
    .A(net732),
    .B(\mem.mem_internal.code_mem[158][1] ));
 sg13g2_nand2_1 _18306_ (.Y(_11679_),
    .A(net1141),
    .B(net380));
 sg13g2_o21ai_1 _18307_ (.B1(_11679_),
    .Y(_00627_),
    .A1(net380),
    .A2(_11678_));
 sg13g2_nand2_1 _18308_ (.Y(_11680_),
    .A(net732),
    .B(\mem.mem_internal.code_mem[158][2] ));
 sg13g2_nand2_1 _18309_ (.Y(_11681_),
    .A(net1140),
    .B(_11675_));
 sg13g2_o21ai_1 _18310_ (.B1(_11681_),
    .Y(_00628_),
    .A1(_11676_),
    .A2(_11680_));
 sg13g2_nand2_1 _18311_ (.Y(_11682_),
    .A(net732),
    .B(\mem.mem_internal.code_mem[158][3] ));
 sg13g2_nand2_1 _18312_ (.Y(_11683_),
    .A(net1139),
    .B(_11675_));
 sg13g2_o21ai_1 _18313_ (.B1(_11683_),
    .Y(_00629_),
    .A1(_11676_),
    .A2(_11682_));
 sg13g2_nand2_1 _18314_ (.Y(_11684_),
    .A(net732),
    .B(\mem.mem_internal.code_mem[158][4] ));
 sg13g2_nand2_1 _18315_ (.Y(_11685_),
    .A(_11601_),
    .B(_11675_));
 sg13g2_o21ai_1 _18316_ (.B1(_11685_),
    .Y(_00630_),
    .A1(net380),
    .A2(_11684_));
 sg13g2_nand2_1 _18317_ (.Y(_11686_),
    .A(net732),
    .B(\mem.mem_internal.code_mem[158][5] ));
 sg13g2_nand2_1 _18318_ (.Y(_11687_),
    .A(_11604_),
    .B(_11675_));
 sg13g2_o21ai_1 _18319_ (.B1(_11687_),
    .Y(_00631_),
    .A1(net380),
    .A2(_11686_));
 sg13g2_nand2_1 _18320_ (.Y(_11688_),
    .A(net732),
    .B(\mem.mem_internal.code_mem[158][6] ));
 sg13g2_nand2_1 _18321_ (.Y(_11689_),
    .A(_11608_),
    .B(_11675_));
 sg13g2_o21ai_1 _18322_ (.B1(_11689_),
    .Y(_00632_),
    .A1(net380),
    .A2(_11688_));
 sg13g2_nand2_1 _18323_ (.Y(_11690_),
    .A(_11666_),
    .B(\mem.mem_internal.code_mem[158][7] ));
 sg13g2_nand2_1 _18324_ (.Y(_11691_),
    .A(net1135),
    .B(_11675_));
 sg13g2_o21ai_1 _18325_ (.B1(_11691_),
    .Y(_00633_),
    .A1(net380),
    .A2(_11690_));
 sg13g2_buf_1 _18326_ (.A(_11058_),
    .X(_11692_));
 sg13g2_nand2_1 _18327_ (.Y(_11693_),
    .A(net846),
    .B(\mem.mem_internal.code_mem[159][0] ));
 sg13g2_nor2_1 _18328_ (.A(net770),
    .B(_11357_),
    .Y(_11694_));
 sg13g2_buf_2 _18329_ (.A(_11694_),
    .X(_11695_));
 sg13g2_buf_1 _18330_ (.A(_11695_),
    .X(_11696_));
 sg13g2_nand2_1 _18331_ (.Y(_11697_),
    .A(net1142),
    .B(net379));
 sg13g2_o21ai_1 _18332_ (.B1(_11697_),
    .Y(_00634_),
    .A1(_11693_),
    .A2(net379));
 sg13g2_buf_1 _18333_ (.A(_11665_),
    .X(_11698_));
 sg13g2_nand2_1 _18334_ (.Y(_11699_),
    .A(net731),
    .B(\mem.mem_internal.code_mem[159][1] ));
 sg13g2_nand2_1 _18335_ (.Y(_11700_),
    .A(net1141),
    .B(net379));
 sg13g2_o21ai_1 _18336_ (.B1(_11700_),
    .Y(_00635_),
    .A1(net379),
    .A2(_11699_));
 sg13g2_nand2_1 _18337_ (.Y(_11701_),
    .A(net731),
    .B(\mem.mem_internal.code_mem[159][2] ));
 sg13g2_nand2_1 _18338_ (.Y(_11702_),
    .A(net1140),
    .B(_11695_));
 sg13g2_o21ai_1 _18339_ (.B1(_11702_),
    .Y(_00636_),
    .A1(_11696_),
    .A2(_11701_));
 sg13g2_nand2_1 _18340_ (.Y(_11703_),
    .A(_11698_),
    .B(\mem.mem_internal.code_mem[159][3] ));
 sg13g2_nand2_1 _18341_ (.Y(_11704_),
    .A(net1139),
    .B(_11695_));
 sg13g2_o21ai_1 _18342_ (.B1(_11704_),
    .Y(_00637_),
    .A1(_11696_),
    .A2(_11703_));
 sg13g2_nand2_1 _18343_ (.Y(_11705_),
    .A(net731),
    .B(\mem.mem_internal.code_mem[159][4] ));
 sg13g2_nand2_1 _18344_ (.Y(_11706_),
    .A(net1138),
    .B(_11695_));
 sg13g2_o21ai_1 _18345_ (.B1(_11706_),
    .Y(_00638_),
    .A1(net379),
    .A2(_11705_));
 sg13g2_nand2_1 _18346_ (.Y(_11707_),
    .A(net731),
    .B(\mem.mem_internal.code_mem[159][5] ));
 sg13g2_nand2_1 _18347_ (.Y(_11708_),
    .A(net1137),
    .B(_11695_));
 sg13g2_o21ai_1 _18348_ (.B1(_11708_),
    .Y(_00639_),
    .A1(net379),
    .A2(_11707_));
 sg13g2_nand2_1 _18349_ (.Y(_11709_),
    .A(net731),
    .B(\mem.mem_internal.code_mem[159][6] ));
 sg13g2_nand2_1 _18350_ (.Y(_11710_),
    .A(net1136),
    .B(_11695_));
 sg13g2_o21ai_1 _18351_ (.B1(_11710_),
    .Y(_00640_),
    .A1(net379),
    .A2(_11709_));
 sg13g2_nand2_1 _18352_ (.Y(_11711_),
    .A(_11698_),
    .B(\mem.mem_internal.code_mem[159][7] ));
 sg13g2_nand2_1 _18353_ (.Y(_11712_),
    .A(_11611_),
    .B(_11695_));
 sg13g2_o21ai_1 _18354_ (.B1(_11712_),
    .Y(_00641_),
    .A1(net379),
    .A2(_11711_));
 sg13g2_nand2_1 _18355_ (.Y(_11713_),
    .A(net846),
    .B(\mem.mem_internal.code_mem[15][0] ));
 sg13g2_nor2_1 _18356_ (.A(net470),
    .B(net770),
    .Y(_11714_));
 sg13g2_buf_2 _18357_ (.A(_11714_),
    .X(_11715_));
 sg13g2_buf_1 _18358_ (.A(_11715_),
    .X(_11716_));
 sg13g2_nand2_1 _18359_ (.Y(_11717_),
    .A(_11589_),
    .B(net248));
 sg13g2_o21ai_1 _18360_ (.B1(_11717_),
    .Y(_00642_),
    .A1(_11713_),
    .A2(net248));
 sg13g2_nand2_1 _18361_ (.Y(_11718_),
    .A(net731),
    .B(\mem.mem_internal.code_mem[15][1] ));
 sg13g2_nand2_1 _18362_ (.Y(_11719_),
    .A(_11592_),
    .B(net248));
 sg13g2_o21ai_1 _18363_ (.B1(_11719_),
    .Y(_00643_),
    .A1(net248),
    .A2(_11718_));
 sg13g2_nand2_1 _18364_ (.Y(_11720_),
    .A(net731),
    .B(\mem.mem_internal.code_mem[15][2] ));
 sg13g2_nand2_1 _18365_ (.Y(_11721_),
    .A(net1140),
    .B(_11715_));
 sg13g2_o21ai_1 _18366_ (.B1(_11721_),
    .Y(_00644_),
    .A1(net248),
    .A2(_11720_));
 sg13g2_nand2_1 _18367_ (.Y(_11722_),
    .A(net731),
    .B(\mem.mem_internal.code_mem[15][3] ));
 sg13g2_nand2_1 _18368_ (.Y(_11723_),
    .A(net1139),
    .B(_11715_));
 sg13g2_o21ai_1 _18369_ (.B1(_11723_),
    .Y(_00645_),
    .A1(net248),
    .A2(_11722_));
 sg13g2_buf_1 _18370_ (.A(_11665_),
    .X(_11724_));
 sg13g2_nand2_1 _18371_ (.Y(_11725_),
    .A(net730),
    .B(\mem.mem_internal.code_mem[15][4] ));
 sg13g2_nand2_1 _18372_ (.Y(_11726_),
    .A(_11601_),
    .B(_11715_));
 sg13g2_o21ai_1 _18373_ (.B1(_11726_),
    .Y(_00646_),
    .A1(net248),
    .A2(_11725_));
 sg13g2_nand2_1 _18374_ (.Y(_11727_),
    .A(net730),
    .B(\mem.mem_internal.code_mem[15][5] ));
 sg13g2_nand2_1 _18375_ (.Y(_11728_),
    .A(_11604_),
    .B(_11715_));
 sg13g2_o21ai_1 _18376_ (.B1(_11728_),
    .Y(_00647_),
    .A1(net248),
    .A2(_11727_));
 sg13g2_nand2_1 _18377_ (.Y(_11729_),
    .A(_11724_),
    .B(\mem.mem_internal.code_mem[15][6] ));
 sg13g2_nand2_1 _18378_ (.Y(_11730_),
    .A(_11608_),
    .B(_11715_));
 sg13g2_o21ai_1 _18379_ (.B1(_11730_),
    .Y(_00648_),
    .A1(_11716_),
    .A2(_11729_));
 sg13g2_nand2_1 _18380_ (.Y(_11731_),
    .A(_11724_),
    .B(\mem.mem_internal.code_mem[15][7] ));
 sg13g2_nand2_1 _18381_ (.Y(_11732_),
    .A(_11611_),
    .B(_11715_));
 sg13g2_o21ai_1 _18382_ (.B1(_11732_),
    .Y(_00649_),
    .A1(_11716_),
    .A2(_11731_));
 sg13g2_nand2_1 _18383_ (.Y(_11733_),
    .A(net846),
    .B(\mem.mem_internal.code_mem[160][0] ));
 sg13g2_nand2_1 _18384_ (.Y(_11734_),
    .A(_10298_),
    .B(_10976_));
 sg13g2_buf_2 _18385_ (.A(_11734_),
    .X(_11735_));
 sg13g2_buf_1 _18386_ (.A(_11735_),
    .X(_11736_));
 sg13g2_nor2_1 _18387_ (.A(net529),
    .B(net465),
    .Y(_11737_));
 sg13g2_buf_2 _18388_ (.A(_11737_),
    .X(_11738_));
 sg13g2_buf_1 _18389_ (.A(_11738_),
    .X(_11739_));
 sg13g2_nand2_1 _18390_ (.Y(_11740_),
    .A(net1142),
    .B(net247));
 sg13g2_o21ai_1 _18391_ (.B1(_11740_),
    .Y(_00650_),
    .A1(_11733_),
    .A2(net247));
 sg13g2_nand2_1 _18392_ (.Y(_11741_),
    .A(net730),
    .B(\mem.mem_internal.code_mem[160][1] ));
 sg13g2_nand2_1 _18393_ (.Y(_11742_),
    .A(net1141),
    .B(_11739_));
 sg13g2_o21ai_1 _18394_ (.B1(_11742_),
    .Y(_00651_),
    .A1(_11739_),
    .A2(_11741_));
 sg13g2_nand2_1 _18395_ (.Y(_11743_),
    .A(net730),
    .B(\mem.mem_internal.code_mem[160][2] ));
 sg13g2_nand2_1 _18396_ (.Y(_11744_),
    .A(net1140),
    .B(_11738_));
 sg13g2_o21ai_1 _18397_ (.B1(_11744_),
    .Y(_00652_),
    .A1(net247),
    .A2(_11743_));
 sg13g2_nand2_1 _18398_ (.Y(_11745_),
    .A(net730),
    .B(\mem.mem_internal.code_mem[160][3] ));
 sg13g2_nand2_1 _18399_ (.Y(_11746_),
    .A(net1139),
    .B(_11738_));
 sg13g2_o21ai_1 _18400_ (.B1(_11746_),
    .Y(_00653_),
    .A1(net247),
    .A2(_11745_));
 sg13g2_nand2_1 _18401_ (.Y(_11747_),
    .A(net730),
    .B(\mem.mem_internal.code_mem[160][4] ));
 sg13g2_nand2_1 _18402_ (.Y(_11748_),
    .A(net1138),
    .B(_11738_));
 sg13g2_o21ai_1 _18403_ (.B1(_11748_),
    .Y(_00654_),
    .A1(net247),
    .A2(_11747_));
 sg13g2_nand2_1 _18404_ (.Y(_11749_),
    .A(net730),
    .B(\mem.mem_internal.code_mem[160][5] ));
 sg13g2_nand2_1 _18405_ (.Y(_11750_),
    .A(net1137),
    .B(_11738_));
 sg13g2_o21ai_1 _18406_ (.B1(_11750_),
    .Y(_00655_),
    .A1(net247),
    .A2(_11749_));
 sg13g2_nand2_1 _18407_ (.Y(_11751_),
    .A(net730),
    .B(\mem.mem_internal.code_mem[160][6] ));
 sg13g2_nand2_1 _18408_ (.Y(_11752_),
    .A(net1136),
    .B(_11738_));
 sg13g2_o21ai_1 _18409_ (.B1(_11752_),
    .Y(_00656_),
    .A1(net247),
    .A2(_11751_));
 sg13g2_buf_1 _18410_ (.A(_11665_),
    .X(_11753_));
 sg13g2_nand2_1 _18411_ (.Y(_11754_),
    .A(_11753_),
    .B(\mem.mem_internal.code_mem[160][7] ));
 sg13g2_nand2_1 _18412_ (.Y(_11755_),
    .A(net1135),
    .B(_11738_));
 sg13g2_o21ai_1 _18413_ (.B1(_11755_),
    .Y(_00657_),
    .A1(net247),
    .A2(_11754_));
 sg13g2_nand2_1 _18414_ (.Y(_11756_),
    .A(_11692_),
    .B(\mem.mem_internal.code_mem[161][0] ));
 sg13g2_nor2_1 _18415_ (.A(net528),
    .B(net465),
    .Y(_11757_));
 sg13g2_buf_2 _18416_ (.A(_11757_),
    .X(_11758_));
 sg13g2_buf_1 _18417_ (.A(_11758_),
    .X(_11759_));
 sg13g2_nand2_1 _18418_ (.Y(_11760_),
    .A(net1142),
    .B(net246));
 sg13g2_o21ai_1 _18419_ (.B1(_11760_),
    .Y(_00658_),
    .A1(_11756_),
    .A2(net246));
 sg13g2_nand2_1 _18420_ (.Y(_11761_),
    .A(net729),
    .B(\mem.mem_internal.code_mem[161][1] ));
 sg13g2_nand2_1 _18421_ (.Y(_11762_),
    .A(net1141),
    .B(net246));
 sg13g2_o21ai_1 _18422_ (.B1(_11762_),
    .Y(_00659_),
    .A1(_11759_),
    .A2(_11761_));
 sg13g2_nand2_1 _18423_ (.Y(_11763_),
    .A(net729),
    .B(\mem.mem_internal.code_mem[161][2] ));
 sg13g2_nand2_1 _18424_ (.Y(_11764_),
    .A(net1140),
    .B(_11758_));
 sg13g2_o21ai_1 _18425_ (.B1(_11764_),
    .Y(_00660_),
    .A1(net246),
    .A2(_11763_));
 sg13g2_nand2_1 _18426_ (.Y(_11765_),
    .A(net729),
    .B(\mem.mem_internal.code_mem[161][3] ));
 sg13g2_nand2_1 _18427_ (.Y(_11766_),
    .A(net1139),
    .B(_11758_));
 sg13g2_o21ai_1 _18428_ (.B1(_11766_),
    .Y(_00661_),
    .A1(net246),
    .A2(_11765_));
 sg13g2_nand2_1 _18429_ (.Y(_11767_),
    .A(net729),
    .B(\mem.mem_internal.code_mem[161][4] ));
 sg13g2_nand2_1 _18430_ (.Y(_11768_),
    .A(net1138),
    .B(_11758_));
 sg13g2_o21ai_1 _18431_ (.B1(_11768_),
    .Y(_00662_),
    .A1(net246),
    .A2(_11767_));
 sg13g2_nand2_1 _18432_ (.Y(_11769_),
    .A(net729),
    .B(\mem.mem_internal.code_mem[161][5] ));
 sg13g2_nand2_1 _18433_ (.Y(_11770_),
    .A(net1137),
    .B(_11758_));
 sg13g2_o21ai_1 _18434_ (.B1(_11770_),
    .Y(_00663_),
    .A1(net246),
    .A2(_11769_));
 sg13g2_nand2_1 _18435_ (.Y(_11771_),
    .A(net729),
    .B(\mem.mem_internal.code_mem[161][6] ));
 sg13g2_nand2_1 _18436_ (.Y(_11772_),
    .A(net1136),
    .B(_11758_));
 sg13g2_o21ai_1 _18437_ (.B1(_11772_),
    .Y(_00664_),
    .A1(net246),
    .A2(_11771_));
 sg13g2_nand2_1 _18438_ (.Y(_11773_),
    .A(_11753_),
    .B(\mem.mem_internal.code_mem[161][7] ));
 sg13g2_nand2_1 _18439_ (.Y(_11774_),
    .A(net1135),
    .B(_11758_));
 sg13g2_o21ai_1 _18440_ (.B1(_11774_),
    .Y(_00665_),
    .A1(_11759_),
    .A2(_11773_));
 sg13g2_nand2_1 _18441_ (.Y(_11775_),
    .A(_11692_),
    .B(\mem.mem_internal.code_mem[162][0] ));
 sg13g2_nor2_1 _18442_ (.A(net527),
    .B(_11736_),
    .Y(_11776_));
 sg13g2_buf_2 _18443_ (.A(_11776_),
    .X(_11777_));
 sg13g2_buf_1 _18444_ (.A(_11777_),
    .X(_11778_));
 sg13g2_nand2_1 _18445_ (.Y(_11779_),
    .A(net1142),
    .B(_11778_));
 sg13g2_o21ai_1 _18446_ (.B1(_11779_),
    .Y(_00666_),
    .A1(_11775_),
    .A2(_11778_));
 sg13g2_nand2_1 _18447_ (.Y(_11780_),
    .A(net729),
    .B(\mem.mem_internal.code_mem[162][1] ));
 sg13g2_nand2_1 _18448_ (.Y(_11781_),
    .A(net1141),
    .B(net245));
 sg13g2_o21ai_1 _18449_ (.B1(_11781_),
    .Y(_00667_),
    .A1(net245),
    .A2(_11780_));
 sg13g2_nand2_1 _18450_ (.Y(_11782_),
    .A(net729),
    .B(\mem.mem_internal.code_mem[162][2] ));
 sg13g2_nand2_1 _18451_ (.Y(_11783_),
    .A(net1140),
    .B(_11777_));
 sg13g2_o21ai_1 _18452_ (.B1(_11783_),
    .Y(_00668_),
    .A1(net245),
    .A2(_11782_));
 sg13g2_buf_1 _18453_ (.A(_11665_),
    .X(_11784_));
 sg13g2_nand2_1 _18454_ (.Y(_11785_),
    .A(net728),
    .B(\mem.mem_internal.code_mem[162][3] ));
 sg13g2_nand2_1 _18455_ (.Y(_11786_),
    .A(net1139),
    .B(_11777_));
 sg13g2_o21ai_1 _18456_ (.B1(_11786_),
    .Y(_00669_),
    .A1(net245),
    .A2(_11785_));
 sg13g2_nand2_1 _18457_ (.Y(_11787_),
    .A(net728),
    .B(\mem.mem_internal.code_mem[162][4] ));
 sg13g2_nand2_1 _18458_ (.Y(_11788_),
    .A(net1138),
    .B(_11777_));
 sg13g2_o21ai_1 _18459_ (.B1(_11788_),
    .Y(_00670_),
    .A1(net245),
    .A2(_11787_));
 sg13g2_nand2_1 _18460_ (.Y(_11789_),
    .A(net728),
    .B(\mem.mem_internal.code_mem[162][5] ));
 sg13g2_nand2_1 _18461_ (.Y(_11790_),
    .A(net1137),
    .B(_11777_));
 sg13g2_o21ai_1 _18462_ (.B1(_11790_),
    .Y(_00671_),
    .A1(net245),
    .A2(_11789_));
 sg13g2_nand2_1 _18463_ (.Y(_11791_),
    .A(net728),
    .B(\mem.mem_internal.code_mem[162][6] ));
 sg13g2_nand2_1 _18464_ (.Y(_11792_),
    .A(net1136),
    .B(_11777_));
 sg13g2_o21ai_1 _18465_ (.B1(_11792_),
    .Y(_00672_),
    .A1(net245),
    .A2(_11791_));
 sg13g2_nand2_1 _18466_ (.Y(_11793_),
    .A(net728),
    .B(\mem.mem_internal.code_mem[162][7] ));
 sg13g2_nand2_1 _18467_ (.Y(_11794_),
    .A(net1135),
    .B(_11777_));
 sg13g2_o21ai_1 _18468_ (.B1(_11794_),
    .Y(_00673_),
    .A1(net245),
    .A2(_11793_));
 sg13g2_nand2_1 _18469_ (.Y(_11795_),
    .A(net846),
    .B(\mem.mem_internal.code_mem[163][0] ));
 sg13g2_nor2_1 _18470_ (.A(net526),
    .B(_11736_),
    .Y(_11796_));
 sg13g2_buf_2 _18471_ (.A(_11796_),
    .X(_11797_));
 sg13g2_buf_1 _18472_ (.A(_11797_),
    .X(_11798_));
 sg13g2_buf_1 _18473_ (.A(_11163_),
    .X(_11799_));
 sg13g2_nand2_1 _18474_ (.Y(_11800_),
    .A(_11799_),
    .B(net244));
 sg13g2_o21ai_1 _18475_ (.B1(_11800_),
    .Y(_00674_),
    .A1(_11795_),
    .A2(net244));
 sg13g2_nand2_1 _18476_ (.Y(_11801_),
    .A(_11784_),
    .B(\mem.mem_internal.code_mem[163][1] ));
 sg13g2_buf_1 _18477_ (.A(_11167_),
    .X(_11802_));
 sg13g2_nand2_1 _18478_ (.Y(_11803_),
    .A(_11802_),
    .B(net244));
 sg13g2_o21ai_1 _18479_ (.B1(_11803_),
    .Y(_00675_),
    .A1(net244),
    .A2(_11801_));
 sg13g2_nand2_1 _18480_ (.Y(_11804_),
    .A(net728),
    .B(\mem.mem_internal.code_mem[163][2] ));
 sg13g2_buf_1 _18481_ (.A(_11171_),
    .X(_11805_));
 sg13g2_nand2_1 _18482_ (.Y(_11806_),
    .A(_11805_),
    .B(_11797_));
 sg13g2_o21ai_1 _18483_ (.B1(_11806_),
    .Y(_00676_),
    .A1(_11798_),
    .A2(_11804_));
 sg13g2_nand2_1 _18484_ (.Y(_11807_),
    .A(net728),
    .B(\mem.mem_internal.code_mem[163][3] ));
 sg13g2_buf_1 _18485_ (.A(_11175_),
    .X(_11808_));
 sg13g2_nand2_1 _18486_ (.Y(_11809_),
    .A(_11808_),
    .B(_11797_));
 sg13g2_o21ai_1 _18487_ (.B1(_11809_),
    .Y(_00677_),
    .A1(_11798_),
    .A2(_11807_));
 sg13g2_nand2_1 _18488_ (.Y(_11810_),
    .A(net728),
    .B(\mem.mem_internal.code_mem[163][4] ));
 sg13g2_buf_1 _18489_ (.A(_11179_),
    .X(_11811_));
 sg13g2_nand2_1 _18490_ (.Y(_11812_),
    .A(_11811_),
    .B(_11797_));
 sg13g2_o21ai_1 _18491_ (.B1(_11812_),
    .Y(_00678_),
    .A1(net244),
    .A2(_11810_));
 sg13g2_nand2_1 _18492_ (.Y(_11813_),
    .A(_11784_),
    .B(\mem.mem_internal.code_mem[163][5] ));
 sg13g2_buf_1 _18493_ (.A(_11183_),
    .X(_11814_));
 sg13g2_nand2_1 _18494_ (.Y(_11815_),
    .A(_11814_),
    .B(_11797_));
 sg13g2_o21ai_1 _18495_ (.B1(_11815_),
    .Y(_00679_),
    .A1(net244),
    .A2(_11813_));
 sg13g2_buf_1 _18496_ (.A(_11665_),
    .X(_11816_));
 sg13g2_nand2_1 _18497_ (.Y(_11817_),
    .A(_11816_),
    .B(\mem.mem_internal.code_mem[163][6] ));
 sg13g2_buf_1 _18498_ (.A(_11188_),
    .X(_11818_));
 sg13g2_nand2_1 _18499_ (.Y(_11819_),
    .A(_11818_),
    .B(_11797_));
 sg13g2_o21ai_1 _18500_ (.B1(_11819_),
    .Y(_00680_),
    .A1(net244),
    .A2(_11817_));
 sg13g2_nand2_1 _18501_ (.Y(_11820_),
    .A(_11816_),
    .B(\mem.mem_internal.code_mem[163][7] ));
 sg13g2_buf_1 _18502_ (.A(_11192_),
    .X(_11821_));
 sg13g2_nand2_1 _18503_ (.Y(_11822_),
    .A(_11821_),
    .B(_11797_));
 sg13g2_o21ai_1 _18504_ (.B1(_11822_),
    .Y(_00681_),
    .A1(net244),
    .A2(_11820_));
 sg13g2_nand2_1 _18505_ (.Y(_11823_),
    .A(net846),
    .B(\mem.mem_internal.code_mem[164][0] ));
 sg13g2_nor2_1 _18506_ (.A(net556),
    .B(net465),
    .Y(_11824_));
 sg13g2_buf_2 _18507_ (.A(_11824_),
    .X(_11825_));
 sg13g2_buf_1 _18508_ (.A(_11825_),
    .X(_11826_));
 sg13g2_nand2_1 _18509_ (.Y(_11827_),
    .A(net1134),
    .B(net243));
 sg13g2_o21ai_1 _18510_ (.B1(_11827_),
    .Y(_00682_),
    .A1(_11823_),
    .A2(net243));
 sg13g2_nand2_1 _18511_ (.Y(_11828_),
    .A(net727),
    .B(\mem.mem_internal.code_mem[164][1] ));
 sg13g2_nand2_1 _18512_ (.Y(_11829_),
    .A(net1133),
    .B(net243));
 sg13g2_o21ai_1 _18513_ (.B1(_11829_),
    .Y(_00683_),
    .A1(_11826_),
    .A2(_11828_));
 sg13g2_nand2_1 _18514_ (.Y(_11830_),
    .A(net727),
    .B(\mem.mem_internal.code_mem[164][2] ));
 sg13g2_nand2_1 _18515_ (.Y(_11831_),
    .A(net1132),
    .B(_11825_));
 sg13g2_o21ai_1 _18516_ (.B1(_11831_),
    .Y(_00684_),
    .A1(_11826_),
    .A2(_11830_));
 sg13g2_nand2_1 _18517_ (.Y(_11832_),
    .A(net727),
    .B(\mem.mem_internal.code_mem[164][3] ));
 sg13g2_nand2_1 _18518_ (.Y(_11833_),
    .A(net1131),
    .B(_11825_));
 sg13g2_o21ai_1 _18519_ (.B1(_11833_),
    .Y(_00685_),
    .A1(net243),
    .A2(_11832_));
 sg13g2_nand2_1 _18520_ (.Y(_11834_),
    .A(net727),
    .B(\mem.mem_internal.code_mem[164][4] ));
 sg13g2_nand2_1 _18521_ (.Y(_11835_),
    .A(net1130),
    .B(_11825_));
 sg13g2_o21ai_1 _18522_ (.B1(_11835_),
    .Y(_00686_),
    .A1(net243),
    .A2(_11834_));
 sg13g2_nand2_1 _18523_ (.Y(_11836_),
    .A(net727),
    .B(\mem.mem_internal.code_mem[164][5] ));
 sg13g2_nand2_1 _18524_ (.Y(_11837_),
    .A(net1129),
    .B(_11825_));
 sg13g2_o21ai_1 _18525_ (.B1(_11837_),
    .Y(_00687_),
    .A1(net243),
    .A2(_11836_));
 sg13g2_nand2_1 _18526_ (.Y(_11838_),
    .A(net727),
    .B(\mem.mem_internal.code_mem[164][6] ));
 sg13g2_nand2_1 _18527_ (.Y(_11839_),
    .A(net1128),
    .B(_11825_));
 sg13g2_o21ai_1 _18528_ (.B1(_11839_),
    .Y(_00688_),
    .A1(net243),
    .A2(_11838_));
 sg13g2_nand2_1 _18529_ (.Y(_11840_),
    .A(net727),
    .B(\mem.mem_internal.code_mem[164][7] ));
 sg13g2_nand2_1 _18530_ (.Y(_11841_),
    .A(net1127),
    .B(_11825_));
 sg13g2_o21ai_1 _18531_ (.B1(_11841_),
    .Y(_00689_),
    .A1(net243),
    .A2(_11840_));
 sg13g2_nand2_1 _18532_ (.Y(_11842_),
    .A(net846),
    .B(\mem.mem_internal.code_mem[165][0] ));
 sg13g2_nor2_1 _18533_ (.A(net555),
    .B(net465),
    .Y(_11843_));
 sg13g2_buf_2 _18534_ (.A(_11843_),
    .X(_11844_));
 sg13g2_buf_1 _18535_ (.A(_11844_),
    .X(_11845_));
 sg13g2_nand2_1 _18536_ (.Y(_11846_),
    .A(net1134),
    .B(_11845_));
 sg13g2_o21ai_1 _18537_ (.B1(_11846_),
    .Y(_00690_),
    .A1(_11842_),
    .A2(_11845_));
 sg13g2_nand2_1 _18538_ (.Y(_11847_),
    .A(net727),
    .B(\mem.mem_internal.code_mem[165][1] ));
 sg13g2_nand2_1 _18539_ (.Y(_11848_),
    .A(net1133),
    .B(net242));
 sg13g2_o21ai_1 _18540_ (.B1(_11848_),
    .Y(_00691_),
    .A1(net242),
    .A2(_11847_));
 sg13g2_buf_1 _18541_ (.A(_11665_),
    .X(_11849_));
 sg13g2_nand2_1 _18542_ (.Y(_11850_),
    .A(net726),
    .B(\mem.mem_internal.code_mem[165][2] ));
 sg13g2_nand2_1 _18543_ (.Y(_11851_),
    .A(net1132),
    .B(_11844_));
 sg13g2_o21ai_1 _18544_ (.B1(_11851_),
    .Y(_00692_),
    .A1(net242),
    .A2(_11850_));
 sg13g2_nand2_1 _18545_ (.Y(_11852_),
    .A(net726),
    .B(\mem.mem_internal.code_mem[165][3] ));
 sg13g2_nand2_1 _18546_ (.Y(_11853_),
    .A(net1131),
    .B(_11844_));
 sg13g2_o21ai_1 _18547_ (.B1(_11853_),
    .Y(_00693_),
    .A1(net242),
    .A2(_11852_));
 sg13g2_nand2_1 _18548_ (.Y(_11854_),
    .A(net726),
    .B(\mem.mem_internal.code_mem[165][4] ));
 sg13g2_nand2_1 _18549_ (.Y(_11855_),
    .A(net1130),
    .B(_11844_));
 sg13g2_o21ai_1 _18550_ (.B1(_11855_),
    .Y(_00694_),
    .A1(net242),
    .A2(_11854_));
 sg13g2_nand2_1 _18551_ (.Y(_11856_),
    .A(net726),
    .B(\mem.mem_internal.code_mem[165][5] ));
 sg13g2_nand2_1 _18552_ (.Y(_11857_),
    .A(net1129),
    .B(_11844_));
 sg13g2_o21ai_1 _18553_ (.B1(_11857_),
    .Y(_00695_),
    .A1(net242),
    .A2(_11856_));
 sg13g2_nand2_1 _18554_ (.Y(_11858_),
    .A(net726),
    .B(\mem.mem_internal.code_mem[165][6] ));
 sg13g2_nand2_1 _18555_ (.Y(_11859_),
    .A(net1128),
    .B(_11844_));
 sg13g2_o21ai_1 _18556_ (.B1(_11859_),
    .Y(_00696_),
    .A1(net242),
    .A2(_11858_));
 sg13g2_nand2_1 _18557_ (.Y(_11860_),
    .A(net726),
    .B(\mem.mem_internal.code_mem[165][7] ));
 sg13g2_nand2_1 _18558_ (.Y(_11861_),
    .A(net1127),
    .B(_11844_));
 sg13g2_o21ai_1 _18559_ (.B1(_11861_),
    .Y(_00697_),
    .A1(net242),
    .A2(_11860_));
 sg13g2_nand2_1 _18560_ (.Y(_11862_),
    .A(net846),
    .B(\mem.mem_internal.code_mem[166][0] ));
 sg13g2_nor2_1 _18561_ (.A(net554),
    .B(net465),
    .Y(_11863_));
 sg13g2_buf_2 _18562_ (.A(_11863_),
    .X(_11864_));
 sg13g2_buf_1 _18563_ (.A(_11864_),
    .X(_11865_));
 sg13g2_nand2_1 _18564_ (.Y(_11866_),
    .A(net1134),
    .B(net241));
 sg13g2_o21ai_1 _18565_ (.B1(_11866_),
    .Y(_00698_),
    .A1(_11862_),
    .A2(net241));
 sg13g2_nand2_1 _18566_ (.Y(_11867_),
    .A(net726),
    .B(\mem.mem_internal.code_mem[166][1] ));
 sg13g2_nand2_1 _18567_ (.Y(_11868_),
    .A(net1133),
    .B(net241));
 sg13g2_o21ai_1 _18568_ (.B1(_11868_),
    .Y(_00699_),
    .A1(_11865_),
    .A2(_11867_));
 sg13g2_nand2_1 _18569_ (.Y(_11869_),
    .A(net726),
    .B(\mem.mem_internal.code_mem[166][2] ));
 sg13g2_nand2_1 _18570_ (.Y(_11870_),
    .A(net1132),
    .B(_11864_));
 sg13g2_o21ai_1 _18571_ (.B1(_11870_),
    .Y(_00700_),
    .A1(_11865_),
    .A2(_11869_));
 sg13g2_nand2_1 _18572_ (.Y(_11871_),
    .A(_11849_),
    .B(\mem.mem_internal.code_mem[166][3] ));
 sg13g2_nand2_1 _18573_ (.Y(_11872_),
    .A(net1131),
    .B(_11864_));
 sg13g2_o21ai_1 _18574_ (.B1(_11872_),
    .Y(_00701_),
    .A1(net241),
    .A2(_11871_));
 sg13g2_nand2_1 _18575_ (.Y(_11873_),
    .A(_11849_),
    .B(\mem.mem_internal.code_mem[166][4] ));
 sg13g2_nand2_1 _18576_ (.Y(_11874_),
    .A(net1130),
    .B(_11864_));
 sg13g2_o21ai_1 _18577_ (.B1(_11874_),
    .Y(_00702_),
    .A1(net241),
    .A2(_11873_));
 sg13g2_buf_2 _18578_ (.A(net1276),
    .X(_11875_));
 sg13g2_buf_1 _18579_ (.A(_11875_),
    .X(_11876_));
 sg13g2_buf_1 _18580_ (.A(_11876_),
    .X(_11877_));
 sg13g2_nand2_1 _18581_ (.Y(_11878_),
    .A(net725),
    .B(\mem.mem_internal.code_mem[166][5] ));
 sg13g2_nand2_1 _18582_ (.Y(_11879_),
    .A(net1129),
    .B(_11864_));
 sg13g2_o21ai_1 _18583_ (.B1(_11879_),
    .Y(_00703_),
    .A1(net241),
    .A2(_11878_));
 sg13g2_nand2_1 _18584_ (.Y(_11880_),
    .A(net725),
    .B(\mem.mem_internal.code_mem[166][6] ));
 sg13g2_nand2_1 _18585_ (.Y(_11881_),
    .A(net1128),
    .B(_11864_));
 sg13g2_o21ai_1 _18586_ (.B1(_11881_),
    .Y(_00704_),
    .A1(net241),
    .A2(_11880_));
 sg13g2_nand2_1 _18587_ (.Y(_11882_),
    .A(_11877_),
    .B(\mem.mem_internal.code_mem[166][7] ));
 sg13g2_nand2_1 _18588_ (.Y(_11883_),
    .A(net1127),
    .B(_11864_));
 sg13g2_o21ai_1 _18589_ (.B1(_11883_),
    .Y(_00705_),
    .A1(net241),
    .A2(_11882_));
 sg13g2_nand2_1 _18590_ (.Y(_11884_),
    .A(net846),
    .B(\mem.mem_internal.code_mem[167][0] ));
 sg13g2_nor2_1 _18591_ (.A(net553),
    .B(net465),
    .Y(_11885_));
 sg13g2_buf_2 _18592_ (.A(_11885_),
    .X(_11886_));
 sg13g2_buf_1 _18593_ (.A(_11886_),
    .X(_11887_));
 sg13g2_nand2_1 _18594_ (.Y(_11888_),
    .A(net1134),
    .B(_11887_));
 sg13g2_o21ai_1 _18595_ (.B1(_11888_),
    .Y(_00706_),
    .A1(_11884_),
    .A2(_11887_));
 sg13g2_nand2_1 _18596_ (.Y(_11889_),
    .A(_11877_),
    .B(\mem.mem_internal.code_mem[167][1] ));
 sg13g2_nand2_1 _18597_ (.Y(_11890_),
    .A(net1133),
    .B(net240));
 sg13g2_o21ai_1 _18598_ (.B1(_11890_),
    .Y(_00707_),
    .A1(net240),
    .A2(_11889_));
 sg13g2_nand2_1 _18599_ (.Y(_11891_),
    .A(net725),
    .B(\mem.mem_internal.code_mem[167][2] ));
 sg13g2_nand2_1 _18600_ (.Y(_11892_),
    .A(net1132),
    .B(_11886_));
 sg13g2_o21ai_1 _18601_ (.B1(_11892_),
    .Y(_00708_),
    .A1(net240),
    .A2(_11891_));
 sg13g2_nand2_1 _18602_ (.Y(_11893_),
    .A(net725),
    .B(\mem.mem_internal.code_mem[167][3] ));
 sg13g2_nand2_1 _18603_ (.Y(_11894_),
    .A(net1131),
    .B(_11886_));
 sg13g2_o21ai_1 _18604_ (.B1(_11894_),
    .Y(_00709_),
    .A1(net240),
    .A2(_11893_));
 sg13g2_nand2_1 _18605_ (.Y(_11895_),
    .A(net725),
    .B(\mem.mem_internal.code_mem[167][4] ));
 sg13g2_nand2_1 _18606_ (.Y(_11896_),
    .A(net1130),
    .B(_11886_));
 sg13g2_o21ai_1 _18607_ (.B1(_11896_),
    .Y(_00710_),
    .A1(net240),
    .A2(_11895_));
 sg13g2_nand2_1 _18608_ (.Y(_11897_),
    .A(net725),
    .B(\mem.mem_internal.code_mem[167][5] ));
 sg13g2_nand2_1 _18609_ (.Y(_11898_),
    .A(net1129),
    .B(_11886_));
 sg13g2_o21ai_1 _18610_ (.B1(_11898_),
    .Y(_00711_),
    .A1(net240),
    .A2(_11897_));
 sg13g2_nand2_1 _18611_ (.Y(_11899_),
    .A(net725),
    .B(\mem.mem_internal.code_mem[167][6] ));
 sg13g2_nand2_1 _18612_ (.Y(_11900_),
    .A(net1128),
    .B(_11886_));
 sg13g2_o21ai_1 _18613_ (.B1(_11900_),
    .Y(_00712_),
    .A1(net240),
    .A2(_11899_));
 sg13g2_nand2_1 _18614_ (.Y(_11901_),
    .A(net725),
    .B(\mem.mem_internal.code_mem[167][7] ));
 sg13g2_nand2_1 _18615_ (.Y(_11902_),
    .A(net1127),
    .B(_11886_));
 sg13g2_o21ai_1 _18616_ (.B1(_11902_),
    .Y(_00713_),
    .A1(net240),
    .A2(_11901_));
 sg13g2_buf_1 _18617_ (.A(_11058_),
    .X(_11903_));
 sg13g2_nand2_1 _18618_ (.Y(_11904_),
    .A(net845),
    .B(\mem.mem_internal.code_mem[168][0] ));
 sg13g2_nor2_1 _18619_ (.A(net552),
    .B(net465),
    .Y(_11905_));
 sg13g2_buf_2 _18620_ (.A(_11905_),
    .X(_11906_));
 sg13g2_buf_1 _18621_ (.A(_11906_),
    .X(_11907_));
 sg13g2_nand2_1 _18622_ (.Y(_11908_),
    .A(net1134),
    .B(net239));
 sg13g2_o21ai_1 _18623_ (.B1(_11908_),
    .Y(_00714_),
    .A1(_11904_),
    .A2(net239));
 sg13g2_buf_1 _18624_ (.A(_11876_),
    .X(_11909_));
 sg13g2_nand2_1 _18625_ (.Y(_11910_),
    .A(net724),
    .B(\mem.mem_internal.code_mem[168][1] ));
 sg13g2_nand2_1 _18626_ (.Y(_11911_),
    .A(net1133),
    .B(net239));
 sg13g2_o21ai_1 _18627_ (.B1(_11911_),
    .Y(_00715_),
    .A1(net239),
    .A2(_11910_));
 sg13g2_nand2_1 _18628_ (.Y(_11912_),
    .A(net724),
    .B(\mem.mem_internal.code_mem[168][2] ));
 sg13g2_nand2_1 _18629_ (.Y(_11913_),
    .A(net1132),
    .B(_11906_));
 sg13g2_o21ai_1 _18630_ (.B1(_11913_),
    .Y(_00716_),
    .A1(net239),
    .A2(_11912_));
 sg13g2_nand2_1 _18631_ (.Y(_11914_),
    .A(net724),
    .B(\mem.mem_internal.code_mem[168][3] ));
 sg13g2_nand2_1 _18632_ (.Y(_11915_),
    .A(net1131),
    .B(_11906_));
 sg13g2_o21ai_1 _18633_ (.B1(_11915_),
    .Y(_00717_),
    .A1(net239),
    .A2(_11914_));
 sg13g2_nand2_1 _18634_ (.Y(_11916_),
    .A(net724),
    .B(\mem.mem_internal.code_mem[168][4] ));
 sg13g2_nand2_1 _18635_ (.Y(_11917_),
    .A(net1130),
    .B(_11906_));
 sg13g2_o21ai_1 _18636_ (.B1(_11917_),
    .Y(_00718_),
    .A1(_11907_),
    .A2(_11916_));
 sg13g2_nand2_1 _18637_ (.Y(_11918_),
    .A(net724),
    .B(\mem.mem_internal.code_mem[168][5] ));
 sg13g2_nand2_1 _18638_ (.Y(_11919_),
    .A(net1129),
    .B(_11906_));
 sg13g2_o21ai_1 _18639_ (.B1(_11919_),
    .Y(_00719_),
    .A1(net239),
    .A2(_11918_));
 sg13g2_nand2_1 _18640_ (.Y(_11920_),
    .A(net724),
    .B(\mem.mem_internal.code_mem[168][6] ));
 sg13g2_nand2_1 _18641_ (.Y(_11921_),
    .A(net1128),
    .B(_11906_));
 sg13g2_o21ai_1 _18642_ (.B1(_11921_),
    .Y(_00720_),
    .A1(net239),
    .A2(_11920_));
 sg13g2_nand2_1 _18643_ (.Y(_11922_),
    .A(_11909_),
    .B(\mem.mem_internal.code_mem[168][7] ));
 sg13g2_nand2_1 _18644_ (.Y(_11923_),
    .A(net1127),
    .B(_11906_));
 sg13g2_o21ai_1 _18645_ (.B1(_11923_),
    .Y(_00721_),
    .A1(_11907_),
    .A2(_11922_));
 sg13g2_nand2_1 _18646_ (.Y(_11924_),
    .A(net845),
    .B(\mem.mem_internal.code_mem[169][0] ));
 sg13g2_nor2_1 _18647_ (.A(net551),
    .B(net465),
    .Y(_11925_));
 sg13g2_buf_2 _18648_ (.A(_11925_),
    .X(_11926_));
 sg13g2_buf_1 _18649_ (.A(_11926_),
    .X(_11927_));
 sg13g2_nand2_1 _18650_ (.Y(_11928_),
    .A(net1134),
    .B(net238));
 sg13g2_o21ai_1 _18651_ (.B1(_11928_),
    .Y(_00722_),
    .A1(_11924_),
    .A2(net238));
 sg13g2_nand2_1 _18652_ (.Y(_11929_),
    .A(net724),
    .B(\mem.mem_internal.code_mem[169][1] ));
 sg13g2_nand2_1 _18653_ (.Y(_11930_),
    .A(net1133),
    .B(net238));
 sg13g2_o21ai_1 _18654_ (.B1(_11930_),
    .Y(_00723_),
    .A1(net238),
    .A2(_11929_));
 sg13g2_nand2_1 _18655_ (.Y(_11931_),
    .A(_11909_),
    .B(\mem.mem_internal.code_mem[169][2] ));
 sg13g2_nand2_1 _18656_ (.Y(_11932_),
    .A(net1132),
    .B(_11926_));
 sg13g2_o21ai_1 _18657_ (.B1(_11932_),
    .Y(_00724_),
    .A1(net238),
    .A2(_11931_));
 sg13g2_nand2_1 _18658_ (.Y(_11933_),
    .A(net724),
    .B(\mem.mem_internal.code_mem[169][3] ));
 sg13g2_nand2_1 _18659_ (.Y(_11934_),
    .A(net1131),
    .B(_11926_));
 sg13g2_o21ai_1 _18660_ (.B1(_11934_),
    .Y(_00725_),
    .A1(net238),
    .A2(_11933_));
 sg13g2_buf_1 _18661_ (.A(_11876_),
    .X(_11935_));
 sg13g2_nand2_1 _18662_ (.Y(_11936_),
    .A(net723),
    .B(\mem.mem_internal.code_mem[169][4] ));
 sg13g2_nand2_1 _18663_ (.Y(_11937_),
    .A(net1130),
    .B(_11926_));
 sg13g2_o21ai_1 _18664_ (.B1(_11937_),
    .Y(_00726_),
    .A1(net238),
    .A2(_11936_));
 sg13g2_nand2_1 _18665_ (.Y(_11938_),
    .A(net723),
    .B(\mem.mem_internal.code_mem[169][5] ));
 sg13g2_nand2_1 _18666_ (.Y(_11939_),
    .A(net1129),
    .B(_11926_));
 sg13g2_o21ai_1 _18667_ (.B1(_11939_),
    .Y(_00727_),
    .A1(_11927_),
    .A2(_11938_));
 sg13g2_nand2_1 _18668_ (.Y(_11940_),
    .A(net723),
    .B(\mem.mem_internal.code_mem[169][6] ));
 sg13g2_nand2_1 _18669_ (.Y(_11941_),
    .A(net1128),
    .B(_11926_));
 sg13g2_o21ai_1 _18670_ (.B1(_11941_),
    .Y(_00728_),
    .A1(_11927_),
    .A2(_11940_));
 sg13g2_nand2_1 _18671_ (.Y(_11942_),
    .A(net723),
    .B(\mem.mem_internal.code_mem[169][7] ));
 sg13g2_nand2_1 _18672_ (.Y(_11943_),
    .A(net1127),
    .B(_11926_));
 sg13g2_o21ai_1 _18673_ (.B1(_11943_),
    .Y(_00729_),
    .A1(net238),
    .A2(_11942_));
 sg13g2_nand2_1 _18674_ (.Y(_11944_),
    .A(_11903_),
    .B(\mem.mem_internal.code_mem[16][0] ));
 sg13g2_nand2_1 _18675_ (.Y(_11945_),
    .A(_10234_),
    .B(_11355_));
 sg13g2_buf_2 _18676_ (.A(_11945_),
    .X(_11946_));
 sg13g2_buf_2 _18677_ (.A(_11946_),
    .X(_11947_));
 sg13g2_nor2_1 _18678_ (.A(net529),
    .B(net464),
    .Y(_11948_));
 sg13g2_buf_2 _18679_ (.A(_11948_),
    .X(_11949_));
 sg13g2_buf_1 _18680_ (.A(_11949_),
    .X(_11950_));
 sg13g2_nand2_1 _18681_ (.Y(_11951_),
    .A(_11799_),
    .B(net237));
 sg13g2_o21ai_1 _18682_ (.B1(_11951_),
    .Y(_00730_),
    .A1(_11944_),
    .A2(_11950_));
 sg13g2_nand2_1 _18683_ (.Y(_11952_),
    .A(net723),
    .B(\mem.mem_internal.code_mem[16][1] ));
 sg13g2_nand2_1 _18684_ (.Y(_11953_),
    .A(_11802_),
    .B(net237));
 sg13g2_o21ai_1 _18685_ (.B1(_11953_),
    .Y(_00731_),
    .A1(net237),
    .A2(_11952_));
 sg13g2_nand2_1 _18686_ (.Y(_11954_),
    .A(net723),
    .B(\mem.mem_internal.code_mem[16][2] ));
 sg13g2_nand2_1 _18687_ (.Y(_11955_),
    .A(_11805_),
    .B(_11949_));
 sg13g2_o21ai_1 _18688_ (.B1(_11955_),
    .Y(_00732_),
    .A1(net237),
    .A2(_11954_));
 sg13g2_nand2_1 _18689_ (.Y(_11956_),
    .A(net723),
    .B(\mem.mem_internal.code_mem[16][3] ));
 sg13g2_nand2_1 _18690_ (.Y(_11957_),
    .A(_11808_),
    .B(_11949_));
 sg13g2_o21ai_1 _18691_ (.B1(_11957_),
    .Y(_00733_),
    .A1(net237),
    .A2(_11956_));
 sg13g2_nand2_1 _18692_ (.Y(_11958_),
    .A(net723),
    .B(\mem.mem_internal.code_mem[16][4] ));
 sg13g2_nand2_1 _18693_ (.Y(_11959_),
    .A(_11811_),
    .B(_11949_));
 sg13g2_o21ai_1 _18694_ (.B1(_11959_),
    .Y(_00734_),
    .A1(net237),
    .A2(_11958_));
 sg13g2_nand2_1 _18695_ (.Y(_11960_),
    .A(_11935_),
    .B(\mem.mem_internal.code_mem[16][5] ));
 sg13g2_nand2_1 _18696_ (.Y(_11961_),
    .A(_11814_),
    .B(_11949_));
 sg13g2_o21ai_1 _18697_ (.B1(_11961_),
    .Y(_00735_),
    .A1(_11950_),
    .A2(_11960_));
 sg13g2_nand2_1 _18698_ (.Y(_11962_),
    .A(_11935_),
    .B(\mem.mem_internal.code_mem[16][6] ));
 sg13g2_nand2_1 _18699_ (.Y(_11963_),
    .A(_11818_),
    .B(_11949_));
 sg13g2_o21ai_1 _18700_ (.B1(_11963_),
    .Y(_00736_),
    .A1(net237),
    .A2(_11962_));
 sg13g2_buf_1 _18701_ (.A(_11876_),
    .X(_11964_));
 sg13g2_nand2_1 _18702_ (.Y(_11965_),
    .A(_11964_),
    .B(\mem.mem_internal.code_mem[16][7] ));
 sg13g2_nand2_1 _18703_ (.Y(_11966_),
    .A(_11821_),
    .B(_11949_));
 sg13g2_o21ai_1 _18704_ (.B1(_11966_),
    .Y(_00737_),
    .A1(net237),
    .A2(_11965_));
 sg13g2_nand2_1 _18705_ (.Y(_11967_),
    .A(net845),
    .B(\mem.mem_internal.code_mem[170][0] ));
 sg13g2_nor2_1 _18706_ (.A(net550),
    .B(_11735_),
    .Y(_11968_));
 sg13g2_buf_2 _18707_ (.A(_11968_),
    .X(_11969_));
 sg13g2_buf_1 _18708_ (.A(_11969_),
    .X(_11970_));
 sg13g2_nand2_1 _18709_ (.Y(_11971_),
    .A(net1134),
    .B(_11970_));
 sg13g2_o21ai_1 _18710_ (.B1(_11971_),
    .Y(_00738_),
    .A1(_11967_),
    .A2(_11970_));
 sg13g2_nand2_1 _18711_ (.Y(_11972_),
    .A(net722),
    .B(\mem.mem_internal.code_mem[170][1] ));
 sg13g2_nand2_1 _18712_ (.Y(_11973_),
    .A(net1133),
    .B(net378));
 sg13g2_o21ai_1 _18713_ (.B1(_11973_),
    .Y(_00739_),
    .A1(net378),
    .A2(_11972_));
 sg13g2_nand2_1 _18714_ (.Y(_11974_),
    .A(net722),
    .B(\mem.mem_internal.code_mem[170][2] ));
 sg13g2_nand2_1 _18715_ (.Y(_11975_),
    .A(net1132),
    .B(_11969_));
 sg13g2_o21ai_1 _18716_ (.B1(_11975_),
    .Y(_00740_),
    .A1(net378),
    .A2(_11974_));
 sg13g2_nand2_1 _18717_ (.Y(_11976_),
    .A(net722),
    .B(\mem.mem_internal.code_mem[170][3] ));
 sg13g2_nand2_1 _18718_ (.Y(_11977_),
    .A(net1131),
    .B(_11969_));
 sg13g2_o21ai_1 _18719_ (.B1(_11977_),
    .Y(_00741_),
    .A1(net378),
    .A2(_11976_));
 sg13g2_nand2_1 _18720_ (.Y(_11978_),
    .A(net722),
    .B(\mem.mem_internal.code_mem[170][4] ));
 sg13g2_nand2_1 _18721_ (.Y(_11979_),
    .A(net1130),
    .B(_11969_));
 sg13g2_o21ai_1 _18722_ (.B1(_11979_),
    .Y(_00742_),
    .A1(net378),
    .A2(_11978_));
 sg13g2_nand2_1 _18723_ (.Y(_11980_),
    .A(_11964_),
    .B(\mem.mem_internal.code_mem[170][5] ));
 sg13g2_nand2_1 _18724_ (.Y(_11981_),
    .A(net1129),
    .B(_11969_));
 sg13g2_o21ai_1 _18725_ (.B1(_11981_),
    .Y(_00743_),
    .A1(net378),
    .A2(_11980_));
 sg13g2_nand2_1 _18726_ (.Y(_11982_),
    .A(net722),
    .B(\mem.mem_internal.code_mem[170][6] ));
 sg13g2_nand2_1 _18727_ (.Y(_11983_),
    .A(net1128),
    .B(_11969_));
 sg13g2_o21ai_1 _18728_ (.B1(_11983_),
    .Y(_00744_),
    .A1(net378),
    .A2(_11982_));
 sg13g2_nand2_1 _18729_ (.Y(_11984_),
    .A(net722),
    .B(\mem.mem_internal.code_mem[170][7] ));
 sg13g2_nand2_1 _18730_ (.Y(_11985_),
    .A(net1127),
    .B(_11969_));
 sg13g2_o21ai_1 _18731_ (.B1(_11985_),
    .Y(_00745_),
    .A1(net378),
    .A2(_11984_));
 sg13g2_nand2_1 _18732_ (.Y(_11986_),
    .A(net845),
    .B(\mem.mem_internal.code_mem[171][0] ));
 sg13g2_nor2_1 _18733_ (.A(net549),
    .B(_11735_),
    .Y(_11987_));
 sg13g2_buf_2 _18734_ (.A(_11987_),
    .X(_11988_));
 sg13g2_buf_1 _18735_ (.A(_11988_),
    .X(_11989_));
 sg13g2_nand2_1 _18736_ (.Y(_11990_),
    .A(net1134),
    .B(net377));
 sg13g2_o21ai_1 _18737_ (.B1(_11990_),
    .Y(_00746_),
    .A1(_11986_),
    .A2(net377));
 sg13g2_nand2_1 _18738_ (.Y(_11991_),
    .A(net722),
    .B(\mem.mem_internal.code_mem[171][1] ));
 sg13g2_nand2_1 _18739_ (.Y(_11992_),
    .A(net1133),
    .B(net377));
 sg13g2_o21ai_1 _18740_ (.B1(_11992_),
    .Y(_00747_),
    .A1(net377),
    .A2(_11991_));
 sg13g2_nand2_1 _18741_ (.Y(_11993_),
    .A(net722),
    .B(\mem.mem_internal.code_mem[171][2] ));
 sg13g2_nand2_1 _18742_ (.Y(_11994_),
    .A(net1132),
    .B(_11988_));
 sg13g2_o21ai_1 _18743_ (.B1(_11994_),
    .Y(_00748_),
    .A1(net377),
    .A2(_11993_));
 sg13g2_buf_1 _18744_ (.A(_11876_),
    .X(_11995_));
 sg13g2_nand2_1 _18745_ (.Y(_11996_),
    .A(net721),
    .B(\mem.mem_internal.code_mem[171][3] ));
 sg13g2_nand2_1 _18746_ (.Y(_11997_),
    .A(net1131),
    .B(_11988_));
 sg13g2_o21ai_1 _18747_ (.B1(_11997_),
    .Y(_00749_),
    .A1(net377),
    .A2(_11996_));
 sg13g2_nand2_1 _18748_ (.Y(_11998_),
    .A(_11995_),
    .B(\mem.mem_internal.code_mem[171][4] ));
 sg13g2_nand2_1 _18749_ (.Y(_11999_),
    .A(net1130),
    .B(_11988_));
 sg13g2_o21ai_1 _18750_ (.B1(_11999_),
    .Y(_00750_),
    .A1(_11989_),
    .A2(_11998_));
 sg13g2_nand2_1 _18751_ (.Y(_12000_),
    .A(_11995_),
    .B(\mem.mem_internal.code_mem[171][5] ));
 sg13g2_nand2_1 _18752_ (.Y(_12001_),
    .A(net1129),
    .B(_11988_));
 sg13g2_o21ai_1 _18753_ (.B1(_12001_),
    .Y(_00751_),
    .A1(_11989_),
    .A2(_12000_));
 sg13g2_nand2_1 _18754_ (.Y(_12002_),
    .A(net721),
    .B(\mem.mem_internal.code_mem[171][6] ));
 sg13g2_nand2_1 _18755_ (.Y(_12003_),
    .A(net1128),
    .B(_11988_));
 sg13g2_o21ai_1 _18756_ (.B1(_12003_),
    .Y(_00752_),
    .A1(net377),
    .A2(_12002_));
 sg13g2_nand2_1 _18757_ (.Y(_12004_),
    .A(net721),
    .B(\mem.mem_internal.code_mem[171][7] ));
 sg13g2_nand2_1 _18758_ (.Y(_12005_),
    .A(net1127),
    .B(_11988_));
 sg13g2_o21ai_1 _18759_ (.B1(_12005_),
    .Y(_00753_),
    .A1(net377),
    .A2(_12004_));
 sg13g2_nand2_1 _18760_ (.Y(_12006_),
    .A(net845),
    .B(\mem.mem_internal.code_mem[172][0] ));
 sg13g2_nor2_1 _18761_ (.A(net773),
    .B(_11735_),
    .Y(_12007_));
 sg13g2_buf_2 _18762_ (.A(_12007_),
    .X(_12008_));
 sg13g2_buf_1 _18763_ (.A(_12008_),
    .X(_12009_));
 sg13g2_buf_1 _18764_ (.A(_11163_),
    .X(_12010_));
 sg13g2_nand2_1 _18765_ (.Y(_12011_),
    .A(net1126),
    .B(net376));
 sg13g2_o21ai_1 _18766_ (.B1(_12011_),
    .Y(_00754_),
    .A1(_12006_),
    .A2(_12009_));
 sg13g2_nand2_1 _18767_ (.Y(_12012_),
    .A(net721),
    .B(\mem.mem_internal.code_mem[172][1] ));
 sg13g2_buf_1 _18768_ (.A(_11167_),
    .X(_12013_));
 sg13g2_nand2_1 _18769_ (.Y(_12014_),
    .A(net1125),
    .B(net376));
 sg13g2_o21ai_1 _18770_ (.B1(_12014_),
    .Y(_00755_),
    .A1(net376),
    .A2(_12012_));
 sg13g2_nand2_1 _18771_ (.Y(_12015_),
    .A(net721),
    .B(\mem.mem_internal.code_mem[172][2] ));
 sg13g2_buf_1 _18772_ (.A(_11171_),
    .X(_12016_));
 sg13g2_nand2_1 _18773_ (.Y(_12017_),
    .A(net1124),
    .B(_12008_));
 sg13g2_o21ai_1 _18774_ (.B1(_12017_),
    .Y(_00756_),
    .A1(net376),
    .A2(_12015_));
 sg13g2_nand2_1 _18775_ (.Y(_12018_),
    .A(net721),
    .B(\mem.mem_internal.code_mem[172][3] ));
 sg13g2_buf_1 _18776_ (.A(_11175_),
    .X(_12019_));
 sg13g2_nand2_1 _18777_ (.Y(_12020_),
    .A(net1123),
    .B(_12008_));
 sg13g2_o21ai_1 _18778_ (.B1(_12020_),
    .Y(_00757_),
    .A1(net376),
    .A2(_12018_));
 sg13g2_nand2_1 _18779_ (.Y(_12021_),
    .A(net721),
    .B(\mem.mem_internal.code_mem[172][4] ));
 sg13g2_buf_1 _18780_ (.A(_11179_),
    .X(_12022_));
 sg13g2_nand2_1 _18781_ (.Y(_12023_),
    .A(net1122),
    .B(_12008_));
 sg13g2_o21ai_1 _18782_ (.B1(_12023_),
    .Y(_00758_),
    .A1(net376),
    .A2(_12021_));
 sg13g2_nand2_1 _18783_ (.Y(_12024_),
    .A(net721),
    .B(\mem.mem_internal.code_mem[172][5] ));
 sg13g2_buf_1 _18784_ (.A(_11183_),
    .X(_12025_));
 sg13g2_nand2_1 _18785_ (.Y(_12026_),
    .A(net1121),
    .B(_12008_));
 sg13g2_o21ai_1 _18786_ (.B1(_12026_),
    .Y(_00759_),
    .A1(net376),
    .A2(_12024_));
 sg13g2_buf_1 _18787_ (.A(_11876_),
    .X(_12027_));
 sg13g2_nand2_1 _18788_ (.Y(_12028_),
    .A(net720),
    .B(\mem.mem_internal.code_mem[172][6] ));
 sg13g2_buf_1 _18789_ (.A(_11188_),
    .X(_12029_));
 sg13g2_nand2_1 _18790_ (.Y(_12030_),
    .A(net1120),
    .B(_12008_));
 sg13g2_o21ai_1 _18791_ (.B1(_12030_),
    .Y(_00760_),
    .A1(net376),
    .A2(_12028_));
 sg13g2_nand2_1 _18792_ (.Y(_12031_),
    .A(net720),
    .B(\mem.mem_internal.code_mem[172][7] ));
 sg13g2_buf_1 _18793_ (.A(_11192_),
    .X(_12032_));
 sg13g2_nand2_1 _18794_ (.Y(_12033_),
    .A(net1119),
    .B(_12008_));
 sg13g2_o21ai_1 _18795_ (.B1(_12033_),
    .Y(_00761_),
    .A1(_12009_),
    .A2(_12031_));
 sg13g2_nand2_1 _18796_ (.Y(_12034_),
    .A(net845),
    .B(\mem.mem_internal.code_mem[173][0] ));
 sg13g2_nor2_1 _18797_ (.A(net548),
    .B(_11735_),
    .Y(_12035_));
 sg13g2_buf_2 _18798_ (.A(_12035_),
    .X(_12036_));
 sg13g2_buf_1 _18799_ (.A(_12036_),
    .X(_12037_));
 sg13g2_nand2_1 _18800_ (.Y(_12038_),
    .A(net1126),
    .B(net375));
 sg13g2_o21ai_1 _18801_ (.B1(_12038_),
    .Y(_00762_),
    .A1(_12034_),
    .A2(net375));
 sg13g2_nand2_1 _18802_ (.Y(_12039_),
    .A(_12027_),
    .B(\mem.mem_internal.code_mem[173][1] ));
 sg13g2_nand2_1 _18803_ (.Y(_12040_),
    .A(net1125),
    .B(net375));
 sg13g2_o21ai_1 _18804_ (.B1(_12040_),
    .Y(_00763_),
    .A1(_12037_),
    .A2(_12039_));
 sg13g2_nand2_1 _18805_ (.Y(_12041_),
    .A(_12027_),
    .B(\mem.mem_internal.code_mem[173][2] ));
 sg13g2_nand2_1 _18806_ (.Y(_12042_),
    .A(net1124),
    .B(_12036_));
 sg13g2_o21ai_1 _18807_ (.B1(_12042_),
    .Y(_00764_),
    .A1(_12037_),
    .A2(_12041_));
 sg13g2_nand2_1 _18808_ (.Y(_12043_),
    .A(net720),
    .B(\mem.mem_internal.code_mem[173][3] ));
 sg13g2_nand2_1 _18809_ (.Y(_12044_),
    .A(net1123),
    .B(_12036_));
 sg13g2_o21ai_1 _18810_ (.B1(_12044_),
    .Y(_00765_),
    .A1(net375),
    .A2(_12043_));
 sg13g2_nand2_1 _18811_ (.Y(_12045_),
    .A(net720),
    .B(\mem.mem_internal.code_mem[173][4] ));
 sg13g2_nand2_1 _18812_ (.Y(_12046_),
    .A(net1122),
    .B(_12036_));
 sg13g2_o21ai_1 _18813_ (.B1(_12046_),
    .Y(_00766_),
    .A1(net375),
    .A2(_12045_));
 sg13g2_nand2_1 _18814_ (.Y(_12047_),
    .A(net720),
    .B(\mem.mem_internal.code_mem[173][5] ));
 sg13g2_nand2_1 _18815_ (.Y(_12048_),
    .A(net1121),
    .B(_12036_));
 sg13g2_o21ai_1 _18816_ (.B1(_12048_),
    .Y(_00767_),
    .A1(net375),
    .A2(_12047_));
 sg13g2_nand2_1 _18817_ (.Y(_12049_),
    .A(net720),
    .B(\mem.mem_internal.code_mem[173][6] ));
 sg13g2_nand2_1 _18818_ (.Y(_12050_),
    .A(net1120),
    .B(_12036_));
 sg13g2_o21ai_1 _18819_ (.B1(_12050_),
    .Y(_00768_),
    .A1(net375),
    .A2(_12049_));
 sg13g2_nand2_1 _18820_ (.Y(_12051_),
    .A(net720),
    .B(\mem.mem_internal.code_mem[173][7] ));
 sg13g2_nand2_1 _18821_ (.Y(_12052_),
    .A(net1119),
    .B(_12036_));
 sg13g2_o21ai_1 _18822_ (.B1(_12052_),
    .Y(_00769_),
    .A1(net375),
    .A2(_12051_));
 sg13g2_nand2_1 _18823_ (.Y(_12053_),
    .A(net845),
    .B(\mem.mem_internal.code_mem[174][0] ));
 sg13g2_nor2_1 _18824_ (.A(net547),
    .B(_11735_),
    .Y(_12054_));
 sg13g2_buf_2 _18825_ (.A(_12054_),
    .X(_12055_));
 sg13g2_buf_1 _18826_ (.A(_12055_),
    .X(_12056_));
 sg13g2_nand2_1 _18827_ (.Y(_12057_),
    .A(net1126),
    .B(net374));
 sg13g2_o21ai_1 _18828_ (.B1(_12057_),
    .Y(_00770_),
    .A1(_12053_),
    .A2(net374));
 sg13g2_nand2_1 _18829_ (.Y(_12058_),
    .A(net720),
    .B(\mem.mem_internal.code_mem[174][1] ));
 sg13g2_nand2_1 _18830_ (.Y(_12059_),
    .A(net1125),
    .B(net374));
 sg13g2_o21ai_1 _18831_ (.B1(_12059_),
    .Y(_00771_),
    .A1(net374),
    .A2(_12058_));
 sg13g2_buf_1 _18832_ (.A(_11876_),
    .X(_12060_));
 sg13g2_nand2_1 _18833_ (.Y(_12061_),
    .A(net719),
    .B(\mem.mem_internal.code_mem[174][2] ));
 sg13g2_nand2_1 _18834_ (.Y(_12062_),
    .A(net1124),
    .B(_12055_));
 sg13g2_o21ai_1 _18835_ (.B1(_12062_),
    .Y(_00772_),
    .A1(_12056_),
    .A2(_12061_));
 sg13g2_nand2_1 _18836_ (.Y(_12063_),
    .A(net719),
    .B(\mem.mem_internal.code_mem[174][3] ));
 sg13g2_nand2_1 _18837_ (.Y(_12064_),
    .A(net1123),
    .B(_12055_));
 sg13g2_o21ai_1 _18838_ (.B1(_12064_),
    .Y(_00773_),
    .A1(_12056_),
    .A2(_12063_));
 sg13g2_nand2_1 _18839_ (.Y(_12065_),
    .A(net719),
    .B(\mem.mem_internal.code_mem[174][4] ));
 sg13g2_nand2_1 _18840_ (.Y(_12066_),
    .A(net1122),
    .B(_12055_));
 sg13g2_o21ai_1 _18841_ (.B1(_12066_),
    .Y(_00774_),
    .A1(net374),
    .A2(_12065_));
 sg13g2_nand2_1 _18842_ (.Y(_12067_),
    .A(net719),
    .B(\mem.mem_internal.code_mem[174][5] ));
 sg13g2_nand2_1 _18843_ (.Y(_12068_),
    .A(net1121),
    .B(_12055_));
 sg13g2_o21ai_1 _18844_ (.B1(_12068_),
    .Y(_00775_),
    .A1(net374),
    .A2(_12067_));
 sg13g2_nand2_1 _18845_ (.Y(_12069_),
    .A(net719),
    .B(\mem.mem_internal.code_mem[174][6] ));
 sg13g2_nand2_1 _18846_ (.Y(_12070_),
    .A(_12029_),
    .B(_12055_));
 sg13g2_o21ai_1 _18847_ (.B1(_12070_),
    .Y(_00776_),
    .A1(net374),
    .A2(_12069_));
 sg13g2_nand2_1 _18848_ (.Y(_12071_),
    .A(net719),
    .B(\mem.mem_internal.code_mem[174][7] ));
 sg13g2_nand2_1 _18849_ (.Y(_12072_),
    .A(net1119),
    .B(_12055_));
 sg13g2_o21ai_1 _18850_ (.B1(_12072_),
    .Y(_00777_),
    .A1(net374),
    .A2(_12071_));
 sg13g2_nand2_1 _18851_ (.Y(_12073_),
    .A(net845),
    .B(\mem.mem_internal.code_mem[175][0] ));
 sg13g2_nor2_1 _18852_ (.A(net770),
    .B(_11735_),
    .Y(_12074_));
 sg13g2_buf_2 _18853_ (.A(_12074_),
    .X(_12075_));
 sg13g2_buf_1 _18854_ (.A(_12075_),
    .X(_12076_));
 sg13g2_nand2_1 _18855_ (.Y(_12077_),
    .A(net1126),
    .B(net373));
 sg13g2_o21ai_1 _18856_ (.B1(_12077_),
    .Y(_00778_),
    .A1(_12073_),
    .A2(net373));
 sg13g2_nand2_1 _18857_ (.Y(_12078_),
    .A(net719),
    .B(\mem.mem_internal.code_mem[175][1] ));
 sg13g2_nand2_1 _18858_ (.Y(_12079_),
    .A(net1125),
    .B(net373));
 sg13g2_o21ai_1 _18859_ (.B1(_12079_),
    .Y(_00779_),
    .A1(net373),
    .A2(_12078_));
 sg13g2_nand2_1 _18860_ (.Y(_12080_),
    .A(_12060_),
    .B(\mem.mem_internal.code_mem[175][2] ));
 sg13g2_nand2_1 _18861_ (.Y(_12081_),
    .A(net1124),
    .B(_12075_));
 sg13g2_o21ai_1 _18862_ (.B1(_12081_),
    .Y(_00780_),
    .A1(_12076_),
    .A2(_12080_));
 sg13g2_nand2_1 _18863_ (.Y(_12082_),
    .A(_12060_),
    .B(\mem.mem_internal.code_mem[175][3] ));
 sg13g2_nand2_1 _18864_ (.Y(_12083_),
    .A(net1123),
    .B(_12075_));
 sg13g2_o21ai_1 _18865_ (.B1(_12083_),
    .Y(_00781_),
    .A1(_12076_),
    .A2(_12082_));
 sg13g2_nand2_1 _18866_ (.Y(_12084_),
    .A(net719),
    .B(\mem.mem_internal.code_mem[175][4] ));
 sg13g2_nand2_1 _18867_ (.Y(_12085_),
    .A(net1122),
    .B(_12075_));
 sg13g2_o21ai_1 _18868_ (.B1(_12085_),
    .Y(_00782_),
    .A1(net373),
    .A2(_12084_));
 sg13g2_buf_1 _18869_ (.A(_11875_),
    .X(_12086_));
 sg13g2_buf_1 _18870_ (.A(_12086_),
    .X(_12087_));
 sg13g2_nand2_1 _18871_ (.Y(_12088_),
    .A(net718),
    .B(\mem.mem_internal.code_mem[175][5] ));
 sg13g2_nand2_1 _18872_ (.Y(_12089_),
    .A(net1121),
    .B(_12075_));
 sg13g2_o21ai_1 _18873_ (.B1(_12089_),
    .Y(_00783_),
    .A1(net373),
    .A2(_12088_));
 sg13g2_nand2_1 _18874_ (.Y(_12090_),
    .A(net718),
    .B(\mem.mem_internal.code_mem[175][6] ));
 sg13g2_nand2_1 _18875_ (.Y(_12091_),
    .A(net1120),
    .B(_12075_));
 sg13g2_o21ai_1 _18876_ (.B1(_12091_),
    .Y(_00784_),
    .A1(net373),
    .A2(_12090_));
 sg13g2_nand2_1 _18877_ (.Y(_12092_),
    .A(net718),
    .B(\mem.mem_internal.code_mem[175][7] ));
 sg13g2_nand2_1 _18878_ (.Y(_12093_),
    .A(_12032_),
    .B(_12075_));
 sg13g2_o21ai_1 _18879_ (.B1(_12093_),
    .Y(_00785_),
    .A1(net373),
    .A2(_12092_));
 sg13g2_nand2_1 _18880_ (.Y(_12094_),
    .A(_10607_),
    .B(_10976_));
 sg13g2_buf_2 _18881_ (.A(_12094_),
    .X(_12095_));
 sg13g2_buf_1 _18882_ (.A(_12095_),
    .X(_12096_));
 sg13g2_nor2_1 _18883_ (.A(net529),
    .B(net463),
    .Y(_12097_));
 sg13g2_buf_2 _18884_ (.A(_12097_),
    .X(_12098_));
 sg13g2_buf_1 _18885_ (.A(_12098_),
    .X(_12099_));
 sg13g2_nand2_1 _18886_ (.Y(_12100_),
    .A(_12087_),
    .B(\mem.mem_internal.code_mem[176][0] ));
 sg13g2_nand2_1 _18887_ (.Y(_12101_),
    .A(net1126),
    .B(net236));
 sg13g2_o21ai_1 _18888_ (.B1(_12101_),
    .Y(_00786_),
    .A1(net236),
    .A2(_12100_));
 sg13g2_nand2_1 _18889_ (.Y(_12102_),
    .A(_12087_),
    .B(\mem.mem_internal.code_mem[176][1] ));
 sg13g2_nand2_1 _18890_ (.Y(_12103_),
    .A(net1125),
    .B(_12099_));
 sg13g2_o21ai_1 _18891_ (.B1(_12103_),
    .Y(_00787_),
    .A1(_12099_),
    .A2(_12102_));
 sg13g2_nand2_1 _18892_ (.Y(_12104_),
    .A(net718),
    .B(\mem.mem_internal.code_mem[176][2] ));
 sg13g2_nand2_1 _18893_ (.Y(_12105_),
    .A(net1124),
    .B(_12098_));
 sg13g2_o21ai_1 _18894_ (.B1(_12105_),
    .Y(_00788_),
    .A1(net236),
    .A2(_12104_));
 sg13g2_nand2_1 _18895_ (.Y(_12106_),
    .A(net718),
    .B(\mem.mem_internal.code_mem[176][3] ));
 sg13g2_nand2_1 _18896_ (.Y(_12107_),
    .A(net1123),
    .B(_12098_));
 sg13g2_o21ai_1 _18897_ (.B1(_12107_),
    .Y(_00789_),
    .A1(net236),
    .A2(_12106_));
 sg13g2_nand2_1 _18898_ (.Y(_12108_),
    .A(net718),
    .B(\mem.mem_internal.code_mem[176][4] ));
 sg13g2_nand2_1 _18899_ (.Y(_12109_),
    .A(net1122),
    .B(_12098_));
 sg13g2_o21ai_1 _18900_ (.B1(_12109_),
    .Y(_00790_),
    .A1(net236),
    .A2(_12108_));
 sg13g2_nand2_1 _18901_ (.Y(_12110_),
    .A(net718),
    .B(\mem.mem_internal.code_mem[176][5] ));
 sg13g2_nand2_1 _18902_ (.Y(_12111_),
    .A(net1121),
    .B(_12098_));
 sg13g2_o21ai_1 _18903_ (.B1(_12111_),
    .Y(_00791_),
    .A1(net236),
    .A2(_12110_));
 sg13g2_nand2_1 _18904_ (.Y(_12112_),
    .A(net718),
    .B(\mem.mem_internal.code_mem[176][6] ));
 sg13g2_nand2_1 _18905_ (.Y(_12113_),
    .A(net1120),
    .B(_12098_));
 sg13g2_o21ai_1 _18906_ (.B1(_12113_),
    .Y(_00792_),
    .A1(net236),
    .A2(_12112_));
 sg13g2_buf_1 _18907_ (.A(_12086_),
    .X(_12114_));
 sg13g2_nand2_1 _18908_ (.Y(_12115_),
    .A(net717),
    .B(\mem.mem_internal.code_mem[176][7] ));
 sg13g2_nand2_1 _18909_ (.Y(_12116_),
    .A(net1119),
    .B(_12098_));
 sg13g2_o21ai_1 _18910_ (.B1(_12116_),
    .Y(_00793_),
    .A1(net236),
    .A2(_12115_));
 sg13g2_nor2_1 _18911_ (.A(net528),
    .B(net463),
    .Y(_12117_));
 sg13g2_buf_2 _18912_ (.A(_12117_),
    .X(_12118_));
 sg13g2_buf_1 _18913_ (.A(_12118_),
    .X(_12119_));
 sg13g2_nand2_1 _18914_ (.Y(_12120_),
    .A(_12114_),
    .B(\mem.mem_internal.code_mem[177][0] ));
 sg13g2_nand2_1 _18915_ (.Y(_12121_),
    .A(net1126),
    .B(net235));
 sg13g2_o21ai_1 _18916_ (.B1(_12121_),
    .Y(_00794_),
    .A1(net235),
    .A2(_12120_));
 sg13g2_nand2_1 _18917_ (.Y(_12122_),
    .A(net717),
    .B(\mem.mem_internal.code_mem[177][1] ));
 sg13g2_nand2_1 _18918_ (.Y(_12123_),
    .A(net1125),
    .B(_12119_));
 sg13g2_o21ai_1 _18919_ (.B1(_12123_),
    .Y(_00795_),
    .A1(_12119_),
    .A2(_12122_));
 sg13g2_nand2_1 _18920_ (.Y(_12124_),
    .A(net717),
    .B(\mem.mem_internal.code_mem[177][2] ));
 sg13g2_nand2_1 _18921_ (.Y(_12125_),
    .A(net1124),
    .B(_12118_));
 sg13g2_o21ai_1 _18922_ (.B1(_12125_),
    .Y(_00796_),
    .A1(net235),
    .A2(_12124_));
 sg13g2_nand2_1 _18923_ (.Y(_12126_),
    .A(net717),
    .B(\mem.mem_internal.code_mem[177][3] ));
 sg13g2_nand2_1 _18924_ (.Y(_12127_),
    .A(net1123),
    .B(_12118_));
 sg13g2_o21ai_1 _18925_ (.B1(_12127_),
    .Y(_00797_),
    .A1(net235),
    .A2(_12126_));
 sg13g2_nand2_1 _18926_ (.Y(_12128_),
    .A(net717),
    .B(\mem.mem_internal.code_mem[177][4] ));
 sg13g2_nand2_1 _18927_ (.Y(_12129_),
    .A(net1122),
    .B(_12118_));
 sg13g2_o21ai_1 _18928_ (.B1(_12129_),
    .Y(_00798_),
    .A1(net235),
    .A2(_12128_));
 sg13g2_nand2_1 _18929_ (.Y(_12130_),
    .A(net717),
    .B(\mem.mem_internal.code_mem[177][5] ));
 sg13g2_nand2_1 _18930_ (.Y(_12131_),
    .A(net1121),
    .B(_12118_));
 sg13g2_o21ai_1 _18931_ (.B1(_12131_),
    .Y(_00799_),
    .A1(net235),
    .A2(_12130_));
 sg13g2_nand2_1 _18932_ (.Y(_12132_),
    .A(net717),
    .B(\mem.mem_internal.code_mem[177][6] ));
 sg13g2_nand2_1 _18933_ (.Y(_12133_),
    .A(net1120),
    .B(_12118_));
 sg13g2_o21ai_1 _18934_ (.B1(_12133_),
    .Y(_00800_),
    .A1(net235),
    .A2(_12132_));
 sg13g2_nand2_1 _18935_ (.Y(_12134_),
    .A(net717),
    .B(\mem.mem_internal.code_mem[177][7] ));
 sg13g2_nand2_1 _18936_ (.Y(_12135_),
    .A(net1119),
    .B(_12118_));
 sg13g2_o21ai_1 _18937_ (.B1(_12135_),
    .Y(_00801_),
    .A1(net235),
    .A2(_12134_));
 sg13g2_nor2_1 _18938_ (.A(net527),
    .B(net463),
    .Y(_12136_));
 sg13g2_buf_2 _18939_ (.A(_12136_),
    .X(_12137_));
 sg13g2_buf_1 _18940_ (.A(_12137_),
    .X(_12138_));
 sg13g2_nand2_1 _18941_ (.Y(_12139_),
    .A(_12114_),
    .B(\mem.mem_internal.code_mem[178][0] ));
 sg13g2_nand2_1 _18942_ (.Y(_12140_),
    .A(net1126),
    .B(net234));
 sg13g2_o21ai_1 _18943_ (.B1(_12140_),
    .Y(_00802_),
    .A1(_12138_),
    .A2(_12139_));
 sg13g2_buf_1 _18944_ (.A(_12086_),
    .X(_12141_));
 sg13g2_nand2_1 _18945_ (.Y(_12142_),
    .A(net716),
    .B(\mem.mem_internal.code_mem[178][1] ));
 sg13g2_nand2_1 _18946_ (.Y(_12143_),
    .A(net1125),
    .B(net234));
 sg13g2_o21ai_1 _18947_ (.B1(_12143_),
    .Y(_00803_),
    .A1(net234),
    .A2(_12142_));
 sg13g2_nand2_1 _18948_ (.Y(_12144_),
    .A(net716),
    .B(\mem.mem_internal.code_mem[178][2] ));
 sg13g2_nand2_1 _18949_ (.Y(_12145_),
    .A(net1124),
    .B(_12137_));
 sg13g2_o21ai_1 _18950_ (.B1(_12145_),
    .Y(_00804_),
    .A1(net234),
    .A2(_12144_));
 sg13g2_nand2_1 _18951_ (.Y(_12146_),
    .A(net716),
    .B(\mem.mem_internal.code_mem[178][3] ));
 sg13g2_nand2_1 _18952_ (.Y(_12147_),
    .A(net1123),
    .B(_12137_));
 sg13g2_o21ai_1 _18953_ (.B1(_12147_),
    .Y(_00805_),
    .A1(net234),
    .A2(_12146_));
 sg13g2_nand2_1 _18954_ (.Y(_12148_),
    .A(net716),
    .B(\mem.mem_internal.code_mem[178][4] ));
 sg13g2_nand2_1 _18955_ (.Y(_12149_),
    .A(net1122),
    .B(_12137_));
 sg13g2_o21ai_1 _18956_ (.B1(_12149_),
    .Y(_00806_),
    .A1(net234),
    .A2(_12148_));
 sg13g2_nand2_1 _18957_ (.Y(_12150_),
    .A(net716),
    .B(\mem.mem_internal.code_mem[178][5] ));
 sg13g2_nand2_1 _18958_ (.Y(_12151_),
    .A(net1121),
    .B(_12137_));
 sg13g2_o21ai_1 _18959_ (.B1(_12151_),
    .Y(_00807_),
    .A1(net234),
    .A2(_12150_));
 sg13g2_nand2_1 _18960_ (.Y(_12152_),
    .A(net716),
    .B(\mem.mem_internal.code_mem[178][6] ));
 sg13g2_nand2_1 _18961_ (.Y(_12153_),
    .A(net1120),
    .B(_12137_));
 sg13g2_o21ai_1 _18962_ (.B1(_12153_),
    .Y(_00808_),
    .A1(net234),
    .A2(_12152_));
 sg13g2_nand2_1 _18963_ (.Y(_12154_),
    .A(net716),
    .B(\mem.mem_internal.code_mem[178][7] ));
 sg13g2_nand2_1 _18964_ (.Y(_12155_),
    .A(net1119),
    .B(_12137_));
 sg13g2_o21ai_1 _18965_ (.B1(_12155_),
    .Y(_00809_),
    .A1(_12138_),
    .A2(_12154_));
 sg13g2_nor2_1 _18966_ (.A(net526),
    .B(net463),
    .Y(_12156_));
 sg13g2_buf_2 _18967_ (.A(_12156_),
    .X(_12157_));
 sg13g2_buf_1 _18968_ (.A(_12157_),
    .X(_12158_));
 sg13g2_nand2_1 _18969_ (.Y(_12159_),
    .A(_12141_),
    .B(\mem.mem_internal.code_mem[179][0] ));
 sg13g2_nand2_1 _18970_ (.Y(_12160_),
    .A(net1126),
    .B(net233));
 sg13g2_o21ai_1 _18971_ (.B1(_12160_),
    .Y(_00810_),
    .A1(net233),
    .A2(_12159_));
 sg13g2_nand2_1 _18972_ (.Y(_12161_),
    .A(_12141_),
    .B(\mem.mem_internal.code_mem[179][1] ));
 sg13g2_nand2_1 _18973_ (.Y(_12162_),
    .A(net1125),
    .B(_12158_));
 sg13g2_o21ai_1 _18974_ (.B1(_12162_),
    .Y(_00811_),
    .A1(_12158_),
    .A2(_12161_));
 sg13g2_nand2_1 _18975_ (.Y(_12163_),
    .A(net716),
    .B(\mem.mem_internal.code_mem[179][2] ));
 sg13g2_nand2_1 _18976_ (.Y(_12164_),
    .A(net1124),
    .B(_12157_));
 sg13g2_o21ai_1 _18977_ (.B1(_12164_),
    .Y(_00812_),
    .A1(net233),
    .A2(_12163_));
 sg13g2_buf_1 _18978_ (.A(_12086_),
    .X(_12165_));
 sg13g2_nand2_1 _18979_ (.Y(_12166_),
    .A(net715),
    .B(\mem.mem_internal.code_mem[179][3] ));
 sg13g2_nand2_1 _18980_ (.Y(_12167_),
    .A(net1123),
    .B(_12157_));
 sg13g2_o21ai_1 _18981_ (.B1(_12167_),
    .Y(_00813_),
    .A1(net233),
    .A2(_12166_));
 sg13g2_nand2_1 _18982_ (.Y(_12168_),
    .A(net715),
    .B(\mem.mem_internal.code_mem[179][4] ));
 sg13g2_nand2_1 _18983_ (.Y(_12169_),
    .A(net1122),
    .B(_12157_));
 sg13g2_o21ai_1 _18984_ (.B1(_12169_),
    .Y(_00814_),
    .A1(net233),
    .A2(_12168_));
 sg13g2_nand2_1 _18985_ (.Y(_12170_),
    .A(net715),
    .B(\mem.mem_internal.code_mem[179][5] ));
 sg13g2_nand2_1 _18986_ (.Y(_12171_),
    .A(net1121),
    .B(_12157_));
 sg13g2_o21ai_1 _18987_ (.B1(_12171_),
    .Y(_00815_),
    .A1(net233),
    .A2(_12170_));
 sg13g2_nand2_1 _18988_ (.Y(_12172_),
    .A(net715),
    .B(\mem.mem_internal.code_mem[179][6] ));
 sg13g2_nand2_1 _18989_ (.Y(_12173_),
    .A(net1120),
    .B(_12157_));
 sg13g2_o21ai_1 _18990_ (.B1(_12173_),
    .Y(_00816_),
    .A1(net233),
    .A2(_12172_));
 sg13g2_nand2_1 _18991_ (.Y(_12174_),
    .A(net715),
    .B(\mem.mem_internal.code_mem[179][7] ));
 sg13g2_nand2_1 _18992_ (.Y(_12175_),
    .A(net1119),
    .B(_12157_));
 sg13g2_o21ai_1 _18993_ (.B1(_12175_),
    .Y(_00817_),
    .A1(net233),
    .A2(_12174_));
 sg13g2_nand2_1 _18994_ (.Y(_12176_),
    .A(_11903_),
    .B(\mem.mem_internal.code_mem[17][0] ));
 sg13g2_nor2_1 _18995_ (.A(net528),
    .B(net464),
    .Y(_12177_));
 sg13g2_buf_2 _18996_ (.A(_12177_),
    .X(_12178_));
 sg13g2_buf_1 _18997_ (.A(_12178_),
    .X(_12179_));
 sg13g2_nand2_1 _18998_ (.Y(_12180_),
    .A(_12010_),
    .B(net232));
 sg13g2_o21ai_1 _18999_ (.B1(_12180_),
    .Y(_00818_),
    .A1(_12176_),
    .A2(net232));
 sg13g2_nand2_1 _19000_ (.Y(_12181_),
    .A(net715),
    .B(\mem.mem_internal.code_mem[17][1] ));
 sg13g2_nand2_1 _19001_ (.Y(_12182_),
    .A(_12013_),
    .B(_12179_));
 sg13g2_o21ai_1 _19002_ (.B1(_12182_),
    .Y(_00819_),
    .A1(_12179_),
    .A2(_12181_));
 sg13g2_nand2_1 _19003_ (.Y(_12183_),
    .A(net715),
    .B(\mem.mem_internal.code_mem[17][2] ));
 sg13g2_nand2_1 _19004_ (.Y(_12184_),
    .A(_12016_),
    .B(_12178_));
 sg13g2_o21ai_1 _19005_ (.B1(_12184_),
    .Y(_00820_),
    .A1(net232),
    .A2(_12183_));
 sg13g2_nand2_1 _19006_ (.Y(_12185_),
    .A(net715),
    .B(\mem.mem_internal.code_mem[17][3] ));
 sg13g2_nand2_1 _19007_ (.Y(_12186_),
    .A(_12019_),
    .B(_12178_));
 sg13g2_o21ai_1 _19008_ (.B1(_12186_),
    .Y(_00821_),
    .A1(net232),
    .A2(_12185_));
 sg13g2_nand2_1 _19009_ (.Y(_12187_),
    .A(_12165_),
    .B(\mem.mem_internal.code_mem[17][4] ));
 sg13g2_nand2_1 _19010_ (.Y(_12188_),
    .A(_12022_),
    .B(_12178_));
 sg13g2_o21ai_1 _19011_ (.B1(_12188_),
    .Y(_00822_),
    .A1(net232),
    .A2(_12187_));
 sg13g2_nand2_1 _19012_ (.Y(_12189_),
    .A(_12165_),
    .B(\mem.mem_internal.code_mem[17][5] ));
 sg13g2_nand2_1 _19013_ (.Y(_12190_),
    .A(_12025_),
    .B(_12178_));
 sg13g2_o21ai_1 _19014_ (.B1(_12190_),
    .Y(_00823_),
    .A1(net232),
    .A2(_12189_));
 sg13g2_buf_1 _19015_ (.A(_12086_),
    .X(_12191_));
 sg13g2_nand2_1 _19016_ (.Y(_12192_),
    .A(_12191_),
    .B(\mem.mem_internal.code_mem[17][6] ));
 sg13g2_nand2_1 _19017_ (.Y(_12193_),
    .A(_12029_),
    .B(_12178_));
 sg13g2_o21ai_1 _19018_ (.B1(_12193_),
    .Y(_00824_),
    .A1(net232),
    .A2(_12192_));
 sg13g2_nand2_1 _19019_ (.Y(_12194_),
    .A(_12191_),
    .B(\mem.mem_internal.code_mem[17][7] ));
 sg13g2_nand2_1 _19020_ (.Y(_12195_),
    .A(_12032_),
    .B(_12178_));
 sg13g2_o21ai_1 _19021_ (.B1(_12195_),
    .Y(_00825_),
    .A1(net232),
    .A2(_12194_));
 sg13g2_nor2_1 _19022_ (.A(net556),
    .B(net463),
    .Y(_12196_));
 sg13g2_buf_2 _19023_ (.A(_12196_),
    .X(_12197_));
 sg13g2_buf_1 _19024_ (.A(_12197_),
    .X(_12198_));
 sg13g2_nand2_1 _19025_ (.Y(_12199_),
    .A(net714),
    .B(\mem.mem_internal.code_mem[180][0] ));
 sg13g2_nand2_1 _19026_ (.Y(_12200_),
    .A(_12010_),
    .B(_12198_));
 sg13g2_o21ai_1 _19027_ (.B1(_12200_),
    .Y(_00826_),
    .A1(_12198_),
    .A2(_12199_));
 sg13g2_nand2_1 _19028_ (.Y(_12201_),
    .A(net714),
    .B(\mem.mem_internal.code_mem[180][1] ));
 sg13g2_nand2_1 _19029_ (.Y(_12202_),
    .A(_12013_),
    .B(net231));
 sg13g2_o21ai_1 _19030_ (.B1(_12202_),
    .Y(_00827_),
    .A1(net231),
    .A2(_12201_));
 sg13g2_nand2_1 _19031_ (.Y(_12203_),
    .A(net714),
    .B(\mem.mem_internal.code_mem[180][2] ));
 sg13g2_nand2_1 _19032_ (.Y(_12204_),
    .A(_12016_),
    .B(_12197_));
 sg13g2_o21ai_1 _19033_ (.B1(_12204_),
    .Y(_00828_),
    .A1(net231),
    .A2(_12203_));
 sg13g2_nand2_1 _19034_ (.Y(_12205_),
    .A(net714),
    .B(\mem.mem_internal.code_mem[180][3] ));
 sg13g2_nand2_1 _19035_ (.Y(_12206_),
    .A(_12019_),
    .B(_12197_));
 sg13g2_o21ai_1 _19036_ (.B1(_12206_),
    .Y(_00829_),
    .A1(net231),
    .A2(_12205_));
 sg13g2_nand2_1 _19037_ (.Y(_12207_),
    .A(net714),
    .B(\mem.mem_internal.code_mem[180][4] ));
 sg13g2_nand2_1 _19038_ (.Y(_12208_),
    .A(_12022_),
    .B(_12197_));
 sg13g2_o21ai_1 _19039_ (.B1(_12208_),
    .Y(_00830_),
    .A1(net231),
    .A2(_12207_));
 sg13g2_nand2_1 _19040_ (.Y(_12209_),
    .A(net714),
    .B(\mem.mem_internal.code_mem[180][5] ));
 sg13g2_nand2_1 _19041_ (.Y(_12210_),
    .A(_12025_),
    .B(_12197_));
 sg13g2_o21ai_1 _19042_ (.B1(_12210_),
    .Y(_00831_),
    .A1(net231),
    .A2(_12209_));
 sg13g2_nand2_1 _19043_ (.Y(_12211_),
    .A(net714),
    .B(\mem.mem_internal.code_mem[180][6] ));
 sg13g2_nand2_1 _19044_ (.Y(_12212_),
    .A(net1120),
    .B(_12197_));
 sg13g2_o21ai_1 _19045_ (.B1(_12212_),
    .Y(_00832_),
    .A1(net231),
    .A2(_12211_));
 sg13g2_nand2_1 _19046_ (.Y(_12213_),
    .A(net714),
    .B(\mem.mem_internal.code_mem[180][7] ));
 sg13g2_nand2_1 _19047_ (.Y(_12214_),
    .A(net1119),
    .B(_12197_));
 sg13g2_o21ai_1 _19048_ (.B1(_12214_),
    .Y(_00833_),
    .A1(net231),
    .A2(_12213_));
 sg13g2_nor2_1 _19049_ (.A(net555),
    .B(_12096_),
    .Y(_12215_));
 sg13g2_buf_2 _19050_ (.A(_12215_),
    .X(_12216_));
 sg13g2_buf_1 _19051_ (.A(_12216_),
    .X(_12217_));
 sg13g2_buf_1 _19052_ (.A(_12086_),
    .X(_12218_));
 sg13g2_nand2_1 _19053_ (.Y(_12219_),
    .A(net713),
    .B(\mem.mem_internal.code_mem[181][0] ));
 sg13g2_buf_1 _19054_ (.A(_11163_),
    .X(_12220_));
 sg13g2_nand2_1 _19055_ (.Y(_12221_),
    .A(net1118),
    .B(net230));
 sg13g2_o21ai_1 _19056_ (.B1(_12221_),
    .Y(_00834_),
    .A1(net230),
    .A2(_12219_));
 sg13g2_nand2_1 _19057_ (.Y(_12222_),
    .A(net713),
    .B(\mem.mem_internal.code_mem[181][1] ));
 sg13g2_buf_1 _19058_ (.A(_11167_),
    .X(_12223_));
 sg13g2_nand2_1 _19059_ (.Y(_12224_),
    .A(net1117),
    .B(net230));
 sg13g2_o21ai_1 _19060_ (.B1(_12224_),
    .Y(_00835_),
    .A1(_12217_),
    .A2(_12222_));
 sg13g2_nand2_1 _19061_ (.Y(_12225_),
    .A(_12218_),
    .B(\mem.mem_internal.code_mem[181][2] ));
 sg13g2_buf_1 _19062_ (.A(_11171_),
    .X(_12226_));
 sg13g2_nand2_1 _19063_ (.Y(_12227_),
    .A(net1116),
    .B(_12216_));
 sg13g2_o21ai_1 _19064_ (.B1(_12227_),
    .Y(_00836_),
    .A1(net230),
    .A2(_12225_));
 sg13g2_nand2_1 _19065_ (.Y(_12228_),
    .A(_12218_),
    .B(\mem.mem_internal.code_mem[181][3] ));
 sg13g2_buf_1 _19066_ (.A(_11175_),
    .X(_12229_));
 sg13g2_nand2_1 _19067_ (.Y(_12230_),
    .A(net1115),
    .B(_12216_));
 sg13g2_o21ai_1 _19068_ (.B1(_12230_),
    .Y(_00837_),
    .A1(net230),
    .A2(_12228_));
 sg13g2_nand2_1 _19069_ (.Y(_12231_),
    .A(net713),
    .B(\mem.mem_internal.code_mem[181][4] ));
 sg13g2_buf_1 _19070_ (.A(_11179_),
    .X(_12232_));
 sg13g2_nand2_1 _19071_ (.Y(_12233_),
    .A(net1114),
    .B(_12216_));
 sg13g2_o21ai_1 _19072_ (.B1(_12233_),
    .Y(_00838_),
    .A1(_12217_),
    .A2(_12231_));
 sg13g2_nand2_1 _19073_ (.Y(_12234_),
    .A(net713),
    .B(\mem.mem_internal.code_mem[181][5] ));
 sg13g2_buf_1 _19074_ (.A(_11183_),
    .X(_12235_));
 sg13g2_nand2_1 _19075_ (.Y(_12236_),
    .A(net1113),
    .B(_12216_));
 sg13g2_o21ai_1 _19076_ (.B1(_12236_),
    .Y(_00839_),
    .A1(net230),
    .A2(_12234_));
 sg13g2_nand2_1 _19077_ (.Y(_12237_),
    .A(net713),
    .B(\mem.mem_internal.code_mem[181][6] ));
 sg13g2_buf_1 _19078_ (.A(_11188_),
    .X(_12238_));
 sg13g2_nand2_1 _19079_ (.Y(_12239_),
    .A(net1112),
    .B(_12216_));
 sg13g2_o21ai_1 _19080_ (.B1(_12239_),
    .Y(_00840_),
    .A1(net230),
    .A2(_12237_));
 sg13g2_nand2_1 _19081_ (.Y(_12240_),
    .A(net713),
    .B(\mem.mem_internal.code_mem[181][7] ));
 sg13g2_buf_1 _19082_ (.A(_11192_),
    .X(_12241_));
 sg13g2_nand2_1 _19083_ (.Y(_12242_),
    .A(net1111),
    .B(_12216_));
 sg13g2_o21ai_1 _19084_ (.B1(_12242_),
    .Y(_00841_),
    .A1(net230),
    .A2(_12240_));
 sg13g2_nor2_1 _19085_ (.A(net554),
    .B(_12096_),
    .Y(_12243_));
 sg13g2_buf_2 _19086_ (.A(_12243_),
    .X(_12244_));
 sg13g2_buf_1 _19087_ (.A(_12244_),
    .X(_12245_));
 sg13g2_nand2_1 _19088_ (.Y(_12246_),
    .A(net713),
    .B(\mem.mem_internal.code_mem[182][0] ));
 sg13g2_nand2_1 _19089_ (.Y(_12247_),
    .A(net1118),
    .B(net229));
 sg13g2_o21ai_1 _19090_ (.B1(_12247_),
    .Y(_00842_),
    .A1(net229),
    .A2(_12246_));
 sg13g2_nand2_1 _19091_ (.Y(_12248_),
    .A(net713),
    .B(\mem.mem_internal.code_mem[182][1] ));
 sg13g2_nand2_1 _19092_ (.Y(_12249_),
    .A(net1117),
    .B(net229));
 sg13g2_o21ai_1 _19093_ (.B1(_12249_),
    .Y(_00843_),
    .A1(_12245_),
    .A2(_12248_));
 sg13g2_buf_1 _19094_ (.A(_12086_),
    .X(_12250_));
 sg13g2_nand2_1 _19095_ (.Y(_12251_),
    .A(net712),
    .B(\mem.mem_internal.code_mem[182][2] ));
 sg13g2_nand2_1 _19096_ (.Y(_12252_),
    .A(net1116),
    .B(_12244_));
 sg13g2_o21ai_1 _19097_ (.B1(_12252_),
    .Y(_00844_),
    .A1(net229),
    .A2(_12251_));
 sg13g2_nand2_1 _19098_ (.Y(_12253_),
    .A(net712),
    .B(\mem.mem_internal.code_mem[182][3] ));
 sg13g2_nand2_1 _19099_ (.Y(_12254_),
    .A(net1115),
    .B(_12244_));
 sg13g2_o21ai_1 _19100_ (.B1(_12254_),
    .Y(_00845_),
    .A1(net229),
    .A2(_12253_));
 sg13g2_nand2_1 _19101_ (.Y(_12255_),
    .A(_12250_),
    .B(\mem.mem_internal.code_mem[182][4] ));
 sg13g2_nand2_1 _19102_ (.Y(_12256_),
    .A(net1114),
    .B(_12244_));
 sg13g2_o21ai_1 _19103_ (.B1(_12256_),
    .Y(_00846_),
    .A1(_12245_),
    .A2(_12255_));
 sg13g2_nand2_1 _19104_ (.Y(_12257_),
    .A(net712),
    .B(\mem.mem_internal.code_mem[182][5] ));
 sg13g2_nand2_1 _19105_ (.Y(_12258_),
    .A(net1113),
    .B(_12244_));
 sg13g2_o21ai_1 _19106_ (.B1(_12258_),
    .Y(_00847_),
    .A1(net229),
    .A2(_12257_));
 sg13g2_nand2_1 _19107_ (.Y(_12259_),
    .A(net712),
    .B(\mem.mem_internal.code_mem[182][6] ));
 sg13g2_nand2_1 _19108_ (.Y(_12260_),
    .A(net1112),
    .B(_12244_));
 sg13g2_o21ai_1 _19109_ (.B1(_12260_),
    .Y(_00848_),
    .A1(net229),
    .A2(_12259_));
 sg13g2_nand2_1 _19110_ (.Y(_12261_),
    .A(net712),
    .B(\mem.mem_internal.code_mem[182][7] ));
 sg13g2_nand2_1 _19111_ (.Y(_12262_),
    .A(net1111),
    .B(_12244_));
 sg13g2_o21ai_1 _19112_ (.B1(_12262_),
    .Y(_00849_),
    .A1(net229),
    .A2(_12261_));
 sg13g2_nor2_1 _19113_ (.A(net553),
    .B(net463),
    .Y(_12263_));
 sg13g2_buf_2 _19114_ (.A(_12263_),
    .X(_12264_));
 sg13g2_buf_1 _19115_ (.A(_12264_),
    .X(_12265_));
 sg13g2_nand2_1 _19116_ (.Y(_12266_),
    .A(_12250_),
    .B(\mem.mem_internal.code_mem[183][0] ));
 sg13g2_nand2_1 _19117_ (.Y(_12267_),
    .A(net1118),
    .B(net228));
 sg13g2_o21ai_1 _19118_ (.B1(_12267_),
    .Y(_00850_),
    .A1(net228),
    .A2(_12266_));
 sg13g2_nand2_1 _19119_ (.Y(_12268_),
    .A(net712),
    .B(\mem.mem_internal.code_mem[183][1] ));
 sg13g2_nand2_1 _19120_ (.Y(_12269_),
    .A(net1117),
    .B(net228));
 sg13g2_o21ai_1 _19121_ (.B1(_12269_),
    .Y(_00851_),
    .A1(_12265_),
    .A2(_12268_));
 sg13g2_nand2_1 _19122_ (.Y(_12270_),
    .A(net712),
    .B(\mem.mem_internal.code_mem[183][2] ));
 sg13g2_nand2_1 _19123_ (.Y(_12271_),
    .A(net1116),
    .B(_12264_));
 sg13g2_o21ai_1 _19124_ (.B1(_12271_),
    .Y(_00852_),
    .A1(_12265_),
    .A2(_12270_));
 sg13g2_nand2_1 _19125_ (.Y(_12272_),
    .A(net712),
    .B(\mem.mem_internal.code_mem[183][3] ));
 sg13g2_nand2_1 _19126_ (.Y(_12273_),
    .A(net1115),
    .B(_12264_));
 sg13g2_o21ai_1 _19127_ (.B1(_12273_),
    .Y(_00853_),
    .A1(net228),
    .A2(_12272_));
 sg13g2_buf_1 _19128_ (.A(_11875_),
    .X(_12274_));
 sg13g2_buf_1 _19129_ (.A(_12274_),
    .X(_12275_));
 sg13g2_nand2_1 _19130_ (.Y(_12276_),
    .A(_12275_),
    .B(\mem.mem_internal.code_mem[183][4] ));
 sg13g2_nand2_1 _19131_ (.Y(_12277_),
    .A(net1114),
    .B(_12264_));
 sg13g2_o21ai_1 _19132_ (.B1(_12277_),
    .Y(_00854_),
    .A1(net228),
    .A2(_12276_));
 sg13g2_nand2_1 _19133_ (.Y(_12278_),
    .A(net711),
    .B(\mem.mem_internal.code_mem[183][5] ));
 sg13g2_nand2_1 _19134_ (.Y(_12279_),
    .A(net1113),
    .B(_12264_));
 sg13g2_o21ai_1 _19135_ (.B1(_12279_),
    .Y(_00855_),
    .A1(net228),
    .A2(_12278_));
 sg13g2_nand2_1 _19136_ (.Y(_12280_),
    .A(net711),
    .B(\mem.mem_internal.code_mem[183][6] ));
 sg13g2_nand2_1 _19137_ (.Y(_12281_),
    .A(net1112),
    .B(_12264_));
 sg13g2_o21ai_1 _19138_ (.B1(_12281_),
    .Y(_00856_),
    .A1(net228),
    .A2(_12280_));
 sg13g2_nand2_1 _19139_ (.Y(_12282_),
    .A(net711),
    .B(\mem.mem_internal.code_mem[183][7] ));
 sg13g2_nand2_1 _19140_ (.Y(_12283_),
    .A(net1111),
    .B(_12264_));
 sg13g2_o21ai_1 _19141_ (.B1(_12283_),
    .Y(_00857_),
    .A1(net228),
    .A2(_12282_));
 sg13g2_nor2_1 _19142_ (.A(net552),
    .B(net463),
    .Y(_12284_));
 sg13g2_buf_2 _19143_ (.A(_12284_),
    .X(_12285_));
 sg13g2_buf_1 _19144_ (.A(_12285_),
    .X(_12286_));
 sg13g2_nand2_1 _19145_ (.Y(_12287_),
    .A(net711),
    .B(\mem.mem_internal.code_mem[184][0] ));
 sg13g2_nand2_1 _19146_ (.Y(_12288_),
    .A(net1118),
    .B(net227));
 sg13g2_o21ai_1 _19147_ (.B1(_12288_),
    .Y(_00858_),
    .A1(_12286_),
    .A2(_12287_));
 sg13g2_nand2_1 _19148_ (.Y(_12289_),
    .A(net711),
    .B(\mem.mem_internal.code_mem[184][1] ));
 sg13g2_nand2_1 _19149_ (.Y(_12290_),
    .A(net1117),
    .B(net227));
 sg13g2_o21ai_1 _19150_ (.B1(_12290_),
    .Y(_00859_),
    .A1(net227),
    .A2(_12289_));
 sg13g2_nand2_1 _19151_ (.Y(_12291_),
    .A(net711),
    .B(\mem.mem_internal.code_mem[184][2] ));
 sg13g2_nand2_1 _19152_ (.Y(_12292_),
    .A(net1116),
    .B(_12285_));
 sg13g2_o21ai_1 _19153_ (.B1(_12292_),
    .Y(_00860_),
    .A1(net227),
    .A2(_12291_));
 sg13g2_nand2_1 _19154_ (.Y(_12293_),
    .A(net711),
    .B(\mem.mem_internal.code_mem[184][3] ));
 sg13g2_nand2_1 _19155_ (.Y(_12294_),
    .A(net1115),
    .B(_12285_));
 sg13g2_o21ai_1 _19156_ (.B1(_12294_),
    .Y(_00861_),
    .A1(_12286_),
    .A2(_12293_));
 sg13g2_nand2_1 _19157_ (.Y(_12295_),
    .A(net711),
    .B(\mem.mem_internal.code_mem[184][4] ));
 sg13g2_nand2_1 _19158_ (.Y(_12296_),
    .A(net1114),
    .B(_12285_));
 sg13g2_o21ai_1 _19159_ (.B1(_12296_),
    .Y(_00862_),
    .A1(net227),
    .A2(_12295_));
 sg13g2_nand2_1 _19160_ (.Y(_12297_),
    .A(_12275_),
    .B(\mem.mem_internal.code_mem[184][5] ));
 sg13g2_nand2_1 _19161_ (.Y(_12298_),
    .A(net1113),
    .B(_12285_));
 sg13g2_o21ai_1 _19162_ (.B1(_12298_),
    .Y(_00863_),
    .A1(net227),
    .A2(_12297_));
 sg13g2_buf_1 _19163_ (.A(_12274_),
    .X(_12299_));
 sg13g2_nand2_1 _19164_ (.Y(_12300_),
    .A(net710),
    .B(\mem.mem_internal.code_mem[184][6] ));
 sg13g2_nand2_1 _19165_ (.Y(_12301_),
    .A(net1112),
    .B(_12285_));
 sg13g2_o21ai_1 _19166_ (.B1(_12301_),
    .Y(_00864_),
    .A1(net227),
    .A2(_12300_));
 sg13g2_nand2_1 _19167_ (.Y(_12302_),
    .A(net710),
    .B(\mem.mem_internal.code_mem[184][7] ));
 sg13g2_nand2_1 _19168_ (.Y(_12303_),
    .A(net1111),
    .B(_12285_));
 sg13g2_o21ai_1 _19169_ (.B1(_12303_),
    .Y(_00865_),
    .A1(net227),
    .A2(_12302_));
 sg13g2_nor2_1 _19170_ (.A(net551),
    .B(net463),
    .Y(_12304_));
 sg13g2_buf_2 _19171_ (.A(_12304_),
    .X(_12305_));
 sg13g2_buf_1 _19172_ (.A(_12305_),
    .X(_12306_));
 sg13g2_nand2_1 _19173_ (.Y(_12307_),
    .A(_12299_),
    .B(\mem.mem_internal.code_mem[185][0] ));
 sg13g2_nand2_1 _19174_ (.Y(_12308_),
    .A(net1118),
    .B(_12306_));
 sg13g2_o21ai_1 _19175_ (.B1(_12308_),
    .Y(_00866_),
    .A1(net226),
    .A2(_12307_));
 sg13g2_nand2_1 _19176_ (.Y(_12309_),
    .A(net710),
    .B(\mem.mem_internal.code_mem[185][1] ));
 sg13g2_nand2_1 _19177_ (.Y(_12310_),
    .A(net1117),
    .B(net226));
 sg13g2_o21ai_1 _19178_ (.B1(_12310_),
    .Y(_00867_),
    .A1(net226),
    .A2(_12309_));
 sg13g2_nand2_1 _19179_ (.Y(_12311_),
    .A(net710),
    .B(\mem.mem_internal.code_mem[185][2] ));
 sg13g2_nand2_1 _19180_ (.Y(_12312_),
    .A(_12226_),
    .B(_12305_));
 sg13g2_o21ai_1 _19181_ (.B1(_12312_),
    .Y(_00868_),
    .A1(net226),
    .A2(_12311_));
 sg13g2_nand2_1 _19182_ (.Y(_12313_),
    .A(_12299_),
    .B(\mem.mem_internal.code_mem[185][3] ));
 sg13g2_nand2_1 _19183_ (.Y(_12314_),
    .A(_12229_),
    .B(_12305_));
 sg13g2_o21ai_1 _19184_ (.B1(_12314_),
    .Y(_00869_),
    .A1(_12306_),
    .A2(_12313_));
 sg13g2_nand2_1 _19185_ (.Y(_12315_),
    .A(net710),
    .B(\mem.mem_internal.code_mem[185][4] ));
 sg13g2_nand2_1 _19186_ (.Y(_12316_),
    .A(net1114),
    .B(_12305_));
 sg13g2_o21ai_1 _19187_ (.B1(_12316_),
    .Y(_00870_),
    .A1(net226),
    .A2(_12315_));
 sg13g2_nand2_1 _19188_ (.Y(_12317_),
    .A(net710),
    .B(\mem.mem_internal.code_mem[185][5] ));
 sg13g2_nand2_1 _19189_ (.Y(_12318_),
    .A(_12235_),
    .B(_12305_));
 sg13g2_o21ai_1 _19190_ (.B1(_12318_),
    .Y(_00871_),
    .A1(net226),
    .A2(_12317_));
 sg13g2_nand2_1 _19191_ (.Y(_12319_),
    .A(net710),
    .B(\mem.mem_internal.code_mem[185][6] ));
 sg13g2_nand2_1 _19192_ (.Y(_12320_),
    .A(_12238_),
    .B(_12305_));
 sg13g2_o21ai_1 _19193_ (.B1(_12320_),
    .Y(_00872_),
    .A1(net226),
    .A2(_12319_));
 sg13g2_nand2_1 _19194_ (.Y(_12321_),
    .A(net710),
    .B(\mem.mem_internal.code_mem[185][7] ));
 sg13g2_nand2_1 _19195_ (.Y(_12322_),
    .A(net1111),
    .B(_12305_));
 sg13g2_o21ai_1 _19196_ (.B1(_12322_),
    .Y(_00873_),
    .A1(net226),
    .A2(_12321_));
 sg13g2_nor2_1 _19197_ (.A(net550),
    .B(_12095_),
    .Y(_12323_));
 sg13g2_buf_2 _19198_ (.A(_12323_),
    .X(_12324_));
 sg13g2_buf_1 _19199_ (.A(_12324_),
    .X(_12325_));
 sg13g2_buf_1 _19200_ (.A(_12274_),
    .X(_12326_));
 sg13g2_nand2_1 _19201_ (.Y(_12327_),
    .A(_12326_),
    .B(\mem.mem_internal.code_mem[186][0] ));
 sg13g2_nand2_1 _19202_ (.Y(_12328_),
    .A(net1118),
    .B(net372));
 sg13g2_o21ai_1 _19203_ (.B1(_12328_),
    .Y(_00874_),
    .A1(_12325_),
    .A2(_12327_));
 sg13g2_nand2_1 _19204_ (.Y(_12329_),
    .A(net709),
    .B(\mem.mem_internal.code_mem[186][1] ));
 sg13g2_nand2_1 _19205_ (.Y(_12330_),
    .A(net1117),
    .B(net372));
 sg13g2_o21ai_1 _19206_ (.B1(_12330_),
    .Y(_00875_),
    .A1(net372),
    .A2(_12329_));
 sg13g2_nand2_1 _19207_ (.Y(_12331_),
    .A(net709),
    .B(\mem.mem_internal.code_mem[186][2] ));
 sg13g2_nand2_1 _19208_ (.Y(_12332_),
    .A(net1116),
    .B(_12324_));
 sg13g2_o21ai_1 _19209_ (.B1(_12332_),
    .Y(_00876_),
    .A1(net372),
    .A2(_12331_));
 sg13g2_nand2_1 _19210_ (.Y(_12333_),
    .A(_12326_),
    .B(\mem.mem_internal.code_mem[186][3] ));
 sg13g2_nand2_1 _19211_ (.Y(_12334_),
    .A(net1115),
    .B(_12324_));
 sg13g2_o21ai_1 _19212_ (.B1(_12334_),
    .Y(_00877_),
    .A1(_12325_),
    .A2(_12333_));
 sg13g2_nand2_1 _19213_ (.Y(_12335_),
    .A(net709),
    .B(\mem.mem_internal.code_mem[186][4] ));
 sg13g2_nand2_1 _19214_ (.Y(_12336_),
    .A(_12232_),
    .B(_12324_));
 sg13g2_o21ai_1 _19215_ (.B1(_12336_),
    .Y(_00878_),
    .A1(net372),
    .A2(_12335_));
 sg13g2_nand2_1 _19216_ (.Y(_12337_),
    .A(net709),
    .B(\mem.mem_internal.code_mem[186][5] ));
 sg13g2_nand2_1 _19217_ (.Y(_12338_),
    .A(net1113),
    .B(_12324_));
 sg13g2_o21ai_1 _19218_ (.B1(_12338_),
    .Y(_00879_),
    .A1(net372),
    .A2(_12337_));
 sg13g2_nand2_1 _19219_ (.Y(_12339_),
    .A(net709),
    .B(\mem.mem_internal.code_mem[186][6] ));
 sg13g2_nand2_1 _19220_ (.Y(_12340_),
    .A(net1112),
    .B(_12324_));
 sg13g2_o21ai_1 _19221_ (.B1(_12340_),
    .Y(_00880_),
    .A1(net372),
    .A2(_12339_));
 sg13g2_nand2_1 _19222_ (.Y(_12341_),
    .A(net709),
    .B(\mem.mem_internal.code_mem[186][7] ));
 sg13g2_nand2_1 _19223_ (.Y(_12342_),
    .A(_12241_),
    .B(_12324_));
 sg13g2_o21ai_1 _19224_ (.B1(_12342_),
    .Y(_00881_),
    .A1(net372),
    .A2(_12341_));
 sg13g2_nor2_1 _19225_ (.A(net549),
    .B(_12095_),
    .Y(_12343_));
 sg13g2_buf_1 _19226_ (.A(_12343_),
    .X(_12344_));
 sg13g2_buf_1 _19227_ (.A(_12344_),
    .X(_12345_));
 sg13g2_nand2_1 _19228_ (.Y(_12346_),
    .A(net709),
    .B(\mem.mem_internal.code_mem[187][0] ));
 sg13g2_nand2_1 _19229_ (.Y(_12347_),
    .A(_12220_),
    .B(net371));
 sg13g2_o21ai_1 _19230_ (.B1(_12347_),
    .Y(_00882_),
    .A1(net371),
    .A2(_12346_));
 sg13g2_nand2_1 _19231_ (.Y(_12348_),
    .A(net709),
    .B(\mem.mem_internal.code_mem[187][1] ));
 sg13g2_nand2_1 _19232_ (.Y(_12349_),
    .A(net1117),
    .B(net371));
 sg13g2_o21ai_1 _19233_ (.B1(_12349_),
    .Y(_00883_),
    .A1(net371),
    .A2(_12348_));
 sg13g2_buf_1 _19234_ (.A(_12274_),
    .X(_12350_));
 sg13g2_nand2_1 _19235_ (.Y(_12351_),
    .A(_12350_),
    .B(\mem.mem_internal.code_mem[187][2] ));
 sg13g2_nand2_1 _19236_ (.Y(_12352_),
    .A(net1116),
    .B(_12344_));
 sg13g2_o21ai_1 _19237_ (.B1(_12352_),
    .Y(_00884_),
    .A1(net371),
    .A2(_12351_));
 sg13g2_nand2_1 _19238_ (.Y(_12353_),
    .A(net708),
    .B(\mem.mem_internal.code_mem[187][3] ));
 sg13g2_nand2_1 _19239_ (.Y(_12354_),
    .A(net1115),
    .B(_12344_));
 sg13g2_o21ai_1 _19240_ (.B1(_12354_),
    .Y(_00885_),
    .A1(_12345_),
    .A2(_12353_));
 sg13g2_nand2_1 _19241_ (.Y(_12355_),
    .A(net708),
    .B(\mem.mem_internal.code_mem[187][4] ));
 sg13g2_nand2_1 _19242_ (.Y(_12356_),
    .A(_12232_),
    .B(_12344_));
 sg13g2_o21ai_1 _19243_ (.B1(_12356_),
    .Y(_00886_),
    .A1(net371),
    .A2(_12355_));
 sg13g2_nand2_1 _19244_ (.Y(_12357_),
    .A(net708),
    .B(\mem.mem_internal.code_mem[187][5] ));
 sg13g2_nand2_1 _19245_ (.Y(_12358_),
    .A(net1113),
    .B(_12344_));
 sg13g2_o21ai_1 _19246_ (.B1(_12358_),
    .Y(_00887_),
    .A1(net371),
    .A2(_12357_));
 sg13g2_nand2_1 _19247_ (.Y(_12359_),
    .A(net708),
    .B(\mem.mem_internal.code_mem[187][6] ));
 sg13g2_nand2_1 _19248_ (.Y(_12360_),
    .A(net1112),
    .B(_12344_));
 sg13g2_o21ai_1 _19249_ (.B1(_12360_),
    .Y(_00888_),
    .A1(net371),
    .A2(_12359_));
 sg13g2_nand2_1 _19250_ (.Y(_12361_),
    .A(net708),
    .B(\mem.mem_internal.code_mem[187][7] ));
 sg13g2_nand2_1 _19251_ (.Y(_12362_),
    .A(_12241_),
    .B(_12344_));
 sg13g2_o21ai_1 _19252_ (.B1(_12362_),
    .Y(_00889_),
    .A1(_12345_),
    .A2(_12361_));
 sg13g2_nor2_1 _19253_ (.A(net773),
    .B(_12095_),
    .Y(_12363_));
 sg13g2_buf_2 _19254_ (.A(_12363_),
    .X(_12364_));
 sg13g2_buf_1 _19255_ (.A(_12364_),
    .X(_12365_));
 sg13g2_nand2_1 _19256_ (.Y(_12366_),
    .A(net708),
    .B(\mem.mem_internal.code_mem[188][0] ));
 sg13g2_nand2_1 _19257_ (.Y(_12367_),
    .A(net1118),
    .B(net370));
 sg13g2_o21ai_1 _19258_ (.B1(_12367_),
    .Y(_00890_),
    .A1(net370),
    .A2(_12366_));
 sg13g2_nand2_1 _19259_ (.Y(_12368_),
    .A(net708),
    .B(\mem.mem_internal.code_mem[188][1] ));
 sg13g2_nand2_1 _19260_ (.Y(_12369_),
    .A(net1117),
    .B(net370));
 sg13g2_o21ai_1 _19261_ (.B1(_12369_),
    .Y(_00891_),
    .A1(net370),
    .A2(_12368_));
 sg13g2_nand2_1 _19262_ (.Y(_12370_),
    .A(net708),
    .B(\mem.mem_internal.code_mem[188][2] ));
 sg13g2_nand2_1 _19263_ (.Y(_12371_),
    .A(net1116),
    .B(_12364_));
 sg13g2_o21ai_1 _19264_ (.B1(_12371_),
    .Y(_00892_),
    .A1(net370),
    .A2(_12370_));
 sg13g2_nand2_1 _19265_ (.Y(_12372_),
    .A(_12350_),
    .B(\mem.mem_internal.code_mem[188][3] ));
 sg13g2_nand2_1 _19266_ (.Y(_12373_),
    .A(net1115),
    .B(_12364_));
 sg13g2_o21ai_1 _19267_ (.B1(_12373_),
    .Y(_00893_),
    .A1(net370),
    .A2(_12372_));
 sg13g2_buf_1 _19268_ (.A(_12274_),
    .X(_12374_));
 sg13g2_nand2_1 _19269_ (.Y(_12375_),
    .A(net707),
    .B(\mem.mem_internal.code_mem[188][4] ));
 sg13g2_nand2_1 _19270_ (.Y(_12376_),
    .A(net1114),
    .B(_12364_));
 sg13g2_o21ai_1 _19271_ (.B1(_12376_),
    .Y(_00894_),
    .A1(net370),
    .A2(_12375_));
 sg13g2_nand2_1 _19272_ (.Y(_12377_),
    .A(net707),
    .B(\mem.mem_internal.code_mem[188][5] ));
 sg13g2_nand2_1 _19273_ (.Y(_12378_),
    .A(_12235_),
    .B(_12364_));
 sg13g2_o21ai_1 _19274_ (.B1(_12378_),
    .Y(_00895_),
    .A1(net370),
    .A2(_12377_));
 sg13g2_nand2_1 _19275_ (.Y(_12379_),
    .A(net707),
    .B(\mem.mem_internal.code_mem[188][6] ));
 sg13g2_nand2_1 _19276_ (.Y(_12380_),
    .A(_12238_),
    .B(_12364_));
 sg13g2_o21ai_1 _19277_ (.B1(_12380_),
    .Y(_00896_),
    .A1(_12365_),
    .A2(_12379_));
 sg13g2_nand2_1 _19278_ (.Y(_12381_),
    .A(net707),
    .B(\mem.mem_internal.code_mem[188][7] ));
 sg13g2_nand2_1 _19279_ (.Y(_12382_),
    .A(net1111),
    .B(_12364_));
 sg13g2_o21ai_1 _19280_ (.B1(_12382_),
    .Y(_00897_),
    .A1(_12365_),
    .A2(_12381_));
 sg13g2_nor2_1 _19281_ (.A(net548),
    .B(_12095_),
    .Y(_12383_));
 sg13g2_buf_2 _19282_ (.A(_12383_),
    .X(_12384_));
 sg13g2_buf_1 _19283_ (.A(_12384_),
    .X(_12385_));
 sg13g2_nand2_1 _19284_ (.Y(_12386_),
    .A(net707),
    .B(\mem.mem_internal.code_mem[189][0] ));
 sg13g2_nand2_1 _19285_ (.Y(_12387_),
    .A(net1118),
    .B(net369));
 sg13g2_o21ai_1 _19286_ (.B1(_12387_),
    .Y(_00898_),
    .A1(net369),
    .A2(_12386_));
 sg13g2_nand2_1 _19287_ (.Y(_12388_),
    .A(net707),
    .B(\mem.mem_internal.code_mem[189][1] ));
 sg13g2_nand2_1 _19288_ (.Y(_12389_),
    .A(_12223_),
    .B(net369));
 sg13g2_o21ai_1 _19289_ (.B1(_12389_),
    .Y(_00899_),
    .A1(net369),
    .A2(_12388_));
 sg13g2_nand2_1 _19290_ (.Y(_12390_),
    .A(net707),
    .B(\mem.mem_internal.code_mem[189][2] ));
 sg13g2_nand2_1 _19291_ (.Y(_12391_),
    .A(net1116),
    .B(_12384_));
 sg13g2_o21ai_1 _19292_ (.B1(_12391_),
    .Y(_00900_),
    .A1(_12385_),
    .A2(_12390_));
 sg13g2_nand2_1 _19293_ (.Y(_12392_),
    .A(net707),
    .B(\mem.mem_internal.code_mem[189][3] ));
 sg13g2_nand2_1 _19294_ (.Y(_12393_),
    .A(net1115),
    .B(_12384_));
 sg13g2_o21ai_1 _19295_ (.B1(_12393_),
    .Y(_00901_),
    .A1(_12385_),
    .A2(_12392_));
 sg13g2_nand2_1 _19296_ (.Y(_12394_),
    .A(_12374_),
    .B(\mem.mem_internal.code_mem[189][4] ));
 sg13g2_nand2_1 _19297_ (.Y(_12395_),
    .A(net1114),
    .B(_12384_));
 sg13g2_o21ai_1 _19298_ (.B1(_12395_),
    .Y(_00902_),
    .A1(net369),
    .A2(_12394_));
 sg13g2_nand2_1 _19299_ (.Y(_12396_),
    .A(_12374_),
    .B(\mem.mem_internal.code_mem[189][5] ));
 sg13g2_nand2_1 _19300_ (.Y(_12397_),
    .A(net1113),
    .B(_12384_));
 sg13g2_o21ai_1 _19301_ (.B1(_12397_),
    .Y(_00903_),
    .A1(net369),
    .A2(_12396_));
 sg13g2_buf_1 _19302_ (.A(_12274_),
    .X(_12398_));
 sg13g2_nand2_1 _19303_ (.Y(_12399_),
    .A(net706),
    .B(\mem.mem_internal.code_mem[189][6] ));
 sg13g2_nand2_1 _19304_ (.Y(_12400_),
    .A(net1112),
    .B(_12384_));
 sg13g2_o21ai_1 _19305_ (.B1(_12400_),
    .Y(_00904_),
    .A1(net369),
    .A2(_12399_));
 sg13g2_nand2_1 _19306_ (.Y(_12401_),
    .A(net706),
    .B(\mem.mem_internal.code_mem[189][7] ));
 sg13g2_nand2_1 _19307_ (.Y(_12402_),
    .A(net1111),
    .B(_12384_));
 sg13g2_o21ai_1 _19308_ (.B1(_12402_),
    .Y(_00905_),
    .A1(net369),
    .A2(_12401_));
 sg13g2_buf_1 _19309_ (.A(_11058_),
    .X(_12403_));
 sg13g2_nand2_1 _19310_ (.Y(_12404_),
    .A(net844),
    .B(\mem.mem_internal.code_mem[18][0] ));
 sg13g2_nor2_1 _19311_ (.A(net527),
    .B(net464),
    .Y(_12405_));
 sg13g2_buf_2 _19312_ (.A(_12405_),
    .X(_12406_));
 sg13g2_buf_1 _19313_ (.A(_12406_),
    .X(_12407_));
 sg13g2_nand2_1 _19314_ (.Y(_12408_),
    .A(_12220_),
    .B(net225));
 sg13g2_o21ai_1 _19315_ (.B1(_12408_),
    .Y(_00906_),
    .A1(_12404_),
    .A2(net225));
 sg13g2_nand2_1 _19316_ (.Y(_12409_),
    .A(net706),
    .B(\mem.mem_internal.code_mem[18][1] ));
 sg13g2_nand2_1 _19317_ (.Y(_12410_),
    .A(_12223_),
    .B(net225));
 sg13g2_o21ai_1 _19318_ (.B1(_12410_),
    .Y(_00907_),
    .A1(net225),
    .A2(_12409_));
 sg13g2_nand2_1 _19319_ (.Y(_12411_),
    .A(net706),
    .B(\mem.mem_internal.code_mem[18][2] ));
 sg13g2_nand2_1 _19320_ (.Y(_12412_),
    .A(_12226_),
    .B(_12406_));
 sg13g2_o21ai_1 _19321_ (.B1(_12412_),
    .Y(_00908_),
    .A1(net225),
    .A2(_12411_));
 sg13g2_nand2_1 _19322_ (.Y(_12413_),
    .A(net706),
    .B(\mem.mem_internal.code_mem[18][3] ));
 sg13g2_nand2_1 _19323_ (.Y(_12414_),
    .A(_12229_),
    .B(_12406_));
 sg13g2_o21ai_1 _19324_ (.B1(_12414_),
    .Y(_00909_),
    .A1(net225),
    .A2(_12413_));
 sg13g2_nand2_1 _19325_ (.Y(_12415_),
    .A(net706),
    .B(\mem.mem_internal.code_mem[18][4] ));
 sg13g2_nand2_1 _19326_ (.Y(_12416_),
    .A(net1114),
    .B(_12406_));
 sg13g2_o21ai_1 _19327_ (.B1(_12416_),
    .Y(_00910_),
    .A1(_12407_),
    .A2(_12415_));
 sg13g2_nand2_1 _19328_ (.Y(_12417_),
    .A(net706),
    .B(\mem.mem_internal.code_mem[18][5] ));
 sg13g2_nand2_1 _19329_ (.Y(_12418_),
    .A(net1113),
    .B(_12406_));
 sg13g2_o21ai_1 _19330_ (.B1(_12418_),
    .Y(_00911_),
    .A1(net225),
    .A2(_12417_));
 sg13g2_nand2_1 _19331_ (.Y(_12419_),
    .A(_12398_),
    .B(\mem.mem_internal.code_mem[18][6] ));
 sg13g2_nand2_1 _19332_ (.Y(_12420_),
    .A(net1112),
    .B(_12406_));
 sg13g2_o21ai_1 _19333_ (.B1(_12420_),
    .Y(_00912_),
    .A1(net225),
    .A2(_12419_));
 sg13g2_nand2_1 _19334_ (.Y(_12421_),
    .A(_12398_),
    .B(\mem.mem_internal.code_mem[18][7] ));
 sg13g2_nand2_1 _19335_ (.Y(_12422_),
    .A(net1111),
    .B(_12406_));
 sg13g2_o21ai_1 _19336_ (.B1(_12422_),
    .Y(_00913_),
    .A1(_12407_),
    .A2(_12421_));
 sg13g2_nor2_1 _19337_ (.A(net547),
    .B(_12095_),
    .Y(_12423_));
 sg13g2_buf_1 _19338_ (.A(_12423_),
    .X(_12424_));
 sg13g2_buf_1 _19339_ (.A(_12424_),
    .X(_12425_));
 sg13g2_nand2_1 _19340_ (.Y(_12426_),
    .A(net706),
    .B(\mem.mem_internal.code_mem[190][0] ));
 sg13g2_buf_1 _19341_ (.A(_11163_),
    .X(_12427_));
 sg13g2_nand2_1 _19342_ (.Y(_12428_),
    .A(net1110),
    .B(net368));
 sg13g2_o21ai_1 _19343_ (.B1(_12428_),
    .Y(_00914_),
    .A1(net368),
    .A2(_12426_));
 sg13g2_buf_1 _19344_ (.A(_12274_),
    .X(_12429_));
 sg13g2_nand2_1 _19345_ (.Y(_12430_),
    .A(net705),
    .B(\mem.mem_internal.code_mem[190][1] ));
 sg13g2_buf_1 _19346_ (.A(_11167_),
    .X(_12431_));
 sg13g2_nand2_1 _19347_ (.Y(_12432_),
    .A(net1109),
    .B(net368));
 sg13g2_o21ai_1 _19348_ (.B1(_12432_),
    .Y(_00915_),
    .A1(net368),
    .A2(_12430_));
 sg13g2_nand2_1 _19349_ (.Y(_12433_),
    .A(net705),
    .B(\mem.mem_internal.code_mem[190][2] ));
 sg13g2_buf_1 _19350_ (.A(_11171_),
    .X(_12434_));
 sg13g2_nand2_1 _19351_ (.Y(_12435_),
    .A(net1108),
    .B(_12424_));
 sg13g2_o21ai_1 _19352_ (.B1(_12435_),
    .Y(_00916_),
    .A1(net368),
    .A2(_12433_));
 sg13g2_nand2_1 _19353_ (.Y(_12436_),
    .A(net705),
    .B(\mem.mem_internal.code_mem[190][3] ));
 sg13g2_buf_1 _19354_ (.A(_11175_),
    .X(_12437_));
 sg13g2_nand2_1 _19355_ (.Y(_12438_),
    .A(net1107),
    .B(_12424_));
 sg13g2_o21ai_1 _19356_ (.B1(_12438_),
    .Y(_00917_),
    .A1(net368),
    .A2(_12436_));
 sg13g2_nand2_1 _19357_ (.Y(_12439_),
    .A(net705),
    .B(\mem.mem_internal.code_mem[190][4] ));
 sg13g2_buf_1 _19358_ (.A(_11179_),
    .X(_12440_));
 sg13g2_nand2_1 _19359_ (.Y(_12441_),
    .A(net1106),
    .B(_12424_));
 sg13g2_o21ai_1 _19360_ (.B1(_12441_),
    .Y(_00918_),
    .A1(_12425_),
    .A2(_12439_));
 sg13g2_nand2_1 _19361_ (.Y(_12442_),
    .A(net705),
    .B(\mem.mem_internal.code_mem[190][5] ));
 sg13g2_buf_1 _19362_ (.A(_11183_),
    .X(_12443_));
 sg13g2_nand2_1 _19363_ (.Y(_12444_),
    .A(net1105),
    .B(_12424_));
 sg13g2_o21ai_1 _19364_ (.B1(_12444_),
    .Y(_00919_),
    .A1(_12425_),
    .A2(_12442_));
 sg13g2_nand2_1 _19365_ (.Y(_12445_),
    .A(_12429_),
    .B(\mem.mem_internal.code_mem[190][6] ));
 sg13g2_buf_1 _19366_ (.A(_11188_),
    .X(_12446_));
 sg13g2_nand2_1 _19367_ (.Y(_12447_),
    .A(net1104),
    .B(_12424_));
 sg13g2_o21ai_1 _19368_ (.B1(_12447_),
    .Y(_00920_),
    .A1(net368),
    .A2(_12445_));
 sg13g2_nand2_1 _19369_ (.Y(_12448_),
    .A(_12429_),
    .B(\mem.mem_internal.code_mem[190][7] ));
 sg13g2_buf_1 _19370_ (.A(_11192_),
    .X(_12449_));
 sg13g2_nand2_1 _19371_ (.Y(_12450_),
    .A(net1103),
    .B(_12424_));
 sg13g2_o21ai_1 _19372_ (.B1(_12450_),
    .Y(_00921_),
    .A1(net368),
    .A2(_12448_));
 sg13g2_nor2_1 _19373_ (.A(net770),
    .B(_12095_),
    .Y(_12451_));
 sg13g2_buf_2 _19374_ (.A(_12451_),
    .X(_12452_));
 sg13g2_buf_1 _19375_ (.A(_12452_),
    .X(_12453_));
 sg13g2_nand2_1 _19376_ (.Y(_12454_),
    .A(net705),
    .B(\mem.mem_internal.code_mem[191][0] ));
 sg13g2_nand2_1 _19377_ (.Y(_12455_),
    .A(net1110),
    .B(net367));
 sg13g2_o21ai_1 _19378_ (.B1(_12455_),
    .Y(_00922_),
    .A1(net367),
    .A2(_12454_));
 sg13g2_nand2_1 _19379_ (.Y(_12456_),
    .A(net705),
    .B(\mem.mem_internal.code_mem[191][1] ));
 sg13g2_nand2_1 _19380_ (.Y(_12457_),
    .A(net1109),
    .B(net367));
 sg13g2_o21ai_1 _19381_ (.B1(_12457_),
    .Y(_00923_),
    .A1(net367),
    .A2(_12456_));
 sg13g2_nand2_1 _19382_ (.Y(_12458_),
    .A(net705),
    .B(\mem.mem_internal.code_mem[191][2] ));
 sg13g2_nand2_1 _19383_ (.Y(_12459_),
    .A(net1108),
    .B(_12452_));
 sg13g2_o21ai_1 _19384_ (.B1(_12459_),
    .Y(_00924_),
    .A1(net367),
    .A2(_12458_));
 sg13g2_buf_1 _19385_ (.A(_11875_),
    .X(_12460_));
 sg13g2_buf_1 _19386_ (.A(_12460_),
    .X(_12461_));
 sg13g2_nand2_1 _19387_ (.Y(_12462_),
    .A(net704),
    .B(\mem.mem_internal.code_mem[191][3] ));
 sg13g2_nand2_1 _19388_ (.Y(_12463_),
    .A(net1107),
    .B(_12452_));
 sg13g2_o21ai_1 _19389_ (.B1(_12463_),
    .Y(_00925_),
    .A1(net367),
    .A2(_12462_));
 sg13g2_nand2_1 _19390_ (.Y(_12464_),
    .A(net704),
    .B(\mem.mem_internal.code_mem[191][4] ));
 sg13g2_nand2_1 _19391_ (.Y(_12465_),
    .A(net1106),
    .B(_12452_));
 sg13g2_o21ai_1 _19392_ (.B1(_12465_),
    .Y(_00926_),
    .A1(net367),
    .A2(_12464_));
 sg13g2_nand2_1 _19393_ (.Y(_12466_),
    .A(net704),
    .B(\mem.mem_internal.code_mem[191][5] ));
 sg13g2_nand2_1 _19394_ (.Y(_12467_),
    .A(net1105),
    .B(_12452_));
 sg13g2_o21ai_1 _19395_ (.B1(_12467_),
    .Y(_00927_),
    .A1(net367),
    .A2(_12466_));
 sg13g2_nand2_1 _19396_ (.Y(_12468_),
    .A(net704),
    .B(\mem.mem_internal.code_mem[191][6] ));
 sg13g2_nand2_1 _19397_ (.Y(_12469_),
    .A(net1104),
    .B(_12452_));
 sg13g2_o21ai_1 _19398_ (.B1(_12469_),
    .Y(_00928_),
    .A1(_12453_),
    .A2(_12468_));
 sg13g2_nand2_1 _19399_ (.Y(_12470_),
    .A(net704),
    .B(\mem.mem_internal.code_mem[191][7] ));
 sg13g2_nand2_1 _19400_ (.Y(_12471_),
    .A(net1103),
    .B(_12452_));
 sg13g2_o21ai_1 _19401_ (.B1(_12471_),
    .Y(_00929_),
    .A1(_12453_),
    .A2(_12470_));
 sg13g2_nand2_1 _19402_ (.Y(_12472_),
    .A(net844),
    .B(\mem.mem_internal.code_mem[192][0] ));
 sg13g2_nand3_1 _19403_ (.B(_10033_),
    .C(_10244_),
    .A(net1297),
    .Y(_12473_));
 sg13g2_buf_2 _19404_ (.A(_12473_),
    .X(_12474_));
 sg13g2_buf_1 _19405_ (.A(_12474_),
    .X(_12475_));
 sg13g2_nor2_1 _19406_ (.A(_10233_),
    .B(net462),
    .Y(_12476_));
 sg13g2_buf_2 _19407_ (.A(_12476_),
    .X(_12477_));
 sg13g2_buf_1 _19408_ (.A(_12477_),
    .X(_12478_));
 sg13g2_nand2_1 _19409_ (.Y(_12479_),
    .A(net1110),
    .B(net224));
 sg13g2_o21ai_1 _19410_ (.B1(_12479_),
    .Y(_00930_),
    .A1(_12472_),
    .A2(net224));
 sg13g2_nand2_1 _19411_ (.Y(_12480_),
    .A(net704),
    .B(\mem.mem_internal.code_mem[192][1] ));
 sg13g2_nand2_1 _19412_ (.Y(_12481_),
    .A(net1109),
    .B(net224));
 sg13g2_o21ai_1 _19413_ (.B1(_12481_),
    .Y(_00931_),
    .A1(net224),
    .A2(_12480_));
 sg13g2_nand2_1 _19414_ (.Y(_12482_),
    .A(net704),
    .B(\mem.mem_internal.code_mem[192][2] ));
 sg13g2_nand2_1 _19415_ (.Y(_12483_),
    .A(net1108),
    .B(_12477_));
 sg13g2_o21ai_1 _19416_ (.B1(_12483_),
    .Y(_00932_),
    .A1(net224),
    .A2(_12482_));
 sg13g2_nand2_1 _19417_ (.Y(_12484_),
    .A(net704),
    .B(\mem.mem_internal.code_mem[192][3] ));
 sg13g2_nand2_1 _19418_ (.Y(_12485_),
    .A(net1107),
    .B(_12477_));
 sg13g2_o21ai_1 _19419_ (.B1(_12485_),
    .Y(_00933_),
    .A1(_12478_),
    .A2(_12484_));
 sg13g2_nand2_1 _19420_ (.Y(_12486_),
    .A(_12461_),
    .B(\mem.mem_internal.code_mem[192][4] ));
 sg13g2_nand2_1 _19421_ (.Y(_12487_),
    .A(net1106),
    .B(_12477_));
 sg13g2_o21ai_1 _19422_ (.B1(_12487_),
    .Y(_00934_),
    .A1(_12478_),
    .A2(_12486_));
 sg13g2_nand2_1 _19423_ (.Y(_12488_),
    .A(_12461_),
    .B(\mem.mem_internal.code_mem[192][5] ));
 sg13g2_nand2_1 _19424_ (.Y(_12489_),
    .A(net1105),
    .B(_12477_));
 sg13g2_o21ai_1 _19425_ (.B1(_12489_),
    .Y(_00935_),
    .A1(net224),
    .A2(_12488_));
 sg13g2_buf_1 _19426_ (.A(_12460_),
    .X(_12490_));
 sg13g2_nand2_1 _19427_ (.Y(_12491_),
    .A(net703),
    .B(\mem.mem_internal.code_mem[192][6] ));
 sg13g2_nand2_1 _19428_ (.Y(_12492_),
    .A(net1104),
    .B(_12477_));
 sg13g2_o21ai_1 _19429_ (.B1(_12492_),
    .Y(_00936_),
    .A1(net224),
    .A2(_12491_));
 sg13g2_nand2_1 _19430_ (.Y(_12493_),
    .A(net703),
    .B(\mem.mem_internal.code_mem[192][7] ));
 sg13g2_nand2_1 _19431_ (.Y(_12494_),
    .A(net1103),
    .B(_12477_));
 sg13g2_o21ai_1 _19432_ (.B1(_12494_),
    .Y(_00937_),
    .A1(net224),
    .A2(_12493_));
 sg13g2_nand2_1 _19433_ (.Y(_12495_),
    .A(net844),
    .B(\mem.mem_internal.code_mem[193][0] ));
 sg13g2_nor2_1 _19434_ (.A(_10632_),
    .B(net462),
    .Y(_12496_));
 sg13g2_buf_2 _19435_ (.A(_12496_),
    .X(_12497_));
 sg13g2_buf_1 _19436_ (.A(_12497_),
    .X(_12498_));
 sg13g2_nand2_1 _19437_ (.Y(_12499_),
    .A(net1110),
    .B(net223));
 sg13g2_o21ai_1 _19438_ (.B1(_12499_),
    .Y(_00938_),
    .A1(_12495_),
    .A2(net223));
 sg13g2_nand2_1 _19439_ (.Y(_12500_),
    .A(net703),
    .B(\mem.mem_internal.code_mem[193][1] ));
 sg13g2_nand2_1 _19440_ (.Y(_12501_),
    .A(net1109),
    .B(net223));
 sg13g2_o21ai_1 _19441_ (.B1(_12501_),
    .Y(_00939_),
    .A1(net223),
    .A2(_12500_));
 sg13g2_nand2_1 _19442_ (.Y(_12502_),
    .A(net703),
    .B(\mem.mem_internal.code_mem[193][2] ));
 sg13g2_nand2_1 _19443_ (.Y(_12503_),
    .A(net1108),
    .B(_12497_));
 sg13g2_o21ai_1 _19444_ (.B1(_12503_),
    .Y(_00940_),
    .A1(net223),
    .A2(_12502_));
 sg13g2_nand2_1 _19445_ (.Y(_12504_),
    .A(_12490_),
    .B(\mem.mem_internal.code_mem[193][3] ));
 sg13g2_nand2_1 _19446_ (.Y(_12505_),
    .A(net1107),
    .B(_12497_));
 sg13g2_o21ai_1 _19447_ (.B1(_12505_),
    .Y(_00941_),
    .A1(net223),
    .A2(_12504_));
 sg13g2_nand2_1 _19448_ (.Y(_12506_),
    .A(net703),
    .B(\mem.mem_internal.code_mem[193][4] ));
 sg13g2_nand2_1 _19449_ (.Y(_12507_),
    .A(net1106),
    .B(_12497_));
 sg13g2_o21ai_1 _19450_ (.B1(_12507_),
    .Y(_00942_),
    .A1(_12498_),
    .A2(_12506_));
 sg13g2_nand2_1 _19451_ (.Y(_12508_),
    .A(net703),
    .B(\mem.mem_internal.code_mem[193][5] ));
 sg13g2_nand2_1 _19452_ (.Y(_12509_),
    .A(net1105),
    .B(_12497_));
 sg13g2_o21ai_1 _19453_ (.B1(_12509_),
    .Y(_00943_),
    .A1(net223),
    .A2(_12508_));
 sg13g2_nand2_1 _19454_ (.Y(_12510_),
    .A(net703),
    .B(\mem.mem_internal.code_mem[193][6] ));
 sg13g2_nand2_1 _19455_ (.Y(_12511_),
    .A(net1104),
    .B(_12497_));
 sg13g2_o21ai_1 _19456_ (.B1(_12511_),
    .Y(_00944_),
    .A1(_12498_),
    .A2(_12510_));
 sg13g2_nand2_1 _19457_ (.Y(_12512_),
    .A(net703),
    .B(\mem.mem_internal.code_mem[193][7] ));
 sg13g2_nand2_1 _19458_ (.Y(_12513_),
    .A(net1103),
    .B(_12497_));
 sg13g2_o21ai_1 _19459_ (.B1(_12513_),
    .Y(_00945_),
    .A1(net223),
    .A2(_12512_));
 sg13g2_nand2_1 _19460_ (.Y(_12514_),
    .A(net844),
    .B(\mem.mem_internal.code_mem[194][0] ));
 sg13g2_nor2_1 _19461_ (.A(_10656_),
    .B(net462),
    .Y(_12515_));
 sg13g2_buf_2 _19462_ (.A(_12515_),
    .X(_12516_));
 sg13g2_buf_1 _19463_ (.A(_12516_),
    .X(_12517_));
 sg13g2_nand2_1 _19464_ (.Y(_12518_),
    .A(net1110),
    .B(net222));
 sg13g2_o21ai_1 _19465_ (.B1(_12518_),
    .Y(_00946_),
    .A1(_12514_),
    .A2(net222));
 sg13g2_nand2_1 _19466_ (.Y(_12519_),
    .A(_12490_),
    .B(\mem.mem_internal.code_mem[194][1] ));
 sg13g2_nand2_1 _19467_ (.Y(_12520_),
    .A(net1109),
    .B(net222));
 sg13g2_o21ai_1 _19468_ (.B1(_12520_),
    .Y(_00947_),
    .A1(net222),
    .A2(_12519_));
 sg13g2_buf_1 _19469_ (.A(_12460_),
    .X(_12521_));
 sg13g2_nand2_1 _19470_ (.Y(_12522_),
    .A(net702),
    .B(\mem.mem_internal.code_mem[194][2] ));
 sg13g2_nand2_1 _19471_ (.Y(_12523_),
    .A(net1108),
    .B(_12516_));
 sg13g2_o21ai_1 _19472_ (.B1(_12523_),
    .Y(_00948_),
    .A1(net222),
    .A2(_12522_));
 sg13g2_nand2_1 _19473_ (.Y(_12524_),
    .A(_12521_),
    .B(\mem.mem_internal.code_mem[194][3] ));
 sg13g2_nand2_1 _19474_ (.Y(_12525_),
    .A(net1107),
    .B(_12516_));
 sg13g2_o21ai_1 _19475_ (.B1(_12525_),
    .Y(_00949_),
    .A1(net222),
    .A2(_12524_));
 sg13g2_nand2_1 _19476_ (.Y(_12526_),
    .A(net702),
    .B(\mem.mem_internal.code_mem[194][4] ));
 sg13g2_nand2_1 _19477_ (.Y(_12527_),
    .A(net1106),
    .B(_12516_));
 sg13g2_o21ai_1 _19478_ (.B1(_12527_),
    .Y(_00950_),
    .A1(_12517_),
    .A2(_12526_));
 sg13g2_nand2_1 _19479_ (.Y(_12528_),
    .A(net702),
    .B(\mem.mem_internal.code_mem[194][5] ));
 sg13g2_nand2_1 _19480_ (.Y(_12529_),
    .A(net1105),
    .B(_12516_));
 sg13g2_o21ai_1 _19481_ (.B1(_12529_),
    .Y(_00951_),
    .A1(net222),
    .A2(_12528_));
 sg13g2_nand2_1 _19482_ (.Y(_12530_),
    .A(net702),
    .B(\mem.mem_internal.code_mem[194][6] ));
 sg13g2_nand2_1 _19483_ (.Y(_12531_),
    .A(net1104),
    .B(_12516_));
 sg13g2_o21ai_1 _19484_ (.B1(_12531_),
    .Y(_00952_),
    .A1(_12517_),
    .A2(_12530_));
 sg13g2_nand2_1 _19485_ (.Y(_12532_),
    .A(net702),
    .B(\mem.mem_internal.code_mem[194][7] ));
 sg13g2_nand2_1 _19486_ (.Y(_12533_),
    .A(net1103),
    .B(_12516_));
 sg13g2_o21ai_1 _19487_ (.B1(_12533_),
    .Y(_00953_),
    .A1(net222),
    .A2(_12532_));
 sg13g2_nand2_1 _19488_ (.Y(_12534_),
    .A(net844),
    .B(\mem.mem_internal.code_mem[195][0] ));
 sg13g2_nor2_1 _19489_ (.A(net526),
    .B(net462),
    .Y(_12535_));
 sg13g2_buf_2 _19490_ (.A(_12535_),
    .X(_12536_));
 sg13g2_buf_1 _19491_ (.A(_12536_),
    .X(_12537_));
 sg13g2_nand2_1 _19492_ (.Y(_12538_),
    .A(net1110),
    .B(net221));
 sg13g2_o21ai_1 _19493_ (.B1(_12538_),
    .Y(_00954_),
    .A1(_12534_),
    .A2(net221));
 sg13g2_nand2_1 _19494_ (.Y(_12539_),
    .A(net702),
    .B(\mem.mem_internal.code_mem[195][1] ));
 sg13g2_nand2_1 _19495_ (.Y(_12540_),
    .A(net1109),
    .B(net221));
 sg13g2_o21ai_1 _19496_ (.B1(_12540_),
    .Y(_00955_),
    .A1(net221),
    .A2(_12539_));
 sg13g2_nand2_1 _19497_ (.Y(_12541_),
    .A(net702),
    .B(\mem.mem_internal.code_mem[195][2] ));
 sg13g2_nand2_1 _19498_ (.Y(_12542_),
    .A(net1108),
    .B(_12536_));
 sg13g2_o21ai_1 _19499_ (.B1(_12542_),
    .Y(_00956_),
    .A1(net221),
    .A2(_12541_));
 sg13g2_nand2_1 _19500_ (.Y(_12543_),
    .A(_12521_),
    .B(\mem.mem_internal.code_mem[195][3] ));
 sg13g2_nand2_1 _19501_ (.Y(_12544_),
    .A(net1107),
    .B(_12536_));
 sg13g2_o21ai_1 _19502_ (.B1(_12544_),
    .Y(_00957_),
    .A1(net221),
    .A2(_12543_));
 sg13g2_nand2_1 _19503_ (.Y(_12545_),
    .A(net702),
    .B(\mem.mem_internal.code_mem[195][4] ));
 sg13g2_nand2_1 _19504_ (.Y(_12546_),
    .A(net1106),
    .B(_12536_));
 sg13g2_o21ai_1 _19505_ (.B1(_12546_),
    .Y(_00958_),
    .A1(_12537_),
    .A2(_12545_));
 sg13g2_buf_1 _19506_ (.A(_12460_),
    .X(_12547_));
 sg13g2_nand2_1 _19507_ (.Y(_12548_),
    .A(net701),
    .B(\mem.mem_internal.code_mem[195][5] ));
 sg13g2_nand2_1 _19508_ (.Y(_12549_),
    .A(net1105),
    .B(_12536_));
 sg13g2_o21ai_1 _19509_ (.B1(_12549_),
    .Y(_00959_),
    .A1(net221),
    .A2(_12548_));
 sg13g2_nand2_1 _19510_ (.Y(_12550_),
    .A(_12547_),
    .B(\mem.mem_internal.code_mem[195][6] ));
 sg13g2_nand2_1 _19511_ (.Y(_12551_),
    .A(net1104),
    .B(_12536_));
 sg13g2_o21ai_1 _19512_ (.B1(_12551_),
    .Y(_00960_),
    .A1(_12537_),
    .A2(_12550_));
 sg13g2_nand2_1 _19513_ (.Y(_12552_),
    .A(net701),
    .B(\mem.mem_internal.code_mem[195][7] ));
 sg13g2_nand2_1 _19514_ (.Y(_12553_),
    .A(net1103),
    .B(_12536_));
 sg13g2_o21ai_1 _19515_ (.B1(_12553_),
    .Y(_00961_),
    .A1(net221),
    .A2(_12552_));
 sg13g2_nand2_1 _19516_ (.Y(_12554_),
    .A(net844),
    .B(\mem.mem_internal.code_mem[196][0] ));
 sg13g2_nor2_1 _19517_ (.A(_10296_),
    .B(net462),
    .Y(_12555_));
 sg13g2_buf_2 _19518_ (.A(_12555_),
    .X(_12556_));
 sg13g2_buf_1 _19519_ (.A(_12556_),
    .X(_12557_));
 sg13g2_nand2_1 _19520_ (.Y(_12558_),
    .A(net1110),
    .B(net220));
 sg13g2_o21ai_1 _19521_ (.B1(_12558_),
    .Y(_00962_),
    .A1(_12554_),
    .A2(net220));
 sg13g2_nand2_1 _19522_ (.Y(_12559_),
    .A(_12547_),
    .B(\mem.mem_internal.code_mem[196][1] ));
 sg13g2_nand2_1 _19523_ (.Y(_12560_),
    .A(net1109),
    .B(net220));
 sg13g2_o21ai_1 _19524_ (.B1(_12560_),
    .Y(_00963_),
    .A1(net220),
    .A2(_12559_));
 sg13g2_nand2_1 _19525_ (.Y(_12561_),
    .A(net701),
    .B(\mem.mem_internal.code_mem[196][2] ));
 sg13g2_nand2_1 _19526_ (.Y(_12562_),
    .A(net1108),
    .B(_12556_));
 sg13g2_o21ai_1 _19527_ (.B1(_12562_),
    .Y(_00964_),
    .A1(_12557_),
    .A2(_12561_));
 sg13g2_nand2_1 _19528_ (.Y(_12563_),
    .A(net701),
    .B(\mem.mem_internal.code_mem[196][3] ));
 sg13g2_nand2_1 _19529_ (.Y(_12564_),
    .A(net1107),
    .B(_12556_));
 sg13g2_o21ai_1 _19530_ (.B1(_12564_),
    .Y(_00965_),
    .A1(_12557_),
    .A2(_12563_));
 sg13g2_nand2_1 _19531_ (.Y(_12565_),
    .A(net701),
    .B(\mem.mem_internal.code_mem[196][4] ));
 sg13g2_nand2_1 _19532_ (.Y(_12566_),
    .A(net1106),
    .B(_12556_));
 sg13g2_o21ai_1 _19533_ (.B1(_12566_),
    .Y(_00966_),
    .A1(net220),
    .A2(_12565_));
 sg13g2_nand2_1 _19534_ (.Y(_12567_),
    .A(net701),
    .B(\mem.mem_internal.code_mem[196][5] ));
 sg13g2_nand2_1 _19535_ (.Y(_12568_),
    .A(net1105),
    .B(_12556_));
 sg13g2_o21ai_1 _19536_ (.B1(_12568_),
    .Y(_00967_),
    .A1(net220),
    .A2(_12567_));
 sg13g2_nand2_1 _19537_ (.Y(_12569_),
    .A(net701),
    .B(\mem.mem_internal.code_mem[196][6] ));
 sg13g2_nand2_1 _19538_ (.Y(_12570_),
    .A(net1104),
    .B(_12556_));
 sg13g2_o21ai_1 _19539_ (.B1(_12570_),
    .Y(_00968_),
    .A1(net220),
    .A2(_12569_));
 sg13g2_nand2_1 _19540_ (.Y(_12571_),
    .A(net701),
    .B(\mem.mem_internal.code_mem[196][7] ));
 sg13g2_nand2_1 _19541_ (.Y(_12572_),
    .A(net1103),
    .B(_12556_));
 sg13g2_o21ai_1 _19542_ (.B1(_12572_),
    .Y(_00969_),
    .A1(net220),
    .A2(_12571_));
 sg13g2_nand2_1 _19543_ (.Y(_12573_),
    .A(net844),
    .B(\mem.mem_internal.code_mem[197][0] ));
 sg13g2_nor2_1 _19544_ (.A(_10326_),
    .B(net462),
    .Y(_12574_));
 sg13g2_buf_2 _19545_ (.A(_12574_),
    .X(_12575_));
 sg13g2_buf_1 _19546_ (.A(_12575_),
    .X(_12576_));
 sg13g2_nand2_1 _19547_ (.Y(_12577_),
    .A(net1110),
    .B(net219));
 sg13g2_o21ai_1 _19548_ (.B1(_12577_),
    .Y(_00970_),
    .A1(_12573_),
    .A2(net219));
 sg13g2_buf_1 _19549_ (.A(_12460_),
    .X(_12578_));
 sg13g2_nand2_1 _19550_ (.Y(_12579_),
    .A(net700),
    .B(\mem.mem_internal.code_mem[197][1] ));
 sg13g2_nand2_1 _19551_ (.Y(_12580_),
    .A(net1109),
    .B(net219));
 sg13g2_o21ai_1 _19552_ (.B1(_12580_),
    .Y(_00971_),
    .A1(net219),
    .A2(_12579_));
 sg13g2_nand2_1 _19553_ (.Y(_12581_),
    .A(net700),
    .B(\mem.mem_internal.code_mem[197][2] ));
 sg13g2_nand2_1 _19554_ (.Y(_12582_),
    .A(net1108),
    .B(_12575_));
 sg13g2_o21ai_1 _19555_ (.B1(_12582_),
    .Y(_00972_),
    .A1(_12576_),
    .A2(_12581_));
 sg13g2_nand2_1 _19556_ (.Y(_12583_),
    .A(net700),
    .B(\mem.mem_internal.code_mem[197][3] ));
 sg13g2_nand2_1 _19557_ (.Y(_12584_),
    .A(net1107),
    .B(_12575_));
 sg13g2_o21ai_1 _19558_ (.B1(_12584_),
    .Y(_00973_),
    .A1(_12576_),
    .A2(_12583_));
 sg13g2_nand2_1 _19559_ (.Y(_12585_),
    .A(net700),
    .B(\mem.mem_internal.code_mem[197][4] ));
 sg13g2_nand2_1 _19560_ (.Y(_12586_),
    .A(net1106),
    .B(_12575_));
 sg13g2_o21ai_1 _19561_ (.B1(_12586_),
    .Y(_00974_),
    .A1(net219),
    .A2(_12585_));
 sg13g2_nand2_1 _19562_ (.Y(_12587_),
    .A(net700),
    .B(\mem.mem_internal.code_mem[197][5] ));
 sg13g2_nand2_1 _19563_ (.Y(_12588_),
    .A(net1105),
    .B(_12575_));
 sg13g2_o21ai_1 _19564_ (.B1(_12588_),
    .Y(_00975_),
    .A1(net219),
    .A2(_12587_));
 sg13g2_nand2_1 _19565_ (.Y(_12589_),
    .A(net700),
    .B(\mem.mem_internal.code_mem[197][6] ));
 sg13g2_nand2_1 _19566_ (.Y(_12590_),
    .A(net1104),
    .B(_12575_));
 sg13g2_o21ai_1 _19567_ (.B1(_12590_),
    .Y(_00976_),
    .A1(net219),
    .A2(_12589_));
 sg13g2_nand2_1 _19568_ (.Y(_12591_),
    .A(net700),
    .B(\mem.mem_internal.code_mem[197][7] ));
 sg13g2_nand2_1 _19569_ (.Y(_12592_),
    .A(net1103),
    .B(_12575_));
 sg13g2_o21ai_1 _19570_ (.B1(_12592_),
    .Y(_00977_),
    .A1(net219),
    .A2(_12591_));
 sg13g2_nand2_1 _19571_ (.Y(_12593_),
    .A(_12403_),
    .B(\mem.mem_internal.code_mem[198][0] ));
 sg13g2_nor2_1 _19572_ (.A(net779),
    .B(net462),
    .Y(_12594_));
 sg13g2_buf_2 _19573_ (.A(_12594_),
    .X(_12595_));
 sg13g2_buf_1 _19574_ (.A(_12595_),
    .X(_12596_));
 sg13g2_nand2_1 _19575_ (.Y(_12597_),
    .A(_12427_),
    .B(net218));
 sg13g2_o21ai_1 _19576_ (.B1(_12597_),
    .Y(_00978_),
    .A1(_12593_),
    .A2(net218));
 sg13g2_nand2_1 _19577_ (.Y(_12598_),
    .A(_12578_),
    .B(\mem.mem_internal.code_mem[198][1] ));
 sg13g2_nand2_1 _19578_ (.Y(_12599_),
    .A(_12431_),
    .B(net218));
 sg13g2_o21ai_1 _19579_ (.B1(_12599_),
    .Y(_00979_),
    .A1(net218),
    .A2(_12598_));
 sg13g2_nand2_1 _19580_ (.Y(_12600_),
    .A(_12578_),
    .B(\mem.mem_internal.code_mem[198][2] ));
 sg13g2_nand2_1 _19581_ (.Y(_12601_),
    .A(_12434_),
    .B(_12595_));
 sg13g2_o21ai_1 _19582_ (.B1(_12601_),
    .Y(_00980_),
    .A1(_12596_),
    .A2(_12600_));
 sg13g2_nand2_1 _19583_ (.Y(_12602_),
    .A(net700),
    .B(\mem.mem_internal.code_mem[198][3] ));
 sg13g2_nand2_1 _19584_ (.Y(_12603_),
    .A(_12437_),
    .B(_12595_));
 sg13g2_o21ai_1 _19585_ (.B1(_12603_),
    .Y(_00981_),
    .A1(_12596_),
    .A2(_12602_));
 sg13g2_buf_1 _19586_ (.A(_12460_),
    .X(_12604_));
 sg13g2_nand2_1 _19587_ (.Y(_12605_),
    .A(net699),
    .B(\mem.mem_internal.code_mem[198][4] ));
 sg13g2_nand2_1 _19588_ (.Y(_12606_),
    .A(_12440_),
    .B(_12595_));
 sg13g2_o21ai_1 _19589_ (.B1(_12606_),
    .Y(_00982_),
    .A1(net218),
    .A2(_12605_));
 sg13g2_nand2_1 _19590_ (.Y(_12607_),
    .A(net699),
    .B(\mem.mem_internal.code_mem[198][5] ));
 sg13g2_nand2_1 _19591_ (.Y(_12608_),
    .A(_12443_),
    .B(_12595_));
 sg13g2_o21ai_1 _19592_ (.B1(_12608_),
    .Y(_00983_),
    .A1(net218),
    .A2(_12607_));
 sg13g2_nand2_1 _19593_ (.Y(_12609_),
    .A(net699),
    .B(\mem.mem_internal.code_mem[198][6] ));
 sg13g2_nand2_1 _19594_ (.Y(_12610_),
    .A(_12446_),
    .B(_12595_));
 sg13g2_o21ai_1 _19595_ (.B1(_12610_),
    .Y(_00984_),
    .A1(net218),
    .A2(_12609_));
 sg13g2_nand2_1 _19596_ (.Y(_12611_),
    .A(net699),
    .B(\mem.mem_internal.code_mem[198][7] ));
 sg13g2_nand2_1 _19597_ (.Y(_12612_),
    .A(_12449_),
    .B(_12595_));
 sg13g2_o21ai_1 _19598_ (.B1(_12612_),
    .Y(_00985_),
    .A1(net218),
    .A2(_12611_));
 sg13g2_nand2_1 _19599_ (.Y(_12613_),
    .A(_12403_),
    .B(\mem.mem_internal.code_mem[199][0] ));
 sg13g2_nor2_1 _19600_ (.A(_10373_),
    .B(net462),
    .Y(_12614_));
 sg13g2_buf_2 _19601_ (.A(_12614_),
    .X(_12615_));
 sg13g2_buf_1 _19602_ (.A(_12615_),
    .X(_12616_));
 sg13g2_nand2_1 _19603_ (.Y(_12617_),
    .A(_12427_),
    .B(net217));
 sg13g2_o21ai_1 _19604_ (.B1(_12617_),
    .Y(_00986_),
    .A1(_12613_),
    .A2(net217));
 sg13g2_nand2_1 _19605_ (.Y(_12618_),
    .A(_12604_),
    .B(\mem.mem_internal.code_mem[199][1] ));
 sg13g2_nand2_1 _19606_ (.Y(_12619_),
    .A(_12431_),
    .B(net217));
 sg13g2_o21ai_1 _19607_ (.B1(_12619_),
    .Y(_00987_),
    .A1(net217),
    .A2(_12618_));
 sg13g2_nand2_1 _19608_ (.Y(_12620_),
    .A(_12604_),
    .B(\mem.mem_internal.code_mem[199][2] ));
 sg13g2_nand2_1 _19609_ (.Y(_12621_),
    .A(_12434_),
    .B(_12615_));
 sg13g2_o21ai_1 _19610_ (.B1(_12621_),
    .Y(_00988_),
    .A1(net217),
    .A2(_12620_));
 sg13g2_nand2_1 _19611_ (.Y(_12622_),
    .A(net699),
    .B(\mem.mem_internal.code_mem[199][3] ));
 sg13g2_nand2_1 _19612_ (.Y(_12623_),
    .A(_12437_),
    .B(_12615_));
 sg13g2_o21ai_1 _19613_ (.B1(_12623_),
    .Y(_00989_),
    .A1(_12616_),
    .A2(_12622_));
 sg13g2_nand2_1 _19614_ (.Y(_12624_),
    .A(net699),
    .B(\mem.mem_internal.code_mem[199][4] ));
 sg13g2_nand2_1 _19615_ (.Y(_12625_),
    .A(_12440_),
    .B(_12615_));
 sg13g2_o21ai_1 _19616_ (.B1(_12625_),
    .Y(_00990_),
    .A1(_12616_),
    .A2(_12624_));
 sg13g2_nand2_1 _19617_ (.Y(_12626_),
    .A(net699),
    .B(\mem.mem_internal.code_mem[199][5] ));
 sg13g2_nand2_1 _19618_ (.Y(_12627_),
    .A(_12443_),
    .B(_12615_));
 sg13g2_o21ai_1 _19619_ (.B1(_12627_),
    .Y(_00991_),
    .A1(net217),
    .A2(_12626_));
 sg13g2_nand2_1 _19620_ (.Y(_12628_),
    .A(net699),
    .B(\mem.mem_internal.code_mem[199][6] ));
 sg13g2_nand2_1 _19621_ (.Y(_12629_),
    .A(_12446_),
    .B(_12615_));
 sg13g2_o21ai_1 _19622_ (.B1(_12629_),
    .Y(_00992_),
    .A1(net217),
    .A2(_12628_));
 sg13g2_buf_1 _19623_ (.A(_12460_),
    .X(_12630_));
 sg13g2_nand2_1 _19624_ (.Y(_12631_),
    .A(_12630_),
    .B(\mem.mem_internal.code_mem[199][7] ));
 sg13g2_nand2_1 _19625_ (.Y(_12632_),
    .A(_12449_),
    .B(_12615_));
 sg13g2_o21ai_1 _19626_ (.B1(_12632_),
    .Y(_00993_),
    .A1(net217),
    .A2(_12631_));
 sg13g2_nand2_1 _19627_ (.Y(_12633_),
    .A(net844),
    .B(\mem.mem_internal.code_mem[19][0] ));
 sg13g2_nor2_1 _19628_ (.A(_10679_),
    .B(net464),
    .Y(_12634_));
 sg13g2_buf_2 _19629_ (.A(_12634_),
    .X(_12635_));
 sg13g2_buf_1 _19630_ (.A(_12635_),
    .X(_12636_));
 sg13g2_buf_1 _19631_ (.A(_10251_),
    .X(_12637_));
 sg13g2_buf_1 _19632_ (.A(_12637_),
    .X(_12638_));
 sg13g2_nand2_1 _19633_ (.Y(_12639_),
    .A(net1102),
    .B(net216));
 sg13g2_o21ai_1 _19634_ (.B1(_12639_),
    .Y(_00994_),
    .A1(_12633_),
    .A2(net216));
 sg13g2_nand2_1 _19635_ (.Y(_12640_),
    .A(net698),
    .B(\mem.mem_internal.code_mem[19][1] ));
 sg13g2_buf_1 _19636_ (.A(_10256_),
    .X(_12641_));
 sg13g2_buf_1 _19637_ (.A(_12641_),
    .X(_12642_));
 sg13g2_nand2_1 _19638_ (.Y(_12643_),
    .A(net1101),
    .B(net216));
 sg13g2_o21ai_1 _19639_ (.B1(_12643_),
    .Y(_00995_),
    .A1(net216),
    .A2(_12640_));
 sg13g2_nand2_1 _19640_ (.Y(_12644_),
    .A(net698),
    .B(\mem.mem_internal.code_mem[19][2] ));
 sg13g2_buf_1 _19641_ (.A(_10262_),
    .X(_12645_));
 sg13g2_buf_1 _19642_ (.A(_12645_),
    .X(_12646_));
 sg13g2_nand2_1 _19643_ (.Y(_12647_),
    .A(net1100),
    .B(_12635_));
 sg13g2_o21ai_1 _19644_ (.B1(_12647_),
    .Y(_00996_),
    .A1(net216),
    .A2(_12644_));
 sg13g2_nand2_1 _19645_ (.Y(_12648_),
    .A(net698),
    .B(\mem.mem_internal.code_mem[19][3] ));
 sg13g2_buf_2 _19646_ (.A(_10267_),
    .X(_12649_));
 sg13g2_buf_1 _19647_ (.A(_12649_),
    .X(_12650_));
 sg13g2_nand2_1 _19648_ (.Y(_12651_),
    .A(net1099),
    .B(_12635_));
 sg13g2_o21ai_1 _19649_ (.B1(_12651_),
    .Y(_00997_),
    .A1(net216),
    .A2(_12648_));
 sg13g2_nand2_1 _19650_ (.Y(_12652_),
    .A(net698),
    .B(\mem.mem_internal.code_mem[19][4] ));
 sg13g2_buf_2 _19651_ (.A(_10272_),
    .X(_12653_));
 sg13g2_buf_1 _19652_ (.A(_12653_),
    .X(_12654_));
 sg13g2_nand2_1 _19653_ (.Y(_12655_),
    .A(net1098),
    .B(_12635_));
 sg13g2_o21ai_1 _19654_ (.B1(_12655_),
    .Y(_00998_),
    .A1(_12636_),
    .A2(_12652_));
 sg13g2_nand2_1 _19655_ (.Y(_12656_),
    .A(net698),
    .B(\mem.mem_internal.code_mem[19][5] ));
 sg13g2_buf_2 _19656_ (.A(_10277_),
    .X(_12657_));
 sg13g2_buf_1 _19657_ (.A(_12657_),
    .X(_12658_));
 sg13g2_nand2_1 _19658_ (.Y(_12659_),
    .A(net1097),
    .B(_12635_));
 sg13g2_o21ai_1 _19659_ (.B1(_12659_),
    .Y(_00999_),
    .A1(net216),
    .A2(_12656_));
 sg13g2_nand2_1 _19660_ (.Y(_12660_),
    .A(net698),
    .B(\mem.mem_internal.code_mem[19][6] ));
 sg13g2_buf_2 _19661_ (.A(_10282_),
    .X(_12661_));
 sg13g2_buf_1 _19662_ (.A(_12661_),
    .X(_12662_));
 sg13g2_nand2_1 _19663_ (.Y(_12663_),
    .A(net1096),
    .B(_12635_));
 sg13g2_o21ai_1 _19664_ (.B1(_12663_),
    .Y(_01000_),
    .A1(_12636_),
    .A2(_12660_));
 sg13g2_nand2_1 _19665_ (.Y(_12664_),
    .A(net698),
    .B(\mem.mem_internal.code_mem[19][7] ));
 sg13g2_buf_1 _19666_ (.A(_10287_),
    .X(_12665_));
 sg13g2_buf_1 _19667_ (.A(_12665_),
    .X(_12666_));
 sg13g2_nand2_1 _19668_ (.Y(_12667_),
    .A(net1095),
    .B(_12635_));
 sg13g2_o21ai_1 _19669_ (.B1(_12667_),
    .Y(_01001_),
    .A1(net216),
    .A2(_12664_));
 sg13g2_buf_1 _19670_ (.A(_11058_),
    .X(_12668_));
 sg13g2_nand2_1 _19671_ (.Y(_12669_),
    .A(_12668_),
    .B(\mem.mem_internal.code_mem[1][0] ));
 sg13g2_nor2_1 _19672_ (.A(_10247_),
    .B(net528),
    .Y(_12670_));
 sg13g2_buf_2 _19673_ (.A(_12670_),
    .X(_12671_));
 sg13g2_buf_1 _19674_ (.A(_12671_),
    .X(_12672_));
 sg13g2_nand2_1 _19675_ (.Y(_12673_),
    .A(net1102),
    .B(net215));
 sg13g2_o21ai_1 _19676_ (.B1(_12673_),
    .Y(_01002_),
    .A1(_12669_),
    .A2(net215));
 sg13g2_nand2_1 _19677_ (.Y(_12674_),
    .A(net698),
    .B(\mem.mem_internal.code_mem[1][1] ));
 sg13g2_nand2_1 _19678_ (.Y(_12675_),
    .A(net1101),
    .B(net215));
 sg13g2_o21ai_1 _19679_ (.B1(_12675_),
    .Y(_01003_),
    .A1(net215),
    .A2(_12674_));
 sg13g2_nand2_1 _19680_ (.Y(_12676_),
    .A(_12630_),
    .B(\mem.mem_internal.code_mem[1][2] ));
 sg13g2_nand2_1 _19681_ (.Y(_12677_),
    .A(net1100),
    .B(_12671_));
 sg13g2_o21ai_1 _19682_ (.B1(_12677_),
    .Y(_01004_),
    .A1(net215),
    .A2(_12676_));
 sg13g2_buf_1 _19683_ (.A(_11875_),
    .X(_12678_));
 sg13g2_buf_1 _19684_ (.A(_12678_),
    .X(_12679_));
 sg13g2_nand2_1 _19685_ (.Y(_12680_),
    .A(net697),
    .B(\mem.mem_internal.code_mem[1][3] ));
 sg13g2_nand2_1 _19686_ (.Y(_12681_),
    .A(net1099),
    .B(_12671_));
 sg13g2_o21ai_1 _19687_ (.B1(_12681_),
    .Y(_01005_),
    .A1(net215),
    .A2(_12680_));
 sg13g2_nand2_1 _19688_ (.Y(_12682_),
    .A(net697),
    .B(\mem.mem_internal.code_mem[1][4] ));
 sg13g2_nand2_1 _19689_ (.Y(_12683_),
    .A(net1098),
    .B(_12671_));
 sg13g2_o21ai_1 _19690_ (.B1(_12683_),
    .Y(_01006_),
    .A1(net215),
    .A2(_12682_));
 sg13g2_nand2_1 _19691_ (.Y(_12684_),
    .A(net697),
    .B(\mem.mem_internal.code_mem[1][5] ));
 sg13g2_nand2_1 _19692_ (.Y(_12685_),
    .A(net1097),
    .B(_12671_));
 sg13g2_o21ai_1 _19693_ (.B1(_12685_),
    .Y(_01007_),
    .A1(net215),
    .A2(_12684_));
 sg13g2_nand2_1 _19694_ (.Y(_12686_),
    .A(net697),
    .B(\mem.mem_internal.code_mem[1][6] ));
 sg13g2_nand2_1 _19695_ (.Y(_12687_),
    .A(net1096),
    .B(_12671_));
 sg13g2_o21ai_1 _19696_ (.B1(_12687_),
    .Y(_01008_),
    .A1(_12672_),
    .A2(_12686_));
 sg13g2_nand2_1 _19697_ (.Y(_12688_),
    .A(net697),
    .B(\mem.mem_internal.code_mem[1][7] ));
 sg13g2_nand2_1 _19698_ (.Y(_12689_),
    .A(net1095),
    .B(_12671_));
 sg13g2_o21ai_1 _19699_ (.B1(_12689_),
    .Y(_01009_),
    .A1(_12672_),
    .A2(_12688_));
 sg13g2_nand2_1 _19700_ (.Y(_12690_),
    .A(net843),
    .B(\mem.mem_internal.code_mem[200][0] ));
 sg13g2_nor2_1 _19701_ (.A(_10398_),
    .B(_12475_),
    .Y(_12691_));
 sg13g2_buf_2 _19702_ (.A(_12691_),
    .X(_12692_));
 sg13g2_buf_1 _19703_ (.A(_12692_),
    .X(_12693_));
 sg13g2_nand2_1 _19704_ (.Y(_12694_),
    .A(net1102),
    .B(net214));
 sg13g2_o21ai_1 _19705_ (.B1(_12694_),
    .Y(_01010_),
    .A1(_12690_),
    .A2(net214));
 sg13g2_nand2_1 _19706_ (.Y(_12695_),
    .A(net697),
    .B(\mem.mem_internal.code_mem[200][1] ));
 sg13g2_nand2_1 _19707_ (.Y(_12696_),
    .A(net1101),
    .B(net214));
 sg13g2_o21ai_1 _19708_ (.B1(_12696_),
    .Y(_01011_),
    .A1(net214),
    .A2(_12695_));
 sg13g2_nand2_1 _19709_ (.Y(_12697_),
    .A(net697),
    .B(\mem.mem_internal.code_mem[200][2] ));
 sg13g2_nand2_1 _19710_ (.Y(_12698_),
    .A(net1100),
    .B(_12692_));
 sg13g2_o21ai_1 _19711_ (.B1(_12698_),
    .Y(_01012_),
    .A1(net214),
    .A2(_12697_));
 sg13g2_nand2_1 _19712_ (.Y(_12699_),
    .A(net697),
    .B(\mem.mem_internal.code_mem[200][3] ));
 sg13g2_nand2_1 _19713_ (.Y(_12700_),
    .A(net1099),
    .B(_12692_));
 sg13g2_o21ai_1 _19714_ (.B1(_12700_),
    .Y(_01013_),
    .A1(net214),
    .A2(_12699_));
 sg13g2_nand2_1 _19715_ (.Y(_12701_),
    .A(_12679_),
    .B(\mem.mem_internal.code_mem[200][4] ));
 sg13g2_nand2_1 _19716_ (.Y(_12702_),
    .A(net1098),
    .B(_12692_));
 sg13g2_o21ai_1 _19717_ (.B1(_12702_),
    .Y(_01014_),
    .A1(net214),
    .A2(_12701_));
 sg13g2_nand2_1 _19718_ (.Y(_12703_),
    .A(_12679_),
    .B(\mem.mem_internal.code_mem[200][5] ));
 sg13g2_nand2_1 _19719_ (.Y(_12704_),
    .A(net1097),
    .B(_12692_));
 sg13g2_o21ai_1 _19720_ (.B1(_12704_),
    .Y(_01015_),
    .A1(net214),
    .A2(_12703_));
 sg13g2_buf_1 _19721_ (.A(_12678_),
    .X(_12705_));
 sg13g2_nand2_1 _19722_ (.Y(_12706_),
    .A(net696),
    .B(\mem.mem_internal.code_mem[200][6] ));
 sg13g2_nand2_1 _19723_ (.Y(_12707_),
    .A(net1096),
    .B(_12692_));
 sg13g2_o21ai_1 _19724_ (.B1(_12707_),
    .Y(_01016_),
    .A1(_12693_),
    .A2(_12706_));
 sg13g2_nand2_1 _19725_ (.Y(_12708_),
    .A(net696),
    .B(\mem.mem_internal.code_mem[200][7] ));
 sg13g2_nand2_1 _19726_ (.Y(_12709_),
    .A(net1095),
    .B(_12692_));
 sg13g2_o21ai_1 _19727_ (.B1(_12709_),
    .Y(_01017_),
    .A1(_12693_),
    .A2(_12708_));
 sg13g2_nand2_1 _19728_ (.Y(_12710_),
    .A(net843),
    .B(\mem.mem_internal.code_mem[201][0] ));
 sg13g2_nor2_1 _19729_ (.A(_10423_),
    .B(_12475_),
    .Y(_12711_));
 sg13g2_buf_2 _19730_ (.A(_12711_),
    .X(_12712_));
 sg13g2_buf_1 _19731_ (.A(_12712_),
    .X(_12713_));
 sg13g2_nand2_1 _19732_ (.Y(_12714_),
    .A(net1102),
    .B(net213));
 sg13g2_o21ai_1 _19733_ (.B1(_12714_),
    .Y(_01018_),
    .A1(_12710_),
    .A2(net213));
 sg13g2_nand2_1 _19734_ (.Y(_12715_),
    .A(net696),
    .B(\mem.mem_internal.code_mem[201][1] ));
 sg13g2_nand2_1 _19735_ (.Y(_12716_),
    .A(net1101),
    .B(net213));
 sg13g2_o21ai_1 _19736_ (.B1(_12716_),
    .Y(_01019_),
    .A1(net213),
    .A2(_12715_));
 sg13g2_nand2_1 _19737_ (.Y(_12717_),
    .A(net696),
    .B(\mem.mem_internal.code_mem[201][2] ));
 sg13g2_nand2_1 _19738_ (.Y(_12718_),
    .A(net1100),
    .B(_12712_));
 sg13g2_o21ai_1 _19739_ (.B1(_12718_),
    .Y(_01020_),
    .A1(net213),
    .A2(_12717_));
 sg13g2_nand2_1 _19740_ (.Y(_12719_),
    .A(net696),
    .B(\mem.mem_internal.code_mem[201][3] ));
 sg13g2_nand2_1 _19741_ (.Y(_12720_),
    .A(net1099),
    .B(_12712_));
 sg13g2_o21ai_1 _19742_ (.B1(_12720_),
    .Y(_01021_),
    .A1(net213),
    .A2(_12719_));
 sg13g2_nand2_1 _19743_ (.Y(_12721_),
    .A(net696),
    .B(\mem.mem_internal.code_mem[201][4] ));
 sg13g2_nand2_1 _19744_ (.Y(_12722_),
    .A(net1098),
    .B(_12712_));
 sg13g2_o21ai_1 _19745_ (.B1(_12722_),
    .Y(_01022_),
    .A1(net213),
    .A2(_12721_));
 sg13g2_nand2_1 _19746_ (.Y(_12723_),
    .A(_12705_),
    .B(\mem.mem_internal.code_mem[201][5] ));
 sg13g2_nand2_1 _19747_ (.Y(_12724_),
    .A(net1097),
    .B(_12712_));
 sg13g2_o21ai_1 _19748_ (.B1(_12724_),
    .Y(_01023_),
    .A1(net213),
    .A2(_12723_));
 sg13g2_nand2_1 _19749_ (.Y(_12725_),
    .A(net696),
    .B(\mem.mem_internal.code_mem[201][6] ));
 sg13g2_nand2_1 _19750_ (.Y(_12726_),
    .A(net1096),
    .B(_12712_));
 sg13g2_o21ai_1 _19751_ (.B1(_12726_),
    .Y(_01024_),
    .A1(_12713_),
    .A2(_12725_));
 sg13g2_nand2_1 _19752_ (.Y(_12727_),
    .A(_12705_),
    .B(\mem.mem_internal.code_mem[201][7] ));
 sg13g2_nand2_1 _19753_ (.Y(_12728_),
    .A(net1095),
    .B(_12712_));
 sg13g2_o21ai_1 _19754_ (.B1(_12728_),
    .Y(_01025_),
    .A1(_12713_),
    .A2(_12727_));
 sg13g2_nand2_1 _19755_ (.Y(_12729_),
    .A(net843),
    .B(\mem.mem_internal.code_mem[202][0] ));
 sg13g2_nor2_1 _19756_ (.A(_10445_),
    .B(_12474_),
    .Y(_12730_));
 sg13g2_buf_2 _19757_ (.A(_12730_),
    .X(_12731_));
 sg13g2_buf_1 _19758_ (.A(_12731_),
    .X(_12732_));
 sg13g2_nand2_1 _19759_ (.Y(_12733_),
    .A(net1102),
    .B(net366));
 sg13g2_o21ai_1 _19760_ (.B1(_12733_),
    .Y(_01026_),
    .A1(_12729_),
    .A2(net366));
 sg13g2_nand2_1 _19761_ (.Y(_12734_),
    .A(net696),
    .B(\mem.mem_internal.code_mem[202][1] ));
 sg13g2_nand2_1 _19762_ (.Y(_12735_),
    .A(net1101),
    .B(net366));
 sg13g2_o21ai_1 _19763_ (.B1(_12735_),
    .Y(_01027_),
    .A1(net366),
    .A2(_12734_));
 sg13g2_buf_1 _19764_ (.A(_12678_),
    .X(_12736_));
 sg13g2_nand2_1 _19765_ (.Y(_12737_),
    .A(net695),
    .B(\mem.mem_internal.code_mem[202][2] ));
 sg13g2_nand2_1 _19766_ (.Y(_12738_),
    .A(net1100),
    .B(_12731_));
 sg13g2_o21ai_1 _19767_ (.B1(_12738_),
    .Y(_01028_),
    .A1(net366),
    .A2(_12737_));
 sg13g2_nand2_1 _19768_ (.Y(_12739_),
    .A(net695),
    .B(\mem.mem_internal.code_mem[202][3] ));
 sg13g2_nand2_1 _19769_ (.Y(_12740_),
    .A(net1099),
    .B(_12731_));
 sg13g2_o21ai_1 _19770_ (.B1(_12740_),
    .Y(_01029_),
    .A1(net366),
    .A2(_12739_));
 sg13g2_nand2_1 _19771_ (.Y(_12741_),
    .A(net695),
    .B(\mem.mem_internal.code_mem[202][4] ));
 sg13g2_nand2_1 _19772_ (.Y(_12742_),
    .A(net1098),
    .B(_12731_));
 sg13g2_o21ai_1 _19773_ (.B1(_12742_),
    .Y(_01030_),
    .A1(net366),
    .A2(_12741_));
 sg13g2_nand2_1 _19774_ (.Y(_12743_),
    .A(_12736_),
    .B(\mem.mem_internal.code_mem[202][5] ));
 sg13g2_nand2_1 _19775_ (.Y(_12744_),
    .A(net1097),
    .B(_12731_));
 sg13g2_o21ai_1 _19776_ (.B1(_12744_),
    .Y(_01031_),
    .A1(net366),
    .A2(_12743_));
 sg13g2_nand2_1 _19777_ (.Y(_12745_),
    .A(net695),
    .B(\mem.mem_internal.code_mem[202][6] ));
 sg13g2_nand2_1 _19778_ (.Y(_12746_),
    .A(net1096),
    .B(_12731_));
 sg13g2_o21ai_1 _19779_ (.B1(_12746_),
    .Y(_01032_),
    .A1(_12732_),
    .A2(_12745_));
 sg13g2_nand2_1 _19780_ (.Y(_12747_),
    .A(net695),
    .B(\mem.mem_internal.code_mem[202][7] ));
 sg13g2_nand2_1 _19781_ (.Y(_12748_),
    .A(net1095),
    .B(_12731_));
 sg13g2_o21ai_1 _19782_ (.B1(_12748_),
    .Y(_01033_),
    .A1(_12732_),
    .A2(_12747_));
 sg13g2_nand2_1 _19783_ (.Y(_12749_),
    .A(net843),
    .B(\mem.mem_internal.code_mem[203][0] ));
 sg13g2_nor2_1 _19784_ (.A(_10468_),
    .B(_12474_),
    .Y(_12750_));
 sg13g2_buf_2 _19785_ (.A(_12750_),
    .X(_12751_));
 sg13g2_buf_1 _19786_ (.A(_12751_),
    .X(_12752_));
 sg13g2_nand2_1 _19787_ (.Y(_12753_),
    .A(net1102),
    .B(net365));
 sg13g2_o21ai_1 _19788_ (.B1(_12753_),
    .Y(_01034_),
    .A1(_12749_),
    .A2(net365));
 sg13g2_nand2_1 _19789_ (.Y(_12754_),
    .A(net695),
    .B(\mem.mem_internal.code_mem[203][1] ));
 sg13g2_nand2_1 _19790_ (.Y(_12755_),
    .A(net1101),
    .B(net365));
 sg13g2_o21ai_1 _19791_ (.B1(_12755_),
    .Y(_01035_),
    .A1(net365),
    .A2(_12754_));
 sg13g2_nand2_1 _19792_ (.Y(_12756_),
    .A(net695),
    .B(\mem.mem_internal.code_mem[203][2] ));
 sg13g2_nand2_1 _19793_ (.Y(_12757_),
    .A(net1100),
    .B(_12751_));
 sg13g2_o21ai_1 _19794_ (.B1(_12757_),
    .Y(_01036_),
    .A1(net365),
    .A2(_12756_));
 sg13g2_nand2_1 _19795_ (.Y(_12758_),
    .A(_12736_),
    .B(\mem.mem_internal.code_mem[203][3] ));
 sg13g2_nand2_1 _19796_ (.Y(_12759_),
    .A(net1099),
    .B(_12751_));
 sg13g2_o21ai_1 _19797_ (.B1(_12759_),
    .Y(_01037_),
    .A1(net365),
    .A2(_12758_));
 sg13g2_nand2_1 _19798_ (.Y(_12760_),
    .A(net695),
    .B(\mem.mem_internal.code_mem[203][4] ));
 sg13g2_nand2_1 _19799_ (.Y(_12761_),
    .A(net1098),
    .B(_12751_));
 sg13g2_o21ai_1 _19800_ (.B1(_12761_),
    .Y(_01038_),
    .A1(net365),
    .A2(_12760_));
 sg13g2_buf_1 _19801_ (.A(_12678_),
    .X(_12762_));
 sg13g2_nand2_1 _19802_ (.Y(_12763_),
    .A(_12762_),
    .B(\mem.mem_internal.code_mem[203][5] ));
 sg13g2_nand2_1 _19803_ (.Y(_12764_),
    .A(net1097),
    .B(_12751_));
 sg13g2_o21ai_1 _19804_ (.B1(_12764_),
    .Y(_01039_),
    .A1(net365),
    .A2(_12763_));
 sg13g2_nand2_1 _19805_ (.Y(_12765_),
    .A(_12762_),
    .B(\mem.mem_internal.code_mem[203][6] ));
 sg13g2_nand2_1 _19806_ (.Y(_12766_),
    .A(net1096),
    .B(_12751_));
 sg13g2_o21ai_1 _19807_ (.B1(_12766_),
    .Y(_01040_),
    .A1(_12752_),
    .A2(_12765_));
 sg13g2_nand2_1 _19808_ (.Y(_12767_),
    .A(net694),
    .B(\mem.mem_internal.code_mem[203][7] ));
 sg13g2_nand2_1 _19809_ (.Y(_12768_),
    .A(net1095),
    .B(_12751_));
 sg13g2_o21ai_1 _19810_ (.B1(_12768_),
    .Y(_01041_),
    .A1(_12752_),
    .A2(_12767_));
 sg13g2_nand2_1 _19811_ (.Y(_12769_),
    .A(net843),
    .B(\mem.mem_internal.code_mem[204][0] ));
 sg13g2_nor2_1 _19812_ (.A(_10492_),
    .B(_12474_),
    .Y(_12770_));
 sg13g2_buf_2 _19813_ (.A(_12770_),
    .X(_12771_));
 sg13g2_buf_1 _19814_ (.A(_12771_),
    .X(_12772_));
 sg13g2_nand2_1 _19815_ (.Y(_12773_),
    .A(net1102),
    .B(net364));
 sg13g2_o21ai_1 _19816_ (.B1(_12773_),
    .Y(_01042_),
    .A1(_12769_),
    .A2(net364));
 sg13g2_nand2_1 _19817_ (.Y(_12774_),
    .A(net694),
    .B(\mem.mem_internal.code_mem[204][1] ));
 sg13g2_nand2_1 _19818_ (.Y(_12775_),
    .A(net1101),
    .B(net364));
 sg13g2_o21ai_1 _19819_ (.B1(_12775_),
    .Y(_01043_),
    .A1(net364),
    .A2(_12774_));
 sg13g2_nand2_1 _19820_ (.Y(_12776_),
    .A(net694),
    .B(\mem.mem_internal.code_mem[204][2] ));
 sg13g2_nand2_1 _19821_ (.Y(_12777_),
    .A(net1100),
    .B(_12771_));
 sg13g2_o21ai_1 _19822_ (.B1(_12777_),
    .Y(_01044_),
    .A1(net364),
    .A2(_12776_));
 sg13g2_nand2_1 _19823_ (.Y(_12778_),
    .A(net694),
    .B(\mem.mem_internal.code_mem[204][3] ));
 sg13g2_nand2_1 _19824_ (.Y(_12779_),
    .A(net1099),
    .B(_12771_));
 sg13g2_o21ai_1 _19825_ (.B1(_12779_),
    .Y(_01045_),
    .A1(_12772_),
    .A2(_12778_));
 sg13g2_nand2_1 _19826_ (.Y(_12780_),
    .A(net694),
    .B(\mem.mem_internal.code_mem[204][4] ));
 sg13g2_nand2_1 _19827_ (.Y(_12781_),
    .A(net1098),
    .B(_12771_));
 sg13g2_o21ai_1 _19828_ (.B1(_12781_),
    .Y(_01046_),
    .A1(_12772_),
    .A2(_12780_));
 sg13g2_nand2_1 _19829_ (.Y(_12782_),
    .A(net694),
    .B(\mem.mem_internal.code_mem[204][5] ));
 sg13g2_nand2_1 _19830_ (.Y(_12783_),
    .A(net1097),
    .B(_12771_));
 sg13g2_o21ai_1 _19831_ (.B1(_12783_),
    .Y(_01047_),
    .A1(net364),
    .A2(_12782_));
 sg13g2_nand2_1 _19832_ (.Y(_12784_),
    .A(net694),
    .B(\mem.mem_internal.code_mem[204][6] ));
 sg13g2_nand2_1 _19833_ (.Y(_12785_),
    .A(net1096),
    .B(_12771_));
 sg13g2_o21ai_1 _19834_ (.B1(_12785_),
    .Y(_01048_),
    .A1(net364),
    .A2(_12784_));
 sg13g2_nand2_1 _19835_ (.Y(_12786_),
    .A(net694),
    .B(\mem.mem_internal.code_mem[204][7] ));
 sg13g2_nand2_1 _19836_ (.Y(_12787_),
    .A(net1095),
    .B(_12771_));
 sg13g2_o21ai_1 _19837_ (.B1(_12787_),
    .Y(_01049_),
    .A1(net364),
    .A2(_12786_));
 sg13g2_nand2_1 _19838_ (.Y(_12788_),
    .A(net843),
    .B(\mem.mem_internal.code_mem[205][0] ));
 sg13g2_nor2_1 _19839_ (.A(_10514_),
    .B(_12474_),
    .Y(_12789_));
 sg13g2_buf_2 _19840_ (.A(_12789_),
    .X(_12790_));
 sg13g2_buf_1 _19841_ (.A(_12790_),
    .X(_12791_));
 sg13g2_nand2_1 _19842_ (.Y(_12792_),
    .A(net1102),
    .B(net363));
 sg13g2_o21ai_1 _19843_ (.B1(_12792_),
    .Y(_01050_),
    .A1(_12788_),
    .A2(net363));
 sg13g2_buf_1 _19844_ (.A(_12678_),
    .X(_12793_));
 sg13g2_nand2_1 _19845_ (.Y(_12794_),
    .A(net693),
    .B(\mem.mem_internal.code_mem[205][1] ));
 sg13g2_nand2_1 _19846_ (.Y(_12795_),
    .A(net1101),
    .B(net363));
 sg13g2_o21ai_1 _19847_ (.B1(_12795_),
    .Y(_01051_),
    .A1(net363),
    .A2(_12794_));
 sg13g2_nand2_1 _19848_ (.Y(_12796_),
    .A(net693),
    .B(\mem.mem_internal.code_mem[205][2] ));
 sg13g2_nand2_1 _19849_ (.Y(_12797_),
    .A(net1100),
    .B(_12790_));
 sg13g2_o21ai_1 _19850_ (.B1(_12797_),
    .Y(_01052_),
    .A1(net363),
    .A2(_12796_));
 sg13g2_nand2_1 _19851_ (.Y(_12798_),
    .A(net693),
    .B(\mem.mem_internal.code_mem[205][3] ));
 sg13g2_nand2_1 _19852_ (.Y(_12799_),
    .A(net1099),
    .B(_12790_));
 sg13g2_o21ai_1 _19853_ (.B1(_12799_),
    .Y(_01053_),
    .A1(net363),
    .A2(_12798_));
 sg13g2_nand2_1 _19854_ (.Y(_12800_),
    .A(_12793_),
    .B(\mem.mem_internal.code_mem[205][4] ));
 sg13g2_nand2_1 _19855_ (.Y(_12801_),
    .A(net1098),
    .B(_12790_));
 sg13g2_o21ai_1 _19856_ (.B1(_12801_),
    .Y(_01054_),
    .A1(net363),
    .A2(_12800_));
 sg13g2_nand2_1 _19857_ (.Y(_12802_),
    .A(net693),
    .B(\mem.mem_internal.code_mem[205][5] ));
 sg13g2_nand2_1 _19858_ (.Y(_12803_),
    .A(net1097),
    .B(_12790_));
 sg13g2_o21ai_1 _19859_ (.B1(_12803_),
    .Y(_01055_),
    .A1(_12791_),
    .A2(_12802_));
 sg13g2_nand2_1 _19860_ (.Y(_12804_),
    .A(net693),
    .B(\mem.mem_internal.code_mem[205][6] ));
 sg13g2_nand2_1 _19861_ (.Y(_12805_),
    .A(net1096),
    .B(_12790_));
 sg13g2_o21ai_1 _19862_ (.B1(_12805_),
    .Y(_01056_),
    .A1(net363),
    .A2(_12804_));
 sg13g2_nand2_1 _19863_ (.Y(_12806_),
    .A(net693),
    .B(\mem.mem_internal.code_mem[205][7] ));
 sg13g2_nand2_1 _19864_ (.Y(_12807_),
    .A(net1095),
    .B(_12790_));
 sg13g2_o21ai_1 _19865_ (.B1(_12807_),
    .Y(_01057_),
    .A1(_12791_),
    .A2(_12806_));
 sg13g2_nand2_1 _19866_ (.Y(_12808_),
    .A(net843),
    .B(\mem.mem_internal.code_mem[206][0] ));
 sg13g2_nor2_1 _19867_ (.A(_10565_),
    .B(_12474_),
    .Y(_12809_));
 sg13g2_buf_2 _19868_ (.A(_12809_),
    .X(_12810_));
 sg13g2_buf_1 _19869_ (.A(_12810_),
    .X(_12811_));
 sg13g2_nand2_1 _19870_ (.Y(_12812_),
    .A(_12638_),
    .B(net362));
 sg13g2_o21ai_1 _19871_ (.B1(_12812_),
    .Y(_01058_),
    .A1(_12808_),
    .A2(net362));
 sg13g2_nand2_1 _19872_ (.Y(_12813_),
    .A(net693),
    .B(\mem.mem_internal.code_mem[206][1] ));
 sg13g2_nand2_1 _19873_ (.Y(_12814_),
    .A(_12642_),
    .B(net362));
 sg13g2_o21ai_1 _19874_ (.B1(_12814_),
    .Y(_01059_),
    .A1(net362),
    .A2(_12813_));
 sg13g2_nand2_1 _19875_ (.Y(_12815_),
    .A(net693),
    .B(\mem.mem_internal.code_mem[206][2] ));
 sg13g2_nand2_1 _19876_ (.Y(_12816_),
    .A(_12646_),
    .B(_12810_));
 sg13g2_o21ai_1 _19877_ (.B1(_12816_),
    .Y(_01060_),
    .A1(net362),
    .A2(_12815_));
 sg13g2_nand2_1 _19878_ (.Y(_12817_),
    .A(_12793_),
    .B(\mem.mem_internal.code_mem[206][3] ));
 sg13g2_nand2_1 _19879_ (.Y(_12818_),
    .A(_12650_),
    .B(_12810_));
 sg13g2_o21ai_1 _19880_ (.B1(_12818_),
    .Y(_01061_),
    .A1(net362),
    .A2(_12817_));
 sg13g2_buf_1 _19881_ (.A(_12678_),
    .X(_12819_));
 sg13g2_nand2_1 _19882_ (.Y(_12820_),
    .A(_12819_),
    .B(\mem.mem_internal.code_mem[206][4] ));
 sg13g2_nand2_1 _19883_ (.Y(_12821_),
    .A(_12654_),
    .B(_12810_));
 sg13g2_o21ai_1 _19884_ (.B1(_12821_),
    .Y(_01062_),
    .A1(net362),
    .A2(_12820_));
 sg13g2_nand2_1 _19885_ (.Y(_12822_),
    .A(net692),
    .B(\mem.mem_internal.code_mem[206][5] ));
 sg13g2_nand2_1 _19886_ (.Y(_12823_),
    .A(_12658_),
    .B(_12810_));
 sg13g2_o21ai_1 _19887_ (.B1(_12823_),
    .Y(_01063_),
    .A1(_12811_),
    .A2(_12822_));
 sg13g2_nand2_1 _19888_ (.Y(_12824_),
    .A(net692),
    .B(\mem.mem_internal.code_mem[206][6] ));
 sg13g2_nand2_1 _19889_ (.Y(_12825_),
    .A(_12662_),
    .B(_12810_));
 sg13g2_o21ai_1 _19890_ (.B1(_12825_),
    .Y(_01064_),
    .A1(net362),
    .A2(_12824_));
 sg13g2_nand2_1 _19891_ (.Y(_12826_),
    .A(net692),
    .B(\mem.mem_internal.code_mem[206][7] ));
 sg13g2_nand2_1 _19892_ (.Y(_12827_),
    .A(_12666_),
    .B(_12810_));
 sg13g2_o21ai_1 _19893_ (.B1(_12827_),
    .Y(_01065_),
    .A1(_12811_),
    .A2(_12826_));
 sg13g2_nand2_1 _19894_ (.Y(_12828_),
    .A(_12668_),
    .B(\mem.mem_internal.code_mem[207][0] ));
 sg13g2_nor2_1 _19895_ (.A(_10587_),
    .B(_12474_),
    .Y(_12829_));
 sg13g2_buf_2 _19896_ (.A(_12829_),
    .X(_12830_));
 sg13g2_buf_1 _19897_ (.A(_12830_),
    .X(_12831_));
 sg13g2_nand2_1 _19898_ (.Y(_12832_),
    .A(_12638_),
    .B(net361));
 sg13g2_o21ai_1 _19899_ (.B1(_12832_),
    .Y(_01066_),
    .A1(_12828_),
    .A2(net361));
 sg13g2_nand2_1 _19900_ (.Y(_12833_),
    .A(net692),
    .B(\mem.mem_internal.code_mem[207][1] ));
 sg13g2_nand2_1 _19901_ (.Y(_12834_),
    .A(_12642_),
    .B(net361));
 sg13g2_o21ai_1 _19902_ (.B1(_12834_),
    .Y(_01067_),
    .A1(net361),
    .A2(_12833_));
 sg13g2_nand2_1 _19903_ (.Y(_12835_),
    .A(net692),
    .B(\mem.mem_internal.code_mem[207][2] ));
 sg13g2_nand2_1 _19904_ (.Y(_12836_),
    .A(_12646_),
    .B(_12830_));
 sg13g2_o21ai_1 _19905_ (.B1(_12836_),
    .Y(_01068_),
    .A1(net361),
    .A2(_12835_));
 sg13g2_nand2_1 _19906_ (.Y(_12837_),
    .A(net692),
    .B(\mem.mem_internal.code_mem[207][3] ));
 sg13g2_nand2_1 _19907_ (.Y(_12838_),
    .A(_12650_),
    .B(_12830_));
 sg13g2_o21ai_1 _19908_ (.B1(_12838_),
    .Y(_01069_),
    .A1(net361),
    .A2(_12837_));
 sg13g2_nand2_1 _19909_ (.Y(_12839_),
    .A(_12819_),
    .B(\mem.mem_internal.code_mem[207][4] ));
 sg13g2_nand2_1 _19910_ (.Y(_12840_),
    .A(_12654_),
    .B(_12830_));
 sg13g2_o21ai_1 _19911_ (.B1(_12840_),
    .Y(_01070_),
    .A1(_12831_),
    .A2(_12839_));
 sg13g2_nand2_1 _19912_ (.Y(_12841_),
    .A(net692),
    .B(\mem.mem_internal.code_mem[207][5] ));
 sg13g2_nand2_1 _19913_ (.Y(_12842_),
    .A(_12658_),
    .B(_12830_));
 sg13g2_o21ai_1 _19914_ (.B1(_12842_),
    .Y(_01071_),
    .A1(net361),
    .A2(_12841_));
 sg13g2_nand2_1 _19915_ (.Y(_12843_),
    .A(net692),
    .B(\mem.mem_internal.code_mem[207][6] ));
 sg13g2_nand2_1 _19916_ (.Y(_12844_),
    .A(_12662_),
    .B(_12830_));
 sg13g2_o21ai_1 _19917_ (.B1(_12844_),
    .Y(_01072_),
    .A1(net361),
    .A2(_12843_));
 sg13g2_buf_1 _19918_ (.A(_12678_),
    .X(_12845_));
 sg13g2_nand2_1 _19919_ (.Y(_12846_),
    .A(net691),
    .B(\mem.mem_internal.code_mem[207][7] ));
 sg13g2_nand2_1 _19920_ (.Y(_12847_),
    .A(_12666_),
    .B(_12830_));
 sg13g2_o21ai_1 _19921_ (.B1(_12847_),
    .Y(_01073_),
    .A1(_12831_),
    .A2(_12846_));
 sg13g2_nand2_1 _19922_ (.Y(_12848_),
    .A(net843),
    .B(\mem.mem_internal.code_mem[208][0] ));
 sg13g2_nand3_1 _19923_ (.B(net1296),
    .C(_11355_),
    .A(net1297),
    .Y(_12849_));
 sg13g2_buf_2 _19924_ (.A(_12849_),
    .X(_12850_));
 sg13g2_buf_1 _19925_ (.A(_12850_),
    .X(_12851_));
 sg13g2_nor2_1 _19926_ (.A(_10232_),
    .B(net461),
    .Y(_12852_));
 sg13g2_buf_2 _19927_ (.A(_12852_),
    .X(_12853_));
 sg13g2_buf_1 _19928_ (.A(_12853_),
    .X(_12854_));
 sg13g2_buf_1 _19929_ (.A(_12637_),
    .X(_12855_));
 sg13g2_nand2_1 _19930_ (.Y(_12856_),
    .A(net1094),
    .B(net212));
 sg13g2_o21ai_1 _19931_ (.B1(_12856_),
    .Y(_01074_),
    .A1(_12848_),
    .A2(net212));
 sg13g2_nand2_1 _19932_ (.Y(_12857_),
    .A(_12845_),
    .B(\mem.mem_internal.code_mem[208][1] ));
 sg13g2_buf_1 _19933_ (.A(_12641_),
    .X(_12858_));
 sg13g2_nand2_1 _19934_ (.Y(_12859_),
    .A(net1093),
    .B(net212));
 sg13g2_o21ai_1 _19935_ (.B1(_12859_),
    .Y(_01075_),
    .A1(net212),
    .A2(_12857_));
 sg13g2_nand2_1 _19936_ (.Y(_12860_),
    .A(net691),
    .B(\mem.mem_internal.code_mem[208][2] ));
 sg13g2_buf_1 _19937_ (.A(_12645_),
    .X(_12861_));
 sg13g2_nand2_1 _19938_ (.Y(_12862_),
    .A(net1092),
    .B(_12853_));
 sg13g2_o21ai_1 _19939_ (.B1(_12862_),
    .Y(_01076_),
    .A1(_12854_),
    .A2(_12860_));
 sg13g2_nand2_1 _19940_ (.Y(_12863_),
    .A(net691),
    .B(\mem.mem_internal.code_mem[208][3] ));
 sg13g2_buf_1 _19941_ (.A(_12649_),
    .X(_12864_));
 sg13g2_nand2_1 _19942_ (.Y(_12865_),
    .A(net1091),
    .B(_12853_));
 sg13g2_o21ai_1 _19943_ (.B1(_12865_),
    .Y(_01077_),
    .A1(net212),
    .A2(_12863_));
 sg13g2_nand2_1 _19944_ (.Y(_12866_),
    .A(net691),
    .B(\mem.mem_internal.code_mem[208][4] ));
 sg13g2_buf_1 _19945_ (.A(_12653_),
    .X(_12867_));
 sg13g2_nand2_1 _19946_ (.Y(_12868_),
    .A(net1090),
    .B(_12853_));
 sg13g2_o21ai_1 _19947_ (.B1(_12868_),
    .Y(_01078_),
    .A1(_12854_),
    .A2(_12866_));
 sg13g2_nand2_1 _19948_ (.Y(_12869_),
    .A(net691),
    .B(\mem.mem_internal.code_mem[208][5] ));
 sg13g2_buf_1 _19949_ (.A(_12657_),
    .X(_12870_));
 sg13g2_nand2_1 _19950_ (.Y(_12871_),
    .A(net1089),
    .B(_12853_));
 sg13g2_o21ai_1 _19951_ (.B1(_12871_),
    .Y(_01079_),
    .A1(net212),
    .A2(_12869_));
 sg13g2_nand2_1 _19952_ (.Y(_12872_),
    .A(net691),
    .B(\mem.mem_internal.code_mem[208][6] ));
 sg13g2_buf_1 _19953_ (.A(_12661_),
    .X(_12873_));
 sg13g2_nand2_1 _19954_ (.Y(_12874_),
    .A(net1088),
    .B(_12853_));
 sg13g2_o21ai_1 _19955_ (.B1(_12874_),
    .Y(_01080_),
    .A1(net212),
    .A2(_12872_));
 sg13g2_nand2_1 _19956_ (.Y(_12875_),
    .A(net691),
    .B(\mem.mem_internal.code_mem[208][7] ));
 sg13g2_buf_1 _19957_ (.A(_12665_),
    .X(_12876_));
 sg13g2_nand2_1 _19958_ (.Y(_12877_),
    .A(net1087),
    .B(_12853_));
 sg13g2_o21ai_1 _19959_ (.B1(_12877_),
    .Y(_01081_),
    .A1(net212),
    .A2(_12875_));
 sg13g2_buf_2 _19960_ (.A(net1273),
    .X(_12878_));
 sg13g2_buf_1 _19961_ (.A(_12878_),
    .X(_12879_));
 sg13g2_nand2_1 _19962_ (.Y(_12880_),
    .A(_12879_),
    .B(\mem.mem_internal.code_mem[209][0] ));
 sg13g2_nor2_1 _19963_ (.A(_10632_),
    .B(net461),
    .Y(_12881_));
 sg13g2_buf_2 _19964_ (.A(_12881_),
    .X(_12882_));
 sg13g2_buf_1 _19965_ (.A(_12882_),
    .X(_12883_));
 sg13g2_nand2_1 _19966_ (.Y(_12884_),
    .A(net1094),
    .B(net211));
 sg13g2_o21ai_1 _19967_ (.B1(_12884_),
    .Y(_01082_),
    .A1(_12880_),
    .A2(net211));
 sg13g2_nand2_1 _19968_ (.Y(_12885_),
    .A(_12845_),
    .B(\mem.mem_internal.code_mem[209][1] ));
 sg13g2_nand2_1 _19969_ (.Y(_12886_),
    .A(net1093),
    .B(net211));
 sg13g2_o21ai_1 _19970_ (.B1(_12886_),
    .Y(_01083_),
    .A1(net211),
    .A2(_12885_));
 sg13g2_nand2_1 _19971_ (.Y(_12887_),
    .A(net691),
    .B(\mem.mem_internal.code_mem[209][2] ));
 sg13g2_nand2_1 _19972_ (.Y(_12888_),
    .A(net1092),
    .B(_12882_));
 sg13g2_o21ai_1 _19973_ (.B1(_12888_),
    .Y(_01084_),
    .A1(net211),
    .A2(_12887_));
 sg13g2_buf_1 _19974_ (.A(_11875_),
    .X(_12889_));
 sg13g2_buf_1 _19975_ (.A(_12889_),
    .X(_12890_));
 sg13g2_nand2_1 _19976_ (.Y(_12891_),
    .A(net690),
    .B(\mem.mem_internal.code_mem[209][3] ));
 sg13g2_nand2_1 _19977_ (.Y(_12892_),
    .A(net1091),
    .B(_12882_));
 sg13g2_o21ai_1 _19978_ (.B1(_12892_),
    .Y(_01085_),
    .A1(_12883_),
    .A2(_12891_));
 sg13g2_nand2_1 _19979_ (.Y(_12893_),
    .A(net690),
    .B(\mem.mem_internal.code_mem[209][4] ));
 sg13g2_nand2_1 _19980_ (.Y(_12894_),
    .A(net1090),
    .B(_12882_));
 sg13g2_o21ai_1 _19981_ (.B1(_12894_),
    .Y(_01086_),
    .A1(net211),
    .A2(_12893_));
 sg13g2_nand2_1 _19982_ (.Y(_12895_),
    .A(net690),
    .B(\mem.mem_internal.code_mem[209][5] ));
 sg13g2_nand2_1 _19983_ (.Y(_12896_),
    .A(net1089),
    .B(_12882_));
 sg13g2_o21ai_1 _19984_ (.B1(_12896_),
    .Y(_01087_),
    .A1(net211),
    .A2(_12895_));
 sg13g2_nand2_1 _19985_ (.Y(_12897_),
    .A(_12890_),
    .B(\mem.mem_internal.code_mem[209][6] ));
 sg13g2_nand2_1 _19986_ (.Y(_12898_),
    .A(net1088),
    .B(_12882_));
 sg13g2_o21ai_1 _19987_ (.B1(_12898_),
    .Y(_01088_),
    .A1(_12883_),
    .A2(_12897_));
 sg13g2_nand2_1 _19988_ (.Y(_12899_),
    .A(_12890_),
    .B(\mem.mem_internal.code_mem[209][7] ));
 sg13g2_nand2_1 _19989_ (.Y(_12900_),
    .A(net1087),
    .B(_12882_));
 sg13g2_o21ai_1 _19990_ (.B1(_12900_),
    .Y(_01089_),
    .A1(net211),
    .A2(_12899_));
 sg13g2_nand2_1 _19991_ (.Y(_12901_),
    .A(net842),
    .B(\mem.mem_internal.code_mem[20][0] ));
 sg13g2_nor2_1 _19992_ (.A(_10295_),
    .B(net464),
    .Y(_12902_));
 sg13g2_buf_2 _19993_ (.A(_12902_),
    .X(_12903_));
 sg13g2_buf_1 _19994_ (.A(_12903_),
    .X(_12904_));
 sg13g2_nand2_1 _19995_ (.Y(_12905_),
    .A(net1094),
    .B(net210));
 sg13g2_o21ai_1 _19996_ (.B1(_12905_),
    .Y(_01090_),
    .A1(_12901_),
    .A2(net210));
 sg13g2_nand2_1 _19997_ (.Y(_12906_),
    .A(net690),
    .B(\mem.mem_internal.code_mem[20][1] ));
 sg13g2_nand2_1 _19998_ (.Y(_12907_),
    .A(net1093),
    .B(_12904_));
 sg13g2_o21ai_1 _19999_ (.B1(_12907_),
    .Y(_01091_),
    .A1(net210),
    .A2(_12906_));
 sg13g2_nand2_1 _20000_ (.Y(_12908_),
    .A(net690),
    .B(\mem.mem_internal.code_mem[20][2] ));
 sg13g2_nand2_1 _20001_ (.Y(_12909_),
    .A(_12861_),
    .B(_12903_));
 sg13g2_o21ai_1 _20002_ (.B1(_12909_),
    .Y(_01092_),
    .A1(net210),
    .A2(_12908_));
 sg13g2_nand2_1 _20003_ (.Y(_12910_),
    .A(net690),
    .B(\mem.mem_internal.code_mem[20][3] ));
 sg13g2_nand2_1 _20004_ (.Y(_12911_),
    .A(_12864_),
    .B(_12903_));
 sg13g2_o21ai_1 _20005_ (.B1(_12911_),
    .Y(_01093_),
    .A1(net210),
    .A2(_12910_));
 sg13g2_nand2_1 _20006_ (.Y(_12912_),
    .A(net690),
    .B(\mem.mem_internal.code_mem[20][4] ));
 sg13g2_nand2_1 _20007_ (.Y(_12913_),
    .A(_12867_),
    .B(_12903_));
 sg13g2_o21ai_1 _20008_ (.B1(_12913_),
    .Y(_01094_),
    .A1(_12904_),
    .A2(_12912_));
 sg13g2_nand2_1 _20009_ (.Y(_12914_),
    .A(net690),
    .B(\mem.mem_internal.code_mem[20][5] ));
 sg13g2_nand2_1 _20010_ (.Y(_12915_),
    .A(net1089),
    .B(_12903_));
 sg13g2_o21ai_1 _20011_ (.B1(_12915_),
    .Y(_01095_),
    .A1(net210),
    .A2(_12914_));
 sg13g2_buf_1 _20012_ (.A(_12889_),
    .X(_12916_));
 sg13g2_nand2_1 _20013_ (.Y(_12917_),
    .A(net689),
    .B(\mem.mem_internal.code_mem[20][6] ));
 sg13g2_nand2_1 _20014_ (.Y(_12918_),
    .A(net1088),
    .B(_12903_));
 sg13g2_o21ai_1 _20015_ (.B1(_12918_),
    .Y(_01096_),
    .A1(net210),
    .A2(_12917_));
 sg13g2_nand2_1 _20016_ (.Y(_12919_),
    .A(net689),
    .B(\mem.mem_internal.code_mem[20][7] ));
 sg13g2_nand2_1 _20017_ (.Y(_12920_),
    .A(_12876_),
    .B(_12903_));
 sg13g2_o21ai_1 _20018_ (.B1(_12920_),
    .Y(_01097_),
    .A1(net210),
    .A2(_12919_));
 sg13g2_nand2_1 _20019_ (.Y(_12921_),
    .A(net842),
    .B(\mem.mem_internal.code_mem[210][0] ));
 sg13g2_nor2_1 _20020_ (.A(_10656_),
    .B(_12851_),
    .Y(_12922_));
 sg13g2_buf_2 _20021_ (.A(_12922_),
    .X(_12923_));
 sg13g2_buf_1 _20022_ (.A(_12923_),
    .X(_12924_));
 sg13g2_nand2_1 _20023_ (.Y(_12925_),
    .A(_12855_),
    .B(net209));
 sg13g2_o21ai_1 _20024_ (.B1(_12925_),
    .Y(_01098_),
    .A1(_12921_),
    .A2(net209));
 sg13g2_nand2_1 _20025_ (.Y(_12926_),
    .A(net689),
    .B(\mem.mem_internal.code_mem[210][1] ));
 sg13g2_nand2_1 _20026_ (.Y(_12927_),
    .A(net1093),
    .B(net209));
 sg13g2_o21ai_1 _20027_ (.B1(_12927_),
    .Y(_01099_),
    .A1(net209),
    .A2(_12926_));
 sg13g2_nand2_1 _20028_ (.Y(_12928_),
    .A(net689),
    .B(\mem.mem_internal.code_mem[210][2] ));
 sg13g2_nand2_1 _20029_ (.Y(_12929_),
    .A(net1092),
    .B(_12923_));
 sg13g2_o21ai_1 _20030_ (.B1(_12929_),
    .Y(_01100_),
    .A1(net209),
    .A2(_12928_));
 sg13g2_nand2_1 _20031_ (.Y(_12930_),
    .A(net689),
    .B(\mem.mem_internal.code_mem[210][3] ));
 sg13g2_nand2_1 _20032_ (.Y(_12931_),
    .A(net1091),
    .B(_12923_));
 sg13g2_o21ai_1 _20033_ (.B1(_12931_),
    .Y(_01101_),
    .A1(_12924_),
    .A2(_12930_));
 sg13g2_nand2_1 _20034_ (.Y(_12932_),
    .A(net689),
    .B(\mem.mem_internal.code_mem[210][4] ));
 sg13g2_nand2_1 _20035_ (.Y(_12933_),
    .A(net1090),
    .B(_12923_));
 sg13g2_o21ai_1 _20036_ (.B1(_12933_),
    .Y(_01102_),
    .A1(net209),
    .A2(_12932_));
 sg13g2_nand2_1 _20037_ (.Y(_12934_),
    .A(net689),
    .B(\mem.mem_internal.code_mem[210][5] ));
 sg13g2_nand2_1 _20038_ (.Y(_12935_),
    .A(net1089),
    .B(_12923_));
 sg13g2_o21ai_1 _20039_ (.B1(_12935_),
    .Y(_01103_),
    .A1(net209),
    .A2(_12934_));
 sg13g2_nand2_1 _20040_ (.Y(_12936_),
    .A(net689),
    .B(\mem.mem_internal.code_mem[210][6] ));
 sg13g2_nand2_1 _20041_ (.Y(_12937_),
    .A(net1088),
    .B(_12923_));
 sg13g2_o21ai_1 _20042_ (.B1(_12937_),
    .Y(_01104_),
    .A1(net209),
    .A2(_12936_));
 sg13g2_nand2_1 _20043_ (.Y(_12938_),
    .A(_12916_),
    .B(\mem.mem_internal.code_mem[210][7] ));
 sg13g2_nand2_1 _20044_ (.Y(_12939_),
    .A(net1087),
    .B(_12923_));
 sg13g2_o21ai_1 _20045_ (.B1(_12939_),
    .Y(_01105_),
    .A1(_12924_),
    .A2(_12938_));
 sg13g2_nand2_1 _20046_ (.Y(_12940_),
    .A(_12879_),
    .B(\mem.mem_internal.code_mem[211][0] ));
 sg13g2_nor2_1 _20047_ (.A(_10679_),
    .B(net461),
    .Y(_12941_));
 sg13g2_buf_2 _20048_ (.A(_12941_),
    .X(_12942_));
 sg13g2_buf_1 _20049_ (.A(_12942_),
    .X(_12943_));
 sg13g2_nand2_1 _20050_ (.Y(_12944_),
    .A(_12855_),
    .B(net208));
 sg13g2_o21ai_1 _20051_ (.B1(_12944_),
    .Y(_01106_),
    .A1(_12940_),
    .A2(net208));
 sg13g2_nand2_1 _20052_ (.Y(_12945_),
    .A(_12916_),
    .B(\mem.mem_internal.code_mem[211][1] ));
 sg13g2_nand2_1 _20053_ (.Y(_12946_),
    .A(net1093),
    .B(_12943_));
 sg13g2_o21ai_1 _20054_ (.B1(_12946_),
    .Y(_01107_),
    .A1(_12943_),
    .A2(_12945_));
 sg13g2_buf_1 _20055_ (.A(_12889_),
    .X(_12947_));
 sg13g2_nand2_1 _20056_ (.Y(_12948_),
    .A(net688),
    .B(\mem.mem_internal.code_mem[211][2] ));
 sg13g2_nand2_1 _20057_ (.Y(_12949_),
    .A(net1092),
    .B(_12942_));
 sg13g2_o21ai_1 _20058_ (.B1(_12949_),
    .Y(_01108_),
    .A1(net208),
    .A2(_12948_));
 sg13g2_nand2_1 _20059_ (.Y(_12950_),
    .A(net688),
    .B(\mem.mem_internal.code_mem[211][3] ));
 sg13g2_nand2_1 _20060_ (.Y(_12951_),
    .A(net1091),
    .B(_12942_));
 sg13g2_o21ai_1 _20061_ (.B1(_12951_),
    .Y(_01109_),
    .A1(net208),
    .A2(_12950_));
 sg13g2_nand2_1 _20062_ (.Y(_12952_),
    .A(net688),
    .B(\mem.mem_internal.code_mem[211][4] ));
 sg13g2_nand2_1 _20063_ (.Y(_12953_),
    .A(net1090),
    .B(_12942_));
 sg13g2_o21ai_1 _20064_ (.B1(_12953_),
    .Y(_01110_),
    .A1(net208),
    .A2(_12952_));
 sg13g2_nand2_1 _20065_ (.Y(_12954_),
    .A(net688),
    .B(\mem.mem_internal.code_mem[211][5] ));
 sg13g2_nand2_1 _20066_ (.Y(_12955_),
    .A(net1089),
    .B(_12942_));
 sg13g2_o21ai_1 _20067_ (.B1(_12955_),
    .Y(_01111_),
    .A1(net208),
    .A2(_12954_));
 sg13g2_nand2_1 _20068_ (.Y(_12956_),
    .A(net688),
    .B(\mem.mem_internal.code_mem[211][6] ));
 sg13g2_nand2_1 _20069_ (.Y(_12957_),
    .A(net1088),
    .B(_12942_));
 sg13g2_o21ai_1 _20070_ (.B1(_12957_),
    .Y(_01112_),
    .A1(net208),
    .A2(_12956_));
 sg13g2_nand2_1 _20071_ (.Y(_12958_),
    .A(net688),
    .B(\mem.mem_internal.code_mem[211][7] ));
 sg13g2_nand2_1 _20072_ (.Y(_12959_),
    .A(net1087),
    .B(_12942_));
 sg13g2_o21ai_1 _20073_ (.B1(_12959_),
    .Y(_01113_),
    .A1(net208),
    .A2(_12958_));
 sg13g2_nand2_1 _20074_ (.Y(_12960_),
    .A(net842),
    .B(\mem.mem_internal.code_mem[212][0] ));
 sg13g2_nor2_1 _20075_ (.A(_10295_),
    .B(net461),
    .Y(_12961_));
 sg13g2_buf_2 _20076_ (.A(_12961_),
    .X(_12962_));
 sg13g2_buf_1 _20077_ (.A(_12962_),
    .X(_12963_));
 sg13g2_nand2_1 _20078_ (.Y(_12964_),
    .A(net1094),
    .B(net207));
 sg13g2_o21ai_1 _20079_ (.B1(_12964_),
    .Y(_01114_),
    .A1(_12960_),
    .A2(net207));
 sg13g2_nand2_1 _20080_ (.Y(_12965_),
    .A(net688),
    .B(\mem.mem_internal.code_mem[212][1] ));
 sg13g2_nand2_1 _20081_ (.Y(_12966_),
    .A(net1093),
    .B(net207));
 sg13g2_o21ai_1 _20082_ (.B1(_12966_),
    .Y(_01115_),
    .A1(net207),
    .A2(_12965_));
 sg13g2_nand2_1 _20083_ (.Y(_12967_),
    .A(net688),
    .B(\mem.mem_internal.code_mem[212][2] ));
 sg13g2_nand2_1 _20084_ (.Y(_12968_),
    .A(net1092),
    .B(_12962_));
 sg13g2_o21ai_1 _20085_ (.B1(_12968_),
    .Y(_01116_),
    .A1(net207),
    .A2(_12967_));
 sg13g2_nand2_1 _20086_ (.Y(_12969_),
    .A(_12947_),
    .B(\mem.mem_internal.code_mem[212][3] ));
 sg13g2_nand2_1 _20087_ (.Y(_12970_),
    .A(net1091),
    .B(_12962_));
 sg13g2_o21ai_1 _20088_ (.B1(_12970_),
    .Y(_01117_),
    .A1(net207),
    .A2(_12969_));
 sg13g2_nand2_1 _20089_ (.Y(_12971_),
    .A(_12947_),
    .B(\mem.mem_internal.code_mem[212][4] ));
 sg13g2_nand2_1 _20090_ (.Y(_12972_),
    .A(net1090),
    .B(_12962_));
 sg13g2_o21ai_1 _20091_ (.B1(_12972_),
    .Y(_01118_),
    .A1(net207),
    .A2(_12971_));
 sg13g2_buf_1 _20092_ (.A(_12889_),
    .X(_12973_));
 sg13g2_nand2_1 _20093_ (.Y(_12974_),
    .A(net687),
    .B(\mem.mem_internal.code_mem[212][5] ));
 sg13g2_nand2_1 _20094_ (.Y(_12975_),
    .A(net1089),
    .B(_12962_));
 sg13g2_o21ai_1 _20095_ (.B1(_12975_),
    .Y(_01119_),
    .A1(_12963_),
    .A2(_12974_));
 sg13g2_nand2_1 _20096_ (.Y(_12976_),
    .A(net687),
    .B(\mem.mem_internal.code_mem[212][6] ));
 sg13g2_nand2_1 _20097_ (.Y(_12977_),
    .A(net1088),
    .B(_12962_));
 sg13g2_o21ai_1 _20098_ (.B1(_12977_),
    .Y(_01120_),
    .A1(_12963_),
    .A2(_12976_));
 sg13g2_nand2_1 _20099_ (.Y(_12978_),
    .A(net687),
    .B(\mem.mem_internal.code_mem[212][7] ));
 sg13g2_nand2_1 _20100_ (.Y(_12979_),
    .A(net1087),
    .B(_12962_));
 sg13g2_o21ai_1 _20101_ (.B1(_12979_),
    .Y(_01121_),
    .A1(net207),
    .A2(_12978_));
 sg13g2_nand2_1 _20102_ (.Y(_12980_),
    .A(net842),
    .B(\mem.mem_internal.code_mem[213][0] ));
 sg13g2_nor2_1 _20103_ (.A(_10325_),
    .B(net461),
    .Y(_12981_));
 sg13g2_buf_2 _20104_ (.A(_12981_),
    .X(_12982_));
 sg13g2_buf_1 _20105_ (.A(_12982_),
    .X(_12983_));
 sg13g2_nand2_1 _20106_ (.Y(_12984_),
    .A(net1094),
    .B(net206));
 sg13g2_o21ai_1 _20107_ (.B1(_12984_),
    .Y(_01122_),
    .A1(_12980_),
    .A2(net206));
 sg13g2_nand2_1 _20108_ (.Y(_12985_),
    .A(net687),
    .B(\mem.mem_internal.code_mem[213][1] ));
 sg13g2_nand2_1 _20109_ (.Y(_12986_),
    .A(net1093),
    .B(net206));
 sg13g2_o21ai_1 _20110_ (.B1(_12986_),
    .Y(_01123_),
    .A1(net206),
    .A2(_12985_));
 sg13g2_nand2_1 _20111_ (.Y(_12987_),
    .A(net687),
    .B(\mem.mem_internal.code_mem[213][2] ));
 sg13g2_nand2_1 _20112_ (.Y(_12988_),
    .A(net1092),
    .B(_12982_));
 sg13g2_o21ai_1 _20113_ (.B1(_12988_),
    .Y(_01124_),
    .A1(net206),
    .A2(_12987_));
 sg13g2_nand2_1 _20114_ (.Y(_12989_),
    .A(net687),
    .B(\mem.mem_internal.code_mem[213][3] ));
 sg13g2_nand2_1 _20115_ (.Y(_12990_),
    .A(net1091),
    .B(_12982_));
 sg13g2_o21ai_1 _20116_ (.B1(_12990_),
    .Y(_01125_),
    .A1(net206),
    .A2(_12989_));
 sg13g2_nand2_1 _20117_ (.Y(_12991_),
    .A(net687),
    .B(\mem.mem_internal.code_mem[213][4] ));
 sg13g2_nand2_1 _20118_ (.Y(_12992_),
    .A(net1090),
    .B(_12982_));
 sg13g2_o21ai_1 _20119_ (.B1(_12992_),
    .Y(_01126_),
    .A1(net206),
    .A2(_12991_));
 sg13g2_nand2_1 _20120_ (.Y(_12993_),
    .A(_12973_),
    .B(\mem.mem_internal.code_mem[213][5] ));
 sg13g2_nand2_1 _20121_ (.Y(_12994_),
    .A(net1089),
    .B(_12982_));
 sg13g2_o21ai_1 _20122_ (.B1(_12994_),
    .Y(_01127_),
    .A1(net206),
    .A2(_12993_));
 sg13g2_nand2_1 _20123_ (.Y(_12995_),
    .A(_12973_),
    .B(\mem.mem_internal.code_mem[213][6] ));
 sg13g2_nand2_1 _20124_ (.Y(_12996_),
    .A(net1088),
    .B(_12982_));
 sg13g2_o21ai_1 _20125_ (.B1(_12996_),
    .Y(_01128_),
    .A1(_12983_),
    .A2(_12995_));
 sg13g2_nand2_1 _20126_ (.Y(_12997_),
    .A(net687),
    .B(\mem.mem_internal.code_mem[213][7] ));
 sg13g2_nand2_1 _20127_ (.Y(_12998_),
    .A(net1087),
    .B(_12982_));
 sg13g2_o21ai_1 _20128_ (.B1(_12998_),
    .Y(_01129_),
    .A1(_12983_),
    .A2(_12997_));
 sg13g2_nand2_1 _20129_ (.Y(_12999_),
    .A(net842),
    .B(\mem.mem_internal.code_mem[214][0] ));
 sg13g2_nor2_1 _20130_ (.A(net779),
    .B(_12851_),
    .Y(_13000_));
 sg13g2_buf_2 _20131_ (.A(_13000_),
    .X(_13001_));
 sg13g2_buf_1 _20132_ (.A(_13001_),
    .X(_13002_));
 sg13g2_nand2_1 _20133_ (.Y(_13003_),
    .A(net1094),
    .B(net205));
 sg13g2_o21ai_1 _20134_ (.B1(_13003_),
    .Y(_01130_),
    .A1(_12999_),
    .A2(net205));
 sg13g2_buf_1 _20135_ (.A(_12889_),
    .X(_13004_));
 sg13g2_nand2_1 _20136_ (.Y(_13005_),
    .A(net686),
    .B(\mem.mem_internal.code_mem[214][1] ));
 sg13g2_nand2_1 _20137_ (.Y(_13006_),
    .A(_12858_),
    .B(net205));
 sg13g2_o21ai_1 _20138_ (.B1(_13006_),
    .Y(_01131_),
    .A1(net205),
    .A2(_13005_));
 sg13g2_nand2_1 _20139_ (.Y(_13007_),
    .A(net686),
    .B(\mem.mem_internal.code_mem[214][2] ));
 sg13g2_nand2_1 _20140_ (.Y(_13008_),
    .A(net1092),
    .B(_13001_));
 sg13g2_o21ai_1 _20141_ (.B1(_13008_),
    .Y(_01132_),
    .A1(net205),
    .A2(_13007_));
 sg13g2_nand2_1 _20142_ (.Y(_13009_),
    .A(net686),
    .B(\mem.mem_internal.code_mem[214][3] ));
 sg13g2_nand2_1 _20143_ (.Y(_13010_),
    .A(net1091),
    .B(_13001_));
 sg13g2_o21ai_1 _20144_ (.B1(_13010_),
    .Y(_01133_),
    .A1(_13002_),
    .A2(_13009_));
 sg13g2_nand2_1 _20145_ (.Y(_13011_),
    .A(net686),
    .B(\mem.mem_internal.code_mem[214][4] ));
 sg13g2_nand2_1 _20146_ (.Y(_13012_),
    .A(net1090),
    .B(_13001_));
 sg13g2_o21ai_1 _20147_ (.B1(_13012_),
    .Y(_01134_),
    .A1(net205),
    .A2(_13011_));
 sg13g2_nand2_1 _20148_ (.Y(_13013_),
    .A(net686),
    .B(\mem.mem_internal.code_mem[214][5] ));
 sg13g2_nand2_1 _20149_ (.Y(_13014_),
    .A(_12870_),
    .B(_13001_));
 sg13g2_o21ai_1 _20150_ (.B1(_13014_),
    .Y(_01135_),
    .A1(net205),
    .A2(_13013_));
 sg13g2_nand2_1 _20151_ (.Y(_13015_),
    .A(_13004_),
    .B(\mem.mem_internal.code_mem[214][6] ));
 sg13g2_nand2_1 _20152_ (.Y(_13016_),
    .A(_12873_),
    .B(_13001_));
 sg13g2_o21ai_1 _20153_ (.B1(_13016_),
    .Y(_01136_),
    .A1(_13002_),
    .A2(_13015_));
 sg13g2_nand2_1 _20154_ (.Y(_13017_),
    .A(net686),
    .B(\mem.mem_internal.code_mem[214][7] ));
 sg13g2_nand2_1 _20155_ (.Y(_13018_),
    .A(_12876_),
    .B(_13001_));
 sg13g2_o21ai_1 _20156_ (.B1(_13018_),
    .Y(_01137_),
    .A1(net205),
    .A2(_13017_));
 sg13g2_nand2_1 _20157_ (.Y(_13019_),
    .A(net842),
    .B(\mem.mem_internal.code_mem[215][0] ));
 sg13g2_nor2_1 _20158_ (.A(_10372_),
    .B(net461),
    .Y(_13020_));
 sg13g2_buf_2 _20159_ (.A(_13020_),
    .X(_13021_));
 sg13g2_buf_1 _20160_ (.A(_13021_),
    .X(_13022_));
 sg13g2_nand2_1 _20161_ (.Y(_13023_),
    .A(net1094),
    .B(net204));
 sg13g2_o21ai_1 _20162_ (.B1(_13023_),
    .Y(_01138_),
    .A1(_13019_),
    .A2(net204));
 sg13g2_nand2_1 _20163_ (.Y(_13024_),
    .A(net686),
    .B(\mem.mem_internal.code_mem[215][1] ));
 sg13g2_nand2_1 _20164_ (.Y(_13025_),
    .A(_12858_),
    .B(net204));
 sg13g2_o21ai_1 _20165_ (.B1(_13025_),
    .Y(_01139_),
    .A1(net204),
    .A2(_13024_));
 sg13g2_nand2_1 _20166_ (.Y(_13026_),
    .A(net686),
    .B(\mem.mem_internal.code_mem[215][2] ));
 sg13g2_nand2_1 _20167_ (.Y(_13027_),
    .A(_12861_),
    .B(_13021_));
 sg13g2_o21ai_1 _20168_ (.B1(_13027_),
    .Y(_01140_),
    .A1(_13022_),
    .A2(_13026_));
 sg13g2_nand2_1 _20169_ (.Y(_13028_),
    .A(_13004_),
    .B(\mem.mem_internal.code_mem[215][3] ));
 sg13g2_nand2_1 _20170_ (.Y(_13029_),
    .A(_12864_),
    .B(_13021_));
 sg13g2_o21ai_1 _20171_ (.B1(_13029_),
    .Y(_01141_),
    .A1(net204),
    .A2(_13028_));
 sg13g2_buf_1 _20172_ (.A(_12889_),
    .X(_13030_));
 sg13g2_nand2_1 _20173_ (.Y(_13031_),
    .A(_13030_),
    .B(\mem.mem_internal.code_mem[215][4] ));
 sg13g2_nand2_1 _20174_ (.Y(_13032_),
    .A(_12867_),
    .B(_13021_));
 sg13g2_o21ai_1 _20175_ (.B1(_13032_),
    .Y(_01142_),
    .A1(net204),
    .A2(_13031_));
 sg13g2_nand2_1 _20176_ (.Y(_13033_),
    .A(_13030_),
    .B(\mem.mem_internal.code_mem[215][5] ));
 sg13g2_nand2_1 _20177_ (.Y(_13034_),
    .A(_12870_),
    .B(_13021_));
 sg13g2_o21ai_1 _20178_ (.B1(_13034_),
    .Y(_01143_),
    .A1(net204),
    .A2(_13033_));
 sg13g2_nand2_1 _20179_ (.Y(_13035_),
    .A(net685),
    .B(\mem.mem_internal.code_mem[215][6] ));
 sg13g2_nand2_1 _20180_ (.Y(_13036_),
    .A(_12873_),
    .B(_13021_));
 sg13g2_o21ai_1 _20181_ (.B1(_13036_),
    .Y(_01144_),
    .A1(_13022_),
    .A2(_13035_));
 sg13g2_nand2_1 _20182_ (.Y(_13037_),
    .A(net685),
    .B(\mem.mem_internal.code_mem[215][7] ));
 sg13g2_nand2_1 _20183_ (.Y(_13038_),
    .A(net1087),
    .B(_13021_));
 sg13g2_o21ai_1 _20184_ (.B1(_13038_),
    .Y(_01145_),
    .A1(net204),
    .A2(_13037_));
 sg13g2_nand2_1 _20185_ (.Y(_13039_),
    .A(net842),
    .B(\mem.mem_internal.code_mem[216][0] ));
 sg13g2_nor2_1 _20186_ (.A(net778),
    .B(net461),
    .Y(_13040_));
 sg13g2_buf_2 _20187_ (.A(_13040_),
    .X(_13041_));
 sg13g2_buf_1 _20188_ (.A(_13041_),
    .X(_13042_));
 sg13g2_nand2_1 _20189_ (.Y(_02779_),
    .A(net1094),
    .B(net203));
 sg13g2_o21ai_1 _20190_ (.B1(_02779_),
    .Y(_01146_),
    .A1(_13039_),
    .A2(net203));
 sg13g2_nand2_1 _20191_ (.Y(_02780_),
    .A(net685),
    .B(\mem.mem_internal.code_mem[216][1] ));
 sg13g2_nand2_1 _20192_ (.Y(_02781_),
    .A(net1093),
    .B(net203));
 sg13g2_o21ai_1 _20193_ (.B1(_02781_),
    .Y(_01147_),
    .A1(net203),
    .A2(_02780_));
 sg13g2_nand2_1 _20194_ (.Y(_02782_),
    .A(net685),
    .B(\mem.mem_internal.code_mem[216][2] ));
 sg13g2_nand2_1 _20195_ (.Y(_02783_),
    .A(net1092),
    .B(_13041_));
 sg13g2_o21ai_1 _20196_ (.B1(_02783_),
    .Y(_01148_),
    .A1(_13042_),
    .A2(_02782_));
 sg13g2_nand2_1 _20197_ (.Y(_02784_),
    .A(net685),
    .B(\mem.mem_internal.code_mem[216][3] ));
 sg13g2_nand2_1 _20198_ (.Y(_02785_),
    .A(net1091),
    .B(_13041_));
 sg13g2_o21ai_1 _20199_ (.B1(_02785_),
    .Y(_01149_),
    .A1(net203),
    .A2(_02784_));
 sg13g2_nand2_1 _20200_ (.Y(_02786_),
    .A(net685),
    .B(\mem.mem_internal.code_mem[216][4] ));
 sg13g2_nand2_1 _20201_ (.Y(_02787_),
    .A(net1090),
    .B(_13041_));
 sg13g2_o21ai_1 _20202_ (.B1(_02787_),
    .Y(_01150_),
    .A1(net203),
    .A2(_02786_));
 sg13g2_nand2_1 _20203_ (.Y(_02788_),
    .A(net685),
    .B(\mem.mem_internal.code_mem[216][5] ));
 sg13g2_nand2_1 _20204_ (.Y(_02789_),
    .A(net1089),
    .B(_13041_));
 sg13g2_o21ai_1 _20205_ (.B1(_02789_),
    .Y(_01151_),
    .A1(net203),
    .A2(_02788_));
 sg13g2_nand2_1 _20206_ (.Y(_02790_),
    .A(net685),
    .B(\mem.mem_internal.code_mem[216][6] ));
 sg13g2_nand2_1 _20207_ (.Y(_02791_),
    .A(net1088),
    .B(_13041_));
 sg13g2_o21ai_1 _20208_ (.B1(_02791_),
    .Y(_01152_),
    .A1(_13042_),
    .A2(_02790_));
 sg13g2_buf_1 _20209_ (.A(_12889_),
    .X(_02792_));
 sg13g2_nand2_1 _20210_ (.Y(_02793_),
    .A(net684),
    .B(\mem.mem_internal.code_mem[216][7] ));
 sg13g2_nand2_1 _20211_ (.Y(_02794_),
    .A(net1087),
    .B(_13041_));
 sg13g2_o21ai_1 _20212_ (.B1(_02794_),
    .Y(_01153_),
    .A1(net203),
    .A2(_02793_));
 sg13g2_nand2_1 _20213_ (.Y(_02795_),
    .A(net842),
    .B(\mem.mem_internal.code_mem[217][0] ));
 sg13g2_nor2_1 _20214_ (.A(_10422_),
    .B(net461),
    .Y(_02796_));
 sg13g2_buf_2 _20215_ (.A(_02796_),
    .X(_02797_));
 sg13g2_buf_1 _20216_ (.A(_02797_),
    .X(_02798_));
 sg13g2_buf_1 _20217_ (.A(_12637_),
    .X(_02799_));
 sg13g2_nand2_1 _20218_ (.Y(_02800_),
    .A(net1086),
    .B(net202));
 sg13g2_o21ai_1 _20219_ (.B1(_02800_),
    .Y(_01154_),
    .A1(_02795_),
    .A2(net202));
 sg13g2_nand2_1 _20220_ (.Y(_02801_),
    .A(_02792_),
    .B(\mem.mem_internal.code_mem[217][1] ));
 sg13g2_buf_1 _20221_ (.A(_12641_),
    .X(_02802_));
 sg13g2_nand2_1 _20222_ (.Y(_02803_),
    .A(net1085),
    .B(_02798_));
 sg13g2_o21ai_1 _20223_ (.B1(_02803_),
    .Y(_01155_),
    .A1(_02798_),
    .A2(_02801_));
 sg13g2_nand2_1 _20224_ (.Y(_02804_),
    .A(net684),
    .B(\mem.mem_internal.code_mem[217][2] ));
 sg13g2_buf_1 _20225_ (.A(_12645_),
    .X(_02805_));
 sg13g2_nand2_1 _20226_ (.Y(_02806_),
    .A(net1084),
    .B(_02797_));
 sg13g2_o21ai_1 _20227_ (.B1(_02806_),
    .Y(_01156_),
    .A1(net202),
    .A2(_02804_));
 sg13g2_nand2_1 _20228_ (.Y(_02807_),
    .A(net684),
    .B(\mem.mem_internal.code_mem[217][3] ));
 sg13g2_buf_1 _20229_ (.A(_12649_),
    .X(_02808_));
 sg13g2_nand2_1 _20230_ (.Y(_02809_),
    .A(net1083),
    .B(_02797_));
 sg13g2_o21ai_1 _20231_ (.B1(_02809_),
    .Y(_01157_),
    .A1(net202),
    .A2(_02807_));
 sg13g2_nand2_1 _20232_ (.Y(_02810_),
    .A(net684),
    .B(\mem.mem_internal.code_mem[217][4] ));
 sg13g2_buf_1 _20233_ (.A(_12653_),
    .X(_02811_));
 sg13g2_nand2_1 _20234_ (.Y(_02812_),
    .A(net1082),
    .B(_02797_));
 sg13g2_o21ai_1 _20235_ (.B1(_02812_),
    .Y(_01158_),
    .A1(net202),
    .A2(_02810_));
 sg13g2_nand2_1 _20236_ (.Y(_02813_),
    .A(net684),
    .B(\mem.mem_internal.code_mem[217][5] ));
 sg13g2_buf_1 _20237_ (.A(_12657_),
    .X(_02814_));
 sg13g2_nand2_1 _20238_ (.Y(_02815_),
    .A(net1081),
    .B(_02797_));
 sg13g2_o21ai_1 _20239_ (.B1(_02815_),
    .Y(_01159_),
    .A1(net202),
    .A2(_02813_));
 sg13g2_nand2_1 _20240_ (.Y(_02816_),
    .A(net684),
    .B(\mem.mem_internal.code_mem[217][6] ));
 sg13g2_buf_1 _20241_ (.A(_12661_),
    .X(_02817_));
 sg13g2_nand2_1 _20242_ (.Y(_02818_),
    .A(net1080),
    .B(_02797_));
 sg13g2_o21ai_1 _20243_ (.B1(_02818_),
    .Y(_01160_),
    .A1(net202),
    .A2(_02816_));
 sg13g2_nand2_1 _20244_ (.Y(_02819_),
    .A(net684),
    .B(\mem.mem_internal.code_mem[217][7] ));
 sg13g2_buf_1 _20245_ (.A(_12665_),
    .X(_02820_));
 sg13g2_nand2_1 _20246_ (.Y(_02821_),
    .A(net1079),
    .B(_02797_));
 sg13g2_o21ai_1 _20247_ (.B1(_02821_),
    .Y(_01161_),
    .A1(net202),
    .A2(_02819_));
 sg13g2_buf_1 _20248_ (.A(_12878_),
    .X(_02822_));
 sg13g2_nand2_1 _20249_ (.Y(_02823_),
    .A(net841),
    .B(\mem.mem_internal.code_mem[218][0] ));
 sg13g2_nor2_1 _20250_ (.A(_10444_),
    .B(_12850_),
    .Y(_02824_));
 sg13g2_buf_2 _20251_ (.A(_02824_),
    .X(_02825_));
 sg13g2_buf_1 _20252_ (.A(_02825_),
    .X(_02826_));
 sg13g2_nand2_1 _20253_ (.Y(_02827_),
    .A(net1086),
    .B(net360));
 sg13g2_o21ai_1 _20254_ (.B1(_02827_),
    .Y(_01162_),
    .A1(_02823_),
    .A2(net360));
 sg13g2_nand2_1 _20255_ (.Y(_02828_),
    .A(_02792_),
    .B(\mem.mem_internal.code_mem[218][1] ));
 sg13g2_nand2_1 _20256_ (.Y(_02829_),
    .A(net1085),
    .B(net360));
 sg13g2_o21ai_1 _20257_ (.B1(_02829_),
    .Y(_01163_),
    .A1(net360),
    .A2(_02828_));
 sg13g2_nand2_1 _20258_ (.Y(_02830_),
    .A(net684),
    .B(\mem.mem_internal.code_mem[218][2] ));
 sg13g2_nand2_1 _20259_ (.Y(_02831_),
    .A(net1084),
    .B(_02825_));
 sg13g2_o21ai_1 _20260_ (.B1(_02831_),
    .Y(_01164_),
    .A1(_02826_),
    .A2(_02830_));
 sg13g2_buf_1 _20261_ (.A(_11875_),
    .X(_02832_));
 sg13g2_buf_1 _20262_ (.A(_02832_),
    .X(_02833_));
 sg13g2_nand2_1 _20263_ (.Y(_02834_),
    .A(_02833_),
    .B(\mem.mem_internal.code_mem[218][3] ));
 sg13g2_nand2_1 _20264_ (.Y(_02835_),
    .A(net1083),
    .B(_02825_));
 sg13g2_o21ai_1 _20265_ (.B1(_02835_),
    .Y(_01165_),
    .A1(net360),
    .A2(_02834_));
 sg13g2_nand2_1 _20266_ (.Y(_02836_),
    .A(net683),
    .B(\mem.mem_internal.code_mem[218][4] ));
 sg13g2_nand2_1 _20267_ (.Y(_02837_),
    .A(net1082),
    .B(_02825_));
 sg13g2_o21ai_1 _20268_ (.B1(_02837_),
    .Y(_01166_),
    .A1(_02826_),
    .A2(_02836_));
 sg13g2_nand2_1 _20269_ (.Y(_02838_),
    .A(net683),
    .B(\mem.mem_internal.code_mem[218][5] ));
 sg13g2_nand2_1 _20270_ (.Y(_02839_),
    .A(net1081),
    .B(_02825_));
 sg13g2_o21ai_1 _20271_ (.B1(_02839_),
    .Y(_01167_),
    .A1(net360),
    .A2(_02838_));
 sg13g2_nand2_1 _20272_ (.Y(_02840_),
    .A(net683),
    .B(\mem.mem_internal.code_mem[218][6] ));
 sg13g2_nand2_1 _20273_ (.Y(_02841_),
    .A(net1080),
    .B(_02825_));
 sg13g2_o21ai_1 _20274_ (.B1(_02841_),
    .Y(_01168_),
    .A1(net360),
    .A2(_02840_));
 sg13g2_nand2_1 _20275_ (.Y(_02842_),
    .A(net683),
    .B(\mem.mem_internal.code_mem[218][7] ));
 sg13g2_nand2_1 _20276_ (.Y(_02843_),
    .A(net1079),
    .B(_02825_));
 sg13g2_o21ai_1 _20277_ (.B1(_02843_),
    .Y(_01169_),
    .A1(net360),
    .A2(_02842_));
 sg13g2_nand2_1 _20278_ (.Y(_02844_),
    .A(net841),
    .B(\mem.mem_internal.code_mem[219][0] ));
 sg13g2_nor2_1 _20279_ (.A(net775),
    .B(_12850_),
    .Y(_02845_));
 sg13g2_buf_2 _20280_ (.A(_02845_),
    .X(_02846_));
 sg13g2_buf_1 _20281_ (.A(_02846_),
    .X(_02847_));
 sg13g2_nand2_1 _20282_ (.Y(_02848_),
    .A(net1086),
    .B(net359));
 sg13g2_o21ai_1 _20283_ (.B1(_02848_),
    .Y(_01170_),
    .A1(_02844_),
    .A2(net359));
 sg13g2_nand2_1 _20284_ (.Y(_02849_),
    .A(net683),
    .B(\mem.mem_internal.code_mem[219][1] ));
 sg13g2_nand2_1 _20285_ (.Y(_02850_),
    .A(net1085),
    .B(net359));
 sg13g2_o21ai_1 _20286_ (.B1(_02850_),
    .Y(_01171_),
    .A1(net359),
    .A2(_02849_));
 sg13g2_nand2_1 _20287_ (.Y(_02851_),
    .A(net683),
    .B(\mem.mem_internal.code_mem[219][2] ));
 sg13g2_nand2_1 _20288_ (.Y(_02852_),
    .A(net1084),
    .B(_02846_));
 sg13g2_o21ai_1 _20289_ (.B1(_02852_),
    .Y(_01172_),
    .A1(net359),
    .A2(_02851_));
 sg13g2_nand2_1 _20290_ (.Y(_02853_),
    .A(net683),
    .B(\mem.mem_internal.code_mem[219][3] ));
 sg13g2_nand2_1 _20291_ (.Y(_02854_),
    .A(net1083),
    .B(_02846_));
 sg13g2_o21ai_1 _20292_ (.B1(_02854_),
    .Y(_01173_),
    .A1(_02847_),
    .A2(_02853_));
 sg13g2_nand2_1 _20293_ (.Y(_02855_),
    .A(net683),
    .B(\mem.mem_internal.code_mem[219][4] ));
 sg13g2_nand2_1 _20294_ (.Y(_02856_),
    .A(net1082),
    .B(_02846_));
 sg13g2_o21ai_1 _20295_ (.B1(_02856_),
    .Y(_01174_),
    .A1(net359),
    .A2(_02855_));
 sg13g2_nand2_1 _20296_ (.Y(_02857_),
    .A(_02833_),
    .B(\mem.mem_internal.code_mem[219][5] ));
 sg13g2_nand2_1 _20297_ (.Y(_02858_),
    .A(net1081),
    .B(_02846_));
 sg13g2_o21ai_1 _20298_ (.B1(_02858_),
    .Y(_01175_),
    .A1(_02847_),
    .A2(_02857_));
 sg13g2_buf_1 _20299_ (.A(_02832_),
    .X(_02859_));
 sg13g2_nand2_1 _20300_ (.Y(_02860_),
    .A(net682),
    .B(\mem.mem_internal.code_mem[219][6] ));
 sg13g2_nand2_1 _20301_ (.Y(_02861_),
    .A(net1080),
    .B(_02846_));
 sg13g2_o21ai_1 _20302_ (.B1(_02861_),
    .Y(_01176_),
    .A1(net359),
    .A2(_02860_));
 sg13g2_nand2_1 _20303_ (.Y(_02862_),
    .A(_02859_),
    .B(\mem.mem_internal.code_mem[219][7] ));
 sg13g2_nand2_1 _20304_ (.Y(_02863_),
    .A(net1079),
    .B(_02846_));
 sg13g2_o21ai_1 _20305_ (.B1(_02863_),
    .Y(_01177_),
    .A1(net359),
    .A2(_02862_));
 sg13g2_nand2_1 _20306_ (.Y(_02864_),
    .A(net841),
    .B(\mem.mem_internal.code_mem[21][0] ));
 sg13g2_nor2_1 _20307_ (.A(_10325_),
    .B(net464),
    .Y(_02865_));
 sg13g2_buf_2 _20308_ (.A(_02865_),
    .X(_02866_));
 sg13g2_buf_1 _20309_ (.A(_02866_),
    .X(_02867_));
 sg13g2_nand2_1 _20310_ (.Y(_02868_),
    .A(net1086),
    .B(net201));
 sg13g2_o21ai_1 _20311_ (.B1(_02868_),
    .Y(_01178_),
    .A1(_02864_),
    .A2(net201));
 sg13g2_nand2_1 _20312_ (.Y(_02869_),
    .A(net682),
    .B(\mem.mem_internal.code_mem[21][1] ));
 sg13g2_nand2_1 _20313_ (.Y(_02870_),
    .A(net1085),
    .B(_02867_));
 sg13g2_o21ai_1 _20314_ (.B1(_02870_),
    .Y(_01179_),
    .A1(net201),
    .A2(_02869_));
 sg13g2_nand2_1 _20315_ (.Y(_02871_),
    .A(net682),
    .B(\mem.mem_internal.code_mem[21][2] ));
 sg13g2_nand2_1 _20316_ (.Y(_02872_),
    .A(net1084),
    .B(_02866_));
 sg13g2_o21ai_1 _20317_ (.B1(_02872_),
    .Y(_01180_),
    .A1(net201),
    .A2(_02871_));
 sg13g2_nand2_1 _20318_ (.Y(_02873_),
    .A(net682),
    .B(\mem.mem_internal.code_mem[21][3] ));
 sg13g2_nand2_1 _20319_ (.Y(_02874_),
    .A(net1083),
    .B(_02866_));
 sg13g2_o21ai_1 _20320_ (.B1(_02874_),
    .Y(_01181_),
    .A1(net201),
    .A2(_02873_));
 sg13g2_nand2_1 _20321_ (.Y(_02875_),
    .A(net682),
    .B(\mem.mem_internal.code_mem[21][4] ));
 sg13g2_nand2_1 _20322_ (.Y(_02876_),
    .A(net1082),
    .B(_02866_));
 sg13g2_o21ai_1 _20323_ (.B1(_02876_),
    .Y(_01182_),
    .A1(net201),
    .A2(_02875_));
 sg13g2_nand2_1 _20324_ (.Y(_02877_),
    .A(net682),
    .B(\mem.mem_internal.code_mem[21][5] ));
 sg13g2_nand2_1 _20325_ (.Y(_02878_),
    .A(net1081),
    .B(_02866_));
 sg13g2_o21ai_1 _20326_ (.B1(_02878_),
    .Y(_01183_),
    .A1(net201),
    .A2(_02877_));
 sg13g2_nand2_1 _20327_ (.Y(_02879_),
    .A(net682),
    .B(\mem.mem_internal.code_mem[21][6] ));
 sg13g2_nand2_1 _20328_ (.Y(_02880_),
    .A(net1080),
    .B(_02866_));
 sg13g2_o21ai_1 _20329_ (.B1(_02880_),
    .Y(_01184_),
    .A1(net201),
    .A2(_02879_));
 sg13g2_nand2_1 _20330_ (.Y(_02881_),
    .A(net682),
    .B(\mem.mem_internal.code_mem[21][7] ));
 sg13g2_nand2_1 _20331_ (.Y(_02882_),
    .A(net1079),
    .B(_02866_));
 sg13g2_o21ai_1 _20332_ (.B1(_02882_),
    .Y(_01185_),
    .A1(_02867_),
    .A2(_02881_));
 sg13g2_nand2_1 _20333_ (.Y(_02883_),
    .A(net841),
    .B(\mem.mem_internal.code_mem[220][0] ));
 sg13g2_nor2_1 _20334_ (.A(_10491_),
    .B(_12850_),
    .Y(_02884_));
 sg13g2_buf_2 _20335_ (.A(_02884_),
    .X(_02885_));
 sg13g2_buf_1 _20336_ (.A(_02885_),
    .X(_02886_));
 sg13g2_nand2_1 _20337_ (.Y(_02887_),
    .A(net1086),
    .B(net358));
 sg13g2_o21ai_1 _20338_ (.B1(_02887_),
    .Y(_01186_),
    .A1(_02883_),
    .A2(net358));
 sg13g2_nand2_1 _20339_ (.Y(_02888_),
    .A(_02859_),
    .B(\mem.mem_internal.code_mem[220][1] ));
 sg13g2_nand2_1 _20340_ (.Y(_02889_),
    .A(net1085),
    .B(net358));
 sg13g2_o21ai_1 _20341_ (.B1(_02889_),
    .Y(_01187_),
    .A1(net358),
    .A2(_02888_));
 sg13g2_buf_1 _20342_ (.A(_02832_),
    .X(_02890_));
 sg13g2_nand2_1 _20343_ (.Y(_02891_),
    .A(net681),
    .B(\mem.mem_internal.code_mem[220][2] ));
 sg13g2_nand2_1 _20344_ (.Y(_02892_),
    .A(net1084),
    .B(_02885_));
 sg13g2_o21ai_1 _20345_ (.B1(_02892_),
    .Y(_01188_),
    .A1(net358),
    .A2(_02891_));
 sg13g2_nand2_1 _20346_ (.Y(_02893_),
    .A(net681),
    .B(\mem.mem_internal.code_mem[220][3] ));
 sg13g2_nand2_1 _20347_ (.Y(_02894_),
    .A(net1083),
    .B(_02885_));
 sg13g2_o21ai_1 _20348_ (.B1(_02894_),
    .Y(_01189_),
    .A1(_02886_),
    .A2(_02893_));
 sg13g2_nand2_1 _20349_ (.Y(_02895_),
    .A(net681),
    .B(\mem.mem_internal.code_mem[220][4] ));
 sg13g2_nand2_1 _20350_ (.Y(_02896_),
    .A(net1082),
    .B(_02885_));
 sg13g2_o21ai_1 _20351_ (.B1(_02896_),
    .Y(_01190_),
    .A1(_02886_),
    .A2(_02895_));
 sg13g2_nand2_1 _20352_ (.Y(_02897_),
    .A(net681),
    .B(\mem.mem_internal.code_mem[220][5] ));
 sg13g2_nand2_1 _20353_ (.Y(_02898_),
    .A(net1081),
    .B(_02885_));
 sg13g2_o21ai_1 _20354_ (.B1(_02898_),
    .Y(_01191_),
    .A1(net358),
    .A2(_02897_));
 sg13g2_nand2_1 _20355_ (.Y(_02899_),
    .A(net681),
    .B(\mem.mem_internal.code_mem[220][6] ));
 sg13g2_nand2_1 _20356_ (.Y(_02900_),
    .A(net1080),
    .B(_02885_));
 sg13g2_o21ai_1 _20357_ (.B1(_02900_),
    .Y(_01192_),
    .A1(net358),
    .A2(_02899_));
 sg13g2_nand2_1 _20358_ (.Y(_02901_),
    .A(net681),
    .B(\mem.mem_internal.code_mem[220][7] ));
 sg13g2_nand2_1 _20359_ (.Y(_02902_),
    .A(net1079),
    .B(_02885_));
 sg13g2_o21ai_1 _20360_ (.B1(_02902_),
    .Y(_01193_),
    .A1(net358),
    .A2(_02901_));
 sg13g2_nand2_1 _20361_ (.Y(_02903_),
    .A(net841),
    .B(\mem.mem_internal.code_mem[221][0] ));
 sg13g2_nor2_1 _20362_ (.A(_10513_),
    .B(_12850_),
    .Y(_02904_));
 sg13g2_buf_2 _20363_ (.A(_02904_),
    .X(_02905_));
 sg13g2_buf_1 _20364_ (.A(_02905_),
    .X(_02906_));
 sg13g2_nand2_1 _20365_ (.Y(_02907_),
    .A(net1086),
    .B(net357));
 sg13g2_o21ai_1 _20366_ (.B1(_02907_),
    .Y(_01194_),
    .A1(_02903_),
    .A2(net357));
 sg13g2_nand2_1 _20367_ (.Y(_02908_),
    .A(_02890_),
    .B(\mem.mem_internal.code_mem[221][1] ));
 sg13g2_nand2_1 _20368_ (.Y(_02909_),
    .A(net1085),
    .B(_02906_));
 sg13g2_o21ai_1 _20369_ (.B1(_02909_),
    .Y(_01195_),
    .A1(net357),
    .A2(_02908_));
 sg13g2_nand2_1 _20370_ (.Y(_02910_),
    .A(_02890_),
    .B(\mem.mem_internal.code_mem[221][2] ));
 sg13g2_nand2_1 _20371_ (.Y(_02911_),
    .A(net1084),
    .B(_02905_));
 sg13g2_o21ai_1 _20372_ (.B1(_02911_),
    .Y(_01196_),
    .A1(net357),
    .A2(_02910_));
 sg13g2_nand2_1 _20373_ (.Y(_02912_),
    .A(net681),
    .B(\mem.mem_internal.code_mem[221][3] ));
 sg13g2_nand2_1 _20374_ (.Y(_02913_),
    .A(net1083),
    .B(_02905_));
 sg13g2_o21ai_1 _20375_ (.B1(_02913_),
    .Y(_01197_),
    .A1(net357),
    .A2(_02912_));
 sg13g2_nand2_1 _20376_ (.Y(_02914_),
    .A(net681),
    .B(\mem.mem_internal.code_mem[221][4] ));
 sg13g2_nand2_1 _20377_ (.Y(_02915_),
    .A(net1082),
    .B(_02905_));
 sg13g2_o21ai_1 _20378_ (.B1(_02915_),
    .Y(_01198_),
    .A1(net357),
    .A2(_02914_));
 sg13g2_buf_1 _20379_ (.A(_02832_),
    .X(_02916_));
 sg13g2_nand2_1 _20380_ (.Y(_02917_),
    .A(net680),
    .B(\mem.mem_internal.code_mem[221][5] ));
 sg13g2_nand2_1 _20381_ (.Y(_02918_),
    .A(net1081),
    .B(_02905_));
 sg13g2_o21ai_1 _20382_ (.B1(_02918_),
    .Y(_01199_),
    .A1(_02906_),
    .A2(_02917_));
 sg13g2_nand2_1 _20383_ (.Y(_02919_),
    .A(net680),
    .B(\mem.mem_internal.code_mem[221][6] ));
 sg13g2_nand2_1 _20384_ (.Y(_02920_),
    .A(net1080),
    .B(_02905_));
 sg13g2_o21ai_1 _20385_ (.B1(_02920_),
    .Y(_01200_),
    .A1(net357),
    .A2(_02919_));
 sg13g2_nand2_1 _20386_ (.Y(_02921_),
    .A(net680),
    .B(\mem.mem_internal.code_mem[221][7] ));
 sg13g2_nand2_1 _20387_ (.Y(_02922_),
    .A(net1079),
    .B(_02905_));
 sg13g2_o21ai_1 _20388_ (.B1(_02922_),
    .Y(_01201_),
    .A1(net357),
    .A2(_02921_));
 sg13g2_nand2_1 _20389_ (.Y(_02923_),
    .A(net841),
    .B(\mem.mem_internal.code_mem[222][0] ));
 sg13g2_nor2_1 _20390_ (.A(_10564_),
    .B(_12850_),
    .Y(_02924_));
 sg13g2_buf_2 _20391_ (.A(_02924_),
    .X(_02925_));
 sg13g2_buf_1 _20392_ (.A(_02925_),
    .X(_02926_));
 sg13g2_nand2_1 _20393_ (.Y(_02927_),
    .A(net1086),
    .B(net356));
 sg13g2_o21ai_1 _20394_ (.B1(_02927_),
    .Y(_01202_),
    .A1(_02923_),
    .A2(net356));
 sg13g2_nand2_1 _20395_ (.Y(_02928_),
    .A(_02916_),
    .B(\mem.mem_internal.code_mem[222][1] ));
 sg13g2_nand2_1 _20396_ (.Y(_02929_),
    .A(_02802_),
    .B(net356));
 sg13g2_o21ai_1 _20397_ (.B1(_02929_),
    .Y(_01203_),
    .A1(net356),
    .A2(_02928_));
 sg13g2_nand2_1 _20398_ (.Y(_02930_),
    .A(_02916_),
    .B(\mem.mem_internal.code_mem[222][2] ));
 sg13g2_nand2_1 _20399_ (.Y(_02931_),
    .A(_02805_),
    .B(_02925_));
 sg13g2_o21ai_1 _20400_ (.B1(_02931_),
    .Y(_01204_),
    .A1(net356),
    .A2(_02930_));
 sg13g2_nand2_1 _20401_ (.Y(_02932_),
    .A(net680),
    .B(\mem.mem_internal.code_mem[222][3] ));
 sg13g2_nand2_1 _20402_ (.Y(_02933_),
    .A(net1083),
    .B(_02925_));
 sg13g2_o21ai_1 _20403_ (.B1(_02933_),
    .Y(_01205_),
    .A1(net356),
    .A2(_02932_));
 sg13g2_nand2_1 _20404_ (.Y(_02934_),
    .A(net680),
    .B(\mem.mem_internal.code_mem[222][4] ));
 sg13g2_nand2_1 _20405_ (.Y(_02935_),
    .A(_02811_),
    .B(_02925_));
 sg13g2_o21ai_1 _20406_ (.B1(_02935_),
    .Y(_01206_),
    .A1(net356),
    .A2(_02934_));
 sg13g2_nand2_1 _20407_ (.Y(_02936_),
    .A(net680),
    .B(\mem.mem_internal.code_mem[222][5] ));
 sg13g2_nand2_1 _20408_ (.Y(_02937_),
    .A(_02814_),
    .B(_02925_));
 sg13g2_o21ai_1 _20409_ (.B1(_02937_),
    .Y(_01207_),
    .A1(_02926_),
    .A2(_02936_));
 sg13g2_nand2_1 _20410_ (.Y(_02938_),
    .A(net680),
    .B(\mem.mem_internal.code_mem[222][6] ));
 sg13g2_nand2_1 _20411_ (.Y(_02939_),
    .A(net1080),
    .B(_02925_));
 sg13g2_o21ai_1 _20412_ (.B1(_02939_),
    .Y(_01208_),
    .A1(_02926_),
    .A2(_02938_));
 sg13g2_nand2_1 _20413_ (.Y(_02940_),
    .A(net680),
    .B(\mem.mem_internal.code_mem[222][7] ));
 sg13g2_nand2_1 _20414_ (.Y(_02941_),
    .A(net1079),
    .B(_02925_));
 sg13g2_o21ai_1 _20415_ (.B1(_02941_),
    .Y(_01209_),
    .A1(net356),
    .A2(_02940_));
 sg13g2_nand2_1 _20416_ (.Y(_02942_),
    .A(net841),
    .B(\mem.mem_internal.code_mem[223][0] ));
 sg13g2_nor2_1 _20417_ (.A(_10586_),
    .B(_12850_),
    .Y(_02943_));
 sg13g2_buf_2 _20418_ (.A(_02943_),
    .X(_02944_));
 sg13g2_buf_1 _20419_ (.A(_02944_),
    .X(_02945_));
 sg13g2_nand2_1 _20420_ (.Y(_02946_),
    .A(_02799_),
    .B(net355));
 sg13g2_o21ai_1 _20421_ (.B1(_02946_),
    .Y(_01210_),
    .A1(_02942_),
    .A2(net355));
 sg13g2_buf_1 _20422_ (.A(_02832_),
    .X(_02947_));
 sg13g2_nand2_1 _20423_ (.Y(_02948_),
    .A(net679),
    .B(\mem.mem_internal.code_mem[223][1] ));
 sg13g2_nand2_1 _20424_ (.Y(_02949_),
    .A(_02802_),
    .B(net355));
 sg13g2_o21ai_1 _20425_ (.B1(_02949_),
    .Y(_01211_),
    .A1(net355),
    .A2(_02948_));
 sg13g2_nand2_1 _20426_ (.Y(_02950_),
    .A(net679),
    .B(\mem.mem_internal.code_mem[223][2] ));
 sg13g2_nand2_1 _20427_ (.Y(_02951_),
    .A(_02805_),
    .B(_02944_));
 sg13g2_o21ai_1 _20428_ (.B1(_02951_),
    .Y(_01212_),
    .A1(net355),
    .A2(_02950_));
 sg13g2_nand2_1 _20429_ (.Y(_02952_),
    .A(net679),
    .B(\mem.mem_internal.code_mem[223][3] ));
 sg13g2_nand2_1 _20430_ (.Y(_02953_),
    .A(net1083),
    .B(_02944_));
 sg13g2_o21ai_1 _20431_ (.B1(_02953_),
    .Y(_01213_),
    .A1(_02945_),
    .A2(_02952_));
 sg13g2_nand2_1 _20432_ (.Y(_02954_),
    .A(net679),
    .B(\mem.mem_internal.code_mem[223][4] ));
 sg13g2_nand2_1 _20433_ (.Y(_02955_),
    .A(_02811_),
    .B(_02944_));
 sg13g2_o21ai_1 _20434_ (.B1(_02955_),
    .Y(_01214_),
    .A1(_02945_),
    .A2(_02954_));
 sg13g2_nand2_1 _20435_ (.Y(_02956_),
    .A(net679),
    .B(\mem.mem_internal.code_mem[223][5] ));
 sg13g2_nand2_1 _20436_ (.Y(_02957_),
    .A(_02814_),
    .B(_02944_));
 sg13g2_o21ai_1 _20437_ (.B1(_02957_),
    .Y(_01215_),
    .A1(net355),
    .A2(_02956_));
 sg13g2_nand2_1 _20438_ (.Y(_02958_),
    .A(_02947_),
    .B(\mem.mem_internal.code_mem[223][6] ));
 sg13g2_nand2_1 _20439_ (.Y(_02959_),
    .A(net1080),
    .B(_02944_));
 sg13g2_o21ai_1 _20440_ (.B1(_02959_),
    .Y(_01216_),
    .A1(net355),
    .A2(_02958_));
 sg13g2_nand2_1 _20441_ (.Y(_02960_),
    .A(_02947_),
    .B(\mem.mem_internal.code_mem[223][7] ));
 sg13g2_nand2_1 _20442_ (.Y(_02961_),
    .A(net1079),
    .B(_02944_));
 sg13g2_o21ai_1 _20443_ (.B1(_02961_),
    .Y(_01217_),
    .A1(net355),
    .A2(_02960_));
 sg13g2_nand2_1 _20444_ (.Y(_02962_),
    .A(net841),
    .B(\mem.mem_internal.code_mem[224][0] ));
 sg13g2_nand3_1 _20445_ (.B(net1296),
    .C(_10298_),
    .A(net1297),
    .Y(_02963_));
 sg13g2_buf_2 _20446_ (.A(_02963_),
    .X(_02964_));
 sg13g2_buf_1 _20447_ (.A(_02964_),
    .X(_02965_));
 sg13g2_nor2_1 _20448_ (.A(_10232_),
    .B(net460),
    .Y(_02966_));
 sg13g2_buf_2 _20449_ (.A(_02966_),
    .X(_02967_));
 sg13g2_buf_1 _20450_ (.A(_02967_),
    .X(_02968_));
 sg13g2_nand2_1 _20451_ (.Y(_02969_),
    .A(net1086),
    .B(net200));
 sg13g2_o21ai_1 _20452_ (.B1(_02969_),
    .Y(_01218_),
    .A1(_02962_),
    .A2(net200));
 sg13g2_nand2_1 _20453_ (.Y(_02970_),
    .A(net679),
    .B(\mem.mem_internal.code_mem[224][1] ));
 sg13g2_nand2_1 _20454_ (.Y(_02971_),
    .A(net1085),
    .B(net200));
 sg13g2_o21ai_1 _20455_ (.B1(_02971_),
    .Y(_01219_),
    .A1(net200),
    .A2(_02970_));
 sg13g2_nand2_1 _20456_ (.Y(_02972_),
    .A(net679),
    .B(\mem.mem_internal.code_mem[224][2] ));
 sg13g2_nand2_1 _20457_ (.Y(_02973_),
    .A(net1084),
    .B(_02967_));
 sg13g2_o21ai_1 _20458_ (.B1(_02973_),
    .Y(_01220_),
    .A1(net200),
    .A2(_02972_));
 sg13g2_nand2_1 _20459_ (.Y(_02974_),
    .A(net679),
    .B(\mem.mem_internal.code_mem[224][3] ));
 sg13g2_nand2_1 _20460_ (.Y(_02975_),
    .A(_02808_),
    .B(_02967_));
 sg13g2_o21ai_1 _20461_ (.B1(_02975_),
    .Y(_01221_),
    .A1(net200),
    .A2(_02974_));
 sg13g2_buf_1 _20462_ (.A(_02832_),
    .X(_02976_));
 sg13g2_nand2_1 _20463_ (.Y(_02977_),
    .A(net678),
    .B(\mem.mem_internal.code_mem[224][4] ));
 sg13g2_nand2_1 _20464_ (.Y(_02978_),
    .A(net1082),
    .B(_02967_));
 sg13g2_o21ai_1 _20465_ (.B1(_02978_),
    .Y(_01222_),
    .A1(net200),
    .A2(_02977_));
 sg13g2_nand2_1 _20466_ (.Y(_02979_),
    .A(net678),
    .B(\mem.mem_internal.code_mem[224][5] ));
 sg13g2_nand2_1 _20467_ (.Y(_02980_),
    .A(net1081),
    .B(_02967_));
 sg13g2_o21ai_1 _20468_ (.B1(_02980_),
    .Y(_01223_),
    .A1(_02968_),
    .A2(_02979_));
 sg13g2_nand2_1 _20469_ (.Y(_02981_),
    .A(net678),
    .B(\mem.mem_internal.code_mem[224][6] ));
 sg13g2_nand2_1 _20470_ (.Y(_02982_),
    .A(_02817_),
    .B(_02967_));
 sg13g2_o21ai_1 _20471_ (.B1(_02982_),
    .Y(_01224_),
    .A1(_02968_),
    .A2(_02981_));
 sg13g2_nand2_1 _20472_ (.Y(_02983_),
    .A(net678),
    .B(\mem.mem_internal.code_mem[224][7] ));
 sg13g2_nand2_1 _20473_ (.Y(_02984_),
    .A(_02820_),
    .B(_02967_));
 sg13g2_o21ai_1 _20474_ (.B1(_02984_),
    .Y(_01225_),
    .A1(net200),
    .A2(_02983_));
 sg13g2_nand2_1 _20475_ (.Y(_02985_),
    .A(_02822_),
    .B(\mem.mem_internal.code_mem[225][0] ));
 sg13g2_nor2_1 _20476_ (.A(_10632_),
    .B(net460),
    .Y(_02986_));
 sg13g2_buf_2 _20477_ (.A(_02986_),
    .X(_02987_));
 sg13g2_buf_1 _20478_ (.A(_02987_),
    .X(_02988_));
 sg13g2_nand2_1 _20479_ (.Y(_02989_),
    .A(_02799_),
    .B(net199));
 sg13g2_o21ai_1 _20480_ (.B1(_02989_),
    .Y(_01226_),
    .A1(_02985_),
    .A2(net199));
 sg13g2_nand2_1 _20481_ (.Y(_02990_),
    .A(net678),
    .B(\mem.mem_internal.code_mem[225][1] ));
 sg13g2_nand2_1 _20482_ (.Y(_02991_),
    .A(net1085),
    .B(net199));
 sg13g2_o21ai_1 _20483_ (.B1(_02991_),
    .Y(_01227_),
    .A1(net199),
    .A2(_02990_));
 sg13g2_nand2_1 _20484_ (.Y(_02992_),
    .A(net678),
    .B(\mem.mem_internal.code_mem[225][2] ));
 sg13g2_nand2_1 _20485_ (.Y(_02993_),
    .A(net1084),
    .B(_02987_));
 sg13g2_o21ai_1 _20486_ (.B1(_02993_),
    .Y(_01228_),
    .A1(net199),
    .A2(_02992_));
 sg13g2_nand2_1 _20487_ (.Y(_02994_),
    .A(net678),
    .B(\mem.mem_internal.code_mem[225][3] ));
 sg13g2_nand2_1 _20488_ (.Y(_02995_),
    .A(_02808_),
    .B(_02987_));
 sg13g2_o21ai_1 _20489_ (.B1(_02995_),
    .Y(_01229_),
    .A1(net199),
    .A2(_02994_));
 sg13g2_nand2_1 _20490_ (.Y(_02996_),
    .A(net678),
    .B(\mem.mem_internal.code_mem[225][4] ));
 sg13g2_nand2_1 _20491_ (.Y(_02997_),
    .A(net1082),
    .B(_02987_));
 sg13g2_o21ai_1 _20492_ (.B1(_02997_),
    .Y(_01230_),
    .A1(net199),
    .A2(_02996_));
 sg13g2_nand2_1 _20493_ (.Y(_02998_),
    .A(_02976_),
    .B(\mem.mem_internal.code_mem[225][5] ));
 sg13g2_nand2_1 _20494_ (.Y(_02999_),
    .A(net1081),
    .B(_02987_));
 sg13g2_o21ai_1 _20495_ (.B1(_02999_),
    .Y(_01231_),
    .A1(_02988_),
    .A2(_02998_));
 sg13g2_nand2_1 _20496_ (.Y(_03000_),
    .A(_02976_),
    .B(\mem.mem_internal.code_mem[225][6] ));
 sg13g2_nand2_1 _20497_ (.Y(_03001_),
    .A(_02817_),
    .B(_02987_));
 sg13g2_o21ai_1 _20498_ (.B1(_03001_),
    .Y(_01232_),
    .A1(_02988_),
    .A2(_03000_));
 sg13g2_buf_1 _20499_ (.A(_02832_),
    .X(_03002_));
 sg13g2_nand2_1 _20500_ (.Y(_03003_),
    .A(_03002_),
    .B(\mem.mem_internal.code_mem[225][7] ));
 sg13g2_nand2_1 _20501_ (.Y(_03004_),
    .A(_02820_),
    .B(_02987_));
 sg13g2_o21ai_1 _20502_ (.B1(_03004_),
    .Y(_01233_),
    .A1(net199),
    .A2(_03003_));
 sg13g2_nand2_1 _20503_ (.Y(_03005_),
    .A(_02822_),
    .B(\mem.mem_internal.code_mem[226][0] ));
 sg13g2_nor2_1 _20504_ (.A(_10656_),
    .B(_02965_),
    .Y(_03006_));
 sg13g2_buf_2 _20505_ (.A(_03006_),
    .X(_03007_));
 sg13g2_buf_1 _20506_ (.A(_03007_),
    .X(_03008_));
 sg13g2_buf_1 _20507_ (.A(_12637_),
    .X(_03009_));
 sg13g2_nand2_1 _20508_ (.Y(_03010_),
    .A(net1078),
    .B(net198));
 sg13g2_o21ai_1 _20509_ (.B1(_03010_),
    .Y(_01234_),
    .A1(_03005_),
    .A2(net198));
 sg13g2_nand2_1 _20510_ (.Y(_03011_),
    .A(net677),
    .B(\mem.mem_internal.code_mem[226][1] ));
 sg13g2_buf_1 _20511_ (.A(_12641_),
    .X(_03012_));
 sg13g2_nand2_1 _20512_ (.Y(_03013_),
    .A(net1077),
    .B(net198));
 sg13g2_o21ai_1 _20513_ (.B1(_03013_),
    .Y(_01235_),
    .A1(net198),
    .A2(_03011_));
 sg13g2_nand2_1 _20514_ (.Y(_03014_),
    .A(_03002_),
    .B(\mem.mem_internal.code_mem[226][2] ));
 sg13g2_buf_1 _20515_ (.A(_12645_),
    .X(_03015_));
 sg13g2_nand2_1 _20516_ (.Y(_03016_),
    .A(net1076),
    .B(_03007_));
 sg13g2_o21ai_1 _20517_ (.B1(_03016_),
    .Y(_01236_),
    .A1(net198),
    .A2(_03014_));
 sg13g2_nand2_1 _20518_ (.Y(_03017_),
    .A(net677),
    .B(\mem.mem_internal.code_mem[226][3] ));
 sg13g2_buf_1 _20519_ (.A(_12649_),
    .X(_03018_));
 sg13g2_nand2_1 _20520_ (.Y(_03019_),
    .A(net1075),
    .B(_03007_));
 sg13g2_o21ai_1 _20521_ (.B1(_03019_),
    .Y(_01237_),
    .A1(net198),
    .A2(_03017_));
 sg13g2_nand2_1 _20522_ (.Y(_03020_),
    .A(net677),
    .B(\mem.mem_internal.code_mem[226][4] ));
 sg13g2_buf_1 _20523_ (.A(_12653_),
    .X(_03021_));
 sg13g2_nand2_1 _20524_ (.Y(_03022_),
    .A(net1074),
    .B(_03007_));
 sg13g2_o21ai_1 _20525_ (.B1(_03022_),
    .Y(_01238_),
    .A1(net198),
    .A2(_03020_));
 sg13g2_nand2_1 _20526_ (.Y(_03023_),
    .A(net677),
    .B(\mem.mem_internal.code_mem[226][5] ));
 sg13g2_buf_1 _20527_ (.A(_12657_),
    .X(_03024_));
 sg13g2_nand2_1 _20528_ (.Y(_03025_),
    .A(net1073),
    .B(_03007_));
 sg13g2_o21ai_1 _20529_ (.B1(_03025_),
    .Y(_01239_),
    .A1(_03008_),
    .A2(_03023_));
 sg13g2_nand2_1 _20530_ (.Y(_03026_),
    .A(net677),
    .B(\mem.mem_internal.code_mem[226][6] ));
 sg13g2_buf_1 _20531_ (.A(_12661_),
    .X(_03027_));
 sg13g2_nand2_1 _20532_ (.Y(_03028_),
    .A(net1072),
    .B(_03007_));
 sg13g2_o21ai_1 _20533_ (.B1(_03028_),
    .Y(_01240_),
    .A1(_03008_),
    .A2(_03026_));
 sg13g2_nand2_1 _20534_ (.Y(_03029_),
    .A(net677),
    .B(\mem.mem_internal.code_mem[226][7] ));
 sg13g2_buf_1 _20535_ (.A(_12665_),
    .X(_03030_));
 sg13g2_nand2_1 _20536_ (.Y(_03031_),
    .A(net1071),
    .B(_03007_));
 sg13g2_o21ai_1 _20537_ (.B1(_03031_),
    .Y(_01241_),
    .A1(net198),
    .A2(_03029_));
 sg13g2_buf_1 _20538_ (.A(_12878_),
    .X(_03032_));
 sg13g2_nand2_1 _20539_ (.Y(_03033_),
    .A(_03032_),
    .B(\mem.mem_internal.code_mem[227][0] ));
 sg13g2_nor2_1 _20540_ (.A(_10679_),
    .B(_02965_),
    .Y(_03034_));
 sg13g2_buf_2 _20541_ (.A(_03034_),
    .X(_03035_));
 sg13g2_buf_1 _20542_ (.A(_03035_),
    .X(_03036_));
 sg13g2_nand2_1 _20543_ (.Y(_03037_),
    .A(net1078),
    .B(net197));
 sg13g2_o21ai_1 _20544_ (.B1(_03037_),
    .Y(_01242_),
    .A1(_03033_),
    .A2(net197));
 sg13g2_nand2_1 _20545_ (.Y(_03038_),
    .A(net677),
    .B(\mem.mem_internal.code_mem[227][1] ));
 sg13g2_nand2_1 _20546_ (.Y(_03039_),
    .A(net1077),
    .B(net197));
 sg13g2_o21ai_1 _20547_ (.B1(_03039_),
    .Y(_01243_),
    .A1(net197),
    .A2(_03038_));
 sg13g2_nand2_1 _20548_ (.Y(_03040_),
    .A(net677),
    .B(\mem.mem_internal.code_mem[227][2] ));
 sg13g2_nand2_1 _20549_ (.Y(_03041_),
    .A(net1076),
    .B(_03035_));
 sg13g2_o21ai_1 _20550_ (.B1(_03041_),
    .Y(_01244_),
    .A1(net197),
    .A2(_03040_));
 sg13g2_buf_2 _20551_ (.A(net1276),
    .X(_03042_));
 sg13g2_buf_1 _20552_ (.A(_03042_),
    .X(_03043_));
 sg13g2_buf_1 _20553_ (.A(_03043_),
    .X(_03044_));
 sg13g2_nand2_1 _20554_ (.Y(_03045_),
    .A(net676),
    .B(\mem.mem_internal.code_mem[227][3] ));
 sg13g2_nand2_1 _20555_ (.Y(_03046_),
    .A(net1075),
    .B(_03035_));
 sg13g2_o21ai_1 _20556_ (.B1(_03046_),
    .Y(_01245_),
    .A1(net197),
    .A2(_03045_));
 sg13g2_nand2_1 _20557_ (.Y(_03047_),
    .A(net676),
    .B(\mem.mem_internal.code_mem[227][4] ));
 sg13g2_nand2_1 _20558_ (.Y(_03048_),
    .A(net1074),
    .B(_03035_));
 sg13g2_o21ai_1 _20559_ (.B1(_03048_),
    .Y(_01246_),
    .A1(net197),
    .A2(_03047_));
 sg13g2_nand2_1 _20560_ (.Y(_03049_),
    .A(net676),
    .B(\mem.mem_internal.code_mem[227][5] ));
 sg13g2_nand2_1 _20561_ (.Y(_03050_),
    .A(net1073),
    .B(_03035_));
 sg13g2_o21ai_1 _20562_ (.B1(_03050_),
    .Y(_01247_),
    .A1(_03036_),
    .A2(_03049_));
 sg13g2_nand2_1 _20563_ (.Y(_03051_),
    .A(_03044_),
    .B(\mem.mem_internal.code_mem[227][6] ));
 sg13g2_nand2_1 _20564_ (.Y(_03052_),
    .A(net1072),
    .B(_03035_));
 sg13g2_o21ai_1 _20565_ (.B1(_03052_),
    .Y(_01248_),
    .A1(_03036_),
    .A2(_03051_));
 sg13g2_nand2_1 _20566_ (.Y(_03053_),
    .A(net676),
    .B(\mem.mem_internal.code_mem[227][7] ));
 sg13g2_nand2_1 _20567_ (.Y(_03054_),
    .A(net1071),
    .B(_03035_));
 sg13g2_o21ai_1 _20568_ (.B1(_03054_),
    .Y(_01249_),
    .A1(net197),
    .A2(_03053_));
 sg13g2_nand2_1 _20569_ (.Y(_03055_),
    .A(net840),
    .B(\mem.mem_internal.code_mem[228][0] ));
 sg13g2_nor2_1 _20570_ (.A(_10295_),
    .B(net460),
    .Y(_03056_));
 sg13g2_buf_2 _20571_ (.A(_03056_),
    .X(_03057_));
 sg13g2_buf_1 _20572_ (.A(_03057_),
    .X(_03058_));
 sg13g2_nand2_1 _20573_ (.Y(_03059_),
    .A(net1078),
    .B(net196));
 sg13g2_o21ai_1 _20574_ (.B1(_03059_),
    .Y(_01250_),
    .A1(_03055_),
    .A2(net196));
 sg13g2_nand2_1 _20575_ (.Y(_03060_),
    .A(net676),
    .B(\mem.mem_internal.code_mem[228][1] ));
 sg13g2_nand2_1 _20576_ (.Y(_03061_),
    .A(net1077),
    .B(net196));
 sg13g2_o21ai_1 _20577_ (.B1(_03061_),
    .Y(_01251_),
    .A1(net196),
    .A2(_03060_));
 sg13g2_nand2_1 _20578_ (.Y(_03062_),
    .A(net676),
    .B(\mem.mem_internal.code_mem[228][2] ));
 sg13g2_nand2_1 _20579_ (.Y(_03063_),
    .A(net1076),
    .B(_03057_));
 sg13g2_o21ai_1 _20580_ (.B1(_03063_),
    .Y(_01252_),
    .A1(net196),
    .A2(_03062_));
 sg13g2_nand2_1 _20581_ (.Y(_03064_),
    .A(net676),
    .B(\mem.mem_internal.code_mem[228][3] ));
 sg13g2_nand2_1 _20582_ (.Y(_03065_),
    .A(net1075),
    .B(_03057_));
 sg13g2_o21ai_1 _20583_ (.B1(_03065_),
    .Y(_01253_),
    .A1(net196),
    .A2(_03064_));
 sg13g2_nand2_1 _20584_ (.Y(_03066_),
    .A(_03044_),
    .B(\mem.mem_internal.code_mem[228][4] ));
 sg13g2_nand2_1 _20585_ (.Y(_03067_),
    .A(net1074),
    .B(_03057_));
 sg13g2_o21ai_1 _20586_ (.B1(_03067_),
    .Y(_01254_),
    .A1(net196),
    .A2(_03066_));
 sg13g2_nand2_1 _20587_ (.Y(_03068_),
    .A(net676),
    .B(\mem.mem_internal.code_mem[228][5] ));
 sg13g2_nand2_1 _20588_ (.Y(_03069_),
    .A(net1073),
    .B(_03057_));
 sg13g2_o21ai_1 _20589_ (.B1(_03069_),
    .Y(_01255_),
    .A1(_03058_),
    .A2(_03068_));
 sg13g2_buf_1 _20590_ (.A(_03043_),
    .X(_03070_));
 sg13g2_nand2_1 _20591_ (.Y(_03071_),
    .A(net675),
    .B(\mem.mem_internal.code_mem[228][6] ));
 sg13g2_nand2_1 _20592_ (.Y(_03072_),
    .A(net1072),
    .B(_03057_));
 sg13g2_o21ai_1 _20593_ (.B1(_03072_),
    .Y(_01256_),
    .A1(_03058_),
    .A2(_03071_));
 sg13g2_nand2_1 _20594_ (.Y(_03073_),
    .A(net675),
    .B(\mem.mem_internal.code_mem[228][7] ));
 sg13g2_nand2_1 _20595_ (.Y(_03074_),
    .A(net1071),
    .B(_03057_));
 sg13g2_o21ai_1 _20596_ (.B1(_03074_),
    .Y(_01257_),
    .A1(net196),
    .A2(_03073_));
 sg13g2_nand2_1 _20597_ (.Y(_03075_),
    .A(net840),
    .B(\mem.mem_internal.code_mem[229][0] ));
 sg13g2_nor2_1 _20598_ (.A(_10325_),
    .B(net460),
    .Y(_03076_));
 sg13g2_buf_2 _20599_ (.A(_03076_),
    .X(_03077_));
 sg13g2_buf_1 _20600_ (.A(_03077_),
    .X(_03078_));
 sg13g2_nand2_1 _20601_ (.Y(_03079_),
    .A(_03009_),
    .B(net195));
 sg13g2_o21ai_1 _20602_ (.B1(_03079_),
    .Y(_01258_),
    .A1(_03075_),
    .A2(net195));
 sg13g2_nand2_1 _20603_ (.Y(_03080_),
    .A(net675),
    .B(\mem.mem_internal.code_mem[229][1] ));
 sg13g2_nand2_1 _20604_ (.Y(_03081_),
    .A(net1077),
    .B(net195));
 sg13g2_o21ai_1 _20605_ (.B1(_03081_),
    .Y(_01259_),
    .A1(net195),
    .A2(_03080_));
 sg13g2_nand2_1 _20606_ (.Y(_03082_),
    .A(net675),
    .B(\mem.mem_internal.code_mem[229][2] ));
 sg13g2_nand2_1 _20607_ (.Y(_03083_),
    .A(net1076),
    .B(_03077_));
 sg13g2_o21ai_1 _20608_ (.B1(_03083_),
    .Y(_01260_),
    .A1(net195),
    .A2(_03082_));
 sg13g2_nand2_1 _20609_ (.Y(_03084_),
    .A(_03070_),
    .B(\mem.mem_internal.code_mem[229][3] ));
 sg13g2_nand2_1 _20610_ (.Y(_03085_),
    .A(net1075),
    .B(_03077_));
 sg13g2_o21ai_1 _20611_ (.B1(_03085_),
    .Y(_01261_),
    .A1(net195),
    .A2(_03084_));
 sg13g2_nand2_1 _20612_ (.Y(_03086_),
    .A(_03070_),
    .B(\mem.mem_internal.code_mem[229][4] ));
 sg13g2_nand2_1 _20613_ (.Y(_03087_),
    .A(net1074),
    .B(_03077_));
 sg13g2_o21ai_1 _20614_ (.B1(_03087_),
    .Y(_01262_),
    .A1(net195),
    .A2(_03086_));
 sg13g2_nand2_1 _20615_ (.Y(_03088_),
    .A(net675),
    .B(\mem.mem_internal.code_mem[229][5] ));
 sg13g2_nand2_1 _20616_ (.Y(_03089_),
    .A(net1073),
    .B(_03077_));
 sg13g2_o21ai_1 _20617_ (.B1(_03089_),
    .Y(_01263_),
    .A1(_03078_),
    .A2(_03088_));
 sg13g2_nand2_1 _20618_ (.Y(_03090_),
    .A(net675),
    .B(\mem.mem_internal.code_mem[229][6] ));
 sg13g2_nand2_1 _20619_ (.Y(_03091_),
    .A(net1072),
    .B(_03077_));
 sg13g2_o21ai_1 _20620_ (.B1(_03091_),
    .Y(_01264_),
    .A1(_03078_),
    .A2(_03090_));
 sg13g2_nand2_1 _20621_ (.Y(_03092_),
    .A(net675),
    .B(\mem.mem_internal.code_mem[229][7] ));
 sg13g2_nand2_1 _20622_ (.Y(_03093_),
    .A(net1071),
    .B(_03077_));
 sg13g2_o21ai_1 _20623_ (.B1(_03093_),
    .Y(_01265_),
    .A1(net195),
    .A2(_03092_));
 sg13g2_nand2_1 _20624_ (.Y(_03094_),
    .A(net840),
    .B(\mem.mem_internal.code_mem[22][0] ));
 sg13g2_nor2_1 _20625_ (.A(net779),
    .B(net464),
    .Y(_03095_));
 sg13g2_buf_2 _20626_ (.A(_03095_),
    .X(_03096_));
 sg13g2_buf_1 _20627_ (.A(_03096_),
    .X(_03097_));
 sg13g2_nand2_1 _20628_ (.Y(_03098_),
    .A(net1078),
    .B(net194));
 sg13g2_o21ai_1 _20629_ (.B1(_03098_),
    .Y(_01266_),
    .A1(_03094_),
    .A2(net194));
 sg13g2_nand2_1 _20630_ (.Y(_03099_),
    .A(net675),
    .B(\mem.mem_internal.code_mem[22][1] ));
 sg13g2_nand2_1 _20631_ (.Y(_03100_),
    .A(net1077),
    .B(net194));
 sg13g2_o21ai_1 _20632_ (.B1(_03100_),
    .Y(_01267_),
    .A1(_03097_),
    .A2(_03099_));
 sg13g2_buf_1 _20633_ (.A(_03043_),
    .X(_03101_));
 sg13g2_nand2_1 _20634_ (.Y(_03102_),
    .A(net674),
    .B(\mem.mem_internal.code_mem[22][2] ));
 sg13g2_nand2_1 _20635_ (.Y(_03103_),
    .A(net1076),
    .B(_03096_));
 sg13g2_o21ai_1 _20636_ (.B1(_03103_),
    .Y(_01268_),
    .A1(net194),
    .A2(_03102_));
 sg13g2_nand2_1 _20637_ (.Y(_03104_),
    .A(net674),
    .B(\mem.mem_internal.code_mem[22][3] ));
 sg13g2_nand2_1 _20638_ (.Y(_03105_),
    .A(net1075),
    .B(_03096_));
 sg13g2_o21ai_1 _20639_ (.B1(_03105_),
    .Y(_01269_),
    .A1(_03097_),
    .A2(_03104_));
 sg13g2_nand2_1 _20640_ (.Y(_03106_),
    .A(net674),
    .B(\mem.mem_internal.code_mem[22][4] ));
 sg13g2_nand2_1 _20641_ (.Y(_03107_),
    .A(net1074),
    .B(_03096_));
 sg13g2_o21ai_1 _20642_ (.B1(_03107_),
    .Y(_01270_),
    .A1(net194),
    .A2(_03106_));
 sg13g2_nand2_1 _20643_ (.Y(_03108_),
    .A(net674),
    .B(\mem.mem_internal.code_mem[22][5] ));
 sg13g2_nand2_1 _20644_ (.Y(_03109_),
    .A(net1073),
    .B(_03096_));
 sg13g2_o21ai_1 _20645_ (.B1(_03109_),
    .Y(_01271_),
    .A1(net194),
    .A2(_03108_));
 sg13g2_nand2_1 _20646_ (.Y(_03110_),
    .A(net674),
    .B(\mem.mem_internal.code_mem[22][6] ));
 sg13g2_nand2_1 _20647_ (.Y(_03111_),
    .A(net1072),
    .B(_03096_));
 sg13g2_o21ai_1 _20648_ (.B1(_03111_),
    .Y(_01272_),
    .A1(net194),
    .A2(_03110_));
 sg13g2_nand2_1 _20649_ (.Y(_03112_),
    .A(net674),
    .B(\mem.mem_internal.code_mem[22][7] ));
 sg13g2_nand2_1 _20650_ (.Y(_03113_),
    .A(net1071),
    .B(_03096_));
 sg13g2_o21ai_1 _20651_ (.B1(_03113_),
    .Y(_01273_),
    .A1(net194),
    .A2(_03112_));
 sg13g2_nand2_1 _20652_ (.Y(_03114_),
    .A(net840),
    .B(\mem.mem_internal.code_mem[230][0] ));
 sg13g2_nor2_1 _20653_ (.A(_10349_),
    .B(net460),
    .Y(_03115_));
 sg13g2_buf_2 _20654_ (.A(_03115_),
    .X(_03116_));
 sg13g2_buf_1 _20655_ (.A(_03116_),
    .X(_03117_));
 sg13g2_nand2_1 _20656_ (.Y(_03118_),
    .A(_03009_),
    .B(net193));
 sg13g2_o21ai_1 _20657_ (.B1(_03118_),
    .Y(_01274_),
    .A1(_03114_),
    .A2(net193));
 sg13g2_nand2_1 _20658_ (.Y(_03119_),
    .A(net674),
    .B(\mem.mem_internal.code_mem[230][1] ));
 sg13g2_nand2_1 _20659_ (.Y(_03120_),
    .A(_03012_),
    .B(net193));
 sg13g2_o21ai_1 _20660_ (.B1(_03120_),
    .Y(_01275_),
    .A1(net193),
    .A2(_03119_));
 sg13g2_nand2_1 _20661_ (.Y(_03121_),
    .A(net674),
    .B(\mem.mem_internal.code_mem[230][2] ));
 sg13g2_nand2_1 _20662_ (.Y(_03122_),
    .A(_03015_),
    .B(_03116_));
 sg13g2_o21ai_1 _20663_ (.B1(_03122_),
    .Y(_01276_),
    .A1(net193),
    .A2(_03121_));
 sg13g2_nand2_1 _20664_ (.Y(_03123_),
    .A(_03101_),
    .B(\mem.mem_internal.code_mem[230][3] ));
 sg13g2_nand2_1 _20665_ (.Y(_03124_),
    .A(_03018_),
    .B(_03116_));
 sg13g2_o21ai_1 _20666_ (.B1(_03124_),
    .Y(_01277_),
    .A1(net193),
    .A2(_03123_));
 sg13g2_nand2_1 _20667_ (.Y(_03125_),
    .A(_03101_),
    .B(\mem.mem_internal.code_mem[230][4] ));
 sg13g2_nand2_1 _20668_ (.Y(_03126_),
    .A(_03021_),
    .B(_03116_));
 sg13g2_o21ai_1 _20669_ (.B1(_03126_),
    .Y(_01278_),
    .A1(_03117_),
    .A2(_03125_));
 sg13g2_buf_1 _20670_ (.A(_03043_),
    .X(_03127_));
 sg13g2_nand2_1 _20671_ (.Y(_03128_),
    .A(net673),
    .B(\mem.mem_internal.code_mem[230][5] ));
 sg13g2_nand2_1 _20672_ (.Y(_03129_),
    .A(_03024_),
    .B(_03116_));
 sg13g2_o21ai_1 _20673_ (.B1(_03129_),
    .Y(_01279_),
    .A1(_03117_),
    .A2(_03128_));
 sg13g2_nand2_1 _20674_ (.Y(_03130_),
    .A(net673),
    .B(\mem.mem_internal.code_mem[230][6] ));
 sg13g2_nand2_1 _20675_ (.Y(_03131_),
    .A(_03027_),
    .B(_03116_));
 sg13g2_o21ai_1 _20676_ (.B1(_03131_),
    .Y(_01280_),
    .A1(net193),
    .A2(_03130_));
 sg13g2_nand2_1 _20677_ (.Y(_03132_),
    .A(net673),
    .B(\mem.mem_internal.code_mem[230][7] ));
 sg13g2_nand2_1 _20678_ (.Y(_03133_),
    .A(_03030_),
    .B(_03116_));
 sg13g2_o21ai_1 _20679_ (.B1(_03133_),
    .Y(_01281_),
    .A1(net193),
    .A2(_03132_));
 sg13g2_nand2_1 _20680_ (.Y(_03134_),
    .A(_03032_),
    .B(\mem.mem_internal.code_mem[231][0] ));
 sg13g2_nor2_1 _20681_ (.A(_10372_),
    .B(net460),
    .Y(_03135_));
 sg13g2_buf_2 _20682_ (.A(_03135_),
    .X(_03136_));
 sg13g2_buf_1 _20683_ (.A(_03136_),
    .X(_03137_));
 sg13g2_nand2_1 _20684_ (.Y(_03138_),
    .A(net1078),
    .B(net192));
 sg13g2_o21ai_1 _20685_ (.B1(_03138_),
    .Y(_01282_),
    .A1(_03134_),
    .A2(net192));
 sg13g2_nand2_1 _20686_ (.Y(_03139_),
    .A(net673),
    .B(\mem.mem_internal.code_mem[231][1] ));
 sg13g2_nand2_1 _20687_ (.Y(_03140_),
    .A(_03012_),
    .B(net192));
 sg13g2_o21ai_1 _20688_ (.B1(_03140_),
    .Y(_01283_),
    .A1(net192),
    .A2(_03139_));
 sg13g2_nand2_1 _20689_ (.Y(_03141_),
    .A(net673),
    .B(\mem.mem_internal.code_mem[231][2] ));
 sg13g2_nand2_1 _20690_ (.Y(_03142_),
    .A(_03015_),
    .B(_03136_));
 sg13g2_o21ai_1 _20691_ (.B1(_03142_),
    .Y(_01284_),
    .A1(net192),
    .A2(_03141_));
 sg13g2_nand2_1 _20692_ (.Y(_03143_),
    .A(net673),
    .B(\mem.mem_internal.code_mem[231][3] ));
 sg13g2_nand2_1 _20693_ (.Y(_03144_),
    .A(_03018_),
    .B(_03136_));
 sg13g2_o21ai_1 _20694_ (.B1(_03144_),
    .Y(_01285_),
    .A1(net192),
    .A2(_03143_));
 sg13g2_nand2_1 _20695_ (.Y(_03145_),
    .A(_03127_),
    .B(\mem.mem_internal.code_mem[231][4] ));
 sg13g2_nand2_1 _20696_ (.Y(_03146_),
    .A(_03021_),
    .B(_03136_));
 sg13g2_o21ai_1 _20697_ (.B1(_03146_),
    .Y(_01286_),
    .A1(_03137_),
    .A2(_03145_));
 sg13g2_nand2_1 _20698_ (.Y(_03147_),
    .A(_03127_),
    .B(\mem.mem_internal.code_mem[231][5] ));
 sg13g2_nand2_1 _20699_ (.Y(_03148_),
    .A(_03024_),
    .B(_03136_));
 sg13g2_o21ai_1 _20700_ (.B1(_03148_),
    .Y(_01287_),
    .A1(_03137_),
    .A2(_03147_));
 sg13g2_nand2_1 _20701_ (.Y(_03149_),
    .A(net673),
    .B(\mem.mem_internal.code_mem[231][6] ));
 sg13g2_nand2_1 _20702_ (.Y(_03150_),
    .A(_03027_),
    .B(_03136_));
 sg13g2_o21ai_1 _20703_ (.B1(_03150_),
    .Y(_01288_),
    .A1(net192),
    .A2(_03149_));
 sg13g2_nand2_1 _20704_ (.Y(_03151_),
    .A(net673),
    .B(\mem.mem_internal.code_mem[231][7] ));
 sg13g2_nand2_1 _20705_ (.Y(_03152_),
    .A(_03030_),
    .B(_03136_));
 sg13g2_o21ai_1 _20706_ (.B1(_03152_),
    .Y(_01289_),
    .A1(net192),
    .A2(_03151_));
 sg13g2_nand2_1 _20707_ (.Y(_03153_),
    .A(net840),
    .B(\mem.mem_internal.code_mem[232][0] ));
 sg13g2_nor2_1 _20708_ (.A(net778),
    .B(net460),
    .Y(_03154_));
 sg13g2_buf_2 _20709_ (.A(_03154_),
    .X(_03155_));
 sg13g2_buf_1 _20710_ (.A(_03155_),
    .X(_03156_));
 sg13g2_nand2_1 _20711_ (.Y(_03157_),
    .A(net1078),
    .B(net191));
 sg13g2_o21ai_1 _20712_ (.B1(_03157_),
    .Y(_01290_),
    .A1(_03153_),
    .A2(net191));
 sg13g2_buf_1 _20713_ (.A(_03043_),
    .X(_03158_));
 sg13g2_nand2_1 _20714_ (.Y(_03159_),
    .A(net672),
    .B(\mem.mem_internal.code_mem[232][1] ));
 sg13g2_nand2_1 _20715_ (.Y(_03160_),
    .A(net1077),
    .B(net191));
 sg13g2_o21ai_1 _20716_ (.B1(_03160_),
    .Y(_01291_),
    .A1(net191),
    .A2(_03159_));
 sg13g2_nand2_1 _20717_ (.Y(_03161_),
    .A(net672),
    .B(\mem.mem_internal.code_mem[232][2] ));
 sg13g2_nand2_1 _20718_ (.Y(_03162_),
    .A(net1076),
    .B(_03155_));
 sg13g2_o21ai_1 _20719_ (.B1(_03162_),
    .Y(_01292_),
    .A1(_03156_),
    .A2(_03161_));
 sg13g2_nand2_1 _20720_ (.Y(_03163_),
    .A(net672),
    .B(\mem.mem_internal.code_mem[232][3] ));
 sg13g2_nand2_1 _20721_ (.Y(_03164_),
    .A(net1075),
    .B(_03155_));
 sg13g2_o21ai_1 _20722_ (.B1(_03164_),
    .Y(_01293_),
    .A1(net191),
    .A2(_03163_));
 sg13g2_nand2_1 _20723_ (.Y(_03165_),
    .A(_03158_),
    .B(\mem.mem_internal.code_mem[232][4] ));
 sg13g2_nand2_1 _20724_ (.Y(_03166_),
    .A(net1074),
    .B(_03155_));
 sg13g2_o21ai_1 _20725_ (.B1(_03166_),
    .Y(_01294_),
    .A1(net191),
    .A2(_03165_));
 sg13g2_nand2_1 _20726_ (.Y(_03167_),
    .A(_03158_),
    .B(\mem.mem_internal.code_mem[232][5] ));
 sg13g2_nand2_1 _20727_ (.Y(_03168_),
    .A(net1073),
    .B(_03155_));
 sg13g2_o21ai_1 _20728_ (.B1(_03168_),
    .Y(_01295_),
    .A1(net191),
    .A2(_03167_));
 sg13g2_nand2_1 _20729_ (.Y(_03169_),
    .A(net672),
    .B(\mem.mem_internal.code_mem[232][6] ));
 sg13g2_nand2_1 _20730_ (.Y(_03170_),
    .A(net1072),
    .B(_03155_));
 sg13g2_o21ai_1 _20731_ (.B1(_03170_),
    .Y(_01296_),
    .A1(_03156_),
    .A2(_03169_));
 sg13g2_nand2_1 _20732_ (.Y(_03171_),
    .A(net672),
    .B(\mem.mem_internal.code_mem[232][7] ));
 sg13g2_nand2_1 _20733_ (.Y(_03172_),
    .A(net1071),
    .B(_03155_));
 sg13g2_o21ai_1 _20734_ (.B1(_03172_),
    .Y(_01297_),
    .A1(net191),
    .A2(_03171_));
 sg13g2_nand2_1 _20735_ (.Y(_03173_),
    .A(net840),
    .B(\mem.mem_internal.code_mem[233][0] ));
 sg13g2_nor2_1 _20736_ (.A(_10422_),
    .B(net460),
    .Y(_03174_));
 sg13g2_buf_2 _20737_ (.A(_03174_),
    .X(_03175_));
 sg13g2_buf_1 _20738_ (.A(_03175_),
    .X(_03176_));
 sg13g2_nand2_1 _20739_ (.Y(_03177_),
    .A(net1078),
    .B(net190));
 sg13g2_o21ai_1 _20740_ (.B1(_03177_),
    .Y(_01298_),
    .A1(_03173_),
    .A2(net190));
 sg13g2_nand2_1 _20741_ (.Y(_03178_),
    .A(net672),
    .B(\mem.mem_internal.code_mem[233][1] ));
 sg13g2_nand2_1 _20742_ (.Y(_03179_),
    .A(net1077),
    .B(net190));
 sg13g2_o21ai_1 _20743_ (.B1(_03179_),
    .Y(_01299_),
    .A1(net190),
    .A2(_03178_));
 sg13g2_nand2_1 _20744_ (.Y(_03180_),
    .A(net672),
    .B(\mem.mem_internal.code_mem[233][2] ));
 sg13g2_nand2_1 _20745_ (.Y(_03181_),
    .A(net1076),
    .B(_03175_));
 sg13g2_o21ai_1 _20746_ (.B1(_03181_),
    .Y(_01300_),
    .A1(_03176_),
    .A2(_03180_));
 sg13g2_nand2_1 _20747_ (.Y(_03182_),
    .A(net672),
    .B(\mem.mem_internal.code_mem[233][3] ));
 sg13g2_nand2_1 _20748_ (.Y(_03183_),
    .A(net1075),
    .B(_03175_));
 sg13g2_o21ai_1 _20749_ (.B1(_03183_),
    .Y(_01301_),
    .A1(net190),
    .A2(_03182_));
 sg13g2_buf_1 _20750_ (.A(_03043_),
    .X(_03184_));
 sg13g2_nand2_1 _20751_ (.Y(_03185_),
    .A(_03184_),
    .B(\mem.mem_internal.code_mem[233][4] ));
 sg13g2_nand2_1 _20752_ (.Y(_03186_),
    .A(net1074),
    .B(_03175_));
 sg13g2_o21ai_1 _20753_ (.B1(_03186_),
    .Y(_01302_),
    .A1(net190),
    .A2(_03185_));
 sg13g2_nand2_1 _20754_ (.Y(_03187_),
    .A(net671),
    .B(\mem.mem_internal.code_mem[233][5] ));
 sg13g2_nand2_1 _20755_ (.Y(_03188_),
    .A(net1073),
    .B(_03175_));
 sg13g2_o21ai_1 _20756_ (.B1(_03188_),
    .Y(_01303_),
    .A1(net190),
    .A2(_03187_));
 sg13g2_nand2_1 _20757_ (.Y(_03189_),
    .A(net671),
    .B(\mem.mem_internal.code_mem[233][6] ));
 sg13g2_nand2_1 _20758_ (.Y(_03190_),
    .A(net1072),
    .B(_03175_));
 sg13g2_o21ai_1 _20759_ (.B1(_03190_),
    .Y(_01304_),
    .A1(_03176_),
    .A2(_03189_));
 sg13g2_nand2_1 _20760_ (.Y(_03191_),
    .A(net671),
    .B(\mem.mem_internal.code_mem[233][7] ));
 sg13g2_nand2_1 _20761_ (.Y(_03192_),
    .A(net1071),
    .B(_03175_));
 sg13g2_o21ai_1 _20762_ (.B1(_03192_),
    .Y(_01305_),
    .A1(net190),
    .A2(_03191_));
 sg13g2_nand2_1 _20763_ (.Y(_03193_),
    .A(net840),
    .B(\mem.mem_internal.code_mem[234][0] ));
 sg13g2_nor2_1 _20764_ (.A(_10444_),
    .B(_02964_),
    .Y(_03194_));
 sg13g2_buf_2 _20765_ (.A(_03194_),
    .X(_03195_));
 sg13g2_buf_1 _20766_ (.A(_03195_),
    .X(_03196_));
 sg13g2_nand2_1 _20767_ (.Y(_03197_),
    .A(net1078),
    .B(_03196_));
 sg13g2_o21ai_1 _20768_ (.B1(_03197_),
    .Y(_01306_),
    .A1(_03193_),
    .A2(_03196_));
 sg13g2_nand2_1 _20769_ (.Y(_03198_),
    .A(net671),
    .B(\mem.mem_internal.code_mem[234][1] ));
 sg13g2_nand2_1 _20770_ (.Y(_03199_),
    .A(net1077),
    .B(net354));
 sg13g2_o21ai_1 _20771_ (.B1(_03199_),
    .Y(_01307_),
    .A1(net354),
    .A2(_03198_));
 sg13g2_nand2_1 _20772_ (.Y(_03200_),
    .A(net671),
    .B(\mem.mem_internal.code_mem[234][2] ));
 sg13g2_nand2_1 _20773_ (.Y(_03201_),
    .A(net1076),
    .B(_03195_));
 sg13g2_o21ai_1 _20774_ (.B1(_03201_),
    .Y(_01308_),
    .A1(net354),
    .A2(_03200_));
 sg13g2_nand2_1 _20775_ (.Y(_03202_),
    .A(net671),
    .B(\mem.mem_internal.code_mem[234][3] ));
 sg13g2_nand2_1 _20776_ (.Y(_03203_),
    .A(net1075),
    .B(_03195_));
 sg13g2_o21ai_1 _20777_ (.B1(_03203_),
    .Y(_01309_),
    .A1(net354),
    .A2(_03202_));
 sg13g2_nand2_1 _20778_ (.Y(_03204_),
    .A(_03184_),
    .B(\mem.mem_internal.code_mem[234][4] ));
 sg13g2_nand2_1 _20779_ (.Y(_03205_),
    .A(net1074),
    .B(_03195_));
 sg13g2_o21ai_1 _20780_ (.B1(_03205_),
    .Y(_01310_),
    .A1(net354),
    .A2(_03204_));
 sg13g2_nand2_1 _20781_ (.Y(_03206_),
    .A(net671),
    .B(\mem.mem_internal.code_mem[234][5] ));
 sg13g2_nand2_1 _20782_ (.Y(_03207_),
    .A(net1073),
    .B(_03195_));
 sg13g2_o21ai_1 _20783_ (.B1(_03207_),
    .Y(_01311_),
    .A1(net354),
    .A2(_03206_));
 sg13g2_nand2_1 _20784_ (.Y(_03208_),
    .A(net671),
    .B(\mem.mem_internal.code_mem[234][6] ));
 sg13g2_nand2_1 _20785_ (.Y(_03209_),
    .A(net1072),
    .B(_03195_));
 sg13g2_o21ai_1 _20786_ (.B1(_03209_),
    .Y(_01312_),
    .A1(net354),
    .A2(_03208_));
 sg13g2_buf_1 _20787_ (.A(_03043_),
    .X(_03210_));
 sg13g2_nand2_1 _20788_ (.Y(_03211_),
    .A(net670),
    .B(\mem.mem_internal.code_mem[234][7] ));
 sg13g2_nand2_1 _20789_ (.Y(_03212_),
    .A(net1071),
    .B(_03195_));
 sg13g2_o21ai_1 _20790_ (.B1(_03212_),
    .Y(_01313_),
    .A1(net354),
    .A2(_03211_));
 sg13g2_nand2_1 _20791_ (.Y(_03213_),
    .A(net840),
    .B(\mem.mem_internal.code_mem[235][0] ));
 sg13g2_nor2_1 _20792_ (.A(net775),
    .B(_02964_),
    .Y(_03214_));
 sg13g2_buf_2 _20793_ (.A(_03214_),
    .X(_03215_));
 sg13g2_buf_1 _20794_ (.A(_03215_),
    .X(_03216_));
 sg13g2_buf_1 _20795_ (.A(_12637_),
    .X(_03217_));
 sg13g2_nand2_1 _20796_ (.Y(_03218_),
    .A(net1070),
    .B(_03216_));
 sg13g2_o21ai_1 _20797_ (.B1(_03218_),
    .Y(_01314_),
    .A1(_03213_),
    .A2(net353));
 sg13g2_nand2_1 _20798_ (.Y(_03219_),
    .A(net670),
    .B(\mem.mem_internal.code_mem[235][1] ));
 sg13g2_buf_1 _20799_ (.A(_12641_),
    .X(_03220_));
 sg13g2_nand2_1 _20800_ (.Y(_03221_),
    .A(net1069),
    .B(net353));
 sg13g2_o21ai_1 _20801_ (.B1(_03221_),
    .Y(_01315_),
    .A1(net353),
    .A2(_03219_));
 sg13g2_nand2_1 _20802_ (.Y(_03222_),
    .A(net670),
    .B(\mem.mem_internal.code_mem[235][2] ));
 sg13g2_buf_1 _20803_ (.A(_12645_),
    .X(_03223_));
 sg13g2_nand2_1 _20804_ (.Y(_03224_),
    .A(net1068),
    .B(_03215_));
 sg13g2_o21ai_1 _20805_ (.B1(_03224_),
    .Y(_01316_),
    .A1(net353),
    .A2(_03222_));
 sg13g2_nand2_1 _20806_ (.Y(_03225_),
    .A(net670),
    .B(\mem.mem_internal.code_mem[235][3] ));
 sg13g2_buf_1 _20807_ (.A(_12649_),
    .X(_03226_));
 sg13g2_nand2_1 _20808_ (.Y(_03227_),
    .A(net1067),
    .B(_03215_));
 sg13g2_o21ai_1 _20809_ (.B1(_03227_),
    .Y(_01317_),
    .A1(net353),
    .A2(_03225_));
 sg13g2_nand2_1 _20810_ (.Y(_03228_),
    .A(_03210_),
    .B(\mem.mem_internal.code_mem[235][4] ));
 sg13g2_buf_1 _20811_ (.A(_12653_),
    .X(_03229_));
 sg13g2_nand2_1 _20812_ (.Y(_03230_),
    .A(net1066),
    .B(_03215_));
 sg13g2_o21ai_1 _20813_ (.B1(_03230_),
    .Y(_01318_),
    .A1(net353),
    .A2(_03228_));
 sg13g2_nand2_1 _20814_ (.Y(_03231_),
    .A(_03210_),
    .B(\mem.mem_internal.code_mem[235][5] ));
 sg13g2_buf_1 _20815_ (.A(_12657_),
    .X(_03232_));
 sg13g2_nand2_1 _20816_ (.Y(_03233_),
    .A(net1065),
    .B(_03215_));
 sg13g2_o21ai_1 _20817_ (.B1(_03233_),
    .Y(_01319_),
    .A1(net353),
    .A2(_03231_));
 sg13g2_nand2_1 _20818_ (.Y(_03234_),
    .A(net670),
    .B(\mem.mem_internal.code_mem[235][6] ));
 sg13g2_buf_1 _20819_ (.A(_12661_),
    .X(_03235_));
 sg13g2_nand2_1 _20820_ (.Y(_03236_),
    .A(net1064),
    .B(_03215_));
 sg13g2_o21ai_1 _20821_ (.B1(_03236_),
    .Y(_01320_),
    .A1(_03216_),
    .A2(_03234_));
 sg13g2_nand2_1 _20822_ (.Y(_03237_),
    .A(net670),
    .B(\mem.mem_internal.code_mem[235][7] ));
 sg13g2_buf_1 _20823_ (.A(_12665_),
    .X(_03238_));
 sg13g2_nand2_1 _20824_ (.Y(_03239_),
    .A(_03238_),
    .B(_03215_));
 sg13g2_o21ai_1 _20825_ (.B1(_03239_),
    .Y(_01321_),
    .A1(net353),
    .A2(_03237_));
 sg13g2_buf_1 _20826_ (.A(_12878_),
    .X(_03240_));
 sg13g2_nand2_1 _20827_ (.Y(_03241_),
    .A(net839),
    .B(\mem.mem_internal.code_mem[236][0] ));
 sg13g2_nor2_1 _20828_ (.A(_10491_),
    .B(_02964_),
    .Y(_03242_));
 sg13g2_buf_2 _20829_ (.A(_03242_),
    .X(_03243_));
 sg13g2_buf_1 _20830_ (.A(_03243_),
    .X(_03244_));
 sg13g2_nand2_1 _20831_ (.Y(_03245_),
    .A(net1070),
    .B(net352));
 sg13g2_o21ai_1 _20832_ (.B1(_03245_),
    .Y(_01322_),
    .A1(_03241_),
    .A2(net352));
 sg13g2_nand2_1 _20833_ (.Y(_03246_),
    .A(net670),
    .B(\mem.mem_internal.code_mem[236][1] ));
 sg13g2_nand2_1 _20834_ (.Y(_03247_),
    .A(net1069),
    .B(net352));
 sg13g2_o21ai_1 _20835_ (.B1(_03247_),
    .Y(_01323_),
    .A1(net352),
    .A2(_03246_));
 sg13g2_nand2_1 _20836_ (.Y(_03248_),
    .A(net670),
    .B(\mem.mem_internal.code_mem[236][2] ));
 sg13g2_nand2_1 _20837_ (.Y(_03249_),
    .A(net1068),
    .B(_03243_));
 sg13g2_o21ai_1 _20838_ (.B1(_03249_),
    .Y(_01324_),
    .A1(_03244_),
    .A2(_03248_));
 sg13g2_buf_1 _20839_ (.A(_03042_),
    .X(_03250_));
 sg13g2_buf_1 _20840_ (.A(_03250_),
    .X(_03251_));
 sg13g2_nand2_1 _20841_ (.Y(_03252_),
    .A(net669),
    .B(\mem.mem_internal.code_mem[236][3] ));
 sg13g2_nand2_1 _20842_ (.Y(_03253_),
    .A(net1067),
    .B(_03243_));
 sg13g2_o21ai_1 _20843_ (.B1(_03253_),
    .Y(_01325_),
    .A1(net352),
    .A2(_03252_));
 sg13g2_nand2_1 _20844_ (.Y(_03254_),
    .A(net669),
    .B(\mem.mem_internal.code_mem[236][4] ));
 sg13g2_nand2_1 _20845_ (.Y(_03255_),
    .A(net1066),
    .B(_03243_));
 sg13g2_o21ai_1 _20846_ (.B1(_03255_),
    .Y(_01326_),
    .A1(net352),
    .A2(_03254_));
 sg13g2_nand2_1 _20847_ (.Y(_03256_),
    .A(net669),
    .B(\mem.mem_internal.code_mem[236][5] ));
 sg13g2_nand2_1 _20848_ (.Y(_03257_),
    .A(net1065),
    .B(_03243_));
 sg13g2_o21ai_1 _20849_ (.B1(_03257_),
    .Y(_01327_),
    .A1(net352),
    .A2(_03256_));
 sg13g2_nand2_1 _20850_ (.Y(_03258_),
    .A(net669),
    .B(\mem.mem_internal.code_mem[236][6] ));
 sg13g2_nand2_1 _20851_ (.Y(_03259_),
    .A(net1064),
    .B(_03243_));
 sg13g2_o21ai_1 _20852_ (.B1(_03259_),
    .Y(_01328_),
    .A1(net352),
    .A2(_03258_));
 sg13g2_nand2_1 _20853_ (.Y(_03260_),
    .A(net669),
    .B(\mem.mem_internal.code_mem[236][7] ));
 sg13g2_nand2_1 _20854_ (.Y(_03261_),
    .A(net1063),
    .B(_03243_));
 sg13g2_o21ai_1 _20855_ (.B1(_03261_),
    .Y(_01329_),
    .A1(_03244_),
    .A2(_03260_));
 sg13g2_nand2_1 _20856_ (.Y(_03262_),
    .A(net839),
    .B(\mem.mem_internal.code_mem[237][0] ));
 sg13g2_nor2_1 _20857_ (.A(_10513_),
    .B(_02964_),
    .Y(_03263_));
 sg13g2_buf_2 _20858_ (.A(_03263_),
    .X(_03264_));
 sg13g2_buf_1 _20859_ (.A(_03264_),
    .X(_03265_));
 sg13g2_nand2_1 _20860_ (.Y(_03266_),
    .A(net1070),
    .B(_03265_));
 sg13g2_o21ai_1 _20861_ (.B1(_03266_),
    .Y(_01330_),
    .A1(_03262_),
    .A2(_03265_));
 sg13g2_nand2_1 _20862_ (.Y(_03267_),
    .A(net669),
    .B(\mem.mem_internal.code_mem[237][1] ));
 sg13g2_nand2_1 _20863_ (.Y(_03268_),
    .A(net1069),
    .B(net351));
 sg13g2_o21ai_1 _20864_ (.B1(_03268_),
    .Y(_01331_),
    .A1(net351),
    .A2(_03267_));
 sg13g2_nand2_1 _20865_ (.Y(_03269_),
    .A(_03251_),
    .B(\mem.mem_internal.code_mem[237][2] ));
 sg13g2_nand2_1 _20866_ (.Y(_03270_),
    .A(net1068),
    .B(_03264_));
 sg13g2_o21ai_1 _20867_ (.B1(_03270_),
    .Y(_01332_),
    .A1(net351),
    .A2(_03269_));
 sg13g2_nand2_1 _20868_ (.Y(_03271_),
    .A(net669),
    .B(\mem.mem_internal.code_mem[237][3] ));
 sg13g2_nand2_1 _20869_ (.Y(_03272_),
    .A(net1067),
    .B(_03264_));
 sg13g2_o21ai_1 _20870_ (.B1(_03272_),
    .Y(_01333_),
    .A1(net351),
    .A2(_03271_));
 sg13g2_nand2_1 _20871_ (.Y(_03273_),
    .A(_03251_),
    .B(\mem.mem_internal.code_mem[237][4] ));
 sg13g2_nand2_1 _20872_ (.Y(_03274_),
    .A(net1066),
    .B(_03264_));
 sg13g2_o21ai_1 _20873_ (.B1(_03274_),
    .Y(_01334_),
    .A1(net351),
    .A2(_03273_));
 sg13g2_nand2_1 _20874_ (.Y(_03275_),
    .A(net669),
    .B(\mem.mem_internal.code_mem[237][5] ));
 sg13g2_nand2_1 _20875_ (.Y(_03276_),
    .A(net1065),
    .B(_03264_));
 sg13g2_o21ai_1 _20876_ (.B1(_03276_),
    .Y(_01335_),
    .A1(net351),
    .A2(_03275_));
 sg13g2_buf_1 _20877_ (.A(_03250_),
    .X(_03277_));
 sg13g2_nand2_1 _20878_ (.Y(_03278_),
    .A(net668),
    .B(\mem.mem_internal.code_mem[237][6] ));
 sg13g2_nand2_1 _20879_ (.Y(_03279_),
    .A(net1064),
    .B(_03264_));
 sg13g2_o21ai_1 _20880_ (.B1(_03279_),
    .Y(_01336_),
    .A1(net351),
    .A2(_03278_));
 sg13g2_nand2_1 _20881_ (.Y(_03280_),
    .A(net668),
    .B(\mem.mem_internal.code_mem[237][7] ));
 sg13g2_nand2_1 _20882_ (.Y(_03281_),
    .A(net1063),
    .B(_03264_));
 sg13g2_o21ai_1 _20883_ (.B1(_03281_),
    .Y(_01337_),
    .A1(net351),
    .A2(_03280_));
 sg13g2_nand2_1 _20884_ (.Y(_03282_),
    .A(net839),
    .B(\mem.mem_internal.code_mem[238][0] ));
 sg13g2_nor2_1 _20885_ (.A(_10564_),
    .B(_02964_),
    .Y(_03283_));
 sg13g2_buf_2 _20886_ (.A(_03283_),
    .X(_03284_));
 sg13g2_buf_1 _20887_ (.A(_03284_),
    .X(_03285_));
 sg13g2_nand2_1 _20888_ (.Y(_03286_),
    .A(net1070),
    .B(net350));
 sg13g2_o21ai_1 _20889_ (.B1(_03286_),
    .Y(_01338_),
    .A1(_03282_),
    .A2(net350));
 sg13g2_nand2_1 _20890_ (.Y(_03287_),
    .A(net668),
    .B(\mem.mem_internal.code_mem[238][1] ));
 sg13g2_nand2_1 _20891_ (.Y(_03288_),
    .A(net1069),
    .B(net350));
 sg13g2_o21ai_1 _20892_ (.B1(_03288_),
    .Y(_01339_),
    .A1(net350),
    .A2(_03287_));
 sg13g2_nand2_1 _20893_ (.Y(_03289_),
    .A(_03277_),
    .B(\mem.mem_internal.code_mem[238][2] ));
 sg13g2_nand2_1 _20894_ (.Y(_03290_),
    .A(net1068),
    .B(_03284_));
 sg13g2_o21ai_1 _20895_ (.B1(_03290_),
    .Y(_01340_),
    .A1(net350),
    .A2(_03289_));
 sg13g2_nand2_1 _20896_ (.Y(_03291_),
    .A(net668),
    .B(\mem.mem_internal.code_mem[238][3] ));
 sg13g2_nand2_1 _20897_ (.Y(_03292_),
    .A(net1067),
    .B(_03284_));
 sg13g2_o21ai_1 _20898_ (.B1(_03292_),
    .Y(_01341_),
    .A1(net350),
    .A2(_03291_));
 sg13g2_nand2_1 _20899_ (.Y(_03293_),
    .A(_03277_),
    .B(\mem.mem_internal.code_mem[238][4] ));
 sg13g2_nand2_1 _20900_ (.Y(_03294_),
    .A(net1066),
    .B(_03284_));
 sg13g2_o21ai_1 _20901_ (.B1(_03294_),
    .Y(_01342_),
    .A1(net350),
    .A2(_03293_));
 sg13g2_nand2_1 _20902_ (.Y(_03295_),
    .A(net668),
    .B(\mem.mem_internal.code_mem[238][5] ));
 sg13g2_nand2_1 _20903_ (.Y(_03296_),
    .A(net1065),
    .B(_03284_));
 sg13g2_o21ai_1 _20904_ (.B1(_03296_),
    .Y(_01343_),
    .A1(net350),
    .A2(_03295_));
 sg13g2_nand2_1 _20905_ (.Y(_03297_),
    .A(net668),
    .B(\mem.mem_internal.code_mem[238][6] ));
 sg13g2_nand2_1 _20906_ (.Y(_03298_),
    .A(net1064),
    .B(_03284_));
 sg13g2_o21ai_1 _20907_ (.B1(_03298_),
    .Y(_01344_),
    .A1(_03285_),
    .A2(_03297_));
 sg13g2_nand2_1 _20908_ (.Y(_03299_),
    .A(net668),
    .B(\mem.mem_internal.code_mem[238][7] ));
 sg13g2_nand2_1 _20909_ (.Y(_03300_),
    .A(net1063),
    .B(_03284_));
 sg13g2_o21ai_1 _20910_ (.B1(_03300_),
    .Y(_01345_),
    .A1(_03285_),
    .A2(_03299_));
 sg13g2_nand2_1 _20911_ (.Y(_03301_),
    .A(net839),
    .B(\mem.mem_internal.code_mem[239][0] ));
 sg13g2_nor2_1 _20912_ (.A(_10586_),
    .B(_02964_),
    .Y(_03302_));
 sg13g2_buf_2 _20913_ (.A(_03302_),
    .X(_03303_));
 sg13g2_buf_1 _20914_ (.A(_03303_),
    .X(_03304_));
 sg13g2_nand2_1 _20915_ (.Y(_03305_),
    .A(net1070),
    .B(net349));
 sg13g2_o21ai_1 _20916_ (.B1(_03305_),
    .Y(_01346_),
    .A1(_03301_),
    .A2(net349));
 sg13g2_nand2_1 _20917_ (.Y(_03306_),
    .A(net668),
    .B(\mem.mem_internal.code_mem[239][1] ));
 sg13g2_nand2_1 _20918_ (.Y(_03307_),
    .A(net1069),
    .B(net349));
 sg13g2_o21ai_1 _20919_ (.B1(_03307_),
    .Y(_01347_),
    .A1(net349),
    .A2(_03306_));
 sg13g2_buf_1 _20920_ (.A(_03250_),
    .X(_03308_));
 sg13g2_nand2_1 _20921_ (.Y(_03309_),
    .A(net667),
    .B(\mem.mem_internal.code_mem[239][2] ));
 sg13g2_nand2_1 _20922_ (.Y(_03310_),
    .A(net1068),
    .B(_03303_));
 sg13g2_o21ai_1 _20923_ (.B1(_03310_),
    .Y(_01348_),
    .A1(net349),
    .A2(_03309_));
 sg13g2_nand2_1 _20924_ (.Y(_03311_),
    .A(net667),
    .B(\mem.mem_internal.code_mem[239][3] ));
 sg13g2_nand2_1 _20925_ (.Y(_03312_),
    .A(net1067),
    .B(_03303_));
 sg13g2_o21ai_1 _20926_ (.B1(_03312_),
    .Y(_01349_),
    .A1(net349),
    .A2(_03311_));
 sg13g2_nand2_1 _20927_ (.Y(_03313_),
    .A(net667),
    .B(\mem.mem_internal.code_mem[239][4] ));
 sg13g2_nand2_1 _20928_ (.Y(_03314_),
    .A(net1066),
    .B(_03303_));
 sg13g2_o21ai_1 _20929_ (.B1(_03314_),
    .Y(_01350_),
    .A1(net349),
    .A2(_03313_));
 sg13g2_nand2_1 _20930_ (.Y(_03315_),
    .A(net667),
    .B(\mem.mem_internal.code_mem[239][5] ));
 sg13g2_nand2_1 _20931_ (.Y(_03316_),
    .A(net1065),
    .B(_03303_));
 sg13g2_o21ai_1 _20932_ (.B1(_03316_),
    .Y(_01351_),
    .A1(net349),
    .A2(_03315_));
 sg13g2_nand2_1 _20933_ (.Y(_03317_),
    .A(net667),
    .B(\mem.mem_internal.code_mem[239][6] ));
 sg13g2_nand2_1 _20934_ (.Y(_03318_),
    .A(_03235_),
    .B(_03303_));
 sg13g2_o21ai_1 _20935_ (.B1(_03318_),
    .Y(_01352_),
    .A1(_03304_),
    .A2(_03317_));
 sg13g2_nand2_1 _20936_ (.Y(_03319_),
    .A(net667),
    .B(\mem.mem_internal.code_mem[239][7] ));
 sg13g2_nand2_1 _20937_ (.Y(_03320_),
    .A(net1063),
    .B(_03303_));
 sg13g2_o21ai_1 _20938_ (.B1(_03320_),
    .Y(_01353_),
    .A1(_03304_),
    .A2(_03319_));
 sg13g2_nand2_1 _20939_ (.Y(_03321_),
    .A(_03240_),
    .B(\mem.mem_internal.code_mem[23][0] ));
 sg13g2_nor2_1 _20940_ (.A(_10372_),
    .B(_11947_),
    .Y(_03322_));
 sg13g2_buf_2 _20941_ (.A(_03322_),
    .X(_03323_));
 sg13g2_buf_1 _20942_ (.A(_03323_),
    .X(_03324_));
 sg13g2_nand2_1 _20943_ (.Y(_03325_),
    .A(net1070),
    .B(net189));
 sg13g2_o21ai_1 _20944_ (.B1(_03325_),
    .Y(_01354_),
    .A1(_03321_),
    .A2(net189));
 sg13g2_nand2_1 _20945_ (.Y(_03326_),
    .A(net667),
    .B(\mem.mem_internal.code_mem[23][1] ));
 sg13g2_nand2_1 _20946_ (.Y(_03327_),
    .A(net1069),
    .B(_03324_));
 sg13g2_o21ai_1 _20947_ (.B1(_03327_),
    .Y(_01355_),
    .A1(net189),
    .A2(_03326_));
 sg13g2_nand2_1 _20948_ (.Y(_03328_),
    .A(net667),
    .B(\mem.mem_internal.code_mem[23][2] ));
 sg13g2_nand2_1 _20949_ (.Y(_03329_),
    .A(net1068),
    .B(_03323_));
 sg13g2_o21ai_1 _20950_ (.B1(_03329_),
    .Y(_01356_),
    .A1(net189),
    .A2(_03328_));
 sg13g2_nand2_1 _20951_ (.Y(_03330_),
    .A(_03308_),
    .B(\mem.mem_internal.code_mem[23][3] ));
 sg13g2_nand2_1 _20952_ (.Y(_03331_),
    .A(net1067),
    .B(_03323_));
 sg13g2_o21ai_1 _20953_ (.B1(_03331_),
    .Y(_01357_),
    .A1(net189),
    .A2(_03330_));
 sg13g2_nand2_1 _20954_ (.Y(_03332_),
    .A(_03308_),
    .B(\mem.mem_internal.code_mem[23][4] ));
 sg13g2_nand2_1 _20955_ (.Y(_03333_),
    .A(net1066),
    .B(_03323_));
 sg13g2_o21ai_1 _20956_ (.B1(_03333_),
    .Y(_01358_),
    .A1(net189),
    .A2(_03332_));
 sg13g2_buf_1 _20957_ (.A(_03250_),
    .X(_03334_));
 sg13g2_nand2_1 _20958_ (.Y(_03335_),
    .A(net666),
    .B(\mem.mem_internal.code_mem[23][5] ));
 sg13g2_nand2_1 _20959_ (.Y(_03336_),
    .A(net1065),
    .B(_03323_));
 sg13g2_o21ai_1 _20960_ (.B1(_03336_),
    .Y(_01359_),
    .A1(net189),
    .A2(_03335_));
 sg13g2_nand2_1 _20961_ (.Y(_03337_),
    .A(net666),
    .B(\mem.mem_internal.code_mem[23][6] ));
 sg13g2_nand2_1 _20962_ (.Y(_03338_),
    .A(net1064),
    .B(_03323_));
 sg13g2_o21ai_1 _20963_ (.B1(_03338_),
    .Y(_01360_),
    .A1(net189),
    .A2(_03337_));
 sg13g2_nand2_1 _20964_ (.Y(_03339_),
    .A(net666),
    .B(\mem.mem_internal.code_mem[23][7] ));
 sg13g2_nand2_1 _20965_ (.Y(_03340_),
    .A(_03238_),
    .B(_03323_));
 sg13g2_o21ai_1 _20966_ (.B1(_03340_),
    .Y(_01361_),
    .A1(_03324_),
    .A2(_03339_));
 sg13g2_nand3_1 _20967_ (.B(net1296),
    .C(_10607_),
    .A(net1297),
    .Y(_03341_));
 sg13g2_buf_2 _20968_ (.A(_03341_),
    .X(_03342_));
 sg13g2_buf_1 _20969_ (.A(_03342_),
    .X(_03343_));
 sg13g2_nor2_1 _20970_ (.A(net529),
    .B(net459),
    .Y(_03344_));
 sg13g2_buf_2 _20971_ (.A(_03344_),
    .X(_03345_));
 sg13g2_buf_1 _20972_ (.A(_03345_),
    .X(_03346_));
 sg13g2_nand2_1 _20973_ (.Y(_03347_),
    .A(net666),
    .B(\mem.mem_internal.code_mem[240][0] ));
 sg13g2_nand2_1 _20974_ (.Y(_03348_),
    .A(net1070),
    .B(net188));
 sg13g2_o21ai_1 _20975_ (.B1(_03348_),
    .Y(_01362_),
    .A1(net188),
    .A2(_03347_));
 sg13g2_nand2_1 _20976_ (.Y(_03349_),
    .A(net666),
    .B(\mem.mem_internal.code_mem[240][1] ));
 sg13g2_nand2_1 _20977_ (.Y(_03350_),
    .A(net1069),
    .B(net188));
 sg13g2_o21ai_1 _20978_ (.B1(_03350_),
    .Y(_01363_),
    .A1(net188),
    .A2(_03349_));
 sg13g2_nand2_1 _20979_ (.Y(_03351_),
    .A(net666),
    .B(\mem.mem_internal.code_mem[240][2] ));
 sg13g2_nand2_1 _20980_ (.Y(_03352_),
    .A(net1068),
    .B(_03345_));
 sg13g2_o21ai_1 _20981_ (.B1(_03352_),
    .Y(_01364_),
    .A1(net188),
    .A2(_03351_));
 sg13g2_nand2_1 _20982_ (.Y(_03353_),
    .A(net666),
    .B(\mem.mem_internal.code_mem[240][3] ));
 sg13g2_nand2_1 _20983_ (.Y(_03354_),
    .A(net1067),
    .B(_03345_));
 sg13g2_o21ai_1 _20984_ (.B1(_03354_),
    .Y(_01365_),
    .A1(net188),
    .A2(_03353_));
 sg13g2_nand2_1 _20985_ (.Y(_03355_),
    .A(net666),
    .B(\mem.mem_internal.code_mem[240][4] ));
 sg13g2_nand2_1 _20986_ (.Y(_03356_),
    .A(net1066),
    .B(_03345_));
 sg13g2_o21ai_1 _20987_ (.B1(_03356_),
    .Y(_01366_),
    .A1(_03346_),
    .A2(_03355_));
 sg13g2_nand2_1 _20988_ (.Y(_03357_),
    .A(_03334_),
    .B(\mem.mem_internal.code_mem[240][5] ));
 sg13g2_nand2_1 _20989_ (.Y(_03358_),
    .A(net1065),
    .B(_03345_));
 sg13g2_o21ai_1 _20990_ (.B1(_03358_),
    .Y(_01367_),
    .A1(net188),
    .A2(_03357_));
 sg13g2_nand2_1 _20991_ (.Y(_03359_),
    .A(_03334_),
    .B(\mem.mem_internal.code_mem[240][6] ));
 sg13g2_nand2_1 _20992_ (.Y(_03360_),
    .A(net1064),
    .B(_03345_));
 sg13g2_o21ai_1 _20993_ (.B1(_03360_),
    .Y(_01368_),
    .A1(_03346_),
    .A2(_03359_));
 sg13g2_buf_1 _20994_ (.A(_03250_),
    .X(_03361_));
 sg13g2_nand2_1 _20995_ (.Y(_03362_),
    .A(net665),
    .B(\mem.mem_internal.code_mem[240][7] ));
 sg13g2_nand2_1 _20996_ (.Y(_03363_),
    .A(net1063),
    .B(_03345_));
 sg13g2_o21ai_1 _20997_ (.B1(_03363_),
    .Y(_01369_),
    .A1(net188),
    .A2(_03362_));
 sg13g2_nor2_1 _20998_ (.A(_10633_),
    .B(net459),
    .Y(_03364_));
 sg13g2_buf_2 _20999_ (.A(_03364_),
    .X(_03365_));
 sg13g2_buf_1 _21000_ (.A(_03365_),
    .X(_03366_));
 sg13g2_nand2_1 _21001_ (.Y(_03367_),
    .A(net665),
    .B(\mem.mem_internal.code_mem[241][0] ));
 sg13g2_nand2_1 _21002_ (.Y(_03368_),
    .A(net1070),
    .B(net187));
 sg13g2_o21ai_1 _21003_ (.B1(_03368_),
    .Y(_01370_),
    .A1(net187),
    .A2(_03367_));
 sg13g2_nand2_1 _21004_ (.Y(_03369_),
    .A(net665),
    .B(\mem.mem_internal.code_mem[241][1] ));
 sg13g2_nand2_1 _21005_ (.Y(_03370_),
    .A(net1069),
    .B(net187));
 sg13g2_o21ai_1 _21006_ (.B1(_03370_),
    .Y(_01371_),
    .A1(net187),
    .A2(_03369_));
 sg13g2_nand2_1 _21007_ (.Y(_03371_),
    .A(net665),
    .B(\mem.mem_internal.code_mem[241][2] ));
 sg13g2_nand2_1 _21008_ (.Y(_03372_),
    .A(net1068),
    .B(_03365_));
 sg13g2_o21ai_1 _21009_ (.B1(_03372_),
    .Y(_01372_),
    .A1(net187),
    .A2(_03371_));
 sg13g2_nand2_1 _21010_ (.Y(_03373_),
    .A(net665),
    .B(\mem.mem_internal.code_mem[241][3] ));
 sg13g2_nand2_1 _21011_ (.Y(_03374_),
    .A(net1067),
    .B(_03365_));
 sg13g2_o21ai_1 _21012_ (.B1(_03374_),
    .Y(_01373_),
    .A1(net187),
    .A2(_03373_));
 sg13g2_nand2_1 _21013_ (.Y(_03375_),
    .A(_03361_),
    .B(\mem.mem_internal.code_mem[241][4] ));
 sg13g2_nand2_1 _21014_ (.Y(_03376_),
    .A(net1066),
    .B(_03365_));
 sg13g2_o21ai_1 _21015_ (.B1(_03376_),
    .Y(_01374_),
    .A1(_03366_),
    .A2(_03375_));
 sg13g2_nand2_1 _21016_ (.Y(_03377_),
    .A(_03361_),
    .B(\mem.mem_internal.code_mem[241][5] ));
 sg13g2_nand2_1 _21017_ (.Y(_03378_),
    .A(net1065),
    .B(_03365_));
 sg13g2_o21ai_1 _21018_ (.B1(_03378_),
    .Y(_01375_),
    .A1(_03366_),
    .A2(_03377_));
 sg13g2_nand2_1 _21019_ (.Y(_03379_),
    .A(net665),
    .B(\mem.mem_internal.code_mem[241][6] ));
 sg13g2_nand2_1 _21020_ (.Y(_03380_),
    .A(net1064),
    .B(_03365_));
 sg13g2_o21ai_1 _21021_ (.B1(_03380_),
    .Y(_01376_),
    .A1(net187),
    .A2(_03379_));
 sg13g2_nand2_1 _21022_ (.Y(_03381_),
    .A(net665),
    .B(\mem.mem_internal.code_mem[241][7] ));
 sg13g2_nand2_1 _21023_ (.Y(_03382_),
    .A(net1063),
    .B(_03365_));
 sg13g2_o21ai_1 _21024_ (.B1(_03382_),
    .Y(_01377_),
    .A1(net187),
    .A2(_03381_));
 sg13g2_nor2_1 _21025_ (.A(_10657_),
    .B(_03343_),
    .Y(_03383_));
 sg13g2_buf_2 _21026_ (.A(_03383_),
    .X(_03384_));
 sg13g2_buf_1 _21027_ (.A(_03384_),
    .X(_03385_));
 sg13g2_nand2_1 _21028_ (.Y(_03386_),
    .A(net665),
    .B(\mem.mem_internal.code_mem[242][0] ));
 sg13g2_nand2_1 _21029_ (.Y(_03387_),
    .A(_03217_),
    .B(net186));
 sg13g2_o21ai_1 _21030_ (.B1(_03387_),
    .Y(_01378_),
    .A1(net186),
    .A2(_03386_));
 sg13g2_buf_1 _21031_ (.A(_03250_),
    .X(_03388_));
 sg13g2_nand2_1 _21032_ (.Y(_03389_),
    .A(net664),
    .B(\mem.mem_internal.code_mem[242][1] ));
 sg13g2_nand2_1 _21033_ (.Y(_03390_),
    .A(_03220_),
    .B(net186));
 sg13g2_o21ai_1 _21034_ (.B1(_03390_),
    .Y(_01379_),
    .A1(net186),
    .A2(_03389_));
 sg13g2_nand2_1 _21035_ (.Y(_03391_),
    .A(net664),
    .B(\mem.mem_internal.code_mem[242][2] ));
 sg13g2_nand2_1 _21036_ (.Y(_03392_),
    .A(_03223_),
    .B(_03384_));
 sg13g2_o21ai_1 _21037_ (.B1(_03392_),
    .Y(_01380_),
    .A1(net186),
    .A2(_03391_));
 sg13g2_nand2_1 _21038_ (.Y(_03393_),
    .A(net664),
    .B(\mem.mem_internal.code_mem[242][3] ));
 sg13g2_nand2_1 _21039_ (.Y(_03394_),
    .A(_03226_),
    .B(_03384_));
 sg13g2_o21ai_1 _21040_ (.B1(_03394_),
    .Y(_01381_),
    .A1(net186),
    .A2(_03393_));
 sg13g2_nand2_1 _21041_ (.Y(_03395_),
    .A(_03388_),
    .B(\mem.mem_internal.code_mem[242][4] ));
 sg13g2_nand2_1 _21042_ (.Y(_03396_),
    .A(_03229_),
    .B(_03384_));
 sg13g2_o21ai_1 _21043_ (.B1(_03396_),
    .Y(_01382_),
    .A1(_03385_),
    .A2(_03395_));
 sg13g2_nand2_1 _21044_ (.Y(_03397_),
    .A(_03388_),
    .B(\mem.mem_internal.code_mem[242][5] ));
 sg13g2_nand2_1 _21045_ (.Y(_03398_),
    .A(_03232_),
    .B(_03384_));
 sg13g2_o21ai_1 _21046_ (.B1(_03398_),
    .Y(_01383_),
    .A1(_03385_),
    .A2(_03397_));
 sg13g2_nand2_1 _21047_ (.Y(_03399_),
    .A(net664),
    .B(\mem.mem_internal.code_mem[242][6] ));
 sg13g2_nand2_1 _21048_ (.Y(_03400_),
    .A(net1064),
    .B(_03384_));
 sg13g2_o21ai_1 _21049_ (.B1(_03400_),
    .Y(_01384_),
    .A1(net186),
    .A2(_03399_));
 sg13g2_nand2_1 _21050_ (.Y(_03401_),
    .A(net664),
    .B(\mem.mem_internal.code_mem[242][7] ));
 sg13g2_nand2_1 _21051_ (.Y(_03402_),
    .A(net1063),
    .B(_03384_));
 sg13g2_o21ai_1 _21052_ (.B1(_03402_),
    .Y(_01385_),
    .A1(net186),
    .A2(_03401_));
 sg13g2_nor2_1 _21053_ (.A(_10680_),
    .B(_03343_),
    .Y(_03403_));
 sg13g2_buf_2 _21054_ (.A(_03403_),
    .X(_03404_));
 sg13g2_buf_1 _21055_ (.A(_03404_),
    .X(_03405_));
 sg13g2_nand2_1 _21056_ (.Y(_03406_),
    .A(net664),
    .B(\mem.mem_internal.code_mem[243][0] ));
 sg13g2_nand2_1 _21057_ (.Y(_03407_),
    .A(_03217_),
    .B(net185));
 sg13g2_o21ai_1 _21058_ (.B1(_03407_),
    .Y(_01386_),
    .A1(net185),
    .A2(_03406_));
 sg13g2_nand2_1 _21059_ (.Y(_03408_),
    .A(net664),
    .B(\mem.mem_internal.code_mem[243][1] ));
 sg13g2_nand2_1 _21060_ (.Y(_03409_),
    .A(_03220_),
    .B(net185));
 sg13g2_o21ai_1 _21061_ (.B1(_03409_),
    .Y(_01387_),
    .A1(net185),
    .A2(_03408_));
 sg13g2_nand2_1 _21062_ (.Y(_03410_),
    .A(net664),
    .B(\mem.mem_internal.code_mem[243][2] ));
 sg13g2_nand2_1 _21063_ (.Y(_03411_),
    .A(_03223_),
    .B(_03404_));
 sg13g2_o21ai_1 _21064_ (.B1(_03411_),
    .Y(_01388_),
    .A1(net185),
    .A2(_03410_));
 sg13g2_buf_1 _21065_ (.A(_03250_),
    .X(_03412_));
 sg13g2_nand2_1 _21066_ (.Y(_03413_),
    .A(net663),
    .B(\mem.mem_internal.code_mem[243][3] ));
 sg13g2_nand2_1 _21067_ (.Y(_03414_),
    .A(_03226_),
    .B(_03404_));
 sg13g2_o21ai_1 _21068_ (.B1(_03414_),
    .Y(_01389_),
    .A1(net185),
    .A2(_03413_));
 sg13g2_nand2_1 _21069_ (.Y(_03415_),
    .A(net663),
    .B(\mem.mem_internal.code_mem[243][4] ));
 sg13g2_nand2_1 _21070_ (.Y(_03416_),
    .A(_03229_),
    .B(_03404_));
 sg13g2_o21ai_1 _21071_ (.B1(_03416_),
    .Y(_01390_),
    .A1(_03405_),
    .A2(_03415_));
 sg13g2_nand2_1 _21072_ (.Y(_03417_),
    .A(_03412_),
    .B(\mem.mem_internal.code_mem[243][5] ));
 sg13g2_nand2_1 _21073_ (.Y(_03418_),
    .A(_03232_),
    .B(_03404_));
 sg13g2_o21ai_1 _21074_ (.B1(_03418_),
    .Y(_01391_),
    .A1(_03405_),
    .A2(_03417_));
 sg13g2_nand2_1 _21075_ (.Y(_03419_),
    .A(_03412_),
    .B(\mem.mem_internal.code_mem[243][6] ));
 sg13g2_nand2_1 _21076_ (.Y(_03420_),
    .A(_03235_),
    .B(_03404_));
 sg13g2_o21ai_1 _21077_ (.B1(_03420_),
    .Y(_01392_),
    .A1(net185),
    .A2(_03419_));
 sg13g2_nand2_1 _21078_ (.Y(_03421_),
    .A(net663),
    .B(\mem.mem_internal.code_mem[243][7] ));
 sg13g2_nand2_1 _21079_ (.Y(_03422_),
    .A(net1063),
    .B(_03404_));
 sg13g2_o21ai_1 _21080_ (.B1(_03422_),
    .Y(_01393_),
    .A1(net185),
    .A2(_03421_));
 sg13g2_nor2_1 _21081_ (.A(net556),
    .B(net459),
    .Y(_03423_));
 sg13g2_buf_2 _21082_ (.A(_03423_),
    .X(_03424_));
 sg13g2_buf_1 _21083_ (.A(_03424_),
    .X(_03425_));
 sg13g2_nand2_1 _21084_ (.Y(_03426_),
    .A(net663),
    .B(\mem.mem_internal.code_mem[244][0] ));
 sg13g2_buf_1 _21085_ (.A(_12637_),
    .X(_03427_));
 sg13g2_nand2_1 _21086_ (.Y(_03428_),
    .A(net1062),
    .B(net184));
 sg13g2_o21ai_1 _21087_ (.B1(_03428_),
    .Y(_01394_),
    .A1(net184),
    .A2(_03426_));
 sg13g2_nand2_1 _21088_ (.Y(_03429_),
    .A(net663),
    .B(\mem.mem_internal.code_mem[244][1] ));
 sg13g2_buf_1 _21089_ (.A(_12641_),
    .X(_03430_));
 sg13g2_nand2_1 _21090_ (.Y(_03431_),
    .A(net1061),
    .B(net184));
 sg13g2_o21ai_1 _21091_ (.B1(_03431_),
    .Y(_01395_),
    .A1(net184),
    .A2(_03429_));
 sg13g2_nand2_1 _21092_ (.Y(_03432_),
    .A(net663),
    .B(\mem.mem_internal.code_mem[244][2] ));
 sg13g2_buf_1 _21093_ (.A(_12645_),
    .X(_03433_));
 sg13g2_nand2_1 _21094_ (.Y(_03434_),
    .A(net1060),
    .B(_03424_));
 sg13g2_o21ai_1 _21095_ (.B1(_03434_),
    .Y(_01396_),
    .A1(net184),
    .A2(_03432_));
 sg13g2_nand2_1 _21096_ (.Y(_03435_),
    .A(net663),
    .B(\mem.mem_internal.code_mem[244][3] ));
 sg13g2_buf_1 _21097_ (.A(_12649_),
    .X(_03436_));
 sg13g2_nand2_1 _21098_ (.Y(_03437_),
    .A(net1059),
    .B(_03424_));
 sg13g2_o21ai_1 _21099_ (.B1(_03437_),
    .Y(_01397_),
    .A1(net184),
    .A2(_03435_));
 sg13g2_nand2_1 _21100_ (.Y(_03438_),
    .A(net663),
    .B(\mem.mem_internal.code_mem[244][4] ));
 sg13g2_buf_1 _21101_ (.A(_12653_),
    .X(_03439_));
 sg13g2_nand2_1 _21102_ (.Y(_03440_),
    .A(net1058),
    .B(_03424_));
 sg13g2_o21ai_1 _21103_ (.B1(_03440_),
    .Y(_01398_),
    .A1(net184),
    .A2(_03438_));
 sg13g2_buf_1 _21104_ (.A(_03042_),
    .X(_03441_));
 sg13g2_buf_1 _21105_ (.A(_03441_),
    .X(_03442_));
 sg13g2_nand2_1 _21106_ (.Y(_03443_),
    .A(net662),
    .B(\mem.mem_internal.code_mem[244][5] ));
 sg13g2_buf_1 _21107_ (.A(_12657_),
    .X(_03444_));
 sg13g2_nand2_1 _21108_ (.Y(_03445_),
    .A(net1057),
    .B(_03424_));
 sg13g2_o21ai_1 _21109_ (.B1(_03445_),
    .Y(_01399_),
    .A1(_03425_),
    .A2(_03443_));
 sg13g2_nand2_1 _21110_ (.Y(_03446_),
    .A(net662),
    .B(\mem.mem_internal.code_mem[244][6] ));
 sg13g2_buf_1 _21111_ (.A(_12661_),
    .X(_03447_));
 sg13g2_nand2_1 _21112_ (.Y(_03448_),
    .A(net1056),
    .B(_03424_));
 sg13g2_o21ai_1 _21113_ (.B1(_03448_),
    .Y(_01400_),
    .A1(_03425_),
    .A2(_03446_));
 sg13g2_nand2_1 _21114_ (.Y(_03449_),
    .A(net662),
    .B(\mem.mem_internal.code_mem[244][7] ));
 sg13g2_buf_1 _21115_ (.A(_12665_),
    .X(_03450_));
 sg13g2_nand2_1 _21116_ (.Y(_03451_),
    .A(net1055),
    .B(_03424_));
 sg13g2_o21ai_1 _21117_ (.B1(_03451_),
    .Y(_01401_),
    .A1(net184),
    .A2(_03449_));
 sg13g2_nor2_1 _21118_ (.A(net555),
    .B(net459),
    .Y(_03452_));
 sg13g2_buf_2 _21119_ (.A(_03452_),
    .X(_03453_));
 sg13g2_buf_1 _21120_ (.A(_03453_),
    .X(_03454_));
 sg13g2_nand2_1 _21121_ (.Y(_03455_),
    .A(net662),
    .B(\mem.mem_internal.code_mem[245][0] ));
 sg13g2_nand2_1 _21122_ (.Y(_03456_),
    .A(net1062),
    .B(net183));
 sg13g2_o21ai_1 _21123_ (.B1(_03456_),
    .Y(_01402_),
    .A1(net183),
    .A2(_03455_));
 sg13g2_nand2_1 _21124_ (.Y(_03457_),
    .A(net662),
    .B(\mem.mem_internal.code_mem[245][1] ));
 sg13g2_nand2_1 _21125_ (.Y(_03458_),
    .A(net1061),
    .B(net183));
 sg13g2_o21ai_1 _21126_ (.B1(_03458_),
    .Y(_01403_),
    .A1(net183),
    .A2(_03457_));
 sg13g2_nand2_1 _21127_ (.Y(_03459_),
    .A(_03442_),
    .B(\mem.mem_internal.code_mem[245][2] ));
 sg13g2_nand2_1 _21128_ (.Y(_03460_),
    .A(net1060),
    .B(_03453_));
 sg13g2_o21ai_1 _21129_ (.B1(_03460_),
    .Y(_01404_),
    .A1(_03454_),
    .A2(_03459_));
 sg13g2_nand2_1 _21130_ (.Y(_03461_),
    .A(_03442_),
    .B(\mem.mem_internal.code_mem[245][3] ));
 sg13g2_nand2_1 _21131_ (.Y(_03462_),
    .A(net1059),
    .B(_03453_));
 sg13g2_o21ai_1 _21132_ (.B1(_03462_),
    .Y(_01405_),
    .A1(net183),
    .A2(_03461_));
 sg13g2_nand2_1 _21133_ (.Y(_03463_),
    .A(net662),
    .B(\mem.mem_internal.code_mem[245][4] ));
 sg13g2_nand2_1 _21134_ (.Y(_03464_),
    .A(net1058),
    .B(_03453_));
 sg13g2_o21ai_1 _21135_ (.B1(_03464_),
    .Y(_01406_),
    .A1(net183),
    .A2(_03463_));
 sg13g2_nand2_1 _21136_ (.Y(_03465_),
    .A(net662),
    .B(\mem.mem_internal.code_mem[245][5] ));
 sg13g2_nand2_1 _21137_ (.Y(_03466_),
    .A(net1057),
    .B(_03453_));
 sg13g2_o21ai_1 _21138_ (.B1(_03466_),
    .Y(_01407_),
    .A1(_03454_),
    .A2(_03465_));
 sg13g2_nand2_1 _21139_ (.Y(_03467_),
    .A(net662),
    .B(\mem.mem_internal.code_mem[245][6] ));
 sg13g2_nand2_1 _21140_ (.Y(_03468_),
    .A(net1056),
    .B(_03453_));
 sg13g2_o21ai_1 _21141_ (.B1(_03468_),
    .Y(_01408_),
    .A1(net183),
    .A2(_03467_));
 sg13g2_buf_1 _21142_ (.A(_03441_),
    .X(_03469_));
 sg13g2_nand2_1 _21143_ (.Y(_03470_),
    .A(net661),
    .B(\mem.mem_internal.code_mem[245][7] ));
 sg13g2_nand2_1 _21144_ (.Y(_03471_),
    .A(net1055),
    .B(_03453_));
 sg13g2_o21ai_1 _21145_ (.B1(_03471_),
    .Y(_01409_),
    .A1(net183),
    .A2(_03470_));
 sg13g2_nor2_1 _21146_ (.A(_10350_),
    .B(net459),
    .Y(_03472_));
 sg13g2_buf_2 _21147_ (.A(_03472_),
    .X(_03473_));
 sg13g2_buf_1 _21148_ (.A(_03473_),
    .X(_03474_));
 sg13g2_nand2_1 _21149_ (.Y(_03475_),
    .A(net661),
    .B(\mem.mem_internal.code_mem[246][0] ));
 sg13g2_nand2_1 _21150_ (.Y(_03476_),
    .A(net1062),
    .B(net182));
 sg13g2_o21ai_1 _21151_ (.B1(_03476_),
    .Y(_01410_),
    .A1(net182),
    .A2(_03475_));
 sg13g2_nand2_1 _21152_ (.Y(_03477_),
    .A(net661),
    .B(\mem.mem_internal.code_mem[246][1] ));
 sg13g2_nand2_1 _21153_ (.Y(_03478_),
    .A(net1061),
    .B(net182));
 sg13g2_o21ai_1 _21154_ (.B1(_03478_),
    .Y(_01411_),
    .A1(net182),
    .A2(_03477_));
 sg13g2_nand2_1 _21155_ (.Y(_03479_),
    .A(net661),
    .B(\mem.mem_internal.code_mem[246][2] ));
 sg13g2_nand2_1 _21156_ (.Y(_03480_),
    .A(_03433_),
    .B(_03473_));
 sg13g2_o21ai_1 _21157_ (.B1(_03480_),
    .Y(_01412_),
    .A1(net182),
    .A2(_03479_));
 sg13g2_nand2_1 _21158_ (.Y(_03481_),
    .A(net661),
    .B(\mem.mem_internal.code_mem[246][3] ));
 sg13g2_nand2_1 _21159_ (.Y(_03482_),
    .A(_03436_),
    .B(_03473_));
 sg13g2_o21ai_1 _21160_ (.B1(_03482_),
    .Y(_01413_),
    .A1(net182),
    .A2(_03481_));
 sg13g2_nand2_1 _21161_ (.Y(_03483_),
    .A(net661),
    .B(\mem.mem_internal.code_mem[246][4] ));
 sg13g2_nand2_1 _21162_ (.Y(_03484_),
    .A(_03439_),
    .B(_03473_));
 sg13g2_o21ai_1 _21163_ (.B1(_03484_),
    .Y(_01414_),
    .A1(net182),
    .A2(_03483_));
 sg13g2_nand2_1 _21164_ (.Y(_03485_),
    .A(_03469_),
    .B(\mem.mem_internal.code_mem[246][5] ));
 sg13g2_nand2_1 _21165_ (.Y(_03486_),
    .A(_03444_),
    .B(_03473_));
 sg13g2_o21ai_1 _21166_ (.B1(_03486_),
    .Y(_01415_),
    .A1(_03474_),
    .A2(_03485_));
 sg13g2_nand2_1 _21167_ (.Y(_03487_),
    .A(_03469_),
    .B(\mem.mem_internal.code_mem[246][6] ));
 sg13g2_nand2_1 _21168_ (.Y(_03488_),
    .A(_03447_),
    .B(_03473_));
 sg13g2_o21ai_1 _21169_ (.B1(_03488_),
    .Y(_01416_),
    .A1(_03474_),
    .A2(_03487_));
 sg13g2_nand2_1 _21170_ (.Y(_03489_),
    .A(net661),
    .B(\mem.mem_internal.code_mem[246][7] ));
 sg13g2_nand2_1 _21171_ (.Y(_03490_),
    .A(_03450_),
    .B(_03473_));
 sg13g2_o21ai_1 _21172_ (.B1(_03490_),
    .Y(_01417_),
    .A1(net182),
    .A2(_03489_));
 sg13g2_nor2_1 _21173_ (.A(net553),
    .B(net459),
    .Y(_03491_));
 sg13g2_buf_2 _21174_ (.A(_03491_),
    .X(_03492_));
 sg13g2_buf_1 _21175_ (.A(_03492_),
    .X(_03493_));
 sg13g2_nand2_1 _21176_ (.Y(_03494_),
    .A(net661),
    .B(\mem.mem_internal.code_mem[247][0] ));
 sg13g2_nand2_1 _21177_ (.Y(_03495_),
    .A(net1062),
    .B(net181));
 sg13g2_o21ai_1 _21178_ (.B1(_03495_),
    .Y(_01418_),
    .A1(net181),
    .A2(_03494_));
 sg13g2_buf_1 _21179_ (.A(_03441_),
    .X(_03496_));
 sg13g2_nand2_1 _21180_ (.Y(_03497_),
    .A(net660),
    .B(\mem.mem_internal.code_mem[247][1] ));
 sg13g2_nand2_1 _21181_ (.Y(_03498_),
    .A(net1061),
    .B(net181));
 sg13g2_o21ai_1 _21182_ (.B1(_03498_),
    .Y(_01419_),
    .A1(net181),
    .A2(_03497_));
 sg13g2_nand2_1 _21183_ (.Y(_03499_),
    .A(net660),
    .B(\mem.mem_internal.code_mem[247][2] ));
 sg13g2_nand2_1 _21184_ (.Y(_03500_),
    .A(_03433_),
    .B(_03492_));
 sg13g2_o21ai_1 _21185_ (.B1(_03500_),
    .Y(_01420_),
    .A1(_03493_),
    .A2(_03499_));
 sg13g2_nand2_1 _21186_ (.Y(_03501_),
    .A(net660),
    .B(\mem.mem_internal.code_mem[247][3] ));
 sg13g2_nand2_1 _21187_ (.Y(_03502_),
    .A(_03436_),
    .B(_03492_));
 sg13g2_o21ai_1 _21188_ (.B1(_03502_),
    .Y(_01421_),
    .A1(net181),
    .A2(_03501_));
 sg13g2_nand2_1 _21189_ (.Y(_03503_),
    .A(net660),
    .B(\mem.mem_internal.code_mem[247][4] ));
 sg13g2_nand2_1 _21190_ (.Y(_03504_),
    .A(_03439_),
    .B(_03492_));
 sg13g2_o21ai_1 _21191_ (.B1(_03504_),
    .Y(_01422_),
    .A1(net181),
    .A2(_03503_));
 sg13g2_nand2_1 _21192_ (.Y(_03505_),
    .A(net660),
    .B(\mem.mem_internal.code_mem[247][5] ));
 sg13g2_nand2_1 _21193_ (.Y(_03506_),
    .A(_03444_),
    .B(_03492_));
 sg13g2_o21ai_1 _21194_ (.B1(_03506_),
    .Y(_01423_),
    .A1(_03493_),
    .A2(_03505_));
 sg13g2_nand2_1 _21195_ (.Y(_03507_),
    .A(_03496_),
    .B(\mem.mem_internal.code_mem[247][6] ));
 sg13g2_nand2_1 _21196_ (.Y(_03508_),
    .A(_03447_),
    .B(_03492_));
 sg13g2_o21ai_1 _21197_ (.B1(_03508_),
    .Y(_01424_),
    .A1(net181),
    .A2(_03507_));
 sg13g2_nand2_1 _21198_ (.Y(_03509_),
    .A(_03496_),
    .B(\mem.mem_internal.code_mem[247][7] ));
 sg13g2_nand2_1 _21199_ (.Y(_03510_),
    .A(_03450_),
    .B(_03492_));
 sg13g2_o21ai_1 _21200_ (.B1(_03510_),
    .Y(_01425_),
    .A1(net181),
    .A2(_03509_));
 sg13g2_nor2_1 _21201_ (.A(net552),
    .B(net459),
    .Y(_03511_));
 sg13g2_buf_2 _21202_ (.A(_03511_),
    .X(_03512_));
 sg13g2_buf_1 _21203_ (.A(_03512_),
    .X(_03513_));
 sg13g2_nand2_1 _21204_ (.Y(_03514_),
    .A(net660),
    .B(\mem.mem_internal.code_mem[248][0] ));
 sg13g2_nand2_1 _21205_ (.Y(_03515_),
    .A(net1062),
    .B(net180));
 sg13g2_o21ai_1 _21206_ (.B1(_03515_),
    .Y(_01426_),
    .A1(net180),
    .A2(_03514_));
 sg13g2_nand2_1 _21207_ (.Y(_03516_),
    .A(net660),
    .B(\mem.mem_internal.code_mem[248][1] ));
 sg13g2_nand2_1 _21208_ (.Y(_03517_),
    .A(_03430_),
    .B(net180));
 sg13g2_o21ai_1 _21209_ (.B1(_03517_),
    .Y(_01427_),
    .A1(net180),
    .A2(_03516_));
 sg13g2_nand2_1 _21210_ (.Y(_03518_),
    .A(net660),
    .B(\mem.mem_internal.code_mem[248][2] ));
 sg13g2_nand2_1 _21211_ (.Y(_03519_),
    .A(net1060),
    .B(_03512_));
 sg13g2_o21ai_1 _21212_ (.B1(_03519_),
    .Y(_01428_),
    .A1(_03513_),
    .A2(_03518_));
 sg13g2_buf_1 _21213_ (.A(_03441_),
    .X(_03520_));
 sg13g2_nand2_1 _21214_ (.Y(_03521_),
    .A(net659),
    .B(\mem.mem_internal.code_mem[248][3] ));
 sg13g2_nand2_1 _21215_ (.Y(_03522_),
    .A(net1059),
    .B(_03512_));
 sg13g2_o21ai_1 _21216_ (.B1(_03522_),
    .Y(_01429_),
    .A1(net180),
    .A2(_03521_));
 sg13g2_nand2_1 _21217_ (.Y(_03523_),
    .A(_03520_),
    .B(\mem.mem_internal.code_mem[248][4] ));
 sg13g2_nand2_1 _21218_ (.Y(_03524_),
    .A(net1058),
    .B(_03512_));
 sg13g2_o21ai_1 _21219_ (.B1(_03524_),
    .Y(_01430_),
    .A1(_03513_),
    .A2(_03523_));
 sg13g2_nand2_1 _21220_ (.Y(_03525_),
    .A(net659),
    .B(\mem.mem_internal.code_mem[248][5] ));
 sg13g2_nand2_1 _21221_ (.Y(_03526_),
    .A(net1057),
    .B(_03512_));
 sg13g2_o21ai_1 _21222_ (.B1(_03526_),
    .Y(_01431_),
    .A1(net180),
    .A2(_03525_));
 sg13g2_nand2_1 _21223_ (.Y(_03527_),
    .A(net659),
    .B(\mem.mem_internal.code_mem[248][6] ));
 sg13g2_nand2_1 _21224_ (.Y(_03528_),
    .A(net1056),
    .B(_03512_));
 sg13g2_o21ai_1 _21225_ (.B1(_03528_),
    .Y(_01432_),
    .A1(net180),
    .A2(_03527_));
 sg13g2_nand2_1 _21226_ (.Y(_03529_),
    .A(net659),
    .B(\mem.mem_internal.code_mem[248][7] ));
 sg13g2_nand2_1 _21227_ (.Y(_03530_),
    .A(net1055),
    .B(_03512_));
 sg13g2_o21ai_1 _21228_ (.B1(_03530_),
    .Y(_01433_),
    .A1(net180),
    .A2(_03529_));
 sg13g2_nor2_1 _21229_ (.A(net551),
    .B(net459),
    .Y(_03531_));
 sg13g2_buf_2 _21230_ (.A(_03531_),
    .X(_03532_));
 sg13g2_buf_1 _21231_ (.A(_03532_),
    .X(_03533_));
 sg13g2_nand2_1 _21232_ (.Y(_03534_),
    .A(net659),
    .B(\mem.mem_internal.code_mem[249][0] ));
 sg13g2_nand2_1 _21233_ (.Y(_03535_),
    .A(_03427_),
    .B(_03533_));
 sg13g2_o21ai_1 _21234_ (.B1(_03535_),
    .Y(_01434_),
    .A1(net179),
    .A2(_03534_));
 sg13g2_nand2_1 _21235_ (.Y(_03536_),
    .A(net659),
    .B(\mem.mem_internal.code_mem[249][1] ));
 sg13g2_nand2_1 _21236_ (.Y(_03537_),
    .A(_03430_),
    .B(net179));
 sg13g2_o21ai_1 _21237_ (.B1(_03537_),
    .Y(_01435_),
    .A1(net179),
    .A2(_03536_));
 sg13g2_nand2_1 _21238_ (.Y(_03538_),
    .A(net659),
    .B(\mem.mem_internal.code_mem[249][2] ));
 sg13g2_nand2_1 _21239_ (.Y(_03539_),
    .A(net1060),
    .B(_03532_));
 sg13g2_o21ai_1 _21240_ (.B1(_03539_),
    .Y(_01436_),
    .A1(_03533_),
    .A2(_03538_));
 sg13g2_nand2_1 _21241_ (.Y(_03540_),
    .A(net659),
    .B(\mem.mem_internal.code_mem[249][3] ));
 sg13g2_nand2_1 _21242_ (.Y(_03541_),
    .A(net1059),
    .B(_03532_));
 sg13g2_o21ai_1 _21243_ (.B1(_03541_),
    .Y(_01437_),
    .A1(net179),
    .A2(_03540_));
 sg13g2_nand2_1 _21244_ (.Y(_03542_),
    .A(_03520_),
    .B(\mem.mem_internal.code_mem[249][4] ));
 sg13g2_nand2_1 _21245_ (.Y(_03543_),
    .A(net1058),
    .B(_03532_));
 sg13g2_o21ai_1 _21246_ (.B1(_03543_),
    .Y(_01438_),
    .A1(net179),
    .A2(_03542_));
 sg13g2_buf_1 _21247_ (.A(_03441_),
    .X(_03544_));
 sg13g2_nand2_1 _21248_ (.Y(_03545_),
    .A(net658),
    .B(\mem.mem_internal.code_mem[249][5] ));
 sg13g2_nand2_1 _21249_ (.Y(_03546_),
    .A(net1057),
    .B(_03532_));
 sg13g2_o21ai_1 _21250_ (.B1(_03546_),
    .Y(_01439_),
    .A1(net179),
    .A2(_03545_));
 sg13g2_nand2_1 _21251_ (.Y(_03547_),
    .A(net658),
    .B(\mem.mem_internal.code_mem[249][6] ));
 sg13g2_nand2_1 _21252_ (.Y(_03548_),
    .A(net1056),
    .B(_03532_));
 sg13g2_o21ai_1 _21253_ (.B1(_03548_),
    .Y(_01440_),
    .A1(net179),
    .A2(_03547_));
 sg13g2_nand2_1 _21254_ (.Y(_03549_),
    .A(net658),
    .B(\mem.mem_internal.code_mem[249][7] ));
 sg13g2_nand2_1 _21255_ (.Y(_03550_),
    .A(net1055),
    .B(_03532_));
 sg13g2_o21ai_1 _21256_ (.B1(_03550_),
    .Y(_01441_),
    .A1(net179),
    .A2(_03549_));
 sg13g2_nand2_1 _21257_ (.Y(_03551_),
    .A(_03240_),
    .B(\mem.mem_internal.code_mem[24][0] ));
 sg13g2_nor2_1 _21258_ (.A(_10397_),
    .B(_11947_),
    .Y(_03552_));
 sg13g2_buf_2 _21259_ (.A(_03552_),
    .X(_03553_));
 sg13g2_buf_1 _21260_ (.A(_03553_),
    .X(_03554_));
 sg13g2_nand2_1 _21261_ (.Y(_03555_),
    .A(_03427_),
    .B(net178));
 sg13g2_o21ai_1 _21262_ (.B1(_03555_),
    .Y(_01442_),
    .A1(_03551_),
    .A2(net178));
 sg13g2_nand2_1 _21263_ (.Y(_03556_),
    .A(net658),
    .B(\mem.mem_internal.code_mem[24][1] ));
 sg13g2_nand2_1 _21264_ (.Y(_03557_),
    .A(net1061),
    .B(net178));
 sg13g2_o21ai_1 _21265_ (.B1(_03557_),
    .Y(_01443_),
    .A1(net178),
    .A2(_03556_));
 sg13g2_nand2_1 _21266_ (.Y(_03558_),
    .A(net658),
    .B(\mem.mem_internal.code_mem[24][2] ));
 sg13g2_nand2_1 _21267_ (.Y(_03559_),
    .A(net1060),
    .B(_03553_));
 sg13g2_o21ai_1 _21268_ (.B1(_03559_),
    .Y(_01444_),
    .A1(net178),
    .A2(_03558_));
 sg13g2_nand2_1 _21269_ (.Y(_03560_),
    .A(net658),
    .B(\mem.mem_internal.code_mem[24][3] ));
 sg13g2_nand2_1 _21270_ (.Y(_03561_),
    .A(net1059),
    .B(_03553_));
 sg13g2_o21ai_1 _21271_ (.B1(_03561_),
    .Y(_01445_),
    .A1(net178),
    .A2(_03560_));
 sg13g2_nand2_1 _21272_ (.Y(_03562_),
    .A(net658),
    .B(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_nand2_1 _21273_ (.Y(_03563_),
    .A(net1058),
    .B(_03553_));
 sg13g2_o21ai_1 _21274_ (.B1(_03563_),
    .Y(_01446_),
    .A1(_03554_),
    .A2(_03562_));
 sg13g2_nand2_1 _21275_ (.Y(_03564_),
    .A(net658),
    .B(\mem.mem_internal.code_mem[24][5] ));
 sg13g2_nand2_1 _21276_ (.Y(_03565_),
    .A(net1057),
    .B(_03553_));
 sg13g2_o21ai_1 _21277_ (.B1(_03565_),
    .Y(_01447_),
    .A1(net178),
    .A2(_03564_));
 sg13g2_nand2_1 _21278_ (.Y(_03566_),
    .A(_03544_),
    .B(\mem.mem_internal.code_mem[24][6] ));
 sg13g2_nand2_1 _21279_ (.Y(_03567_),
    .A(net1056),
    .B(_03553_));
 sg13g2_o21ai_1 _21280_ (.B1(_03567_),
    .Y(_01448_),
    .A1(_03554_),
    .A2(_03566_));
 sg13g2_nand2_1 _21281_ (.Y(_03568_),
    .A(_03544_),
    .B(\mem.mem_internal.code_mem[24][7] ));
 sg13g2_nand2_1 _21282_ (.Y(_03569_),
    .A(net1055),
    .B(_03553_));
 sg13g2_o21ai_1 _21283_ (.B1(_03569_),
    .Y(_01449_),
    .A1(net178),
    .A2(_03568_));
 sg13g2_nor2_1 _21284_ (.A(_10445_),
    .B(_03342_),
    .Y(_03570_));
 sg13g2_buf_2 _21285_ (.A(_03570_),
    .X(_03571_));
 sg13g2_buf_1 _21286_ (.A(_03571_),
    .X(_03572_));
 sg13g2_buf_1 _21287_ (.A(_03441_),
    .X(_03573_));
 sg13g2_nand2_1 _21288_ (.Y(_03574_),
    .A(net657),
    .B(\mem.mem_internal.code_mem[250][0] ));
 sg13g2_nand2_1 _21289_ (.Y(_03575_),
    .A(net1062),
    .B(net348));
 sg13g2_o21ai_1 _21290_ (.B1(_03575_),
    .Y(_01450_),
    .A1(net348),
    .A2(_03574_));
 sg13g2_nand2_1 _21291_ (.Y(_03576_),
    .A(net657),
    .B(\mem.mem_internal.code_mem[250][1] ));
 sg13g2_nand2_1 _21292_ (.Y(_03577_),
    .A(net1061),
    .B(net348));
 sg13g2_o21ai_1 _21293_ (.B1(_03577_),
    .Y(_01451_),
    .A1(net348),
    .A2(_03576_));
 sg13g2_nand2_1 _21294_ (.Y(_03578_),
    .A(net657),
    .B(\mem.mem_internal.code_mem[250][2] ));
 sg13g2_nand2_1 _21295_ (.Y(_03579_),
    .A(net1060),
    .B(_03571_));
 sg13g2_o21ai_1 _21296_ (.B1(_03579_),
    .Y(_01452_),
    .A1(_03572_),
    .A2(_03578_));
 sg13g2_nand2_1 _21297_ (.Y(_03580_),
    .A(net657),
    .B(\mem.mem_internal.code_mem[250][3] ));
 sg13g2_nand2_1 _21298_ (.Y(_03581_),
    .A(net1059),
    .B(_03571_));
 sg13g2_o21ai_1 _21299_ (.B1(_03581_),
    .Y(_01453_),
    .A1(net348),
    .A2(_03580_));
 sg13g2_nand2_1 _21300_ (.Y(_03582_),
    .A(_03573_),
    .B(\mem.mem_internal.code_mem[250][4] ));
 sg13g2_nand2_1 _21301_ (.Y(_03583_),
    .A(net1058),
    .B(_03571_));
 sg13g2_o21ai_1 _21302_ (.B1(_03583_),
    .Y(_01454_),
    .A1(_03572_),
    .A2(_03582_));
 sg13g2_nand2_1 _21303_ (.Y(_03584_),
    .A(net657),
    .B(\mem.mem_internal.code_mem[250][5] ));
 sg13g2_nand2_1 _21304_ (.Y(_03585_),
    .A(net1057),
    .B(_03571_));
 sg13g2_o21ai_1 _21305_ (.B1(_03585_),
    .Y(_01455_),
    .A1(net348),
    .A2(_03584_));
 sg13g2_nand2_1 _21306_ (.Y(_03586_),
    .A(net657),
    .B(\mem.mem_internal.code_mem[250][6] ));
 sg13g2_nand2_1 _21307_ (.Y(_03587_),
    .A(net1056),
    .B(_03571_));
 sg13g2_o21ai_1 _21308_ (.B1(_03587_),
    .Y(_01456_),
    .A1(net348),
    .A2(_03586_));
 sg13g2_nand2_1 _21309_ (.Y(_03588_),
    .A(net657),
    .B(\mem.mem_internal.code_mem[250][7] ));
 sg13g2_nand2_1 _21310_ (.Y(_03589_),
    .A(net1055),
    .B(_03571_));
 sg13g2_o21ai_1 _21311_ (.B1(_03589_),
    .Y(_01457_),
    .A1(net348),
    .A2(_03588_));
 sg13g2_nor2_1 _21312_ (.A(_10468_),
    .B(_03342_),
    .Y(_03590_));
 sg13g2_buf_2 _21313_ (.A(_03590_),
    .X(_03591_));
 sg13g2_buf_1 _21314_ (.A(_03591_),
    .X(_03592_));
 sg13g2_nand2_1 _21315_ (.Y(_03593_),
    .A(net657),
    .B(\mem.mem_internal.code_mem[251][0] ));
 sg13g2_nand2_1 _21316_ (.Y(_03594_),
    .A(net1062),
    .B(_03592_));
 sg13g2_o21ai_1 _21317_ (.B1(_03594_),
    .Y(_01458_),
    .A1(net347),
    .A2(_03593_));
 sg13g2_nand2_1 _21318_ (.Y(_03595_),
    .A(_03573_),
    .B(\mem.mem_internal.code_mem[251][1] ));
 sg13g2_nand2_1 _21319_ (.Y(_03596_),
    .A(net1061),
    .B(net347));
 sg13g2_o21ai_1 _21320_ (.B1(_03596_),
    .Y(_01459_),
    .A1(net347),
    .A2(_03595_));
 sg13g2_buf_1 _21321_ (.A(_03441_),
    .X(_03597_));
 sg13g2_nand2_1 _21322_ (.Y(_03598_),
    .A(net656),
    .B(\mem.mem_internal.code_mem[251][2] ));
 sg13g2_nand2_1 _21323_ (.Y(_03599_),
    .A(net1060),
    .B(_03591_));
 sg13g2_o21ai_1 _21324_ (.B1(_03599_),
    .Y(_01460_),
    .A1(_03592_),
    .A2(_03598_));
 sg13g2_nand2_1 _21325_ (.Y(_03600_),
    .A(net656),
    .B(\mem.mem_internal.code_mem[251][3] ));
 sg13g2_nand2_1 _21326_ (.Y(_03601_),
    .A(net1059),
    .B(_03591_));
 sg13g2_o21ai_1 _21327_ (.B1(_03601_),
    .Y(_01461_),
    .A1(net347),
    .A2(_03600_));
 sg13g2_nand2_1 _21328_ (.Y(_03602_),
    .A(net656),
    .B(\mem.mem_internal.code_mem[251][4] ));
 sg13g2_nand2_1 _21329_ (.Y(_03603_),
    .A(net1058),
    .B(_03591_));
 sg13g2_o21ai_1 _21330_ (.B1(_03603_),
    .Y(_01462_),
    .A1(net347),
    .A2(_03602_));
 sg13g2_nand2_1 _21331_ (.Y(_03604_),
    .A(net656),
    .B(\mem.mem_internal.code_mem[251][5] ));
 sg13g2_nand2_1 _21332_ (.Y(_03605_),
    .A(net1057),
    .B(_03591_));
 sg13g2_o21ai_1 _21333_ (.B1(_03605_),
    .Y(_01463_),
    .A1(net347),
    .A2(_03604_));
 sg13g2_nand2_1 _21334_ (.Y(_03606_),
    .A(net656),
    .B(\mem.mem_internal.code_mem[251][6] ));
 sg13g2_nand2_1 _21335_ (.Y(_03607_),
    .A(net1056),
    .B(_03591_));
 sg13g2_o21ai_1 _21336_ (.B1(_03607_),
    .Y(_01464_),
    .A1(net347),
    .A2(_03606_));
 sg13g2_nand2_1 _21337_ (.Y(_03608_),
    .A(net656),
    .B(\mem.mem_internal.code_mem[251][7] ));
 sg13g2_nand2_1 _21338_ (.Y(_03609_),
    .A(net1055),
    .B(_03591_));
 sg13g2_o21ai_1 _21339_ (.B1(_03609_),
    .Y(_01465_),
    .A1(net347),
    .A2(_03608_));
 sg13g2_nor2_1 _21340_ (.A(net773),
    .B(_03342_),
    .Y(_03610_));
 sg13g2_buf_2 _21341_ (.A(_03610_),
    .X(_03611_));
 sg13g2_buf_1 _21342_ (.A(_03611_),
    .X(_03612_));
 sg13g2_nand2_1 _21343_ (.Y(_03613_),
    .A(net656),
    .B(\mem.mem_internal.code_mem[252][0] ));
 sg13g2_nand2_1 _21344_ (.Y(_03614_),
    .A(net1062),
    .B(net346));
 sg13g2_o21ai_1 _21345_ (.B1(_03614_),
    .Y(_01466_),
    .A1(_03612_),
    .A2(_03613_));
 sg13g2_nand2_1 _21346_ (.Y(_03615_),
    .A(_03597_),
    .B(\mem.mem_internal.code_mem[252][1] ));
 sg13g2_nand2_1 _21347_ (.Y(_03616_),
    .A(net1061),
    .B(_03612_));
 sg13g2_o21ai_1 _21348_ (.B1(_03616_),
    .Y(_01467_),
    .A1(net346),
    .A2(_03615_));
 sg13g2_nand2_1 _21349_ (.Y(_03617_),
    .A(_03597_),
    .B(\mem.mem_internal.code_mem[252][2] ));
 sg13g2_nand2_1 _21350_ (.Y(_03618_),
    .A(net1060),
    .B(_03611_));
 sg13g2_o21ai_1 _21351_ (.B1(_03618_),
    .Y(_01468_),
    .A1(net346),
    .A2(_03617_));
 sg13g2_nand2_1 _21352_ (.Y(_03619_),
    .A(net656),
    .B(\mem.mem_internal.code_mem[252][3] ));
 sg13g2_nand2_1 _21353_ (.Y(_03620_),
    .A(net1059),
    .B(_03611_));
 sg13g2_o21ai_1 _21354_ (.B1(_03620_),
    .Y(_01469_),
    .A1(net346),
    .A2(_03619_));
 sg13g2_buf_2 _21355_ (.A(_03042_),
    .X(_03621_));
 sg13g2_buf_1 _21356_ (.A(_03621_),
    .X(_03622_));
 sg13g2_nand2_1 _21357_ (.Y(_03623_),
    .A(net655),
    .B(\mem.mem_internal.code_mem[252][4] ));
 sg13g2_nand2_1 _21358_ (.Y(_03624_),
    .A(net1058),
    .B(_03611_));
 sg13g2_o21ai_1 _21359_ (.B1(_03624_),
    .Y(_01470_),
    .A1(net346),
    .A2(_03623_));
 sg13g2_nand2_1 _21360_ (.Y(_03625_),
    .A(net655),
    .B(\mem.mem_internal.code_mem[252][5] ));
 sg13g2_nand2_1 _21361_ (.Y(_03626_),
    .A(net1057),
    .B(_03611_));
 sg13g2_o21ai_1 _21362_ (.B1(_03626_),
    .Y(_01471_),
    .A1(net346),
    .A2(_03625_));
 sg13g2_nand2_1 _21363_ (.Y(_03627_),
    .A(net655),
    .B(\mem.mem_internal.code_mem[252][6] ));
 sg13g2_nand2_1 _21364_ (.Y(_03628_),
    .A(net1056),
    .B(_03611_));
 sg13g2_o21ai_1 _21365_ (.B1(_03628_),
    .Y(_01472_),
    .A1(net346),
    .A2(_03627_));
 sg13g2_nand2_1 _21366_ (.Y(_03629_),
    .A(net655),
    .B(\mem.mem_internal.code_mem[252][7] ));
 sg13g2_nand2_1 _21367_ (.Y(_03630_),
    .A(net1055),
    .B(_03611_));
 sg13g2_o21ai_1 _21368_ (.B1(_03630_),
    .Y(_01473_),
    .A1(net346),
    .A2(_03629_));
 sg13g2_nor2_1 _21369_ (.A(_10514_),
    .B(_03342_),
    .Y(_03631_));
 sg13g2_buf_2 _21370_ (.A(_03631_),
    .X(_03632_));
 sg13g2_buf_1 _21371_ (.A(_03632_),
    .X(_03633_));
 sg13g2_nand2_1 _21372_ (.Y(_03634_),
    .A(_03622_),
    .B(\mem.mem_internal.code_mem[253][0] ));
 sg13g2_buf_1 _21373_ (.A(_12637_),
    .X(_03635_));
 sg13g2_nand2_1 _21374_ (.Y(_03636_),
    .A(net1054),
    .B(net345));
 sg13g2_o21ai_1 _21375_ (.B1(_03636_),
    .Y(_01474_),
    .A1(net345),
    .A2(_03634_));
 sg13g2_nand2_1 _21376_ (.Y(_03637_),
    .A(net655),
    .B(\mem.mem_internal.code_mem[253][1] ));
 sg13g2_buf_1 _21377_ (.A(_12641_),
    .X(_03638_));
 sg13g2_nand2_1 _21378_ (.Y(_03639_),
    .A(net1053),
    .B(_03633_));
 sg13g2_o21ai_1 _21379_ (.B1(_03639_),
    .Y(_01475_),
    .A1(_03633_),
    .A2(_03637_));
 sg13g2_nand2_1 _21380_ (.Y(_03640_),
    .A(net655),
    .B(\mem.mem_internal.code_mem[253][2] ));
 sg13g2_buf_1 _21381_ (.A(_12645_),
    .X(_03641_));
 sg13g2_nand2_1 _21382_ (.Y(_03642_),
    .A(net1052),
    .B(_03632_));
 sg13g2_o21ai_1 _21383_ (.B1(_03642_),
    .Y(_01476_),
    .A1(net345),
    .A2(_03640_));
 sg13g2_nand2_1 _21384_ (.Y(_03643_),
    .A(net655),
    .B(\mem.mem_internal.code_mem[253][3] ));
 sg13g2_buf_1 _21385_ (.A(_12649_),
    .X(_03644_));
 sg13g2_nand2_1 _21386_ (.Y(_03645_),
    .A(net1051),
    .B(_03632_));
 sg13g2_o21ai_1 _21387_ (.B1(_03645_),
    .Y(_01477_),
    .A1(net345),
    .A2(_03643_));
 sg13g2_nand2_1 _21388_ (.Y(_03646_),
    .A(_03622_),
    .B(\mem.mem_internal.code_mem[253][4] ));
 sg13g2_buf_1 _21389_ (.A(_12653_),
    .X(_03647_));
 sg13g2_nand2_1 _21390_ (.Y(_03648_),
    .A(net1050),
    .B(_03632_));
 sg13g2_o21ai_1 _21391_ (.B1(_03648_),
    .Y(_01478_),
    .A1(net345),
    .A2(_03646_));
 sg13g2_nand2_1 _21392_ (.Y(_03649_),
    .A(net655),
    .B(\mem.mem_internal.code_mem[253][5] ));
 sg13g2_buf_1 _21393_ (.A(_12657_),
    .X(_03650_));
 sg13g2_nand2_1 _21394_ (.Y(_03651_),
    .A(net1049),
    .B(_03632_));
 sg13g2_o21ai_1 _21395_ (.B1(_03651_),
    .Y(_01479_),
    .A1(net345),
    .A2(_03649_));
 sg13g2_buf_1 _21396_ (.A(_03621_),
    .X(_03652_));
 sg13g2_nand2_1 _21397_ (.Y(_03653_),
    .A(net654),
    .B(\mem.mem_internal.code_mem[253][6] ));
 sg13g2_buf_1 _21398_ (.A(_12661_),
    .X(_03654_));
 sg13g2_nand2_1 _21399_ (.Y(_03655_),
    .A(net1048),
    .B(_03632_));
 sg13g2_o21ai_1 _21400_ (.B1(_03655_),
    .Y(_01480_),
    .A1(net345),
    .A2(_03653_));
 sg13g2_nand2_1 _21401_ (.Y(_03656_),
    .A(net654),
    .B(\mem.mem_internal.code_mem[253][7] ));
 sg13g2_buf_1 _21402_ (.A(_12665_),
    .X(_03657_));
 sg13g2_nand2_1 _21403_ (.Y(_03658_),
    .A(net1047),
    .B(_03632_));
 sg13g2_o21ai_1 _21404_ (.B1(_03658_),
    .Y(_01481_),
    .A1(net345),
    .A2(_03656_));
 sg13g2_nor2_1 _21405_ (.A(_10565_),
    .B(_03342_),
    .Y(_03659_));
 sg13g2_buf_2 _21406_ (.A(_03659_),
    .X(_03660_));
 sg13g2_buf_1 _21407_ (.A(_03660_),
    .X(_03661_));
 sg13g2_nand2_1 _21408_ (.Y(_03662_),
    .A(_03652_),
    .B(\mem.mem_internal.code_mem[254][0] ));
 sg13g2_nand2_1 _21409_ (.Y(_03663_),
    .A(_03635_),
    .B(net344));
 sg13g2_o21ai_1 _21410_ (.B1(_03663_),
    .Y(_01482_),
    .A1(net344),
    .A2(_03662_));
 sg13g2_nand2_1 _21411_ (.Y(_03664_),
    .A(_03652_),
    .B(\mem.mem_internal.code_mem[254][1] ));
 sg13g2_nand2_1 _21412_ (.Y(_03665_),
    .A(_03638_),
    .B(_03661_));
 sg13g2_o21ai_1 _21413_ (.B1(_03665_),
    .Y(_01483_),
    .A1(_03661_),
    .A2(_03664_));
 sg13g2_nand2_1 _21414_ (.Y(_03666_),
    .A(net654),
    .B(\mem.mem_internal.code_mem[254][2] ));
 sg13g2_nand2_1 _21415_ (.Y(_03667_),
    .A(_03641_),
    .B(_03660_));
 sg13g2_o21ai_1 _21416_ (.B1(_03667_),
    .Y(_01484_),
    .A1(net344),
    .A2(_03666_));
 sg13g2_nand2_1 _21417_ (.Y(_03668_),
    .A(net654),
    .B(\mem.mem_internal.code_mem[254][3] ));
 sg13g2_nand2_1 _21418_ (.Y(_03669_),
    .A(_03644_),
    .B(_03660_));
 sg13g2_o21ai_1 _21419_ (.B1(_03669_),
    .Y(_01485_),
    .A1(net344),
    .A2(_03668_));
 sg13g2_nand2_1 _21420_ (.Y(_03670_),
    .A(net654),
    .B(\mem.mem_internal.code_mem[254][4] ));
 sg13g2_nand2_1 _21421_ (.Y(_03671_),
    .A(_03647_),
    .B(_03660_));
 sg13g2_o21ai_1 _21422_ (.B1(_03671_),
    .Y(_01486_),
    .A1(net344),
    .A2(_03670_));
 sg13g2_nand2_1 _21423_ (.Y(_03672_),
    .A(net654),
    .B(\mem.mem_internal.code_mem[254][5] ));
 sg13g2_nand2_1 _21424_ (.Y(_03673_),
    .A(_03650_),
    .B(_03660_));
 sg13g2_o21ai_1 _21425_ (.B1(_03673_),
    .Y(_01487_),
    .A1(net344),
    .A2(_03672_));
 sg13g2_nand2_1 _21426_ (.Y(_03674_),
    .A(net654),
    .B(\mem.mem_internal.code_mem[254][6] ));
 sg13g2_nand2_1 _21427_ (.Y(_03675_),
    .A(_03654_),
    .B(_03660_));
 sg13g2_o21ai_1 _21428_ (.B1(_03675_),
    .Y(_01488_),
    .A1(net344),
    .A2(_03674_));
 sg13g2_nand2_1 _21429_ (.Y(_03676_),
    .A(net654),
    .B(\mem.mem_internal.code_mem[254][7] ));
 sg13g2_nand2_1 _21430_ (.Y(_03677_),
    .A(_03657_),
    .B(_03660_));
 sg13g2_o21ai_1 _21431_ (.B1(_03677_),
    .Y(_01489_),
    .A1(net344),
    .A2(_03676_));
 sg13g2_nor2_1 _21432_ (.A(_10587_),
    .B(_03342_),
    .Y(_03678_));
 sg13g2_buf_2 _21433_ (.A(_03678_),
    .X(_03679_));
 sg13g2_buf_1 _21434_ (.A(_03679_),
    .X(_03680_));
 sg13g2_buf_1 _21435_ (.A(_03621_),
    .X(_03681_));
 sg13g2_nand2_1 _21436_ (.Y(_03682_),
    .A(net653),
    .B(\mem.mem_internal.code_mem[255][0] ));
 sg13g2_nand2_1 _21437_ (.Y(_03683_),
    .A(_03635_),
    .B(net343));
 sg13g2_o21ai_1 _21438_ (.B1(_03683_),
    .Y(_01490_),
    .A1(net343),
    .A2(_03682_));
 sg13g2_nand2_1 _21439_ (.Y(_03684_),
    .A(net653),
    .B(\mem.mem_internal.code_mem[255][1] ));
 sg13g2_nand2_1 _21440_ (.Y(_03685_),
    .A(_03638_),
    .B(_03680_));
 sg13g2_o21ai_1 _21441_ (.B1(_03685_),
    .Y(_01491_),
    .A1(_03680_),
    .A2(_03684_));
 sg13g2_nand2_1 _21442_ (.Y(_03686_),
    .A(net653),
    .B(\mem.mem_internal.code_mem[255][2] ));
 sg13g2_nand2_1 _21443_ (.Y(_03687_),
    .A(_03641_),
    .B(_03679_));
 sg13g2_o21ai_1 _21444_ (.B1(_03687_),
    .Y(_01492_),
    .A1(net343),
    .A2(_03686_));
 sg13g2_nand2_1 _21445_ (.Y(_03688_),
    .A(net653),
    .B(\mem.mem_internal.code_mem[255][3] ));
 sg13g2_nand2_1 _21446_ (.Y(_03689_),
    .A(_03644_),
    .B(_03679_));
 sg13g2_o21ai_1 _21447_ (.B1(_03689_),
    .Y(_01493_),
    .A1(net343),
    .A2(_03688_));
 sg13g2_nand2_1 _21448_ (.Y(_03690_),
    .A(net653),
    .B(\mem.mem_internal.code_mem[255][4] ));
 sg13g2_nand2_1 _21449_ (.Y(_03691_),
    .A(_03647_),
    .B(_03679_));
 sg13g2_o21ai_1 _21450_ (.B1(_03691_),
    .Y(_01494_),
    .A1(net343),
    .A2(_03690_));
 sg13g2_nand2_1 _21451_ (.Y(_03692_),
    .A(net653),
    .B(\mem.mem_internal.code_mem[255][5] ));
 sg13g2_nand2_1 _21452_ (.Y(_03693_),
    .A(_03650_),
    .B(_03679_));
 sg13g2_o21ai_1 _21453_ (.B1(_03693_),
    .Y(_01495_),
    .A1(net343),
    .A2(_03692_));
 sg13g2_nand2_1 _21454_ (.Y(_03694_),
    .A(_03681_),
    .B(\mem.mem_internal.code_mem[255][6] ));
 sg13g2_nand2_1 _21455_ (.Y(_03695_),
    .A(_03654_),
    .B(_03679_));
 sg13g2_o21ai_1 _21456_ (.B1(_03695_),
    .Y(_01496_),
    .A1(net343),
    .A2(_03694_));
 sg13g2_nand2_1 _21457_ (.Y(_03696_),
    .A(_03681_),
    .B(\mem.mem_internal.code_mem[255][7] ));
 sg13g2_nand2_1 _21458_ (.Y(_03697_),
    .A(_03657_),
    .B(_03679_));
 sg13g2_o21ai_1 _21459_ (.B1(_03697_),
    .Y(_01497_),
    .A1(net343),
    .A2(_03696_));
 sg13g2_nand2_1 _21460_ (.Y(_03698_),
    .A(net839),
    .B(\mem.mem_internal.code_mem[25][0] ));
 sg13g2_nor2_1 _21461_ (.A(_10422_),
    .B(net464),
    .Y(_03699_));
 sg13g2_buf_2 _21462_ (.A(_03699_),
    .X(_03700_));
 sg13g2_buf_1 _21463_ (.A(_03700_),
    .X(_03701_));
 sg13g2_nand2_1 _21464_ (.Y(_03702_),
    .A(net1054),
    .B(net177));
 sg13g2_o21ai_1 _21465_ (.B1(_03702_),
    .Y(_01498_),
    .A1(_03698_),
    .A2(net177));
 sg13g2_nand2_1 _21466_ (.Y(_03703_),
    .A(net653),
    .B(\mem.mem_internal.code_mem[25][1] ));
 sg13g2_nand2_1 _21467_ (.Y(_03704_),
    .A(net1053),
    .B(net177));
 sg13g2_o21ai_1 _21468_ (.B1(_03704_),
    .Y(_01499_),
    .A1(_03701_),
    .A2(_03703_));
 sg13g2_nand2_1 _21469_ (.Y(_03705_),
    .A(net653),
    .B(\mem.mem_internal.code_mem[25][2] ));
 sg13g2_nand2_1 _21470_ (.Y(_03706_),
    .A(net1052),
    .B(_03700_));
 sg13g2_o21ai_1 _21471_ (.B1(_03706_),
    .Y(_01500_),
    .A1(_03701_),
    .A2(_03705_));
 sg13g2_buf_1 _21472_ (.A(_03621_),
    .X(_03707_));
 sg13g2_nand2_1 _21473_ (.Y(_03708_),
    .A(net652),
    .B(\mem.mem_internal.code_mem[25][3] ));
 sg13g2_nand2_1 _21474_ (.Y(_03709_),
    .A(net1051),
    .B(_03700_));
 sg13g2_o21ai_1 _21475_ (.B1(_03709_),
    .Y(_01501_),
    .A1(net177),
    .A2(_03708_));
 sg13g2_nand2_1 _21476_ (.Y(_03710_),
    .A(net652),
    .B(\mem.mem_internal.code_mem[25][4] ));
 sg13g2_nand2_1 _21477_ (.Y(_03711_),
    .A(net1050),
    .B(_03700_));
 sg13g2_o21ai_1 _21478_ (.B1(_03711_),
    .Y(_01502_),
    .A1(net177),
    .A2(_03710_));
 sg13g2_nand2_1 _21479_ (.Y(_03712_),
    .A(_03707_),
    .B(\mem.mem_internal.code_mem[25][5] ));
 sg13g2_nand2_1 _21480_ (.Y(_03713_),
    .A(net1049),
    .B(_03700_));
 sg13g2_o21ai_1 _21481_ (.B1(_03713_),
    .Y(_01503_),
    .A1(net177),
    .A2(_03712_));
 sg13g2_nand2_1 _21482_ (.Y(_03714_),
    .A(net652),
    .B(\mem.mem_internal.code_mem[25][6] ));
 sg13g2_nand2_1 _21483_ (.Y(_03715_),
    .A(net1048),
    .B(_03700_));
 sg13g2_o21ai_1 _21484_ (.B1(_03715_),
    .Y(_01504_),
    .A1(net177),
    .A2(_03714_));
 sg13g2_nand2_1 _21485_ (.Y(_03716_),
    .A(net652),
    .B(\mem.mem_internal.code_mem[25][7] ));
 sg13g2_nand2_1 _21486_ (.Y(_03717_),
    .A(net1047),
    .B(_03700_));
 sg13g2_o21ai_1 _21487_ (.B1(_03717_),
    .Y(_01505_),
    .A1(net177),
    .A2(_03716_));
 sg13g2_nand2_1 _21488_ (.Y(_03718_),
    .A(net839),
    .B(\mem.mem_internal.code_mem[26][0] ));
 sg13g2_nor2_1 _21489_ (.A(_10444_),
    .B(_11946_),
    .Y(_03719_));
 sg13g2_buf_2 _21490_ (.A(_03719_),
    .X(_03720_));
 sg13g2_buf_1 _21491_ (.A(_03720_),
    .X(_03721_));
 sg13g2_nand2_1 _21492_ (.Y(_03722_),
    .A(net1054),
    .B(net342));
 sg13g2_o21ai_1 _21493_ (.B1(_03722_),
    .Y(_01506_),
    .A1(_03718_),
    .A2(net342));
 sg13g2_nand2_1 _21494_ (.Y(_03723_),
    .A(net652),
    .B(\mem.mem_internal.code_mem[26][1] ));
 sg13g2_nand2_1 _21495_ (.Y(_03724_),
    .A(net1053),
    .B(_03721_));
 sg13g2_o21ai_1 _21496_ (.B1(_03724_),
    .Y(_01507_),
    .A1(_03721_),
    .A2(_03723_));
 sg13g2_nand2_1 _21497_ (.Y(_03725_),
    .A(net652),
    .B(\mem.mem_internal.code_mem[26][2] ));
 sg13g2_nand2_1 _21498_ (.Y(_03726_),
    .A(net1052),
    .B(_03720_));
 sg13g2_o21ai_1 _21499_ (.B1(_03726_),
    .Y(_01508_),
    .A1(net342),
    .A2(_03725_));
 sg13g2_nand2_1 _21500_ (.Y(_03727_),
    .A(net652),
    .B(\mem.mem_internal.code_mem[26][3] ));
 sg13g2_nand2_1 _21501_ (.Y(_03728_),
    .A(net1051),
    .B(_03720_));
 sg13g2_o21ai_1 _21502_ (.B1(_03728_),
    .Y(_01509_),
    .A1(net342),
    .A2(_03727_));
 sg13g2_nand2_1 _21503_ (.Y(_03729_),
    .A(net652),
    .B(\mem.mem_internal.code_mem[26][4] ));
 sg13g2_nand2_1 _21504_ (.Y(_03730_),
    .A(net1050),
    .B(_03720_));
 sg13g2_o21ai_1 _21505_ (.B1(_03730_),
    .Y(_01510_),
    .A1(net342),
    .A2(_03729_));
 sg13g2_nand2_1 _21506_ (.Y(_03731_),
    .A(_03707_),
    .B(\mem.mem_internal.code_mem[26][5] ));
 sg13g2_nand2_1 _21507_ (.Y(_03732_),
    .A(net1049),
    .B(_03720_));
 sg13g2_o21ai_1 _21508_ (.B1(_03732_),
    .Y(_01511_),
    .A1(net342),
    .A2(_03731_));
 sg13g2_buf_1 _21509_ (.A(_03621_),
    .X(_03733_));
 sg13g2_nand2_1 _21510_ (.Y(_03734_),
    .A(net651),
    .B(\mem.mem_internal.code_mem[26][6] ));
 sg13g2_nand2_1 _21511_ (.Y(_03735_),
    .A(net1048),
    .B(_03720_));
 sg13g2_o21ai_1 _21512_ (.B1(_03735_),
    .Y(_01512_),
    .A1(net342),
    .A2(_03734_));
 sg13g2_nand2_1 _21513_ (.Y(_03736_),
    .A(net651),
    .B(\mem.mem_internal.code_mem[26][7] ));
 sg13g2_nand2_1 _21514_ (.Y(_03737_),
    .A(net1047),
    .B(_03720_));
 sg13g2_o21ai_1 _21515_ (.B1(_03737_),
    .Y(_01513_),
    .A1(net342),
    .A2(_03736_));
 sg13g2_nand2_1 _21516_ (.Y(_03738_),
    .A(net839),
    .B(\mem.mem_internal.code_mem[27][0] ));
 sg13g2_nor2_1 _21517_ (.A(_10467_),
    .B(_11946_),
    .Y(_03739_));
 sg13g2_buf_2 _21518_ (.A(_03739_),
    .X(_03740_));
 sg13g2_buf_1 _21519_ (.A(_03740_),
    .X(_03741_));
 sg13g2_nand2_1 _21520_ (.Y(_03742_),
    .A(net1054),
    .B(net341));
 sg13g2_o21ai_1 _21521_ (.B1(_03742_),
    .Y(_01514_),
    .A1(_03738_),
    .A2(net341));
 sg13g2_nand2_1 _21522_ (.Y(_03743_),
    .A(_03733_),
    .B(\mem.mem_internal.code_mem[27][1] ));
 sg13g2_nand2_1 _21523_ (.Y(_03744_),
    .A(net1053),
    .B(net341));
 sg13g2_o21ai_1 _21524_ (.B1(_03744_),
    .Y(_01515_),
    .A1(_03741_),
    .A2(_03743_));
 sg13g2_nand2_1 _21525_ (.Y(_03745_),
    .A(net651),
    .B(\mem.mem_internal.code_mem[27][2] ));
 sg13g2_nand2_1 _21526_ (.Y(_03746_),
    .A(net1052),
    .B(_03740_));
 sg13g2_o21ai_1 _21527_ (.B1(_03746_),
    .Y(_01516_),
    .A1(_03741_),
    .A2(_03745_));
 sg13g2_nand2_1 _21528_ (.Y(_03747_),
    .A(net651),
    .B(\mem.mem_internal.code_mem[27][3] ));
 sg13g2_nand2_1 _21529_ (.Y(_03748_),
    .A(net1051),
    .B(_03740_));
 sg13g2_o21ai_1 _21530_ (.B1(_03748_),
    .Y(_01517_),
    .A1(net341),
    .A2(_03747_));
 sg13g2_nand2_1 _21531_ (.Y(_03749_),
    .A(net651),
    .B(\mem.mem_internal.code_mem[27][4] ));
 sg13g2_nand2_1 _21532_ (.Y(_03750_),
    .A(net1050),
    .B(_03740_));
 sg13g2_o21ai_1 _21533_ (.B1(_03750_),
    .Y(_01518_),
    .A1(net341),
    .A2(_03749_));
 sg13g2_nand2_1 _21534_ (.Y(_03751_),
    .A(net651),
    .B(\mem.mem_internal.code_mem[27][5] ));
 sg13g2_nand2_1 _21535_ (.Y(_03752_),
    .A(net1049),
    .B(_03740_));
 sg13g2_o21ai_1 _21536_ (.B1(_03752_),
    .Y(_01519_),
    .A1(net341),
    .A2(_03751_));
 sg13g2_nand2_1 _21537_ (.Y(_03753_),
    .A(net651),
    .B(\mem.mem_internal.code_mem[27][6] ));
 sg13g2_nand2_1 _21538_ (.Y(_03754_),
    .A(net1048),
    .B(_03740_));
 sg13g2_o21ai_1 _21539_ (.B1(_03754_),
    .Y(_01520_),
    .A1(net341),
    .A2(_03753_));
 sg13g2_nand2_1 _21540_ (.Y(_03755_),
    .A(_03733_),
    .B(\mem.mem_internal.code_mem[27][7] ));
 sg13g2_nand2_1 _21541_ (.Y(_03756_),
    .A(net1047),
    .B(_03740_));
 sg13g2_o21ai_1 _21542_ (.B1(_03756_),
    .Y(_01521_),
    .A1(net341),
    .A2(_03755_));
 sg13g2_nand2_1 _21543_ (.Y(_03757_),
    .A(net839),
    .B(\mem.mem_internal.code_mem[28][0] ));
 sg13g2_nor2_1 _21544_ (.A(_10491_),
    .B(_11946_),
    .Y(_03758_));
 sg13g2_buf_1 _21545_ (.A(_03758_),
    .X(_03759_));
 sg13g2_buf_1 _21546_ (.A(_03759_),
    .X(_03760_));
 sg13g2_nand2_1 _21547_ (.Y(_03761_),
    .A(net1054),
    .B(net340));
 sg13g2_o21ai_1 _21548_ (.B1(_03761_),
    .Y(_01522_),
    .A1(_03757_),
    .A2(net340));
 sg13g2_nand2_1 _21549_ (.Y(_03762_),
    .A(net651),
    .B(\mem.mem_internal.code_mem[28][1] ));
 sg13g2_nand2_1 _21550_ (.Y(_03763_),
    .A(net1053),
    .B(_03760_));
 sg13g2_o21ai_1 _21551_ (.B1(_03763_),
    .Y(_01523_),
    .A1(_03760_),
    .A2(_03762_));
 sg13g2_buf_1 _21552_ (.A(_03621_),
    .X(_03764_));
 sg13g2_nand2_1 _21553_ (.Y(_03765_),
    .A(net650),
    .B(\mem.mem_internal.code_mem[28][2] ));
 sg13g2_nand2_1 _21554_ (.Y(_03766_),
    .A(net1052),
    .B(_03759_));
 sg13g2_o21ai_1 _21555_ (.B1(_03766_),
    .Y(_01524_),
    .A1(net340),
    .A2(_03765_));
 sg13g2_nand2_1 _21556_ (.Y(_03767_),
    .A(net650),
    .B(\mem.mem_internal.code_mem[28][3] ));
 sg13g2_nand2_1 _21557_ (.Y(_03768_),
    .A(net1051),
    .B(_03759_));
 sg13g2_o21ai_1 _21558_ (.B1(_03768_),
    .Y(_01525_),
    .A1(net340),
    .A2(_03767_));
 sg13g2_nand2_1 _21559_ (.Y(_03769_),
    .A(net650),
    .B(\mem.mem_internal.code_mem[28][4] ));
 sg13g2_nand2_1 _21560_ (.Y(_03770_),
    .A(net1050),
    .B(_03759_));
 sg13g2_o21ai_1 _21561_ (.B1(_03770_),
    .Y(_01526_),
    .A1(net340),
    .A2(_03769_));
 sg13g2_nand2_1 _21562_ (.Y(_03771_),
    .A(net650),
    .B(\mem.mem_internal.code_mem[28][5] ));
 sg13g2_nand2_1 _21563_ (.Y(_03772_),
    .A(net1049),
    .B(_03759_));
 sg13g2_o21ai_1 _21564_ (.B1(_03772_),
    .Y(_01527_),
    .A1(net340),
    .A2(_03771_));
 sg13g2_nand2_1 _21565_ (.Y(_03773_),
    .A(net650),
    .B(\mem.mem_internal.code_mem[28][6] ));
 sg13g2_nand2_1 _21566_ (.Y(_03774_),
    .A(net1048),
    .B(_03759_));
 sg13g2_o21ai_1 _21567_ (.B1(_03774_),
    .Y(_01528_),
    .A1(net340),
    .A2(_03773_));
 sg13g2_nand2_1 _21568_ (.Y(_03775_),
    .A(_03764_),
    .B(\mem.mem_internal.code_mem[28][7] ));
 sg13g2_nand2_1 _21569_ (.Y(_03776_),
    .A(net1047),
    .B(_03759_));
 sg13g2_o21ai_1 _21570_ (.B1(_03776_),
    .Y(_01529_),
    .A1(net340),
    .A2(_03775_));
 sg13g2_buf_1 _21571_ (.A(_12878_),
    .X(_03777_));
 sg13g2_nand2_1 _21572_ (.Y(_03778_),
    .A(net838),
    .B(\mem.mem_internal.code_mem[29][0] ));
 sg13g2_nor2_1 _21573_ (.A(_10513_),
    .B(_11946_),
    .Y(_03779_));
 sg13g2_buf_2 _21574_ (.A(_03779_),
    .X(_03780_));
 sg13g2_buf_1 _21575_ (.A(_03780_),
    .X(_03781_));
 sg13g2_nand2_1 _21576_ (.Y(_03782_),
    .A(net1054),
    .B(net339));
 sg13g2_o21ai_1 _21577_ (.B1(_03782_),
    .Y(_01530_),
    .A1(_03778_),
    .A2(net339));
 sg13g2_nand2_1 _21578_ (.Y(_03783_),
    .A(net650),
    .B(\mem.mem_internal.code_mem[29][1] ));
 sg13g2_nand2_1 _21579_ (.Y(_03784_),
    .A(net1053),
    .B(net339));
 sg13g2_o21ai_1 _21580_ (.B1(_03784_),
    .Y(_01531_),
    .A1(net339),
    .A2(_03783_));
 sg13g2_nand2_1 _21581_ (.Y(_03785_),
    .A(net650),
    .B(\mem.mem_internal.code_mem[29][2] ));
 sg13g2_nand2_1 _21582_ (.Y(_03786_),
    .A(net1052),
    .B(_03780_));
 sg13g2_o21ai_1 _21583_ (.B1(_03786_),
    .Y(_01532_),
    .A1(net339),
    .A2(_03785_));
 sg13g2_nand2_1 _21584_ (.Y(_03787_),
    .A(net650),
    .B(\mem.mem_internal.code_mem[29][3] ));
 sg13g2_nand2_1 _21585_ (.Y(_03788_),
    .A(net1051),
    .B(_03780_));
 sg13g2_o21ai_1 _21586_ (.B1(_03788_),
    .Y(_01533_),
    .A1(net339),
    .A2(_03787_));
 sg13g2_nand2_1 _21587_ (.Y(_03789_),
    .A(_03764_),
    .B(\mem.mem_internal.code_mem[29][4] ));
 sg13g2_nand2_1 _21588_ (.Y(_03790_),
    .A(net1050),
    .B(_03780_));
 sg13g2_o21ai_1 _21589_ (.B1(_03790_),
    .Y(_01534_),
    .A1(net339),
    .A2(_03789_));
 sg13g2_buf_1 _21590_ (.A(_03621_),
    .X(_03791_));
 sg13g2_nand2_1 _21591_ (.Y(_03792_),
    .A(_03791_),
    .B(\mem.mem_internal.code_mem[29][5] ));
 sg13g2_nand2_1 _21592_ (.Y(_03793_),
    .A(net1049),
    .B(_03780_));
 sg13g2_o21ai_1 _21593_ (.B1(_03793_),
    .Y(_01535_),
    .A1(_03781_),
    .A2(_03792_));
 sg13g2_nand2_1 _21594_ (.Y(_03794_),
    .A(_03791_),
    .B(\mem.mem_internal.code_mem[29][6] ));
 sg13g2_nand2_1 _21595_ (.Y(_03795_),
    .A(net1048),
    .B(_03780_));
 sg13g2_o21ai_1 _21596_ (.B1(_03795_),
    .Y(_01536_),
    .A1(_03781_),
    .A2(_03794_));
 sg13g2_nand2_1 _21597_ (.Y(_03796_),
    .A(net649),
    .B(\mem.mem_internal.code_mem[29][7] ));
 sg13g2_nand2_1 _21598_ (.Y(_03797_),
    .A(net1047),
    .B(_03780_));
 sg13g2_o21ai_1 _21599_ (.B1(_03797_),
    .Y(_01537_),
    .A1(net339),
    .A2(_03796_));
 sg13g2_nand2_1 _21600_ (.Y(_03798_),
    .A(net838),
    .B(\mem.mem_internal.code_mem[2][0] ));
 sg13g2_nor2_1 _21601_ (.A(net470),
    .B(net527),
    .Y(_03799_));
 sg13g2_buf_2 _21602_ (.A(_03799_),
    .X(_03800_));
 sg13g2_buf_1 _21603_ (.A(_03800_),
    .X(_03801_));
 sg13g2_nand2_1 _21604_ (.Y(_03802_),
    .A(net1054),
    .B(net176));
 sg13g2_o21ai_1 _21605_ (.B1(_03802_),
    .Y(_01538_),
    .A1(_03798_),
    .A2(net176));
 sg13g2_nand2_1 _21606_ (.Y(_03803_),
    .A(net649),
    .B(\mem.mem_internal.code_mem[2][1] ));
 sg13g2_nand2_1 _21607_ (.Y(_03804_),
    .A(net1053),
    .B(net176));
 sg13g2_o21ai_1 _21608_ (.B1(_03804_),
    .Y(_01539_),
    .A1(net176),
    .A2(_03803_));
 sg13g2_nand2_1 _21609_ (.Y(_03805_),
    .A(net649),
    .B(\mem.mem_internal.code_mem[2][2] ));
 sg13g2_nand2_1 _21610_ (.Y(_03806_),
    .A(net1052),
    .B(_03800_));
 sg13g2_o21ai_1 _21611_ (.B1(_03806_),
    .Y(_01540_),
    .A1(net176),
    .A2(_03805_));
 sg13g2_nand2_1 _21612_ (.Y(_03807_),
    .A(net649),
    .B(\mem.mem_internal.code_mem[2][3] ));
 sg13g2_nand2_1 _21613_ (.Y(_03808_),
    .A(net1051),
    .B(_03800_));
 sg13g2_o21ai_1 _21614_ (.B1(_03808_),
    .Y(_01541_),
    .A1(net176),
    .A2(_03807_));
 sg13g2_nand2_1 _21615_ (.Y(_03809_),
    .A(net649),
    .B(\mem.mem_internal.code_mem[2][4] ));
 sg13g2_nand2_1 _21616_ (.Y(_03810_),
    .A(net1050),
    .B(_03800_));
 sg13g2_o21ai_1 _21617_ (.B1(_03810_),
    .Y(_01542_),
    .A1(net176),
    .A2(_03809_));
 sg13g2_nand2_1 _21618_ (.Y(_03811_),
    .A(net649),
    .B(\mem.mem_internal.code_mem[2][5] ));
 sg13g2_nand2_1 _21619_ (.Y(_03812_),
    .A(net1049),
    .B(_03800_));
 sg13g2_o21ai_1 _21620_ (.B1(_03812_),
    .Y(_01543_),
    .A1(_03801_),
    .A2(_03811_));
 sg13g2_nand2_1 _21621_ (.Y(_03813_),
    .A(net649),
    .B(\mem.mem_internal.code_mem[2][6] ));
 sg13g2_nand2_1 _21622_ (.Y(_03814_),
    .A(net1048),
    .B(_03800_));
 sg13g2_o21ai_1 _21623_ (.B1(_03814_),
    .Y(_01544_),
    .A1(_03801_),
    .A2(_03813_));
 sg13g2_nand2_1 _21624_ (.Y(_03815_),
    .A(net649),
    .B(\mem.mem_internal.code_mem[2][7] ));
 sg13g2_nand2_1 _21625_ (.Y(_03816_),
    .A(net1047),
    .B(_03800_));
 sg13g2_o21ai_1 _21626_ (.B1(_03816_),
    .Y(_01545_),
    .A1(net176),
    .A2(_03815_));
 sg13g2_nand2_1 _21627_ (.Y(_03817_),
    .A(_03777_),
    .B(\mem.mem_internal.code_mem[30][0] ));
 sg13g2_nor2_1 _21628_ (.A(_10564_),
    .B(_11946_),
    .Y(_03818_));
 sg13g2_buf_2 _21629_ (.A(_03818_),
    .X(_03819_));
 sg13g2_buf_1 _21630_ (.A(_03819_),
    .X(_03820_));
 sg13g2_nand2_1 _21631_ (.Y(_03821_),
    .A(net1054),
    .B(net338));
 sg13g2_o21ai_1 _21632_ (.B1(_03821_),
    .Y(_01546_),
    .A1(_03817_),
    .A2(net338));
 sg13g2_buf_1 _21633_ (.A(_03042_),
    .X(_03822_));
 sg13g2_buf_1 _21634_ (.A(_03822_),
    .X(_03823_));
 sg13g2_nand2_1 _21635_ (.Y(_03824_),
    .A(net648),
    .B(\mem.mem_internal.code_mem[30][1] ));
 sg13g2_nand2_1 _21636_ (.Y(_03825_),
    .A(net1053),
    .B(net338));
 sg13g2_o21ai_1 _21637_ (.B1(_03825_),
    .Y(_01547_),
    .A1(net338),
    .A2(_03824_));
 sg13g2_nand2_1 _21638_ (.Y(_03826_),
    .A(net648),
    .B(\mem.mem_internal.code_mem[30][2] ));
 sg13g2_nand2_1 _21639_ (.Y(_03827_),
    .A(net1052),
    .B(_03819_));
 sg13g2_o21ai_1 _21640_ (.B1(_03827_),
    .Y(_01548_),
    .A1(net338),
    .A2(_03826_));
 sg13g2_nand2_1 _21641_ (.Y(_03828_),
    .A(net648),
    .B(\mem.mem_internal.code_mem[30][3] ));
 sg13g2_nand2_1 _21642_ (.Y(_03829_),
    .A(net1051),
    .B(_03819_));
 sg13g2_o21ai_1 _21643_ (.B1(_03829_),
    .Y(_01549_),
    .A1(net338),
    .A2(_03828_));
 sg13g2_nand2_1 _21644_ (.Y(_03830_),
    .A(net648),
    .B(\mem.mem_internal.code_mem[30][4] ));
 sg13g2_nand2_1 _21645_ (.Y(_03831_),
    .A(net1050),
    .B(_03819_));
 sg13g2_o21ai_1 _21646_ (.B1(_03831_),
    .Y(_01550_),
    .A1(net338),
    .A2(_03830_));
 sg13g2_nand2_1 _21647_ (.Y(_03832_),
    .A(net648),
    .B(\mem.mem_internal.code_mem[30][5] ));
 sg13g2_nand2_1 _21648_ (.Y(_03833_),
    .A(net1049),
    .B(_03819_));
 sg13g2_o21ai_1 _21649_ (.B1(_03833_),
    .Y(_01551_),
    .A1(_03820_),
    .A2(_03832_));
 sg13g2_nand2_1 _21650_ (.Y(_03834_),
    .A(_03823_),
    .B(\mem.mem_internal.code_mem[30][6] ));
 sg13g2_nand2_1 _21651_ (.Y(_03835_),
    .A(net1048),
    .B(_03819_));
 sg13g2_o21ai_1 _21652_ (.B1(_03835_),
    .Y(_01552_),
    .A1(_03820_),
    .A2(_03834_));
 sg13g2_nand2_1 _21653_ (.Y(_03836_),
    .A(_03823_),
    .B(\mem.mem_internal.code_mem[30][7] ));
 sg13g2_nand2_1 _21654_ (.Y(_03837_),
    .A(net1047),
    .B(_03819_));
 sg13g2_o21ai_1 _21655_ (.B1(_03837_),
    .Y(_01553_),
    .A1(net338),
    .A2(_03836_));
 sg13g2_nand2_1 _21656_ (.Y(_03838_),
    .A(_03777_),
    .B(\mem.mem_internal.code_mem[31][0] ));
 sg13g2_nor2_1 _21657_ (.A(_10586_),
    .B(_11946_),
    .Y(_03839_));
 sg13g2_buf_2 _21658_ (.A(_03839_),
    .X(_03840_));
 sg13g2_buf_1 _21659_ (.A(_03840_),
    .X(_03841_));
 sg13g2_buf_2 _21660_ (.A(_10251_),
    .X(_03842_));
 sg13g2_buf_1 _21661_ (.A(_03842_),
    .X(_03843_));
 sg13g2_nand2_1 _21662_ (.Y(_03844_),
    .A(_03843_),
    .B(_03841_));
 sg13g2_o21ai_1 _21663_ (.B1(_03844_),
    .Y(_01554_),
    .A1(_03838_),
    .A2(_03841_));
 sg13g2_nand2_1 _21664_ (.Y(_03845_),
    .A(net648),
    .B(\mem.mem_internal.code_mem[31][1] ));
 sg13g2_buf_2 _21665_ (.A(_10256_),
    .X(_03846_));
 sg13g2_buf_1 _21666_ (.A(_03846_),
    .X(_03847_));
 sg13g2_nand2_1 _21667_ (.Y(_03848_),
    .A(_03847_),
    .B(net337));
 sg13g2_o21ai_1 _21668_ (.B1(_03848_),
    .Y(_01555_),
    .A1(net337),
    .A2(_03845_));
 sg13g2_nand2_1 _21669_ (.Y(_03849_),
    .A(net648),
    .B(\mem.mem_internal.code_mem[31][2] ));
 sg13g2_buf_2 _21670_ (.A(_10262_),
    .X(_03850_));
 sg13g2_buf_1 _21671_ (.A(_03850_),
    .X(_03851_));
 sg13g2_nand2_1 _21672_ (.Y(_03852_),
    .A(_03851_),
    .B(_03840_));
 sg13g2_o21ai_1 _21673_ (.B1(_03852_),
    .Y(_01556_),
    .A1(net337),
    .A2(_03849_));
 sg13g2_nand2_1 _21674_ (.Y(_03853_),
    .A(net648),
    .B(\mem.mem_internal.code_mem[31][3] ));
 sg13g2_buf_2 _21675_ (.A(_10267_),
    .X(_03854_));
 sg13g2_buf_1 _21676_ (.A(_03854_),
    .X(_03855_));
 sg13g2_nand2_1 _21677_ (.Y(_03856_),
    .A(_03855_),
    .B(_03840_));
 sg13g2_o21ai_1 _21678_ (.B1(_03856_),
    .Y(_01557_),
    .A1(net337),
    .A2(_03853_));
 sg13g2_buf_1 _21679_ (.A(_03822_),
    .X(_03857_));
 sg13g2_nand2_1 _21680_ (.Y(_03858_),
    .A(net647),
    .B(\mem.mem_internal.code_mem[31][4] ));
 sg13g2_buf_2 _21681_ (.A(_10272_),
    .X(_03859_));
 sg13g2_buf_1 _21682_ (.A(_03859_),
    .X(_03860_));
 sg13g2_nand2_1 _21683_ (.Y(_03861_),
    .A(_03860_),
    .B(_03840_));
 sg13g2_o21ai_1 _21684_ (.B1(_03861_),
    .Y(_01558_),
    .A1(net337),
    .A2(_03858_));
 sg13g2_nand2_1 _21685_ (.Y(_03862_),
    .A(net647),
    .B(\mem.mem_internal.code_mem[31][5] ));
 sg13g2_buf_2 _21686_ (.A(_10277_),
    .X(_03863_));
 sg13g2_buf_1 _21687_ (.A(_03863_),
    .X(_03864_));
 sg13g2_nand2_1 _21688_ (.Y(_03865_),
    .A(_03864_),
    .B(_03840_));
 sg13g2_o21ai_1 _21689_ (.B1(_03865_),
    .Y(_01559_),
    .A1(net337),
    .A2(_03862_));
 sg13g2_nand2_1 _21690_ (.Y(_03866_),
    .A(_03857_),
    .B(\mem.mem_internal.code_mem[31][6] ));
 sg13g2_buf_2 _21691_ (.A(_10282_),
    .X(_03867_));
 sg13g2_buf_1 _21692_ (.A(_03867_),
    .X(_03868_));
 sg13g2_nand2_1 _21693_ (.Y(_03869_),
    .A(_03868_),
    .B(_03840_));
 sg13g2_o21ai_1 _21694_ (.B1(_03869_),
    .Y(_01560_),
    .A1(net337),
    .A2(_03866_));
 sg13g2_nand2_1 _21695_ (.Y(_03870_),
    .A(_03857_),
    .B(\mem.mem_internal.code_mem[31][7] ));
 sg13g2_buf_2 _21696_ (.A(_10287_),
    .X(_03871_));
 sg13g2_buf_1 _21697_ (.A(_03871_),
    .X(_03872_));
 sg13g2_nand2_1 _21698_ (.Y(_03873_),
    .A(_03872_),
    .B(_03840_));
 sg13g2_o21ai_1 _21699_ (.B1(_03873_),
    .Y(_01561_),
    .A1(net337),
    .A2(_03870_));
 sg13g2_nand2_1 _21700_ (.Y(_03874_),
    .A(net838),
    .B(\mem.mem_internal.code_mem[32][0] ));
 sg13g2_nand2_1 _21701_ (.Y(_03875_),
    .A(_10234_),
    .B(_10298_));
 sg13g2_buf_2 _21702_ (.A(_03875_),
    .X(_03876_));
 sg13g2_buf_1 _21703_ (.A(_03876_),
    .X(_03877_));
 sg13g2_nor2_1 _21704_ (.A(_10232_),
    .B(net458),
    .Y(_03878_));
 sg13g2_buf_2 _21705_ (.A(_03878_),
    .X(_03879_));
 sg13g2_buf_1 _21706_ (.A(_03879_),
    .X(_03880_));
 sg13g2_nand2_1 _21707_ (.Y(_03881_),
    .A(net1046),
    .B(net175));
 sg13g2_o21ai_1 _21708_ (.B1(_03881_),
    .Y(_01562_),
    .A1(_03874_),
    .A2(net175));
 sg13g2_nand2_1 _21709_ (.Y(_03882_),
    .A(net647),
    .B(\mem.mem_internal.code_mem[32][1] ));
 sg13g2_nand2_1 _21710_ (.Y(_03883_),
    .A(net1045),
    .B(net175));
 sg13g2_o21ai_1 _21711_ (.B1(_03883_),
    .Y(_01563_),
    .A1(net175),
    .A2(_03882_));
 sg13g2_nand2_1 _21712_ (.Y(_03884_),
    .A(net647),
    .B(\mem.mem_internal.code_mem[32][2] ));
 sg13g2_nand2_1 _21713_ (.Y(_03885_),
    .A(net1044),
    .B(_03879_));
 sg13g2_o21ai_1 _21714_ (.B1(_03885_),
    .Y(_01564_),
    .A1(_03880_),
    .A2(_03884_));
 sg13g2_nand2_1 _21715_ (.Y(_03886_),
    .A(net647),
    .B(\mem.mem_internal.code_mem[32][3] ));
 sg13g2_nand2_1 _21716_ (.Y(_03887_),
    .A(net1043),
    .B(_03879_));
 sg13g2_o21ai_1 _21717_ (.B1(_03887_),
    .Y(_01565_),
    .A1(_03880_),
    .A2(_03886_));
 sg13g2_nand2_1 _21718_ (.Y(_03888_),
    .A(net647),
    .B(\mem.mem_internal.code_mem[32][4] ));
 sg13g2_nand2_1 _21719_ (.Y(_03889_),
    .A(net1042),
    .B(_03879_));
 sg13g2_o21ai_1 _21720_ (.B1(_03889_),
    .Y(_01566_),
    .A1(net175),
    .A2(_03888_));
 sg13g2_nand2_1 _21721_ (.Y(_03890_),
    .A(net647),
    .B(\mem.mem_internal.code_mem[32][5] ));
 sg13g2_nand2_1 _21722_ (.Y(_03891_),
    .A(net1041),
    .B(_03879_));
 sg13g2_o21ai_1 _21723_ (.B1(_03891_),
    .Y(_01567_),
    .A1(net175),
    .A2(_03890_));
 sg13g2_nand2_1 _21724_ (.Y(_03892_),
    .A(net647),
    .B(\mem.mem_internal.code_mem[32][6] ));
 sg13g2_nand2_1 _21725_ (.Y(_03893_),
    .A(net1040),
    .B(_03879_));
 sg13g2_o21ai_1 _21726_ (.B1(_03893_),
    .Y(_01568_),
    .A1(net175),
    .A2(_03892_));
 sg13g2_buf_1 _21727_ (.A(_03822_),
    .X(_03894_));
 sg13g2_nand2_1 _21728_ (.Y(_03895_),
    .A(net646),
    .B(\mem.mem_internal.code_mem[32][7] ));
 sg13g2_nand2_1 _21729_ (.Y(_03896_),
    .A(net1039),
    .B(_03879_));
 sg13g2_o21ai_1 _21730_ (.B1(_03896_),
    .Y(_01569_),
    .A1(net175),
    .A2(_03895_));
 sg13g2_nand2_1 _21731_ (.Y(_03897_),
    .A(net838),
    .B(\mem.mem_internal.code_mem[33][0] ));
 sg13g2_nor2_1 _21732_ (.A(_10632_),
    .B(net458),
    .Y(_03898_));
 sg13g2_buf_2 _21733_ (.A(_03898_),
    .X(_03899_));
 sg13g2_buf_1 _21734_ (.A(_03899_),
    .X(_03900_));
 sg13g2_nand2_1 _21735_ (.Y(_03901_),
    .A(net1046),
    .B(net174));
 sg13g2_o21ai_1 _21736_ (.B1(_03901_),
    .Y(_01570_),
    .A1(_03897_),
    .A2(net174));
 sg13g2_nand2_1 _21737_ (.Y(_03902_),
    .A(net646),
    .B(\mem.mem_internal.code_mem[33][1] ));
 sg13g2_nand2_1 _21738_ (.Y(_03903_),
    .A(net1045),
    .B(net174));
 sg13g2_o21ai_1 _21739_ (.B1(_03903_),
    .Y(_01571_),
    .A1(net174),
    .A2(_03902_));
 sg13g2_nand2_1 _21740_ (.Y(_03904_),
    .A(net646),
    .B(\mem.mem_internal.code_mem[33][2] ));
 sg13g2_nand2_1 _21741_ (.Y(_03905_),
    .A(net1044),
    .B(_03899_));
 sg13g2_o21ai_1 _21742_ (.B1(_03905_),
    .Y(_01572_),
    .A1(net174),
    .A2(_03904_));
 sg13g2_nand2_1 _21743_ (.Y(_03906_),
    .A(net646),
    .B(\mem.mem_internal.code_mem[33][3] ));
 sg13g2_nand2_1 _21744_ (.Y(_03907_),
    .A(net1043),
    .B(_03899_));
 sg13g2_o21ai_1 _21745_ (.B1(_03907_),
    .Y(_01573_),
    .A1(net174),
    .A2(_03906_));
 sg13g2_nand2_1 _21746_ (.Y(_03908_),
    .A(net646),
    .B(\mem.mem_internal.code_mem[33][4] ));
 sg13g2_nand2_1 _21747_ (.Y(_03909_),
    .A(net1042),
    .B(_03899_));
 sg13g2_o21ai_1 _21748_ (.B1(_03909_),
    .Y(_01574_),
    .A1(net174),
    .A2(_03908_));
 sg13g2_nand2_1 _21749_ (.Y(_03910_),
    .A(net646),
    .B(\mem.mem_internal.code_mem[33][5] ));
 sg13g2_nand2_1 _21750_ (.Y(_03911_),
    .A(net1041),
    .B(_03899_));
 sg13g2_o21ai_1 _21751_ (.B1(_03911_),
    .Y(_01575_),
    .A1(net174),
    .A2(_03910_));
 sg13g2_nand2_1 _21752_ (.Y(_03912_),
    .A(_03894_),
    .B(\mem.mem_internal.code_mem[33][6] ));
 sg13g2_nand2_1 _21753_ (.Y(_03913_),
    .A(net1040),
    .B(_03899_));
 sg13g2_o21ai_1 _21754_ (.B1(_03913_),
    .Y(_01576_),
    .A1(_03900_),
    .A2(_03912_));
 sg13g2_nand2_1 _21755_ (.Y(_03914_),
    .A(_03894_),
    .B(\mem.mem_internal.code_mem[33][7] ));
 sg13g2_nand2_1 _21756_ (.Y(_03915_),
    .A(net1039),
    .B(_03899_));
 sg13g2_o21ai_1 _21757_ (.B1(_03915_),
    .Y(_01577_),
    .A1(_03900_),
    .A2(_03914_));
 sg13g2_nand2_1 _21758_ (.Y(_03916_),
    .A(net838),
    .B(\mem.mem_internal.code_mem[34][0] ));
 sg13g2_nor2_1 _21759_ (.A(_10656_),
    .B(_03877_),
    .Y(_03917_));
 sg13g2_buf_2 _21760_ (.A(_03917_),
    .X(_03918_));
 sg13g2_buf_1 _21761_ (.A(_03918_),
    .X(_03919_));
 sg13g2_nand2_1 _21762_ (.Y(_03920_),
    .A(net1046),
    .B(net173));
 sg13g2_o21ai_1 _21763_ (.B1(_03920_),
    .Y(_01578_),
    .A1(_03916_),
    .A2(net173));
 sg13g2_nand2_1 _21764_ (.Y(_03921_),
    .A(net646),
    .B(\mem.mem_internal.code_mem[34][1] ));
 sg13g2_nand2_1 _21765_ (.Y(_03922_),
    .A(net1045),
    .B(net173));
 sg13g2_o21ai_1 _21766_ (.B1(_03922_),
    .Y(_01579_),
    .A1(net173),
    .A2(_03921_));
 sg13g2_nand2_1 _21767_ (.Y(_03923_),
    .A(net646),
    .B(\mem.mem_internal.code_mem[34][2] ));
 sg13g2_nand2_1 _21768_ (.Y(_03924_),
    .A(net1044),
    .B(_03918_));
 sg13g2_o21ai_1 _21769_ (.B1(_03924_),
    .Y(_01580_),
    .A1(net173),
    .A2(_03923_));
 sg13g2_buf_1 _21770_ (.A(_03822_),
    .X(_03925_));
 sg13g2_nand2_1 _21771_ (.Y(_03926_),
    .A(net645),
    .B(\mem.mem_internal.code_mem[34][3] ));
 sg13g2_nand2_1 _21772_ (.Y(_03927_),
    .A(net1043),
    .B(_03918_));
 sg13g2_o21ai_1 _21773_ (.B1(_03927_),
    .Y(_01581_),
    .A1(net173),
    .A2(_03926_));
 sg13g2_nand2_1 _21774_ (.Y(_03928_),
    .A(net645),
    .B(\mem.mem_internal.code_mem[34][4] ));
 sg13g2_nand2_1 _21775_ (.Y(_03929_),
    .A(net1042),
    .B(_03918_));
 sg13g2_o21ai_1 _21776_ (.B1(_03929_),
    .Y(_01582_),
    .A1(net173),
    .A2(_03928_));
 sg13g2_nand2_1 _21777_ (.Y(_03930_),
    .A(net645),
    .B(\mem.mem_internal.code_mem[34][5] ));
 sg13g2_nand2_1 _21778_ (.Y(_03931_),
    .A(net1041),
    .B(_03918_));
 sg13g2_o21ai_1 _21779_ (.B1(_03931_),
    .Y(_01583_),
    .A1(net173),
    .A2(_03930_));
 sg13g2_nand2_1 _21780_ (.Y(_03932_),
    .A(net645),
    .B(\mem.mem_internal.code_mem[34][6] ));
 sg13g2_nand2_1 _21781_ (.Y(_03933_),
    .A(net1040),
    .B(_03918_));
 sg13g2_o21ai_1 _21782_ (.B1(_03933_),
    .Y(_01584_),
    .A1(_03919_),
    .A2(_03932_));
 sg13g2_nand2_1 _21783_ (.Y(_03934_),
    .A(net645),
    .B(\mem.mem_internal.code_mem[34][7] ));
 sg13g2_nand2_1 _21784_ (.Y(_03935_),
    .A(net1039),
    .B(_03918_));
 sg13g2_o21ai_1 _21785_ (.B1(_03935_),
    .Y(_01585_),
    .A1(_03919_),
    .A2(_03934_));
 sg13g2_nand2_1 _21786_ (.Y(_03936_),
    .A(net838),
    .B(\mem.mem_internal.code_mem[35][0] ));
 sg13g2_nor2_1 _21787_ (.A(_10679_),
    .B(_03877_),
    .Y(_03937_));
 sg13g2_buf_2 _21788_ (.A(_03937_),
    .X(_03938_));
 sg13g2_buf_1 _21789_ (.A(_03938_),
    .X(_03939_));
 sg13g2_nand2_1 _21790_ (.Y(_03940_),
    .A(net1046),
    .B(net172));
 sg13g2_o21ai_1 _21791_ (.B1(_03940_),
    .Y(_01586_),
    .A1(_03936_),
    .A2(net172));
 sg13g2_nand2_1 _21792_ (.Y(_03941_),
    .A(net645),
    .B(\mem.mem_internal.code_mem[35][1] ));
 sg13g2_nand2_1 _21793_ (.Y(_03942_),
    .A(net1045),
    .B(net172));
 sg13g2_o21ai_1 _21794_ (.B1(_03942_),
    .Y(_01587_),
    .A1(net172),
    .A2(_03941_));
 sg13g2_nand2_1 _21795_ (.Y(_03943_),
    .A(_03925_),
    .B(\mem.mem_internal.code_mem[35][2] ));
 sg13g2_nand2_1 _21796_ (.Y(_03944_),
    .A(net1044),
    .B(_03938_));
 sg13g2_o21ai_1 _21797_ (.B1(_03944_),
    .Y(_01588_),
    .A1(_03939_),
    .A2(_03943_));
 sg13g2_nand2_1 _21798_ (.Y(_03945_),
    .A(_03925_),
    .B(\mem.mem_internal.code_mem[35][3] ));
 sg13g2_nand2_1 _21799_ (.Y(_03946_),
    .A(net1043),
    .B(_03938_));
 sg13g2_o21ai_1 _21800_ (.B1(_03946_),
    .Y(_01589_),
    .A1(net172),
    .A2(_03945_));
 sg13g2_nand2_1 _21801_ (.Y(_03947_),
    .A(net645),
    .B(\mem.mem_internal.code_mem[35][4] ));
 sg13g2_nand2_1 _21802_ (.Y(_03948_),
    .A(net1042),
    .B(_03938_));
 sg13g2_o21ai_1 _21803_ (.B1(_03948_),
    .Y(_01590_),
    .A1(net172),
    .A2(_03947_));
 sg13g2_nand2_1 _21804_ (.Y(_03949_),
    .A(net645),
    .B(\mem.mem_internal.code_mem[35][5] ));
 sg13g2_nand2_1 _21805_ (.Y(_03950_),
    .A(net1041),
    .B(_03938_));
 sg13g2_o21ai_1 _21806_ (.B1(_03950_),
    .Y(_01591_),
    .A1(_03939_),
    .A2(_03949_));
 sg13g2_buf_1 _21807_ (.A(_03822_),
    .X(_03951_));
 sg13g2_nand2_1 _21808_ (.Y(_03952_),
    .A(_03951_),
    .B(\mem.mem_internal.code_mem[35][6] ));
 sg13g2_nand2_1 _21809_ (.Y(_03953_),
    .A(net1040),
    .B(_03938_));
 sg13g2_o21ai_1 _21810_ (.B1(_03953_),
    .Y(_01592_),
    .A1(net172),
    .A2(_03952_));
 sg13g2_nand2_1 _21811_ (.Y(_03954_),
    .A(_03951_),
    .B(\mem.mem_internal.code_mem[35][7] ));
 sg13g2_nand2_1 _21812_ (.Y(_03955_),
    .A(net1039),
    .B(_03938_));
 sg13g2_o21ai_1 _21813_ (.B1(_03955_),
    .Y(_01593_),
    .A1(net172),
    .A2(_03954_));
 sg13g2_nand2_1 _21814_ (.Y(_03956_),
    .A(net838),
    .B(\mem.mem_internal.code_mem[36][0] ));
 sg13g2_nor2_1 _21815_ (.A(_10295_),
    .B(net458),
    .Y(_03957_));
 sg13g2_buf_2 _21816_ (.A(_03957_),
    .X(_03958_));
 sg13g2_buf_1 _21817_ (.A(_03958_),
    .X(_03959_));
 sg13g2_nand2_1 _21818_ (.Y(_03960_),
    .A(net1046),
    .B(net171));
 sg13g2_o21ai_1 _21819_ (.B1(_03960_),
    .Y(_01594_),
    .A1(_03956_),
    .A2(net171));
 sg13g2_nand2_1 _21820_ (.Y(_03961_),
    .A(net644),
    .B(\mem.mem_internal.code_mem[36][1] ));
 sg13g2_nand2_1 _21821_ (.Y(_03962_),
    .A(net1045),
    .B(net171));
 sg13g2_o21ai_1 _21822_ (.B1(_03962_),
    .Y(_01595_),
    .A1(_03959_),
    .A2(_03961_));
 sg13g2_nand2_1 _21823_ (.Y(_03963_),
    .A(net644),
    .B(\mem.mem_internal.code_mem[36][2] ));
 sg13g2_nand2_1 _21824_ (.Y(_03964_),
    .A(net1044),
    .B(_03958_));
 sg13g2_o21ai_1 _21825_ (.B1(_03964_),
    .Y(_01596_),
    .A1(net171),
    .A2(_03963_));
 sg13g2_nand2_1 _21826_ (.Y(_03965_),
    .A(net644),
    .B(\mem.mem_internal.code_mem[36][3] ));
 sg13g2_nand2_1 _21827_ (.Y(_03966_),
    .A(net1043),
    .B(_03958_));
 sg13g2_o21ai_1 _21828_ (.B1(_03966_),
    .Y(_01597_),
    .A1(net171),
    .A2(_03965_));
 sg13g2_nand2_1 _21829_ (.Y(_03967_),
    .A(net644),
    .B(\mem.mem_internal.code_mem[36][4] ));
 sg13g2_nand2_1 _21830_ (.Y(_03968_),
    .A(net1042),
    .B(_03958_));
 sg13g2_o21ai_1 _21831_ (.B1(_03968_),
    .Y(_01598_),
    .A1(net171),
    .A2(_03967_));
 sg13g2_nand2_1 _21832_ (.Y(_03969_),
    .A(net644),
    .B(\mem.mem_internal.code_mem[36][5] ));
 sg13g2_nand2_1 _21833_ (.Y(_03970_),
    .A(net1041),
    .B(_03958_));
 sg13g2_o21ai_1 _21834_ (.B1(_03970_),
    .Y(_01599_),
    .A1(_03959_),
    .A2(_03969_));
 sg13g2_nand2_1 _21835_ (.Y(_03971_),
    .A(net644),
    .B(\mem.mem_internal.code_mem[36][6] ));
 sg13g2_nand2_1 _21836_ (.Y(_03972_),
    .A(net1040),
    .B(_03958_));
 sg13g2_o21ai_1 _21837_ (.B1(_03972_),
    .Y(_01600_),
    .A1(net171),
    .A2(_03971_));
 sg13g2_nand2_1 _21838_ (.Y(_03973_),
    .A(net644),
    .B(\mem.mem_internal.code_mem[36][7] ));
 sg13g2_nand2_1 _21839_ (.Y(_03974_),
    .A(net1039),
    .B(_03958_));
 sg13g2_o21ai_1 _21840_ (.B1(_03974_),
    .Y(_01601_),
    .A1(net171),
    .A2(_03973_));
 sg13g2_nand2_1 _21841_ (.Y(_03975_),
    .A(net838),
    .B(\mem.mem_internal.code_mem[37][0] ));
 sg13g2_nor2_1 _21842_ (.A(_10325_),
    .B(net458),
    .Y(_03976_));
 sg13g2_buf_2 _21843_ (.A(_03976_),
    .X(_03977_));
 sg13g2_buf_1 _21844_ (.A(_03977_),
    .X(_03978_));
 sg13g2_nand2_1 _21845_ (.Y(_03979_),
    .A(net1046),
    .B(net170));
 sg13g2_o21ai_1 _21846_ (.B1(_03979_),
    .Y(_01602_),
    .A1(_03975_),
    .A2(net170));
 sg13g2_nand2_1 _21847_ (.Y(_03980_),
    .A(net644),
    .B(\mem.mem_internal.code_mem[37][1] ));
 sg13g2_nand2_1 _21848_ (.Y(_03981_),
    .A(net1045),
    .B(net170));
 sg13g2_o21ai_1 _21849_ (.B1(_03981_),
    .Y(_01603_),
    .A1(_03978_),
    .A2(_03980_));
 sg13g2_buf_1 _21850_ (.A(_03822_),
    .X(_03982_));
 sg13g2_nand2_1 _21851_ (.Y(_03983_),
    .A(_03982_),
    .B(\mem.mem_internal.code_mem[37][2] ));
 sg13g2_nand2_1 _21852_ (.Y(_03984_),
    .A(net1044),
    .B(_03977_));
 sg13g2_o21ai_1 _21853_ (.B1(_03984_),
    .Y(_01604_),
    .A1(net170),
    .A2(_03983_));
 sg13g2_nand2_1 _21854_ (.Y(_03985_),
    .A(net643),
    .B(\mem.mem_internal.code_mem[37][3] ));
 sg13g2_nand2_1 _21855_ (.Y(_03986_),
    .A(net1043),
    .B(_03977_));
 sg13g2_o21ai_1 _21856_ (.B1(_03986_),
    .Y(_01605_),
    .A1(net170),
    .A2(_03985_));
 sg13g2_nand2_1 _21857_ (.Y(_03987_),
    .A(net643),
    .B(\mem.mem_internal.code_mem[37][4] ));
 sg13g2_nand2_1 _21858_ (.Y(_03988_),
    .A(net1042),
    .B(_03977_));
 sg13g2_o21ai_1 _21859_ (.B1(_03988_),
    .Y(_01606_),
    .A1(net170),
    .A2(_03987_));
 sg13g2_nand2_1 _21860_ (.Y(_03989_),
    .A(_03982_),
    .B(\mem.mem_internal.code_mem[37][5] ));
 sg13g2_nand2_1 _21861_ (.Y(_03990_),
    .A(net1041),
    .B(_03977_));
 sg13g2_o21ai_1 _21862_ (.B1(_03990_),
    .Y(_01607_),
    .A1(_03978_),
    .A2(_03989_));
 sg13g2_nand2_1 _21863_ (.Y(_03991_),
    .A(net643),
    .B(\mem.mem_internal.code_mem[37][6] ));
 sg13g2_nand2_1 _21864_ (.Y(_03992_),
    .A(net1040),
    .B(_03977_));
 sg13g2_o21ai_1 _21865_ (.B1(_03992_),
    .Y(_01608_),
    .A1(net170),
    .A2(_03991_));
 sg13g2_nand2_1 _21866_ (.Y(_03993_),
    .A(net643),
    .B(\mem.mem_internal.code_mem[37][7] ));
 sg13g2_nand2_1 _21867_ (.Y(_03994_),
    .A(net1039),
    .B(_03977_));
 sg13g2_o21ai_1 _21868_ (.B1(_03994_),
    .Y(_01609_),
    .A1(net170),
    .A2(_03993_));
 sg13g2_buf_1 _21869_ (.A(_12878_),
    .X(_03995_));
 sg13g2_nand2_1 _21870_ (.Y(_03996_),
    .A(net837),
    .B(\mem.mem_internal.code_mem[38][0] ));
 sg13g2_nor2_1 _21871_ (.A(net779),
    .B(net458),
    .Y(_03997_));
 sg13g2_buf_2 _21872_ (.A(_03997_),
    .X(_03998_));
 sg13g2_buf_1 _21873_ (.A(_03998_),
    .X(_03999_));
 sg13g2_nand2_1 _21874_ (.Y(_04000_),
    .A(net1046),
    .B(net169));
 sg13g2_o21ai_1 _21875_ (.B1(_04000_),
    .Y(_01610_),
    .A1(_03996_),
    .A2(_03999_));
 sg13g2_nand2_1 _21876_ (.Y(_04001_),
    .A(net643),
    .B(\mem.mem_internal.code_mem[38][1] ));
 sg13g2_nand2_1 _21877_ (.Y(_04002_),
    .A(net1045),
    .B(net169));
 sg13g2_o21ai_1 _21878_ (.B1(_04002_),
    .Y(_01611_),
    .A1(net169),
    .A2(_04001_));
 sg13g2_nand2_1 _21879_ (.Y(_04003_),
    .A(net643),
    .B(\mem.mem_internal.code_mem[38][2] ));
 sg13g2_nand2_1 _21880_ (.Y(_04004_),
    .A(net1044),
    .B(_03998_));
 sg13g2_o21ai_1 _21881_ (.B1(_04004_),
    .Y(_01612_),
    .A1(net169),
    .A2(_04003_));
 sg13g2_nand2_1 _21882_ (.Y(_04005_),
    .A(net643),
    .B(\mem.mem_internal.code_mem[38][3] ));
 sg13g2_nand2_1 _21883_ (.Y(_04006_),
    .A(net1043),
    .B(_03998_));
 sg13g2_o21ai_1 _21884_ (.B1(_04006_),
    .Y(_01613_),
    .A1(net169),
    .A2(_04005_));
 sg13g2_nand2_1 _21885_ (.Y(_04007_),
    .A(net643),
    .B(\mem.mem_internal.code_mem[38][4] ));
 sg13g2_nand2_1 _21886_ (.Y(_04008_),
    .A(net1042),
    .B(_03998_));
 sg13g2_o21ai_1 _21887_ (.B1(_04008_),
    .Y(_01614_),
    .A1(net169),
    .A2(_04007_));
 sg13g2_buf_1 _21888_ (.A(_03822_),
    .X(_04009_));
 sg13g2_nand2_1 _21889_ (.Y(_04010_),
    .A(_04009_),
    .B(\mem.mem_internal.code_mem[38][5] ));
 sg13g2_nand2_1 _21890_ (.Y(_04011_),
    .A(net1041),
    .B(_03998_));
 sg13g2_o21ai_1 _21891_ (.B1(_04011_),
    .Y(_01615_),
    .A1(_03999_),
    .A2(_04010_));
 sg13g2_nand2_1 _21892_ (.Y(_04012_),
    .A(net642),
    .B(\mem.mem_internal.code_mem[38][6] ));
 sg13g2_nand2_1 _21893_ (.Y(_04013_),
    .A(net1040),
    .B(_03998_));
 sg13g2_o21ai_1 _21894_ (.B1(_04013_),
    .Y(_01616_),
    .A1(net169),
    .A2(_04012_));
 sg13g2_nand2_1 _21895_ (.Y(_04014_),
    .A(net642),
    .B(\mem.mem_internal.code_mem[38][7] ));
 sg13g2_nand2_1 _21896_ (.Y(_04015_),
    .A(net1039),
    .B(_03998_));
 sg13g2_o21ai_1 _21897_ (.B1(_04015_),
    .Y(_01617_),
    .A1(net169),
    .A2(_04014_));
 sg13g2_nand2_1 _21898_ (.Y(_04016_),
    .A(_03995_),
    .B(\mem.mem_internal.code_mem[39][0] ));
 sg13g2_nor2_1 _21899_ (.A(_10372_),
    .B(net458),
    .Y(_04017_));
 sg13g2_buf_2 _21900_ (.A(_04017_),
    .X(_04018_));
 sg13g2_buf_1 _21901_ (.A(_04018_),
    .X(_04019_));
 sg13g2_nand2_1 _21902_ (.Y(_04020_),
    .A(net1046),
    .B(net168));
 sg13g2_o21ai_1 _21903_ (.B1(_04020_),
    .Y(_01618_),
    .A1(_04016_),
    .A2(_04019_));
 sg13g2_nand2_1 _21904_ (.Y(_04021_),
    .A(net642),
    .B(\mem.mem_internal.code_mem[39][1] ));
 sg13g2_nand2_1 _21905_ (.Y(_04022_),
    .A(net1045),
    .B(net168));
 sg13g2_o21ai_1 _21906_ (.B1(_04022_),
    .Y(_01619_),
    .A1(net168),
    .A2(_04021_));
 sg13g2_nand2_1 _21907_ (.Y(_04023_),
    .A(net642),
    .B(\mem.mem_internal.code_mem[39][2] ));
 sg13g2_nand2_1 _21908_ (.Y(_04024_),
    .A(net1044),
    .B(_04018_));
 sg13g2_o21ai_1 _21909_ (.B1(_04024_),
    .Y(_01620_),
    .A1(net168),
    .A2(_04023_));
 sg13g2_nand2_1 _21910_ (.Y(_04025_),
    .A(net642),
    .B(\mem.mem_internal.code_mem[39][3] ));
 sg13g2_nand2_1 _21911_ (.Y(_04026_),
    .A(net1043),
    .B(_04018_));
 sg13g2_o21ai_1 _21912_ (.B1(_04026_),
    .Y(_01621_),
    .A1(net168),
    .A2(_04025_));
 sg13g2_nand2_1 _21913_ (.Y(_04027_),
    .A(net642),
    .B(\mem.mem_internal.code_mem[39][4] ));
 sg13g2_nand2_1 _21914_ (.Y(_04028_),
    .A(net1042),
    .B(_04018_));
 sg13g2_o21ai_1 _21915_ (.B1(_04028_),
    .Y(_01622_),
    .A1(net168),
    .A2(_04027_));
 sg13g2_nand2_1 _21916_ (.Y(_04029_),
    .A(_04009_),
    .B(\mem.mem_internal.code_mem[39][5] ));
 sg13g2_nand2_1 _21917_ (.Y(_04030_),
    .A(net1041),
    .B(_04018_));
 sg13g2_o21ai_1 _21918_ (.B1(_04030_),
    .Y(_01623_),
    .A1(_04019_),
    .A2(_04029_));
 sg13g2_nand2_1 _21919_ (.Y(_04031_),
    .A(net642),
    .B(\mem.mem_internal.code_mem[39][6] ));
 sg13g2_nand2_1 _21920_ (.Y(_04032_),
    .A(net1040),
    .B(_04018_));
 sg13g2_o21ai_1 _21921_ (.B1(_04032_),
    .Y(_01624_),
    .A1(net168),
    .A2(_04031_));
 sg13g2_nand2_1 _21922_ (.Y(_04033_),
    .A(net642),
    .B(\mem.mem_internal.code_mem[39][7] ));
 sg13g2_nand2_1 _21923_ (.Y(_04034_),
    .A(net1039),
    .B(_04018_));
 sg13g2_o21ai_1 _21924_ (.B1(_04034_),
    .Y(_01625_),
    .A1(net168),
    .A2(_04033_));
 sg13g2_nand2_1 _21925_ (.Y(_04035_),
    .A(_03995_),
    .B(\mem.mem_internal.code_mem[3][0] ));
 sg13g2_nor2_1 _21926_ (.A(net470),
    .B(net526),
    .Y(_04036_));
 sg13g2_buf_2 _21927_ (.A(_04036_),
    .X(_04037_));
 sg13g2_buf_1 _21928_ (.A(_04037_),
    .X(_04038_));
 sg13g2_nand2_1 _21929_ (.Y(_04039_),
    .A(_03843_),
    .B(net167));
 sg13g2_o21ai_1 _21930_ (.B1(_04039_),
    .Y(_01626_),
    .A1(_04035_),
    .A2(net167));
 sg13g2_buf_1 _21931_ (.A(_03042_),
    .X(_04040_));
 sg13g2_buf_1 _21932_ (.A(_04040_),
    .X(_04041_));
 sg13g2_nand2_1 _21933_ (.Y(_04042_),
    .A(net641),
    .B(\mem.mem_internal.code_mem[3][1] ));
 sg13g2_nand2_1 _21934_ (.Y(_04043_),
    .A(_03847_),
    .B(_04038_));
 sg13g2_o21ai_1 _21935_ (.B1(_04043_),
    .Y(_01627_),
    .A1(_04038_),
    .A2(_04042_));
 sg13g2_nand2_1 _21936_ (.Y(_04044_),
    .A(net641),
    .B(\mem.mem_internal.code_mem[3][2] ));
 sg13g2_nand2_1 _21937_ (.Y(_04045_),
    .A(_03851_),
    .B(_04037_));
 sg13g2_o21ai_1 _21938_ (.B1(_04045_),
    .Y(_01628_),
    .A1(net167),
    .A2(_04044_));
 sg13g2_nand2_1 _21939_ (.Y(_04046_),
    .A(net641),
    .B(\mem.mem_internal.code_mem[3][3] ));
 sg13g2_nand2_1 _21940_ (.Y(_04047_),
    .A(_03855_),
    .B(_04037_));
 sg13g2_o21ai_1 _21941_ (.B1(_04047_),
    .Y(_01629_),
    .A1(net167),
    .A2(_04046_));
 sg13g2_nand2_1 _21942_ (.Y(_04048_),
    .A(net641),
    .B(\mem.mem_internal.code_mem[3][4] ));
 sg13g2_nand2_1 _21943_ (.Y(_04049_),
    .A(_03860_),
    .B(_04037_));
 sg13g2_o21ai_1 _21944_ (.B1(_04049_),
    .Y(_01630_),
    .A1(net167),
    .A2(_04048_));
 sg13g2_nand2_1 _21945_ (.Y(_04050_),
    .A(net641),
    .B(\mem.mem_internal.code_mem[3][5] ));
 sg13g2_nand2_1 _21946_ (.Y(_04051_),
    .A(_03864_),
    .B(_04037_));
 sg13g2_o21ai_1 _21947_ (.B1(_04051_),
    .Y(_01631_),
    .A1(net167),
    .A2(_04050_));
 sg13g2_nand2_1 _21948_ (.Y(_04052_),
    .A(_04041_),
    .B(\mem.mem_internal.code_mem[3][6] ));
 sg13g2_nand2_1 _21949_ (.Y(_04053_),
    .A(_03868_),
    .B(_04037_));
 sg13g2_o21ai_1 _21950_ (.B1(_04053_),
    .Y(_01632_),
    .A1(net167),
    .A2(_04052_));
 sg13g2_nand2_1 _21951_ (.Y(_04054_),
    .A(_04041_),
    .B(\mem.mem_internal.code_mem[3][7] ));
 sg13g2_nand2_1 _21952_ (.Y(_04055_),
    .A(_03872_),
    .B(_04037_));
 sg13g2_o21ai_1 _21953_ (.B1(_04055_),
    .Y(_01633_),
    .A1(net167),
    .A2(_04054_));
 sg13g2_nand2_1 _21954_ (.Y(_04056_),
    .A(net837),
    .B(\mem.mem_internal.code_mem[40][0] ));
 sg13g2_nor2_1 _21955_ (.A(net778),
    .B(net458),
    .Y(_04057_));
 sg13g2_buf_2 _21956_ (.A(_04057_),
    .X(_04058_));
 sg13g2_buf_1 _21957_ (.A(_04058_),
    .X(_04059_));
 sg13g2_buf_1 _21958_ (.A(_03842_),
    .X(_04060_));
 sg13g2_nand2_1 _21959_ (.Y(_04061_),
    .A(_04060_),
    .B(net166));
 sg13g2_o21ai_1 _21960_ (.B1(_04061_),
    .Y(_01634_),
    .A1(_04056_),
    .A2(net166));
 sg13g2_nand2_1 _21961_ (.Y(_04062_),
    .A(net641),
    .B(\mem.mem_internal.code_mem[40][1] ));
 sg13g2_buf_1 _21962_ (.A(_03846_),
    .X(_04063_));
 sg13g2_nand2_1 _21963_ (.Y(_04064_),
    .A(_04063_),
    .B(net166));
 sg13g2_o21ai_1 _21964_ (.B1(_04064_),
    .Y(_01635_),
    .A1(net166),
    .A2(_04062_));
 sg13g2_nand2_1 _21965_ (.Y(_04065_),
    .A(net641),
    .B(\mem.mem_internal.code_mem[40][2] ));
 sg13g2_buf_1 _21966_ (.A(_03850_),
    .X(_04066_));
 sg13g2_nand2_1 _21967_ (.Y(_04067_),
    .A(net1036),
    .B(_04058_));
 sg13g2_o21ai_1 _21968_ (.B1(_04067_),
    .Y(_01636_),
    .A1(net166),
    .A2(_04065_));
 sg13g2_nand2_1 _21969_ (.Y(_04068_),
    .A(net641),
    .B(\mem.mem_internal.code_mem[40][3] ));
 sg13g2_buf_1 _21970_ (.A(_03854_),
    .X(_04069_));
 sg13g2_nand2_1 _21971_ (.Y(_04070_),
    .A(net1035),
    .B(_04058_));
 sg13g2_o21ai_1 _21972_ (.B1(_04070_),
    .Y(_01637_),
    .A1(net166),
    .A2(_04068_));
 sg13g2_buf_1 _21973_ (.A(_04040_),
    .X(_04071_));
 sg13g2_nand2_1 _21974_ (.Y(_04072_),
    .A(net640),
    .B(\mem.mem_internal.code_mem[40][4] ));
 sg13g2_buf_1 _21975_ (.A(_03859_),
    .X(_04073_));
 sg13g2_nand2_1 _21976_ (.Y(_04074_),
    .A(net1034),
    .B(_04058_));
 sg13g2_o21ai_1 _21977_ (.B1(_04074_),
    .Y(_01638_),
    .A1(_04059_),
    .A2(_04072_));
 sg13g2_nand2_1 _21978_ (.Y(_04075_),
    .A(net640),
    .B(\mem.mem_internal.code_mem[40][5] ));
 sg13g2_buf_1 _21979_ (.A(_03863_),
    .X(_04076_));
 sg13g2_nand2_1 _21980_ (.Y(_04077_),
    .A(net1033),
    .B(_04058_));
 sg13g2_o21ai_1 _21981_ (.B1(_04077_),
    .Y(_01639_),
    .A1(_04059_),
    .A2(_04075_));
 sg13g2_nand2_1 _21982_ (.Y(_04078_),
    .A(net640),
    .B(\mem.mem_internal.code_mem[40][6] ));
 sg13g2_buf_1 _21983_ (.A(_03867_),
    .X(_04079_));
 sg13g2_nand2_1 _21984_ (.Y(_04080_),
    .A(net1032),
    .B(_04058_));
 sg13g2_o21ai_1 _21985_ (.B1(_04080_),
    .Y(_01640_),
    .A1(net166),
    .A2(_04078_));
 sg13g2_nand2_1 _21986_ (.Y(_04081_),
    .A(net640),
    .B(\mem.mem_internal.code_mem[40][7] ));
 sg13g2_buf_1 _21987_ (.A(_03871_),
    .X(_04082_));
 sg13g2_nand2_1 _21988_ (.Y(_04083_),
    .A(net1031),
    .B(_04058_));
 sg13g2_o21ai_1 _21989_ (.B1(_04083_),
    .Y(_01641_),
    .A1(net166),
    .A2(_04081_));
 sg13g2_nand2_1 _21990_ (.Y(_04084_),
    .A(net837),
    .B(\mem.mem_internal.code_mem[41][0] ));
 sg13g2_nor2_1 _21991_ (.A(_10422_),
    .B(net458),
    .Y(_04085_));
 sg13g2_buf_2 _21992_ (.A(_04085_),
    .X(_04086_));
 sg13g2_buf_1 _21993_ (.A(_04086_),
    .X(_04087_));
 sg13g2_nand2_1 _21994_ (.Y(_04088_),
    .A(net1038),
    .B(net165));
 sg13g2_o21ai_1 _21995_ (.B1(_04088_),
    .Y(_01642_),
    .A1(_04084_),
    .A2(net165));
 sg13g2_nand2_1 _21996_ (.Y(_04089_),
    .A(_04071_),
    .B(\mem.mem_internal.code_mem[41][1] ));
 sg13g2_nand2_1 _21997_ (.Y(_04090_),
    .A(net1037),
    .B(net165));
 sg13g2_o21ai_1 _21998_ (.B1(_04090_),
    .Y(_01643_),
    .A1(net165),
    .A2(_04089_));
 sg13g2_nand2_1 _21999_ (.Y(_04091_),
    .A(net640),
    .B(\mem.mem_internal.code_mem[41][2] ));
 sg13g2_nand2_1 _22000_ (.Y(_04092_),
    .A(net1036),
    .B(_04086_));
 sg13g2_o21ai_1 _22001_ (.B1(_04092_),
    .Y(_01644_),
    .A1(net165),
    .A2(_04091_));
 sg13g2_nand2_1 _22002_ (.Y(_04093_),
    .A(net640),
    .B(\mem.mem_internal.code_mem[41][3] ));
 sg13g2_nand2_1 _22003_ (.Y(_04094_),
    .A(_04069_),
    .B(_04086_));
 sg13g2_o21ai_1 _22004_ (.B1(_04094_),
    .Y(_01645_),
    .A1(net165),
    .A2(_04093_));
 sg13g2_nand2_1 _22005_ (.Y(_04095_),
    .A(_04071_),
    .B(\mem.mem_internal.code_mem[41][4] ));
 sg13g2_nand2_1 _22006_ (.Y(_04096_),
    .A(net1034),
    .B(_04086_));
 sg13g2_o21ai_1 _22007_ (.B1(_04096_),
    .Y(_01646_),
    .A1(_04087_),
    .A2(_04095_));
 sg13g2_nand2_1 _22008_ (.Y(_04097_),
    .A(net640),
    .B(\mem.mem_internal.code_mem[41][5] ));
 sg13g2_nand2_1 _22009_ (.Y(_04098_),
    .A(net1033),
    .B(_04086_));
 sg13g2_o21ai_1 _22010_ (.B1(_04098_),
    .Y(_01647_),
    .A1(_04087_),
    .A2(_04097_));
 sg13g2_nand2_1 _22011_ (.Y(_04099_),
    .A(net640),
    .B(\mem.mem_internal.code_mem[41][6] ));
 sg13g2_nand2_1 _22012_ (.Y(_04100_),
    .A(net1032),
    .B(_04086_));
 sg13g2_o21ai_1 _22013_ (.B1(_04100_),
    .Y(_01648_),
    .A1(net165),
    .A2(_04099_));
 sg13g2_buf_1 _22014_ (.A(_04040_),
    .X(_04101_));
 sg13g2_nand2_1 _22015_ (.Y(_04102_),
    .A(net639),
    .B(\mem.mem_internal.code_mem[41][7] ));
 sg13g2_nand2_1 _22016_ (.Y(_04103_),
    .A(net1031),
    .B(_04086_));
 sg13g2_o21ai_1 _22017_ (.B1(_04103_),
    .Y(_01649_),
    .A1(net165),
    .A2(_04102_));
 sg13g2_nand2_1 _22018_ (.Y(_04104_),
    .A(net837),
    .B(\mem.mem_internal.code_mem[42][0] ));
 sg13g2_nor2_1 _22019_ (.A(_10444_),
    .B(_03876_),
    .Y(_04105_));
 sg13g2_buf_2 _22020_ (.A(_04105_),
    .X(_04106_));
 sg13g2_buf_1 _22021_ (.A(_04106_),
    .X(_04107_));
 sg13g2_nand2_1 _22022_ (.Y(_04108_),
    .A(net1038),
    .B(net336));
 sg13g2_o21ai_1 _22023_ (.B1(_04108_),
    .Y(_01650_),
    .A1(_04104_),
    .A2(net336));
 sg13g2_nand2_1 _22024_ (.Y(_04109_),
    .A(net639),
    .B(\mem.mem_internal.code_mem[42][1] ));
 sg13g2_nand2_1 _22025_ (.Y(_04110_),
    .A(net1037),
    .B(net336));
 sg13g2_o21ai_1 _22026_ (.B1(_04110_),
    .Y(_01651_),
    .A1(net336),
    .A2(_04109_));
 sg13g2_nand2_1 _22027_ (.Y(_04111_),
    .A(_04101_),
    .B(\mem.mem_internal.code_mem[42][2] ));
 sg13g2_nand2_1 _22028_ (.Y(_04112_),
    .A(_04066_),
    .B(_04106_));
 sg13g2_o21ai_1 _22029_ (.B1(_04112_),
    .Y(_01652_),
    .A1(net336),
    .A2(_04111_));
 sg13g2_nand2_1 _22030_ (.Y(_04113_),
    .A(net639),
    .B(\mem.mem_internal.code_mem[42][3] ));
 sg13g2_nand2_1 _22031_ (.Y(_04114_),
    .A(_04069_),
    .B(_04106_));
 sg13g2_o21ai_1 _22032_ (.B1(_04114_),
    .Y(_01653_),
    .A1(_04107_),
    .A2(_04113_));
 sg13g2_nand2_1 _22033_ (.Y(_04115_),
    .A(net639),
    .B(\mem.mem_internal.code_mem[42][4] ));
 sg13g2_nand2_1 _22034_ (.Y(_04116_),
    .A(_04073_),
    .B(_04106_));
 sg13g2_o21ai_1 _22035_ (.B1(_04116_),
    .Y(_01654_),
    .A1(_04107_),
    .A2(_04115_));
 sg13g2_nand2_1 _22036_ (.Y(_04117_),
    .A(net639),
    .B(\mem.mem_internal.code_mem[42][5] ));
 sg13g2_nand2_1 _22037_ (.Y(_04118_),
    .A(_04076_),
    .B(_04106_));
 sg13g2_o21ai_1 _22038_ (.B1(_04118_),
    .Y(_01655_),
    .A1(net336),
    .A2(_04117_));
 sg13g2_nand2_1 _22039_ (.Y(_04119_),
    .A(net639),
    .B(\mem.mem_internal.code_mem[42][6] ));
 sg13g2_nand2_1 _22040_ (.Y(_04120_),
    .A(_04079_),
    .B(_04106_));
 sg13g2_o21ai_1 _22041_ (.B1(_04120_),
    .Y(_01656_),
    .A1(net336),
    .A2(_04119_));
 sg13g2_nand2_1 _22042_ (.Y(_04121_),
    .A(net639),
    .B(\mem.mem_internal.code_mem[42][7] ));
 sg13g2_nand2_1 _22043_ (.Y(_04122_),
    .A(_04082_),
    .B(_04106_));
 sg13g2_o21ai_1 _22044_ (.B1(_04122_),
    .Y(_01657_),
    .A1(net336),
    .A2(_04121_));
 sg13g2_nand2_1 _22045_ (.Y(_04123_),
    .A(net837),
    .B(\mem.mem_internal.code_mem[43][0] ));
 sg13g2_nor2_1 _22046_ (.A(net775),
    .B(_03876_),
    .Y(_04124_));
 sg13g2_buf_2 _22047_ (.A(_04124_),
    .X(_04125_));
 sg13g2_buf_1 _22048_ (.A(_04125_),
    .X(_04126_));
 sg13g2_nand2_1 _22049_ (.Y(_04127_),
    .A(_04060_),
    .B(net335));
 sg13g2_o21ai_1 _22050_ (.B1(_04127_),
    .Y(_01658_),
    .A1(_04123_),
    .A2(net335));
 sg13g2_nand2_1 _22051_ (.Y(_04128_),
    .A(net639),
    .B(\mem.mem_internal.code_mem[43][1] ));
 sg13g2_nand2_1 _22052_ (.Y(_04129_),
    .A(_04063_),
    .B(net335));
 sg13g2_o21ai_1 _22053_ (.B1(_04129_),
    .Y(_01659_),
    .A1(net335),
    .A2(_04128_));
 sg13g2_nand2_1 _22054_ (.Y(_04130_),
    .A(_04101_),
    .B(\mem.mem_internal.code_mem[43][2] ));
 sg13g2_nand2_1 _22055_ (.Y(_04131_),
    .A(_04066_),
    .B(_04125_));
 sg13g2_o21ai_1 _22056_ (.B1(_04131_),
    .Y(_01660_),
    .A1(net335),
    .A2(_04130_));
 sg13g2_buf_1 _22057_ (.A(_04040_),
    .X(_04132_));
 sg13g2_nand2_1 _22058_ (.Y(_04133_),
    .A(net638),
    .B(\mem.mem_internal.code_mem[43][3] ));
 sg13g2_nand2_1 _22059_ (.Y(_04134_),
    .A(net1035),
    .B(_04125_));
 sg13g2_o21ai_1 _22060_ (.B1(_04134_),
    .Y(_01661_),
    .A1(_04126_),
    .A2(_04133_));
 sg13g2_nand2_1 _22061_ (.Y(_04135_),
    .A(net638),
    .B(\mem.mem_internal.code_mem[43][4] ));
 sg13g2_nand2_1 _22062_ (.Y(_04136_),
    .A(_04073_),
    .B(_04125_));
 sg13g2_o21ai_1 _22063_ (.B1(_04136_),
    .Y(_01662_),
    .A1(_04126_),
    .A2(_04135_));
 sg13g2_nand2_1 _22064_ (.Y(_04137_),
    .A(net638),
    .B(\mem.mem_internal.code_mem[43][5] ));
 sg13g2_nand2_1 _22065_ (.Y(_04138_),
    .A(_04076_),
    .B(_04125_));
 sg13g2_o21ai_1 _22066_ (.B1(_04138_),
    .Y(_01663_),
    .A1(net335),
    .A2(_04137_));
 sg13g2_nand2_1 _22067_ (.Y(_04139_),
    .A(_04132_),
    .B(\mem.mem_internal.code_mem[43][6] ));
 sg13g2_nand2_1 _22068_ (.Y(_04140_),
    .A(_04079_),
    .B(_04125_));
 sg13g2_o21ai_1 _22069_ (.B1(_04140_),
    .Y(_01664_),
    .A1(net335),
    .A2(_04139_));
 sg13g2_nand2_1 _22070_ (.Y(_04141_),
    .A(_04132_),
    .B(\mem.mem_internal.code_mem[43][7] ));
 sg13g2_nand2_1 _22071_ (.Y(_04142_),
    .A(_04082_),
    .B(_04125_));
 sg13g2_o21ai_1 _22072_ (.B1(_04142_),
    .Y(_01665_),
    .A1(net335),
    .A2(_04141_));
 sg13g2_nand2_1 _22073_ (.Y(_04143_),
    .A(net837),
    .B(\mem.mem_internal.code_mem[44][0] ));
 sg13g2_nor2_1 _22074_ (.A(_10491_),
    .B(_03876_),
    .Y(_04144_));
 sg13g2_buf_2 _22075_ (.A(_04144_),
    .X(_04145_));
 sg13g2_buf_1 _22076_ (.A(_04145_),
    .X(_04146_));
 sg13g2_nand2_1 _22077_ (.Y(_04147_),
    .A(net1038),
    .B(net334));
 sg13g2_o21ai_1 _22078_ (.B1(_04147_),
    .Y(_01666_),
    .A1(_04143_),
    .A2(net334));
 sg13g2_nand2_1 _22079_ (.Y(_04148_),
    .A(net638),
    .B(\mem.mem_internal.code_mem[44][1] ));
 sg13g2_nand2_1 _22080_ (.Y(_04149_),
    .A(net1037),
    .B(net334));
 sg13g2_o21ai_1 _22081_ (.B1(_04149_),
    .Y(_01667_),
    .A1(net334),
    .A2(_04148_));
 sg13g2_nand2_1 _22082_ (.Y(_04150_),
    .A(net638),
    .B(\mem.mem_internal.code_mem[44][2] ));
 sg13g2_nand2_1 _22083_ (.Y(_04151_),
    .A(net1036),
    .B(_04145_));
 sg13g2_o21ai_1 _22084_ (.B1(_04151_),
    .Y(_01668_),
    .A1(_04146_),
    .A2(_04150_));
 sg13g2_nand2_1 _22085_ (.Y(_04152_),
    .A(net638),
    .B(\mem.mem_internal.code_mem[44][3] ));
 sg13g2_nand2_1 _22086_ (.Y(_04153_),
    .A(net1035),
    .B(_04145_));
 sg13g2_o21ai_1 _22087_ (.B1(_04153_),
    .Y(_01669_),
    .A1(net334),
    .A2(_04152_));
 sg13g2_nand2_1 _22088_ (.Y(_04154_),
    .A(net638),
    .B(\mem.mem_internal.code_mem[44][4] ));
 sg13g2_nand2_1 _22089_ (.Y(_04155_),
    .A(net1034),
    .B(_04145_));
 sg13g2_o21ai_1 _22090_ (.B1(_04155_),
    .Y(_01670_),
    .A1(_04146_),
    .A2(_04154_));
 sg13g2_nand2_1 _22091_ (.Y(_04156_),
    .A(net638),
    .B(\mem.mem_internal.code_mem[44][5] ));
 sg13g2_nand2_1 _22092_ (.Y(_04157_),
    .A(net1033),
    .B(_04145_));
 sg13g2_o21ai_1 _22093_ (.B1(_04157_),
    .Y(_01671_),
    .A1(net334),
    .A2(_04156_));
 sg13g2_buf_1 _22094_ (.A(_04040_),
    .X(_04158_));
 sg13g2_nand2_1 _22095_ (.Y(_04159_),
    .A(net637),
    .B(\mem.mem_internal.code_mem[44][6] ));
 sg13g2_nand2_1 _22096_ (.Y(_04160_),
    .A(net1032),
    .B(_04145_));
 sg13g2_o21ai_1 _22097_ (.B1(_04160_),
    .Y(_01672_),
    .A1(net334),
    .A2(_04159_));
 sg13g2_nand2_1 _22098_ (.Y(_04161_),
    .A(net637),
    .B(\mem.mem_internal.code_mem[44][7] ));
 sg13g2_nand2_1 _22099_ (.Y(_04162_),
    .A(net1031),
    .B(_04145_));
 sg13g2_o21ai_1 _22100_ (.B1(_04162_),
    .Y(_01673_),
    .A1(net334),
    .A2(_04161_));
 sg13g2_nand2_1 _22101_ (.Y(_04163_),
    .A(net837),
    .B(\mem.mem_internal.code_mem[45][0] ));
 sg13g2_nor2_1 _22102_ (.A(_10513_),
    .B(_03876_),
    .Y(_04164_));
 sg13g2_buf_2 _22103_ (.A(_04164_),
    .X(_04165_));
 sg13g2_buf_1 _22104_ (.A(_04165_),
    .X(_04166_));
 sg13g2_nand2_1 _22105_ (.Y(_04167_),
    .A(net1038),
    .B(net333));
 sg13g2_o21ai_1 _22106_ (.B1(_04167_),
    .Y(_01674_),
    .A1(_04163_),
    .A2(net333));
 sg13g2_nand2_1 _22107_ (.Y(_04168_),
    .A(net637),
    .B(\mem.mem_internal.code_mem[45][1] ));
 sg13g2_nand2_1 _22108_ (.Y(_04169_),
    .A(net1037),
    .B(net333));
 sg13g2_o21ai_1 _22109_ (.B1(_04169_),
    .Y(_01675_),
    .A1(net333),
    .A2(_04168_));
 sg13g2_nand2_1 _22110_ (.Y(_04170_),
    .A(net637),
    .B(\mem.mem_internal.code_mem[45][2] ));
 sg13g2_nand2_1 _22111_ (.Y(_04171_),
    .A(net1036),
    .B(_04165_));
 sg13g2_o21ai_1 _22112_ (.B1(_04171_),
    .Y(_01676_),
    .A1(net333),
    .A2(_04170_));
 sg13g2_nand2_1 _22113_ (.Y(_04172_),
    .A(net637),
    .B(\mem.mem_internal.code_mem[45][3] ));
 sg13g2_nand2_1 _22114_ (.Y(_04173_),
    .A(net1035),
    .B(_04165_));
 sg13g2_o21ai_1 _22115_ (.B1(_04173_),
    .Y(_01677_),
    .A1(net333),
    .A2(_04172_));
 sg13g2_nand2_1 _22116_ (.Y(_04174_),
    .A(_04158_),
    .B(\mem.mem_internal.code_mem[45][4] ));
 sg13g2_nand2_1 _22117_ (.Y(_04175_),
    .A(net1034),
    .B(_04165_));
 sg13g2_o21ai_1 _22118_ (.B1(_04175_),
    .Y(_01678_),
    .A1(net333),
    .A2(_04174_));
 sg13g2_nand2_1 _22119_ (.Y(_04176_),
    .A(_04158_),
    .B(\mem.mem_internal.code_mem[45][5] ));
 sg13g2_nand2_1 _22120_ (.Y(_04177_),
    .A(net1033),
    .B(_04165_));
 sg13g2_o21ai_1 _22121_ (.B1(_04177_),
    .Y(_01679_),
    .A1(_04166_),
    .A2(_04176_));
 sg13g2_nand2_1 _22122_ (.Y(_04178_),
    .A(net637),
    .B(\mem.mem_internal.code_mem[45][6] ));
 sg13g2_nand2_1 _22123_ (.Y(_04179_),
    .A(net1032),
    .B(_04165_));
 sg13g2_o21ai_1 _22124_ (.B1(_04179_),
    .Y(_01680_),
    .A1(net333),
    .A2(_04178_));
 sg13g2_nand2_1 _22125_ (.Y(_04180_),
    .A(net637),
    .B(\mem.mem_internal.code_mem[45][7] ));
 sg13g2_nand2_1 _22126_ (.Y(_04181_),
    .A(net1031),
    .B(_04165_));
 sg13g2_o21ai_1 _22127_ (.B1(_04181_),
    .Y(_01681_),
    .A1(_04166_),
    .A2(_04180_));
 sg13g2_nand2_1 _22128_ (.Y(_04182_),
    .A(net837),
    .B(\mem.mem_internal.code_mem[46][0] ));
 sg13g2_nor2_1 _22129_ (.A(_10564_),
    .B(_03876_),
    .Y(_04183_));
 sg13g2_buf_2 _22130_ (.A(_04183_),
    .X(_04184_));
 sg13g2_buf_1 _22131_ (.A(_04184_),
    .X(_04185_));
 sg13g2_nand2_1 _22132_ (.Y(_04186_),
    .A(net1038),
    .B(net332));
 sg13g2_o21ai_1 _22133_ (.B1(_04186_),
    .Y(_01682_),
    .A1(_04182_),
    .A2(_04185_));
 sg13g2_nand2_1 _22134_ (.Y(_04187_),
    .A(net637),
    .B(\mem.mem_internal.code_mem[46][1] ));
 sg13g2_nand2_1 _22135_ (.Y(_04188_),
    .A(net1037),
    .B(net332));
 sg13g2_o21ai_1 _22136_ (.B1(_04188_),
    .Y(_01683_),
    .A1(net332),
    .A2(_04187_));
 sg13g2_buf_1 _22137_ (.A(_04040_),
    .X(_04189_));
 sg13g2_nand2_1 _22138_ (.Y(_04190_),
    .A(net636),
    .B(\mem.mem_internal.code_mem[46][2] ));
 sg13g2_nand2_1 _22139_ (.Y(_04191_),
    .A(net1036),
    .B(_04184_));
 sg13g2_o21ai_1 _22140_ (.B1(_04191_),
    .Y(_01684_),
    .A1(net332),
    .A2(_04190_));
 sg13g2_nand2_1 _22141_ (.Y(_04192_),
    .A(net636),
    .B(\mem.mem_internal.code_mem[46][3] ));
 sg13g2_nand2_1 _22142_ (.Y(_04193_),
    .A(net1035),
    .B(_04184_));
 sg13g2_o21ai_1 _22143_ (.B1(_04193_),
    .Y(_01685_),
    .A1(net332),
    .A2(_04192_));
 sg13g2_nand2_1 _22144_ (.Y(_04194_),
    .A(_04189_),
    .B(\mem.mem_internal.code_mem[46][4] ));
 sg13g2_nand2_1 _22145_ (.Y(_04195_),
    .A(net1034),
    .B(_04184_));
 sg13g2_o21ai_1 _22146_ (.B1(_04195_),
    .Y(_01686_),
    .A1(net332),
    .A2(_04194_));
 sg13g2_nand2_1 _22147_ (.Y(_04196_),
    .A(net636),
    .B(\mem.mem_internal.code_mem[46][5] ));
 sg13g2_nand2_1 _22148_ (.Y(_04197_),
    .A(net1033),
    .B(_04184_));
 sg13g2_o21ai_1 _22149_ (.B1(_04197_),
    .Y(_01687_),
    .A1(net332),
    .A2(_04196_));
 sg13g2_nand2_1 _22150_ (.Y(_04198_),
    .A(net636),
    .B(\mem.mem_internal.code_mem[46][6] ));
 sg13g2_nand2_1 _22151_ (.Y(_04199_),
    .A(net1032),
    .B(_04184_));
 sg13g2_o21ai_1 _22152_ (.B1(_04199_),
    .Y(_01688_),
    .A1(net332),
    .A2(_04198_));
 sg13g2_nand2_1 _22153_ (.Y(_04200_),
    .A(net636),
    .B(\mem.mem_internal.code_mem[46][7] ));
 sg13g2_nand2_1 _22154_ (.Y(_04201_),
    .A(net1031),
    .B(_04184_));
 sg13g2_o21ai_1 _22155_ (.B1(_04201_),
    .Y(_01689_),
    .A1(_04185_),
    .A2(_04200_));
 sg13g2_buf_1 _22156_ (.A(_12878_),
    .X(_04202_));
 sg13g2_nand2_1 _22157_ (.Y(_04203_),
    .A(_04202_),
    .B(\mem.mem_internal.code_mem[47][0] ));
 sg13g2_nor2_1 _22158_ (.A(_10586_),
    .B(_03876_),
    .Y(_04204_));
 sg13g2_buf_2 _22159_ (.A(_04204_),
    .X(_04205_));
 sg13g2_buf_1 _22160_ (.A(_04205_),
    .X(_04206_));
 sg13g2_nand2_1 _22161_ (.Y(_04207_),
    .A(net1038),
    .B(_04206_));
 sg13g2_o21ai_1 _22162_ (.B1(_04207_),
    .Y(_01690_),
    .A1(_04203_),
    .A2(_04206_));
 sg13g2_nand2_1 _22163_ (.Y(_04208_),
    .A(net636),
    .B(\mem.mem_internal.code_mem[47][1] ));
 sg13g2_nand2_1 _22164_ (.Y(_04209_),
    .A(net1037),
    .B(net331));
 sg13g2_o21ai_1 _22165_ (.B1(_04209_),
    .Y(_01691_),
    .A1(net331),
    .A2(_04208_));
 sg13g2_nand2_1 _22166_ (.Y(_04210_),
    .A(net636),
    .B(\mem.mem_internal.code_mem[47][2] ));
 sg13g2_nand2_1 _22167_ (.Y(_04211_),
    .A(net1036),
    .B(_04205_));
 sg13g2_o21ai_1 _22168_ (.B1(_04211_),
    .Y(_01692_),
    .A1(net331),
    .A2(_04210_));
 sg13g2_nand2_1 _22169_ (.Y(_04212_),
    .A(net636),
    .B(\mem.mem_internal.code_mem[47][3] ));
 sg13g2_nand2_1 _22170_ (.Y(_04213_),
    .A(net1035),
    .B(_04205_));
 sg13g2_o21ai_1 _22171_ (.B1(_04213_),
    .Y(_01693_),
    .A1(net331),
    .A2(_04212_));
 sg13g2_nand2_1 _22172_ (.Y(_04214_),
    .A(_04189_),
    .B(\mem.mem_internal.code_mem[47][4] ));
 sg13g2_nand2_1 _22173_ (.Y(_04215_),
    .A(net1034),
    .B(_04205_));
 sg13g2_o21ai_1 _22174_ (.B1(_04215_),
    .Y(_01694_),
    .A1(net331),
    .A2(_04214_));
 sg13g2_buf_1 _22175_ (.A(_04040_),
    .X(_04216_));
 sg13g2_nand2_1 _22176_ (.Y(_04217_),
    .A(net635),
    .B(\mem.mem_internal.code_mem[47][5] ));
 sg13g2_nand2_1 _22177_ (.Y(_04218_),
    .A(net1033),
    .B(_04205_));
 sg13g2_o21ai_1 _22178_ (.B1(_04218_),
    .Y(_01695_),
    .A1(net331),
    .A2(_04217_));
 sg13g2_nand2_1 _22179_ (.Y(_04219_),
    .A(net635),
    .B(\mem.mem_internal.code_mem[47][6] ));
 sg13g2_nand2_1 _22180_ (.Y(_04220_),
    .A(net1032),
    .B(_04205_));
 sg13g2_o21ai_1 _22181_ (.B1(_04220_),
    .Y(_01696_),
    .A1(net331),
    .A2(_04219_));
 sg13g2_nand2_1 _22182_ (.Y(_04221_),
    .A(net635),
    .B(\mem.mem_internal.code_mem[47][7] ));
 sg13g2_nand2_1 _22183_ (.Y(_04222_),
    .A(net1031),
    .B(_04205_));
 sg13g2_o21ai_1 _22184_ (.B1(_04222_),
    .Y(_01697_),
    .A1(net331),
    .A2(_04221_));
 sg13g2_nand3_1 _22185_ (.B(_10034_),
    .C(_10234_),
    .A(_10113_),
    .Y(_04223_));
 sg13g2_buf_2 _22186_ (.A(_04223_),
    .X(_04224_));
 sg13g2_inv_1 _22187_ (.Y(_04225_),
    .A(_04224_));
 sg13g2_nand2b_1 _22188_ (.Y(_04226_),
    .B(_04225_),
    .A_N(_10243_));
 sg13g2_buf_1 _22189_ (.A(_04226_),
    .X(_04227_));
 sg13g2_buf_1 _22190_ (.A(_04227_),
    .X(_04228_));
 sg13g2_nor2_1 _22191_ (.A(net529),
    .B(net482),
    .Y(_04229_));
 sg13g2_buf_2 _22192_ (.A(_04229_),
    .X(_04230_));
 sg13g2_buf_1 _22193_ (.A(_04230_),
    .X(_04231_));
 sg13g2_nand2_1 _22194_ (.Y(_04232_),
    .A(_04216_),
    .B(\mem.mem_internal.code_mem[48][0] ));
 sg13g2_nand2_1 _22195_ (.Y(_04233_),
    .A(net1038),
    .B(_04231_));
 sg13g2_o21ai_1 _22196_ (.B1(_04233_),
    .Y(_01698_),
    .A1(_04231_),
    .A2(_04232_));
 sg13g2_nand2_1 _22197_ (.Y(_04234_),
    .A(net635),
    .B(\mem.mem_internal.code_mem[48][1] ));
 sg13g2_nand2_1 _22198_ (.Y(_04235_),
    .A(net1037),
    .B(net330));
 sg13g2_o21ai_1 _22199_ (.B1(_04235_),
    .Y(_01699_),
    .A1(net330),
    .A2(_04234_));
 sg13g2_nand2_1 _22200_ (.Y(_04236_),
    .A(_04216_),
    .B(\mem.mem_internal.code_mem[48][2] ));
 sg13g2_nand2_1 _22201_ (.Y(_04237_),
    .A(net1036),
    .B(_04230_));
 sg13g2_o21ai_1 _22202_ (.B1(_04237_),
    .Y(_01700_),
    .A1(net330),
    .A2(_04236_));
 sg13g2_nand2_1 _22203_ (.Y(_04238_),
    .A(net635),
    .B(\mem.mem_internal.code_mem[48][3] ));
 sg13g2_nand2_1 _22204_ (.Y(_04239_),
    .A(net1035),
    .B(_04230_));
 sg13g2_o21ai_1 _22205_ (.B1(_04239_),
    .Y(_01701_),
    .A1(net330),
    .A2(_04238_));
 sg13g2_nand2_1 _22206_ (.Y(_04240_),
    .A(net635),
    .B(\mem.mem_internal.code_mem[48][4] ));
 sg13g2_nand2_1 _22207_ (.Y(_04241_),
    .A(net1034),
    .B(_04230_));
 sg13g2_o21ai_1 _22208_ (.B1(_04241_),
    .Y(_01702_),
    .A1(net330),
    .A2(_04240_));
 sg13g2_nand2_1 _22209_ (.Y(_04242_),
    .A(net635),
    .B(\mem.mem_internal.code_mem[48][5] ));
 sg13g2_nand2_1 _22210_ (.Y(_04243_),
    .A(net1033),
    .B(_04230_));
 sg13g2_o21ai_1 _22211_ (.B1(_04243_),
    .Y(_01703_),
    .A1(net330),
    .A2(_04242_));
 sg13g2_nand2_1 _22212_ (.Y(_04244_),
    .A(net635),
    .B(\mem.mem_internal.code_mem[48][6] ));
 sg13g2_nand2_1 _22213_ (.Y(_04245_),
    .A(net1032),
    .B(_04230_));
 sg13g2_o21ai_1 _22214_ (.B1(_04245_),
    .Y(_01704_),
    .A1(net330),
    .A2(_04244_));
 sg13g2_buf_1 _22215_ (.A(_03042_),
    .X(_04246_));
 sg13g2_buf_1 _22216_ (.A(_04246_),
    .X(_04247_));
 sg13g2_nand2_1 _22217_ (.Y(_04248_),
    .A(net634),
    .B(\mem.mem_internal.code_mem[48][7] ));
 sg13g2_nand2_1 _22218_ (.Y(_04249_),
    .A(net1031),
    .B(_04230_));
 sg13g2_o21ai_1 _22219_ (.B1(_04249_),
    .Y(_01705_),
    .A1(net330),
    .A2(_04248_));
 sg13g2_nor2_1 _22220_ (.A(net528),
    .B(net482),
    .Y(_04250_));
 sg13g2_buf_2 _22221_ (.A(_04250_),
    .X(_04251_));
 sg13g2_buf_1 _22222_ (.A(_04251_),
    .X(_04252_));
 sg13g2_nand2_1 _22223_ (.Y(_04253_),
    .A(_04247_),
    .B(\mem.mem_internal.code_mem[49][0] ));
 sg13g2_nand2_1 _22224_ (.Y(_04254_),
    .A(net1038),
    .B(_04252_));
 sg13g2_o21ai_1 _22225_ (.B1(_04254_),
    .Y(_01706_),
    .A1(_04252_),
    .A2(_04253_));
 sg13g2_nand2_1 _22226_ (.Y(_04255_),
    .A(net634),
    .B(\mem.mem_internal.code_mem[49][1] ));
 sg13g2_nand2_1 _22227_ (.Y(_04256_),
    .A(net1037),
    .B(net329));
 sg13g2_o21ai_1 _22228_ (.B1(_04256_),
    .Y(_01707_),
    .A1(net329),
    .A2(_04255_));
 sg13g2_nand2_1 _22229_ (.Y(_04257_),
    .A(net634),
    .B(\mem.mem_internal.code_mem[49][2] ));
 sg13g2_nand2_1 _22230_ (.Y(_04258_),
    .A(net1036),
    .B(_04251_));
 sg13g2_o21ai_1 _22231_ (.B1(_04258_),
    .Y(_01708_),
    .A1(net329),
    .A2(_04257_));
 sg13g2_nand2_1 _22232_ (.Y(_04259_),
    .A(net634),
    .B(\mem.mem_internal.code_mem[49][3] ));
 sg13g2_nand2_1 _22233_ (.Y(_04260_),
    .A(net1035),
    .B(_04251_));
 sg13g2_o21ai_1 _22234_ (.B1(_04260_),
    .Y(_01709_),
    .A1(net329),
    .A2(_04259_));
 sg13g2_nand2_1 _22235_ (.Y(_04261_),
    .A(net634),
    .B(\mem.mem_internal.code_mem[49][4] ));
 sg13g2_nand2_1 _22236_ (.Y(_04262_),
    .A(net1034),
    .B(_04251_));
 sg13g2_o21ai_1 _22237_ (.B1(_04262_),
    .Y(_01710_),
    .A1(net329),
    .A2(_04261_));
 sg13g2_nand2_1 _22238_ (.Y(_04263_),
    .A(net634),
    .B(\mem.mem_internal.code_mem[49][5] ));
 sg13g2_nand2_1 _22239_ (.Y(_04264_),
    .A(net1033),
    .B(_04251_));
 sg13g2_o21ai_1 _22240_ (.B1(_04264_),
    .Y(_01711_),
    .A1(net329),
    .A2(_04263_));
 sg13g2_nand2_1 _22241_ (.Y(_04265_),
    .A(net634),
    .B(\mem.mem_internal.code_mem[49][6] ));
 sg13g2_nand2_1 _22242_ (.Y(_04266_),
    .A(net1032),
    .B(_04251_));
 sg13g2_o21ai_1 _22243_ (.B1(_04266_),
    .Y(_01712_),
    .A1(net329),
    .A2(_04265_));
 sg13g2_nand2_1 _22244_ (.Y(_04267_),
    .A(net634),
    .B(\mem.mem_internal.code_mem[49][7] ));
 sg13g2_nand2_1 _22245_ (.Y(_04268_),
    .A(net1031),
    .B(_04251_));
 sg13g2_o21ai_1 _22246_ (.B1(_04268_),
    .Y(_01713_),
    .A1(net329),
    .A2(_04267_));
 sg13g2_nand2_1 _22247_ (.Y(_04269_),
    .A(net836),
    .B(\mem.mem_internal.code_mem[4][0] ));
 sg13g2_nor2_1 _22248_ (.A(_10246_),
    .B(net556),
    .Y(_04270_));
 sg13g2_buf_2 _22249_ (.A(_04270_),
    .X(_04271_));
 sg13g2_buf_1 _22250_ (.A(_04271_),
    .X(_04272_));
 sg13g2_buf_1 _22251_ (.A(_03842_),
    .X(_04273_));
 sg13g2_nand2_1 _22252_ (.Y(_04274_),
    .A(_04273_),
    .B(net328));
 sg13g2_o21ai_1 _22253_ (.B1(_04274_),
    .Y(_01714_),
    .A1(_04269_),
    .A2(net328));
 sg13g2_nand2_1 _22254_ (.Y(_04275_),
    .A(_04247_),
    .B(\mem.mem_internal.code_mem[4][1] ));
 sg13g2_buf_1 _22255_ (.A(_03846_),
    .X(_04276_));
 sg13g2_nand2_1 _22256_ (.Y(_04277_),
    .A(_04276_),
    .B(net328));
 sg13g2_o21ai_1 _22257_ (.B1(_04277_),
    .Y(_01715_),
    .A1(net328),
    .A2(_04275_));
 sg13g2_buf_1 _22258_ (.A(_04246_),
    .X(_04278_));
 sg13g2_nand2_1 _22259_ (.Y(_04279_),
    .A(net633),
    .B(\mem.mem_internal.code_mem[4][2] ));
 sg13g2_buf_1 _22260_ (.A(_03850_),
    .X(_04280_));
 sg13g2_nand2_1 _22261_ (.Y(_04281_),
    .A(_04280_),
    .B(_04271_));
 sg13g2_o21ai_1 _22262_ (.B1(_04281_),
    .Y(_01716_),
    .A1(net328),
    .A2(_04279_));
 sg13g2_nand2_1 _22263_ (.Y(_04282_),
    .A(net633),
    .B(\mem.mem_internal.code_mem[4][3] ));
 sg13g2_buf_1 _22264_ (.A(_03854_),
    .X(_04283_));
 sg13g2_nand2_1 _22265_ (.Y(_04284_),
    .A(_04283_),
    .B(_04271_));
 sg13g2_o21ai_1 _22266_ (.B1(_04284_),
    .Y(_01717_),
    .A1(net328),
    .A2(_04282_));
 sg13g2_nand2_1 _22267_ (.Y(_04285_),
    .A(net633),
    .B(\mem.mem_internal.code_mem[4][4] ));
 sg13g2_buf_1 _22268_ (.A(_03859_),
    .X(_04286_));
 sg13g2_nand2_1 _22269_ (.Y(_04287_),
    .A(_04286_),
    .B(_04271_));
 sg13g2_o21ai_1 _22270_ (.B1(_04287_),
    .Y(_01718_),
    .A1(net328),
    .A2(_04285_));
 sg13g2_nand2_1 _22271_ (.Y(_04288_),
    .A(net633),
    .B(\mem.mem_internal.code_mem[4][5] ));
 sg13g2_buf_1 _22272_ (.A(_03863_),
    .X(_04289_));
 sg13g2_nand2_1 _22273_ (.Y(_04290_),
    .A(_04289_),
    .B(_04271_));
 sg13g2_o21ai_1 _22274_ (.B1(_04290_),
    .Y(_01719_),
    .A1(net328),
    .A2(_04288_));
 sg13g2_nand2_1 _22275_ (.Y(_04291_),
    .A(_04278_),
    .B(\mem.mem_internal.code_mem[4][6] ));
 sg13g2_buf_1 _22276_ (.A(_03867_),
    .X(_04292_));
 sg13g2_nand2_1 _22277_ (.Y(_04293_),
    .A(_04292_),
    .B(_04271_));
 sg13g2_o21ai_1 _22278_ (.B1(_04293_),
    .Y(_01720_),
    .A1(_04272_),
    .A2(_04291_));
 sg13g2_nand2_1 _22279_ (.Y(_04294_),
    .A(_04278_),
    .B(\mem.mem_internal.code_mem[4][7] ));
 sg13g2_buf_1 _22280_ (.A(_03871_),
    .X(_04295_));
 sg13g2_nand2_1 _22281_ (.Y(_04296_),
    .A(_04295_),
    .B(_04271_));
 sg13g2_o21ai_1 _22282_ (.B1(_04296_),
    .Y(_01721_),
    .A1(_04272_),
    .A2(_04294_));
 sg13g2_nor2_1 _22283_ (.A(net527),
    .B(net482),
    .Y(_04297_));
 sg13g2_buf_2 _22284_ (.A(_04297_),
    .X(_04298_));
 sg13g2_buf_1 _22285_ (.A(_04298_),
    .X(_04299_));
 sg13g2_nand2_1 _22286_ (.Y(_04300_),
    .A(net633),
    .B(\mem.mem_internal.code_mem[50][0] ));
 sg13g2_nand2_1 _22287_ (.Y(_04301_),
    .A(net1030),
    .B(_04299_));
 sg13g2_o21ai_1 _22288_ (.B1(_04301_),
    .Y(_01722_),
    .A1(_04299_),
    .A2(_04300_));
 sg13g2_nand2_1 _22289_ (.Y(_04302_),
    .A(net633),
    .B(\mem.mem_internal.code_mem[50][1] ));
 sg13g2_nand2_1 _22290_ (.Y(_04303_),
    .A(net1029),
    .B(net327));
 sg13g2_o21ai_1 _22291_ (.B1(_04303_),
    .Y(_01723_),
    .A1(net327),
    .A2(_04302_));
 sg13g2_nand2_1 _22292_ (.Y(_04304_),
    .A(net633),
    .B(\mem.mem_internal.code_mem[50][2] ));
 sg13g2_nand2_1 _22293_ (.Y(_04305_),
    .A(net1028),
    .B(_04298_));
 sg13g2_o21ai_1 _22294_ (.B1(_04305_),
    .Y(_01724_),
    .A1(net327),
    .A2(_04304_));
 sg13g2_nand2_1 _22295_ (.Y(_04306_),
    .A(net633),
    .B(\mem.mem_internal.code_mem[50][3] ));
 sg13g2_nand2_1 _22296_ (.Y(_04307_),
    .A(net1027),
    .B(_04298_));
 sg13g2_o21ai_1 _22297_ (.B1(_04307_),
    .Y(_01725_),
    .A1(net327),
    .A2(_04306_));
 sg13g2_buf_1 _22298_ (.A(_04246_),
    .X(_04308_));
 sg13g2_nand2_1 _22299_ (.Y(_04309_),
    .A(net632),
    .B(\mem.mem_internal.code_mem[50][4] ));
 sg13g2_nand2_1 _22300_ (.Y(_04310_),
    .A(net1026),
    .B(_04298_));
 sg13g2_o21ai_1 _22301_ (.B1(_04310_),
    .Y(_01726_),
    .A1(net327),
    .A2(_04309_));
 sg13g2_nand2_1 _22302_ (.Y(_04311_),
    .A(net632),
    .B(\mem.mem_internal.code_mem[50][5] ));
 sg13g2_nand2_1 _22303_ (.Y(_04312_),
    .A(net1025),
    .B(_04298_));
 sg13g2_o21ai_1 _22304_ (.B1(_04312_),
    .Y(_01727_),
    .A1(net327),
    .A2(_04311_));
 sg13g2_nand2_1 _22305_ (.Y(_04313_),
    .A(net632),
    .B(\mem.mem_internal.code_mem[50][6] ));
 sg13g2_nand2_1 _22306_ (.Y(_04314_),
    .A(net1024),
    .B(_04298_));
 sg13g2_o21ai_1 _22307_ (.B1(_04314_),
    .Y(_01728_),
    .A1(net327),
    .A2(_04313_));
 sg13g2_nand2_1 _22308_ (.Y(_04315_),
    .A(_04308_),
    .B(\mem.mem_internal.code_mem[50][7] ));
 sg13g2_nand2_1 _22309_ (.Y(_04316_),
    .A(net1023),
    .B(_04298_));
 sg13g2_o21ai_1 _22310_ (.B1(_04316_),
    .Y(_01729_),
    .A1(net327),
    .A2(_04315_));
 sg13g2_nor2_1 _22311_ (.A(net526),
    .B(net482),
    .Y(_04317_));
 sg13g2_buf_2 _22312_ (.A(_04317_),
    .X(_04318_));
 sg13g2_buf_1 _22313_ (.A(_04318_),
    .X(_04319_));
 sg13g2_nand2_1 _22314_ (.Y(_04320_),
    .A(net632),
    .B(\mem.mem_internal.code_mem[51][0] ));
 sg13g2_nand2_1 _22315_ (.Y(_04321_),
    .A(net1030),
    .B(net326));
 sg13g2_o21ai_1 _22316_ (.B1(_04321_),
    .Y(_01730_),
    .A1(net326),
    .A2(_04320_));
 sg13g2_nand2_1 _22317_ (.Y(_04322_),
    .A(net632),
    .B(\mem.mem_internal.code_mem[51][1] ));
 sg13g2_nand2_1 _22318_ (.Y(_04323_),
    .A(net1029),
    .B(net326));
 sg13g2_o21ai_1 _22319_ (.B1(_04323_),
    .Y(_01731_),
    .A1(net326),
    .A2(_04322_));
 sg13g2_nand2_1 _22320_ (.Y(_04324_),
    .A(_04308_),
    .B(\mem.mem_internal.code_mem[51][2] ));
 sg13g2_nand2_1 _22321_ (.Y(_04325_),
    .A(net1028),
    .B(_04318_));
 sg13g2_o21ai_1 _22322_ (.B1(_04325_),
    .Y(_01732_),
    .A1(_04319_),
    .A2(_04324_));
 sg13g2_nand2_1 _22323_ (.Y(_04326_),
    .A(net632),
    .B(\mem.mem_internal.code_mem[51][3] ));
 sg13g2_nand2_1 _22324_ (.Y(_04327_),
    .A(net1027),
    .B(_04318_));
 sg13g2_o21ai_1 _22325_ (.B1(_04327_),
    .Y(_01733_),
    .A1(net326),
    .A2(_04326_));
 sg13g2_nand2_1 _22326_ (.Y(_04328_),
    .A(net632),
    .B(\mem.mem_internal.code_mem[51][4] ));
 sg13g2_nand2_1 _22327_ (.Y(_04329_),
    .A(net1026),
    .B(_04318_));
 sg13g2_o21ai_1 _22328_ (.B1(_04329_),
    .Y(_01734_),
    .A1(_04319_),
    .A2(_04328_));
 sg13g2_nand2_1 _22329_ (.Y(_04330_),
    .A(net632),
    .B(\mem.mem_internal.code_mem[51][5] ));
 sg13g2_nand2_1 _22330_ (.Y(_04331_),
    .A(net1025),
    .B(_04318_));
 sg13g2_o21ai_1 _22331_ (.B1(_04331_),
    .Y(_01735_),
    .A1(net326),
    .A2(_04330_));
 sg13g2_buf_1 _22332_ (.A(_04246_),
    .X(_04332_));
 sg13g2_nand2_1 _22333_ (.Y(_04333_),
    .A(net631),
    .B(\mem.mem_internal.code_mem[51][6] ));
 sg13g2_nand2_1 _22334_ (.Y(_04334_),
    .A(net1024),
    .B(_04318_));
 sg13g2_o21ai_1 _22335_ (.B1(_04334_),
    .Y(_01736_),
    .A1(net326),
    .A2(_04333_));
 sg13g2_nand2_1 _22336_ (.Y(_04335_),
    .A(_04332_),
    .B(\mem.mem_internal.code_mem[51][7] ));
 sg13g2_nand2_1 _22337_ (.Y(_04336_),
    .A(net1023),
    .B(_04318_));
 sg13g2_o21ai_1 _22338_ (.B1(_04336_),
    .Y(_01737_),
    .A1(net326),
    .A2(_04335_));
 sg13g2_nor2_1 _22339_ (.A(net556),
    .B(net482),
    .Y(_04337_));
 sg13g2_buf_2 _22340_ (.A(_04337_),
    .X(_04338_));
 sg13g2_buf_1 _22341_ (.A(_04338_),
    .X(_04339_));
 sg13g2_nand2_1 _22342_ (.Y(_04340_),
    .A(net631),
    .B(\mem.mem_internal.code_mem[52][0] ));
 sg13g2_nand2_1 _22343_ (.Y(_04341_),
    .A(net1030),
    .B(_04339_));
 sg13g2_o21ai_1 _22344_ (.B1(_04341_),
    .Y(_01738_),
    .A1(net325),
    .A2(_04340_));
 sg13g2_nand2_1 _22345_ (.Y(_04342_),
    .A(net631),
    .B(\mem.mem_internal.code_mem[52][1] ));
 sg13g2_nand2_1 _22346_ (.Y(_04343_),
    .A(net1029),
    .B(net325));
 sg13g2_o21ai_1 _22347_ (.B1(_04343_),
    .Y(_01739_),
    .A1(net325),
    .A2(_04342_));
 sg13g2_nand2_1 _22348_ (.Y(_04344_),
    .A(net631),
    .B(\mem.mem_internal.code_mem[52][2] ));
 sg13g2_nand2_1 _22349_ (.Y(_04345_),
    .A(net1028),
    .B(_04338_));
 sg13g2_o21ai_1 _22350_ (.B1(_04345_),
    .Y(_01740_),
    .A1(net325),
    .A2(_04344_));
 sg13g2_nand2_1 _22351_ (.Y(_04346_),
    .A(net631),
    .B(\mem.mem_internal.code_mem[52][3] ));
 sg13g2_nand2_1 _22352_ (.Y(_04347_),
    .A(net1027),
    .B(_04338_));
 sg13g2_o21ai_1 _22353_ (.B1(_04347_),
    .Y(_01741_),
    .A1(net325),
    .A2(_04346_));
 sg13g2_nand2_1 _22354_ (.Y(_04348_),
    .A(net631),
    .B(\mem.mem_internal.code_mem[52][4] ));
 sg13g2_nand2_1 _22355_ (.Y(_04349_),
    .A(net1026),
    .B(_04338_));
 sg13g2_o21ai_1 _22356_ (.B1(_04349_),
    .Y(_01742_),
    .A1(net325),
    .A2(_04348_));
 sg13g2_nand2_1 _22357_ (.Y(_04350_),
    .A(net631),
    .B(\mem.mem_internal.code_mem[52][5] ));
 sg13g2_nand2_1 _22358_ (.Y(_04351_),
    .A(net1025),
    .B(_04338_));
 sg13g2_o21ai_1 _22359_ (.B1(_04351_),
    .Y(_01743_),
    .A1(net325),
    .A2(_04350_));
 sg13g2_nand2_1 _22360_ (.Y(_04352_),
    .A(_04332_),
    .B(\mem.mem_internal.code_mem[52][6] ));
 sg13g2_nand2_1 _22361_ (.Y(_04353_),
    .A(net1024),
    .B(_04338_));
 sg13g2_o21ai_1 _22362_ (.B1(_04353_),
    .Y(_01744_),
    .A1(_04339_),
    .A2(_04352_));
 sg13g2_nand2_1 _22363_ (.Y(_04354_),
    .A(net631),
    .B(\mem.mem_internal.code_mem[52][7] ));
 sg13g2_nand2_1 _22364_ (.Y(_04355_),
    .A(net1023),
    .B(_04338_));
 sg13g2_o21ai_1 _22365_ (.B1(_04355_),
    .Y(_01745_),
    .A1(net325),
    .A2(_04354_));
 sg13g2_nor2_1 _22366_ (.A(net555),
    .B(net482),
    .Y(_04356_));
 sg13g2_buf_2 _22367_ (.A(_04356_),
    .X(_04357_));
 sg13g2_buf_1 _22368_ (.A(_04357_),
    .X(_04358_));
 sg13g2_buf_1 _22369_ (.A(_04246_),
    .X(_04359_));
 sg13g2_nand2_1 _22370_ (.Y(_04360_),
    .A(net630),
    .B(\mem.mem_internal.code_mem[53][0] ));
 sg13g2_nand2_1 _22371_ (.Y(_04361_),
    .A(net1030),
    .B(_04358_));
 sg13g2_o21ai_1 _22372_ (.B1(_04361_),
    .Y(_01746_),
    .A1(net324),
    .A2(_04360_));
 sg13g2_nand2_1 _22373_ (.Y(_04362_),
    .A(net630),
    .B(\mem.mem_internal.code_mem[53][1] ));
 sg13g2_nand2_1 _22374_ (.Y(_04363_),
    .A(net1029),
    .B(net324));
 sg13g2_o21ai_1 _22375_ (.B1(_04363_),
    .Y(_01747_),
    .A1(net324),
    .A2(_04362_));
 sg13g2_nand2_1 _22376_ (.Y(_04364_),
    .A(net630),
    .B(\mem.mem_internal.code_mem[53][2] ));
 sg13g2_nand2_1 _22377_ (.Y(_04365_),
    .A(net1028),
    .B(_04357_));
 sg13g2_o21ai_1 _22378_ (.B1(_04365_),
    .Y(_01748_),
    .A1(net324),
    .A2(_04364_));
 sg13g2_nand2_1 _22379_ (.Y(_04366_),
    .A(net630),
    .B(\mem.mem_internal.code_mem[53][3] ));
 sg13g2_nand2_1 _22380_ (.Y(_04367_),
    .A(net1027),
    .B(_04357_));
 sg13g2_o21ai_1 _22381_ (.B1(_04367_),
    .Y(_01749_),
    .A1(net324),
    .A2(_04366_));
 sg13g2_nand2_1 _22382_ (.Y(_04368_),
    .A(net630),
    .B(\mem.mem_internal.code_mem[53][4] ));
 sg13g2_nand2_1 _22383_ (.Y(_04369_),
    .A(net1026),
    .B(_04357_));
 sg13g2_o21ai_1 _22384_ (.B1(_04369_),
    .Y(_01750_),
    .A1(net324),
    .A2(_04368_));
 sg13g2_nand2_1 _22385_ (.Y(_04370_),
    .A(net630),
    .B(\mem.mem_internal.code_mem[53][5] ));
 sg13g2_nand2_1 _22386_ (.Y(_04371_),
    .A(net1025),
    .B(_04357_));
 sg13g2_o21ai_1 _22387_ (.B1(_04371_),
    .Y(_01751_),
    .A1(net324),
    .A2(_04370_));
 sg13g2_nand2_1 _22388_ (.Y(_04372_),
    .A(_04359_),
    .B(\mem.mem_internal.code_mem[53][6] ));
 sg13g2_nand2_1 _22389_ (.Y(_04373_),
    .A(net1024),
    .B(_04357_));
 sg13g2_o21ai_1 _22390_ (.B1(_04373_),
    .Y(_01752_),
    .A1(_04358_),
    .A2(_04372_));
 sg13g2_nand2_1 _22391_ (.Y(_04374_),
    .A(_04359_),
    .B(\mem.mem_internal.code_mem[53][7] ));
 sg13g2_nand2_1 _22392_ (.Y(_04375_),
    .A(net1023),
    .B(_04357_));
 sg13g2_o21ai_1 _22393_ (.B1(_04375_),
    .Y(_01753_),
    .A1(net324),
    .A2(_04374_));
 sg13g2_nor2_1 _22394_ (.A(net554),
    .B(net482),
    .Y(_04376_));
 sg13g2_buf_2 _22395_ (.A(_04376_),
    .X(_04377_));
 sg13g2_buf_1 _22396_ (.A(_04377_),
    .X(_04378_));
 sg13g2_nand2_1 _22397_ (.Y(_04379_),
    .A(net630),
    .B(\mem.mem_internal.code_mem[54][0] ));
 sg13g2_nand2_1 _22398_ (.Y(_04380_),
    .A(net1030),
    .B(_04378_));
 sg13g2_o21ai_1 _22399_ (.B1(_04380_),
    .Y(_01754_),
    .A1(net323),
    .A2(_04379_));
 sg13g2_nand2_1 _22400_ (.Y(_04381_),
    .A(net630),
    .B(\mem.mem_internal.code_mem[54][1] ));
 sg13g2_nand2_1 _22401_ (.Y(_04382_),
    .A(net1029),
    .B(net323));
 sg13g2_o21ai_1 _22402_ (.B1(_04382_),
    .Y(_01755_),
    .A1(net323),
    .A2(_04381_));
 sg13g2_buf_1 _22403_ (.A(_04246_),
    .X(_04383_));
 sg13g2_nand2_1 _22404_ (.Y(_04384_),
    .A(net629),
    .B(\mem.mem_internal.code_mem[54][2] ));
 sg13g2_nand2_1 _22405_ (.Y(_04385_),
    .A(net1028),
    .B(_04377_));
 sg13g2_o21ai_1 _22406_ (.B1(_04385_),
    .Y(_01756_),
    .A1(net323),
    .A2(_04384_));
 sg13g2_nand2_1 _22407_ (.Y(_04386_),
    .A(net629),
    .B(\mem.mem_internal.code_mem[54][3] ));
 sg13g2_nand2_1 _22408_ (.Y(_04387_),
    .A(net1027),
    .B(_04377_));
 sg13g2_o21ai_1 _22409_ (.B1(_04387_),
    .Y(_01757_),
    .A1(net323),
    .A2(_04386_));
 sg13g2_nand2_1 _22410_ (.Y(_04388_),
    .A(net629),
    .B(\mem.mem_internal.code_mem[54][4] ));
 sg13g2_nand2_1 _22411_ (.Y(_04389_),
    .A(net1026),
    .B(_04377_));
 sg13g2_o21ai_1 _22412_ (.B1(_04389_),
    .Y(_01758_),
    .A1(net323),
    .A2(_04388_));
 sg13g2_nand2_1 _22413_ (.Y(_04390_),
    .A(net629),
    .B(\mem.mem_internal.code_mem[54][5] ));
 sg13g2_nand2_1 _22414_ (.Y(_04391_),
    .A(net1025),
    .B(_04377_));
 sg13g2_o21ai_1 _22415_ (.B1(_04391_),
    .Y(_01759_),
    .A1(net323),
    .A2(_04390_));
 sg13g2_nand2_1 _22416_ (.Y(_04392_),
    .A(net629),
    .B(\mem.mem_internal.code_mem[54][6] ));
 sg13g2_nand2_1 _22417_ (.Y(_04393_),
    .A(net1024),
    .B(_04377_));
 sg13g2_o21ai_1 _22418_ (.B1(_04393_),
    .Y(_01760_),
    .A1(net323),
    .A2(_04392_));
 sg13g2_nand2_1 _22419_ (.Y(_04394_),
    .A(_04383_),
    .B(\mem.mem_internal.code_mem[54][7] ));
 sg13g2_nand2_1 _22420_ (.Y(_04395_),
    .A(net1023),
    .B(_04377_));
 sg13g2_o21ai_1 _22421_ (.B1(_04395_),
    .Y(_01761_),
    .A1(_04378_),
    .A2(_04394_));
 sg13g2_nor2_1 _22422_ (.A(net553),
    .B(net482),
    .Y(_04396_));
 sg13g2_buf_2 _22423_ (.A(_04396_),
    .X(_04397_));
 sg13g2_buf_1 _22424_ (.A(_04397_),
    .X(_04398_));
 sg13g2_nand2_1 _22425_ (.Y(_04399_),
    .A(_04383_),
    .B(\mem.mem_internal.code_mem[55][0] ));
 sg13g2_nand2_1 _22426_ (.Y(_04400_),
    .A(net1030),
    .B(_04398_));
 sg13g2_o21ai_1 _22427_ (.B1(_04400_),
    .Y(_01762_),
    .A1(net322),
    .A2(_04399_));
 sg13g2_nand2_1 _22428_ (.Y(_04401_),
    .A(net629),
    .B(\mem.mem_internal.code_mem[55][1] ));
 sg13g2_nand2_1 _22429_ (.Y(_04402_),
    .A(net1029),
    .B(net322));
 sg13g2_o21ai_1 _22430_ (.B1(_04402_),
    .Y(_01763_),
    .A1(net322),
    .A2(_04401_));
 sg13g2_nand2_1 _22431_ (.Y(_04403_),
    .A(net629),
    .B(\mem.mem_internal.code_mem[55][2] ));
 sg13g2_nand2_1 _22432_ (.Y(_04404_),
    .A(net1028),
    .B(_04397_));
 sg13g2_o21ai_1 _22433_ (.B1(_04404_),
    .Y(_01764_),
    .A1(net322),
    .A2(_04403_));
 sg13g2_nand2_1 _22434_ (.Y(_04405_),
    .A(net629),
    .B(\mem.mem_internal.code_mem[55][3] ));
 sg13g2_nand2_1 _22435_ (.Y(_04406_),
    .A(net1027),
    .B(_04397_));
 sg13g2_o21ai_1 _22436_ (.B1(_04406_),
    .Y(_01765_),
    .A1(net322),
    .A2(_04405_));
 sg13g2_buf_1 _22437_ (.A(_04246_),
    .X(_04407_));
 sg13g2_nand2_1 _22438_ (.Y(_04408_),
    .A(net628),
    .B(\mem.mem_internal.code_mem[55][4] ));
 sg13g2_nand2_1 _22439_ (.Y(_04409_),
    .A(net1026),
    .B(_04397_));
 sg13g2_o21ai_1 _22440_ (.B1(_04409_),
    .Y(_01766_),
    .A1(net322),
    .A2(_04408_));
 sg13g2_nand2_1 _22441_ (.Y(_04410_),
    .A(net628),
    .B(\mem.mem_internal.code_mem[55][5] ));
 sg13g2_nand2_1 _22442_ (.Y(_04411_),
    .A(net1025),
    .B(_04397_));
 sg13g2_o21ai_1 _22443_ (.B1(_04411_),
    .Y(_01767_),
    .A1(net322),
    .A2(_04410_));
 sg13g2_nand2_1 _22444_ (.Y(_04412_),
    .A(net628),
    .B(\mem.mem_internal.code_mem[55][6] ));
 sg13g2_nand2_1 _22445_ (.Y(_04413_),
    .A(net1024),
    .B(_04397_));
 sg13g2_o21ai_1 _22446_ (.B1(_04413_),
    .Y(_01768_),
    .A1(net322),
    .A2(_04412_));
 sg13g2_nand2_1 _22447_ (.Y(_04414_),
    .A(net628),
    .B(\mem.mem_internal.code_mem[55][7] ));
 sg13g2_nand2_1 _22448_ (.Y(_04415_),
    .A(net1023),
    .B(_04397_));
 sg13g2_o21ai_1 _22449_ (.B1(_04415_),
    .Y(_01769_),
    .A1(_04398_),
    .A2(_04414_));
 sg13g2_nor2_1 _22450_ (.A(net552),
    .B(_04228_),
    .Y(_04416_));
 sg13g2_buf_2 _22451_ (.A(_04416_),
    .X(_04417_));
 sg13g2_buf_1 _22452_ (.A(_04417_),
    .X(_04418_));
 sg13g2_nand2_1 _22453_ (.Y(_04419_),
    .A(net628),
    .B(\mem.mem_internal.code_mem[56][0] ));
 sg13g2_nand2_1 _22454_ (.Y(_04420_),
    .A(net1030),
    .B(net321));
 sg13g2_o21ai_1 _22455_ (.B1(_04420_),
    .Y(_01770_),
    .A1(net321),
    .A2(_04419_));
 sg13g2_nand2_1 _22456_ (.Y(_04421_),
    .A(net628),
    .B(\mem.mem_internal.code_mem[56][1] ));
 sg13g2_nand2_1 _22457_ (.Y(_04422_),
    .A(net1029),
    .B(net321));
 sg13g2_o21ai_1 _22458_ (.B1(_04422_),
    .Y(_01771_),
    .A1(net321),
    .A2(_04421_));
 sg13g2_nand2_1 _22459_ (.Y(_04423_),
    .A(net628),
    .B(\mem.mem_internal.code_mem[56][2] ));
 sg13g2_nand2_1 _22460_ (.Y(_04424_),
    .A(net1028),
    .B(_04417_));
 sg13g2_o21ai_1 _22461_ (.B1(_04424_),
    .Y(_01772_),
    .A1(_04418_),
    .A2(_04423_));
 sg13g2_nand2_1 _22462_ (.Y(_04425_),
    .A(net628),
    .B(\mem.mem_internal.code_mem[56][3] ));
 sg13g2_nand2_1 _22463_ (.Y(_04426_),
    .A(net1027),
    .B(_04417_));
 sg13g2_o21ai_1 _22464_ (.B1(_04426_),
    .Y(_01773_),
    .A1(_04418_),
    .A2(_04425_));
 sg13g2_nand2_1 _22465_ (.Y(_04427_),
    .A(_04407_),
    .B(\mem.mem_internal.code_mem[56][4] ));
 sg13g2_nand2_1 _22466_ (.Y(_04428_),
    .A(net1026),
    .B(_04417_));
 sg13g2_o21ai_1 _22467_ (.B1(_04428_),
    .Y(_01774_),
    .A1(net321),
    .A2(_04427_));
 sg13g2_nand2_1 _22468_ (.Y(_04429_),
    .A(_04407_),
    .B(\mem.mem_internal.code_mem[56][5] ));
 sg13g2_nand2_1 _22469_ (.Y(_04430_),
    .A(net1025),
    .B(_04417_));
 sg13g2_o21ai_1 _22470_ (.B1(_04430_),
    .Y(_01775_),
    .A1(net321),
    .A2(_04429_));
 sg13g2_buf_2 _22471_ (.A(net1276),
    .X(_04431_));
 sg13g2_buf_1 _22472_ (.A(_04431_),
    .X(_04432_));
 sg13g2_buf_1 _22473_ (.A(_04432_),
    .X(_04433_));
 sg13g2_nand2_1 _22474_ (.Y(_04434_),
    .A(net627),
    .B(\mem.mem_internal.code_mem[56][6] ));
 sg13g2_nand2_1 _22475_ (.Y(_04435_),
    .A(net1024),
    .B(_04417_));
 sg13g2_o21ai_1 _22476_ (.B1(_04435_),
    .Y(_01776_),
    .A1(net321),
    .A2(_04434_));
 sg13g2_nand2_1 _22477_ (.Y(_04436_),
    .A(net627),
    .B(\mem.mem_internal.code_mem[56][7] ));
 sg13g2_nand2_1 _22478_ (.Y(_04437_),
    .A(net1023),
    .B(_04417_));
 sg13g2_o21ai_1 _22479_ (.B1(_04437_),
    .Y(_01777_),
    .A1(net321),
    .A2(_04436_));
 sg13g2_nor2_1 _22480_ (.A(net551),
    .B(_04228_),
    .Y(_04438_));
 sg13g2_buf_2 _22481_ (.A(_04438_),
    .X(_04439_));
 sg13g2_buf_1 _22482_ (.A(_04439_),
    .X(_04440_));
 sg13g2_nand2_1 _22483_ (.Y(_04441_),
    .A(net627),
    .B(\mem.mem_internal.code_mem[57][0] ));
 sg13g2_nand2_1 _22484_ (.Y(_04442_),
    .A(net1030),
    .B(net320));
 sg13g2_o21ai_1 _22485_ (.B1(_04442_),
    .Y(_01778_),
    .A1(net320),
    .A2(_04441_));
 sg13g2_nand2_1 _22486_ (.Y(_04443_),
    .A(_04433_),
    .B(\mem.mem_internal.code_mem[57][1] ));
 sg13g2_nand2_1 _22487_ (.Y(_04444_),
    .A(net1029),
    .B(_04440_));
 sg13g2_o21ai_1 _22488_ (.B1(_04444_),
    .Y(_01779_),
    .A1(_04440_),
    .A2(_04443_));
 sg13g2_nand2_1 _22489_ (.Y(_04445_),
    .A(net627),
    .B(\mem.mem_internal.code_mem[57][2] ));
 sg13g2_nand2_1 _22490_ (.Y(_04446_),
    .A(net1028),
    .B(_04439_));
 sg13g2_o21ai_1 _22491_ (.B1(_04446_),
    .Y(_01780_),
    .A1(net320),
    .A2(_04445_));
 sg13g2_nand2_1 _22492_ (.Y(_04447_),
    .A(net627),
    .B(\mem.mem_internal.code_mem[57][3] ));
 sg13g2_nand2_1 _22493_ (.Y(_04448_),
    .A(net1027),
    .B(_04439_));
 sg13g2_o21ai_1 _22494_ (.B1(_04448_),
    .Y(_01781_),
    .A1(net320),
    .A2(_04447_));
 sg13g2_nand2_1 _22495_ (.Y(_04449_),
    .A(_04433_),
    .B(\mem.mem_internal.code_mem[57][4] ));
 sg13g2_nand2_1 _22496_ (.Y(_04450_),
    .A(net1026),
    .B(_04439_));
 sg13g2_o21ai_1 _22497_ (.B1(_04450_),
    .Y(_01782_),
    .A1(net320),
    .A2(_04449_));
 sg13g2_nand2_1 _22498_ (.Y(_04451_),
    .A(net627),
    .B(\mem.mem_internal.code_mem[57][5] ));
 sg13g2_nand2_1 _22499_ (.Y(_04452_),
    .A(net1025),
    .B(_04439_));
 sg13g2_o21ai_1 _22500_ (.B1(_04452_),
    .Y(_01783_),
    .A1(net320),
    .A2(_04451_));
 sg13g2_nand2_1 _22501_ (.Y(_04453_),
    .A(net627),
    .B(\mem.mem_internal.code_mem[57][6] ));
 sg13g2_nand2_1 _22502_ (.Y(_04454_),
    .A(net1024),
    .B(_04439_));
 sg13g2_o21ai_1 _22503_ (.B1(_04454_),
    .Y(_01784_),
    .A1(net320),
    .A2(_04453_));
 sg13g2_nand2_1 _22504_ (.Y(_04455_),
    .A(net627),
    .B(\mem.mem_internal.code_mem[57][7] ));
 sg13g2_nand2_1 _22505_ (.Y(_04456_),
    .A(net1023),
    .B(_04439_));
 sg13g2_o21ai_1 _22506_ (.B1(_04456_),
    .Y(_01785_),
    .A1(net320),
    .A2(_04455_));
 sg13g2_nor2_1 _22507_ (.A(net550),
    .B(_04227_),
    .Y(_04457_));
 sg13g2_buf_2 _22508_ (.A(_04457_),
    .X(_04458_));
 sg13g2_buf_1 _22509_ (.A(_04458_),
    .X(_04459_));
 sg13g2_buf_1 _22510_ (.A(_04432_),
    .X(_04460_));
 sg13g2_nand2_1 _22511_ (.Y(_04461_),
    .A(net626),
    .B(\mem.mem_internal.code_mem[58][0] ));
 sg13g2_nand2_1 _22512_ (.Y(_04462_),
    .A(_04273_),
    .B(net444));
 sg13g2_o21ai_1 _22513_ (.B1(_04462_),
    .Y(_01786_),
    .A1(net444),
    .A2(_04461_));
 sg13g2_nand2_1 _22514_ (.Y(_04463_),
    .A(_04460_),
    .B(\mem.mem_internal.code_mem[58][1] ));
 sg13g2_nand2_1 _22515_ (.Y(_04464_),
    .A(_04276_),
    .B(net444));
 sg13g2_o21ai_1 _22516_ (.B1(_04464_),
    .Y(_01787_),
    .A1(net444),
    .A2(_04463_));
 sg13g2_nand2_1 _22517_ (.Y(_04465_),
    .A(net626),
    .B(\mem.mem_internal.code_mem[58][2] ));
 sg13g2_nand2_1 _22518_ (.Y(_04466_),
    .A(_04280_),
    .B(_04458_));
 sg13g2_o21ai_1 _22519_ (.B1(_04466_),
    .Y(_01788_),
    .A1(net444),
    .A2(_04465_));
 sg13g2_nand2_1 _22520_ (.Y(_04467_),
    .A(net626),
    .B(\mem.mem_internal.code_mem[58][3] ));
 sg13g2_nand2_1 _22521_ (.Y(_04468_),
    .A(_04283_),
    .B(_04458_));
 sg13g2_o21ai_1 _22522_ (.B1(_04468_),
    .Y(_01789_),
    .A1(_04459_),
    .A2(_04467_));
 sg13g2_nand2_1 _22523_ (.Y(_04469_),
    .A(net626),
    .B(\mem.mem_internal.code_mem[58][4] ));
 sg13g2_nand2_1 _22524_ (.Y(_04470_),
    .A(_04286_),
    .B(_04458_));
 sg13g2_o21ai_1 _22525_ (.B1(_04470_),
    .Y(_01790_),
    .A1(_04459_),
    .A2(_04469_));
 sg13g2_nand2_1 _22526_ (.Y(_04471_),
    .A(net626),
    .B(\mem.mem_internal.code_mem[58][5] ));
 sg13g2_nand2_1 _22527_ (.Y(_04472_),
    .A(_04289_),
    .B(_04458_));
 sg13g2_o21ai_1 _22528_ (.B1(_04472_),
    .Y(_01791_),
    .A1(net444),
    .A2(_04471_));
 sg13g2_nand2_1 _22529_ (.Y(_04473_),
    .A(net626),
    .B(\mem.mem_internal.code_mem[58][6] ));
 sg13g2_nand2_1 _22530_ (.Y(_04474_),
    .A(_04292_),
    .B(_04458_));
 sg13g2_o21ai_1 _22531_ (.B1(_04474_),
    .Y(_01792_),
    .A1(net444),
    .A2(_04473_));
 sg13g2_nand2_1 _22532_ (.Y(_04475_),
    .A(net626),
    .B(\mem.mem_internal.code_mem[58][7] ));
 sg13g2_nand2_1 _22533_ (.Y(_04476_),
    .A(_04295_),
    .B(_04458_));
 sg13g2_o21ai_1 _22534_ (.B1(_04476_),
    .Y(_01793_),
    .A1(net444),
    .A2(_04475_));
 sg13g2_nor2_1 _22535_ (.A(net549),
    .B(_04227_),
    .Y(_04477_));
 sg13g2_buf_2 _22536_ (.A(_04477_),
    .X(_04478_));
 sg13g2_buf_1 _22537_ (.A(_04478_),
    .X(_04479_));
 sg13g2_nand2_1 _22538_ (.Y(_04480_),
    .A(net626),
    .B(\mem.mem_internal.code_mem[59][0] ));
 sg13g2_buf_1 _22539_ (.A(_03842_),
    .X(_04481_));
 sg13g2_nand2_1 _22540_ (.Y(_04482_),
    .A(net1022),
    .B(net443));
 sg13g2_o21ai_1 _22541_ (.B1(_04482_),
    .Y(_01794_),
    .A1(net443),
    .A2(_04480_));
 sg13g2_nand2_1 _22542_ (.Y(_04483_),
    .A(_04460_),
    .B(\mem.mem_internal.code_mem[59][1] ));
 sg13g2_buf_1 _22543_ (.A(_03846_),
    .X(_04484_));
 sg13g2_nand2_1 _22544_ (.Y(_04485_),
    .A(net1021),
    .B(net443));
 sg13g2_o21ai_1 _22545_ (.B1(_04485_),
    .Y(_01795_),
    .A1(net443),
    .A2(_04483_));
 sg13g2_buf_1 _22546_ (.A(_04432_),
    .X(_04486_));
 sg13g2_nand2_1 _22547_ (.Y(_04487_),
    .A(net625),
    .B(\mem.mem_internal.code_mem[59][2] ));
 sg13g2_buf_1 _22548_ (.A(_03850_),
    .X(_04488_));
 sg13g2_nand2_1 _22549_ (.Y(_04489_),
    .A(_04488_),
    .B(_04478_));
 sg13g2_o21ai_1 _22550_ (.B1(_04489_),
    .Y(_01796_),
    .A1(net443),
    .A2(_04487_));
 sg13g2_nand2_1 _22551_ (.Y(_04490_),
    .A(net625),
    .B(\mem.mem_internal.code_mem[59][3] ));
 sg13g2_buf_1 _22552_ (.A(_03854_),
    .X(_04491_));
 sg13g2_nand2_1 _22553_ (.Y(_04492_),
    .A(_04491_),
    .B(_04478_));
 sg13g2_o21ai_1 _22554_ (.B1(_04492_),
    .Y(_01797_),
    .A1(net443),
    .A2(_04490_));
 sg13g2_nand2_1 _22555_ (.Y(_04493_),
    .A(net625),
    .B(\mem.mem_internal.code_mem[59][4] ));
 sg13g2_buf_1 _22556_ (.A(_03859_),
    .X(_04494_));
 sg13g2_nand2_1 _22557_ (.Y(_04495_),
    .A(net1018),
    .B(_04478_));
 sg13g2_o21ai_1 _22558_ (.B1(_04495_),
    .Y(_01798_),
    .A1(net443),
    .A2(_04493_));
 sg13g2_nand2_1 _22559_ (.Y(_04496_),
    .A(net625),
    .B(\mem.mem_internal.code_mem[59][5] ));
 sg13g2_buf_1 _22560_ (.A(_03863_),
    .X(_04497_));
 sg13g2_nand2_1 _22561_ (.Y(_04498_),
    .A(net1017),
    .B(_04478_));
 sg13g2_o21ai_1 _22562_ (.B1(_04498_),
    .Y(_01799_),
    .A1(net443),
    .A2(_04496_));
 sg13g2_nand2_1 _22563_ (.Y(_04499_),
    .A(net625),
    .B(\mem.mem_internal.code_mem[59][6] ));
 sg13g2_buf_1 _22564_ (.A(_03867_),
    .X(_04500_));
 sg13g2_nand2_1 _22565_ (.Y(_04501_),
    .A(net1016),
    .B(_04478_));
 sg13g2_o21ai_1 _22566_ (.B1(_04501_),
    .Y(_01800_),
    .A1(_04479_),
    .A2(_04499_));
 sg13g2_nand2_1 _22567_ (.Y(_04502_),
    .A(net625),
    .B(\mem.mem_internal.code_mem[59][7] ));
 sg13g2_buf_1 _22568_ (.A(_03871_),
    .X(_04503_));
 sg13g2_nand2_1 _22569_ (.Y(_04504_),
    .A(net1015),
    .B(_04478_));
 sg13g2_o21ai_1 _22570_ (.B1(_04504_),
    .Y(_01801_),
    .A1(_04479_),
    .A2(_04502_));
 sg13g2_nand2_1 _22571_ (.Y(_04505_),
    .A(net836),
    .B(\mem.mem_internal.code_mem[5][0] ));
 sg13g2_nor2_1 _22572_ (.A(_10246_),
    .B(net555),
    .Y(_04506_));
 sg13g2_buf_1 _22573_ (.A(_04506_),
    .X(_04507_));
 sg13g2_buf_1 _22574_ (.A(_04507_),
    .X(_04508_));
 sg13g2_nand2_1 _22575_ (.Y(_04509_),
    .A(net1022),
    .B(net319));
 sg13g2_o21ai_1 _22576_ (.B1(_04509_),
    .Y(_01802_),
    .A1(_04505_),
    .A2(net319));
 sg13g2_nand2_1 _22577_ (.Y(_04510_),
    .A(net625),
    .B(\mem.mem_internal.code_mem[5][1] ));
 sg13g2_nand2_1 _22578_ (.Y(_04511_),
    .A(net1021),
    .B(net319));
 sg13g2_o21ai_1 _22579_ (.B1(_04511_),
    .Y(_01803_),
    .A1(net319),
    .A2(_04510_));
 sg13g2_nand2_1 _22580_ (.Y(_04512_),
    .A(net625),
    .B(\mem.mem_internal.code_mem[5][2] ));
 sg13g2_nand2_1 _22581_ (.Y(_04513_),
    .A(net1020),
    .B(_04507_));
 sg13g2_o21ai_1 _22582_ (.B1(_04513_),
    .Y(_01804_),
    .A1(net319),
    .A2(_04512_));
 sg13g2_nand2_1 _22583_ (.Y(_04514_),
    .A(_04486_),
    .B(\mem.mem_internal.code_mem[5][3] ));
 sg13g2_nand2_1 _22584_ (.Y(_04515_),
    .A(net1019),
    .B(_04507_));
 sg13g2_o21ai_1 _22585_ (.B1(_04515_),
    .Y(_01805_),
    .A1(_04508_),
    .A2(_04514_));
 sg13g2_nand2_1 _22586_ (.Y(_04516_),
    .A(_04486_),
    .B(\mem.mem_internal.code_mem[5][4] ));
 sg13g2_nand2_1 _22587_ (.Y(_04517_),
    .A(net1018),
    .B(_04507_));
 sg13g2_o21ai_1 _22588_ (.B1(_04517_),
    .Y(_01806_),
    .A1(_04508_),
    .A2(_04516_));
 sg13g2_buf_1 _22589_ (.A(_04432_),
    .X(_04518_));
 sg13g2_nand2_1 _22590_ (.Y(_04519_),
    .A(_04518_),
    .B(\mem.mem_internal.code_mem[5][5] ));
 sg13g2_nand2_1 _22591_ (.Y(_04520_),
    .A(net1017),
    .B(_04507_));
 sg13g2_o21ai_1 _22592_ (.B1(_04520_),
    .Y(_01807_),
    .A1(net319),
    .A2(_04519_));
 sg13g2_nand2_1 _22593_ (.Y(_04521_),
    .A(net624),
    .B(\mem.mem_internal.code_mem[5][6] ));
 sg13g2_nand2_1 _22594_ (.Y(_04522_),
    .A(net1016),
    .B(_04507_));
 sg13g2_o21ai_1 _22595_ (.B1(_04522_),
    .Y(_01808_),
    .A1(net319),
    .A2(_04521_));
 sg13g2_nand2_1 _22596_ (.Y(_04523_),
    .A(_04518_),
    .B(\mem.mem_internal.code_mem[5][7] ));
 sg13g2_nand2_1 _22597_ (.Y(_04524_),
    .A(net1015),
    .B(_04507_));
 sg13g2_o21ai_1 _22598_ (.B1(_04524_),
    .Y(_01809_),
    .A1(net319),
    .A2(_04523_));
 sg13g2_nor2_1 _22599_ (.A(net773),
    .B(_04227_),
    .Y(_04525_));
 sg13g2_buf_2 _22600_ (.A(_04525_),
    .X(_04526_));
 sg13g2_buf_1 _22601_ (.A(_04526_),
    .X(_04527_));
 sg13g2_nand2_1 _22602_ (.Y(_04528_),
    .A(net624),
    .B(\mem.mem_internal.code_mem[60][0] ));
 sg13g2_nand2_1 _22603_ (.Y(_04529_),
    .A(net1022),
    .B(net442));
 sg13g2_o21ai_1 _22604_ (.B1(_04529_),
    .Y(_01810_),
    .A1(net442),
    .A2(_04528_));
 sg13g2_nand2_1 _22605_ (.Y(_04530_),
    .A(net624),
    .B(\mem.mem_internal.code_mem[60][1] ));
 sg13g2_nand2_1 _22606_ (.Y(_04531_),
    .A(net1021),
    .B(net442));
 sg13g2_o21ai_1 _22607_ (.B1(_04531_),
    .Y(_01811_),
    .A1(net442),
    .A2(_04530_));
 sg13g2_nand2_1 _22608_ (.Y(_04532_),
    .A(net624),
    .B(\mem.mem_internal.code_mem[60][2] ));
 sg13g2_nand2_1 _22609_ (.Y(_04533_),
    .A(net1020),
    .B(_04526_));
 sg13g2_o21ai_1 _22610_ (.B1(_04533_),
    .Y(_01812_),
    .A1(net442),
    .A2(_04532_));
 sg13g2_nand2_1 _22611_ (.Y(_04534_),
    .A(net624),
    .B(\mem.mem_internal.code_mem[60][3] ));
 sg13g2_nand2_1 _22612_ (.Y(_04535_),
    .A(net1019),
    .B(_04526_));
 sg13g2_o21ai_1 _22613_ (.B1(_04535_),
    .Y(_01813_),
    .A1(net442),
    .A2(_04534_));
 sg13g2_nand2_1 _22614_ (.Y(_04536_),
    .A(net624),
    .B(\mem.mem_internal.code_mem[60][4] ));
 sg13g2_nand2_1 _22615_ (.Y(_04537_),
    .A(net1018),
    .B(_04526_));
 sg13g2_o21ai_1 _22616_ (.B1(_04537_),
    .Y(_01814_),
    .A1(net442),
    .A2(_04536_));
 sg13g2_nand2_1 _22617_ (.Y(_04538_),
    .A(net624),
    .B(\mem.mem_internal.code_mem[60][5] ));
 sg13g2_nand2_1 _22618_ (.Y(_04539_),
    .A(net1017),
    .B(_04526_));
 sg13g2_o21ai_1 _22619_ (.B1(_04539_),
    .Y(_01815_),
    .A1(_04527_),
    .A2(_04538_));
 sg13g2_nand2_1 _22620_ (.Y(_04540_),
    .A(net624),
    .B(\mem.mem_internal.code_mem[60][6] ));
 sg13g2_nand2_1 _22621_ (.Y(_04541_),
    .A(net1016),
    .B(_04526_));
 sg13g2_o21ai_1 _22622_ (.B1(_04541_),
    .Y(_01816_),
    .A1(_04527_),
    .A2(_04540_));
 sg13g2_buf_1 _22623_ (.A(_04432_),
    .X(_04542_));
 sg13g2_nand2_1 _22624_ (.Y(_04543_),
    .A(net623),
    .B(\mem.mem_internal.code_mem[60][7] ));
 sg13g2_nand2_1 _22625_ (.Y(_04544_),
    .A(net1015),
    .B(_04526_));
 sg13g2_o21ai_1 _22626_ (.B1(_04544_),
    .Y(_01817_),
    .A1(net442),
    .A2(_04543_));
 sg13g2_nor2_1 _22627_ (.A(net548),
    .B(_04227_),
    .Y(_04545_));
 sg13g2_buf_2 _22628_ (.A(_04545_),
    .X(_04546_));
 sg13g2_buf_1 _22629_ (.A(_04546_),
    .X(_04547_));
 sg13g2_nand2_1 _22630_ (.Y(_04548_),
    .A(net623),
    .B(\mem.mem_internal.code_mem[61][0] ));
 sg13g2_nand2_1 _22631_ (.Y(_04549_),
    .A(net1022),
    .B(net441));
 sg13g2_o21ai_1 _22632_ (.B1(_04549_),
    .Y(_01818_),
    .A1(net441),
    .A2(_04548_));
 sg13g2_nand2_1 _22633_ (.Y(_04550_),
    .A(net623),
    .B(\mem.mem_internal.code_mem[61][1] ));
 sg13g2_nand2_1 _22634_ (.Y(_04551_),
    .A(net1021),
    .B(net441));
 sg13g2_o21ai_1 _22635_ (.B1(_04551_),
    .Y(_01819_),
    .A1(net441),
    .A2(_04550_));
 sg13g2_nand2_1 _22636_ (.Y(_04552_),
    .A(net623),
    .B(\mem.mem_internal.code_mem[61][2] ));
 sg13g2_nand2_1 _22637_ (.Y(_04553_),
    .A(net1020),
    .B(_04546_));
 sg13g2_o21ai_1 _22638_ (.B1(_04553_),
    .Y(_01820_),
    .A1(net441),
    .A2(_04552_));
 sg13g2_nand2_1 _22639_ (.Y(_04554_),
    .A(net623),
    .B(\mem.mem_internal.code_mem[61][3] ));
 sg13g2_nand2_1 _22640_ (.Y(_04555_),
    .A(net1019),
    .B(_04546_));
 sg13g2_o21ai_1 _22641_ (.B1(_04555_),
    .Y(_01821_),
    .A1(net441),
    .A2(_04554_));
 sg13g2_nand2_1 _22642_ (.Y(_04556_),
    .A(net623),
    .B(\mem.mem_internal.code_mem[61][4] ));
 sg13g2_nand2_1 _22643_ (.Y(_04557_),
    .A(net1018),
    .B(_04546_));
 sg13g2_o21ai_1 _22644_ (.B1(_04557_),
    .Y(_01822_),
    .A1(net441),
    .A2(_04556_));
 sg13g2_nand2_1 _22645_ (.Y(_04558_),
    .A(_04542_),
    .B(\mem.mem_internal.code_mem[61][5] ));
 sg13g2_nand2_1 _22646_ (.Y(_04559_),
    .A(net1017),
    .B(_04546_));
 sg13g2_o21ai_1 _22647_ (.B1(_04559_),
    .Y(_01823_),
    .A1(_04547_),
    .A2(_04558_));
 sg13g2_nand2_1 _22648_ (.Y(_04560_),
    .A(net623),
    .B(\mem.mem_internal.code_mem[61][6] ));
 sg13g2_nand2_1 _22649_ (.Y(_04561_),
    .A(net1016),
    .B(_04546_));
 sg13g2_o21ai_1 _22650_ (.B1(_04561_),
    .Y(_01824_),
    .A1(_04547_),
    .A2(_04560_));
 sg13g2_nand2_1 _22651_ (.Y(_04562_),
    .A(_04542_),
    .B(\mem.mem_internal.code_mem[61][7] ));
 sg13g2_nand2_1 _22652_ (.Y(_04563_),
    .A(net1015),
    .B(_04546_));
 sg13g2_o21ai_1 _22653_ (.B1(_04563_),
    .Y(_01825_),
    .A1(net441),
    .A2(_04562_));
 sg13g2_nor2_1 _22654_ (.A(net547),
    .B(_04227_),
    .Y(_04564_));
 sg13g2_buf_2 _22655_ (.A(_04564_),
    .X(_04565_));
 sg13g2_buf_1 _22656_ (.A(_04565_),
    .X(_04566_));
 sg13g2_nand2_1 _22657_ (.Y(_04567_),
    .A(net623),
    .B(\mem.mem_internal.code_mem[62][0] ));
 sg13g2_nand2_1 _22658_ (.Y(_04568_),
    .A(net1022),
    .B(net440));
 sg13g2_o21ai_1 _22659_ (.B1(_04568_),
    .Y(_01826_),
    .A1(net440),
    .A2(_04567_));
 sg13g2_buf_1 _22660_ (.A(_04432_),
    .X(_04569_));
 sg13g2_nand2_1 _22661_ (.Y(_04570_),
    .A(net622),
    .B(\mem.mem_internal.code_mem[62][1] ));
 sg13g2_nand2_1 _22662_ (.Y(_04571_),
    .A(net1021),
    .B(net440));
 sg13g2_o21ai_1 _22663_ (.B1(_04571_),
    .Y(_01827_),
    .A1(net440),
    .A2(_04570_));
 sg13g2_nand2_1 _22664_ (.Y(_04572_),
    .A(net622),
    .B(\mem.mem_internal.code_mem[62][2] ));
 sg13g2_nand2_1 _22665_ (.Y(_04573_),
    .A(net1020),
    .B(_04565_));
 sg13g2_o21ai_1 _22666_ (.B1(_04573_),
    .Y(_01828_),
    .A1(net440),
    .A2(_04572_));
 sg13g2_nand2_1 _22667_ (.Y(_04574_),
    .A(net622),
    .B(\mem.mem_internal.code_mem[62][3] ));
 sg13g2_nand2_1 _22668_ (.Y(_04575_),
    .A(net1019),
    .B(_04565_));
 sg13g2_o21ai_1 _22669_ (.B1(_04575_),
    .Y(_01829_),
    .A1(net440),
    .A2(_04574_));
 sg13g2_nand2_1 _22670_ (.Y(_04576_),
    .A(net622),
    .B(\mem.mem_internal.code_mem[62][4] ));
 sg13g2_nand2_1 _22671_ (.Y(_04577_),
    .A(_04494_),
    .B(_04565_));
 sg13g2_o21ai_1 _22672_ (.B1(_04577_),
    .Y(_01830_),
    .A1(net440),
    .A2(_04576_));
 sg13g2_nand2_1 _22673_ (.Y(_04578_),
    .A(net622),
    .B(\mem.mem_internal.code_mem[62][5] ));
 sg13g2_nand2_1 _22674_ (.Y(_04579_),
    .A(_04497_),
    .B(_04565_));
 sg13g2_o21ai_1 _22675_ (.B1(_04579_),
    .Y(_01831_),
    .A1(_04566_),
    .A2(_04578_));
 sg13g2_nand2_1 _22676_ (.Y(_04580_),
    .A(_04569_),
    .B(\mem.mem_internal.code_mem[62][6] ));
 sg13g2_nand2_1 _22677_ (.Y(_04581_),
    .A(net1016),
    .B(_04565_));
 sg13g2_o21ai_1 _22678_ (.B1(_04581_),
    .Y(_01832_),
    .A1(_04566_),
    .A2(_04580_));
 sg13g2_nand2_1 _22679_ (.Y(_04582_),
    .A(_04569_),
    .B(\mem.mem_internal.code_mem[62][7] ));
 sg13g2_nand2_1 _22680_ (.Y(_04583_),
    .A(net1015),
    .B(_04565_));
 sg13g2_o21ai_1 _22681_ (.B1(_04583_),
    .Y(_01833_),
    .A1(net440),
    .A2(_04582_));
 sg13g2_nor2_1 _22682_ (.A(net770),
    .B(_04227_),
    .Y(_04584_));
 sg13g2_buf_2 _22683_ (.A(_04584_),
    .X(_04585_));
 sg13g2_buf_1 _22684_ (.A(_04585_),
    .X(_04586_));
 sg13g2_nand2_1 _22685_ (.Y(_04587_),
    .A(net622),
    .B(\mem.mem_internal.code_mem[63][0] ));
 sg13g2_nand2_1 _22686_ (.Y(_04588_),
    .A(net1022),
    .B(net439));
 sg13g2_o21ai_1 _22687_ (.B1(_04588_),
    .Y(_01834_),
    .A1(net439),
    .A2(_04587_));
 sg13g2_nand2_1 _22688_ (.Y(_04589_),
    .A(net622),
    .B(\mem.mem_internal.code_mem[63][1] ));
 sg13g2_nand2_1 _22689_ (.Y(_04590_),
    .A(net1021),
    .B(net439));
 sg13g2_o21ai_1 _22690_ (.B1(_04590_),
    .Y(_01835_),
    .A1(net439),
    .A2(_04589_));
 sg13g2_nand2_1 _22691_ (.Y(_04591_),
    .A(net622),
    .B(\mem.mem_internal.code_mem[63][2] ));
 sg13g2_nand2_1 _22692_ (.Y(_04592_),
    .A(net1020),
    .B(_04585_));
 sg13g2_o21ai_1 _22693_ (.B1(_04592_),
    .Y(_01836_),
    .A1(net439),
    .A2(_04591_));
 sg13g2_buf_1 _22694_ (.A(_04432_),
    .X(_04593_));
 sg13g2_nand2_1 _22695_ (.Y(_04594_),
    .A(net621),
    .B(\mem.mem_internal.code_mem[63][3] ));
 sg13g2_nand2_1 _22696_ (.Y(_04595_),
    .A(net1019),
    .B(_04585_));
 sg13g2_o21ai_1 _22697_ (.B1(_04595_),
    .Y(_01837_),
    .A1(net439),
    .A2(_04594_));
 sg13g2_nand2_1 _22698_ (.Y(_04596_),
    .A(net621),
    .B(\mem.mem_internal.code_mem[63][4] ));
 sg13g2_nand2_1 _22699_ (.Y(_04597_),
    .A(_04494_),
    .B(_04585_));
 sg13g2_o21ai_1 _22700_ (.B1(_04597_),
    .Y(_01838_),
    .A1(net439),
    .A2(_04596_));
 sg13g2_nand2_1 _22701_ (.Y(_04598_),
    .A(net621),
    .B(\mem.mem_internal.code_mem[63][5] ));
 sg13g2_nand2_1 _22702_ (.Y(_04599_),
    .A(_04497_),
    .B(_04585_));
 sg13g2_o21ai_1 _22703_ (.B1(_04599_),
    .Y(_01839_),
    .A1(net439),
    .A2(_04598_));
 sg13g2_nand2_1 _22704_ (.Y(_04600_),
    .A(net621),
    .B(\mem.mem_internal.code_mem[63][6] ));
 sg13g2_nand2_1 _22705_ (.Y(_04601_),
    .A(net1016),
    .B(_04585_));
 sg13g2_o21ai_1 _22706_ (.B1(_04601_),
    .Y(_01840_),
    .A1(_04586_),
    .A2(_04600_));
 sg13g2_nand2_1 _22707_ (.Y(_04602_),
    .A(net621),
    .B(\mem.mem_internal.code_mem[63][7] ));
 sg13g2_nand2_1 _22708_ (.Y(_04603_),
    .A(net1015),
    .B(_04585_));
 sg13g2_o21ai_1 _22709_ (.B1(_04603_),
    .Y(_01841_),
    .A1(_04586_),
    .A2(_04602_));
 sg13g2_nand2_1 _22710_ (.Y(_04604_),
    .A(net836),
    .B(\mem.mem_internal.code_mem[64][0] ));
 sg13g2_nand2_1 _22711_ (.Y(_04605_),
    .A(_10244_),
    .B(_10297_));
 sg13g2_buf_2 _22712_ (.A(_04605_),
    .X(_04606_));
 sg13g2_buf_1 _22713_ (.A(_04606_),
    .X(_04607_));
 sg13g2_nor2_1 _22714_ (.A(_10232_),
    .B(net457),
    .Y(_04608_));
 sg13g2_buf_2 _22715_ (.A(_04608_),
    .X(_04609_));
 sg13g2_buf_1 _22716_ (.A(_04609_),
    .X(_04610_));
 sg13g2_nand2_1 _22717_ (.Y(_04611_),
    .A(net1022),
    .B(net164));
 sg13g2_o21ai_1 _22718_ (.B1(_04611_),
    .Y(_01842_),
    .A1(_04604_),
    .A2(net164));
 sg13g2_nand2_1 _22719_ (.Y(_04612_),
    .A(_04593_),
    .B(\mem.mem_internal.code_mem[64][1] ));
 sg13g2_nand2_1 _22720_ (.Y(_04613_),
    .A(net1021),
    .B(net164));
 sg13g2_o21ai_1 _22721_ (.B1(_04613_),
    .Y(_01843_),
    .A1(net164),
    .A2(_04612_));
 sg13g2_nand2_1 _22722_ (.Y(_04614_),
    .A(_04593_),
    .B(\mem.mem_internal.code_mem[64][2] ));
 sg13g2_nand2_1 _22723_ (.Y(_04615_),
    .A(net1020),
    .B(_04609_));
 sg13g2_o21ai_1 _22724_ (.B1(_04615_),
    .Y(_01844_),
    .A1(net164),
    .A2(_04614_));
 sg13g2_nand2_1 _22725_ (.Y(_04616_),
    .A(net621),
    .B(\mem.mem_internal.code_mem[64][3] ));
 sg13g2_nand2_1 _22726_ (.Y(_04617_),
    .A(net1019),
    .B(_04609_));
 sg13g2_o21ai_1 _22727_ (.B1(_04617_),
    .Y(_01845_),
    .A1(net164),
    .A2(_04616_));
 sg13g2_nand2_1 _22728_ (.Y(_04618_),
    .A(net621),
    .B(\mem.mem_internal.code_mem[64][4] ));
 sg13g2_nand2_1 _22729_ (.Y(_04619_),
    .A(net1018),
    .B(_04609_));
 sg13g2_o21ai_1 _22730_ (.B1(_04619_),
    .Y(_01846_),
    .A1(_04610_),
    .A2(_04618_));
 sg13g2_nand2_1 _22731_ (.Y(_04620_),
    .A(net621),
    .B(\mem.mem_internal.code_mem[64][5] ));
 sg13g2_nand2_1 _22732_ (.Y(_04621_),
    .A(net1017),
    .B(_04609_));
 sg13g2_o21ai_1 _22733_ (.B1(_04621_),
    .Y(_01847_),
    .A1(_04610_),
    .A2(_04620_));
 sg13g2_buf_1 _22734_ (.A(_04431_),
    .X(_04622_));
 sg13g2_buf_1 _22735_ (.A(_04622_),
    .X(_04623_));
 sg13g2_nand2_1 _22736_ (.Y(_04624_),
    .A(net620),
    .B(\mem.mem_internal.code_mem[64][6] ));
 sg13g2_nand2_1 _22737_ (.Y(_04625_),
    .A(net1016),
    .B(_04609_));
 sg13g2_o21ai_1 _22738_ (.B1(_04625_),
    .Y(_01848_),
    .A1(net164),
    .A2(_04624_));
 sg13g2_nand2_1 _22739_ (.Y(_04626_),
    .A(net620),
    .B(\mem.mem_internal.code_mem[64][7] ));
 sg13g2_nand2_1 _22740_ (.Y(_04627_),
    .A(net1015),
    .B(_04609_));
 sg13g2_o21ai_1 _22741_ (.B1(_04627_),
    .Y(_01849_),
    .A1(net164),
    .A2(_04626_));
 sg13g2_nand2_1 _22742_ (.Y(_04628_),
    .A(net836),
    .B(\mem.mem_internal.code_mem[65][0] ));
 sg13g2_nor2_1 _22743_ (.A(_10632_),
    .B(net457),
    .Y(_04629_));
 sg13g2_buf_2 _22744_ (.A(_04629_),
    .X(_04630_));
 sg13g2_buf_1 _22745_ (.A(_04630_),
    .X(_04631_));
 sg13g2_nand2_1 _22746_ (.Y(_04632_),
    .A(net1022),
    .B(net163));
 sg13g2_o21ai_1 _22747_ (.B1(_04632_),
    .Y(_01850_),
    .A1(_04628_),
    .A2(net163));
 sg13g2_nand2_1 _22748_ (.Y(_04633_),
    .A(net620),
    .B(\mem.mem_internal.code_mem[65][1] ));
 sg13g2_nand2_1 _22749_ (.Y(_04634_),
    .A(net1021),
    .B(net163));
 sg13g2_o21ai_1 _22750_ (.B1(_04634_),
    .Y(_01851_),
    .A1(net163),
    .A2(_04633_));
 sg13g2_nand2_1 _22751_ (.Y(_04635_),
    .A(net620),
    .B(\mem.mem_internal.code_mem[65][2] ));
 sg13g2_nand2_1 _22752_ (.Y(_04636_),
    .A(net1020),
    .B(_04630_));
 sg13g2_o21ai_1 _22753_ (.B1(_04636_),
    .Y(_01852_),
    .A1(net163),
    .A2(_04635_));
 sg13g2_nand2_1 _22754_ (.Y(_04637_),
    .A(net620),
    .B(\mem.mem_internal.code_mem[65][3] ));
 sg13g2_nand2_1 _22755_ (.Y(_04638_),
    .A(net1019),
    .B(_04630_));
 sg13g2_o21ai_1 _22756_ (.B1(_04638_),
    .Y(_01853_),
    .A1(net163),
    .A2(_04637_));
 sg13g2_nand2_1 _22757_ (.Y(_04639_),
    .A(net620),
    .B(\mem.mem_internal.code_mem[65][4] ));
 sg13g2_nand2_1 _22758_ (.Y(_04640_),
    .A(net1018),
    .B(_04630_));
 sg13g2_o21ai_1 _22759_ (.B1(_04640_),
    .Y(_01854_),
    .A1(net163),
    .A2(_04639_));
 sg13g2_nand2_1 _22760_ (.Y(_04641_),
    .A(_04623_),
    .B(\mem.mem_internal.code_mem[65][5] ));
 sg13g2_nand2_1 _22761_ (.Y(_04642_),
    .A(net1017),
    .B(_04630_));
 sg13g2_o21ai_1 _22762_ (.B1(_04642_),
    .Y(_01855_),
    .A1(_04631_),
    .A2(_04641_));
 sg13g2_nand2_1 _22763_ (.Y(_04643_),
    .A(_04623_),
    .B(\mem.mem_internal.code_mem[65][6] ));
 sg13g2_nand2_1 _22764_ (.Y(_04644_),
    .A(net1016),
    .B(_04630_));
 sg13g2_o21ai_1 _22765_ (.B1(_04644_),
    .Y(_01856_),
    .A1(_04631_),
    .A2(_04643_));
 sg13g2_nand2_1 _22766_ (.Y(_04645_),
    .A(net620),
    .B(\mem.mem_internal.code_mem[65][7] ));
 sg13g2_nand2_1 _22767_ (.Y(_04646_),
    .A(net1015),
    .B(_04630_));
 sg13g2_o21ai_1 _22768_ (.B1(_04646_),
    .Y(_01857_),
    .A1(net163),
    .A2(_04645_));
 sg13g2_nand2_1 _22769_ (.Y(_04647_),
    .A(net836),
    .B(\mem.mem_internal.code_mem[66][0] ));
 sg13g2_nor2_1 _22770_ (.A(_10656_),
    .B(net457),
    .Y(_04648_));
 sg13g2_buf_2 _22771_ (.A(_04648_),
    .X(_04649_));
 sg13g2_buf_1 _22772_ (.A(_04649_),
    .X(_04650_));
 sg13g2_nand2_1 _22773_ (.Y(_04651_),
    .A(_04481_),
    .B(net162));
 sg13g2_o21ai_1 _22774_ (.B1(_04651_),
    .Y(_01858_),
    .A1(_04647_),
    .A2(net162));
 sg13g2_nand2_1 _22775_ (.Y(_04652_),
    .A(net620),
    .B(\mem.mem_internal.code_mem[66][1] ));
 sg13g2_nand2_1 _22776_ (.Y(_04653_),
    .A(_04484_),
    .B(net162));
 sg13g2_o21ai_1 _22777_ (.B1(_04653_),
    .Y(_01859_),
    .A1(net162),
    .A2(_04652_));
 sg13g2_buf_1 _22778_ (.A(_04622_),
    .X(_04654_));
 sg13g2_nand2_1 _22779_ (.Y(_04655_),
    .A(net619),
    .B(\mem.mem_internal.code_mem[66][2] ));
 sg13g2_nand2_1 _22780_ (.Y(_04656_),
    .A(_04488_),
    .B(_04649_));
 sg13g2_o21ai_1 _22781_ (.B1(_04656_),
    .Y(_01860_),
    .A1(net162),
    .A2(_04655_));
 sg13g2_nand2_1 _22782_ (.Y(_04657_),
    .A(_04654_),
    .B(\mem.mem_internal.code_mem[66][3] ));
 sg13g2_nand2_1 _22783_ (.Y(_04658_),
    .A(_04491_),
    .B(_04649_));
 sg13g2_o21ai_1 _22784_ (.B1(_04658_),
    .Y(_01861_),
    .A1(net162),
    .A2(_04657_));
 sg13g2_nand2_1 _22785_ (.Y(_04659_),
    .A(net619),
    .B(\mem.mem_internal.code_mem[66][4] ));
 sg13g2_nand2_1 _22786_ (.Y(_04660_),
    .A(net1018),
    .B(_04649_));
 sg13g2_o21ai_1 _22787_ (.B1(_04660_),
    .Y(_01862_),
    .A1(net162),
    .A2(_04659_));
 sg13g2_nand2_1 _22788_ (.Y(_04661_),
    .A(net619),
    .B(\mem.mem_internal.code_mem[66][5] ));
 sg13g2_nand2_1 _22789_ (.Y(_04662_),
    .A(net1017),
    .B(_04649_));
 sg13g2_o21ai_1 _22790_ (.B1(_04662_),
    .Y(_01863_),
    .A1(_04650_),
    .A2(_04661_));
 sg13g2_nand2_1 _22791_ (.Y(_04663_),
    .A(_04654_),
    .B(\mem.mem_internal.code_mem[66][6] ));
 sg13g2_nand2_1 _22792_ (.Y(_04664_),
    .A(_04500_),
    .B(_04649_));
 sg13g2_o21ai_1 _22793_ (.B1(_04664_),
    .Y(_01864_),
    .A1(_04650_),
    .A2(_04663_));
 sg13g2_nand2_1 _22794_ (.Y(_04665_),
    .A(net619),
    .B(\mem.mem_internal.code_mem[66][7] ));
 sg13g2_nand2_1 _22795_ (.Y(_04666_),
    .A(_04503_),
    .B(_04649_));
 sg13g2_o21ai_1 _22796_ (.B1(_04666_),
    .Y(_01865_),
    .A1(net162),
    .A2(_04665_));
 sg13g2_nand2_1 _22797_ (.Y(_04667_),
    .A(net836),
    .B(\mem.mem_internal.code_mem[67][0] ));
 sg13g2_nor2_1 _22798_ (.A(_10679_),
    .B(net457),
    .Y(_04668_));
 sg13g2_buf_2 _22799_ (.A(_04668_),
    .X(_04669_));
 sg13g2_buf_1 _22800_ (.A(_04669_),
    .X(_04670_));
 sg13g2_nand2_1 _22801_ (.Y(_04671_),
    .A(_04481_),
    .B(net161));
 sg13g2_o21ai_1 _22802_ (.B1(_04671_),
    .Y(_01866_),
    .A1(_04667_),
    .A2(net161));
 sg13g2_nand2_1 _22803_ (.Y(_04672_),
    .A(net619),
    .B(\mem.mem_internal.code_mem[67][1] ));
 sg13g2_nand2_1 _22804_ (.Y(_04673_),
    .A(_04484_),
    .B(net161));
 sg13g2_o21ai_1 _22805_ (.B1(_04673_),
    .Y(_01867_),
    .A1(net161),
    .A2(_04672_));
 sg13g2_nand2_1 _22806_ (.Y(_04674_),
    .A(net619),
    .B(\mem.mem_internal.code_mem[67][2] ));
 sg13g2_nand2_1 _22807_ (.Y(_04675_),
    .A(net1020),
    .B(_04669_));
 sg13g2_o21ai_1 _22808_ (.B1(_04675_),
    .Y(_01868_),
    .A1(net161),
    .A2(_04674_));
 sg13g2_nand2_1 _22809_ (.Y(_04676_),
    .A(net619),
    .B(\mem.mem_internal.code_mem[67][3] ));
 sg13g2_nand2_1 _22810_ (.Y(_04677_),
    .A(net1019),
    .B(_04669_));
 sg13g2_o21ai_1 _22811_ (.B1(_04677_),
    .Y(_01869_),
    .A1(net161),
    .A2(_04676_));
 sg13g2_nand2_1 _22812_ (.Y(_04678_),
    .A(net619),
    .B(\mem.mem_internal.code_mem[67][4] ));
 sg13g2_nand2_1 _22813_ (.Y(_04679_),
    .A(net1018),
    .B(_04669_));
 sg13g2_o21ai_1 _22814_ (.B1(_04679_),
    .Y(_01870_),
    .A1(net161),
    .A2(_04678_));
 sg13g2_buf_1 _22815_ (.A(_04622_),
    .X(_04680_));
 sg13g2_nand2_1 _22816_ (.Y(_04681_),
    .A(net618),
    .B(\mem.mem_internal.code_mem[67][5] ));
 sg13g2_nand2_1 _22817_ (.Y(_04682_),
    .A(net1017),
    .B(_04669_));
 sg13g2_o21ai_1 _22818_ (.B1(_04682_),
    .Y(_01871_),
    .A1(_04670_),
    .A2(_04681_));
 sg13g2_nand2_1 _22819_ (.Y(_04683_),
    .A(net618),
    .B(\mem.mem_internal.code_mem[67][6] ));
 sg13g2_nand2_1 _22820_ (.Y(_04684_),
    .A(_04500_),
    .B(_04669_));
 sg13g2_o21ai_1 _22821_ (.B1(_04684_),
    .Y(_01872_),
    .A1(_04670_),
    .A2(_04683_));
 sg13g2_nand2_1 _22822_ (.Y(_04685_),
    .A(net618),
    .B(\mem.mem_internal.code_mem[67][7] ));
 sg13g2_nand2_1 _22823_ (.Y(_04686_),
    .A(_04503_),
    .B(_04669_));
 sg13g2_o21ai_1 _22824_ (.B1(_04686_),
    .Y(_01873_),
    .A1(net161),
    .A2(_04685_));
 sg13g2_nand2_1 _22825_ (.Y(_04687_),
    .A(net836),
    .B(\mem.mem_internal.code_mem[68][0] ));
 sg13g2_nor2_1 _22826_ (.A(_10295_),
    .B(net457),
    .Y(_04688_));
 sg13g2_buf_2 _22827_ (.A(_04688_),
    .X(_04689_));
 sg13g2_buf_1 _22828_ (.A(_04689_),
    .X(_04690_));
 sg13g2_buf_1 _22829_ (.A(_03842_),
    .X(_04691_));
 sg13g2_nand2_1 _22830_ (.Y(_04692_),
    .A(net1014),
    .B(net160));
 sg13g2_o21ai_1 _22831_ (.B1(_04692_),
    .Y(_01874_),
    .A1(_04687_),
    .A2(net160));
 sg13g2_nand2_1 _22832_ (.Y(_04693_),
    .A(net618),
    .B(\mem.mem_internal.code_mem[68][1] ));
 sg13g2_buf_1 _22833_ (.A(_03846_),
    .X(_04694_));
 sg13g2_nand2_1 _22834_ (.Y(_04695_),
    .A(net1013),
    .B(net160));
 sg13g2_o21ai_1 _22835_ (.B1(_04695_),
    .Y(_01875_),
    .A1(net160),
    .A2(_04693_));
 sg13g2_nand2_1 _22836_ (.Y(_04696_),
    .A(net618),
    .B(\mem.mem_internal.code_mem[68][2] ));
 sg13g2_buf_1 _22837_ (.A(_03850_),
    .X(_04697_));
 sg13g2_nand2_1 _22838_ (.Y(_04698_),
    .A(net1012),
    .B(_04689_));
 sg13g2_o21ai_1 _22839_ (.B1(_04698_),
    .Y(_01876_),
    .A1(net160),
    .A2(_04696_));
 sg13g2_nand2_1 _22840_ (.Y(_04699_),
    .A(net618),
    .B(\mem.mem_internal.code_mem[68][3] ));
 sg13g2_buf_1 _22841_ (.A(_03854_),
    .X(_04700_));
 sg13g2_nand2_1 _22842_ (.Y(_04701_),
    .A(net1011),
    .B(_04689_));
 sg13g2_o21ai_1 _22843_ (.B1(_04701_),
    .Y(_01877_),
    .A1(net160),
    .A2(_04699_));
 sg13g2_nand2_1 _22844_ (.Y(_04702_),
    .A(net618),
    .B(\mem.mem_internal.code_mem[68][4] ));
 sg13g2_buf_1 _22845_ (.A(_03859_),
    .X(_04703_));
 sg13g2_nand2_1 _22846_ (.Y(_04704_),
    .A(net1010),
    .B(_04689_));
 sg13g2_o21ai_1 _22847_ (.B1(_04704_),
    .Y(_01878_),
    .A1(net160),
    .A2(_04702_));
 sg13g2_nand2_1 _22848_ (.Y(_04705_),
    .A(_04680_),
    .B(\mem.mem_internal.code_mem[68][5] ));
 sg13g2_buf_1 _22849_ (.A(_03863_),
    .X(_04706_));
 sg13g2_nand2_1 _22850_ (.Y(_04707_),
    .A(net1009),
    .B(_04689_));
 sg13g2_o21ai_1 _22851_ (.B1(_04707_),
    .Y(_01879_),
    .A1(_04690_),
    .A2(_04705_));
 sg13g2_nand2_1 _22852_ (.Y(_04708_),
    .A(_04680_),
    .B(\mem.mem_internal.code_mem[68][6] ));
 sg13g2_buf_1 _22853_ (.A(_03867_),
    .X(_04709_));
 sg13g2_nand2_1 _22854_ (.Y(_04710_),
    .A(net1008),
    .B(_04689_));
 sg13g2_o21ai_1 _22855_ (.B1(_04710_),
    .Y(_01880_),
    .A1(_04690_),
    .A2(_04708_));
 sg13g2_nand2_1 _22856_ (.Y(_04711_),
    .A(net618),
    .B(\mem.mem_internal.code_mem[68][7] ));
 sg13g2_buf_1 _22857_ (.A(_03871_),
    .X(_04712_));
 sg13g2_nand2_1 _22858_ (.Y(_04713_),
    .A(net1007),
    .B(_04689_));
 sg13g2_o21ai_1 _22859_ (.B1(_04713_),
    .Y(_01881_),
    .A1(net160),
    .A2(_04711_));
 sg13g2_nand2_1 _22860_ (.Y(_04714_),
    .A(net836),
    .B(\mem.mem_internal.code_mem[69][0] ));
 sg13g2_nor2_1 _22861_ (.A(_10325_),
    .B(_04607_),
    .Y(_04715_));
 sg13g2_buf_2 _22862_ (.A(_04715_),
    .X(_04716_));
 sg13g2_buf_1 _22863_ (.A(_04716_),
    .X(_04717_));
 sg13g2_nand2_1 _22864_ (.Y(_04718_),
    .A(net1014),
    .B(net159));
 sg13g2_o21ai_1 _22865_ (.B1(_04718_),
    .Y(_01882_),
    .A1(_04714_),
    .A2(net159));
 sg13g2_buf_1 _22866_ (.A(_04622_),
    .X(_04719_));
 sg13g2_nand2_1 _22867_ (.Y(_04720_),
    .A(net617),
    .B(\mem.mem_internal.code_mem[69][1] ));
 sg13g2_nand2_1 _22868_ (.Y(_04721_),
    .A(net1013),
    .B(net159));
 sg13g2_o21ai_1 _22869_ (.B1(_04721_),
    .Y(_01883_),
    .A1(net159),
    .A2(_04720_));
 sg13g2_nand2_1 _22870_ (.Y(_04722_),
    .A(net617),
    .B(\mem.mem_internal.code_mem[69][2] ));
 sg13g2_nand2_1 _22871_ (.Y(_04723_),
    .A(net1012),
    .B(_04716_));
 sg13g2_o21ai_1 _22872_ (.B1(_04723_),
    .Y(_01884_),
    .A1(net159),
    .A2(_04722_));
 sg13g2_nand2_1 _22873_ (.Y(_04724_),
    .A(net617),
    .B(\mem.mem_internal.code_mem[69][3] ));
 sg13g2_nand2_1 _22874_ (.Y(_04725_),
    .A(net1011),
    .B(_04716_));
 sg13g2_o21ai_1 _22875_ (.B1(_04725_),
    .Y(_01885_),
    .A1(net159),
    .A2(_04724_));
 sg13g2_nand2_1 _22876_ (.Y(_04726_),
    .A(net617),
    .B(\mem.mem_internal.code_mem[69][4] ));
 sg13g2_nand2_1 _22877_ (.Y(_04727_),
    .A(net1010),
    .B(_04716_));
 sg13g2_o21ai_1 _22878_ (.B1(_04727_),
    .Y(_01886_),
    .A1(net159),
    .A2(_04726_));
 sg13g2_nand2_1 _22879_ (.Y(_04728_),
    .A(_04719_),
    .B(\mem.mem_internal.code_mem[69][5] ));
 sg13g2_nand2_1 _22880_ (.Y(_04729_),
    .A(net1009),
    .B(_04716_));
 sg13g2_o21ai_1 _22881_ (.B1(_04729_),
    .Y(_01887_),
    .A1(_04717_),
    .A2(_04728_));
 sg13g2_nand2_1 _22882_ (.Y(_04730_),
    .A(_04719_),
    .B(\mem.mem_internal.code_mem[69][6] ));
 sg13g2_nand2_1 _22883_ (.Y(_04731_),
    .A(net1008),
    .B(_04716_));
 sg13g2_o21ai_1 _22884_ (.B1(_04731_),
    .Y(_01888_),
    .A1(_04717_),
    .A2(_04730_));
 sg13g2_nand2_1 _22885_ (.Y(_04732_),
    .A(net617),
    .B(\mem.mem_internal.code_mem[69][7] ));
 sg13g2_nand2_1 _22886_ (.Y(_04733_),
    .A(net1007),
    .B(_04716_));
 sg13g2_o21ai_1 _22887_ (.B1(_04733_),
    .Y(_01889_),
    .A1(net159),
    .A2(_04732_));
 sg13g2_nand2_1 _22888_ (.Y(_04734_),
    .A(_04202_),
    .B(\mem.mem_internal.code_mem[6][0] ));
 sg13g2_nor2_1 _22889_ (.A(_10246_),
    .B(net554),
    .Y(_04735_));
 sg13g2_buf_2 _22890_ (.A(_04735_),
    .X(_04736_));
 sg13g2_buf_1 _22891_ (.A(_04736_),
    .X(_04737_));
 sg13g2_nand2_1 _22892_ (.Y(_04738_),
    .A(net1014),
    .B(net318));
 sg13g2_o21ai_1 _22893_ (.B1(_04738_),
    .Y(_01890_),
    .A1(_04734_),
    .A2(net318));
 sg13g2_nand2_1 _22894_ (.Y(_04739_),
    .A(net617),
    .B(\mem.mem_internal.code_mem[6][1] ));
 sg13g2_nand2_1 _22895_ (.Y(_04740_),
    .A(net1013),
    .B(net318));
 sg13g2_o21ai_1 _22896_ (.B1(_04740_),
    .Y(_01891_),
    .A1(net318),
    .A2(_04739_));
 sg13g2_nand2_1 _22897_ (.Y(_04741_),
    .A(net617),
    .B(\mem.mem_internal.code_mem[6][2] ));
 sg13g2_nand2_1 _22898_ (.Y(_04742_),
    .A(net1012),
    .B(_04736_));
 sg13g2_o21ai_1 _22899_ (.B1(_04742_),
    .Y(_01892_),
    .A1(_04737_),
    .A2(_04741_));
 sg13g2_nand2_1 _22900_ (.Y(_04743_),
    .A(net617),
    .B(\mem.mem_internal.code_mem[6][3] ));
 sg13g2_nand2_1 _22901_ (.Y(_04744_),
    .A(net1011),
    .B(_04736_));
 sg13g2_o21ai_1 _22902_ (.B1(_04744_),
    .Y(_01893_),
    .A1(_04737_),
    .A2(_04743_));
 sg13g2_buf_1 _22903_ (.A(_04622_),
    .X(_04745_));
 sg13g2_nand2_1 _22904_ (.Y(_04746_),
    .A(net616),
    .B(\mem.mem_internal.code_mem[6][4] ));
 sg13g2_nand2_1 _22905_ (.Y(_04747_),
    .A(net1010),
    .B(_04736_));
 sg13g2_o21ai_1 _22906_ (.B1(_04747_),
    .Y(_01894_),
    .A1(net318),
    .A2(_04746_));
 sg13g2_nand2_1 _22907_ (.Y(_04748_),
    .A(net616),
    .B(\mem.mem_internal.code_mem[6][5] ));
 sg13g2_nand2_1 _22908_ (.Y(_04749_),
    .A(net1009),
    .B(_04736_));
 sg13g2_o21ai_1 _22909_ (.B1(_04749_),
    .Y(_01895_),
    .A1(net318),
    .A2(_04748_));
 sg13g2_nand2_1 _22910_ (.Y(_04750_),
    .A(net616),
    .B(\mem.mem_internal.code_mem[6][6] ));
 sg13g2_nand2_1 _22911_ (.Y(_04751_),
    .A(net1008),
    .B(_04736_));
 sg13g2_o21ai_1 _22912_ (.B1(_04751_),
    .Y(_01896_),
    .A1(net318),
    .A2(_04750_));
 sg13g2_nand2_1 _22913_ (.Y(_04752_),
    .A(net616),
    .B(\mem.mem_internal.code_mem[6][7] ));
 sg13g2_nand2_1 _22914_ (.Y(_04753_),
    .A(net1007),
    .B(_04736_));
 sg13g2_o21ai_1 _22915_ (.B1(_04753_),
    .Y(_01897_),
    .A1(net318),
    .A2(_04752_));
 sg13g2_buf_1 _22916_ (.A(net1192),
    .X(_04754_));
 sg13g2_nand2_1 _22917_ (.Y(_04755_),
    .A(net835),
    .B(\mem.mem_internal.code_mem[70][0] ));
 sg13g2_nor2_1 _22918_ (.A(net779),
    .B(net457),
    .Y(_04756_));
 sg13g2_buf_2 _22919_ (.A(_04756_),
    .X(_04757_));
 sg13g2_buf_1 _22920_ (.A(_04757_),
    .X(_04758_));
 sg13g2_nand2_1 _22921_ (.Y(_04759_),
    .A(net1014),
    .B(net158));
 sg13g2_o21ai_1 _22922_ (.B1(_04759_),
    .Y(_01898_),
    .A1(_04755_),
    .A2(net158));
 sg13g2_nand2_1 _22923_ (.Y(_04760_),
    .A(net616),
    .B(\mem.mem_internal.code_mem[70][1] ));
 sg13g2_nand2_1 _22924_ (.Y(_04761_),
    .A(net1013),
    .B(net158));
 sg13g2_o21ai_1 _22925_ (.B1(_04761_),
    .Y(_01899_),
    .A1(net158),
    .A2(_04760_));
 sg13g2_nand2_1 _22926_ (.Y(_04762_),
    .A(net616),
    .B(\mem.mem_internal.code_mem[70][2] ));
 sg13g2_nand2_1 _22927_ (.Y(_04763_),
    .A(net1012),
    .B(_04757_));
 sg13g2_o21ai_1 _22928_ (.B1(_04763_),
    .Y(_01900_),
    .A1(net158),
    .A2(_04762_));
 sg13g2_nand2_1 _22929_ (.Y(_04764_),
    .A(net616),
    .B(\mem.mem_internal.code_mem[70][3] ));
 sg13g2_nand2_1 _22930_ (.Y(_04765_),
    .A(net1011),
    .B(_04757_));
 sg13g2_o21ai_1 _22931_ (.B1(_04765_),
    .Y(_01901_),
    .A1(net158),
    .A2(_04764_));
 sg13g2_nand2_1 _22932_ (.Y(_04766_),
    .A(net616),
    .B(\mem.mem_internal.code_mem[70][4] ));
 sg13g2_nand2_1 _22933_ (.Y(_04767_),
    .A(net1010),
    .B(_04757_));
 sg13g2_o21ai_1 _22934_ (.B1(_04767_),
    .Y(_01902_),
    .A1(_04758_),
    .A2(_04766_));
 sg13g2_nand2_1 _22935_ (.Y(_04768_),
    .A(_04745_),
    .B(\mem.mem_internal.code_mem[70][5] ));
 sg13g2_nand2_1 _22936_ (.Y(_04769_),
    .A(net1009),
    .B(_04757_));
 sg13g2_o21ai_1 _22937_ (.B1(_04769_),
    .Y(_01903_),
    .A1(_04758_),
    .A2(_04768_));
 sg13g2_nand2_1 _22938_ (.Y(_04770_),
    .A(_04745_),
    .B(\mem.mem_internal.code_mem[70][6] ));
 sg13g2_nand2_1 _22939_ (.Y(_04771_),
    .A(net1008),
    .B(_04757_));
 sg13g2_o21ai_1 _22940_ (.B1(_04771_),
    .Y(_01904_),
    .A1(net158),
    .A2(_04770_));
 sg13g2_buf_1 _22941_ (.A(_04622_),
    .X(_04772_));
 sg13g2_nand2_1 _22942_ (.Y(_04773_),
    .A(net615),
    .B(\mem.mem_internal.code_mem[70][7] ));
 sg13g2_nand2_1 _22943_ (.Y(_04774_),
    .A(net1007),
    .B(_04757_));
 sg13g2_o21ai_1 _22944_ (.B1(_04774_),
    .Y(_01905_),
    .A1(net158),
    .A2(_04773_));
 sg13g2_nand2_1 _22945_ (.Y(_04775_),
    .A(net835),
    .B(\mem.mem_internal.code_mem[71][0] ));
 sg13g2_nor2_1 _22946_ (.A(_10372_),
    .B(net457),
    .Y(_04776_));
 sg13g2_buf_2 _22947_ (.A(_04776_),
    .X(_04777_));
 sg13g2_buf_1 _22948_ (.A(_04777_),
    .X(_04778_));
 sg13g2_nand2_1 _22949_ (.Y(_04779_),
    .A(net1014),
    .B(net157));
 sg13g2_o21ai_1 _22950_ (.B1(_04779_),
    .Y(_01906_),
    .A1(_04775_),
    .A2(net157));
 sg13g2_nand2_1 _22951_ (.Y(_04780_),
    .A(net615),
    .B(\mem.mem_internal.code_mem[71][1] ));
 sg13g2_nand2_1 _22952_ (.Y(_04781_),
    .A(net1013),
    .B(net157));
 sg13g2_o21ai_1 _22953_ (.B1(_04781_),
    .Y(_01907_),
    .A1(net157),
    .A2(_04780_));
 sg13g2_nand2_1 _22954_ (.Y(_04782_),
    .A(net615),
    .B(\mem.mem_internal.code_mem[71][2] ));
 sg13g2_nand2_1 _22955_ (.Y(_04783_),
    .A(net1012),
    .B(_04777_));
 sg13g2_o21ai_1 _22956_ (.B1(_04783_),
    .Y(_01908_),
    .A1(net157),
    .A2(_04782_));
 sg13g2_nand2_1 _22957_ (.Y(_04784_),
    .A(net615),
    .B(\mem.mem_internal.code_mem[71][3] ));
 sg13g2_nand2_1 _22958_ (.Y(_04785_),
    .A(net1011),
    .B(_04777_));
 sg13g2_o21ai_1 _22959_ (.B1(_04785_),
    .Y(_01909_),
    .A1(net157),
    .A2(_04784_));
 sg13g2_nand2_1 _22960_ (.Y(_04786_),
    .A(net615),
    .B(\mem.mem_internal.code_mem[71][4] ));
 sg13g2_nand2_1 _22961_ (.Y(_04787_),
    .A(net1010),
    .B(_04777_));
 sg13g2_o21ai_1 _22962_ (.B1(_04787_),
    .Y(_01910_),
    .A1(net157),
    .A2(_04786_));
 sg13g2_nand2_1 _22963_ (.Y(_04788_),
    .A(_04772_),
    .B(\mem.mem_internal.code_mem[71][5] ));
 sg13g2_nand2_1 _22964_ (.Y(_04789_),
    .A(net1009),
    .B(_04777_));
 sg13g2_o21ai_1 _22965_ (.B1(_04789_),
    .Y(_01911_),
    .A1(_04778_),
    .A2(_04788_));
 sg13g2_nand2_1 _22966_ (.Y(_04790_),
    .A(_04772_),
    .B(\mem.mem_internal.code_mem[71][6] ));
 sg13g2_nand2_1 _22967_ (.Y(_04791_),
    .A(net1008),
    .B(_04777_));
 sg13g2_o21ai_1 _22968_ (.B1(_04791_),
    .Y(_01912_),
    .A1(_04778_),
    .A2(_04790_));
 sg13g2_nand2_1 _22969_ (.Y(_04792_),
    .A(net615),
    .B(\mem.mem_internal.code_mem[71][7] ));
 sg13g2_nand2_1 _22970_ (.Y(_04793_),
    .A(net1007),
    .B(_04777_));
 sg13g2_o21ai_1 _22971_ (.B1(_04793_),
    .Y(_01913_),
    .A1(net157),
    .A2(_04792_));
 sg13g2_nand2_1 _22972_ (.Y(_04794_),
    .A(net835),
    .B(\mem.mem_internal.code_mem[72][0] ));
 sg13g2_nor2_1 _22973_ (.A(net778),
    .B(net457),
    .Y(_04795_));
 sg13g2_buf_2 _22974_ (.A(_04795_),
    .X(_04796_));
 sg13g2_buf_1 _22975_ (.A(_04796_),
    .X(_04797_));
 sg13g2_nand2_1 _22976_ (.Y(_04798_),
    .A(_04691_),
    .B(net156));
 sg13g2_o21ai_1 _22977_ (.B1(_04798_),
    .Y(_01914_),
    .A1(_04794_),
    .A2(net156));
 sg13g2_nand2_1 _22978_ (.Y(_04799_),
    .A(net615),
    .B(\mem.mem_internal.code_mem[72][1] ));
 sg13g2_nand2_1 _22979_ (.Y(_04800_),
    .A(net1013),
    .B(net156));
 sg13g2_o21ai_1 _22980_ (.B1(_04800_),
    .Y(_01915_),
    .A1(net156),
    .A2(_04799_));
 sg13g2_nand2_1 _22981_ (.Y(_04801_),
    .A(net615),
    .B(\mem.mem_internal.code_mem[72][2] ));
 sg13g2_nand2_1 _22982_ (.Y(_04802_),
    .A(net1012),
    .B(_04796_));
 sg13g2_o21ai_1 _22983_ (.B1(_04802_),
    .Y(_01916_),
    .A1(net156),
    .A2(_04801_));
 sg13g2_buf_1 _22984_ (.A(_04622_),
    .X(_04803_));
 sg13g2_nand2_1 _22985_ (.Y(_04804_),
    .A(_04803_),
    .B(\mem.mem_internal.code_mem[72][3] ));
 sg13g2_nand2_1 _22986_ (.Y(_04805_),
    .A(_04700_),
    .B(_04796_));
 sg13g2_o21ai_1 _22987_ (.B1(_04805_),
    .Y(_01917_),
    .A1(net156),
    .A2(_04804_));
 sg13g2_nand2_1 _22988_ (.Y(_04806_),
    .A(net614),
    .B(\mem.mem_internal.code_mem[72][4] ));
 sg13g2_nand2_1 _22989_ (.Y(_04807_),
    .A(_04703_),
    .B(_04796_));
 sg13g2_o21ai_1 _22990_ (.B1(_04807_),
    .Y(_01918_),
    .A1(net156),
    .A2(_04806_));
 sg13g2_nand2_1 _22991_ (.Y(_04808_),
    .A(net614),
    .B(\mem.mem_internal.code_mem[72][5] ));
 sg13g2_nand2_1 _22992_ (.Y(_04809_),
    .A(_04706_),
    .B(_04796_));
 sg13g2_o21ai_1 _22993_ (.B1(_04809_),
    .Y(_01919_),
    .A1(_04797_),
    .A2(_04808_));
 sg13g2_nand2_1 _22994_ (.Y(_04810_),
    .A(_04803_),
    .B(\mem.mem_internal.code_mem[72][6] ));
 sg13g2_nand2_1 _22995_ (.Y(_04811_),
    .A(net1008),
    .B(_04796_));
 sg13g2_o21ai_1 _22996_ (.B1(_04811_),
    .Y(_01920_),
    .A1(_04797_),
    .A2(_04810_));
 sg13g2_nand2_1 _22997_ (.Y(_04812_),
    .A(net614),
    .B(\mem.mem_internal.code_mem[72][7] ));
 sg13g2_nand2_1 _22998_ (.Y(_04813_),
    .A(net1007),
    .B(_04796_));
 sg13g2_o21ai_1 _22999_ (.B1(_04813_),
    .Y(_01921_),
    .A1(net156),
    .A2(_04812_));
 sg13g2_nand2_1 _23000_ (.Y(_04814_),
    .A(net835),
    .B(\mem.mem_internal.code_mem[73][0] ));
 sg13g2_nor2_1 _23001_ (.A(_10422_),
    .B(_04607_),
    .Y(_04815_));
 sg13g2_buf_2 _23002_ (.A(_04815_),
    .X(_04816_));
 sg13g2_buf_1 _23003_ (.A(_04816_),
    .X(_04817_));
 sg13g2_nand2_1 _23004_ (.Y(_04818_),
    .A(net1014),
    .B(net155));
 sg13g2_o21ai_1 _23005_ (.B1(_04818_),
    .Y(_01922_),
    .A1(_04814_),
    .A2(net155));
 sg13g2_nand2_1 _23006_ (.Y(_04819_),
    .A(net614),
    .B(\mem.mem_internal.code_mem[73][1] ));
 sg13g2_nand2_1 _23007_ (.Y(_04820_),
    .A(net1013),
    .B(net155));
 sg13g2_o21ai_1 _23008_ (.B1(_04820_),
    .Y(_01923_),
    .A1(net155),
    .A2(_04819_));
 sg13g2_nand2_1 _23009_ (.Y(_04821_),
    .A(net614),
    .B(\mem.mem_internal.code_mem[73][2] ));
 sg13g2_nand2_1 _23010_ (.Y(_04822_),
    .A(net1012),
    .B(_04816_));
 sg13g2_o21ai_1 _23011_ (.B1(_04822_),
    .Y(_01924_),
    .A1(net155),
    .A2(_04821_));
 sg13g2_nand2_1 _23012_ (.Y(_04823_),
    .A(net614),
    .B(\mem.mem_internal.code_mem[73][3] ));
 sg13g2_nand2_1 _23013_ (.Y(_04824_),
    .A(net1011),
    .B(_04816_));
 sg13g2_o21ai_1 _23014_ (.B1(_04824_),
    .Y(_01925_),
    .A1(net155),
    .A2(_04823_));
 sg13g2_nand2_1 _23015_ (.Y(_04825_),
    .A(net614),
    .B(\mem.mem_internal.code_mem[73][4] ));
 sg13g2_nand2_1 _23016_ (.Y(_04826_),
    .A(net1010),
    .B(_04816_));
 sg13g2_o21ai_1 _23017_ (.B1(_04826_),
    .Y(_01926_),
    .A1(net155),
    .A2(_04825_));
 sg13g2_nand2_1 _23018_ (.Y(_04827_),
    .A(net614),
    .B(\mem.mem_internal.code_mem[73][5] ));
 sg13g2_nand2_1 _23019_ (.Y(_04828_),
    .A(net1009),
    .B(_04816_));
 sg13g2_o21ai_1 _23020_ (.B1(_04828_),
    .Y(_01927_),
    .A1(net155),
    .A2(_04827_));
 sg13g2_buf_1 _23021_ (.A(_04431_),
    .X(_04829_));
 sg13g2_buf_1 _23022_ (.A(_04829_),
    .X(_04830_));
 sg13g2_nand2_1 _23023_ (.Y(_04831_),
    .A(_04830_),
    .B(\mem.mem_internal.code_mem[73][6] ));
 sg13g2_nand2_1 _23024_ (.Y(_04832_),
    .A(net1008),
    .B(_04816_));
 sg13g2_o21ai_1 _23025_ (.B1(_04832_),
    .Y(_01928_),
    .A1(_04817_),
    .A2(_04831_));
 sg13g2_nand2_1 _23026_ (.Y(_04833_),
    .A(net613),
    .B(\mem.mem_internal.code_mem[73][7] ));
 sg13g2_nand2_1 _23027_ (.Y(_04834_),
    .A(net1007),
    .B(_04816_));
 sg13g2_o21ai_1 _23028_ (.B1(_04834_),
    .Y(_01929_),
    .A1(_04817_),
    .A2(_04833_));
 sg13g2_nand2_1 _23029_ (.Y(_04835_),
    .A(net835),
    .B(\mem.mem_internal.code_mem[74][0] ));
 sg13g2_nor2_1 _23030_ (.A(_10444_),
    .B(_04606_),
    .Y(_04836_));
 sg13g2_buf_2 _23031_ (.A(_04836_),
    .X(_04837_));
 sg13g2_buf_1 _23032_ (.A(_04837_),
    .X(_04838_));
 sg13g2_nand2_1 _23033_ (.Y(_04839_),
    .A(net1014),
    .B(net317));
 sg13g2_o21ai_1 _23034_ (.B1(_04839_),
    .Y(_01930_),
    .A1(_04835_),
    .A2(net317));
 sg13g2_nand2_1 _23035_ (.Y(_04840_),
    .A(net613),
    .B(\mem.mem_internal.code_mem[74][1] ));
 sg13g2_nand2_1 _23036_ (.Y(_04841_),
    .A(net1013),
    .B(net317));
 sg13g2_o21ai_1 _23037_ (.B1(_04841_),
    .Y(_01931_),
    .A1(net317),
    .A2(_04840_));
 sg13g2_nand2_1 _23038_ (.Y(_04842_),
    .A(net613),
    .B(\mem.mem_internal.code_mem[74][2] ));
 sg13g2_nand2_1 _23039_ (.Y(_04843_),
    .A(net1012),
    .B(_04837_));
 sg13g2_o21ai_1 _23040_ (.B1(_04843_),
    .Y(_01932_),
    .A1(net317),
    .A2(_04842_));
 sg13g2_nand2_1 _23041_ (.Y(_04844_),
    .A(net613),
    .B(\mem.mem_internal.code_mem[74][3] ));
 sg13g2_nand2_1 _23042_ (.Y(_04845_),
    .A(net1011),
    .B(_04837_));
 sg13g2_o21ai_1 _23043_ (.B1(_04845_),
    .Y(_01933_),
    .A1(net317),
    .A2(_04844_));
 sg13g2_nand2_1 _23044_ (.Y(_04846_),
    .A(net613),
    .B(\mem.mem_internal.code_mem[74][4] ));
 sg13g2_nand2_1 _23045_ (.Y(_04847_),
    .A(net1010),
    .B(_04837_));
 sg13g2_o21ai_1 _23046_ (.B1(_04847_),
    .Y(_01934_),
    .A1(net317),
    .A2(_04846_));
 sg13g2_nand2_1 _23047_ (.Y(_04848_),
    .A(net613),
    .B(\mem.mem_internal.code_mem[74][5] ));
 sg13g2_nand2_1 _23048_ (.Y(_04849_),
    .A(net1009),
    .B(_04837_));
 sg13g2_o21ai_1 _23049_ (.B1(_04849_),
    .Y(_01935_),
    .A1(net317),
    .A2(_04848_));
 sg13g2_nand2_1 _23050_ (.Y(_04850_),
    .A(_04830_),
    .B(\mem.mem_internal.code_mem[74][6] ));
 sg13g2_nand2_1 _23051_ (.Y(_04851_),
    .A(net1008),
    .B(_04837_));
 sg13g2_o21ai_1 _23052_ (.B1(_04851_),
    .Y(_01936_),
    .A1(_04838_),
    .A2(_04850_));
 sg13g2_nand2_1 _23053_ (.Y(_04852_),
    .A(net613),
    .B(\mem.mem_internal.code_mem[74][7] ));
 sg13g2_nand2_1 _23054_ (.Y(_04853_),
    .A(net1007),
    .B(_04837_));
 sg13g2_o21ai_1 _23055_ (.B1(_04853_),
    .Y(_01937_),
    .A1(_04838_),
    .A2(_04852_));
 sg13g2_nand2_1 _23056_ (.Y(_04854_),
    .A(net835),
    .B(\mem.mem_internal.code_mem[75][0] ));
 sg13g2_nor2_1 _23057_ (.A(net775),
    .B(_04606_),
    .Y(_04855_));
 sg13g2_buf_2 _23058_ (.A(_04855_),
    .X(_04856_));
 sg13g2_buf_1 _23059_ (.A(_04856_),
    .X(_04857_));
 sg13g2_nand2_1 _23060_ (.Y(_04858_),
    .A(_04691_),
    .B(net316));
 sg13g2_o21ai_1 _23061_ (.B1(_04858_),
    .Y(_01938_),
    .A1(_04854_),
    .A2(net316));
 sg13g2_nand2_1 _23062_ (.Y(_04859_),
    .A(net613),
    .B(\mem.mem_internal.code_mem[75][1] ));
 sg13g2_nand2_1 _23063_ (.Y(_04860_),
    .A(_04694_),
    .B(net316));
 sg13g2_o21ai_1 _23064_ (.B1(_04860_),
    .Y(_01939_),
    .A1(net316),
    .A2(_04859_));
 sg13g2_buf_1 _23065_ (.A(_04829_),
    .X(_04861_));
 sg13g2_nand2_1 _23066_ (.Y(_04862_),
    .A(net612),
    .B(\mem.mem_internal.code_mem[75][2] ));
 sg13g2_nand2_1 _23067_ (.Y(_04863_),
    .A(_04697_),
    .B(_04856_));
 sg13g2_o21ai_1 _23068_ (.B1(_04863_),
    .Y(_01940_),
    .A1(net316),
    .A2(_04862_));
 sg13g2_nand2_1 _23069_ (.Y(_04864_),
    .A(net612),
    .B(\mem.mem_internal.code_mem[75][3] ));
 sg13g2_nand2_1 _23070_ (.Y(_04865_),
    .A(net1011),
    .B(_04856_));
 sg13g2_o21ai_1 _23071_ (.B1(_04865_),
    .Y(_01941_),
    .A1(net316),
    .A2(_04864_));
 sg13g2_nand2_1 _23072_ (.Y(_04866_),
    .A(net612),
    .B(\mem.mem_internal.code_mem[75][4] ));
 sg13g2_nand2_1 _23073_ (.Y(_04867_),
    .A(_04703_),
    .B(_04856_));
 sg13g2_o21ai_1 _23074_ (.B1(_04867_),
    .Y(_01942_),
    .A1(net316),
    .A2(_04866_));
 sg13g2_nand2_1 _23075_ (.Y(_04868_),
    .A(net612),
    .B(\mem.mem_internal.code_mem[75][5] ));
 sg13g2_nand2_1 _23076_ (.Y(_04869_),
    .A(_04706_),
    .B(_04856_));
 sg13g2_o21ai_1 _23077_ (.B1(_04869_),
    .Y(_01943_),
    .A1(_04857_),
    .A2(_04868_));
 sg13g2_nand2_1 _23078_ (.Y(_04870_),
    .A(_04861_),
    .B(\mem.mem_internal.code_mem[75][6] ));
 sg13g2_nand2_1 _23079_ (.Y(_04871_),
    .A(_04709_),
    .B(_04856_));
 sg13g2_o21ai_1 _23080_ (.B1(_04871_),
    .Y(_01944_),
    .A1(_04857_),
    .A2(_04870_));
 sg13g2_nand2_1 _23081_ (.Y(_04872_),
    .A(net612),
    .B(\mem.mem_internal.code_mem[75][7] ));
 sg13g2_nand2_1 _23082_ (.Y(_04873_),
    .A(_04712_),
    .B(_04856_));
 sg13g2_o21ai_1 _23083_ (.B1(_04873_),
    .Y(_01945_),
    .A1(net316),
    .A2(_04872_));
 sg13g2_nand2_1 _23084_ (.Y(_04874_),
    .A(net835),
    .B(\mem.mem_internal.code_mem[76][0] ));
 sg13g2_nor2_1 _23085_ (.A(_10491_),
    .B(_04606_),
    .Y(_04875_));
 sg13g2_buf_2 _23086_ (.A(_04875_),
    .X(_04876_));
 sg13g2_buf_1 _23087_ (.A(_04876_),
    .X(_04877_));
 sg13g2_nand2_1 _23088_ (.Y(_04878_),
    .A(net1014),
    .B(net315));
 sg13g2_o21ai_1 _23089_ (.B1(_04878_),
    .Y(_01946_),
    .A1(_04874_),
    .A2(net315));
 sg13g2_nand2_1 _23090_ (.Y(_04879_),
    .A(net612),
    .B(\mem.mem_internal.code_mem[76][1] ));
 sg13g2_nand2_1 _23091_ (.Y(_04880_),
    .A(_04694_),
    .B(net315));
 sg13g2_o21ai_1 _23092_ (.B1(_04880_),
    .Y(_01947_),
    .A1(net315),
    .A2(_04879_));
 sg13g2_nand2_1 _23093_ (.Y(_04881_),
    .A(net612),
    .B(\mem.mem_internal.code_mem[76][2] ));
 sg13g2_nand2_1 _23094_ (.Y(_04882_),
    .A(_04697_),
    .B(_04876_));
 sg13g2_o21ai_1 _23095_ (.B1(_04882_),
    .Y(_01948_),
    .A1(net315),
    .A2(_04881_));
 sg13g2_nand2_1 _23096_ (.Y(_04883_),
    .A(net612),
    .B(\mem.mem_internal.code_mem[76][3] ));
 sg13g2_nand2_1 _23097_ (.Y(_04884_),
    .A(_04700_),
    .B(_04876_));
 sg13g2_o21ai_1 _23098_ (.B1(_04884_),
    .Y(_01949_),
    .A1(net315),
    .A2(_04883_));
 sg13g2_nand2_1 _23099_ (.Y(_04885_),
    .A(_04861_),
    .B(\mem.mem_internal.code_mem[76][4] ));
 sg13g2_nand2_1 _23100_ (.Y(_04886_),
    .A(net1010),
    .B(_04876_));
 sg13g2_o21ai_1 _23101_ (.B1(_04886_),
    .Y(_01950_),
    .A1(net315),
    .A2(_04885_));
 sg13g2_buf_1 _23102_ (.A(_04829_),
    .X(_04887_));
 sg13g2_nand2_1 _23103_ (.Y(_04888_),
    .A(net611),
    .B(\mem.mem_internal.code_mem[76][5] ));
 sg13g2_nand2_1 _23104_ (.Y(_04889_),
    .A(net1009),
    .B(_04876_));
 sg13g2_o21ai_1 _23105_ (.B1(_04889_),
    .Y(_01951_),
    .A1(_04877_),
    .A2(_04888_));
 sg13g2_nand2_1 _23106_ (.Y(_04890_),
    .A(net611),
    .B(\mem.mem_internal.code_mem[76][6] ));
 sg13g2_nand2_1 _23107_ (.Y(_04891_),
    .A(_04709_),
    .B(_04876_));
 sg13g2_o21ai_1 _23108_ (.B1(_04891_),
    .Y(_01952_),
    .A1(_04877_),
    .A2(_04890_));
 sg13g2_nand2_1 _23109_ (.Y(_04892_),
    .A(net611),
    .B(\mem.mem_internal.code_mem[76][7] ));
 sg13g2_nand2_1 _23110_ (.Y(_04893_),
    .A(_04712_),
    .B(_04876_));
 sg13g2_o21ai_1 _23111_ (.B1(_04893_),
    .Y(_01953_),
    .A1(net315),
    .A2(_04892_));
 sg13g2_nand2_1 _23112_ (.Y(_04894_),
    .A(net835),
    .B(\mem.mem_internal.code_mem[77][0] ));
 sg13g2_nor2_1 _23113_ (.A(_10513_),
    .B(_04606_),
    .Y(_04895_));
 sg13g2_buf_2 _23114_ (.A(_04895_),
    .X(_04896_));
 sg13g2_buf_1 _23115_ (.A(_04896_),
    .X(_04897_));
 sg13g2_buf_1 _23116_ (.A(_03842_),
    .X(_04898_));
 sg13g2_nand2_1 _23117_ (.Y(_04899_),
    .A(net1006),
    .B(net314));
 sg13g2_o21ai_1 _23118_ (.B1(_04899_),
    .Y(_01954_),
    .A1(_04894_),
    .A2(net314));
 sg13g2_nand2_1 _23119_ (.Y(_04900_),
    .A(net611),
    .B(\mem.mem_internal.code_mem[77][1] ));
 sg13g2_buf_1 _23120_ (.A(_03846_),
    .X(_04901_));
 sg13g2_nand2_1 _23121_ (.Y(_04902_),
    .A(net1005),
    .B(net314));
 sg13g2_o21ai_1 _23122_ (.B1(_04902_),
    .Y(_01955_),
    .A1(net314),
    .A2(_04900_));
 sg13g2_nand2_1 _23123_ (.Y(_04903_),
    .A(net611),
    .B(\mem.mem_internal.code_mem[77][2] ));
 sg13g2_buf_1 _23124_ (.A(_03850_),
    .X(_04904_));
 sg13g2_nand2_1 _23125_ (.Y(_04905_),
    .A(net1004),
    .B(_04896_));
 sg13g2_o21ai_1 _23126_ (.B1(_04905_),
    .Y(_01956_),
    .A1(net314),
    .A2(_04903_));
 sg13g2_nand2_1 _23127_ (.Y(_04906_),
    .A(net611),
    .B(\mem.mem_internal.code_mem[77][3] ));
 sg13g2_buf_1 _23128_ (.A(_03854_),
    .X(_04907_));
 sg13g2_nand2_1 _23129_ (.Y(_04908_),
    .A(net1003),
    .B(_04896_));
 sg13g2_o21ai_1 _23130_ (.B1(_04908_),
    .Y(_01957_),
    .A1(net314),
    .A2(_04906_));
 sg13g2_nand2_1 _23131_ (.Y(_04909_),
    .A(net611),
    .B(\mem.mem_internal.code_mem[77][4] ));
 sg13g2_buf_1 _23132_ (.A(_03859_),
    .X(_04910_));
 sg13g2_nand2_1 _23133_ (.Y(_04911_),
    .A(net1002),
    .B(_04896_));
 sg13g2_o21ai_1 _23134_ (.B1(_04911_),
    .Y(_01958_),
    .A1(net314),
    .A2(_04909_));
 sg13g2_nand2_1 _23135_ (.Y(_04912_),
    .A(_04887_),
    .B(\mem.mem_internal.code_mem[77][5] ));
 sg13g2_buf_1 _23136_ (.A(_03863_),
    .X(_04913_));
 sg13g2_nand2_1 _23137_ (.Y(_04914_),
    .A(net1001),
    .B(_04896_));
 sg13g2_o21ai_1 _23138_ (.B1(_04914_),
    .Y(_01959_),
    .A1(_04897_),
    .A2(_04912_));
 sg13g2_nand2_1 _23139_ (.Y(_04915_),
    .A(_04887_),
    .B(\mem.mem_internal.code_mem[77][6] ));
 sg13g2_buf_1 _23140_ (.A(_03867_),
    .X(_04916_));
 sg13g2_nand2_1 _23141_ (.Y(_04917_),
    .A(net1000),
    .B(_04896_));
 sg13g2_o21ai_1 _23142_ (.B1(_04917_),
    .Y(_01960_),
    .A1(_04897_),
    .A2(_04915_));
 sg13g2_nand2_1 _23143_ (.Y(_04918_),
    .A(net611),
    .B(\mem.mem_internal.code_mem[77][7] ));
 sg13g2_buf_1 _23144_ (.A(_03871_),
    .X(_04919_));
 sg13g2_nand2_1 _23145_ (.Y(_04920_),
    .A(net999),
    .B(_04896_));
 sg13g2_o21ai_1 _23146_ (.B1(_04920_),
    .Y(_01961_),
    .A1(net314),
    .A2(_04918_));
 sg13g2_nand2_1 _23147_ (.Y(_04921_),
    .A(_04754_),
    .B(\mem.mem_internal.code_mem[78][0] ));
 sg13g2_nor2_1 _23148_ (.A(_10564_),
    .B(_04606_),
    .Y(_04922_));
 sg13g2_buf_2 _23149_ (.A(_04922_),
    .X(_04923_));
 sg13g2_buf_1 _23150_ (.A(_04923_),
    .X(_04924_));
 sg13g2_nand2_1 _23151_ (.Y(_04925_),
    .A(net1006),
    .B(net313));
 sg13g2_o21ai_1 _23152_ (.B1(_04925_),
    .Y(_01962_),
    .A1(_04921_),
    .A2(net313));
 sg13g2_buf_1 _23153_ (.A(_04829_),
    .X(_04926_));
 sg13g2_nand2_1 _23154_ (.Y(_04927_),
    .A(net610),
    .B(\mem.mem_internal.code_mem[78][1] ));
 sg13g2_nand2_1 _23155_ (.Y(_04928_),
    .A(net1005),
    .B(net313));
 sg13g2_o21ai_1 _23156_ (.B1(_04928_),
    .Y(_01963_),
    .A1(net313),
    .A2(_04927_));
 sg13g2_nand2_1 _23157_ (.Y(_04929_),
    .A(net610),
    .B(\mem.mem_internal.code_mem[78][2] ));
 sg13g2_nand2_1 _23158_ (.Y(_04930_),
    .A(net1004),
    .B(_04923_));
 sg13g2_o21ai_1 _23159_ (.B1(_04930_),
    .Y(_01964_),
    .A1(net313),
    .A2(_04929_));
 sg13g2_nand2_1 _23160_ (.Y(_04931_),
    .A(net610),
    .B(\mem.mem_internal.code_mem[78][3] ));
 sg13g2_nand2_1 _23161_ (.Y(_04932_),
    .A(net1003),
    .B(_04923_));
 sg13g2_o21ai_1 _23162_ (.B1(_04932_),
    .Y(_01965_),
    .A1(net313),
    .A2(_04931_));
 sg13g2_nand2_1 _23163_ (.Y(_04933_),
    .A(net610),
    .B(\mem.mem_internal.code_mem[78][4] ));
 sg13g2_nand2_1 _23164_ (.Y(_04934_),
    .A(_04910_),
    .B(_04923_));
 sg13g2_o21ai_1 _23165_ (.B1(_04934_),
    .Y(_01966_),
    .A1(net313),
    .A2(_04933_));
 sg13g2_nand2_1 _23166_ (.Y(_04935_),
    .A(_04926_),
    .B(\mem.mem_internal.code_mem[78][5] ));
 sg13g2_nand2_1 _23167_ (.Y(_04936_),
    .A(_04913_),
    .B(_04923_));
 sg13g2_o21ai_1 _23168_ (.B1(_04936_),
    .Y(_01967_),
    .A1(_04924_),
    .A2(_04935_));
 sg13g2_nand2_1 _23169_ (.Y(_04937_),
    .A(_04926_),
    .B(\mem.mem_internal.code_mem[78][6] ));
 sg13g2_nand2_1 _23170_ (.Y(_04938_),
    .A(_04916_),
    .B(_04923_));
 sg13g2_o21ai_1 _23171_ (.B1(_04938_),
    .Y(_01968_),
    .A1(_04924_),
    .A2(_04937_));
 sg13g2_nand2_1 _23172_ (.Y(_04939_),
    .A(net610),
    .B(\mem.mem_internal.code_mem[78][7] ));
 sg13g2_nand2_1 _23173_ (.Y(_04940_),
    .A(net999),
    .B(_04923_));
 sg13g2_o21ai_1 _23174_ (.B1(_04940_),
    .Y(_01969_),
    .A1(net313),
    .A2(_04939_));
 sg13g2_nand2_1 _23175_ (.Y(_04941_),
    .A(_04754_),
    .B(\mem.mem_internal.code_mem[79][0] ));
 sg13g2_nor2_1 _23176_ (.A(_10586_),
    .B(_04606_),
    .Y(_04942_));
 sg13g2_buf_2 _23177_ (.A(_04942_),
    .X(_04943_));
 sg13g2_buf_1 _23178_ (.A(_04943_),
    .X(_04944_));
 sg13g2_nand2_1 _23179_ (.Y(_04945_),
    .A(net1006),
    .B(net312));
 sg13g2_o21ai_1 _23180_ (.B1(_04945_),
    .Y(_01970_),
    .A1(_04941_),
    .A2(net312));
 sg13g2_nand2_1 _23181_ (.Y(_04946_),
    .A(net610),
    .B(\mem.mem_internal.code_mem[79][1] ));
 sg13g2_nand2_1 _23182_ (.Y(_04947_),
    .A(net1005),
    .B(net312));
 sg13g2_o21ai_1 _23183_ (.B1(_04947_),
    .Y(_01971_),
    .A1(net312),
    .A2(_04946_));
 sg13g2_nand2_1 _23184_ (.Y(_04948_),
    .A(net610),
    .B(\mem.mem_internal.code_mem[79][2] ));
 sg13g2_nand2_1 _23185_ (.Y(_04949_),
    .A(net1004),
    .B(_04943_));
 sg13g2_o21ai_1 _23186_ (.B1(_04949_),
    .Y(_01972_),
    .A1(net312),
    .A2(_04948_));
 sg13g2_nand2_1 _23187_ (.Y(_04950_),
    .A(net610),
    .B(\mem.mem_internal.code_mem[79][3] ));
 sg13g2_nand2_1 _23188_ (.Y(_04951_),
    .A(net1003),
    .B(_04943_));
 sg13g2_o21ai_1 _23189_ (.B1(_04951_),
    .Y(_01973_),
    .A1(net312),
    .A2(_04950_));
 sg13g2_buf_1 _23190_ (.A(_04829_),
    .X(_04952_));
 sg13g2_nand2_1 _23191_ (.Y(_04953_),
    .A(net609),
    .B(\mem.mem_internal.code_mem[79][4] ));
 sg13g2_nand2_1 _23192_ (.Y(_04954_),
    .A(_04910_),
    .B(_04943_));
 sg13g2_o21ai_1 _23193_ (.B1(_04954_),
    .Y(_01974_),
    .A1(net312),
    .A2(_04953_));
 sg13g2_nand2_1 _23194_ (.Y(_04955_),
    .A(net609),
    .B(\mem.mem_internal.code_mem[79][5] ));
 sg13g2_nand2_1 _23195_ (.Y(_04956_),
    .A(_04913_),
    .B(_04943_));
 sg13g2_o21ai_1 _23196_ (.B1(_04956_),
    .Y(_01975_),
    .A1(net312),
    .A2(_04955_));
 sg13g2_nand2_1 _23197_ (.Y(_04957_),
    .A(_04952_),
    .B(\mem.mem_internal.code_mem[79][6] ));
 sg13g2_nand2_1 _23198_ (.Y(_04958_),
    .A(_04916_),
    .B(_04943_));
 sg13g2_o21ai_1 _23199_ (.B1(_04958_),
    .Y(_01976_),
    .A1(_04944_),
    .A2(_04957_));
 sg13g2_nand2_1 _23200_ (.Y(_04959_),
    .A(_04952_),
    .B(\mem.mem_internal.code_mem[79][7] ));
 sg13g2_nand2_1 _23201_ (.Y(_04960_),
    .A(net999),
    .B(_04943_));
 sg13g2_o21ai_1 _23202_ (.B1(_04960_),
    .Y(_01977_),
    .A1(_04944_),
    .A2(_04959_));
 sg13g2_buf_1 _23203_ (.A(net1192),
    .X(_04961_));
 sg13g2_nand2_1 _23204_ (.Y(_04962_),
    .A(_04961_),
    .B(\mem.mem_internal.code_mem[7][0] ));
 sg13g2_nor2_1 _23205_ (.A(_10246_),
    .B(net553),
    .Y(_04963_));
 sg13g2_buf_1 _23206_ (.A(_04963_),
    .X(_04964_));
 sg13g2_buf_1 _23207_ (.A(_04964_),
    .X(_04965_));
 sg13g2_nand2_1 _23208_ (.Y(_04966_),
    .A(net1006),
    .B(_04965_));
 sg13g2_o21ai_1 _23209_ (.B1(_04966_),
    .Y(_01978_),
    .A1(_04962_),
    .A2(net311));
 sg13g2_nand2_1 _23210_ (.Y(_04967_),
    .A(net609),
    .B(\mem.mem_internal.code_mem[7][1] ));
 sg13g2_nand2_1 _23211_ (.Y(_04968_),
    .A(net1005),
    .B(_04965_));
 sg13g2_o21ai_1 _23212_ (.B1(_04968_),
    .Y(_01979_),
    .A1(net311),
    .A2(_04967_));
 sg13g2_nand2_1 _23213_ (.Y(_04969_),
    .A(net609),
    .B(\mem.mem_internal.code_mem[7][2] ));
 sg13g2_nand2_1 _23214_ (.Y(_04970_),
    .A(net1004),
    .B(_04964_));
 sg13g2_o21ai_1 _23215_ (.B1(_04970_),
    .Y(_01980_),
    .A1(net311),
    .A2(_04969_));
 sg13g2_nand2_1 _23216_ (.Y(_04971_),
    .A(net609),
    .B(\mem.mem_internal.code_mem[7][3] ));
 sg13g2_nand2_1 _23217_ (.Y(_04972_),
    .A(net1003),
    .B(_04964_));
 sg13g2_o21ai_1 _23218_ (.B1(_04972_),
    .Y(_01981_),
    .A1(net311),
    .A2(_04971_));
 sg13g2_nand2_1 _23219_ (.Y(_04973_),
    .A(net609),
    .B(\mem.mem_internal.code_mem[7][4] ));
 sg13g2_nand2_1 _23220_ (.Y(_04974_),
    .A(net1002),
    .B(_04964_));
 sg13g2_o21ai_1 _23221_ (.B1(_04974_),
    .Y(_01982_),
    .A1(net311),
    .A2(_04973_));
 sg13g2_nand2_1 _23222_ (.Y(_04975_),
    .A(net609),
    .B(\mem.mem_internal.code_mem[7][5] ));
 sg13g2_nand2_1 _23223_ (.Y(_04976_),
    .A(net1001),
    .B(_04964_));
 sg13g2_o21ai_1 _23224_ (.B1(_04976_),
    .Y(_01983_),
    .A1(net311),
    .A2(_04975_));
 sg13g2_nand2_1 _23225_ (.Y(_04977_),
    .A(net609),
    .B(\mem.mem_internal.code_mem[7][6] ));
 sg13g2_nand2_1 _23226_ (.Y(_04978_),
    .A(net1000),
    .B(_04964_));
 sg13g2_o21ai_1 _23227_ (.B1(_04978_),
    .Y(_01984_),
    .A1(net311),
    .A2(_04977_));
 sg13g2_buf_1 _23228_ (.A(_04829_),
    .X(_04979_));
 sg13g2_nand2_1 _23229_ (.Y(_04980_),
    .A(net608),
    .B(\mem.mem_internal.code_mem[7][7] ));
 sg13g2_nand2_1 _23230_ (.Y(_04981_),
    .A(net999),
    .B(_04964_));
 sg13g2_o21ai_1 _23231_ (.B1(_04981_),
    .Y(_01985_),
    .A1(net311),
    .A2(_04980_));
 sg13g2_nand2_1 _23232_ (.Y(_04982_),
    .A(net834),
    .B(\mem.mem_internal.code_mem[80][0] ));
 sg13g2_nand2_1 _23233_ (.Y(_04983_),
    .A(_10297_),
    .B(_11355_));
 sg13g2_buf_2 _23234_ (.A(_04983_),
    .X(_04984_));
 sg13g2_buf_1 _23235_ (.A(_04984_),
    .X(_04985_));
 sg13g2_nor2_1 _23236_ (.A(_10232_),
    .B(net456),
    .Y(_04986_));
 sg13g2_buf_2 _23237_ (.A(_04986_),
    .X(_04987_));
 sg13g2_buf_1 _23238_ (.A(_04987_),
    .X(_04988_));
 sg13g2_nand2_1 _23239_ (.Y(_04989_),
    .A(net1006),
    .B(net154));
 sg13g2_o21ai_1 _23240_ (.B1(_04989_),
    .Y(_01986_),
    .A1(_04982_),
    .A2(net154));
 sg13g2_nand2_1 _23241_ (.Y(_04990_),
    .A(net608),
    .B(\mem.mem_internal.code_mem[80][1] ));
 sg13g2_nand2_1 _23242_ (.Y(_04991_),
    .A(net1005),
    .B(_04988_));
 sg13g2_o21ai_1 _23243_ (.B1(_04991_),
    .Y(_01987_),
    .A1(_04988_),
    .A2(_04990_));
 sg13g2_nand2_1 _23244_ (.Y(_04992_),
    .A(net608),
    .B(\mem.mem_internal.code_mem[80][2] ));
 sg13g2_nand2_1 _23245_ (.Y(_04993_),
    .A(net1004),
    .B(_04987_));
 sg13g2_o21ai_1 _23246_ (.B1(_04993_),
    .Y(_01988_),
    .A1(net154),
    .A2(_04992_));
 sg13g2_nand2_1 _23247_ (.Y(_04994_),
    .A(net608),
    .B(\mem.mem_internal.code_mem[80][3] ));
 sg13g2_nand2_1 _23248_ (.Y(_04995_),
    .A(net1003),
    .B(_04987_));
 sg13g2_o21ai_1 _23249_ (.B1(_04995_),
    .Y(_01989_),
    .A1(net154),
    .A2(_04994_));
 sg13g2_nand2_1 _23250_ (.Y(_04996_),
    .A(net608),
    .B(\mem.mem_internal.code_mem[80][4] ));
 sg13g2_nand2_1 _23251_ (.Y(_04997_),
    .A(net1002),
    .B(_04987_));
 sg13g2_o21ai_1 _23252_ (.B1(_04997_),
    .Y(_01990_),
    .A1(net154),
    .A2(_04996_));
 sg13g2_nand2_1 _23253_ (.Y(_04998_),
    .A(net608),
    .B(\mem.mem_internal.code_mem[80][5] ));
 sg13g2_nand2_1 _23254_ (.Y(_04999_),
    .A(net1001),
    .B(_04987_));
 sg13g2_o21ai_1 _23255_ (.B1(_04999_),
    .Y(_01991_),
    .A1(net154),
    .A2(_04998_));
 sg13g2_nand2_1 _23256_ (.Y(_05000_),
    .A(net608),
    .B(\mem.mem_internal.code_mem[80][6] ));
 sg13g2_nand2_1 _23257_ (.Y(_05001_),
    .A(net1000),
    .B(_04987_));
 sg13g2_o21ai_1 _23258_ (.B1(_05001_),
    .Y(_01992_),
    .A1(net154),
    .A2(_05000_));
 sg13g2_nand2_1 _23259_ (.Y(_05002_),
    .A(_04979_),
    .B(\mem.mem_internal.code_mem[80][7] ));
 sg13g2_nand2_1 _23260_ (.Y(_05003_),
    .A(_04919_),
    .B(_04987_));
 sg13g2_o21ai_1 _23261_ (.B1(_05003_),
    .Y(_01993_),
    .A1(net154),
    .A2(_05002_));
 sg13g2_nand2_1 _23262_ (.Y(_05004_),
    .A(net834),
    .B(\mem.mem_internal.code_mem[81][0] ));
 sg13g2_nor2_1 _23263_ (.A(_10632_),
    .B(net456),
    .Y(_05005_));
 sg13g2_buf_2 _23264_ (.A(_05005_),
    .X(_05006_));
 sg13g2_buf_1 _23265_ (.A(_05006_),
    .X(_05007_));
 sg13g2_nand2_1 _23266_ (.Y(_05008_),
    .A(net1006),
    .B(net153));
 sg13g2_o21ai_1 _23267_ (.B1(_05008_),
    .Y(_01994_),
    .A1(_05004_),
    .A2(net153));
 sg13g2_nand2_1 _23268_ (.Y(_05009_),
    .A(net608),
    .B(\mem.mem_internal.code_mem[81][1] ));
 sg13g2_nand2_1 _23269_ (.Y(_05010_),
    .A(net1005),
    .B(net153));
 sg13g2_o21ai_1 _23270_ (.B1(_05010_),
    .Y(_01995_),
    .A1(_05007_),
    .A2(_05009_));
 sg13g2_nand2_1 _23271_ (.Y(_05011_),
    .A(_04979_),
    .B(\mem.mem_internal.code_mem[81][2] ));
 sg13g2_nand2_1 _23272_ (.Y(_05012_),
    .A(net1004),
    .B(_05006_));
 sg13g2_o21ai_1 _23273_ (.B1(_05012_),
    .Y(_01996_),
    .A1(net153),
    .A2(_05011_));
 sg13g2_buf_1 _23274_ (.A(_04829_),
    .X(_05013_));
 sg13g2_nand2_1 _23275_ (.Y(_05014_),
    .A(net607),
    .B(\mem.mem_internal.code_mem[81][3] ));
 sg13g2_nand2_1 _23276_ (.Y(_05015_),
    .A(net1003),
    .B(_05006_));
 sg13g2_o21ai_1 _23277_ (.B1(_05015_),
    .Y(_01997_),
    .A1(net153),
    .A2(_05014_));
 sg13g2_nand2_1 _23278_ (.Y(_05016_),
    .A(net607),
    .B(\mem.mem_internal.code_mem[81][4] ));
 sg13g2_nand2_1 _23279_ (.Y(_05017_),
    .A(net1002),
    .B(_05006_));
 sg13g2_o21ai_1 _23280_ (.B1(_05017_),
    .Y(_01998_),
    .A1(net153),
    .A2(_05016_));
 sg13g2_nand2_1 _23281_ (.Y(_05018_),
    .A(net607),
    .B(\mem.mem_internal.code_mem[81][5] ));
 sg13g2_nand2_1 _23282_ (.Y(_05019_),
    .A(net1001),
    .B(_05006_));
 sg13g2_o21ai_1 _23283_ (.B1(_05019_),
    .Y(_01999_),
    .A1(net153),
    .A2(_05018_));
 sg13g2_nand2_1 _23284_ (.Y(_05020_),
    .A(net607),
    .B(\mem.mem_internal.code_mem[81][6] ));
 sg13g2_nand2_1 _23285_ (.Y(_05021_),
    .A(net1000),
    .B(_05006_));
 sg13g2_o21ai_1 _23286_ (.B1(_05021_),
    .Y(_02000_),
    .A1(net153),
    .A2(_05020_));
 sg13g2_nand2_1 _23287_ (.Y(_05022_),
    .A(_05013_),
    .B(\mem.mem_internal.code_mem[81][7] ));
 sg13g2_nand2_1 _23288_ (.Y(_05023_),
    .A(net999),
    .B(_05006_));
 sg13g2_o21ai_1 _23289_ (.B1(_05023_),
    .Y(_02001_),
    .A1(_05007_),
    .A2(_05022_));
 sg13g2_nand2_1 _23290_ (.Y(_05024_),
    .A(net834),
    .B(\mem.mem_internal.code_mem[82][0] ));
 sg13g2_nor2_1 _23291_ (.A(_10656_),
    .B(net456),
    .Y(_05025_));
 sg13g2_buf_2 _23292_ (.A(_05025_),
    .X(_05026_));
 sg13g2_buf_1 _23293_ (.A(_05026_),
    .X(_05027_));
 sg13g2_nand2_1 _23294_ (.Y(_05028_),
    .A(net1006),
    .B(net152));
 sg13g2_o21ai_1 _23295_ (.B1(_05028_),
    .Y(_02002_),
    .A1(_05024_),
    .A2(net152));
 sg13g2_nand2_1 _23296_ (.Y(_05029_),
    .A(_05013_),
    .B(\mem.mem_internal.code_mem[82][1] ));
 sg13g2_nand2_1 _23297_ (.Y(_05030_),
    .A(net1005),
    .B(_05027_));
 sg13g2_o21ai_1 _23298_ (.B1(_05030_),
    .Y(_02003_),
    .A1(_05027_),
    .A2(_05029_));
 sg13g2_nand2_1 _23299_ (.Y(_05031_),
    .A(net607),
    .B(\mem.mem_internal.code_mem[82][2] ));
 sg13g2_nand2_1 _23300_ (.Y(_05032_),
    .A(net1004),
    .B(_05026_));
 sg13g2_o21ai_1 _23301_ (.B1(_05032_),
    .Y(_02004_),
    .A1(net152),
    .A2(_05031_));
 sg13g2_nand2_1 _23302_ (.Y(_05033_),
    .A(net607),
    .B(\mem.mem_internal.code_mem[82][3] ));
 sg13g2_nand2_1 _23303_ (.Y(_05034_),
    .A(net1003),
    .B(_05026_));
 sg13g2_o21ai_1 _23304_ (.B1(_05034_),
    .Y(_02005_),
    .A1(net152),
    .A2(_05033_));
 sg13g2_nand2_1 _23305_ (.Y(_05035_),
    .A(net607),
    .B(\mem.mem_internal.code_mem[82][4] ));
 sg13g2_nand2_1 _23306_ (.Y(_05036_),
    .A(net1002),
    .B(_05026_));
 sg13g2_o21ai_1 _23307_ (.B1(_05036_),
    .Y(_02006_),
    .A1(net152),
    .A2(_05035_));
 sg13g2_nand2_1 _23308_ (.Y(_05037_),
    .A(net607),
    .B(\mem.mem_internal.code_mem[82][5] ));
 sg13g2_nand2_1 _23309_ (.Y(_05038_),
    .A(net1001),
    .B(_05026_));
 sg13g2_o21ai_1 _23310_ (.B1(_05038_),
    .Y(_02007_),
    .A1(net152),
    .A2(_05037_));
 sg13g2_buf_1 _23311_ (.A(_04431_),
    .X(_05039_));
 sg13g2_buf_1 _23312_ (.A(_05039_),
    .X(_05040_));
 sg13g2_nand2_1 _23313_ (.Y(_05041_),
    .A(net606),
    .B(\mem.mem_internal.code_mem[82][6] ));
 sg13g2_nand2_1 _23314_ (.Y(_05042_),
    .A(net1000),
    .B(_05026_));
 sg13g2_o21ai_1 _23315_ (.B1(_05042_),
    .Y(_02008_),
    .A1(net152),
    .A2(_05041_));
 sg13g2_nand2_1 _23316_ (.Y(_05043_),
    .A(net606),
    .B(\mem.mem_internal.code_mem[82][7] ));
 sg13g2_nand2_1 _23317_ (.Y(_05044_),
    .A(net999),
    .B(_05026_));
 sg13g2_o21ai_1 _23318_ (.B1(_05044_),
    .Y(_02009_),
    .A1(net152),
    .A2(_05043_));
 sg13g2_nand2_1 _23319_ (.Y(_05045_),
    .A(net834),
    .B(\mem.mem_internal.code_mem[83][0] ));
 sg13g2_nor2_1 _23320_ (.A(_10679_),
    .B(net456),
    .Y(_05046_));
 sg13g2_buf_2 _23321_ (.A(_05046_),
    .X(_05047_));
 sg13g2_buf_1 _23322_ (.A(_05047_),
    .X(_05048_));
 sg13g2_nand2_1 _23323_ (.Y(_05049_),
    .A(net1006),
    .B(net151));
 sg13g2_o21ai_1 _23324_ (.B1(_05049_),
    .Y(_02010_),
    .A1(_05045_),
    .A2(net151));
 sg13g2_nand2_1 _23325_ (.Y(_05050_),
    .A(net606),
    .B(\mem.mem_internal.code_mem[83][1] ));
 sg13g2_nand2_1 _23326_ (.Y(_05051_),
    .A(net1005),
    .B(_05048_));
 sg13g2_o21ai_1 _23327_ (.B1(_05051_),
    .Y(_02011_),
    .A1(_05048_),
    .A2(_05050_));
 sg13g2_nand2_1 _23328_ (.Y(_05052_),
    .A(_05040_),
    .B(\mem.mem_internal.code_mem[83][2] ));
 sg13g2_nand2_1 _23329_ (.Y(_05053_),
    .A(net1004),
    .B(_05047_));
 sg13g2_o21ai_1 _23330_ (.B1(_05053_),
    .Y(_02012_),
    .A1(net151),
    .A2(_05052_));
 sg13g2_nand2_1 _23331_ (.Y(_05054_),
    .A(net606),
    .B(\mem.mem_internal.code_mem[83][3] ));
 sg13g2_nand2_1 _23332_ (.Y(_05055_),
    .A(net1003),
    .B(_05047_));
 sg13g2_o21ai_1 _23333_ (.B1(_05055_),
    .Y(_02013_),
    .A1(net151),
    .A2(_05054_));
 sg13g2_nand2_1 _23334_ (.Y(_05056_),
    .A(net606),
    .B(\mem.mem_internal.code_mem[83][4] ));
 sg13g2_nand2_1 _23335_ (.Y(_05057_),
    .A(net1002),
    .B(_05047_));
 sg13g2_o21ai_1 _23336_ (.B1(_05057_),
    .Y(_02014_),
    .A1(net151),
    .A2(_05056_));
 sg13g2_nand2_1 _23337_ (.Y(_05058_),
    .A(net606),
    .B(\mem.mem_internal.code_mem[83][5] ));
 sg13g2_nand2_1 _23338_ (.Y(_05059_),
    .A(net1001),
    .B(_05047_));
 sg13g2_o21ai_1 _23339_ (.B1(_05059_),
    .Y(_02015_),
    .A1(net151),
    .A2(_05058_));
 sg13g2_nand2_1 _23340_ (.Y(_05060_),
    .A(net606),
    .B(\mem.mem_internal.code_mem[83][6] ));
 sg13g2_nand2_1 _23341_ (.Y(_05061_),
    .A(net1000),
    .B(_05047_));
 sg13g2_o21ai_1 _23342_ (.B1(_05061_),
    .Y(_02016_),
    .A1(net151),
    .A2(_05060_));
 sg13g2_nand2_1 _23343_ (.Y(_05062_),
    .A(net606),
    .B(\mem.mem_internal.code_mem[83][7] ));
 sg13g2_nand2_1 _23344_ (.Y(_05063_),
    .A(_04919_),
    .B(_05047_));
 sg13g2_o21ai_1 _23345_ (.B1(_05063_),
    .Y(_02017_),
    .A1(net151),
    .A2(_05062_));
 sg13g2_nand2_1 _23346_ (.Y(_05064_),
    .A(net834),
    .B(\mem.mem_internal.code_mem[84][0] ));
 sg13g2_nor2_1 _23347_ (.A(_10295_),
    .B(net456),
    .Y(_05065_));
 sg13g2_buf_2 _23348_ (.A(_05065_),
    .X(_05066_));
 sg13g2_buf_1 _23349_ (.A(_05066_),
    .X(_05067_));
 sg13g2_nand2_1 _23350_ (.Y(_05068_),
    .A(_04898_),
    .B(net150));
 sg13g2_o21ai_1 _23351_ (.B1(_05068_),
    .Y(_02018_),
    .A1(_05064_),
    .A2(net150));
 sg13g2_nand2_1 _23352_ (.Y(_05069_),
    .A(_05040_),
    .B(\mem.mem_internal.code_mem[84][1] ));
 sg13g2_nand2_1 _23353_ (.Y(_05070_),
    .A(_04901_),
    .B(net150));
 sg13g2_o21ai_1 _23354_ (.B1(_05070_),
    .Y(_02019_),
    .A1(net150),
    .A2(_05069_));
 sg13g2_buf_1 _23355_ (.A(_05039_),
    .X(_05071_));
 sg13g2_nand2_1 _23356_ (.Y(_05072_),
    .A(net605),
    .B(\mem.mem_internal.code_mem[84][2] ));
 sg13g2_nand2_1 _23357_ (.Y(_05073_),
    .A(_04904_),
    .B(_05066_));
 sg13g2_o21ai_1 _23358_ (.B1(_05073_),
    .Y(_02020_),
    .A1(net150),
    .A2(_05072_));
 sg13g2_nand2_1 _23359_ (.Y(_05074_),
    .A(net605),
    .B(\mem.mem_internal.code_mem[84][3] ));
 sg13g2_nand2_1 _23360_ (.Y(_05075_),
    .A(_04907_),
    .B(_05066_));
 sg13g2_o21ai_1 _23361_ (.B1(_05075_),
    .Y(_02021_),
    .A1(net150),
    .A2(_05074_));
 sg13g2_nand2_1 _23362_ (.Y(_05076_),
    .A(net605),
    .B(\mem.mem_internal.code_mem[84][4] ));
 sg13g2_nand2_1 _23363_ (.Y(_05077_),
    .A(net1002),
    .B(_05066_));
 sg13g2_o21ai_1 _23364_ (.B1(_05077_),
    .Y(_02022_),
    .A1(net150),
    .A2(_05076_));
 sg13g2_nand2_1 _23365_ (.Y(_05078_),
    .A(net605),
    .B(\mem.mem_internal.code_mem[84][5] ));
 sg13g2_nand2_1 _23366_ (.Y(_05079_),
    .A(net1001),
    .B(_05066_));
 sg13g2_o21ai_1 _23367_ (.B1(_05079_),
    .Y(_02023_),
    .A1(_05067_),
    .A2(_05078_));
 sg13g2_nand2_1 _23368_ (.Y(_05080_),
    .A(net605),
    .B(\mem.mem_internal.code_mem[84][6] ));
 sg13g2_nand2_1 _23369_ (.Y(_05081_),
    .A(net1000),
    .B(_05066_));
 sg13g2_o21ai_1 _23370_ (.B1(_05081_),
    .Y(_02024_),
    .A1(_05067_),
    .A2(_05080_));
 sg13g2_nand2_1 _23371_ (.Y(_05082_),
    .A(net605),
    .B(\mem.mem_internal.code_mem[84][7] ));
 sg13g2_nand2_1 _23372_ (.Y(_05083_),
    .A(net999),
    .B(_05066_));
 sg13g2_o21ai_1 _23373_ (.B1(_05083_),
    .Y(_02025_),
    .A1(net150),
    .A2(_05082_));
 sg13g2_nand2_1 _23374_ (.Y(_05084_),
    .A(net834),
    .B(\mem.mem_internal.code_mem[85][0] ));
 sg13g2_nor2_1 _23375_ (.A(_10325_),
    .B(net456),
    .Y(_05085_));
 sg13g2_buf_2 _23376_ (.A(_05085_),
    .X(_05086_));
 sg13g2_buf_1 _23377_ (.A(_05086_),
    .X(_05087_));
 sg13g2_nand2_1 _23378_ (.Y(_05088_),
    .A(_04898_),
    .B(net149));
 sg13g2_o21ai_1 _23379_ (.B1(_05088_),
    .Y(_02026_),
    .A1(_05084_),
    .A2(net149));
 sg13g2_nand2_1 _23380_ (.Y(_05089_),
    .A(net605),
    .B(\mem.mem_internal.code_mem[85][1] ));
 sg13g2_nand2_1 _23381_ (.Y(_05090_),
    .A(_04901_),
    .B(net149));
 sg13g2_o21ai_1 _23382_ (.B1(_05090_),
    .Y(_02027_),
    .A1(net149),
    .A2(_05089_));
 sg13g2_nand2_1 _23383_ (.Y(_05091_),
    .A(net605),
    .B(\mem.mem_internal.code_mem[85][2] ));
 sg13g2_nand2_1 _23384_ (.Y(_05092_),
    .A(_04904_),
    .B(_05086_));
 sg13g2_o21ai_1 _23385_ (.B1(_05092_),
    .Y(_02028_),
    .A1(net149),
    .A2(_05091_));
 sg13g2_nand2_1 _23386_ (.Y(_05093_),
    .A(_05071_),
    .B(\mem.mem_internal.code_mem[85][3] ));
 sg13g2_nand2_1 _23387_ (.Y(_05094_),
    .A(_04907_),
    .B(_05086_));
 sg13g2_o21ai_1 _23388_ (.B1(_05094_),
    .Y(_02029_),
    .A1(net149),
    .A2(_05093_));
 sg13g2_nand2_1 _23389_ (.Y(_05095_),
    .A(_05071_),
    .B(\mem.mem_internal.code_mem[85][4] ));
 sg13g2_nand2_1 _23390_ (.Y(_05096_),
    .A(net1002),
    .B(_05086_));
 sg13g2_o21ai_1 _23391_ (.B1(_05096_),
    .Y(_02030_),
    .A1(net149),
    .A2(_05095_));
 sg13g2_buf_1 _23392_ (.A(_05039_),
    .X(_05097_));
 sg13g2_nand2_1 _23393_ (.Y(_05098_),
    .A(_05097_),
    .B(\mem.mem_internal.code_mem[85][5] ));
 sg13g2_nand2_1 _23394_ (.Y(_05099_),
    .A(net1001),
    .B(_05086_));
 sg13g2_o21ai_1 _23395_ (.B1(_05099_),
    .Y(_02031_),
    .A1(_05087_),
    .A2(_05098_));
 sg13g2_nand2_1 _23396_ (.Y(_05100_),
    .A(_05097_),
    .B(\mem.mem_internal.code_mem[85][6] ));
 sg13g2_nand2_1 _23397_ (.Y(_05101_),
    .A(net1000),
    .B(_05086_));
 sg13g2_o21ai_1 _23398_ (.B1(_05101_),
    .Y(_02032_),
    .A1(_05087_),
    .A2(_05100_));
 sg13g2_nand2_1 _23399_ (.Y(_05102_),
    .A(net604),
    .B(\mem.mem_internal.code_mem[85][7] ));
 sg13g2_nand2_1 _23400_ (.Y(_05103_),
    .A(net999),
    .B(_05086_));
 sg13g2_o21ai_1 _23401_ (.B1(_05103_),
    .Y(_02033_),
    .A1(net149),
    .A2(_05102_));
 sg13g2_nand2_1 _23402_ (.Y(_05104_),
    .A(net834),
    .B(\mem.mem_internal.code_mem[86][0] ));
 sg13g2_nor2_1 _23403_ (.A(net779),
    .B(net456),
    .Y(_05105_));
 sg13g2_buf_2 _23404_ (.A(_05105_),
    .X(_05106_));
 sg13g2_buf_1 _23405_ (.A(_05106_),
    .X(_05107_));
 sg13g2_buf_1 _23406_ (.A(_03842_),
    .X(_05108_));
 sg13g2_nand2_1 _23407_ (.Y(_05109_),
    .A(net998),
    .B(net148));
 sg13g2_o21ai_1 _23408_ (.B1(_05109_),
    .Y(_02034_),
    .A1(_05104_),
    .A2(net148));
 sg13g2_nand2_1 _23409_ (.Y(_05110_),
    .A(net604),
    .B(\mem.mem_internal.code_mem[86][1] ));
 sg13g2_buf_1 _23410_ (.A(_03846_),
    .X(_05111_));
 sg13g2_nand2_1 _23411_ (.Y(_05112_),
    .A(net997),
    .B(net148));
 sg13g2_o21ai_1 _23412_ (.B1(_05112_),
    .Y(_02035_),
    .A1(net148),
    .A2(_05110_));
 sg13g2_nand2_1 _23413_ (.Y(_05113_),
    .A(net604),
    .B(\mem.mem_internal.code_mem[86][2] ));
 sg13g2_buf_1 _23414_ (.A(_03850_),
    .X(_05114_));
 sg13g2_nand2_1 _23415_ (.Y(_05115_),
    .A(net996),
    .B(_05106_));
 sg13g2_o21ai_1 _23416_ (.B1(_05115_),
    .Y(_02036_),
    .A1(net148),
    .A2(_05113_));
 sg13g2_nand2_1 _23417_ (.Y(_05116_),
    .A(net604),
    .B(\mem.mem_internal.code_mem[86][3] ));
 sg13g2_buf_1 _23418_ (.A(_03854_),
    .X(_05117_));
 sg13g2_nand2_1 _23419_ (.Y(_05118_),
    .A(net995),
    .B(_05106_));
 sg13g2_o21ai_1 _23420_ (.B1(_05118_),
    .Y(_02037_),
    .A1(net148),
    .A2(_05116_));
 sg13g2_nand2_1 _23421_ (.Y(_05119_),
    .A(net604),
    .B(\mem.mem_internal.code_mem[86][4] ));
 sg13g2_buf_1 _23422_ (.A(_03859_),
    .X(_05120_));
 sg13g2_nand2_1 _23423_ (.Y(_05121_),
    .A(net994),
    .B(_05106_));
 sg13g2_o21ai_1 _23424_ (.B1(_05121_),
    .Y(_02038_),
    .A1(net148),
    .A2(_05119_));
 sg13g2_nand2_1 _23425_ (.Y(_05122_),
    .A(net604),
    .B(\mem.mem_internal.code_mem[86][5] ));
 sg13g2_buf_1 _23426_ (.A(_03863_),
    .X(_05123_));
 sg13g2_nand2_1 _23427_ (.Y(_05124_),
    .A(net993),
    .B(_05106_));
 sg13g2_o21ai_1 _23428_ (.B1(_05124_),
    .Y(_02039_),
    .A1(net148),
    .A2(_05122_));
 sg13g2_nand2_1 _23429_ (.Y(_05125_),
    .A(net604),
    .B(\mem.mem_internal.code_mem[86][6] ));
 sg13g2_buf_1 _23430_ (.A(_03867_),
    .X(_05126_));
 sg13g2_nand2_1 _23431_ (.Y(_05127_),
    .A(net992),
    .B(_05106_));
 sg13g2_o21ai_1 _23432_ (.B1(_05127_),
    .Y(_02040_),
    .A1(_05107_),
    .A2(_05125_));
 sg13g2_nand2_1 _23433_ (.Y(_05128_),
    .A(net604),
    .B(\mem.mem_internal.code_mem[86][7] ));
 sg13g2_buf_1 _23434_ (.A(_03871_),
    .X(_05129_));
 sg13g2_nand2_1 _23435_ (.Y(_05130_),
    .A(net991),
    .B(_05106_));
 sg13g2_o21ai_1 _23436_ (.B1(_05130_),
    .Y(_02041_),
    .A1(_05107_),
    .A2(_05128_));
 sg13g2_nand2_1 _23437_ (.Y(_05131_),
    .A(_04961_),
    .B(\mem.mem_internal.code_mem[87][0] ));
 sg13g2_nor2_1 _23438_ (.A(_10372_),
    .B(net456),
    .Y(_05132_));
 sg13g2_buf_2 _23439_ (.A(_05132_),
    .X(_05133_));
 sg13g2_buf_1 _23440_ (.A(_05133_),
    .X(_05134_));
 sg13g2_nand2_1 _23441_ (.Y(_05135_),
    .A(net998),
    .B(net147));
 sg13g2_o21ai_1 _23442_ (.B1(_05135_),
    .Y(_02042_),
    .A1(_05131_),
    .A2(net147));
 sg13g2_buf_1 _23443_ (.A(_05039_),
    .X(_05136_));
 sg13g2_nand2_1 _23444_ (.Y(_05137_),
    .A(net603),
    .B(\mem.mem_internal.code_mem[87][1] ));
 sg13g2_nand2_1 _23445_ (.Y(_05138_),
    .A(net997),
    .B(net147));
 sg13g2_o21ai_1 _23446_ (.B1(_05138_),
    .Y(_02043_),
    .A1(net147),
    .A2(_05137_));
 sg13g2_nand2_1 _23447_ (.Y(_05139_),
    .A(_05136_),
    .B(\mem.mem_internal.code_mem[87][2] ));
 sg13g2_nand2_1 _23448_ (.Y(_05140_),
    .A(net996),
    .B(_05133_));
 sg13g2_o21ai_1 _23449_ (.B1(_05140_),
    .Y(_02044_),
    .A1(_05134_),
    .A2(_05139_));
 sg13g2_nand2_1 _23450_ (.Y(_05141_),
    .A(net603),
    .B(\mem.mem_internal.code_mem[87][3] ));
 sg13g2_nand2_1 _23451_ (.Y(_05142_),
    .A(net995),
    .B(_05133_));
 sg13g2_o21ai_1 _23452_ (.B1(_05142_),
    .Y(_02045_),
    .A1(net147),
    .A2(_05141_));
 sg13g2_nand2_1 _23453_ (.Y(_05143_),
    .A(net603),
    .B(\mem.mem_internal.code_mem[87][4] ));
 sg13g2_nand2_1 _23454_ (.Y(_05144_),
    .A(net994),
    .B(_05133_));
 sg13g2_o21ai_1 _23455_ (.B1(_05144_),
    .Y(_02046_),
    .A1(net147),
    .A2(_05143_));
 sg13g2_nand2_1 _23456_ (.Y(_05145_),
    .A(net603),
    .B(\mem.mem_internal.code_mem[87][5] ));
 sg13g2_nand2_1 _23457_ (.Y(_05146_),
    .A(net993),
    .B(_05133_));
 sg13g2_o21ai_1 _23458_ (.B1(_05146_),
    .Y(_02047_),
    .A1(net147),
    .A2(_05145_));
 sg13g2_nand2_1 _23459_ (.Y(_05147_),
    .A(_05136_),
    .B(\mem.mem_internal.code_mem[87][6] ));
 sg13g2_nand2_1 _23460_ (.Y(_05148_),
    .A(net992),
    .B(_05133_));
 sg13g2_o21ai_1 _23461_ (.B1(_05148_),
    .Y(_02048_),
    .A1(_05134_),
    .A2(_05147_));
 sg13g2_nand2_1 _23462_ (.Y(_05149_),
    .A(net603),
    .B(\mem.mem_internal.code_mem[87][7] ));
 sg13g2_nand2_1 _23463_ (.Y(_05150_),
    .A(net991),
    .B(_05133_));
 sg13g2_o21ai_1 _23464_ (.B1(_05150_),
    .Y(_02049_),
    .A1(net147),
    .A2(_05149_));
 sg13g2_nand2_1 _23465_ (.Y(_05151_),
    .A(net834),
    .B(\mem.mem_internal.code_mem[88][0] ));
 sg13g2_nor2_1 _23466_ (.A(_10397_),
    .B(_04985_),
    .Y(_05152_));
 sg13g2_buf_2 _23467_ (.A(_05152_),
    .X(_05153_));
 sg13g2_buf_1 _23468_ (.A(_05153_),
    .X(_05154_));
 sg13g2_nand2_1 _23469_ (.Y(_05155_),
    .A(net998),
    .B(net146));
 sg13g2_o21ai_1 _23470_ (.B1(_05155_),
    .Y(_02050_),
    .A1(_05151_),
    .A2(net146));
 sg13g2_nand2_1 _23471_ (.Y(_05156_),
    .A(net603),
    .B(\mem.mem_internal.code_mem[88][1] ));
 sg13g2_nand2_1 _23472_ (.Y(_05157_),
    .A(net997),
    .B(net146));
 sg13g2_o21ai_1 _23473_ (.B1(_05157_),
    .Y(_02051_),
    .A1(net146),
    .A2(_05156_));
 sg13g2_nand2_1 _23474_ (.Y(_05158_),
    .A(net603),
    .B(\mem.mem_internal.code_mem[88][2] ));
 sg13g2_nand2_1 _23475_ (.Y(_05159_),
    .A(net996),
    .B(_05153_));
 sg13g2_o21ai_1 _23476_ (.B1(_05159_),
    .Y(_02052_),
    .A1(net146),
    .A2(_05158_));
 sg13g2_nand2_1 _23477_ (.Y(_05160_),
    .A(net603),
    .B(\mem.mem_internal.code_mem[88][3] ));
 sg13g2_nand2_1 _23478_ (.Y(_05161_),
    .A(net995),
    .B(_05153_));
 sg13g2_o21ai_1 _23479_ (.B1(_05161_),
    .Y(_02053_),
    .A1(net146),
    .A2(_05160_));
 sg13g2_buf_1 _23480_ (.A(_05039_),
    .X(_05162_));
 sg13g2_nand2_1 _23481_ (.Y(_05163_),
    .A(net602),
    .B(\mem.mem_internal.code_mem[88][4] ));
 sg13g2_nand2_1 _23482_ (.Y(_05164_),
    .A(net994),
    .B(_05153_));
 sg13g2_o21ai_1 _23483_ (.B1(_05164_),
    .Y(_02054_),
    .A1(net146),
    .A2(_05163_));
 sg13g2_nand2_1 _23484_ (.Y(_05165_),
    .A(net602),
    .B(\mem.mem_internal.code_mem[88][5] ));
 sg13g2_nand2_1 _23485_ (.Y(_05166_),
    .A(net993),
    .B(_05153_));
 sg13g2_o21ai_1 _23486_ (.B1(_05166_),
    .Y(_02055_),
    .A1(_05154_),
    .A2(_05165_));
 sg13g2_nand2_1 _23487_ (.Y(_05167_),
    .A(net602),
    .B(\mem.mem_internal.code_mem[88][6] ));
 sg13g2_nand2_1 _23488_ (.Y(_05168_),
    .A(net992),
    .B(_05153_));
 sg13g2_o21ai_1 _23489_ (.B1(_05168_),
    .Y(_02056_),
    .A1(_05154_),
    .A2(_05167_));
 sg13g2_nand2_1 _23490_ (.Y(_05169_),
    .A(net602),
    .B(\mem.mem_internal.code_mem[88][7] ));
 sg13g2_nand2_1 _23491_ (.Y(_05170_),
    .A(net991),
    .B(_05153_));
 sg13g2_o21ai_1 _23492_ (.B1(_05170_),
    .Y(_02057_),
    .A1(net146),
    .A2(_05169_));
 sg13g2_buf_1 _23493_ (.A(net1192),
    .X(_05171_));
 sg13g2_nand2_1 _23494_ (.Y(_05172_),
    .A(net833),
    .B(\mem.mem_internal.code_mem[89][0] ));
 sg13g2_nor2_1 _23495_ (.A(_10422_),
    .B(_04985_),
    .Y(_05173_));
 sg13g2_buf_2 _23496_ (.A(_05173_),
    .X(_05174_));
 sg13g2_buf_1 _23497_ (.A(_05174_),
    .X(_05175_));
 sg13g2_nand2_1 _23498_ (.Y(_05176_),
    .A(_05108_),
    .B(net145));
 sg13g2_o21ai_1 _23499_ (.B1(_05176_),
    .Y(_02058_),
    .A1(_05172_),
    .A2(net145));
 sg13g2_nand2_1 _23500_ (.Y(_05177_),
    .A(net602),
    .B(\mem.mem_internal.code_mem[89][1] ));
 sg13g2_nand2_1 _23501_ (.Y(_05178_),
    .A(net997),
    .B(net145));
 sg13g2_o21ai_1 _23502_ (.B1(_05178_),
    .Y(_02059_),
    .A1(net145),
    .A2(_05177_));
 sg13g2_nand2_1 _23503_ (.Y(_05179_),
    .A(net602),
    .B(\mem.mem_internal.code_mem[89][2] ));
 sg13g2_nand2_1 _23504_ (.Y(_05180_),
    .A(net996),
    .B(_05174_));
 sg13g2_o21ai_1 _23505_ (.B1(_05180_),
    .Y(_02060_),
    .A1(net145),
    .A2(_05179_));
 sg13g2_nand2_1 _23506_ (.Y(_05181_),
    .A(net602),
    .B(\mem.mem_internal.code_mem[89][3] ));
 sg13g2_nand2_1 _23507_ (.Y(_05182_),
    .A(net995),
    .B(_05174_));
 sg13g2_o21ai_1 _23508_ (.B1(_05182_),
    .Y(_02061_),
    .A1(net145),
    .A2(_05181_));
 sg13g2_nand2_1 _23509_ (.Y(_05183_),
    .A(net602),
    .B(\mem.mem_internal.code_mem[89][4] ));
 sg13g2_nand2_1 _23510_ (.Y(_05184_),
    .A(net994),
    .B(_05174_));
 sg13g2_o21ai_1 _23511_ (.B1(_05184_),
    .Y(_02062_),
    .A1(net145),
    .A2(_05183_));
 sg13g2_nand2_1 _23512_ (.Y(_05185_),
    .A(_05162_),
    .B(\mem.mem_internal.code_mem[89][5] ));
 sg13g2_nand2_1 _23513_ (.Y(_05186_),
    .A(net993),
    .B(_05174_));
 sg13g2_o21ai_1 _23514_ (.B1(_05186_),
    .Y(_02063_),
    .A1(_05175_),
    .A2(_05185_));
 sg13g2_nand2_1 _23515_ (.Y(_05187_),
    .A(_05162_),
    .B(\mem.mem_internal.code_mem[89][6] ));
 sg13g2_nand2_1 _23516_ (.Y(_05188_),
    .A(net992),
    .B(_05174_));
 sg13g2_o21ai_1 _23517_ (.B1(_05188_),
    .Y(_02064_),
    .A1(_05175_),
    .A2(_05187_));
 sg13g2_buf_1 _23518_ (.A(_05039_),
    .X(_05189_));
 sg13g2_nand2_1 _23519_ (.Y(_05190_),
    .A(_05189_),
    .B(\mem.mem_internal.code_mem[89][7] ));
 sg13g2_nand2_1 _23520_ (.Y(_05191_),
    .A(net991),
    .B(_05174_));
 sg13g2_o21ai_1 _23521_ (.B1(_05191_),
    .Y(_02065_),
    .A1(net145),
    .A2(_05190_));
 sg13g2_nand2_1 _23522_ (.Y(_05192_),
    .A(net833),
    .B(\mem.mem_internal.code_mem[8][0] ));
 sg13g2_nor2_1 _23523_ (.A(_10246_),
    .B(_10398_),
    .Y(_05193_));
 sg13g2_buf_1 _23524_ (.A(_05193_),
    .X(_05194_));
 sg13g2_buf_1 _23525_ (.A(_05194_),
    .X(_05195_));
 sg13g2_nand2_1 _23526_ (.Y(_05196_),
    .A(net998),
    .B(net310));
 sg13g2_o21ai_1 _23527_ (.B1(_05196_),
    .Y(_02066_),
    .A1(_05192_),
    .A2(_05195_));
 sg13g2_nand2_1 _23528_ (.Y(_05197_),
    .A(net601),
    .B(\mem.mem_internal.code_mem[8][1] ));
 sg13g2_nand2_1 _23529_ (.Y(_05198_),
    .A(net997),
    .B(_05195_));
 sg13g2_o21ai_1 _23530_ (.B1(_05198_),
    .Y(_02067_),
    .A1(net310),
    .A2(_05197_));
 sg13g2_nand2_1 _23531_ (.Y(_05199_),
    .A(net601),
    .B(\mem.mem_internal.code_mem[8][2] ));
 sg13g2_nand2_1 _23532_ (.Y(_05200_),
    .A(net996),
    .B(_05194_));
 sg13g2_o21ai_1 _23533_ (.B1(_05200_),
    .Y(_02068_),
    .A1(net310),
    .A2(_05199_));
 sg13g2_nand2_1 _23534_ (.Y(_05201_),
    .A(net601),
    .B(\mem.mem_internal.code_mem[8][3] ));
 sg13g2_nand2_1 _23535_ (.Y(_05202_),
    .A(net995),
    .B(_05194_));
 sg13g2_o21ai_1 _23536_ (.B1(_05202_),
    .Y(_02069_),
    .A1(net310),
    .A2(_05201_));
 sg13g2_nand2_1 _23537_ (.Y(_05203_),
    .A(net601),
    .B(\mem.mem_internal.code_mem[8][4] ));
 sg13g2_nand2_1 _23538_ (.Y(_05204_),
    .A(net994),
    .B(_05194_));
 sg13g2_o21ai_1 _23539_ (.B1(_05204_),
    .Y(_02070_),
    .A1(net310),
    .A2(_05203_));
 sg13g2_nand2_1 _23540_ (.Y(_05205_),
    .A(net601),
    .B(\mem.mem_internal.code_mem[8][5] ));
 sg13g2_nand2_1 _23541_ (.Y(_05206_),
    .A(net993),
    .B(_05194_));
 sg13g2_o21ai_1 _23542_ (.B1(_05206_),
    .Y(_02071_),
    .A1(net310),
    .A2(_05205_));
 sg13g2_nand2_1 _23543_ (.Y(_05207_),
    .A(net601),
    .B(\mem.mem_internal.code_mem[8][6] ));
 sg13g2_nand2_1 _23544_ (.Y(_05208_),
    .A(net992),
    .B(_05194_));
 sg13g2_o21ai_1 _23545_ (.B1(_05208_),
    .Y(_02072_),
    .A1(net310),
    .A2(_05207_));
 sg13g2_nand2_1 _23546_ (.Y(_05209_),
    .A(net601),
    .B(\mem.mem_internal.code_mem[8][7] ));
 sg13g2_nand2_1 _23547_ (.Y(_05210_),
    .A(net991),
    .B(_05194_));
 sg13g2_o21ai_1 _23548_ (.B1(_05210_),
    .Y(_02073_),
    .A1(net310),
    .A2(_05209_));
 sg13g2_nand2_1 _23549_ (.Y(_05211_),
    .A(net833),
    .B(\mem.mem_internal.code_mem[90][0] ));
 sg13g2_nor2_1 _23550_ (.A(_10444_),
    .B(_04984_),
    .Y(_05212_));
 sg13g2_buf_2 _23551_ (.A(_05212_),
    .X(_05213_));
 sg13g2_buf_1 _23552_ (.A(_05213_),
    .X(_05214_));
 sg13g2_nand2_1 _23553_ (.Y(_05215_),
    .A(_05108_),
    .B(net309));
 sg13g2_o21ai_1 _23554_ (.B1(_05215_),
    .Y(_02074_),
    .A1(_05211_),
    .A2(net309));
 sg13g2_nand2_1 _23555_ (.Y(_05216_),
    .A(net601),
    .B(\mem.mem_internal.code_mem[90][1] ));
 sg13g2_nand2_1 _23556_ (.Y(_05217_),
    .A(_05111_),
    .B(net309));
 sg13g2_o21ai_1 _23557_ (.B1(_05217_),
    .Y(_02075_),
    .A1(net309),
    .A2(_05216_));
 sg13g2_nand2_1 _23558_ (.Y(_05218_),
    .A(_05189_),
    .B(\mem.mem_internal.code_mem[90][2] ));
 sg13g2_nand2_1 _23559_ (.Y(_05219_),
    .A(_05114_),
    .B(_05213_));
 sg13g2_o21ai_1 _23560_ (.B1(_05219_),
    .Y(_02076_),
    .A1(net309),
    .A2(_05218_));
 sg13g2_buf_1 _23561_ (.A(_05039_),
    .X(_05220_));
 sg13g2_nand2_1 _23562_ (.Y(_05221_),
    .A(net600),
    .B(\mem.mem_internal.code_mem[90][3] ));
 sg13g2_nand2_1 _23563_ (.Y(_05222_),
    .A(_05117_),
    .B(_05213_));
 sg13g2_o21ai_1 _23564_ (.B1(_05222_),
    .Y(_02077_),
    .A1(net309),
    .A2(_05221_));
 sg13g2_nand2_1 _23565_ (.Y(_05223_),
    .A(net600),
    .B(\mem.mem_internal.code_mem[90][4] ));
 sg13g2_nand2_1 _23566_ (.Y(_05224_),
    .A(_05120_),
    .B(_05213_));
 sg13g2_o21ai_1 _23567_ (.B1(_05224_),
    .Y(_02078_),
    .A1(net309),
    .A2(_05223_));
 sg13g2_nand2_1 _23568_ (.Y(_05225_),
    .A(net600),
    .B(\mem.mem_internal.code_mem[90][5] ));
 sg13g2_nand2_1 _23569_ (.Y(_05226_),
    .A(_05123_),
    .B(_05213_));
 sg13g2_o21ai_1 _23570_ (.B1(_05226_),
    .Y(_02079_),
    .A1(_05214_),
    .A2(_05225_));
 sg13g2_nand2_1 _23571_ (.Y(_05227_),
    .A(net600),
    .B(\mem.mem_internal.code_mem[90][6] ));
 sg13g2_nand2_1 _23572_ (.Y(_05228_),
    .A(_05126_),
    .B(_05213_));
 sg13g2_o21ai_1 _23573_ (.B1(_05228_),
    .Y(_02080_),
    .A1(_05214_),
    .A2(_05227_));
 sg13g2_nand2_1 _23574_ (.Y(_05229_),
    .A(net600),
    .B(\mem.mem_internal.code_mem[90][7] ));
 sg13g2_nand2_1 _23575_ (.Y(_05230_),
    .A(_05129_),
    .B(_05213_));
 sg13g2_o21ai_1 _23576_ (.B1(_05230_),
    .Y(_02081_),
    .A1(net309),
    .A2(_05229_));
 sg13g2_nand2_1 _23577_ (.Y(_05231_),
    .A(net833),
    .B(\mem.mem_internal.code_mem[91][0] ));
 sg13g2_nor2_1 _23578_ (.A(_10467_),
    .B(_04984_),
    .Y(_05232_));
 sg13g2_buf_2 _23579_ (.A(_05232_),
    .X(_05233_));
 sg13g2_buf_1 _23580_ (.A(_05233_),
    .X(_05234_));
 sg13g2_nand2_1 _23581_ (.Y(_05235_),
    .A(net998),
    .B(net308));
 sg13g2_o21ai_1 _23582_ (.B1(_05235_),
    .Y(_02082_),
    .A1(_05231_),
    .A2(net308));
 sg13g2_nand2_1 _23583_ (.Y(_05236_),
    .A(net600),
    .B(\mem.mem_internal.code_mem[91][1] ));
 sg13g2_nand2_1 _23584_ (.Y(_05237_),
    .A(_05111_),
    .B(net308));
 sg13g2_o21ai_1 _23585_ (.B1(_05237_),
    .Y(_02083_),
    .A1(net308),
    .A2(_05236_));
 sg13g2_nand2_1 _23586_ (.Y(_05238_),
    .A(net600),
    .B(\mem.mem_internal.code_mem[91][2] ));
 sg13g2_nand2_1 _23587_ (.Y(_05239_),
    .A(_05114_),
    .B(_05233_));
 sg13g2_o21ai_1 _23588_ (.B1(_05239_),
    .Y(_02084_),
    .A1(net308),
    .A2(_05238_));
 sg13g2_nand2_1 _23589_ (.Y(_05240_),
    .A(net600),
    .B(\mem.mem_internal.code_mem[91][3] ));
 sg13g2_nand2_1 _23590_ (.Y(_05241_),
    .A(_05117_),
    .B(_05233_));
 sg13g2_o21ai_1 _23591_ (.B1(_05241_),
    .Y(_02085_),
    .A1(net308),
    .A2(_05240_));
 sg13g2_nand2_1 _23592_ (.Y(_05242_),
    .A(_05220_),
    .B(\mem.mem_internal.code_mem[91][4] ));
 sg13g2_nand2_1 _23593_ (.Y(_05243_),
    .A(_05120_),
    .B(_05233_));
 sg13g2_o21ai_1 _23594_ (.B1(_05243_),
    .Y(_02086_),
    .A1(net308),
    .A2(_05242_));
 sg13g2_nand2_1 _23595_ (.Y(_05244_),
    .A(_05220_),
    .B(\mem.mem_internal.code_mem[91][5] ));
 sg13g2_nand2_1 _23596_ (.Y(_05245_),
    .A(_05123_),
    .B(_05233_));
 sg13g2_o21ai_1 _23597_ (.B1(_05245_),
    .Y(_02087_),
    .A1(_05234_),
    .A2(_05244_));
 sg13g2_buf_1 _23598_ (.A(_04431_),
    .X(_05246_));
 sg13g2_buf_1 _23599_ (.A(_05246_),
    .X(_05247_));
 sg13g2_nand2_1 _23600_ (.Y(_05248_),
    .A(net599),
    .B(\mem.mem_internal.code_mem[91][6] ));
 sg13g2_nand2_1 _23601_ (.Y(_05249_),
    .A(_05126_),
    .B(_05233_));
 sg13g2_o21ai_1 _23602_ (.B1(_05249_),
    .Y(_02088_),
    .A1(_05234_),
    .A2(_05248_));
 sg13g2_nand2_1 _23603_ (.Y(_05250_),
    .A(net599),
    .B(\mem.mem_internal.code_mem[91][7] ));
 sg13g2_nand2_1 _23604_ (.Y(_05251_),
    .A(_05129_),
    .B(_05233_));
 sg13g2_o21ai_1 _23605_ (.B1(_05251_),
    .Y(_02089_),
    .A1(net308),
    .A2(_05250_));
 sg13g2_nand2_1 _23606_ (.Y(_05252_),
    .A(net833),
    .B(\mem.mem_internal.code_mem[92][0] ));
 sg13g2_nor2_1 _23607_ (.A(_10491_),
    .B(_04984_),
    .Y(_05253_));
 sg13g2_buf_2 _23608_ (.A(_05253_),
    .X(_05254_));
 sg13g2_buf_1 _23609_ (.A(_05254_),
    .X(_05255_));
 sg13g2_nand2_1 _23610_ (.Y(_05256_),
    .A(net998),
    .B(net307));
 sg13g2_o21ai_1 _23611_ (.B1(_05256_),
    .Y(_02090_),
    .A1(_05252_),
    .A2(net307));
 sg13g2_nand2_1 _23612_ (.Y(_05257_),
    .A(net599),
    .B(\mem.mem_internal.code_mem[92][1] ));
 sg13g2_nand2_1 _23613_ (.Y(_05258_),
    .A(net997),
    .B(net307));
 sg13g2_o21ai_1 _23614_ (.B1(_05258_),
    .Y(_02091_),
    .A1(net307),
    .A2(_05257_));
 sg13g2_nand2_1 _23615_ (.Y(_05259_),
    .A(net599),
    .B(\mem.mem_internal.code_mem[92][2] ));
 sg13g2_nand2_1 _23616_ (.Y(_05260_),
    .A(net996),
    .B(_05254_));
 sg13g2_o21ai_1 _23617_ (.B1(_05260_),
    .Y(_02092_),
    .A1(net307),
    .A2(_05259_));
 sg13g2_nand2_1 _23618_ (.Y(_05261_),
    .A(net599),
    .B(\mem.mem_internal.code_mem[92][3] ));
 sg13g2_nand2_1 _23619_ (.Y(_05262_),
    .A(net995),
    .B(_05254_));
 sg13g2_o21ai_1 _23620_ (.B1(_05262_),
    .Y(_02093_),
    .A1(net307),
    .A2(_05261_));
 sg13g2_nand2_1 _23621_ (.Y(_05263_),
    .A(net599),
    .B(\mem.mem_internal.code_mem[92][4] ));
 sg13g2_nand2_1 _23622_ (.Y(_05264_),
    .A(net994),
    .B(_05254_));
 sg13g2_o21ai_1 _23623_ (.B1(_05264_),
    .Y(_02094_),
    .A1(net307),
    .A2(_05263_));
 sg13g2_nand2_1 _23624_ (.Y(_05265_),
    .A(_05247_),
    .B(\mem.mem_internal.code_mem[92][5] ));
 sg13g2_nand2_1 _23625_ (.Y(_05266_),
    .A(net993),
    .B(_05254_));
 sg13g2_o21ai_1 _23626_ (.B1(_05266_),
    .Y(_02095_),
    .A1(_05255_),
    .A2(_05265_));
 sg13g2_nand2_1 _23627_ (.Y(_05267_),
    .A(_05247_),
    .B(\mem.mem_internal.code_mem[92][6] ));
 sg13g2_nand2_1 _23628_ (.Y(_05268_),
    .A(net992),
    .B(_05254_));
 sg13g2_o21ai_1 _23629_ (.B1(_05268_),
    .Y(_02096_),
    .A1(_05255_),
    .A2(_05267_));
 sg13g2_nand2_1 _23630_ (.Y(_05269_),
    .A(net599),
    .B(\mem.mem_internal.code_mem[92][7] ));
 sg13g2_nand2_1 _23631_ (.Y(_05270_),
    .A(net991),
    .B(_05254_));
 sg13g2_o21ai_1 _23632_ (.B1(_05270_),
    .Y(_02097_),
    .A1(net307),
    .A2(_05269_));
 sg13g2_nand2_1 _23633_ (.Y(_05271_),
    .A(_05171_),
    .B(\mem.mem_internal.code_mem[93][0] ));
 sg13g2_nor2_1 _23634_ (.A(_10513_),
    .B(_04984_),
    .Y(_05272_));
 sg13g2_buf_2 _23635_ (.A(_05272_),
    .X(_05273_));
 sg13g2_buf_1 _23636_ (.A(_05273_),
    .X(_05274_));
 sg13g2_nand2_1 _23637_ (.Y(_05275_),
    .A(net998),
    .B(net306));
 sg13g2_o21ai_1 _23638_ (.B1(_05275_),
    .Y(_02098_),
    .A1(_05271_),
    .A2(net306));
 sg13g2_nand2_1 _23639_ (.Y(_05276_),
    .A(net599),
    .B(\mem.mem_internal.code_mem[93][1] ));
 sg13g2_nand2_1 _23640_ (.Y(_05277_),
    .A(net997),
    .B(net306));
 sg13g2_o21ai_1 _23641_ (.B1(_05277_),
    .Y(_02099_),
    .A1(net306),
    .A2(_05276_));
 sg13g2_buf_1 _23642_ (.A(_05246_),
    .X(_05278_));
 sg13g2_nand2_1 _23643_ (.Y(_05279_),
    .A(net598),
    .B(\mem.mem_internal.code_mem[93][2] ));
 sg13g2_nand2_1 _23644_ (.Y(_05280_),
    .A(net996),
    .B(_05273_));
 sg13g2_o21ai_1 _23645_ (.B1(_05280_),
    .Y(_02100_),
    .A1(net306),
    .A2(_05279_));
 sg13g2_nand2_1 _23646_ (.Y(_05281_),
    .A(net598),
    .B(\mem.mem_internal.code_mem[93][3] ));
 sg13g2_nand2_1 _23647_ (.Y(_05282_),
    .A(net995),
    .B(_05273_));
 sg13g2_o21ai_1 _23648_ (.B1(_05282_),
    .Y(_02101_),
    .A1(net306),
    .A2(_05281_));
 sg13g2_nand2_1 _23649_ (.Y(_05283_),
    .A(net598),
    .B(\mem.mem_internal.code_mem[93][4] ));
 sg13g2_nand2_1 _23650_ (.Y(_05284_),
    .A(net994),
    .B(_05273_));
 sg13g2_o21ai_1 _23651_ (.B1(_05284_),
    .Y(_02102_),
    .A1(net306),
    .A2(_05283_));
 sg13g2_nand2_1 _23652_ (.Y(_05285_),
    .A(_05278_),
    .B(\mem.mem_internal.code_mem[93][5] ));
 sg13g2_nand2_1 _23653_ (.Y(_05286_),
    .A(net993),
    .B(_05273_));
 sg13g2_o21ai_1 _23654_ (.B1(_05286_),
    .Y(_02103_),
    .A1(_05274_),
    .A2(_05285_));
 sg13g2_nand2_1 _23655_ (.Y(_05287_),
    .A(net598),
    .B(\mem.mem_internal.code_mem[93][6] ));
 sg13g2_nand2_1 _23656_ (.Y(_05288_),
    .A(net992),
    .B(_05273_));
 sg13g2_o21ai_1 _23657_ (.B1(_05288_),
    .Y(_02104_),
    .A1(_05274_),
    .A2(_05287_));
 sg13g2_nand2_1 _23658_ (.Y(_05289_),
    .A(net598),
    .B(\mem.mem_internal.code_mem[93][7] ));
 sg13g2_nand2_1 _23659_ (.Y(_05290_),
    .A(net991),
    .B(_05273_));
 sg13g2_o21ai_1 _23660_ (.B1(_05290_),
    .Y(_02105_),
    .A1(net306),
    .A2(_05289_));
 sg13g2_nand2_1 _23661_ (.Y(_05291_),
    .A(_05171_),
    .B(\mem.mem_internal.code_mem[94][0] ));
 sg13g2_nor2_1 _23662_ (.A(_10564_),
    .B(_04984_),
    .Y(_05292_));
 sg13g2_buf_2 _23663_ (.A(_05292_),
    .X(_05293_));
 sg13g2_buf_1 _23664_ (.A(_05293_),
    .X(_05294_));
 sg13g2_nand2_1 _23665_ (.Y(_05295_),
    .A(net998),
    .B(net305));
 sg13g2_o21ai_1 _23666_ (.B1(_05295_),
    .Y(_02106_),
    .A1(_05291_),
    .A2(net305));
 sg13g2_nand2_1 _23667_ (.Y(_05296_),
    .A(net598),
    .B(\mem.mem_internal.code_mem[94][1] ));
 sg13g2_nand2_1 _23668_ (.Y(_05297_),
    .A(net997),
    .B(net305));
 sg13g2_o21ai_1 _23669_ (.B1(_05297_),
    .Y(_02107_),
    .A1(net305),
    .A2(_05296_));
 sg13g2_nand2_1 _23670_ (.Y(_05298_),
    .A(net598),
    .B(\mem.mem_internal.code_mem[94][2] ));
 sg13g2_nand2_1 _23671_ (.Y(_05299_),
    .A(net996),
    .B(_05293_));
 sg13g2_o21ai_1 _23672_ (.B1(_05299_),
    .Y(_02108_),
    .A1(net305),
    .A2(_05298_));
 sg13g2_nand2_1 _23673_ (.Y(_05300_),
    .A(net598),
    .B(\mem.mem_internal.code_mem[94][3] ));
 sg13g2_nand2_1 _23674_ (.Y(_05301_),
    .A(net995),
    .B(_05293_));
 sg13g2_o21ai_1 _23675_ (.B1(_05301_),
    .Y(_02109_),
    .A1(net305),
    .A2(_05300_));
 sg13g2_nand2_1 _23676_ (.Y(_05302_),
    .A(_05278_),
    .B(\mem.mem_internal.code_mem[94][4] ));
 sg13g2_nand2_1 _23677_ (.Y(_05303_),
    .A(net994),
    .B(_05293_));
 sg13g2_o21ai_1 _23678_ (.B1(_05303_),
    .Y(_02110_),
    .A1(net305),
    .A2(_05302_));
 sg13g2_buf_1 _23679_ (.A(_05246_),
    .X(_05304_));
 sg13g2_nand2_1 _23680_ (.Y(_05305_),
    .A(_05304_),
    .B(\mem.mem_internal.code_mem[94][5] ));
 sg13g2_nand2_1 _23681_ (.Y(_05306_),
    .A(net993),
    .B(_05293_));
 sg13g2_o21ai_1 _23682_ (.B1(_05306_),
    .Y(_02111_),
    .A1(_05294_),
    .A2(_05305_));
 sg13g2_nand2_1 _23683_ (.Y(_05307_),
    .A(_05304_),
    .B(\mem.mem_internal.code_mem[94][6] ));
 sg13g2_nand2_1 _23684_ (.Y(_05308_),
    .A(net992),
    .B(_05293_));
 sg13g2_o21ai_1 _23685_ (.B1(_05308_),
    .Y(_02112_),
    .A1(_05294_),
    .A2(_05307_));
 sg13g2_nand2_1 _23686_ (.Y(_05309_),
    .A(net597),
    .B(\mem.mem_internal.code_mem[94][7] ));
 sg13g2_nand2_1 _23687_ (.Y(_05310_),
    .A(net991),
    .B(_05293_));
 sg13g2_o21ai_1 _23688_ (.B1(_05310_),
    .Y(_02113_),
    .A1(net305),
    .A2(_05309_));
 sg13g2_nand2_1 _23689_ (.Y(_05311_),
    .A(net833),
    .B(\mem.mem_internal.code_mem[95][0] ));
 sg13g2_nor2_1 _23690_ (.A(_10586_),
    .B(_04984_),
    .Y(_05312_));
 sg13g2_buf_1 _23691_ (.A(_05312_),
    .X(_05313_));
 sg13g2_buf_1 _23692_ (.A(_05313_),
    .X(_05314_));
 sg13g2_nand2_1 _23693_ (.Y(_05315_),
    .A(_10252_),
    .B(net304));
 sg13g2_o21ai_1 _23694_ (.B1(_05315_),
    .Y(_02114_),
    .A1(_05311_),
    .A2(net304));
 sg13g2_nand2_1 _23695_ (.Y(_05316_),
    .A(net597),
    .B(\mem.mem_internal.code_mem[95][1] ));
 sg13g2_nand2_1 _23696_ (.Y(_05317_),
    .A(net1267),
    .B(net304));
 sg13g2_o21ai_1 _23697_ (.B1(_05317_),
    .Y(_02115_),
    .A1(net304),
    .A2(_05316_));
 sg13g2_nand2_1 _23698_ (.Y(_05318_),
    .A(net597),
    .B(\mem.mem_internal.code_mem[95][2] ));
 sg13g2_nand2_1 _23699_ (.Y(_05319_),
    .A(_10263_),
    .B(_05313_));
 sg13g2_o21ai_1 _23700_ (.B1(_05319_),
    .Y(_02116_),
    .A1(net304),
    .A2(_05318_));
 sg13g2_nand2_1 _23701_ (.Y(_05320_),
    .A(net597),
    .B(\mem.mem_internal.code_mem[95][3] ));
 sg13g2_nand2_1 _23702_ (.Y(_05321_),
    .A(_10268_),
    .B(_05313_));
 sg13g2_o21ai_1 _23703_ (.B1(_05321_),
    .Y(_02117_),
    .A1(net304),
    .A2(_05320_));
 sg13g2_nand2_1 _23704_ (.Y(_05322_),
    .A(net597),
    .B(\mem.mem_internal.code_mem[95][4] ));
 sg13g2_nand2_1 _23705_ (.Y(_05323_),
    .A(_10273_),
    .B(_05313_));
 sg13g2_o21ai_1 _23706_ (.B1(_05323_),
    .Y(_02118_),
    .A1(net304),
    .A2(_05322_));
 sg13g2_nand2_1 _23707_ (.Y(_05324_),
    .A(net597),
    .B(\mem.mem_internal.code_mem[95][5] ));
 sg13g2_nand2_1 _23708_ (.Y(_05325_),
    .A(_10278_),
    .B(_05313_));
 sg13g2_o21ai_1 _23709_ (.B1(_05325_),
    .Y(_02119_),
    .A1(_05314_),
    .A2(_05324_));
 sg13g2_nand2_1 _23710_ (.Y(_05326_),
    .A(net597),
    .B(\mem.mem_internal.code_mem[95][6] ));
 sg13g2_nand2_1 _23711_ (.Y(_05327_),
    .A(_10283_),
    .B(_05313_));
 sg13g2_o21ai_1 _23712_ (.B1(_05327_),
    .Y(_02120_),
    .A1(_05314_),
    .A2(_05326_));
 sg13g2_nand2_1 _23713_ (.Y(_05328_),
    .A(net597),
    .B(\mem.mem_internal.code_mem[95][7] ));
 sg13g2_nand2_1 _23714_ (.Y(_05329_),
    .A(_10288_),
    .B(_05313_));
 sg13g2_o21ai_1 _23715_ (.B1(_05329_),
    .Y(_02121_),
    .A1(net304),
    .A2(_05328_));
 sg13g2_nand2_1 _23716_ (.Y(_05330_),
    .A(net833),
    .B(\mem.mem_internal.code_mem[96][0] ));
 sg13g2_nor2_1 _23717_ (.A(_10232_),
    .B(_10301_),
    .Y(_05331_));
 sg13g2_buf_2 _23718_ (.A(_05331_),
    .X(_05332_));
 sg13g2_buf_1 _23719_ (.A(_05332_),
    .X(_05333_));
 sg13g2_nand2_1 _23720_ (.Y(_05334_),
    .A(net1268),
    .B(_05333_));
 sg13g2_o21ai_1 _23721_ (.B1(_05334_),
    .Y(_02122_),
    .A1(_05330_),
    .A2(_05333_));
 sg13g2_buf_1 _23722_ (.A(_05246_),
    .X(_05335_));
 sg13g2_nand2_1 _23723_ (.Y(_05336_),
    .A(net596),
    .B(\mem.mem_internal.code_mem[96][1] ));
 sg13g2_nand2_1 _23724_ (.Y(_05337_),
    .A(net1267),
    .B(net144));
 sg13g2_o21ai_1 _23725_ (.B1(_05337_),
    .Y(_02123_),
    .A1(net144),
    .A2(_05336_));
 sg13g2_nand2_1 _23726_ (.Y(_05338_),
    .A(_05335_),
    .B(\mem.mem_internal.code_mem[96][2] ));
 sg13g2_nand2_1 _23727_ (.Y(_05339_),
    .A(net1266),
    .B(_05332_));
 sg13g2_o21ai_1 _23728_ (.B1(_05339_),
    .Y(_02124_),
    .A1(net144),
    .A2(_05338_));
 sg13g2_nand2_1 _23729_ (.Y(_05340_),
    .A(net596),
    .B(\mem.mem_internal.code_mem[96][3] ));
 sg13g2_nand2_1 _23730_ (.Y(_05341_),
    .A(net1265),
    .B(_05332_));
 sg13g2_o21ai_1 _23731_ (.B1(_05341_),
    .Y(_02125_),
    .A1(net144),
    .A2(_05340_));
 sg13g2_nand2_1 _23732_ (.Y(_05342_),
    .A(net596),
    .B(\mem.mem_internal.code_mem[96][4] ));
 sg13g2_nand2_1 _23733_ (.Y(_05343_),
    .A(net1264),
    .B(_05332_));
 sg13g2_o21ai_1 _23734_ (.B1(_05343_),
    .Y(_02126_),
    .A1(net144),
    .A2(_05342_));
 sg13g2_nand2_1 _23735_ (.Y(_05344_),
    .A(net596),
    .B(\mem.mem_internal.code_mem[96][5] ));
 sg13g2_nand2_1 _23736_ (.Y(_05345_),
    .A(net1263),
    .B(_05332_));
 sg13g2_o21ai_1 _23737_ (.B1(_05345_),
    .Y(_02127_),
    .A1(net144),
    .A2(_05344_));
 sg13g2_nand2_1 _23738_ (.Y(_05346_),
    .A(net596),
    .B(\mem.mem_internal.code_mem[96][6] ));
 sg13g2_nand2_1 _23739_ (.Y(_05347_),
    .A(net1262),
    .B(_05332_));
 sg13g2_o21ai_1 _23740_ (.B1(_05347_),
    .Y(_02128_),
    .A1(net144),
    .A2(_05346_));
 sg13g2_nand2_1 _23741_ (.Y(_05348_),
    .A(net596),
    .B(\mem.mem_internal.code_mem[96][7] ));
 sg13g2_nand2_1 _23742_ (.Y(_05349_),
    .A(net1261),
    .B(_05332_));
 sg13g2_o21ai_1 _23743_ (.B1(_05349_),
    .Y(_02129_),
    .A1(net144),
    .A2(_05348_));
 sg13g2_nand2_1 _23744_ (.Y(_05350_),
    .A(net833),
    .B(\mem.mem_internal.code_mem[97][0] ));
 sg13g2_nor2_1 _23745_ (.A(_10300_),
    .B(net528),
    .Y(_05351_));
 sg13g2_buf_2 _23746_ (.A(_05351_),
    .X(_05352_));
 sg13g2_buf_1 _23747_ (.A(_05352_),
    .X(_05353_));
 sg13g2_nand2_1 _23748_ (.Y(_05354_),
    .A(net1268),
    .B(_05353_));
 sg13g2_o21ai_1 _23749_ (.B1(_05354_),
    .Y(_02130_),
    .A1(_05350_),
    .A2(net303));
 sg13g2_nand2_1 _23750_ (.Y(_05355_),
    .A(net596),
    .B(\mem.mem_internal.code_mem[97][1] ));
 sg13g2_nand2_1 _23751_ (.Y(_05356_),
    .A(net1267),
    .B(net303));
 sg13g2_o21ai_1 _23752_ (.B1(_05356_),
    .Y(_02131_),
    .A1(net303),
    .A2(_05355_));
 sg13g2_nand2_1 _23753_ (.Y(_05357_),
    .A(_05335_),
    .B(\mem.mem_internal.code_mem[97][2] ));
 sg13g2_nand2_1 _23754_ (.Y(_05358_),
    .A(net1266),
    .B(_05352_));
 sg13g2_o21ai_1 _23755_ (.B1(_05358_),
    .Y(_02132_),
    .A1(net303),
    .A2(_05357_));
 sg13g2_nand2_1 _23756_ (.Y(_05359_),
    .A(net596),
    .B(\mem.mem_internal.code_mem[97][3] ));
 sg13g2_nand2_1 _23757_ (.Y(_05360_),
    .A(net1265),
    .B(_05352_));
 sg13g2_o21ai_1 _23758_ (.B1(_05360_),
    .Y(_02133_),
    .A1(net303),
    .A2(_05359_));
 sg13g2_buf_1 _23759_ (.A(_05246_),
    .X(_05361_));
 sg13g2_nand2_1 _23760_ (.Y(_05362_),
    .A(net595),
    .B(\mem.mem_internal.code_mem[97][4] ));
 sg13g2_nand2_1 _23761_ (.Y(_05363_),
    .A(net1264),
    .B(_05352_));
 sg13g2_o21ai_1 _23762_ (.B1(_05363_),
    .Y(_02134_),
    .A1(net303),
    .A2(_05362_));
 sg13g2_nand2_1 _23763_ (.Y(_05364_),
    .A(_05361_),
    .B(\mem.mem_internal.code_mem[97][5] ));
 sg13g2_nand2_1 _23764_ (.Y(_05365_),
    .A(net1263),
    .B(_05352_));
 sg13g2_o21ai_1 _23765_ (.B1(_05365_),
    .Y(_02135_),
    .A1(_05353_),
    .A2(_05364_));
 sg13g2_nand2_1 _23766_ (.Y(_05366_),
    .A(net595),
    .B(\mem.mem_internal.code_mem[97][6] ));
 sg13g2_nand2_1 _23767_ (.Y(_05367_),
    .A(net1262),
    .B(_05352_));
 sg13g2_o21ai_1 _23768_ (.B1(_05367_),
    .Y(_02136_),
    .A1(net303),
    .A2(_05366_));
 sg13g2_nand2_1 _23769_ (.Y(_05368_),
    .A(net595),
    .B(\mem.mem_internal.code_mem[97][7] ));
 sg13g2_nand2_1 _23770_ (.Y(_05369_),
    .A(net1261),
    .B(_05352_));
 sg13g2_o21ai_1 _23771_ (.B1(_05369_),
    .Y(_02137_),
    .A1(net303),
    .A2(_05368_));
 sg13g2_nand2_1 _23772_ (.Y(_05370_),
    .A(net1193),
    .B(\mem.mem_internal.code_mem[98][0] ));
 sg13g2_nor2_1 _23773_ (.A(_10300_),
    .B(net527),
    .Y(_05371_));
 sg13g2_buf_2 _23774_ (.A(_05371_),
    .X(_05372_));
 sg13g2_buf_1 _23775_ (.A(_05372_),
    .X(_05373_));
 sg13g2_nand2_1 _23776_ (.Y(_05374_),
    .A(_10252_),
    .B(_05373_));
 sg13g2_o21ai_1 _23777_ (.B1(_05374_),
    .Y(_02138_),
    .A1(_05370_),
    .A2(net302));
 sg13g2_nand2_1 _23778_ (.Y(_05375_),
    .A(net595),
    .B(\mem.mem_internal.code_mem[98][1] ));
 sg13g2_nand2_1 _23779_ (.Y(_05376_),
    .A(_10257_),
    .B(net302));
 sg13g2_o21ai_1 _23780_ (.B1(_05376_),
    .Y(_02139_),
    .A1(net302),
    .A2(_05375_));
 sg13g2_nand2_1 _23781_ (.Y(_05377_),
    .A(net595),
    .B(\mem.mem_internal.code_mem[98][2] ));
 sg13g2_nand2_1 _23782_ (.Y(_05378_),
    .A(net1266),
    .B(_05372_));
 sg13g2_o21ai_1 _23783_ (.B1(_05378_),
    .Y(_02140_),
    .A1(net302),
    .A2(_05377_));
 sg13g2_nand2_1 _23784_ (.Y(_05379_),
    .A(net595),
    .B(\mem.mem_internal.code_mem[98][3] ));
 sg13g2_nand2_1 _23785_ (.Y(_05380_),
    .A(_10268_),
    .B(_05372_));
 sg13g2_o21ai_1 _23786_ (.B1(_05380_),
    .Y(_02141_),
    .A1(net302),
    .A2(_05379_));
 sg13g2_nand2_1 _23787_ (.Y(_05381_),
    .A(net595),
    .B(\mem.mem_internal.code_mem[98][4] ));
 sg13g2_nand2_1 _23788_ (.Y(_05382_),
    .A(_10273_),
    .B(_05372_));
 sg13g2_o21ai_1 _23789_ (.B1(_05382_),
    .Y(_02142_),
    .A1(net302),
    .A2(_05381_));
 sg13g2_nand2_1 _23790_ (.Y(_05383_),
    .A(_05361_),
    .B(\mem.mem_internal.code_mem[98][5] ));
 sg13g2_nand2_1 _23791_ (.Y(_05384_),
    .A(_10278_),
    .B(_05372_));
 sg13g2_o21ai_1 _23792_ (.B1(_05384_),
    .Y(_02143_),
    .A1(_05373_),
    .A2(_05383_));
 sg13g2_nand2_1 _23793_ (.Y(_05385_),
    .A(net595),
    .B(\mem.mem_internal.code_mem[98][6] ));
 sg13g2_nand2_1 _23794_ (.Y(_05386_),
    .A(_10283_),
    .B(_05372_));
 sg13g2_o21ai_1 _23795_ (.B1(_05386_),
    .Y(_02144_),
    .A1(net302),
    .A2(_05385_));
 sg13g2_buf_1 _23796_ (.A(_05246_),
    .X(_05387_));
 sg13g2_nand2_1 _23797_ (.Y(_05388_),
    .A(net594),
    .B(\mem.mem_internal.code_mem[98][7] ));
 sg13g2_nand2_1 _23798_ (.Y(_05389_),
    .A(_10288_),
    .B(_05372_));
 sg13g2_o21ai_1 _23799_ (.B1(_05389_),
    .Y(_02145_),
    .A1(net302),
    .A2(_05388_));
 sg13g2_nand2_1 _23800_ (.Y(_05390_),
    .A(net1193),
    .B(\mem.mem_internal.code_mem[99][0] ));
 sg13g2_nor2_1 _23801_ (.A(_10300_),
    .B(net526),
    .Y(_05391_));
 sg13g2_buf_2 _23802_ (.A(_05391_),
    .X(_05392_));
 sg13g2_buf_1 _23803_ (.A(_05392_),
    .X(_05393_));
 sg13g2_nand2_1 _23804_ (.Y(_05394_),
    .A(net1268),
    .B(_05393_));
 sg13g2_o21ai_1 _23805_ (.B1(_05394_),
    .Y(_02146_),
    .A1(_05390_),
    .A2(_05393_));
 sg13g2_nand2_1 _23806_ (.Y(_05395_),
    .A(net594),
    .B(\mem.mem_internal.code_mem[99][1] ));
 sg13g2_nand2_1 _23807_ (.Y(_05396_),
    .A(_10257_),
    .B(net301));
 sg13g2_o21ai_1 _23808_ (.B1(_05396_),
    .Y(_02147_),
    .A1(net301),
    .A2(_05395_));
 sg13g2_nand2_1 _23809_ (.Y(_05397_),
    .A(net594),
    .B(\mem.mem_internal.code_mem[99][2] ));
 sg13g2_nand2_1 _23810_ (.Y(_05398_),
    .A(_10263_),
    .B(_05392_));
 sg13g2_o21ai_1 _23811_ (.B1(_05398_),
    .Y(_02148_),
    .A1(net301),
    .A2(_05397_));
 sg13g2_nand2_1 _23812_ (.Y(_05399_),
    .A(_05387_),
    .B(\mem.mem_internal.code_mem[99][3] ));
 sg13g2_nand2_1 _23813_ (.Y(_05400_),
    .A(net1265),
    .B(_05392_));
 sg13g2_o21ai_1 _23814_ (.B1(_05400_),
    .Y(_02149_),
    .A1(net301),
    .A2(_05399_));
 sg13g2_nand2_1 _23815_ (.Y(_05401_),
    .A(net594),
    .B(\mem.mem_internal.code_mem[99][4] ));
 sg13g2_nand2_1 _23816_ (.Y(_05402_),
    .A(net1264),
    .B(_05392_));
 sg13g2_o21ai_1 _23817_ (.B1(_05402_),
    .Y(_02150_),
    .A1(net301),
    .A2(_05401_));
 sg13g2_nand2_1 _23818_ (.Y(_05403_),
    .A(_05387_),
    .B(\mem.mem_internal.code_mem[99][5] ));
 sg13g2_nand2_1 _23819_ (.Y(_05404_),
    .A(net1263),
    .B(_05392_));
 sg13g2_o21ai_1 _23820_ (.B1(_05404_),
    .Y(_02151_),
    .A1(net301),
    .A2(_05403_));
 sg13g2_nand2_1 _23821_ (.Y(_05405_),
    .A(net594),
    .B(\mem.mem_internal.code_mem[99][6] ));
 sg13g2_nand2_1 _23822_ (.Y(_05406_),
    .A(net1262),
    .B(_05392_));
 sg13g2_o21ai_1 _23823_ (.B1(_05406_),
    .Y(_02152_),
    .A1(net301),
    .A2(_05405_));
 sg13g2_nand2_1 _23824_ (.Y(_05407_),
    .A(net594),
    .B(\mem.mem_internal.code_mem[99][7] ));
 sg13g2_nand2_1 _23825_ (.Y(_05408_),
    .A(net1261),
    .B(_05392_));
 sg13g2_o21ai_1 _23826_ (.B1(_05408_),
    .Y(_02153_),
    .A1(net301),
    .A2(_05407_));
 sg13g2_nand2_1 _23827_ (.Y(_05409_),
    .A(net1193),
    .B(\mem.mem_internal.code_mem[9][0] ));
 sg13g2_nor2_1 _23828_ (.A(_10246_),
    .B(_10423_),
    .Y(_05410_));
 sg13g2_buf_2 _23829_ (.A(_05410_),
    .X(_05411_));
 sg13g2_buf_1 _23830_ (.A(_05411_),
    .X(_05412_));
 sg13g2_nand2_1 _23831_ (.Y(_05413_),
    .A(net1268),
    .B(net300));
 sg13g2_o21ai_1 _23832_ (.B1(_05413_),
    .Y(_02154_),
    .A1(_05409_),
    .A2(_05412_));
 sg13g2_nand2_1 _23833_ (.Y(_05414_),
    .A(net594),
    .B(\mem.mem_internal.code_mem[9][1] ));
 sg13g2_nand2_1 _23834_ (.Y(_05415_),
    .A(net1267),
    .B(net300));
 sg13g2_o21ai_1 _23835_ (.B1(_05415_),
    .Y(_02155_),
    .A1(net300),
    .A2(_05414_));
 sg13g2_nand2_1 _23836_ (.Y(_05416_),
    .A(net594),
    .B(\mem.mem_internal.code_mem[9][2] ));
 sg13g2_nand2_1 _23837_ (.Y(_05417_),
    .A(net1266),
    .B(_05411_));
 sg13g2_o21ai_1 _23838_ (.B1(_05417_),
    .Y(_02156_),
    .A1(net300),
    .A2(_05416_));
 sg13g2_buf_1 _23839_ (.A(_05246_),
    .X(_05418_));
 sg13g2_nand2_1 _23840_ (.Y(_05419_),
    .A(net593),
    .B(\mem.mem_internal.code_mem[9][3] ));
 sg13g2_nand2_1 _23841_ (.Y(_05420_),
    .A(net1265),
    .B(_05411_));
 sg13g2_o21ai_1 _23842_ (.B1(_05420_),
    .Y(_02157_),
    .A1(_05412_),
    .A2(_05419_));
 sg13g2_nand2_1 _23843_ (.Y(_05421_),
    .A(net593),
    .B(\mem.mem_internal.code_mem[9][4] ));
 sg13g2_nand2_1 _23844_ (.Y(_05422_),
    .A(net1264),
    .B(_05411_));
 sg13g2_o21ai_1 _23845_ (.B1(_05422_),
    .Y(_02158_),
    .A1(net300),
    .A2(_05421_));
 sg13g2_nand2_1 _23846_ (.Y(_05423_),
    .A(net593),
    .B(\mem.mem_internal.code_mem[9][5] ));
 sg13g2_nand2_1 _23847_ (.Y(_05424_),
    .A(net1263),
    .B(_05411_));
 sg13g2_o21ai_1 _23848_ (.B1(_05424_),
    .Y(_02159_),
    .A1(net300),
    .A2(_05423_));
 sg13g2_nand2_1 _23849_ (.Y(_05425_),
    .A(_05418_),
    .B(\mem.mem_internal.code_mem[9][6] ));
 sg13g2_nand2_1 _23850_ (.Y(_05426_),
    .A(net1262),
    .B(_05411_));
 sg13g2_o21ai_1 _23851_ (.B1(_05426_),
    .Y(_02160_),
    .A1(net300),
    .A2(_05425_));
 sg13g2_nand2_1 _23852_ (.Y(_05427_),
    .A(_05418_),
    .B(\mem.mem_internal.code_mem[9][7] ));
 sg13g2_nand2_1 _23853_ (.Y(_05428_),
    .A(net1261),
    .B(_05411_));
 sg13g2_o21ai_1 _23854_ (.B1(_05428_),
    .Y(_02161_),
    .A1(net300),
    .A2(_05427_));
 sg13g2_nand2_1 _23855_ (.Y(_05429_),
    .A(_10114_),
    .B(_10229_));
 sg13g2_inv_1 _23856_ (.Y(_05430_),
    .A(_00070_));
 sg13g2_nor3_1 _23857_ (.A(net1296),
    .B(_10034_),
    .C(_10032_),
    .Y(_05431_));
 sg13g2_buf_1 _23858_ (.A(_05431_),
    .X(_05432_));
 sg13g2_and3_1 _23859_ (.X(_05433_),
    .A(_05430_),
    .B(_10241_),
    .C(_05432_));
 sg13g2_buf_1 _23860_ (.A(_05433_),
    .X(_05434_));
 sg13g2_nand2_1 _23861_ (.Y(_05435_),
    .A(_10230_),
    .B(_05434_));
 sg13g2_buf_2 _23862_ (.A(_05435_),
    .X(_05436_));
 sg13g2_nor2_1 _23863_ (.A(_05429_),
    .B(_05436_),
    .Y(_05437_));
 sg13g2_buf_1 _23864_ (.A(_05437_),
    .X(_05438_));
 sg13g2_buf_1 _23865_ (.A(_05438_),
    .X(_05439_));
 sg13g2_nand2_1 _23866_ (.Y(_05440_),
    .A(net593),
    .B(\mem.mem_internal.data_mem[0][0] ));
 sg13g2_buf_1 _23867_ (.A(\mem.data_in[0] ),
    .X(_05441_));
 sg13g2_buf_1 _23868_ (.A(net1292),
    .X(_05442_));
 sg13g2_nand2_1 _23869_ (.Y(_05443_),
    .A(net1260),
    .B(net438));
 sg13g2_o21ai_1 _23870_ (.B1(_05443_),
    .Y(_02164_),
    .A1(net438),
    .A2(_05440_));
 sg13g2_nand2_1 _23871_ (.Y(_05444_),
    .A(net593),
    .B(\mem.mem_internal.data_mem[0][1] ));
 sg13g2_buf_1 _23872_ (.A(\mem.data_in[1] ),
    .X(_05445_));
 sg13g2_buf_1 _23873_ (.A(_05445_),
    .X(_05446_));
 sg13g2_nand2_1 _23874_ (.Y(_05447_),
    .A(net1259),
    .B(net438));
 sg13g2_o21ai_1 _23875_ (.B1(_05447_),
    .Y(_02165_),
    .A1(net438),
    .A2(_05444_));
 sg13g2_nand2_1 _23876_ (.Y(_05448_),
    .A(net593),
    .B(\mem.mem_internal.data_mem[0][2] ));
 sg13g2_buf_1 _23877_ (.A(\mem.data_in[2] ),
    .X(_05449_));
 sg13g2_buf_1 _23878_ (.A(net1290),
    .X(_05450_));
 sg13g2_nand2_1 _23879_ (.Y(_05451_),
    .A(net1258),
    .B(_05438_));
 sg13g2_o21ai_1 _23880_ (.B1(_05451_),
    .Y(_02166_),
    .A1(_05439_),
    .A2(_05448_));
 sg13g2_nand2_1 _23881_ (.Y(_05452_),
    .A(net593),
    .B(\mem.mem_internal.data_mem[0][3] ));
 sg13g2_buf_1 _23882_ (.A(\mem.data_in[3] ),
    .X(_05453_));
 sg13g2_buf_1 _23883_ (.A(net1289),
    .X(_05454_));
 sg13g2_nand2_1 _23884_ (.Y(_05455_),
    .A(net1257),
    .B(_05438_));
 sg13g2_o21ai_1 _23885_ (.B1(_05455_),
    .Y(_02167_),
    .A1(net438),
    .A2(_05452_));
 sg13g2_nand2_1 _23886_ (.Y(_05456_),
    .A(net593),
    .B(\mem.mem_internal.data_mem[0][4] ));
 sg13g2_buf_1 _23887_ (.A(\mem.data_in[4] ),
    .X(_05457_));
 sg13g2_buf_1 _23888_ (.A(net1288),
    .X(_05458_));
 sg13g2_nand2_1 _23889_ (.Y(_05459_),
    .A(net1256),
    .B(_05438_));
 sg13g2_o21ai_1 _23890_ (.B1(_05459_),
    .Y(_02168_),
    .A1(net438),
    .A2(_05456_));
 sg13g2_buf_1 _23891_ (.A(_04431_),
    .X(_05460_));
 sg13g2_buf_1 _23892_ (.A(_05460_),
    .X(_05461_));
 sg13g2_nand2_1 _23893_ (.Y(_05462_),
    .A(net592),
    .B(\mem.mem_internal.data_mem[0][5] ));
 sg13g2_buf_1 _23894_ (.A(\mem.data_in[5] ),
    .X(_05463_));
 sg13g2_buf_1 _23895_ (.A(net1287),
    .X(_05464_));
 sg13g2_nand2_1 _23896_ (.Y(_05465_),
    .A(net1255),
    .B(_05438_));
 sg13g2_o21ai_1 _23897_ (.B1(_05465_),
    .Y(_02169_),
    .A1(net438),
    .A2(_05462_));
 sg13g2_nand2_1 _23898_ (.Y(_05466_),
    .A(net592),
    .B(\mem.mem_internal.data_mem[0][6] ));
 sg13g2_buf_1 _23899_ (.A(\mem.data_in[6] ),
    .X(_05467_));
 sg13g2_buf_1 _23900_ (.A(net1286),
    .X(_05468_));
 sg13g2_nand2_1 _23901_ (.Y(_05469_),
    .A(net1254),
    .B(_05438_));
 sg13g2_o21ai_1 _23902_ (.B1(_05469_),
    .Y(_02170_),
    .A1(net438),
    .A2(_05466_));
 sg13g2_nand2_1 _23903_ (.Y(_05470_),
    .A(net592),
    .B(\mem.mem_internal.data_mem[0][7] ));
 sg13g2_buf_2 _23904_ (.A(\mem.data_in[7] ),
    .X(_05471_));
 sg13g2_buf_1 _23905_ (.A(net1285),
    .X(_05472_));
 sg13g2_nand2_1 _23906_ (.Y(_05473_),
    .A(net1253),
    .B(_05438_));
 sg13g2_o21ai_1 _23907_ (.B1(_05473_),
    .Y(_02171_),
    .A1(_05439_),
    .A2(_05470_));
 sg13g2_nand2b_1 _23908_ (.Y(_05474_),
    .B(net1271),
    .A_N(net1293));
 sg13g2_buf_1 _23909_ (.A(_05474_),
    .X(_05475_));
 sg13g2_nand2_1 _23910_ (.Y(_05476_),
    .A(_10347_),
    .B(_05434_));
 sg13g2_buf_2 _23911_ (.A(_05476_),
    .X(_05477_));
 sg13g2_nor3_1 _23912_ (.A(net1269),
    .B(_05475_),
    .C(_05477_),
    .Y(_05478_));
 sg13g2_buf_2 _23913_ (.A(_05478_),
    .X(_05479_));
 sg13g2_buf_1 _23914_ (.A(_05479_),
    .X(_05480_));
 sg13g2_nand2_1 _23915_ (.Y(_05481_),
    .A(net592),
    .B(\mem.mem_internal.data_mem[10][0] ));
 sg13g2_nand2_1 _23916_ (.Y(_05482_),
    .A(net1260),
    .B(net437));
 sg13g2_o21ai_1 _23917_ (.B1(_05482_),
    .Y(_02172_),
    .A1(net437),
    .A2(_05481_));
 sg13g2_nand2_1 _23918_ (.Y(_05483_),
    .A(net592),
    .B(\mem.mem_internal.data_mem[10][1] ));
 sg13g2_nand2_1 _23919_ (.Y(_05484_),
    .A(_05446_),
    .B(net437));
 sg13g2_o21ai_1 _23920_ (.B1(_05484_),
    .Y(_02173_),
    .A1(_05480_),
    .A2(_05483_));
 sg13g2_nand2_1 _23921_ (.Y(_05485_),
    .A(net592),
    .B(\mem.mem_internal.data_mem[10][2] ));
 sg13g2_nand2_1 _23922_ (.Y(_05486_),
    .A(net1258),
    .B(_05479_));
 sg13g2_o21ai_1 _23923_ (.B1(_05486_),
    .Y(_02174_),
    .A1(net437),
    .A2(_05485_));
 sg13g2_nand2_1 _23924_ (.Y(_05487_),
    .A(_05461_),
    .B(\mem.mem_internal.data_mem[10][3] ));
 sg13g2_nand2_1 _23925_ (.Y(_05488_),
    .A(net1257),
    .B(_05479_));
 sg13g2_o21ai_1 _23926_ (.B1(_05488_),
    .Y(_02175_),
    .A1(net437),
    .A2(_05487_));
 sg13g2_nand2_1 _23927_ (.Y(_05489_),
    .A(net592),
    .B(\mem.mem_internal.data_mem[10][4] ));
 sg13g2_nand2_1 _23928_ (.Y(_05490_),
    .A(_05458_),
    .B(_05479_));
 sg13g2_o21ai_1 _23929_ (.B1(_05490_),
    .Y(_02176_),
    .A1(net437),
    .A2(_05489_));
 sg13g2_nand2_1 _23930_ (.Y(_05491_),
    .A(net592),
    .B(\mem.mem_internal.data_mem[10][5] ));
 sg13g2_nand2_1 _23931_ (.Y(_05492_),
    .A(_05464_),
    .B(_05479_));
 sg13g2_o21ai_1 _23932_ (.B1(_05492_),
    .Y(_02177_),
    .A1(_05480_),
    .A2(_05491_));
 sg13g2_nand2_1 _23933_ (.Y(_05493_),
    .A(_05461_),
    .B(\mem.mem_internal.data_mem[10][6] ));
 sg13g2_nand2_1 _23934_ (.Y(_05494_),
    .A(net1254),
    .B(_05479_));
 sg13g2_o21ai_1 _23935_ (.B1(_05494_),
    .Y(_02178_),
    .A1(net437),
    .A2(_05493_));
 sg13g2_buf_1 _23936_ (.A(_05460_),
    .X(_05495_));
 sg13g2_nand2_1 _23937_ (.Y(_05496_),
    .A(net591),
    .B(\mem.mem_internal.data_mem[10][7] ));
 sg13g2_nand2_1 _23938_ (.Y(_05497_),
    .A(net1253),
    .B(_05479_));
 sg13g2_o21ai_1 _23939_ (.B1(_05497_),
    .Y(_02179_),
    .A1(net437),
    .A2(_05496_));
 sg13g2_nand3_1 _23940_ (.B(net1294),
    .C(_05434_),
    .A(net1295),
    .Y(_05498_));
 sg13g2_buf_2 _23941_ (.A(_05498_),
    .X(_05499_));
 sg13g2_nor3_1 _23942_ (.A(net1269),
    .B(_05475_),
    .C(_05499_),
    .Y(_05500_));
 sg13g2_buf_2 _23943_ (.A(_05500_),
    .X(_05501_));
 sg13g2_buf_1 _23944_ (.A(_05501_),
    .X(_05502_));
 sg13g2_nand2_1 _23945_ (.Y(_05503_),
    .A(net591),
    .B(\mem.mem_internal.data_mem[11][0] ));
 sg13g2_nand2_1 _23946_ (.Y(_05504_),
    .A(net1260),
    .B(net436));
 sg13g2_o21ai_1 _23947_ (.B1(_05504_),
    .Y(_02180_),
    .A1(_05502_),
    .A2(_05503_));
 sg13g2_nand2_1 _23948_ (.Y(_05505_),
    .A(net591),
    .B(\mem.mem_internal.data_mem[11][1] ));
 sg13g2_nand2_1 _23949_ (.Y(_05506_),
    .A(net1259),
    .B(net436));
 sg13g2_o21ai_1 _23950_ (.B1(_05506_),
    .Y(_02181_),
    .A1(net436),
    .A2(_05505_));
 sg13g2_nand2_1 _23951_ (.Y(_05507_),
    .A(net591),
    .B(\mem.mem_internal.data_mem[11][2] ));
 sg13g2_nand2_1 _23952_ (.Y(_05508_),
    .A(net1258),
    .B(_05501_));
 sg13g2_o21ai_1 _23953_ (.B1(_05508_),
    .Y(_02182_),
    .A1(net436),
    .A2(_05507_));
 sg13g2_nand2_1 _23954_ (.Y(_05509_),
    .A(net591),
    .B(\mem.mem_internal.data_mem[11][3] ));
 sg13g2_nand2_1 _23955_ (.Y(_05510_),
    .A(_05454_),
    .B(_05501_));
 sg13g2_o21ai_1 _23956_ (.B1(_05510_),
    .Y(_02183_),
    .A1(net436),
    .A2(_05509_));
 sg13g2_nand2_1 _23957_ (.Y(_05511_),
    .A(net591),
    .B(\mem.mem_internal.data_mem[11][4] ));
 sg13g2_nand2_1 _23958_ (.Y(_05512_),
    .A(_05458_),
    .B(_05501_));
 sg13g2_o21ai_1 _23959_ (.B1(_05512_),
    .Y(_02184_),
    .A1(net436),
    .A2(_05511_));
 sg13g2_nand2_1 _23960_ (.Y(_05513_),
    .A(_05495_),
    .B(\mem.mem_internal.data_mem[11][5] ));
 sg13g2_nand2_1 _23961_ (.Y(_05514_),
    .A(_05464_),
    .B(_05501_));
 sg13g2_o21ai_1 _23962_ (.B1(_05514_),
    .Y(_02185_),
    .A1(net436),
    .A2(_05513_));
 sg13g2_nand2_1 _23963_ (.Y(_05515_),
    .A(_05495_),
    .B(\mem.mem_internal.data_mem[11][6] ));
 sg13g2_nand2_1 _23964_ (.Y(_05516_),
    .A(net1254),
    .B(_05501_));
 sg13g2_o21ai_1 _23965_ (.B1(_05516_),
    .Y(_02186_),
    .A1(_05502_),
    .A2(_05515_));
 sg13g2_nand2_1 _23966_ (.Y(_05517_),
    .A(net591),
    .B(\mem.mem_internal.data_mem[11][7] ));
 sg13g2_nand2_1 _23967_ (.Y(_05518_),
    .A(_05472_),
    .B(_05501_));
 sg13g2_o21ai_1 _23968_ (.B1(_05518_),
    .Y(_02187_),
    .A1(net436),
    .A2(_05517_));
 sg13g2_inv_1 _23969_ (.Y(_05519_),
    .A(_00071_));
 sg13g2_nand3_1 _23970_ (.B(net1271),
    .C(_05519_),
    .A(_10114_),
    .Y(_05520_));
 sg13g2_buf_1 _23971_ (.A(_05520_),
    .X(_05521_));
 sg13g2_nor2_1 _23972_ (.A(_05436_),
    .B(_05521_),
    .Y(_05522_));
 sg13g2_buf_2 _23973_ (.A(_05522_),
    .X(_05523_));
 sg13g2_buf_1 _23974_ (.A(_05523_),
    .X(_05524_));
 sg13g2_nand2_1 _23975_ (.Y(_05525_),
    .A(net591),
    .B(\mem.mem_internal.data_mem[12][0] ));
 sg13g2_nand2_1 _23976_ (.Y(_05526_),
    .A(net1260),
    .B(net435));
 sg13g2_o21ai_1 _23977_ (.B1(_05526_),
    .Y(_02188_),
    .A1(net435),
    .A2(_05525_));
 sg13g2_buf_1 _23978_ (.A(_05460_),
    .X(_05527_));
 sg13g2_nand2_1 _23979_ (.Y(_05528_),
    .A(net590),
    .B(\mem.mem_internal.data_mem[12][1] ));
 sg13g2_nand2_1 _23980_ (.Y(_05529_),
    .A(net1259),
    .B(_05524_));
 sg13g2_o21ai_1 _23981_ (.B1(_05529_),
    .Y(_02189_),
    .A1(_05524_),
    .A2(_05528_));
 sg13g2_nand2_1 _23982_ (.Y(_05530_),
    .A(net590),
    .B(\mem.mem_internal.data_mem[12][2] ));
 sg13g2_nand2_1 _23983_ (.Y(_05531_),
    .A(net1258),
    .B(_05523_));
 sg13g2_o21ai_1 _23984_ (.B1(_05531_),
    .Y(_02190_),
    .A1(net435),
    .A2(_05530_));
 sg13g2_nand2_1 _23985_ (.Y(_05532_),
    .A(net590),
    .B(\mem.mem_internal.data_mem[12][3] ));
 sg13g2_nand2_1 _23986_ (.Y(_05533_),
    .A(net1257),
    .B(_05523_));
 sg13g2_o21ai_1 _23987_ (.B1(_05533_),
    .Y(_02191_),
    .A1(net435),
    .A2(_05532_));
 sg13g2_nand2_1 _23988_ (.Y(_05534_),
    .A(net590),
    .B(\mem.mem_internal.data_mem[12][4] ));
 sg13g2_nand2_1 _23989_ (.Y(_05535_),
    .A(net1256),
    .B(_05523_));
 sg13g2_o21ai_1 _23990_ (.B1(_05535_),
    .Y(_02192_),
    .A1(net435),
    .A2(_05534_));
 sg13g2_nand2_1 _23991_ (.Y(_05536_),
    .A(_05527_),
    .B(\mem.mem_internal.data_mem[12][5] ));
 sg13g2_nand2_1 _23992_ (.Y(_05537_),
    .A(net1255),
    .B(_05523_));
 sg13g2_o21ai_1 _23993_ (.B1(_05537_),
    .Y(_02193_),
    .A1(net435),
    .A2(_05536_));
 sg13g2_nand2_1 _23994_ (.Y(_05538_),
    .A(net590),
    .B(\mem.mem_internal.data_mem[12][6] ));
 sg13g2_nand2_1 _23995_ (.Y(_05539_),
    .A(net1254),
    .B(_05523_));
 sg13g2_o21ai_1 _23996_ (.B1(_05539_),
    .Y(_02194_),
    .A1(net435),
    .A2(_05538_));
 sg13g2_nand2_1 _23997_ (.Y(_05540_),
    .A(net590),
    .B(\mem.mem_internal.data_mem[12][7] ));
 sg13g2_nand2_1 _23998_ (.Y(_05541_),
    .A(net1253),
    .B(_05523_));
 sg13g2_o21ai_1 _23999_ (.B1(_05541_),
    .Y(_02195_),
    .A1(net435),
    .A2(_05540_));
 sg13g2_nand2_1 _24000_ (.Y(_05542_),
    .A(_10323_),
    .B(_05434_));
 sg13g2_buf_2 _24001_ (.A(_05542_),
    .X(_05543_));
 sg13g2_nor2_1 _24002_ (.A(_05521_),
    .B(_05543_),
    .Y(_05544_));
 sg13g2_buf_2 _24003_ (.A(_05544_),
    .X(_05545_));
 sg13g2_buf_1 _24004_ (.A(_05545_),
    .X(_05546_));
 sg13g2_nand2_1 _24005_ (.Y(_05547_),
    .A(net590),
    .B(\mem.mem_internal.data_mem[13][0] ));
 sg13g2_nand2_1 _24006_ (.Y(_05548_),
    .A(net1260),
    .B(net434));
 sg13g2_o21ai_1 _24007_ (.B1(_05548_),
    .Y(_02196_),
    .A1(net434),
    .A2(_05547_));
 sg13g2_nand2_1 _24008_ (.Y(_05549_),
    .A(net590),
    .B(\mem.mem_internal.data_mem[13][1] ));
 sg13g2_nand2_1 _24009_ (.Y(_05550_),
    .A(net1259),
    .B(_05546_));
 sg13g2_o21ai_1 _24010_ (.B1(_05550_),
    .Y(_02197_),
    .A1(_05546_),
    .A2(_05549_));
 sg13g2_nand2_1 _24011_ (.Y(_05551_),
    .A(_05527_),
    .B(\mem.mem_internal.data_mem[13][2] ));
 sg13g2_nand2_1 _24012_ (.Y(_05552_),
    .A(net1258),
    .B(_05545_));
 sg13g2_o21ai_1 _24013_ (.B1(_05552_),
    .Y(_02198_),
    .A1(net434),
    .A2(_05551_));
 sg13g2_buf_1 _24014_ (.A(_05460_),
    .X(_05553_));
 sg13g2_nand2_1 _24015_ (.Y(_05554_),
    .A(net589),
    .B(\mem.mem_internal.data_mem[13][3] ));
 sg13g2_nand2_1 _24016_ (.Y(_05555_),
    .A(net1257),
    .B(_05545_));
 sg13g2_o21ai_1 _24017_ (.B1(_05555_),
    .Y(_02199_),
    .A1(net434),
    .A2(_05554_));
 sg13g2_nand2_1 _24018_ (.Y(_05556_),
    .A(net589),
    .B(\mem.mem_internal.data_mem[13][4] ));
 sg13g2_nand2_1 _24019_ (.Y(_05557_),
    .A(net1256),
    .B(_05545_));
 sg13g2_o21ai_1 _24020_ (.B1(_05557_),
    .Y(_02200_),
    .A1(net434),
    .A2(_05556_));
 sg13g2_nand2_1 _24021_ (.Y(_05558_),
    .A(net589),
    .B(\mem.mem_internal.data_mem[13][5] ));
 sg13g2_nand2_1 _24022_ (.Y(_05559_),
    .A(net1255),
    .B(_05545_));
 sg13g2_o21ai_1 _24023_ (.B1(_05559_),
    .Y(_02201_),
    .A1(net434),
    .A2(_05558_));
 sg13g2_nand2_1 _24024_ (.Y(_05560_),
    .A(net589),
    .B(\mem.mem_internal.data_mem[13][6] ));
 sg13g2_nand2_1 _24025_ (.Y(_05561_),
    .A(net1254),
    .B(_05545_));
 sg13g2_o21ai_1 _24026_ (.B1(_05561_),
    .Y(_02202_),
    .A1(net434),
    .A2(_05560_));
 sg13g2_nand2_1 _24027_ (.Y(_05562_),
    .A(net589),
    .B(\mem.mem_internal.data_mem[13][7] ));
 sg13g2_nand2_1 _24028_ (.Y(_05563_),
    .A(net1253),
    .B(_05545_));
 sg13g2_o21ai_1 _24029_ (.B1(_05563_),
    .Y(_02203_),
    .A1(net434),
    .A2(_05562_));
 sg13g2_nor2_1 _24030_ (.A(_05477_),
    .B(_05521_),
    .Y(_05564_));
 sg13g2_buf_2 _24031_ (.A(_05564_),
    .X(_05565_));
 sg13g2_buf_1 _24032_ (.A(_05565_),
    .X(_05566_));
 sg13g2_nand2_1 _24033_ (.Y(_05567_),
    .A(net589),
    .B(\mem.mem_internal.data_mem[14][0] ));
 sg13g2_nand2_1 _24034_ (.Y(_05568_),
    .A(_05442_),
    .B(net433));
 sg13g2_o21ai_1 _24035_ (.B1(_05568_),
    .Y(_02204_),
    .A1(net433),
    .A2(_05567_));
 sg13g2_nand2_1 _24036_ (.Y(_05569_),
    .A(net589),
    .B(\mem.mem_internal.data_mem[14][1] ));
 sg13g2_nand2_1 _24037_ (.Y(_05570_),
    .A(net1259),
    .B(net433));
 sg13g2_o21ai_1 _24038_ (.B1(_05570_),
    .Y(_02205_),
    .A1(net433),
    .A2(_05569_));
 sg13g2_nand2_1 _24039_ (.Y(_05571_),
    .A(_05553_),
    .B(\mem.mem_internal.data_mem[14][2] ));
 sg13g2_nand2_1 _24040_ (.Y(_05572_),
    .A(_05450_),
    .B(_05565_));
 sg13g2_o21ai_1 _24041_ (.B1(_05572_),
    .Y(_02206_),
    .A1(_05566_),
    .A2(_05571_));
 sg13g2_nand2_1 _24042_ (.Y(_05573_),
    .A(_05553_),
    .B(\mem.mem_internal.data_mem[14][3] ));
 sg13g2_nand2_1 _24043_ (.Y(_05574_),
    .A(_05454_),
    .B(_05565_));
 sg13g2_o21ai_1 _24044_ (.B1(_05574_),
    .Y(_02207_),
    .A1(net433),
    .A2(_05573_));
 sg13g2_nand2_1 _24045_ (.Y(_05575_),
    .A(net589),
    .B(\mem.mem_internal.data_mem[14][4] ));
 sg13g2_nand2_1 _24046_ (.Y(_05576_),
    .A(net1256),
    .B(_05565_));
 sg13g2_o21ai_1 _24047_ (.B1(_05576_),
    .Y(_02208_),
    .A1(net433),
    .A2(_05575_));
 sg13g2_buf_1 _24048_ (.A(_05460_),
    .X(_05577_));
 sg13g2_nand2_1 _24049_ (.Y(_05578_),
    .A(net588),
    .B(\mem.mem_internal.data_mem[14][5] ));
 sg13g2_nand2_1 _24050_ (.Y(_05579_),
    .A(net1255),
    .B(_05565_));
 sg13g2_o21ai_1 _24051_ (.B1(_05579_),
    .Y(_02209_),
    .A1(_05566_),
    .A2(_05578_));
 sg13g2_nand2_1 _24052_ (.Y(_05580_),
    .A(net588),
    .B(\mem.mem_internal.data_mem[14][6] ));
 sg13g2_nand2_1 _24053_ (.Y(_05581_),
    .A(_05468_),
    .B(_05565_));
 sg13g2_o21ai_1 _24054_ (.B1(_05581_),
    .Y(_02210_),
    .A1(net433),
    .A2(_05580_));
 sg13g2_nand2_1 _24055_ (.Y(_05582_),
    .A(net588),
    .B(\mem.mem_internal.data_mem[14][7] ));
 sg13g2_nand2_1 _24056_ (.Y(_05583_),
    .A(net1253),
    .B(_05565_));
 sg13g2_o21ai_1 _24057_ (.B1(_05583_),
    .Y(_02211_),
    .A1(net433),
    .A2(_05582_));
 sg13g2_nor2_1 _24058_ (.A(_05499_),
    .B(_05521_),
    .Y(_05584_));
 sg13g2_buf_2 _24059_ (.A(_05584_),
    .X(_05585_));
 sg13g2_buf_1 _24060_ (.A(_05585_),
    .X(_05586_));
 sg13g2_nand2_1 _24061_ (.Y(_05587_),
    .A(net588),
    .B(\mem.mem_internal.data_mem[15][0] ));
 sg13g2_nand2_1 _24062_ (.Y(_05588_),
    .A(_05442_),
    .B(net432));
 sg13g2_o21ai_1 _24063_ (.B1(_05588_),
    .Y(_02212_),
    .A1(net432),
    .A2(_05587_));
 sg13g2_nand2_1 _24064_ (.Y(_05589_),
    .A(net588),
    .B(\mem.mem_internal.data_mem[15][1] ));
 sg13g2_nand2_1 _24065_ (.Y(_05590_),
    .A(net1259),
    .B(_05586_));
 sg13g2_o21ai_1 _24066_ (.B1(_05590_),
    .Y(_02213_),
    .A1(_05586_),
    .A2(_05589_));
 sg13g2_nand2_1 _24067_ (.Y(_05591_),
    .A(net588),
    .B(\mem.mem_internal.data_mem[15][2] ));
 sg13g2_nand2_1 _24068_ (.Y(_05592_),
    .A(_05450_),
    .B(_05585_));
 sg13g2_o21ai_1 _24069_ (.B1(_05592_),
    .Y(_02214_),
    .A1(net432),
    .A2(_05591_));
 sg13g2_nand2_1 _24070_ (.Y(_05593_),
    .A(_05577_),
    .B(\mem.mem_internal.data_mem[15][3] ));
 sg13g2_nand2_1 _24071_ (.Y(_05594_),
    .A(net1257),
    .B(_05585_));
 sg13g2_o21ai_1 _24072_ (.B1(_05594_),
    .Y(_02215_),
    .A1(net432),
    .A2(_05593_));
 sg13g2_nand2_1 _24073_ (.Y(_05595_),
    .A(net588),
    .B(\mem.mem_internal.data_mem[15][4] ));
 sg13g2_nand2_1 _24074_ (.Y(_05596_),
    .A(net1256),
    .B(_05585_));
 sg13g2_o21ai_1 _24075_ (.B1(_05596_),
    .Y(_02216_),
    .A1(net432),
    .A2(_05595_));
 sg13g2_nand2_1 _24076_ (.Y(_05597_),
    .A(_05577_),
    .B(\mem.mem_internal.data_mem[15][5] ));
 sg13g2_nand2_1 _24077_ (.Y(_05598_),
    .A(net1255),
    .B(_05585_));
 sg13g2_o21ai_1 _24078_ (.B1(_05598_),
    .Y(_02217_),
    .A1(net432),
    .A2(_05597_));
 sg13g2_nand2_1 _24079_ (.Y(_05599_),
    .A(net588),
    .B(\mem.mem_internal.data_mem[15][6] ));
 sg13g2_nand2_1 _24080_ (.Y(_05600_),
    .A(_05468_),
    .B(_05585_));
 sg13g2_o21ai_1 _24081_ (.B1(_05600_),
    .Y(_02218_),
    .A1(net432),
    .A2(_05599_));
 sg13g2_buf_1 _24082_ (.A(_05460_),
    .X(_05601_));
 sg13g2_nand2_1 _24083_ (.Y(_05602_),
    .A(net587),
    .B(\mem.mem_internal.data_mem[15][7] ));
 sg13g2_nand2_1 _24084_ (.Y(_05603_),
    .A(net1253),
    .B(_05585_));
 sg13g2_o21ai_1 _24085_ (.B1(_05603_),
    .Y(_02219_),
    .A1(net432),
    .A2(_05602_));
 sg13g2_nand2_1 _24086_ (.Y(_05604_),
    .A(net1269),
    .B(_10229_));
 sg13g2_nor2_1 _24087_ (.A(_05436_),
    .B(_05604_),
    .Y(_05605_));
 sg13g2_buf_2 _24088_ (.A(_05605_),
    .X(_05606_));
 sg13g2_buf_1 _24089_ (.A(_05606_),
    .X(_05607_));
 sg13g2_nand2_1 _24090_ (.Y(_05608_),
    .A(_05601_),
    .B(\mem.mem_internal.data_mem[16][0] ));
 sg13g2_nand2_1 _24091_ (.Y(_05609_),
    .A(net1260),
    .B(_05607_));
 sg13g2_o21ai_1 _24092_ (.B1(_05609_),
    .Y(_02220_),
    .A1(_05607_),
    .A2(_05608_));
 sg13g2_nand2_1 _24093_ (.Y(_05610_),
    .A(net587),
    .B(\mem.mem_internal.data_mem[16][1] ));
 sg13g2_nand2_1 _24094_ (.Y(_05611_),
    .A(net1259),
    .B(net431));
 sg13g2_o21ai_1 _24095_ (.B1(_05611_),
    .Y(_02221_),
    .A1(net431),
    .A2(_05610_));
 sg13g2_nand2_1 _24096_ (.Y(_05612_),
    .A(net587),
    .B(\mem.mem_internal.data_mem[16][2] ));
 sg13g2_nand2_1 _24097_ (.Y(_05613_),
    .A(net1258),
    .B(_05606_));
 sg13g2_o21ai_1 _24098_ (.B1(_05613_),
    .Y(_02222_),
    .A1(net431),
    .A2(_05612_));
 sg13g2_nand2_1 _24099_ (.Y(_05614_),
    .A(net587),
    .B(\mem.mem_internal.data_mem[16][3] ));
 sg13g2_nand2_1 _24100_ (.Y(_05615_),
    .A(net1257),
    .B(_05606_));
 sg13g2_o21ai_1 _24101_ (.B1(_05615_),
    .Y(_02223_),
    .A1(net431),
    .A2(_05614_));
 sg13g2_nand2_1 _24102_ (.Y(_05616_),
    .A(net587),
    .B(\mem.mem_internal.data_mem[16][4] ));
 sg13g2_nand2_1 _24103_ (.Y(_05617_),
    .A(net1256),
    .B(_05606_));
 sg13g2_o21ai_1 _24104_ (.B1(_05617_),
    .Y(_02224_),
    .A1(net431),
    .A2(_05616_));
 sg13g2_nand2_1 _24105_ (.Y(_05618_),
    .A(net587),
    .B(\mem.mem_internal.data_mem[16][5] ));
 sg13g2_nand2_1 _24106_ (.Y(_05619_),
    .A(net1255),
    .B(_05606_));
 sg13g2_o21ai_1 _24107_ (.B1(_05619_),
    .Y(_02225_),
    .A1(net431),
    .A2(_05618_));
 sg13g2_nand2_1 _24108_ (.Y(_05620_),
    .A(_05601_),
    .B(\mem.mem_internal.data_mem[16][6] ));
 sg13g2_nand2_1 _24109_ (.Y(_05621_),
    .A(net1254),
    .B(_05606_));
 sg13g2_o21ai_1 _24110_ (.B1(_05621_),
    .Y(_02226_),
    .A1(net431),
    .A2(_05620_));
 sg13g2_nand2_1 _24111_ (.Y(_05622_),
    .A(net587),
    .B(\mem.mem_internal.data_mem[16][7] ));
 sg13g2_nand2_1 _24112_ (.Y(_05623_),
    .A(net1253),
    .B(_05606_));
 sg13g2_o21ai_1 _24113_ (.B1(_05623_),
    .Y(_02227_),
    .A1(net431),
    .A2(_05622_));
 sg13g2_nor2_1 _24114_ (.A(_05543_),
    .B(_05604_),
    .Y(_05624_));
 sg13g2_buf_2 _24115_ (.A(_05624_),
    .X(_05625_));
 sg13g2_buf_1 _24116_ (.A(_05625_),
    .X(_05626_));
 sg13g2_nand2_1 _24117_ (.Y(_05627_),
    .A(net587),
    .B(\mem.mem_internal.data_mem[17][0] ));
 sg13g2_nand2_1 _24118_ (.Y(_05628_),
    .A(net1260),
    .B(_05626_));
 sg13g2_o21ai_1 _24119_ (.B1(_05628_),
    .Y(_02228_),
    .A1(_05626_),
    .A2(_05627_));
 sg13g2_buf_1 _24120_ (.A(_05460_),
    .X(_05629_));
 sg13g2_nand2_1 _24121_ (.Y(_05630_),
    .A(net586),
    .B(\mem.mem_internal.data_mem[17][1] ));
 sg13g2_nand2_1 _24122_ (.Y(_05631_),
    .A(net1259),
    .B(net430));
 sg13g2_o21ai_1 _24123_ (.B1(_05631_),
    .Y(_02229_),
    .A1(net430),
    .A2(_05630_));
 sg13g2_nand2_1 _24124_ (.Y(_05632_),
    .A(net586),
    .B(\mem.mem_internal.data_mem[17][2] ));
 sg13g2_nand2_1 _24125_ (.Y(_05633_),
    .A(net1258),
    .B(_05625_));
 sg13g2_o21ai_1 _24126_ (.B1(_05633_),
    .Y(_02230_),
    .A1(net430),
    .A2(_05632_));
 sg13g2_nand2_1 _24127_ (.Y(_05634_),
    .A(net586),
    .B(\mem.mem_internal.data_mem[17][3] ));
 sg13g2_nand2_1 _24128_ (.Y(_05635_),
    .A(net1257),
    .B(_05625_));
 sg13g2_o21ai_1 _24129_ (.B1(_05635_),
    .Y(_02231_),
    .A1(net430),
    .A2(_05634_));
 sg13g2_nand2_1 _24130_ (.Y(_05636_),
    .A(net586),
    .B(\mem.mem_internal.data_mem[17][4] ));
 sg13g2_nand2_1 _24131_ (.Y(_05637_),
    .A(net1256),
    .B(_05625_));
 sg13g2_o21ai_1 _24132_ (.B1(_05637_),
    .Y(_02232_),
    .A1(net430),
    .A2(_05636_));
 sg13g2_nand2_1 _24133_ (.Y(_05638_),
    .A(net586),
    .B(\mem.mem_internal.data_mem[17][5] ));
 sg13g2_nand2_1 _24134_ (.Y(_05639_),
    .A(net1255),
    .B(_05625_));
 sg13g2_o21ai_1 _24135_ (.B1(_05639_),
    .Y(_02233_),
    .A1(net430),
    .A2(_05638_));
 sg13g2_nand2_1 _24136_ (.Y(_05640_),
    .A(_05629_),
    .B(\mem.mem_internal.data_mem[17][6] ));
 sg13g2_nand2_1 _24137_ (.Y(_05641_),
    .A(net1254),
    .B(_05625_));
 sg13g2_o21ai_1 _24138_ (.B1(_05641_),
    .Y(_02234_),
    .A1(net430),
    .A2(_05640_));
 sg13g2_nand2_1 _24139_ (.Y(_05642_),
    .A(net586),
    .B(\mem.mem_internal.data_mem[17][7] ));
 sg13g2_nand2_1 _24140_ (.Y(_05643_),
    .A(net1253),
    .B(_05625_));
 sg13g2_o21ai_1 _24141_ (.B1(_05643_),
    .Y(_02235_),
    .A1(net430),
    .A2(_05642_));
 sg13g2_nor2_1 _24142_ (.A(_05477_),
    .B(_05604_),
    .Y(_05644_));
 sg13g2_buf_2 _24143_ (.A(_05644_),
    .X(_05645_));
 sg13g2_buf_1 _24144_ (.A(_05645_),
    .X(_05646_));
 sg13g2_nand2_1 _24145_ (.Y(_05647_),
    .A(net586),
    .B(\mem.mem_internal.data_mem[18][0] ));
 sg13g2_nand2_1 _24146_ (.Y(_05648_),
    .A(net1260),
    .B(net429));
 sg13g2_o21ai_1 _24147_ (.B1(_05648_),
    .Y(_02236_),
    .A1(net429),
    .A2(_05647_));
 sg13g2_nand2_1 _24148_ (.Y(_05649_),
    .A(net586),
    .B(\mem.mem_internal.data_mem[18][1] ));
 sg13g2_buf_1 _24149_ (.A(net1291),
    .X(_05650_));
 sg13g2_nand2_1 _24150_ (.Y(_05651_),
    .A(_05650_),
    .B(net429));
 sg13g2_o21ai_1 _24151_ (.B1(_05651_),
    .Y(_02237_),
    .A1(net429),
    .A2(_05649_));
 sg13g2_nand2_1 _24152_ (.Y(_05652_),
    .A(_05629_),
    .B(\mem.mem_internal.data_mem[18][2] ));
 sg13g2_nand2_1 _24153_ (.Y(_05653_),
    .A(net1258),
    .B(_05645_));
 sg13g2_o21ai_1 _24154_ (.B1(_05653_),
    .Y(_02238_),
    .A1(net429),
    .A2(_05652_));
 sg13g2_buf_1 _24155_ (.A(_04431_),
    .X(_05654_));
 sg13g2_buf_1 _24156_ (.A(_05654_),
    .X(_05655_));
 sg13g2_nand2_1 _24157_ (.Y(_05656_),
    .A(_05655_),
    .B(\mem.mem_internal.data_mem[18][3] ));
 sg13g2_nand2_1 _24158_ (.Y(_05657_),
    .A(net1257),
    .B(_05645_));
 sg13g2_o21ai_1 _24159_ (.B1(_05657_),
    .Y(_02239_),
    .A1(_05646_),
    .A2(_05656_));
 sg13g2_nand2_1 _24160_ (.Y(_05658_),
    .A(net585),
    .B(\mem.mem_internal.data_mem[18][4] ));
 sg13g2_nand2_1 _24161_ (.Y(_05659_),
    .A(net1256),
    .B(_05645_));
 sg13g2_o21ai_1 _24162_ (.B1(_05659_),
    .Y(_02240_),
    .A1(net429),
    .A2(_05658_));
 sg13g2_nand2_1 _24163_ (.Y(_05660_),
    .A(net585),
    .B(\mem.mem_internal.data_mem[18][5] ));
 sg13g2_nand2_1 _24164_ (.Y(_05661_),
    .A(net1255),
    .B(_05645_));
 sg13g2_o21ai_1 _24165_ (.B1(_05661_),
    .Y(_02241_),
    .A1(net429),
    .A2(_05660_));
 sg13g2_nand2_1 _24166_ (.Y(_05662_),
    .A(_05655_),
    .B(\mem.mem_internal.data_mem[18][6] ));
 sg13g2_nand2_1 _24167_ (.Y(_05663_),
    .A(net1254),
    .B(_05645_));
 sg13g2_o21ai_1 _24168_ (.B1(_05663_),
    .Y(_02242_),
    .A1(_05646_),
    .A2(_05662_));
 sg13g2_nand2_1 _24169_ (.Y(_05664_),
    .A(net585),
    .B(\mem.mem_internal.data_mem[18][7] ));
 sg13g2_nand2_1 _24170_ (.Y(_05665_),
    .A(_05472_),
    .B(_05645_));
 sg13g2_o21ai_1 _24171_ (.B1(_05665_),
    .Y(_02243_),
    .A1(net429),
    .A2(_05664_));
 sg13g2_nor2_1 _24172_ (.A(_05499_),
    .B(_05604_),
    .Y(_05666_));
 sg13g2_buf_2 _24173_ (.A(_05666_),
    .X(_05667_));
 sg13g2_buf_1 _24174_ (.A(_05667_),
    .X(_05668_));
 sg13g2_nand2_1 _24175_ (.Y(_05669_),
    .A(net585),
    .B(\mem.mem_internal.data_mem[19][0] ));
 sg13g2_buf_1 _24176_ (.A(net1292),
    .X(_05670_));
 sg13g2_nand2_1 _24177_ (.Y(_05671_),
    .A(net1251),
    .B(net428));
 sg13g2_o21ai_1 _24178_ (.B1(_05671_),
    .Y(_02244_),
    .A1(net428),
    .A2(_05669_));
 sg13g2_nand2_1 _24179_ (.Y(_05672_),
    .A(net585),
    .B(\mem.mem_internal.data_mem[19][1] ));
 sg13g2_nand2_1 _24180_ (.Y(_05673_),
    .A(_05650_),
    .B(net428));
 sg13g2_o21ai_1 _24181_ (.B1(_05673_),
    .Y(_02245_),
    .A1(net428),
    .A2(_05672_));
 sg13g2_nand2_1 _24182_ (.Y(_05674_),
    .A(net585),
    .B(\mem.mem_internal.data_mem[19][2] ));
 sg13g2_buf_1 _24183_ (.A(net1290),
    .X(_05675_));
 sg13g2_nand2_1 _24184_ (.Y(_05676_),
    .A(net1250),
    .B(_05667_));
 sg13g2_o21ai_1 _24185_ (.B1(_05676_),
    .Y(_02246_),
    .A1(net428),
    .A2(_05674_));
 sg13g2_nand2_1 _24186_ (.Y(_05677_),
    .A(net585),
    .B(\mem.mem_internal.data_mem[19][3] ));
 sg13g2_buf_1 _24187_ (.A(net1289),
    .X(_05678_));
 sg13g2_nand2_1 _24188_ (.Y(_05679_),
    .A(net1249),
    .B(_05667_));
 sg13g2_o21ai_1 _24189_ (.B1(_05679_),
    .Y(_02247_),
    .A1(net428),
    .A2(_05677_));
 sg13g2_nand2_1 _24190_ (.Y(_05680_),
    .A(net585),
    .B(\mem.mem_internal.data_mem[19][4] ));
 sg13g2_buf_1 _24191_ (.A(net1288),
    .X(_05681_));
 sg13g2_nand2_1 _24192_ (.Y(_05682_),
    .A(_05681_),
    .B(_05667_));
 sg13g2_o21ai_1 _24193_ (.B1(_05682_),
    .Y(_02248_),
    .A1(net428),
    .A2(_05680_));
 sg13g2_buf_1 _24194_ (.A(_05654_),
    .X(_05683_));
 sg13g2_nand2_1 _24195_ (.Y(_05684_),
    .A(net584),
    .B(\mem.mem_internal.data_mem[19][5] ));
 sg13g2_buf_1 _24196_ (.A(net1287),
    .X(_05685_));
 sg13g2_nand2_1 _24197_ (.Y(_05686_),
    .A(_05685_),
    .B(_05667_));
 sg13g2_o21ai_1 _24198_ (.B1(_05686_),
    .Y(_02249_),
    .A1(_05668_),
    .A2(_05684_));
 sg13g2_nand2_1 _24199_ (.Y(_05687_),
    .A(net584),
    .B(\mem.mem_internal.data_mem[19][6] ));
 sg13g2_buf_1 _24200_ (.A(net1286),
    .X(_05688_));
 sg13g2_nand2_1 _24201_ (.Y(_05689_),
    .A(net1246),
    .B(_05667_));
 sg13g2_o21ai_1 _24202_ (.B1(_05689_),
    .Y(_02250_),
    .A1(_05668_),
    .A2(_05687_));
 sg13g2_nand2_1 _24203_ (.Y(_05690_),
    .A(net584),
    .B(\mem.mem_internal.data_mem[19][7] ));
 sg13g2_buf_1 _24204_ (.A(net1285),
    .X(_05691_));
 sg13g2_nand2_1 _24205_ (.Y(_05692_),
    .A(net1245),
    .B(_05667_));
 sg13g2_o21ai_1 _24206_ (.B1(_05692_),
    .Y(_02251_),
    .A1(net428),
    .A2(_05690_));
 sg13g2_nor2_1 _24207_ (.A(_05429_),
    .B(_05543_),
    .Y(_05693_));
 sg13g2_buf_1 _24208_ (.A(_05693_),
    .X(_05694_));
 sg13g2_buf_1 _24209_ (.A(_05694_),
    .X(_05695_));
 sg13g2_nand2_1 _24210_ (.Y(_05696_),
    .A(net584),
    .B(\mem.mem_internal.data_mem[1][0] ));
 sg13g2_nand2_1 _24211_ (.Y(_05697_),
    .A(net1251),
    .B(net427));
 sg13g2_o21ai_1 _24212_ (.B1(_05697_),
    .Y(_02252_),
    .A1(net427),
    .A2(_05696_));
 sg13g2_nand2_1 _24213_ (.Y(_05698_),
    .A(_05683_),
    .B(\mem.mem_internal.data_mem[1][1] ));
 sg13g2_nand2_1 _24214_ (.Y(_05699_),
    .A(net1252),
    .B(net427));
 sg13g2_o21ai_1 _24215_ (.B1(_05699_),
    .Y(_02253_),
    .A1(net427),
    .A2(_05698_));
 sg13g2_nand2_1 _24216_ (.Y(_05700_),
    .A(net584),
    .B(\mem.mem_internal.data_mem[1][2] ));
 sg13g2_nand2_1 _24217_ (.Y(_05701_),
    .A(net1250),
    .B(_05694_));
 sg13g2_o21ai_1 _24218_ (.B1(_05701_),
    .Y(_02254_),
    .A1(_05695_),
    .A2(_05700_));
 sg13g2_nand2_1 _24219_ (.Y(_05702_),
    .A(net584),
    .B(\mem.mem_internal.data_mem[1][3] ));
 sg13g2_nand2_1 _24220_ (.Y(_05703_),
    .A(net1249),
    .B(_05694_));
 sg13g2_o21ai_1 _24221_ (.B1(_05703_),
    .Y(_02255_),
    .A1(net427),
    .A2(_05702_));
 sg13g2_nand2_1 _24222_ (.Y(_05704_),
    .A(net584),
    .B(\mem.mem_internal.data_mem[1][4] ));
 sg13g2_nand2_1 _24223_ (.Y(_05705_),
    .A(_05681_),
    .B(_05694_));
 sg13g2_o21ai_1 _24224_ (.B1(_05705_),
    .Y(_02256_),
    .A1(net427),
    .A2(_05704_));
 sg13g2_nand2_1 _24225_ (.Y(_05706_),
    .A(net584),
    .B(\mem.mem_internal.data_mem[1][5] ));
 sg13g2_nand2_1 _24226_ (.Y(_05707_),
    .A(net1247),
    .B(_05694_));
 sg13g2_o21ai_1 _24227_ (.B1(_05707_),
    .Y(_02257_),
    .A1(_05695_),
    .A2(_05706_));
 sg13g2_nand2_1 _24228_ (.Y(_05708_),
    .A(_05683_),
    .B(\mem.mem_internal.data_mem[1][6] ));
 sg13g2_nand2_1 _24229_ (.Y(_05709_),
    .A(net1246),
    .B(_05694_));
 sg13g2_o21ai_1 _24230_ (.B1(_05709_),
    .Y(_02258_),
    .A1(net427),
    .A2(_05708_));
 sg13g2_buf_1 _24231_ (.A(_05654_),
    .X(_05710_));
 sg13g2_nand2_1 _24232_ (.Y(_05711_),
    .A(_05710_),
    .B(\mem.mem_internal.data_mem[1][7] ));
 sg13g2_nand2_1 _24233_ (.Y(_05712_),
    .A(net1245),
    .B(_05694_));
 sg13g2_o21ai_1 _24234_ (.B1(_05712_),
    .Y(_02259_),
    .A1(net427),
    .A2(_05711_));
 sg13g2_nor2_1 _24235_ (.A(net1271),
    .B(_00071_),
    .Y(_05713_));
 sg13g2_nand2_2 _24236_ (.Y(_05714_),
    .A(net1269),
    .B(_05713_));
 sg13g2_nor2_1 _24237_ (.A(_05436_),
    .B(_05714_),
    .Y(_05715_));
 sg13g2_buf_2 _24238_ (.A(_05715_),
    .X(_05716_));
 sg13g2_buf_1 _24239_ (.A(_05716_),
    .X(_05717_));
 sg13g2_nand2_1 _24240_ (.Y(_05718_),
    .A(net583),
    .B(\mem.mem_internal.data_mem[20][0] ));
 sg13g2_nand2_1 _24241_ (.Y(_05719_),
    .A(net1251),
    .B(net426));
 sg13g2_o21ai_1 _24242_ (.B1(_05719_),
    .Y(_02260_),
    .A1(net426),
    .A2(_05718_));
 sg13g2_nand2_1 _24243_ (.Y(_05720_),
    .A(net583),
    .B(\mem.mem_internal.data_mem[20][1] ));
 sg13g2_nand2_1 _24244_ (.Y(_05721_),
    .A(net1252),
    .B(net426));
 sg13g2_o21ai_1 _24245_ (.B1(_05721_),
    .Y(_02261_),
    .A1(net426),
    .A2(_05720_));
 sg13g2_nand2_1 _24246_ (.Y(_05722_),
    .A(net583),
    .B(\mem.mem_internal.data_mem[20][2] ));
 sg13g2_nand2_1 _24247_ (.Y(_05723_),
    .A(_05675_),
    .B(_05716_));
 sg13g2_o21ai_1 _24248_ (.B1(_05723_),
    .Y(_02262_),
    .A1(net426),
    .A2(_05722_));
 sg13g2_nand2_1 _24249_ (.Y(_05724_),
    .A(net583),
    .B(\mem.mem_internal.data_mem[20][3] ));
 sg13g2_nand2_1 _24250_ (.Y(_05725_),
    .A(_05678_),
    .B(_05716_));
 sg13g2_o21ai_1 _24251_ (.B1(_05725_),
    .Y(_02263_),
    .A1(net426),
    .A2(_05724_));
 sg13g2_nand2_1 _24252_ (.Y(_05726_),
    .A(net583),
    .B(\mem.mem_internal.data_mem[20][4] ));
 sg13g2_nand2_1 _24253_ (.Y(_05727_),
    .A(net1248),
    .B(_05716_));
 sg13g2_o21ai_1 _24254_ (.B1(_05727_),
    .Y(_02264_),
    .A1(_05717_),
    .A2(_05726_));
 sg13g2_nand2_1 _24255_ (.Y(_05728_),
    .A(net583),
    .B(\mem.mem_internal.data_mem[20][5] ));
 sg13g2_nand2_1 _24256_ (.Y(_05729_),
    .A(_05685_),
    .B(_05716_));
 sg13g2_o21ai_1 _24257_ (.B1(_05729_),
    .Y(_02265_),
    .A1(net426),
    .A2(_05728_));
 sg13g2_nand2_1 _24258_ (.Y(_05730_),
    .A(net583),
    .B(\mem.mem_internal.data_mem[20][6] ));
 sg13g2_nand2_1 _24259_ (.Y(_05731_),
    .A(_05688_),
    .B(_05716_));
 sg13g2_o21ai_1 _24260_ (.B1(_05731_),
    .Y(_02266_),
    .A1(net426),
    .A2(_05730_));
 sg13g2_nand2_1 _24261_ (.Y(_05732_),
    .A(_05710_),
    .B(\mem.mem_internal.data_mem[20][7] ));
 sg13g2_nand2_1 _24262_ (.Y(_05733_),
    .A(_05691_),
    .B(_05716_));
 sg13g2_o21ai_1 _24263_ (.B1(_05733_),
    .Y(_02267_),
    .A1(_05717_),
    .A2(_05732_));
 sg13g2_nor2_1 _24264_ (.A(_05543_),
    .B(_05714_),
    .Y(_05734_));
 sg13g2_buf_2 _24265_ (.A(_05734_),
    .X(_05735_));
 sg13g2_buf_1 _24266_ (.A(_05735_),
    .X(_05736_));
 sg13g2_nand2_1 _24267_ (.Y(_05737_),
    .A(net583),
    .B(\mem.mem_internal.data_mem[21][0] ));
 sg13g2_nand2_1 _24268_ (.Y(_05738_),
    .A(_05670_),
    .B(net425));
 sg13g2_o21ai_1 _24269_ (.B1(_05738_),
    .Y(_02268_),
    .A1(net425),
    .A2(_05737_));
 sg13g2_buf_1 _24270_ (.A(_05654_),
    .X(_05739_));
 sg13g2_nand2_1 _24271_ (.Y(_05740_),
    .A(net582),
    .B(\mem.mem_internal.data_mem[21][1] ));
 sg13g2_nand2_1 _24272_ (.Y(_05741_),
    .A(net1252),
    .B(net425));
 sg13g2_o21ai_1 _24273_ (.B1(_05741_),
    .Y(_02269_),
    .A1(net425),
    .A2(_05740_));
 sg13g2_nand2_1 _24274_ (.Y(_05742_),
    .A(_05739_),
    .B(\mem.mem_internal.data_mem[21][2] ));
 sg13g2_nand2_1 _24275_ (.Y(_05743_),
    .A(_05675_),
    .B(_05735_));
 sg13g2_o21ai_1 _24276_ (.B1(_05743_),
    .Y(_02270_),
    .A1(_05736_),
    .A2(_05742_));
 sg13g2_nand2_1 _24277_ (.Y(_05744_),
    .A(net582),
    .B(\mem.mem_internal.data_mem[21][3] ));
 sg13g2_nand2_1 _24278_ (.Y(_05745_),
    .A(_05678_),
    .B(_05735_));
 sg13g2_o21ai_1 _24279_ (.B1(_05745_),
    .Y(_02271_),
    .A1(net425),
    .A2(_05744_));
 sg13g2_nand2_1 _24280_ (.Y(_05746_),
    .A(net582),
    .B(\mem.mem_internal.data_mem[21][4] ));
 sg13g2_nand2_1 _24281_ (.Y(_05747_),
    .A(net1248),
    .B(_05735_));
 sg13g2_o21ai_1 _24282_ (.B1(_05747_),
    .Y(_02272_),
    .A1(_05736_),
    .A2(_05746_));
 sg13g2_nand2_1 _24283_ (.Y(_05748_),
    .A(net582),
    .B(\mem.mem_internal.data_mem[21][5] ));
 sg13g2_nand2_1 _24284_ (.Y(_05749_),
    .A(net1247),
    .B(_05735_));
 sg13g2_o21ai_1 _24285_ (.B1(_05749_),
    .Y(_02273_),
    .A1(net425),
    .A2(_05748_));
 sg13g2_nand2_1 _24286_ (.Y(_05750_),
    .A(net582),
    .B(\mem.mem_internal.data_mem[21][6] ));
 sg13g2_nand2_1 _24287_ (.Y(_05751_),
    .A(_05688_),
    .B(_05735_));
 sg13g2_o21ai_1 _24288_ (.B1(_05751_),
    .Y(_02274_),
    .A1(net425),
    .A2(_05750_));
 sg13g2_nand2_1 _24289_ (.Y(_05752_),
    .A(_05739_),
    .B(\mem.mem_internal.data_mem[21][7] ));
 sg13g2_nand2_1 _24290_ (.Y(_05753_),
    .A(_05691_),
    .B(_05735_));
 sg13g2_o21ai_1 _24291_ (.B1(_05753_),
    .Y(_02275_),
    .A1(net425),
    .A2(_05752_));
 sg13g2_nor2_1 _24292_ (.A(_05477_),
    .B(_05714_),
    .Y(_05754_));
 sg13g2_buf_1 _24293_ (.A(_05754_),
    .X(_05755_));
 sg13g2_buf_1 _24294_ (.A(_05755_),
    .X(_05756_));
 sg13g2_nand2_1 _24295_ (.Y(_05757_),
    .A(net582),
    .B(\mem.mem_internal.data_mem[22][0] ));
 sg13g2_nand2_1 _24296_ (.Y(_05758_),
    .A(_05670_),
    .B(net424));
 sg13g2_o21ai_1 _24297_ (.B1(_05758_),
    .Y(_02276_),
    .A1(net424),
    .A2(_05757_));
 sg13g2_nand2_1 _24298_ (.Y(_05759_),
    .A(net582),
    .B(\mem.mem_internal.data_mem[22][1] ));
 sg13g2_nand2_1 _24299_ (.Y(_05760_),
    .A(net1252),
    .B(net424));
 sg13g2_o21ai_1 _24300_ (.B1(_05760_),
    .Y(_02277_),
    .A1(net424),
    .A2(_05759_));
 sg13g2_nand2_1 _24301_ (.Y(_05761_),
    .A(net582),
    .B(\mem.mem_internal.data_mem[22][2] ));
 sg13g2_nand2_1 _24302_ (.Y(_05762_),
    .A(net1250),
    .B(_05755_));
 sg13g2_o21ai_1 _24303_ (.B1(_05762_),
    .Y(_02278_),
    .A1(net424),
    .A2(_05761_));
 sg13g2_buf_1 _24304_ (.A(_05654_),
    .X(_05763_));
 sg13g2_nand2_1 _24305_ (.Y(_05764_),
    .A(net581),
    .B(\mem.mem_internal.data_mem[22][3] ));
 sg13g2_nand2_1 _24306_ (.Y(_05765_),
    .A(net1249),
    .B(_05755_));
 sg13g2_o21ai_1 _24307_ (.B1(_05765_),
    .Y(_02279_),
    .A1(net424),
    .A2(_05764_));
 sg13g2_nand2_1 _24308_ (.Y(_05766_),
    .A(net581),
    .B(\mem.mem_internal.data_mem[22][4] ));
 sg13g2_nand2_1 _24309_ (.Y(_05767_),
    .A(net1248),
    .B(_05755_));
 sg13g2_o21ai_1 _24310_ (.B1(_05767_),
    .Y(_02280_),
    .A1(_05756_),
    .A2(_05766_));
 sg13g2_nand2_1 _24311_ (.Y(_05768_),
    .A(net581),
    .B(\mem.mem_internal.data_mem[22][5] ));
 sg13g2_nand2_1 _24312_ (.Y(_05769_),
    .A(net1247),
    .B(_05755_));
 sg13g2_o21ai_1 _24313_ (.B1(_05769_),
    .Y(_02281_),
    .A1(net424),
    .A2(_05768_));
 sg13g2_nand2_1 _24314_ (.Y(_05770_),
    .A(net581),
    .B(\mem.mem_internal.data_mem[22][6] ));
 sg13g2_nand2_1 _24315_ (.Y(_05771_),
    .A(net1246),
    .B(_05755_));
 sg13g2_o21ai_1 _24316_ (.B1(_05771_),
    .Y(_02282_),
    .A1(_05756_),
    .A2(_05770_));
 sg13g2_nand2_1 _24317_ (.Y(_05772_),
    .A(_05763_),
    .B(\mem.mem_internal.data_mem[22][7] ));
 sg13g2_nand2_1 _24318_ (.Y(_05773_),
    .A(net1245),
    .B(_05755_));
 sg13g2_o21ai_1 _24319_ (.B1(_05773_),
    .Y(_02283_),
    .A1(net424),
    .A2(_05772_));
 sg13g2_nor2_1 _24320_ (.A(_05499_),
    .B(_05714_),
    .Y(_05774_));
 sg13g2_buf_2 _24321_ (.A(_05774_),
    .X(_05775_));
 sg13g2_buf_1 _24322_ (.A(_05775_),
    .X(_05776_));
 sg13g2_nand2_1 _24323_ (.Y(_05777_),
    .A(net581),
    .B(\mem.mem_internal.data_mem[23][0] ));
 sg13g2_nand2_1 _24324_ (.Y(_05778_),
    .A(net1251),
    .B(net423));
 sg13g2_o21ai_1 _24325_ (.B1(_05778_),
    .Y(_02284_),
    .A1(net423),
    .A2(_05777_));
 sg13g2_nand2_1 _24326_ (.Y(_05779_),
    .A(net581),
    .B(\mem.mem_internal.data_mem[23][1] ));
 sg13g2_nand2_1 _24327_ (.Y(_05780_),
    .A(net1252),
    .B(net423));
 sg13g2_o21ai_1 _24328_ (.B1(_05780_),
    .Y(_02285_),
    .A1(net423),
    .A2(_05779_));
 sg13g2_nand2_1 _24329_ (.Y(_05781_),
    .A(net581),
    .B(\mem.mem_internal.data_mem[23][2] ));
 sg13g2_nand2_1 _24330_ (.Y(_05782_),
    .A(net1250),
    .B(_05775_));
 sg13g2_o21ai_1 _24331_ (.B1(_05782_),
    .Y(_02286_),
    .A1(net423),
    .A2(_05781_));
 sg13g2_nand2_1 _24332_ (.Y(_05783_),
    .A(net581),
    .B(\mem.mem_internal.data_mem[23][3] ));
 sg13g2_nand2_1 _24333_ (.Y(_05784_),
    .A(net1249),
    .B(_05775_));
 sg13g2_o21ai_1 _24334_ (.B1(_05784_),
    .Y(_02287_),
    .A1(net423),
    .A2(_05783_));
 sg13g2_nand2_1 _24335_ (.Y(_05785_),
    .A(_05763_),
    .B(\mem.mem_internal.data_mem[23][4] ));
 sg13g2_nand2_1 _24336_ (.Y(_05786_),
    .A(net1248),
    .B(_05775_));
 sg13g2_o21ai_1 _24337_ (.B1(_05786_),
    .Y(_02288_),
    .A1(_05776_),
    .A2(_05785_));
 sg13g2_buf_1 _24338_ (.A(_05654_),
    .X(_05787_));
 sg13g2_nand2_1 _24339_ (.Y(_05788_),
    .A(net580),
    .B(\mem.mem_internal.data_mem[23][5] ));
 sg13g2_nand2_1 _24340_ (.Y(_05789_),
    .A(net1247),
    .B(_05775_));
 sg13g2_o21ai_1 _24341_ (.B1(_05789_),
    .Y(_02289_),
    .A1(net423),
    .A2(_05788_));
 sg13g2_nand2_1 _24342_ (.Y(_05790_),
    .A(_05787_),
    .B(\mem.mem_internal.data_mem[23][6] ));
 sg13g2_nand2_1 _24343_ (.Y(_05791_),
    .A(net1246),
    .B(_05775_));
 sg13g2_o21ai_1 _24344_ (.B1(_05791_),
    .Y(_02290_),
    .A1(_05776_),
    .A2(_05790_));
 sg13g2_nand2_1 _24345_ (.Y(_05792_),
    .A(net580),
    .B(\mem.mem_internal.data_mem[23][7] ));
 sg13g2_nand2_1 _24346_ (.Y(_05793_),
    .A(net1245),
    .B(_05775_));
 sg13g2_o21ai_1 _24347_ (.B1(_05793_),
    .Y(_02291_),
    .A1(net423),
    .A2(_05792_));
 sg13g2_nand2_2 _24348_ (.Y(_05794_),
    .A(net1269),
    .B(_10395_));
 sg13g2_nor2_1 _24349_ (.A(_05436_),
    .B(_05794_),
    .Y(_05795_));
 sg13g2_buf_2 _24350_ (.A(_05795_),
    .X(_05796_));
 sg13g2_buf_1 _24351_ (.A(_05796_),
    .X(_05797_));
 sg13g2_nand2_1 _24352_ (.Y(_05798_),
    .A(net580),
    .B(\mem.mem_internal.data_mem[24][0] ));
 sg13g2_nand2_1 _24353_ (.Y(_05799_),
    .A(net1251),
    .B(net422));
 sg13g2_o21ai_1 _24354_ (.B1(_05799_),
    .Y(_02292_),
    .A1(net422),
    .A2(_05798_));
 sg13g2_nand2_1 _24355_ (.Y(_05800_),
    .A(net580),
    .B(\mem.mem_internal.data_mem[24][1] ));
 sg13g2_nand2_1 _24356_ (.Y(_05801_),
    .A(net1252),
    .B(net422));
 sg13g2_o21ai_1 _24357_ (.B1(_05801_),
    .Y(_02293_),
    .A1(net422),
    .A2(_05800_));
 sg13g2_nand2_1 _24358_ (.Y(_05802_),
    .A(net580),
    .B(\mem.mem_internal.data_mem[24][2] ));
 sg13g2_nand2_1 _24359_ (.Y(_05803_),
    .A(net1250),
    .B(_05796_));
 sg13g2_o21ai_1 _24360_ (.B1(_05803_),
    .Y(_02294_),
    .A1(net422),
    .A2(_05802_));
 sg13g2_nand2_1 _24361_ (.Y(_05804_),
    .A(net580),
    .B(\mem.mem_internal.data_mem[24][3] ));
 sg13g2_nand2_1 _24362_ (.Y(_05805_),
    .A(net1249),
    .B(_05796_));
 sg13g2_o21ai_1 _24363_ (.B1(_05805_),
    .Y(_02295_),
    .A1(net422),
    .A2(_05804_));
 sg13g2_nand2_1 _24364_ (.Y(_05806_),
    .A(_05787_),
    .B(\mem.mem_internal.data_mem[24][4] ));
 sg13g2_nand2_1 _24365_ (.Y(_05807_),
    .A(net1248),
    .B(_05796_));
 sg13g2_o21ai_1 _24366_ (.B1(_05807_),
    .Y(_02296_),
    .A1(net422),
    .A2(_05806_));
 sg13g2_nand2_1 _24367_ (.Y(_05808_),
    .A(net580),
    .B(\mem.mem_internal.data_mem[24][5] ));
 sg13g2_nand2_1 _24368_ (.Y(_05809_),
    .A(net1247),
    .B(_05796_));
 sg13g2_o21ai_1 _24369_ (.B1(_05809_),
    .Y(_02297_),
    .A1(net422),
    .A2(_05808_));
 sg13g2_nand2_1 _24370_ (.Y(_05810_),
    .A(net580),
    .B(\mem.mem_internal.data_mem[24][6] ));
 sg13g2_nand2_1 _24371_ (.Y(_05811_),
    .A(net1246),
    .B(_05796_));
 sg13g2_o21ai_1 _24372_ (.B1(_05811_),
    .Y(_02298_),
    .A1(_05797_),
    .A2(_05810_));
 sg13g2_buf_1 _24373_ (.A(_05654_),
    .X(_05812_));
 sg13g2_nand2_1 _24374_ (.Y(_05813_),
    .A(net579),
    .B(\mem.mem_internal.data_mem[24][7] ));
 sg13g2_nand2_1 _24375_ (.Y(_05814_),
    .A(net1245),
    .B(_05796_));
 sg13g2_o21ai_1 _24376_ (.B1(_05814_),
    .Y(_02299_),
    .A1(_05797_),
    .A2(_05813_));
 sg13g2_nor2_1 _24377_ (.A(_05543_),
    .B(_05794_),
    .Y(_05815_));
 sg13g2_buf_2 _24378_ (.A(_05815_),
    .X(_05816_));
 sg13g2_buf_1 _24379_ (.A(_05816_),
    .X(_05817_));
 sg13g2_nand2_1 _24380_ (.Y(_05818_),
    .A(net579),
    .B(\mem.mem_internal.data_mem[25][0] ));
 sg13g2_nand2_1 _24381_ (.Y(_05819_),
    .A(net1251),
    .B(net421));
 sg13g2_o21ai_1 _24382_ (.B1(_05819_),
    .Y(_02300_),
    .A1(net421),
    .A2(_05818_));
 sg13g2_nand2_1 _24383_ (.Y(_05820_),
    .A(net579),
    .B(\mem.mem_internal.data_mem[25][1] ));
 sg13g2_nand2_1 _24384_ (.Y(_05821_),
    .A(net1252),
    .B(net421));
 sg13g2_o21ai_1 _24385_ (.B1(_05821_),
    .Y(_02301_),
    .A1(net421),
    .A2(_05820_));
 sg13g2_nand2_1 _24386_ (.Y(_05822_),
    .A(net579),
    .B(\mem.mem_internal.data_mem[25][2] ));
 sg13g2_nand2_1 _24387_ (.Y(_05823_),
    .A(net1250),
    .B(_05816_));
 sg13g2_o21ai_1 _24388_ (.B1(_05823_),
    .Y(_02302_),
    .A1(net421),
    .A2(_05822_));
 sg13g2_nand2_1 _24389_ (.Y(_05824_),
    .A(net579),
    .B(\mem.mem_internal.data_mem[25][3] ));
 sg13g2_nand2_1 _24390_ (.Y(_05825_),
    .A(net1249),
    .B(_05816_));
 sg13g2_o21ai_1 _24391_ (.B1(_05825_),
    .Y(_02303_),
    .A1(net421),
    .A2(_05824_));
 sg13g2_nand2_1 _24392_ (.Y(_05826_),
    .A(net579),
    .B(\mem.mem_internal.data_mem[25][4] ));
 sg13g2_nand2_1 _24393_ (.Y(_05827_),
    .A(net1248),
    .B(_05816_));
 sg13g2_o21ai_1 _24394_ (.B1(_05827_),
    .Y(_02304_),
    .A1(net421),
    .A2(_05826_));
 sg13g2_nand2_1 _24395_ (.Y(_05828_),
    .A(net579),
    .B(\mem.mem_internal.data_mem[25][5] ));
 sg13g2_nand2_1 _24396_ (.Y(_05829_),
    .A(net1247),
    .B(_05816_));
 sg13g2_o21ai_1 _24397_ (.B1(_05829_),
    .Y(_02305_),
    .A1(net421),
    .A2(_05828_));
 sg13g2_nand2_1 _24398_ (.Y(_05830_),
    .A(_05812_),
    .B(\mem.mem_internal.data_mem[25][6] ));
 sg13g2_nand2_1 _24399_ (.Y(_05831_),
    .A(net1246),
    .B(_05816_));
 sg13g2_o21ai_1 _24400_ (.B1(_05831_),
    .Y(_02306_),
    .A1(_05817_),
    .A2(_05830_));
 sg13g2_nand2_1 _24401_ (.Y(_05832_),
    .A(_05812_),
    .B(\mem.mem_internal.data_mem[25][7] ));
 sg13g2_nand2_1 _24402_ (.Y(_05833_),
    .A(net1245),
    .B(_05816_));
 sg13g2_o21ai_1 _24403_ (.B1(_05833_),
    .Y(_02307_),
    .A1(_05817_),
    .A2(_05832_));
 sg13g2_nor2_1 _24404_ (.A(_05477_),
    .B(_05794_),
    .Y(_05834_));
 sg13g2_buf_2 _24405_ (.A(_05834_),
    .X(_05835_));
 sg13g2_buf_1 _24406_ (.A(_05835_),
    .X(_05836_));
 sg13g2_nand2_1 _24407_ (.Y(_05837_),
    .A(net579),
    .B(\mem.mem_internal.data_mem[26][0] ));
 sg13g2_nand2_1 _24408_ (.Y(_05838_),
    .A(net1251),
    .B(net420));
 sg13g2_o21ai_1 _24409_ (.B1(_05838_),
    .Y(_02308_),
    .A1(net420),
    .A2(_05837_));
 sg13g2_buf_1 _24410_ (.A(net1273),
    .X(_05839_));
 sg13g2_buf_1 _24411_ (.A(_05839_),
    .X(_05840_));
 sg13g2_nand2_1 _24412_ (.Y(_05841_),
    .A(net831),
    .B(\mem.mem_internal.data_mem[26][1] ));
 sg13g2_nand2_1 _24413_ (.Y(_05842_),
    .A(net1252),
    .B(net420));
 sg13g2_o21ai_1 _24414_ (.B1(_05842_),
    .Y(_02309_),
    .A1(net420),
    .A2(_05841_));
 sg13g2_nand2_1 _24415_ (.Y(_05843_),
    .A(net831),
    .B(\mem.mem_internal.data_mem[26][2] ));
 sg13g2_nand2_1 _24416_ (.Y(_05844_),
    .A(net1250),
    .B(_05835_));
 sg13g2_o21ai_1 _24417_ (.B1(_05844_),
    .Y(_02310_),
    .A1(net420),
    .A2(_05843_));
 sg13g2_nand2_1 _24418_ (.Y(_05845_),
    .A(net831),
    .B(\mem.mem_internal.data_mem[26][3] ));
 sg13g2_nand2_1 _24419_ (.Y(_05846_),
    .A(net1249),
    .B(_05835_));
 sg13g2_o21ai_1 _24420_ (.B1(_05846_),
    .Y(_02311_),
    .A1(net420),
    .A2(_05845_));
 sg13g2_nand2_1 _24421_ (.Y(_05847_),
    .A(net831),
    .B(\mem.mem_internal.data_mem[26][4] ));
 sg13g2_nand2_1 _24422_ (.Y(_05848_),
    .A(net1248),
    .B(_05835_));
 sg13g2_o21ai_1 _24423_ (.B1(_05848_),
    .Y(_02312_),
    .A1(net420),
    .A2(_05847_));
 sg13g2_nand2_1 _24424_ (.Y(_05849_),
    .A(net831),
    .B(\mem.mem_internal.data_mem[26][5] ));
 sg13g2_nand2_1 _24425_ (.Y(_05850_),
    .A(net1247),
    .B(_05835_));
 sg13g2_o21ai_1 _24426_ (.B1(_05850_),
    .Y(_02313_),
    .A1(net420),
    .A2(_05849_));
 sg13g2_nand2_1 _24427_ (.Y(_05851_),
    .A(_05840_),
    .B(\mem.mem_internal.data_mem[26][6] ));
 sg13g2_nand2_1 _24428_ (.Y(_05852_),
    .A(net1246),
    .B(_05835_));
 sg13g2_o21ai_1 _24429_ (.B1(_05852_),
    .Y(_02314_),
    .A1(_05836_),
    .A2(_05851_));
 sg13g2_nand2_1 _24430_ (.Y(_05853_),
    .A(_05840_),
    .B(\mem.mem_internal.data_mem[26][7] ));
 sg13g2_nand2_1 _24431_ (.Y(_05854_),
    .A(net1245),
    .B(_05835_));
 sg13g2_o21ai_1 _24432_ (.B1(_05854_),
    .Y(_02315_),
    .A1(_05836_),
    .A2(_05853_));
 sg13g2_nor2_1 _24433_ (.A(_05499_),
    .B(_05794_),
    .Y(_05855_));
 sg13g2_buf_2 _24434_ (.A(_05855_),
    .X(_05856_));
 sg13g2_buf_1 _24435_ (.A(_05856_),
    .X(_05857_));
 sg13g2_nand2_1 _24436_ (.Y(_05858_),
    .A(net831),
    .B(\mem.mem_internal.data_mem[27][0] ));
 sg13g2_nand2_1 _24437_ (.Y(_05859_),
    .A(net1251),
    .B(net419));
 sg13g2_o21ai_1 _24438_ (.B1(_05859_),
    .Y(_02316_),
    .A1(net419),
    .A2(_05858_));
 sg13g2_nand2_1 _24439_ (.Y(_05860_),
    .A(net831),
    .B(\mem.mem_internal.data_mem[27][1] ));
 sg13g2_buf_1 _24440_ (.A(net1291),
    .X(_05861_));
 sg13g2_nand2_1 _24441_ (.Y(_05862_),
    .A(net1244),
    .B(net419));
 sg13g2_o21ai_1 _24442_ (.B1(_05862_),
    .Y(_02317_),
    .A1(net419),
    .A2(_05860_));
 sg13g2_nand2_1 _24443_ (.Y(_05863_),
    .A(net831),
    .B(\mem.mem_internal.data_mem[27][2] ));
 sg13g2_nand2_1 _24444_ (.Y(_05864_),
    .A(net1250),
    .B(_05856_));
 sg13g2_o21ai_1 _24445_ (.B1(_05864_),
    .Y(_02318_),
    .A1(net419),
    .A2(_05863_));
 sg13g2_buf_1 _24446_ (.A(_05839_),
    .X(_05865_));
 sg13g2_nand2_1 _24447_ (.Y(_05866_),
    .A(net830),
    .B(\mem.mem_internal.data_mem[27][3] ));
 sg13g2_nand2_1 _24448_ (.Y(_05867_),
    .A(net1249),
    .B(_05856_));
 sg13g2_o21ai_1 _24449_ (.B1(_05867_),
    .Y(_02319_),
    .A1(net419),
    .A2(_05866_));
 sg13g2_nand2_1 _24450_ (.Y(_05868_),
    .A(net830),
    .B(\mem.mem_internal.data_mem[27][4] ));
 sg13g2_nand2_1 _24451_ (.Y(_05869_),
    .A(net1248),
    .B(_05856_));
 sg13g2_o21ai_1 _24452_ (.B1(_05869_),
    .Y(_02320_),
    .A1(_05857_),
    .A2(_05868_));
 sg13g2_nand2_1 _24453_ (.Y(_05870_),
    .A(net830),
    .B(\mem.mem_internal.data_mem[27][5] ));
 sg13g2_nand2_1 _24454_ (.Y(_05871_),
    .A(net1247),
    .B(_05856_));
 sg13g2_o21ai_1 _24455_ (.B1(_05871_),
    .Y(_02321_),
    .A1(net419),
    .A2(_05870_));
 sg13g2_nand2_1 _24456_ (.Y(_05872_),
    .A(net830),
    .B(\mem.mem_internal.data_mem[27][6] ));
 sg13g2_nand2_1 _24457_ (.Y(_05873_),
    .A(net1246),
    .B(_05856_));
 sg13g2_o21ai_1 _24458_ (.B1(_05873_),
    .Y(_02322_),
    .A1(net419),
    .A2(_05872_));
 sg13g2_nand2_1 _24459_ (.Y(_05874_),
    .A(net830),
    .B(\mem.mem_internal.data_mem[27][7] ));
 sg13g2_nand2_1 _24460_ (.Y(_05875_),
    .A(net1245),
    .B(_05856_));
 sg13g2_o21ai_1 _24461_ (.B1(_05875_),
    .Y(_02323_),
    .A1(_05857_),
    .A2(_05874_));
 sg13g2_nand3_1 _24462_ (.B(net1271),
    .C(_05519_),
    .A(net1269),
    .Y(_05876_));
 sg13g2_buf_1 _24463_ (.A(_05876_),
    .X(_05877_));
 sg13g2_nor2_1 _24464_ (.A(_05436_),
    .B(_05877_),
    .Y(_05878_));
 sg13g2_buf_2 _24465_ (.A(_05878_),
    .X(_05879_));
 sg13g2_buf_1 _24466_ (.A(_05879_),
    .X(_05880_));
 sg13g2_nand2_1 _24467_ (.Y(_05881_),
    .A(net830),
    .B(\mem.mem_internal.data_mem[28][0] ));
 sg13g2_buf_1 _24468_ (.A(net1292),
    .X(_05882_));
 sg13g2_nand2_1 _24469_ (.Y(_05883_),
    .A(net1243),
    .B(net418));
 sg13g2_o21ai_1 _24470_ (.B1(_05883_),
    .Y(_02324_),
    .A1(_05880_),
    .A2(_05881_));
 sg13g2_nand2_1 _24471_ (.Y(_05884_),
    .A(net830),
    .B(\mem.mem_internal.data_mem[28][1] ));
 sg13g2_nand2_1 _24472_ (.Y(_05885_),
    .A(net1244),
    .B(net418));
 sg13g2_o21ai_1 _24473_ (.B1(_05885_),
    .Y(_02325_),
    .A1(net418),
    .A2(_05884_));
 sg13g2_nand2_1 _24474_ (.Y(_05886_),
    .A(net830),
    .B(\mem.mem_internal.data_mem[28][2] ));
 sg13g2_buf_1 _24475_ (.A(net1290),
    .X(_05887_));
 sg13g2_nand2_1 _24476_ (.Y(_05888_),
    .A(net1242),
    .B(_05879_));
 sg13g2_o21ai_1 _24477_ (.B1(_05888_),
    .Y(_02326_),
    .A1(net418),
    .A2(_05886_));
 sg13g2_nand2_1 _24478_ (.Y(_05889_),
    .A(_05865_),
    .B(\mem.mem_internal.data_mem[28][3] ));
 sg13g2_buf_1 _24479_ (.A(net1289),
    .X(_05890_));
 sg13g2_nand2_1 _24480_ (.Y(_05891_),
    .A(net1241),
    .B(_05879_));
 sg13g2_o21ai_1 _24481_ (.B1(_05891_),
    .Y(_02327_),
    .A1(net418),
    .A2(_05889_));
 sg13g2_nand2_1 _24482_ (.Y(_05892_),
    .A(_05865_),
    .B(\mem.mem_internal.data_mem[28][4] ));
 sg13g2_buf_1 _24483_ (.A(net1288),
    .X(_05893_));
 sg13g2_nand2_1 _24484_ (.Y(_05894_),
    .A(net1240),
    .B(_05879_));
 sg13g2_o21ai_1 _24485_ (.B1(_05894_),
    .Y(_02328_),
    .A1(net418),
    .A2(_05892_));
 sg13g2_buf_1 _24486_ (.A(_05839_),
    .X(_05895_));
 sg13g2_nand2_1 _24487_ (.Y(_05896_),
    .A(net829),
    .B(\mem.mem_internal.data_mem[28][5] ));
 sg13g2_buf_1 _24488_ (.A(net1287),
    .X(_05897_));
 sg13g2_nand2_1 _24489_ (.Y(_05898_),
    .A(net1239),
    .B(_05879_));
 sg13g2_o21ai_1 _24490_ (.B1(_05898_),
    .Y(_02329_),
    .A1(net418),
    .A2(_05896_));
 sg13g2_nand2_1 _24491_ (.Y(_05899_),
    .A(net829),
    .B(\mem.mem_internal.data_mem[28][6] ));
 sg13g2_buf_1 _24492_ (.A(net1286),
    .X(_05900_));
 sg13g2_nand2_1 _24493_ (.Y(_05901_),
    .A(net1238),
    .B(_05879_));
 sg13g2_o21ai_1 _24494_ (.B1(_05901_),
    .Y(_02330_),
    .A1(net418),
    .A2(_05899_));
 sg13g2_nand2_1 _24495_ (.Y(_05902_),
    .A(net829),
    .B(\mem.mem_internal.data_mem[28][7] ));
 sg13g2_buf_1 _24496_ (.A(net1285),
    .X(_05903_));
 sg13g2_nand2_1 _24497_ (.Y(_05904_),
    .A(net1237),
    .B(_05879_));
 sg13g2_o21ai_1 _24498_ (.B1(_05904_),
    .Y(_02331_),
    .A1(_05880_),
    .A2(_05902_));
 sg13g2_nor2_1 _24499_ (.A(_05543_),
    .B(_05877_),
    .Y(_05905_));
 sg13g2_buf_2 _24500_ (.A(_05905_),
    .X(_05906_));
 sg13g2_buf_1 _24501_ (.A(_05906_),
    .X(_05907_));
 sg13g2_nand2_1 _24502_ (.Y(_05908_),
    .A(_05895_),
    .B(\mem.mem_internal.data_mem[29][0] ));
 sg13g2_nand2_1 _24503_ (.Y(_05909_),
    .A(net1243),
    .B(_05907_));
 sg13g2_o21ai_1 _24504_ (.B1(_05909_),
    .Y(_02332_),
    .A1(_05907_),
    .A2(_05908_));
 sg13g2_nand2_1 _24505_ (.Y(_05910_),
    .A(_05895_),
    .B(\mem.mem_internal.data_mem[29][1] ));
 sg13g2_nand2_1 _24506_ (.Y(_05911_),
    .A(net1244),
    .B(net417));
 sg13g2_o21ai_1 _24507_ (.B1(_05911_),
    .Y(_02333_),
    .A1(net417),
    .A2(_05910_));
 sg13g2_nand2_1 _24508_ (.Y(_05912_),
    .A(net829),
    .B(\mem.mem_internal.data_mem[29][2] ));
 sg13g2_nand2_1 _24509_ (.Y(_05913_),
    .A(net1242),
    .B(_05906_));
 sg13g2_o21ai_1 _24510_ (.B1(_05913_),
    .Y(_02334_),
    .A1(net417),
    .A2(_05912_));
 sg13g2_nand2_1 _24511_ (.Y(_05914_),
    .A(net829),
    .B(\mem.mem_internal.data_mem[29][3] ));
 sg13g2_nand2_1 _24512_ (.Y(_05915_),
    .A(net1241),
    .B(_05906_));
 sg13g2_o21ai_1 _24513_ (.B1(_05915_),
    .Y(_02335_),
    .A1(net417),
    .A2(_05914_));
 sg13g2_nand2_1 _24514_ (.Y(_05916_),
    .A(net829),
    .B(\mem.mem_internal.data_mem[29][4] ));
 sg13g2_nand2_1 _24515_ (.Y(_05917_),
    .A(net1240),
    .B(_05906_));
 sg13g2_o21ai_1 _24516_ (.B1(_05917_),
    .Y(_02336_),
    .A1(net417),
    .A2(_05916_));
 sg13g2_nand2_1 _24517_ (.Y(_05918_),
    .A(net829),
    .B(\mem.mem_internal.data_mem[29][5] ));
 sg13g2_nand2_1 _24518_ (.Y(_05919_),
    .A(net1239),
    .B(_05906_));
 sg13g2_o21ai_1 _24519_ (.B1(_05919_),
    .Y(_02337_),
    .A1(net417),
    .A2(_05918_));
 sg13g2_nand2_1 _24520_ (.Y(_05920_),
    .A(net829),
    .B(\mem.mem_internal.data_mem[29][6] ));
 sg13g2_nand2_1 _24521_ (.Y(_05921_),
    .A(net1238),
    .B(_05906_));
 sg13g2_o21ai_1 _24522_ (.B1(_05921_),
    .Y(_02338_),
    .A1(net417),
    .A2(_05920_));
 sg13g2_buf_1 _24523_ (.A(_05839_),
    .X(_05922_));
 sg13g2_nand2_1 _24524_ (.Y(_05923_),
    .A(net828),
    .B(\mem.mem_internal.data_mem[29][7] ));
 sg13g2_nand2_1 _24525_ (.Y(_05924_),
    .A(net1237),
    .B(_05906_));
 sg13g2_o21ai_1 _24526_ (.B1(_05924_),
    .Y(_02339_),
    .A1(net417),
    .A2(_05923_));
 sg13g2_nor2_1 _24527_ (.A(_05429_),
    .B(_05477_),
    .Y(_05925_));
 sg13g2_buf_2 _24528_ (.A(_05925_),
    .X(_05926_));
 sg13g2_buf_1 _24529_ (.A(_05926_),
    .X(_05927_));
 sg13g2_nand2_1 _24530_ (.Y(_05928_),
    .A(net828),
    .B(\mem.mem_internal.data_mem[2][0] ));
 sg13g2_nand2_1 _24531_ (.Y(_05929_),
    .A(_05882_),
    .B(net416));
 sg13g2_o21ai_1 _24532_ (.B1(_05929_),
    .Y(_02340_),
    .A1(net416),
    .A2(_05928_));
 sg13g2_nand2_1 _24533_ (.Y(_05930_),
    .A(net828),
    .B(\mem.mem_internal.data_mem[2][1] ));
 sg13g2_nand2_1 _24534_ (.Y(_05931_),
    .A(_05861_),
    .B(net416));
 sg13g2_o21ai_1 _24535_ (.B1(_05931_),
    .Y(_02341_),
    .A1(net416),
    .A2(_05930_));
 sg13g2_nand2_1 _24536_ (.Y(_05932_),
    .A(net828),
    .B(\mem.mem_internal.data_mem[2][2] ));
 sg13g2_nand2_1 _24537_ (.Y(_05933_),
    .A(_05887_),
    .B(_05926_));
 sg13g2_o21ai_1 _24538_ (.B1(_05933_),
    .Y(_02342_),
    .A1(net416),
    .A2(_05932_));
 sg13g2_nand2_1 _24539_ (.Y(_05934_),
    .A(net828),
    .B(\mem.mem_internal.data_mem[2][3] ));
 sg13g2_nand2_1 _24540_ (.Y(_05935_),
    .A(net1241),
    .B(_05926_));
 sg13g2_o21ai_1 _24541_ (.B1(_05935_),
    .Y(_02343_),
    .A1(_05927_),
    .A2(_05934_));
 sg13g2_nand2_1 _24542_ (.Y(_05936_),
    .A(net828),
    .B(\mem.mem_internal.data_mem[2][4] ));
 sg13g2_nand2_1 _24543_ (.Y(_05937_),
    .A(net1240),
    .B(_05926_));
 sg13g2_o21ai_1 _24544_ (.B1(_05937_),
    .Y(_02344_),
    .A1(_05927_),
    .A2(_05936_));
 sg13g2_nand2_1 _24545_ (.Y(_05938_),
    .A(net828),
    .B(\mem.mem_internal.data_mem[2][5] ));
 sg13g2_nand2_1 _24546_ (.Y(_05939_),
    .A(net1239),
    .B(_05926_));
 sg13g2_o21ai_1 _24547_ (.B1(_05939_),
    .Y(_02345_),
    .A1(net416),
    .A2(_05938_));
 sg13g2_nand2_1 _24548_ (.Y(_05940_),
    .A(_05922_),
    .B(\mem.mem_internal.data_mem[2][6] ));
 sg13g2_nand2_1 _24549_ (.Y(_05941_),
    .A(net1238),
    .B(_05926_));
 sg13g2_o21ai_1 _24550_ (.B1(_05941_),
    .Y(_02346_),
    .A1(net416),
    .A2(_05940_));
 sg13g2_nand2_1 _24551_ (.Y(_05942_),
    .A(_05922_),
    .B(\mem.mem_internal.data_mem[2][7] ));
 sg13g2_nand2_1 _24552_ (.Y(_05943_),
    .A(_05903_),
    .B(_05926_));
 sg13g2_o21ai_1 _24553_ (.B1(_05943_),
    .Y(_02347_),
    .A1(net416),
    .A2(_05942_));
 sg13g2_nor2_1 _24554_ (.A(_05477_),
    .B(_05877_),
    .Y(_05944_));
 sg13g2_buf_2 _24555_ (.A(_05944_),
    .X(_05945_));
 sg13g2_buf_1 _24556_ (.A(_05945_),
    .X(_05946_));
 sg13g2_nand2_1 _24557_ (.Y(_05947_),
    .A(net828),
    .B(\mem.mem_internal.data_mem[30][0] ));
 sg13g2_nand2_1 _24558_ (.Y(_05948_),
    .A(net1243),
    .B(net415));
 sg13g2_o21ai_1 _24559_ (.B1(_05948_),
    .Y(_02348_),
    .A1(_05946_),
    .A2(_05947_));
 sg13g2_buf_1 _24560_ (.A(_05839_),
    .X(_05949_));
 sg13g2_nand2_1 _24561_ (.Y(_05950_),
    .A(_05949_),
    .B(\mem.mem_internal.data_mem[30][1] ));
 sg13g2_nand2_1 _24562_ (.Y(_05951_),
    .A(net1244),
    .B(net415));
 sg13g2_o21ai_1 _24563_ (.B1(_05951_),
    .Y(_02349_),
    .A1(_05946_),
    .A2(_05950_));
 sg13g2_nand2_1 _24564_ (.Y(_05952_),
    .A(net827),
    .B(\mem.mem_internal.data_mem[30][2] ));
 sg13g2_nand2_1 _24565_ (.Y(_05953_),
    .A(net1242),
    .B(_05945_));
 sg13g2_o21ai_1 _24566_ (.B1(_05953_),
    .Y(_02350_),
    .A1(net415),
    .A2(_05952_));
 sg13g2_nand2_1 _24567_ (.Y(_05954_),
    .A(net827),
    .B(\mem.mem_internal.data_mem[30][3] ));
 sg13g2_nand2_1 _24568_ (.Y(_05955_),
    .A(net1241),
    .B(_05945_));
 sg13g2_o21ai_1 _24569_ (.B1(_05955_),
    .Y(_02351_),
    .A1(net415),
    .A2(_05954_));
 sg13g2_nand2_1 _24570_ (.Y(_05956_),
    .A(net827),
    .B(\mem.mem_internal.data_mem[30][4] ));
 sg13g2_nand2_1 _24571_ (.Y(_05957_),
    .A(net1240),
    .B(_05945_));
 sg13g2_o21ai_1 _24572_ (.B1(_05957_),
    .Y(_02352_),
    .A1(net415),
    .A2(_05956_));
 sg13g2_nand2_1 _24573_ (.Y(_05958_),
    .A(net827),
    .B(\mem.mem_internal.data_mem[30][5] ));
 sg13g2_nand2_1 _24574_ (.Y(_05959_),
    .A(net1239),
    .B(_05945_));
 sg13g2_o21ai_1 _24575_ (.B1(_05959_),
    .Y(_02353_),
    .A1(net415),
    .A2(_05958_));
 sg13g2_nand2_1 _24576_ (.Y(_05960_),
    .A(net827),
    .B(\mem.mem_internal.data_mem[30][6] ));
 sg13g2_nand2_1 _24577_ (.Y(_05961_),
    .A(net1238),
    .B(_05945_));
 sg13g2_o21ai_1 _24578_ (.B1(_05961_),
    .Y(_02354_),
    .A1(net415),
    .A2(_05960_));
 sg13g2_nand2_1 _24579_ (.Y(_05962_),
    .A(net827),
    .B(\mem.mem_internal.data_mem[30][7] ));
 sg13g2_nand2_1 _24580_ (.Y(_05963_),
    .A(net1237),
    .B(_05945_));
 sg13g2_o21ai_1 _24581_ (.B1(_05963_),
    .Y(_02355_),
    .A1(net415),
    .A2(_05962_));
 sg13g2_nor2_1 _24582_ (.A(_05499_),
    .B(_05877_),
    .Y(_05964_));
 sg13g2_buf_2 _24583_ (.A(_05964_),
    .X(_05965_));
 sg13g2_buf_1 _24584_ (.A(_05965_),
    .X(_05966_));
 sg13g2_nand2_1 _24585_ (.Y(_05967_),
    .A(net827),
    .B(\mem.mem_internal.data_mem[31][0] ));
 sg13g2_nand2_1 _24586_ (.Y(_05968_),
    .A(net1243),
    .B(_05966_));
 sg13g2_o21ai_1 _24587_ (.B1(_05968_),
    .Y(_02356_),
    .A1(_05966_),
    .A2(_05967_));
 sg13g2_nand2_1 _24588_ (.Y(_05969_),
    .A(_05949_),
    .B(\mem.mem_internal.data_mem[31][1] ));
 sg13g2_nand2_1 _24589_ (.Y(_05970_),
    .A(net1244),
    .B(net414));
 sg13g2_o21ai_1 _24590_ (.B1(_05970_),
    .Y(_02357_),
    .A1(net414),
    .A2(_05969_));
 sg13g2_nand2_1 _24591_ (.Y(_05971_),
    .A(net827),
    .B(\mem.mem_internal.data_mem[31][2] ));
 sg13g2_nand2_1 _24592_ (.Y(_05972_),
    .A(net1242),
    .B(_05965_));
 sg13g2_o21ai_1 _24593_ (.B1(_05972_),
    .Y(_02358_),
    .A1(net414),
    .A2(_05971_));
 sg13g2_buf_1 _24594_ (.A(_05839_),
    .X(_05973_));
 sg13g2_nand2_1 _24595_ (.Y(_05974_),
    .A(net826),
    .B(\mem.mem_internal.data_mem[31][3] ));
 sg13g2_nand2_1 _24596_ (.Y(_05975_),
    .A(net1241),
    .B(_05965_));
 sg13g2_o21ai_1 _24597_ (.B1(_05975_),
    .Y(_02359_),
    .A1(net414),
    .A2(_05974_));
 sg13g2_nand2_1 _24598_ (.Y(_05976_),
    .A(net826),
    .B(\mem.mem_internal.data_mem[31][4] ));
 sg13g2_nand2_1 _24599_ (.Y(_05977_),
    .A(net1240),
    .B(_05965_));
 sg13g2_o21ai_1 _24600_ (.B1(_05977_),
    .Y(_02360_),
    .A1(net414),
    .A2(_05976_));
 sg13g2_nand2_1 _24601_ (.Y(_05978_),
    .A(net826),
    .B(\mem.mem_internal.data_mem[31][5] ));
 sg13g2_nand2_1 _24602_ (.Y(_05979_),
    .A(net1239),
    .B(_05965_));
 sg13g2_o21ai_1 _24603_ (.B1(_05979_),
    .Y(_02361_),
    .A1(net414),
    .A2(_05978_));
 sg13g2_nand2_1 _24604_ (.Y(_05980_),
    .A(net826),
    .B(\mem.mem_internal.data_mem[31][6] ));
 sg13g2_nand2_1 _24605_ (.Y(_05981_),
    .A(net1238),
    .B(_05965_));
 sg13g2_o21ai_1 _24606_ (.B1(_05981_),
    .Y(_02362_),
    .A1(net414),
    .A2(_05980_));
 sg13g2_nand2_1 _24607_ (.Y(_05982_),
    .A(net826),
    .B(\mem.mem_internal.data_mem[31][7] ));
 sg13g2_nand2_1 _24608_ (.Y(_05983_),
    .A(net1237),
    .B(_05965_));
 sg13g2_o21ai_1 _24609_ (.B1(_05983_),
    .Y(_02363_),
    .A1(net414),
    .A2(_05982_));
 sg13g2_nor2_1 _24610_ (.A(_05429_),
    .B(_05499_),
    .Y(_05984_));
 sg13g2_buf_1 _24611_ (.A(_05984_),
    .X(_05985_));
 sg13g2_buf_1 _24612_ (.A(_05985_),
    .X(_05986_));
 sg13g2_nand2_1 _24613_ (.Y(_05987_),
    .A(net826),
    .B(\mem.mem_internal.data_mem[3][0] ));
 sg13g2_nand2_1 _24614_ (.Y(_05988_),
    .A(_05882_),
    .B(net413));
 sg13g2_o21ai_1 _24615_ (.B1(_05988_),
    .Y(_02364_),
    .A1(net413),
    .A2(_05987_));
 sg13g2_nand2_1 _24616_ (.Y(_05989_),
    .A(net826),
    .B(\mem.mem_internal.data_mem[3][1] ));
 sg13g2_nand2_1 _24617_ (.Y(_05990_),
    .A(_05861_),
    .B(net413));
 sg13g2_o21ai_1 _24618_ (.B1(_05990_),
    .Y(_02365_),
    .A1(net413),
    .A2(_05989_));
 sg13g2_nand2_1 _24619_ (.Y(_05991_),
    .A(net826),
    .B(\mem.mem_internal.data_mem[3][2] ));
 sg13g2_nand2_1 _24620_ (.Y(_05992_),
    .A(_05887_),
    .B(_05985_));
 sg13g2_o21ai_1 _24621_ (.B1(_05992_),
    .Y(_02366_),
    .A1(net413),
    .A2(_05991_));
 sg13g2_nand2_1 _24622_ (.Y(_05993_),
    .A(_05973_),
    .B(\mem.mem_internal.data_mem[3][3] ));
 sg13g2_nand2_1 _24623_ (.Y(_05994_),
    .A(net1241),
    .B(_05985_));
 sg13g2_o21ai_1 _24624_ (.B1(_05994_),
    .Y(_02367_),
    .A1(_05986_),
    .A2(_05993_));
 sg13g2_nand2_1 _24625_ (.Y(_05995_),
    .A(_05973_),
    .B(\mem.mem_internal.data_mem[3][4] ));
 sg13g2_nand2_1 _24626_ (.Y(_05996_),
    .A(net1240),
    .B(_05985_));
 sg13g2_o21ai_1 _24627_ (.B1(_05996_),
    .Y(_02368_),
    .A1(_05986_),
    .A2(_05995_));
 sg13g2_buf_1 _24628_ (.A(_05839_),
    .X(_05997_));
 sg13g2_nand2_1 _24629_ (.Y(_05998_),
    .A(_05997_),
    .B(\mem.mem_internal.data_mem[3][5] ));
 sg13g2_nand2_1 _24630_ (.Y(_05999_),
    .A(net1239),
    .B(_05985_));
 sg13g2_o21ai_1 _24631_ (.B1(_05999_),
    .Y(_02369_),
    .A1(net413),
    .A2(_05998_));
 sg13g2_nand2_1 _24632_ (.Y(_06000_),
    .A(net825),
    .B(\mem.mem_internal.data_mem[3][6] ));
 sg13g2_nand2_1 _24633_ (.Y(_06001_),
    .A(net1238),
    .B(_05985_));
 sg13g2_o21ai_1 _24634_ (.B1(_06001_),
    .Y(_02370_),
    .A1(net413),
    .A2(_06000_));
 sg13g2_nand2_1 _24635_ (.Y(_06002_),
    .A(_05997_),
    .B(\mem.mem_internal.data_mem[3][7] ));
 sg13g2_nand2_1 _24636_ (.Y(_06003_),
    .A(_05903_),
    .B(_05985_));
 sg13g2_o21ai_1 _24637_ (.B1(_06003_),
    .Y(_02371_),
    .A1(net413),
    .A2(_06002_));
 sg13g2_nand2_1 _24638_ (.Y(_06004_),
    .A(_10114_),
    .B(_05713_));
 sg13g2_nor2_1 _24639_ (.A(_05436_),
    .B(_06004_),
    .Y(_06005_));
 sg13g2_buf_2 _24640_ (.A(_06005_),
    .X(_06006_));
 sg13g2_buf_1 _24641_ (.A(_06006_),
    .X(_06007_));
 sg13g2_nand2_1 _24642_ (.Y(_06008_),
    .A(net825),
    .B(\mem.mem_internal.data_mem[4][0] ));
 sg13g2_nand2_1 _24643_ (.Y(_06009_),
    .A(net1243),
    .B(net412));
 sg13g2_o21ai_1 _24644_ (.B1(_06009_),
    .Y(_02372_),
    .A1(net412),
    .A2(_06008_));
 sg13g2_nand2_1 _24645_ (.Y(_06010_),
    .A(net825),
    .B(\mem.mem_internal.data_mem[4][1] ));
 sg13g2_nand2_1 _24646_ (.Y(_06011_),
    .A(net1244),
    .B(net412));
 sg13g2_o21ai_1 _24647_ (.B1(_06011_),
    .Y(_02373_),
    .A1(net412),
    .A2(_06010_));
 sg13g2_nand2_1 _24648_ (.Y(_06012_),
    .A(net825),
    .B(\mem.mem_internal.data_mem[4][2] ));
 sg13g2_nand2_1 _24649_ (.Y(_06013_),
    .A(net1242),
    .B(_06006_));
 sg13g2_o21ai_1 _24650_ (.B1(_06013_),
    .Y(_02374_),
    .A1(net412),
    .A2(_06012_));
 sg13g2_nand2_1 _24651_ (.Y(_06014_),
    .A(net825),
    .B(\mem.mem_internal.data_mem[4][3] ));
 sg13g2_nand2_1 _24652_ (.Y(_06015_),
    .A(net1241),
    .B(_06006_));
 sg13g2_o21ai_1 _24653_ (.B1(_06015_),
    .Y(_02375_),
    .A1(net412),
    .A2(_06014_));
 sg13g2_nand2_1 _24654_ (.Y(_06016_),
    .A(net825),
    .B(\mem.mem_internal.data_mem[4][4] ));
 sg13g2_nand2_1 _24655_ (.Y(_06017_),
    .A(net1240),
    .B(_06006_));
 sg13g2_o21ai_1 _24656_ (.B1(_06017_),
    .Y(_02376_),
    .A1(net412),
    .A2(_06016_));
 sg13g2_nand2_1 _24657_ (.Y(_06018_),
    .A(net825),
    .B(\mem.mem_internal.data_mem[4][5] ));
 sg13g2_nand2_1 _24658_ (.Y(_06019_),
    .A(net1239),
    .B(_06006_));
 sg13g2_o21ai_1 _24659_ (.B1(_06019_),
    .Y(_02377_),
    .A1(_06007_),
    .A2(_06018_));
 sg13g2_nand2_1 _24660_ (.Y(_06020_),
    .A(net825),
    .B(\mem.mem_internal.data_mem[4][6] ));
 sg13g2_nand2_1 _24661_ (.Y(_06021_),
    .A(net1238),
    .B(_06006_));
 sg13g2_o21ai_1 _24662_ (.B1(_06021_),
    .Y(_02378_),
    .A1(_06007_),
    .A2(_06020_));
 sg13g2_buf_1 _24663_ (.A(_10070_),
    .X(_06022_));
 sg13g2_nand2_1 _24664_ (.Y(_06023_),
    .A(net824),
    .B(\mem.mem_internal.data_mem[4][7] ));
 sg13g2_nand2_1 _24665_ (.Y(_06024_),
    .A(net1237),
    .B(_06006_));
 sg13g2_o21ai_1 _24666_ (.B1(_06024_),
    .Y(_02379_),
    .A1(net412),
    .A2(_06023_));
 sg13g2_nor2_1 _24667_ (.A(_05543_),
    .B(_06004_),
    .Y(_06025_));
 sg13g2_buf_2 _24668_ (.A(_06025_),
    .X(_06026_));
 sg13g2_buf_1 _24669_ (.A(_06026_),
    .X(_06027_));
 sg13g2_nand2_1 _24670_ (.Y(_06028_),
    .A(net824),
    .B(\mem.mem_internal.data_mem[5][0] ));
 sg13g2_nand2_1 _24671_ (.Y(_06029_),
    .A(net1243),
    .B(net411));
 sg13g2_o21ai_1 _24672_ (.B1(_06029_),
    .Y(_02380_),
    .A1(net411),
    .A2(_06028_));
 sg13g2_nand2_1 _24673_ (.Y(_06030_),
    .A(net824),
    .B(\mem.mem_internal.data_mem[5][1] ));
 sg13g2_nand2_1 _24674_ (.Y(_06031_),
    .A(net1244),
    .B(net411));
 sg13g2_o21ai_1 _24675_ (.B1(_06031_),
    .Y(_02381_),
    .A1(net411),
    .A2(_06030_));
 sg13g2_nand2_1 _24676_ (.Y(_06032_),
    .A(net824),
    .B(\mem.mem_internal.data_mem[5][2] ));
 sg13g2_nand2_1 _24677_ (.Y(_06033_),
    .A(net1242),
    .B(_06026_));
 sg13g2_o21ai_1 _24678_ (.B1(_06033_),
    .Y(_02382_),
    .A1(net411),
    .A2(_06032_));
 sg13g2_nand2_1 _24679_ (.Y(_06034_),
    .A(net824),
    .B(\mem.mem_internal.data_mem[5][3] ));
 sg13g2_nand2_1 _24680_ (.Y(_06035_),
    .A(net1241),
    .B(_06026_));
 sg13g2_o21ai_1 _24681_ (.B1(_06035_),
    .Y(_02383_),
    .A1(net411),
    .A2(_06034_));
 sg13g2_nand2_1 _24682_ (.Y(_06036_),
    .A(net824),
    .B(\mem.mem_internal.data_mem[5][4] ));
 sg13g2_nand2_1 _24683_ (.Y(_06037_),
    .A(_05893_),
    .B(_06026_));
 sg13g2_o21ai_1 _24684_ (.B1(_06037_),
    .Y(_02384_),
    .A1(net411),
    .A2(_06036_));
 sg13g2_nand2_1 _24685_ (.Y(_06038_),
    .A(net824),
    .B(\mem.mem_internal.data_mem[5][5] ));
 sg13g2_nand2_1 _24686_ (.Y(_06039_),
    .A(_05897_),
    .B(_06026_));
 sg13g2_o21ai_1 _24687_ (.B1(_06039_),
    .Y(_02385_),
    .A1(net411),
    .A2(_06038_));
 sg13g2_nand2_1 _24688_ (.Y(_06040_),
    .A(_06022_),
    .B(\mem.mem_internal.data_mem[5][6] ));
 sg13g2_nand2_1 _24689_ (.Y(_06041_),
    .A(net1238),
    .B(_06026_));
 sg13g2_o21ai_1 _24690_ (.B1(_06041_),
    .Y(_02386_),
    .A1(_06027_),
    .A2(_06040_));
 sg13g2_nand2_1 _24691_ (.Y(_06042_),
    .A(_06022_),
    .B(\mem.mem_internal.data_mem[5][7] ));
 sg13g2_nand2_1 _24692_ (.Y(_06043_),
    .A(net1237),
    .B(_06026_));
 sg13g2_o21ai_1 _24693_ (.B1(_06043_),
    .Y(_02387_),
    .A1(_06027_),
    .A2(_06042_));
 sg13g2_nor2_1 _24694_ (.A(_05477_),
    .B(_06004_),
    .Y(_06044_));
 sg13g2_buf_2 _24695_ (.A(_06044_),
    .X(_06045_));
 sg13g2_buf_1 _24696_ (.A(_06045_),
    .X(_06046_));
 sg13g2_nand2_1 _24697_ (.Y(_06047_),
    .A(net824),
    .B(\mem.mem_internal.data_mem[6][0] ));
 sg13g2_nand2_1 _24698_ (.Y(_06048_),
    .A(net1243),
    .B(net410));
 sg13g2_o21ai_1 _24699_ (.B1(_06048_),
    .Y(_02388_),
    .A1(net410),
    .A2(_06047_));
 sg13g2_buf_1 _24700_ (.A(_10070_),
    .X(_06049_));
 sg13g2_nand2_1 _24701_ (.Y(_06050_),
    .A(net823),
    .B(\mem.mem_internal.data_mem[6][1] ));
 sg13g2_nand2_1 _24702_ (.Y(_06051_),
    .A(net1244),
    .B(net410));
 sg13g2_o21ai_1 _24703_ (.B1(_06051_),
    .Y(_02389_),
    .A1(_06046_),
    .A2(_06050_));
 sg13g2_nand2_1 _24704_ (.Y(_06052_),
    .A(net823),
    .B(\mem.mem_internal.data_mem[6][2] ));
 sg13g2_nand2_1 _24705_ (.Y(_06053_),
    .A(net1242),
    .B(_06045_));
 sg13g2_o21ai_1 _24706_ (.B1(_06053_),
    .Y(_02390_),
    .A1(net410),
    .A2(_06052_));
 sg13g2_nand2_1 _24707_ (.Y(_06054_),
    .A(net823),
    .B(\mem.mem_internal.data_mem[6][3] ));
 sg13g2_nand2_1 _24708_ (.Y(_06055_),
    .A(_05890_),
    .B(_06045_));
 sg13g2_o21ai_1 _24709_ (.B1(_06055_),
    .Y(_02391_),
    .A1(net410),
    .A2(_06054_));
 sg13g2_nand2_1 _24710_ (.Y(_06056_),
    .A(net823),
    .B(\mem.mem_internal.data_mem[6][4] ));
 sg13g2_nand2_1 _24711_ (.Y(_06057_),
    .A(_05893_),
    .B(_06045_));
 sg13g2_o21ai_1 _24712_ (.B1(_06057_),
    .Y(_02392_),
    .A1(net410),
    .A2(_06056_));
 sg13g2_nand2_1 _24713_ (.Y(_06058_),
    .A(_06049_),
    .B(\mem.mem_internal.data_mem[6][5] ));
 sg13g2_nand2_1 _24714_ (.Y(_06059_),
    .A(_05897_),
    .B(_06045_));
 sg13g2_o21ai_1 _24715_ (.B1(_06059_),
    .Y(_02393_),
    .A1(net410),
    .A2(_06058_));
 sg13g2_nand2_1 _24716_ (.Y(_06060_),
    .A(_06049_),
    .B(\mem.mem_internal.data_mem[6][6] ));
 sg13g2_nand2_1 _24717_ (.Y(_06061_),
    .A(_05900_),
    .B(_06045_));
 sg13g2_o21ai_1 _24718_ (.B1(_06061_),
    .Y(_02394_),
    .A1(_06046_),
    .A2(_06060_));
 sg13g2_nand2_1 _24719_ (.Y(_06062_),
    .A(net823),
    .B(\mem.mem_internal.data_mem[6][7] ));
 sg13g2_nand2_1 _24720_ (.Y(_06063_),
    .A(net1237),
    .B(_06045_));
 sg13g2_o21ai_1 _24721_ (.B1(_06063_),
    .Y(_02395_),
    .A1(net410),
    .A2(_06062_));
 sg13g2_nor2_1 _24722_ (.A(_05499_),
    .B(_06004_),
    .Y(_06064_));
 sg13g2_buf_2 _24723_ (.A(_06064_),
    .X(_06065_));
 sg13g2_buf_1 _24724_ (.A(_06065_),
    .X(_06066_));
 sg13g2_nand2_1 _24725_ (.Y(_06067_),
    .A(net823),
    .B(\mem.mem_internal.data_mem[7][0] ));
 sg13g2_nand2_1 _24726_ (.Y(_06068_),
    .A(net1243),
    .B(net409));
 sg13g2_o21ai_1 _24727_ (.B1(_06068_),
    .Y(_02396_),
    .A1(net409),
    .A2(_06067_));
 sg13g2_nand2_1 _24728_ (.Y(_06069_),
    .A(net823),
    .B(\mem.mem_internal.data_mem[7][1] ));
 sg13g2_nand2_1 _24729_ (.Y(_06070_),
    .A(net1291),
    .B(net409));
 sg13g2_o21ai_1 _24730_ (.B1(_06070_),
    .Y(_02397_),
    .A1(net409),
    .A2(_06069_));
 sg13g2_nand2_1 _24731_ (.Y(_06071_),
    .A(net823),
    .B(\mem.mem_internal.data_mem[7][2] ));
 sg13g2_nand2_1 _24732_ (.Y(_06072_),
    .A(net1242),
    .B(_06065_));
 sg13g2_o21ai_1 _24733_ (.B1(_06072_),
    .Y(_02398_),
    .A1(net409),
    .A2(_06071_));
 sg13g2_buf_1 _24734_ (.A(_10070_),
    .X(_06073_));
 sg13g2_nand2_1 _24735_ (.Y(_06074_),
    .A(net822),
    .B(\mem.mem_internal.data_mem[7][3] ));
 sg13g2_nand2_1 _24736_ (.Y(_06075_),
    .A(_05890_),
    .B(_06065_));
 sg13g2_o21ai_1 _24737_ (.B1(_06075_),
    .Y(_02399_),
    .A1(_06066_),
    .A2(_06074_));
 sg13g2_nand2_1 _24738_ (.Y(_06076_),
    .A(net822),
    .B(\mem.mem_internal.data_mem[7][4] ));
 sg13g2_nand2_1 _24739_ (.Y(_06077_),
    .A(net1240),
    .B(_06065_));
 sg13g2_o21ai_1 _24740_ (.B1(_06077_),
    .Y(_02400_),
    .A1(net409),
    .A2(_06076_));
 sg13g2_nand2_1 _24741_ (.Y(_06078_),
    .A(net822),
    .B(\mem.mem_internal.data_mem[7][5] ));
 sg13g2_nand2_1 _24742_ (.Y(_06079_),
    .A(net1239),
    .B(_06065_));
 sg13g2_o21ai_1 _24743_ (.B1(_06079_),
    .Y(_02401_),
    .A1(net409),
    .A2(_06078_));
 sg13g2_nand2_1 _24744_ (.Y(_06080_),
    .A(net822),
    .B(\mem.mem_internal.data_mem[7][6] ));
 sg13g2_nand2_1 _24745_ (.Y(_06081_),
    .A(_05900_),
    .B(_06065_));
 sg13g2_o21ai_1 _24746_ (.B1(_06081_),
    .Y(_02402_),
    .A1(_06066_),
    .A2(_06080_));
 sg13g2_nand2_1 _24747_ (.Y(_06082_),
    .A(net822),
    .B(\mem.mem_internal.data_mem[7][7] ));
 sg13g2_nand2_1 _24748_ (.Y(_06083_),
    .A(net1237),
    .B(_06065_));
 sg13g2_o21ai_1 _24749_ (.B1(_06083_),
    .Y(_02403_),
    .A1(net409),
    .A2(_06082_));
 sg13g2_nor3_1 _24750_ (.A(net1269),
    .B(_05475_),
    .C(_05436_),
    .Y(_06084_));
 sg13g2_buf_2 _24751_ (.A(_06084_),
    .X(_06085_));
 sg13g2_buf_1 _24752_ (.A(_06085_),
    .X(_06086_));
 sg13g2_nand2_1 _24753_ (.Y(_06087_),
    .A(net822),
    .B(\mem.mem_internal.data_mem[8][0] ));
 sg13g2_nand2_1 _24754_ (.Y(_06088_),
    .A(net1292),
    .B(net408));
 sg13g2_o21ai_1 _24755_ (.B1(_06088_),
    .Y(_02404_),
    .A1(net408),
    .A2(_06087_));
 sg13g2_nand2_1 _24756_ (.Y(_06089_),
    .A(net822),
    .B(\mem.mem_internal.data_mem[8][1] ));
 sg13g2_nand2_1 _24757_ (.Y(_06090_),
    .A(net1291),
    .B(net408));
 sg13g2_o21ai_1 _24758_ (.B1(_06090_),
    .Y(_02405_),
    .A1(_06086_),
    .A2(_06089_));
 sg13g2_nand2_1 _24759_ (.Y(_06091_),
    .A(net822),
    .B(\mem.mem_internal.data_mem[8][2] ));
 sg13g2_nand2_1 _24760_ (.Y(_06092_),
    .A(net1290),
    .B(_06085_));
 sg13g2_o21ai_1 _24761_ (.B1(_06092_),
    .Y(_02406_),
    .A1(net408),
    .A2(_06091_));
 sg13g2_nand2_1 _24762_ (.Y(_06093_),
    .A(_06073_),
    .B(\mem.mem_internal.data_mem[8][3] ));
 sg13g2_nand2_1 _24763_ (.Y(_06094_),
    .A(net1289),
    .B(_06085_));
 sg13g2_o21ai_1 _24764_ (.B1(_06094_),
    .Y(_02407_),
    .A1(net408),
    .A2(_06093_));
 sg13g2_nand2_1 _24765_ (.Y(_06095_),
    .A(_06073_),
    .B(\mem.mem_internal.data_mem[8][4] ));
 sg13g2_nand2_1 _24766_ (.Y(_06096_),
    .A(net1288),
    .B(_06085_));
 sg13g2_o21ai_1 _24767_ (.B1(_06096_),
    .Y(_02408_),
    .A1(net408),
    .A2(_06095_));
 sg13g2_buf_1 _24768_ (.A(_10070_),
    .X(_06097_));
 sg13g2_nand2_1 _24769_ (.Y(_06098_),
    .A(_06097_),
    .B(\mem.mem_internal.data_mem[8][5] ));
 sg13g2_nand2_1 _24770_ (.Y(_06099_),
    .A(net1287),
    .B(_06085_));
 sg13g2_o21ai_1 _24771_ (.B1(_06099_),
    .Y(_02409_),
    .A1(_06086_),
    .A2(_06098_));
 sg13g2_nand2_1 _24772_ (.Y(_06100_),
    .A(net821),
    .B(\mem.mem_internal.data_mem[8][6] ));
 sg13g2_nand2_1 _24773_ (.Y(_06101_),
    .A(net1286),
    .B(_06085_));
 sg13g2_o21ai_1 _24774_ (.B1(_06101_),
    .Y(_02410_),
    .A1(net408),
    .A2(_06100_));
 sg13g2_nand2_1 _24775_ (.Y(_06102_),
    .A(net821),
    .B(\mem.mem_internal.data_mem[8][7] ));
 sg13g2_nand2_1 _24776_ (.Y(_06103_),
    .A(net1285),
    .B(_06085_));
 sg13g2_o21ai_1 _24777_ (.B1(_06103_),
    .Y(_02411_),
    .A1(net408),
    .A2(_06102_));
 sg13g2_nor3_1 _24778_ (.A(net1269),
    .B(_05475_),
    .C(_05543_),
    .Y(_06104_));
 sg13g2_buf_2 _24779_ (.A(_06104_),
    .X(_06105_));
 sg13g2_buf_1 _24780_ (.A(_06105_),
    .X(_06106_));
 sg13g2_nand2_1 _24781_ (.Y(_06107_),
    .A(net821),
    .B(\mem.mem_internal.data_mem[9][0] ));
 sg13g2_nand2_1 _24782_ (.Y(_06108_),
    .A(net1292),
    .B(net407));
 sg13g2_o21ai_1 _24783_ (.B1(_06108_),
    .Y(_02412_),
    .A1(net407),
    .A2(_06107_));
 sg13g2_nand2_1 _24784_ (.Y(_06109_),
    .A(net821),
    .B(\mem.mem_internal.data_mem[9][1] ));
 sg13g2_nand2_1 _24785_ (.Y(_06110_),
    .A(net1291),
    .B(net407));
 sg13g2_o21ai_1 _24786_ (.B1(_06110_),
    .Y(_02413_),
    .A1(net407),
    .A2(_06109_));
 sg13g2_nand2_1 _24787_ (.Y(_06111_),
    .A(net821),
    .B(\mem.mem_internal.data_mem[9][2] ));
 sg13g2_nand2_1 _24788_ (.Y(_06112_),
    .A(net1290),
    .B(_06105_));
 sg13g2_o21ai_1 _24789_ (.B1(_06112_),
    .Y(_02414_),
    .A1(net407),
    .A2(_06111_));
 sg13g2_nand2_1 _24790_ (.Y(_06113_),
    .A(net821),
    .B(\mem.mem_internal.data_mem[9][3] ));
 sg13g2_nand2_1 _24791_ (.Y(_06114_),
    .A(net1289),
    .B(_06105_));
 sg13g2_o21ai_1 _24792_ (.B1(_06114_),
    .Y(_02415_),
    .A1(net407),
    .A2(_06113_));
 sg13g2_nand2_1 _24793_ (.Y(_06115_),
    .A(net821),
    .B(\mem.mem_internal.data_mem[9][4] ));
 sg13g2_nand2_1 _24794_ (.Y(_06116_),
    .A(net1288),
    .B(_06105_));
 sg13g2_o21ai_1 _24795_ (.B1(_06116_),
    .Y(_02416_),
    .A1(net407),
    .A2(_06115_));
 sg13g2_nand2_1 _24796_ (.Y(_06117_),
    .A(_06097_),
    .B(\mem.mem_internal.data_mem[9][5] ));
 sg13g2_nand2_1 _24797_ (.Y(_06118_),
    .A(net1287),
    .B(_06105_));
 sg13g2_o21ai_1 _24798_ (.B1(_06118_),
    .Y(_02417_),
    .A1(_06106_),
    .A2(_06117_));
 sg13g2_nand2_1 _24799_ (.Y(_06119_),
    .A(net821),
    .B(\mem.mem_internal.data_mem[9][6] ));
 sg13g2_nand2_1 _24800_ (.Y(_06120_),
    .A(net1286),
    .B(_06105_));
 sg13g2_o21ai_1 _24801_ (.B1(_06120_),
    .Y(_02418_),
    .A1(_06106_),
    .A2(_06119_));
 sg13g2_nand2_1 _24802_ (.Y(_06121_),
    .A(_10226_),
    .B(\mem.mem_internal.data_mem[9][7] ));
 sg13g2_nand2_1 _24803_ (.Y(_06122_),
    .A(net1285),
    .B(_06105_));
 sg13g2_o21ai_1 _24804_ (.B1(_06122_),
    .Y(_02419_),
    .A1(net407),
    .A2(_06121_));
 sg13g2_o21ai_1 _24805_ (.B1(_09991_),
    .Y(_06123_),
    .A1(_10032_),
    .A2(_10035_));
 sg13g2_nor3_1 _24806_ (.A(_10237_),
    .B(_10238_),
    .C(_10236_),
    .Y(_06124_));
 sg13g2_o21ai_1 _24807_ (.B1(net1276),
    .Y(_06125_),
    .A1(_06123_),
    .A2(_06124_));
 sg13g2_buf_2 _24808_ (.A(_06125_),
    .X(_06126_));
 sg13g2_buf_1 _24809_ (.A(_06126_),
    .X(_06127_));
 sg13g2_buf_2 _24810_ (.A(_00000_),
    .X(_06128_));
 sg13g2_buf_1 _24811_ (.A(_06128_),
    .X(_06129_));
 sg13g2_buf_2 _24812_ (.A(_06129_),
    .X(_06130_));
 sg13g2_buf_1 _24813_ (.A(net990),
    .X(_06131_));
 sg13g2_buf_4 _24814_ (.X(_06132_),
    .A(net820));
 sg13g2_buf_2 _24815_ (.A(_06132_),
    .X(_06133_));
 sg13g2_buf_1 _24816_ (.A(_00001_),
    .X(_06134_));
 sg13g2_buf_2 _24817_ (.A(_06134_),
    .X(_06135_));
 sg13g2_buf_1 _24818_ (.A(_06135_),
    .X(_06136_));
 sg13g2_buf_1 _24819_ (.A(net989),
    .X(_06137_));
 sg13g2_buf_1 _24820_ (.A(net819),
    .X(_06138_));
 sg13g2_buf_1 _24821_ (.A(net578),
    .X(_06139_));
 sg13g2_mux4_1 _24822_ (.S0(net545),
    .A0(\mem.mem_internal.data_mem[0][0] ),
    .A1(\mem.mem_internal.data_mem[1][0] ),
    .A2(\mem.mem_internal.data_mem[2][0] ),
    .A3(\mem.mem_internal.data_mem[3][0] ),
    .S1(net544),
    .X(_06140_));
 sg13g2_mux4_1 _24823_ (.S0(net545),
    .A0(\mem.mem_internal.data_mem[4][0] ),
    .A1(\mem.mem_internal.data_mem[5][0] ),
    .A2(\mem.mem_internal.data_mem[6][0] ),
    .A3(\mem.mem_internal.data_mem[7][0] ),
    .S1(net544),
    .X(_06141_));
 sg13g2_buf_2 _24824_ (.A(net820),
    .X(_06142_));
 sg13g2_buf_1 _24825_ (.A(net578),
    .X(_06143_));
 sg13g2_mux4_1 _24826_ (.S0(net577),
    .A0(\mem.mem_internal.data_mem[16][0] ),
    .A1(\mem.mem_internal.data_mem[17][0] ),
    .A2(\mem.mem_internal.data_mem[18][0] ),
    .A3(\mem.mem_internal.data_mem[19][0] ),
    .S1(net543),
    .X(_06144_));
 sg13g2_buf_2 _24827_ (.A(_06132_),
    .X(_06145_));
 sg13g2_buf_1 _24828_ (.A(net578),
    .X(_06146_));
 sg13g2_mux4_1 _24829_ (.S0(net542),
    .A0(\mem.mem_internal.data_mem[20][0] ),
    .A1(\mem.mem_internal.data_mem[21][0] ),
    .A2(\mem.mem_internal.data_mem[22][0] ),
    .A3(\mem.mem_internal.data_mem[23][0] ),
    .S1(net541),
    .X(_06147_));
 sg13g2_buf_1 _24830_ (.A(_00002_),
    .X(_06148_));
 sg13g2_buf_1 _24831_ (.A(_06148_),
    .X(_06149_));
 sg13g2_buf_2 _24832_ (.A(net1236),
    .X(_06150_));
 sg13g2_buf_2 _24833_ (.A(net988),
    .X(_06151_));
 sg13g2_buf_1 _24834_ (.A(_00004_),
    .X(_06152_));
 sg13g2_buf_2 _24835_ (.A(_06152_),
    .X(_06153_));
 sg13g2_buf_1 _24836_ (.A(_06153_),
    .X(_06154_));
 sg13g2_buf_1 _24837_ (.A(net987),
    .X(_06155_));
 sg13g2_mux4_1 _24838_ (.S0(net818),
    .A0(_06140_),
    .A1(_06141_),
    .A2(_06144_),
    .A3(_06147_),
    .S1(net817),
    .X(_06156_));
 sg13g2_buf_2 _24839_ (.A(_06132_),
    .X(_06157_));
 sg13g2_buf_1 _24840_ (.A(net578),
    .X(_06158_));
 sg13g2_mux4_1 _24841_ (.S0(net540),
    .A0(\mem.mem_internal.data_mem[8][0] ),
    .A1(\mem.mem_internal.data_mem[9][0] ),
    .A2(\mem.mem_internal.data_mem[10][0] ),
    .A3(\mem.mem_internal.data_mem[11][0] ),
    .S1(net539),
    .X(_06159_));
 sg13g2_buf_2 _24842_ (.A(_06132_),
    .X(_06160_));
 sg13g2_buf_1 _24843_ (.A(_06138_),
    .X(_06161_));
 sg13g2_mux4_1 _24844_ (.S0(_06160_),
    .A0(\mem.mem_internal.data_mem[12][0] ),
    .A1(\mem.mem_internal.data_mem[13][0] ),
    .A2(\mem.mem_internal.data_mem[14][0] ),
    .A3(\mem.mem_internal.data_mem[15][0] ),
    .S1(_06161_),
    .X(_06162_));
 sg13g2_buf_2 _24845_ (.A(net820),
    .X(_06163_));
 sg13g2_buf_1 _24846_ (.A(net819),
    .X(_06164_));
 sg13g2_mux4_1 _24847_ (.S0(net576),
    .A0(\mem.mem_internal.data_mem[24][0] ),
    .A1(\mem.mem_internal.data_mem[25][0] ),
    .A2(\mem.mem_internal.data_mem[26][0] ),
    .A3(\mem.mem_internal.data_mem[27][0] ),
    .S1(net575),
    .X(_06165_));
 sg13g2_mux4_1 _24848_ (.S0(net577),
    .A0(\mem.mem_internal.data_mem[28][0] ),
    .A1(\mem.mem_internal.data_mem[29][0] ),
    .A2(\mem.mem_internal.data_mem[30][0] ),
    .A3(\mem.mem_internal.data_mem[31][0] ),
    .S1(net543),
    .X(_06166_));
 sg13g2_mux4_1 _24849_ (.S0(net818),
    .A0(_06159_),
    .A1(_06162_),
    .A2(_06165_),
    .A3(_06166_),
    .S1(net817),
    .X(_06167_));
 sg13g2_buf_4 _24850_ (.X(_06168_),
    .A(_00003_));
 sg13g2_buf_2 _24851_ (.A(_06168_),
    .X(_06169_));
 sg13g2_buf_1 _24852_ (.A(net1235),
    .X(_06170_));
 sg13g2_mux2_1 _24853_ (.A0(_06156_),
    .A1(_06167_),
    .S(net986),
    .X(_06171_));
 sg13g2_buf_2 _24854_ (.A(_06128_),
    .X(_06172_));
 sg13g2_buf_2 _24855_ (.A(_06172_),
    .X(_06173_));
 sg13g2_buf_2 _24856_ (.A(_06135_),
    .X(_06174_));
 sg13g2_buf_1 _24857_ (.A(_06174_),
    .X(_06175_));
 sg13g2_mux4_1 _24858_ (.S0(net985),
    .A0(\mem.mem_internal.code_mem[0][0] ),
    .A1(\mem.mem_internal.code_mem[1][0] ),
    .A2(\mem.mem_internal.code_mem[2][0] ),
    .A3(\mem.mem_internal.code_mem[3][0] ),
    .S1(net816),
    .X(_06176_));
 sg13g2_buf_1 _24859_ (.A(_06128_),
    .X(_06177_));
 sg13g2_buf_2 _24860_ (.A(_06177_),
    .X(_06178_));
 sg13g2_buf_1 _24861_ (.A(_06174_),
    .X(_06179_));
 sg13g2_mux4_1 _24862_ (.S0(net984),
    .A0(\mem.mem_internal.code_mem[4][0] ),
    .A1(\mem.mem_internal.code_mem[5][0] ),
    .A2(\mem.mem_internal.code_mem[6][0] ),
    .A3(\mem.mem_internal.code_mem[7][0] ),
    .S1(net815),
    .X(_06180_));
 sg13g2_buf_1 _24863_ (.A(_06128_),
    .X(_06181_));
 sg13g2_buf_2 _24864_ (.A(_06181_),
    .X(_06182_));
 sg13g2_buf_1 _24865_ (.A(_06134_),
    .X(_06183_));
 sg13g2_buf_1 _24866_ (.A(_06183_),
    .X(_06184_));
 sg13g2_mux4_1 _24867_ (.S0(net983),
    .A0(\mem.mem_internal.code_mem[16][0] ),
    .A1(\mem.mem_internal.code_mem[17][0] ),
    .A2(\mem.mem_internal.code_mem[18][0] ),
    .A3(\mem.mem_internal.code_mem[19][0] ),
    .S1(net982),
    .X(_06185_));
 sg13g2_buf_2 _24868_ (.A(_06181_),
    .X(_06186_));
 sg13g2_buf_2 _24869_ (.A(_06134_),
    .X(_06187_));
 sg13g2_buf_2 _24870_ (.A(_06187_),
    .X(_06188_));
 sg13g2_mux4_1 _24871_ (.S0(net981),
    .A0(\mem.mem_internal.code_mem[20][0] ),
    .A1(\mem.mem_internal.code_mem[21][0] ),
    .A2(\mem.mem_internal.code_mem[22][0] ),
    .A3(\mem.mem_internal.code_mem[23][0] ),
    .S1(_06188_),
    .X(_06189_));
 sg13g2_buf_2 _24872_ (.A(net1236),
    .X(_06190_));
 sg13g2_buf_1 _24873_ (.A(_06153_),
    .X(_06191_));
 sg13g2_mux4_1 _24874_ (.S0(net979),
    .A0(_06176_),
    .A1(_06180_),
    .A2(_06185_),
    .A3(_06189_),
    .S1(net978),
    .X(_06192_));
 sg13g2_mux4_1 _24875_ (.S0(_06178_),
    .A0(\mem.mem_internal.code_mem[8][0] ),
    .A1(\mem.mem_internal.code_mem[9][0] ),
    .A2(\mem.mem_internal.code_mem[10][0] ),
    .A3(\mem.mem_internal.code_mem[11][0] ),
    .S1(_06179_),
    .X(_06193_));
 sg13g2_mux4_1 _24876_ (.S0(_06178_),
    .A0(\mem.mem_internal.code_mem[12][0] ),
    .A1(\mem.mem_internal.code_mem[13][0] ),
    .A2(\mem.mem_internal.code_mem[14][0] ),
    .A3(\mem.mem_internal.code_mem[15][0] ),
    .S1(_06179_),
    .X(_06194_));
 sg13g2_buf_2 _24877_ (.A(_06181_),
    .X(_06195_));
 sg13g2_buf_2 _24878_ (.A(_06187_),
    .X(_06196_));
 sg13g2_mux4_1 _24879_ (.S0(net977),
    .A0(\mem.mem_internal.code_mem[24][0] ),
    .A1(\mem.mem_internal.code_mem[25][0] ),
    .A2(\mem.mem_internal.code_mem[26][0] ),
    .A3(\mem.mem_internal.code_mem[27][0] ),
    .S1(net976),
    .X(_06197_));
 sg13g2_mux4_1 _24880_ (.S0(net977),
    .A0(\mem.mem_internal.code_mem[28][0] ),
    .A1(\mem.mem_internal.code_mem[29][0] ),
    .A2(\mem.mem_internal.code_mem[30][0] ),
    .A3(\mem.mem_internal.code_mem[31][0] ),
    .S1(net976),
    .X(_06198_));
 sg13g2_mux4_1 _24881_ (.S0(net979),
    .A0(_06193_),
    .A1(_06194_),
    .A2(_06197_),
    .A3(_06198_),
    .S1(_06191_),
    .X(_06199_));
 sg13g2_mux4_1 _24882_ (.S0(net983),
    .A0(\mem.mem_internal.code_mem[128][0] ),
    .A1(\mem.mem_internal.code_mem[129][0] ),
    .A2(\mem.mem_internal.code_mem[130][0] ),
    .A3(\mem.mem_internal.code_mem[131][0] ),
    .S1(_06184_),
    .X(_06200_));
 sg13g2_mux4_1 _24883_ (.S0(_06186_),
    .A0(\mem.mem_internal.code_mem[132][0] ),
    .A1(\mem.mem_internal.code_mem[133][0] ),
    .A2(\mem.mem_internal.code_mem[134][0] ),
    .A3(\mem.mem_internal.code_mem[135][0] ),
    .S1(net976),
    .X(_06201_));
 sg13g2_buf_2 _24884_ (.A(_06129_),
    .X(_06202_));
 sg13g2_buf_2 _24885_ (.A(_06134_),
    .X(_06203_));
 sg13g2_buf_1 _24886_ (.A(_06203_),
    .X(_06204_));
 sg13g2_mux4_1 _24887_ (.S0(net975),
    .A0(\mem.mem_internal.code_mem[144][0] ),
    .A1(\mem.mem_internal.code_mem[145][0] ),
    .A2(\mem.mem_internal.code_mem[146][0] ),
    .A3(\mem.mem_internal.code_mem[147][0] ),
    .S1(net974),
    .X(_06205_));
 sg13g2_buf_2 _24888_ (.A(_06128_),
    .X(_06206_));
 sg13g2_buf_2 _24889_ (.A(_06206_),
    .X(_06207_));
 sg13g2_buf_1 _24890_ (.A(_06203_),
    .X(_06208_));
 sg13g2_mux4_1 _24891_ (.S0(net973),
    .A0(\mem.mem_internal.code_mem[148][0] ),
    .A1(\mem.mem_internal.code_mem[149][0] ),
    .A2(\mem.mem_internal.code_mem[150][0] ),
    .A3(\mem.mem_internal.code_mem[151][0] ),
    .S1(net972),
    .X(_06209_));
 sg13g2_buf_1 _24892_ (.A(_06148_),
    .X(_06210_));
 sg13g2_buf_2 _24893_ (.A(_06210_),
    .X(_06211_));
 sg13g2_buf_2 _24894_ (.A(_06152_),
    .X(_06212_));
 sg13g2_buf_1 _24895_ (.A(_06212_),
    .X(_06213_));
 sg13g2_mux4_1 _24896_ (.S0(net971),
    .A0(_06200_),
    .A1(_06201_),
    .A2(_06205_),
    .A3(_06209_),
    .S1(net970),
    .X(_06214_));
 sg13g2_mux4_1 _24897_ (.S0(net981),
    .A0(\mem.mem_internal.code_mem[136][0] ),
    .A1(\mem.mem_internal.code_mem[137][0] ),
    .A2(\mem.mem_internal.code_mem[138][0] ),
    .A3(\mem.mem_internal.code_mem[139][0] ),
    .S1(net980),
    .X(_06215_));
 sg13g2_mux4_1 _24898_ (.S0(net977),
    .A0(\mem.mem_internal.code_mem[140][0] ),
    .A1(\mem.mem_internal.code_mem[141][0] ),
    .A2(\mem.mem_internal.code_mem[142][0] ),
    .A3(\mem.mem_internal.code_mem[143][0] ),
    .S1(_06196_),
    .X(_06216_));
 sg13g2_mux4_1 _24899_ (.S0(net973),
    .A0(\mem.mem_internal.code_mem[152][0] ),
    .A1(\mem.mem_internal.code_mem[153][0] ),
    .A2(\mem.mem_internal.code_mem[154][0] ),
    .A3(\mem.mem_internal.code_mem[155][0] ),
    .S1(net972),
    .X(_06217_));
 sg13g2_buf_2 _24900_ (.A(_06206_),
    .X(_06218_));
 sg13g2_buf_2 _24901_ (.A(_06203_),
    .X(_06219_));
 sg13g2_mux4_1 _24902_ (.S0(net969),
    .A0(\mem.mem_internal.code_mem[156][0] ),
    .A1(\mem.mem_internal.code_mem[157][0] ),
    .A2(\mem.mem_internal.code_mem[158][0] ),
    .A3(\mem.mem_internal.code_mem[159][0] ),
    .S1(net968),
    .X(_06220_));
 sg13g2_buf_2 _24903_ (.A(_06210_),
    .X(_06221_));
 sg13g2_mux4_1 _24904_ (.S0(net967),
    .A0(_06215_),
    .A1(_06216_),
    .A2(_06217_),
    .A3(_06220_),
    .S1(net970),
    .X(_06222_));
 sg13g2_buf_2 _24905_ (.A(_06168_),
    .X(_06223_));
 sg13g2_buf_1 _24906_ (.A(_00007_),
    .X(_06224_));
 sg13g2_buf_1 _24907_ (.A(_06224_),
    .X(_06225_));
 sg13g2_mux4_1 _24908_ (.S0(net1234),
    .A0(_06192_),
    .A1(_06199_),
    .A2(_06214_),
    .A3(_06222_),
    .S1(net1233),
    .X(_06226_));
 sg13g2_mux4_1 _24909_ (.S0(net984),
    .A0(\mem.mem_internal.code_mem[32][0] ),
    .A1(\mem.mem_internal.code_mem[33][0] ),
    .A2(\mem.mem_internal.code_mem[34][0] ),
    .A3(\mem.mem_internal.code_mem[35][0] ),
    .S1(net815),
    .X(_06227_));
 sg13g2_mux4_1 _24910_ (.S0(net984),
    .A0(\mem.mem_internal.code_mem[36][0] ),
    .A1(\mem.mem_internal.code_mem[37][0] ),
    .A2(\mem.mem_internal.code_mem[38][0] ),
    .A3(\mem.mem_internal.code_mem[39][0] ),
    .S1(net815),
    .X(_06228_));
 sg13g2_mux4_1 _24911_ (.S0(net981),
    .A0(\mem.mem_internal.code_mem[48][0] ),
    .A1(\mem.mem_internal.code_mem[49][0] ),
    .A2(\mem.mem_internal.code_mem[50][0] ),
    .A3(\mem.mem_internal.code_mem[51][0] ),
    .S1(net976),
    .X(_06229_));
 sg13g2_mux4_1 _24912_ (.S0(net977),
    .A0(\mem.mem_internal.code_mem[52][0] ),
    .A1(\mem.mem_internal.code_mem[53][0] ),
    .A2(\mem.mem_internal.code_mem[54][0] ),
    .A3(\mem.mem_internal.code_mem[55][0] ),
    .S1(net976),
    .X(_06230_));
 sg13g2_mux4_1 _24913_ (.S0(net979),
    .A0(_06227_),
    .A1(_06228_),
    .A2(_06229_),
    .A3(_06230_),
    .S1(net978),
    .X(_06231_));
 sg13g2_buf_1 _24914_ (.A(_06174_),
    .X(_06232_));
 sg13g2_mux4_1 _24915_ (.S0(net984),
    .A0(\mem.mem_internal.code_mem[40][0] ),
    .A1(\mem.mem_internal.code_mem[41][0] ),
    .A2(\mem.mem_internal.code_mem[42][0] ),
    .A3(\mem.mem_internal.code_mem[43][0] ),
    .S1(net814),
    .X(_06233_));
 sg13g2_mux4_1 _24916_ (.S0(net984),
    .A0(\mem.mem_internal.code_mem[44][0] ),
    .A1(\mem.mem_internal.code_mem[45][0] ),
    .A2(\mem.mem_internal.code_mem[46][0] ),
    .A3(\mem.mem_internal.code_mem[47][0] ),
    .S1(net814),
    .X(_06234_));
 sg13g2_buf_2 _24917_ (.A(_06187_),
    .X(_06235_));
 sg13g2_mux4_1 _24918_ (.S0(net977),
    .A0(\mem.mem_internal.code_mem[56][0] ),
    .A1(\mem.mem_internal.code_mem[57][0] ),
    .A2(\mem.mem_internal.code_mem[58][0] ),
    .A3(\mem.mem_internal.code_mem[59][0] ),
    .S1(net966),
    .X(_06236_));
 sg13g2_buf_1 _24919_ (.A(_06128_),
    .X(_06237_));
 sg13g2_buf_2 _24920_ (.A(_06237_),
    .X(_06238_));
 sg13g2_mux4_1 _24921_ (.S0(net965),
    .A0(\mem.mem_internal.code_mem[60][0] ),
    .A1(\mem.mem_internal.code_mem[61][0] ),
    .A2(\mem.mem_internal.code_mem[62][0] ),
    .A3(\mem.mem_internal.code_mem[63][0] ),
    .S1(net966),
    .X(_06239_));
 sg13g2_mux4_1 _24922_ (.S0(net979),
    .A0(_06233_),
    .A1(_06234_),
    .A2(_06236_),
    .A3(_06239_),
    .S1(net978),
    .X(_06240_));
 sg13g2_mux4_1 _24923_ (.S0(net977),
    .A0(\mem.mem_internal.code_mem[160][0] ),
    .A1(\mem.mem_internal.code_mem[161][0] ),
    .A2(\mem.mem_internal.code_mem[162][0] ),
    .A3(\mem.mem_internal.code_mem[163][0] ),
    .S1(net976),
    .X(_06241_));
 sg13g2_mux4_1 _24924_ (.S0(net965),
    .A0(\mem.mem_internal.code_mem[164][0] ),
    .A1(\mem.mem_internal.code_mem[165][0] ),
    .A2(\mem.mem_internal.code_mem[166][0] ),
    .A3(\mem.mem_internal.code_mem[167][0] ),
    .S1(net966),
    .X(_06242_));
 sg13g2_mux4_1 _24925_ (.S0(net973),
    .A0(\mem.mem_internal.code_mem[176][0] ),
    .A1(\mem.mem_internal.code_mem[177][0] ),
    .A2(\mem.mem_internal.code_mem[178][0] ),
    .A3(\mem.mem_internal.code_mem[179][0] ),
    .S1(net968),
    .X(_06243_));
 sg13g2_buf_2 _24926_ (.A(_06203_),
    .X(_06244_));
 sg13g2_mux4_1 _24927_ (.S0(net969),
    .A0(\mem.mem_internal.code_mem[180][0] ),
    .A1(\mem.mem_internal.code_mem[181][0] ),
    .A2(\mem.mem_internal.code_mem[182][0] ),
    .A3(\mem.mem_internal.code_mem[183][0] ),
    .S1(net964),
    .X(_06245_));
 sg13g2_mux4_1 _24928_ (.S0(net967),
    .A0(_06241_),
    .A1(_06242_),
    .A2(_06243_),
    .A3(_06245_),
    .S1(net970),
    .X(_06246_));
 sg13g2_mux4_1 _24929_ (.S0(net977),
    .A0(\mem.mem_internal.code_mem[168][0] ),
    .A1(\mem.mem_internal.code_mem[169][0] ),
    .A2(\mem.mem_internal.code_mem[170][0] ),
    .A3(\mem.mem_internal.code_mem[171][0] ),
    .S1(net976),
    .X(_06247_));
 sg13g2_mux4_1 _24930_ (.S0(net965),
    .A0(\mem.mem_internal.code_mem[172][0] ),
    .A1(\mem.mem_internal.code_mem[173][0] ),
    .A2(\mem.mem_internal.code_mem[174][0] ),
    .A3(\mem.mem_internal.code_mem[175][0] ),
    .S1(net966),
    .X(_06248_));
 sg13g2_mux4_1 _24931_ (.S0(net969),
    .A0(\mem.mem_internal.code_mem[184][0] ),
    .A1(\mem.mem_internal.code_mem[185][0] ),
    .A2(\mem.mem_internal.code_mem[186][0] ),
    .A3(\mem.mem_internal.code_mem[187][0] ),
    .S1(net968),
    .X(_06249_));
 sg13g2_buf_2 _24932_ (.A(_06206_),
    .X(_06250_));
 sg13g2_mux4_1 _24933_ (.S0(net963),
    .A0(\mem.mem_internal.code_mem[188][0] ),
    .A1(\mem.mem_internal.code_mem[189][0] ),
    .A2(\mem.mem_internal.code_mem[190][0] ),
    .A3(\mem.mem_internal.code_mem[191][0] ),
    .S1(net964),
    .X(_06251_));
 sg13g2_mux4_1 _24934_ (.S0(net967),
    .A0(_06247_),
    .A1(_06248_),
    .A2(_06249_),
    .A3(_06251_),
    .S1(net970),
    .X(_06252_));
 sg13g2_mux4_1 _24935_ (.S0(net1234),
    .A0(_06231_),
    .A1(_06240_),
    .A2(_06246_),
    .A3(_06252_),
    .S1(net1233),
    .X(_06253_));
 sg13g2_buf_2 _24936_ (.A(_06181_),
    .X(_06254_));
 sg13g2_mux4_1 _24937_ (.S0(_06254_),
    .A0(\mem.mem_internal.code_mem[64][0] ),
    .A1(\mem.mem_internal.code_mem[65][0] ),
    .A2(\mem.mem_internal.code_mem[66][0] ),
    .A3(\mem.mem_internal.code_mem[67][0] ),
    .S1(net982),
    .X(_06255_));
 sg13g2_mux4_1 _24938_ (.S0(net981),
    .A0(\mem.mem_internal.code_mem[68][0] ),
    .A1(\mem.mem_internal.code_mem[69][0] ),
    .A2(\mem.mem_internal.code_mem[70][0] ),
    .A3(\mem.mem_internal.code_mem[71][0] ),
    .S1(net980),
    .X(_06256_));
 sg13g2_mux4_1 _24939_ (.S0(net975),
    .A0(\mem.mem_internal.code_mem[80][0] ),
    .A1(\mem.mem_internal.code_mem[81][0] ),
    .A2(\mem.mem_internal.code_mem[82][0] ),
    .A3(\mem.mem_internal.code_mem[83][0] ),
    .S1(net974),
    .X(_06257_));
 sg13g2_mux4_1 _24940_ (.S0(net973),
    .A0(\mem.mem_internal.code_mem[84][0] ),
    .A1(\mem.mem_internal.code_mem[85][0] ),
    .A2(\mem.mem_internal.code_mem[86][0] ),
    .A3(\mem.mem_internal.code_mem[87][0] ),
    .S1(net972),
    .X(_06258_));
 sg13g2_mux4_1 _24941_ (.S0(net971),
    .A0(_06255_),
    .A1(_06256_),
    .A2(_06257_),
    .A3(_06258_),
    .S1(net970),
    .X(_06259_));
 sg13g2_mux4_1 _24942_ (.S0(net981),
    .A0(\mem.mem_internal.code_mem[72][0] ),
    .A1(\mem.mem_internal.code_mem[73][0] ),
    .A2(\mem.mem_internal.code_mem[74][0] ),
    .A3(\mem.mem_internal.code_mem[75][0] ),
    .S1(net980),
    .X(_06260_));
 sg13g2_mux4_1 _24943_ (.S0(_06195_),
    .A0(\mem.mem_internal.code_mem[76][0] ),
    .A1(\mem.mem_internal.code_mem[77][0] ),
    .A2(\mem.mem_internal.code_mem[78][0] ),
    .A3(\mem.mem_internal.code_mem[79][0] ),
    .S1(_06235_),
    .X(_06261_));
 sg13g2_mux4_1 _24944_ (.S0(_06207_),
    .A0(\mem.mem_internal.code_mem[88][0] ),
    .A1(\mem.mem_internal.code_mem[89][0] ),
    .A2(\mem.mem_internal.code_mem[90][0] ),
    .A3(\mem.mem_internal.code_mem[91][0] ),
    .S1(_06219_),
    .X(_06262_));
 sg13g2_mux4_1 _24945_ (.S0(_06218_),
    .A0(\mem.mem_internal.code_mem[92][0] ),
    .A1(\mem.mem_internal.code_mem[93][0] ),
    .A2(\mem.mem_internal.code_mem[94][0] ),
    .A3(\mem.mem_internal.code_mem[95][0] ),
    .S1(net968),
    .X(_06263_));
 sg13g2_mux4_1 _24946_ (.S0(net967),
    .A0(_06260_),
    .A1(_06261_),
    .A2(_06262_),
    .A3(_06263_),
    .S1(net970),
    .X(_06264_));
 sg13g2_mux4_1 _24947_ (.S0(net975),
    .A0(\mem.mem_internal.code_mem[192][0] ),
    .A1(\mem.mem_internal.code_mem[193][0] ),
    .A2(\mem.mem_internal.code_mem[194][0] ),
    .A3(\mem.mem_internal.code_mem[195][0] ),
    .S1(net974),
    .X(_06265_));
 sg13g2_mux4_1 _24948_ (.S0(net973),
    .A0(\mem.mem_internal.code_mem[196][0] ),
    .A1(\mem.mem_internal.code_mem[197][0] ),
    .A2(\mem.mem_internal.code_mem[198][0] ),
    .A3(\mem.mem_internal.code_mem[199][0] ),
    .S1(net972),
    .X(_06266_));
 sg13g2_mux4_1 _24949_ (.S0(net990),
    .A0(\mem.mem_internal.code_mem[208][0] ),
    .A1(\mem.mem_internal.code_mem[209][0] ),
    .A2(\mem.mem_internal.code_mem[210][0] ),
    .A3(\mem.mem_internal.code_mem[211][0] ),
    .S1(net989),
    .X(_06267_));
 sg13g2_mux4_1 _24950_ (.S0(net990),
    .A0(\mem.mem_internal.code_mem[212][0] ),
    .A1(\mem.mem_internal.code_mem[213][0] ),
    .A2(\mem.mem_internal.code_mem[214][0] ),
    .A3(\mem.mem_internal.code_mem[215][0] ),
    .S1(net989),
    .X(_06268_));
 sg13g2_mux4_1 _24951_ (.S0(net1236),
    .A0(_06265_),
    .A1(_06266_),
    .A2(_06267_),
    .A3(_06268_),
    .S1(_06153_),
    .X(_06269_));
 sg13g2_mux4_1 _24952_ (.S0(net973),
    .A0(\mem.mem_internal.code_mem[200][0] ),
    .A1(\mem.mem_internal.code_mem[201][0] ),
    .A2(\mem.mem_internal.code_mem[202][0] ),
    .A3(\mem.mem_internal.code_mem[203][0] ),
    .S1(net972),
    .X(_06270_));
 sg13g2_mux4_1 _24953_ (.S0(net969),
    .A0(\mem.mem_internal.code_mem[204][0] ),
    .A1(\mem.mem_internal.code_mem[205][0] ),
    .A2(\mem.mem_internal.code_mem[206][0] ),
    .A3(\mem.mem_internal.code_mem[207][0] ),
    .S1(net968),
    .X(_06271_));
 sg13g2_mux4_1 _24954_ (.S0(net990),
    .A0(\mem.mem_internal.code_mem[216][0] ),
    .A1(\mem.mem_internal.code_mem[217][0] ),
    .A2(\mem.mem_internal.code_mem[218][0] ),
    .A3(\mem.mem_internal.code_mem[219][0] ),
    .S1(net989),
    .X(_06272_));
 sg13g2_buf_1 _24955_ (.A(_06135_),
    .X(_06273_));
 sg13g2_mux4_1 _24956_ (.S0(net990),
    .A0(\mem.mem_internal.code_mem[220][0] ),
    .A1(\mem.mem_internal.code_mem[221][0] ),
    .A2(\mem.mem_internal.code_mem[222][0] ),
    .A3(\mem.mem_internal.code_mem[223][0] ),
    .S1(_06273_),
    .X(_06274_));
 sg13g2_buf_1 _24957_ (.A(_06212_),
    .X(_06275_));
 sg13g2_mux4_1 _24958_ (.S0(net1236),
    .A0(_06270_),
    .A1(_06271_),
    .A2(_06272_),
    .A3(_06274_),
    .S1(net960),
    .X(_06276_));
 sg13g2_mux4_1 _24959_ (.S0(_06168_),
    .A0(_06259_),
    .A1(_06264_),
    .A2(_06269_),
    .A3(_06276_),
    .S1(_06224_),
    .X(_06277_));
 sg13g2_mux4_1 _24960_ (.S0(_06186_),
    .A0(\mem.mem_internal.code_mem[96][0] ),
    .A1(\mem.mem_internal.code_mem[97][0] ),
    .A2(\mem.mem_internal.code_mem[98][0] ),
    .A3(\mem.mem_internal.code_mem[99][0] ),
    .S1(_06188_),
    .X(_06278_));
 sg13g2_mux4_1 _24961_ (.S0(_06195_),
    .A0(\mem.mem_internal.code_mem[100][0] ),
    .A1(\mem.mem_internal.code_mem[101][0] ),
    .A2(\mem.mem_internal.code_mem[102][0] ),
    .A3(\mem.mem_internal.code_mem[103][0] ),
    .S1(_06196_),
    .X(_06279_));
 sg13g2_mux4_1 _24962_ (.S0(net973),
    .A0(\mem.mem_internal.code_mem[112][0] ),
    .A1(\mem.mem_internal.code_mem[113][0] ),
    .A2(\mem.mem_internal.code_mem[114][0] ),
    .A3(\mem.mem_internal.code_mem[115][0] ),
    .S1(net972),
    .X(_06280_));
 sg13g2_mux4_1 _24963_ (.S0(net969),
    .A0(\mem.mem_internal.code_mem[116][0] ),
    .A1(\mem.mem_internal.code_mem[117][0] ),
    .A2(\mem.mem_internal.code_mem[118][0] ),
    .A3(\mem.mem_internal.code_mem[119][0] ),
    .S1(net968),
    .X(_06281_));
 sg13g2_mux4_1 _24964_ (.S0(net971),
    .A0(_06278_),
    .A1(_06279_),
    .A2(_06280_),
    .A3(_06281_),
    .S1(_06213_),
    .X(_06282_));
 sg13g2_mux4_1 _24965_ (.S0(net977),
    .A0(\mem.mem_internal.code_mem[104][0] ),
    .A1(\mem.mem_internal.code_mem[105][0] ),
    .A2(\mem.mem_internal.code_mem[106][0] ),
    .A3(\mem.mem_internal.code_mem[107][0] ),
    .S1(net976),
    .X(_06283_));
 sg13g2_mux4_1 _24966_ (.S0(_06238_),
    .A0(\mem.mem_internal.code_mem[108][0] ),
    .A1(\mem.mem_internal.code_mem[109][0] ),
    .A2(\mem.mem_internal.code_mem[110][0] ),
    .A3(\mem.mem_internal.code_mem[111][0] ),
    .S1(_06235_),
    .X(_06284_));
 sg13g2_mux4_1 _24967_ (.S0(net969),
    .A0(\mem.mem_internal.code_mem[120][0] ),
    .A1(\mem.mem_internal.code_mem[121][0] ),
    .A2(\mem.mem_internal.code_mem[122][0] ),
    .A3(\mem.mem_internal.code_mem[123][0] ),
    .S1(net968),
    .X(_06285_));
 sg13g2_mux4_1 _24968_ (.S0(net963),
    .A0(\mem.mem_internal.code_mem[124][0] ),
    .A1(\mem.mem_internal.code_mem[125][0] ),
    .A2(\mem.mem_internal.code_mem[126][0] ),
    .A3(\mem.mem_internal.code_mem[127][0] ),
    .S1(_06244_),
    .X(_06286_));
 sg13g2_mux4_1 _24969_ (.S0(net967),
    .A0(_06283_),
    .A1(_06284_),
    .A2(_06285_),
    .A3(_06286_),
    .S1(_06213_),
    .X(_06287_));
 sg13g2_mux4_1 _24970_ (.S0(net973),
    .A0(\mem.mem_internal.code_mem[224][0] ),
    .A1(\mem.mem_internal.code_mem[225][0] ),
    .A2(\mem.mem_internal.code_mem[226][0] ),
    .A3(\mem.mem_internal.code_mem[227][0] ),
    .S1(net972),
    .X(_06288_));
 sg13g2_mux4_1 _24971_ (.S0(net969),
    .A0(\mem.mem_internal.code_mem[228][0] ),
    .A1(\mem.mem_internal.code_mem[229][0] ),
    .A2(\mem.mem_internal.code_mem[230][0] ),
    .A3(\mem.mem_internal.code_mem[231][0] ),
    .S1(net968),
    .X(_06289_));
 sg13g2_mux4_1 _24972_ (.S0(net990),
    .A0(\mem.mem_internal.code_mem[240][0] ),
    .A1(\mem.mem_internal.code_mem[241][0] ),
    .A2(\mem.mem_internal.code_mem[242][0] ),
    .A3(\mem.mem_internal.code_mem[243][0] ),
    .S1(_06136_),
    .X(_06290_));
 sg13g2_buf_2 _24973_ (.A(_06129_),
    .X(_06291_));
 sg13g2_mux4_1 _24974_ (.S0(net959),
    .A0(\mem.mem_internal.code_mem[244][0] ),
    .A1(\mem.mem_internal.code_mem[245][0] ),
    .A2(\mem.mem_internal.code_mem[246][0] ),
    .A3(\mem.mem_internal.code_mem[247][0] ),
    .S1(net961),
    .X(_06292_));
 sg13g2_mux4_1 _24975_ (.S0(net1236),
    .A0(_06288_),
    .A1(_06289_),
    .A2(_06290_),
    .A3(_06292_),
    .S1(net960),
    .X(_06293_));
 sg13g2_mux4_1 _24976_ (.S0(net969),
    .A0(\mem.mem_internal.code_mem[232][0] ),
    .A1(\mem.mem_internal.code_mem[233][0] ),
    .A2(\mem.mem_internal.code_mem[234][0] ),
    .A3(\mem.mem_internal.code_mem[235][0] ),
    .S1(_06219_),
    .X(_06294_));
 sg13g2_mux4_1 _24977_ (.S0(_06218_),
    .A0(\mem.mem_internal.code_mem[236][0] ),
    .A1(\mem.mem_internal.code_mem[237][0] ),
    .A2(\mem.mem_internal.code_mem[238][0] ),
    .A3(\mem.mem_internal.code_mem[239][0] ),
    .S1(_06244_),
    .X(_06295_));
 sg13g2_mux4_1 _24978_ (.S0(_06130_),
    .A0(\mem.mem_internal.code_mem[248][0] ),
    .A1(\mem.mem_internal.code_mem[249][0] ),
    .A2(\mem.mem_internal.code_mem[250][0] ),
    .A3(\mem.mem_internal.code_mem[251][0] ),
    .S1(net961),
    .X(_06296_));
 sg13g2_mux4_1 _24979_ (.S0(net959),
    .A0(\mem.mem_internal.code_mem[252][0] ),
    .A1(\mem.mem_internal.code_mem[253][0] ),
    .A2(\mem.mem_internal.code_mem[254][0] ),
    .A3(\mem.mem_internal.code_mem[255][0] ),
    .S1(net961),
    .X(_06297_));
 sg13g2_mux4_1 _24980_ (.S0(net1236),
    .A0(_06294_),
    .A1(_06295_),
    .A2(_06296_),
    .A3(_06297_),
    .S1(net960),
    .X(_06298_));
 sg13g2_mux4_1 _24981_ (.S0(_06168_),
    .A0(_06282_),
    .A1(_06287_),
    .A2(_06293_),
    .A3(_06298_),
    .S1(_06224_),
    .X(_06299_));
 sg13g2_buf_4 _24982_ (.X(_06300_),
    .A(_00005_));
 sg13g2_buf_4 _24983_ (.X(_06301_),
    .A(_00006_));
 sg13g2_mux4_1 _24984_ (.S0(_06300_),
    .A0(_06226_),
    .A1(_06253_),
    .A2(_06277_),
    .A3(_06299_),
    .S1(_06301_),
    .X(_06302_));
 sg13g2_nand2b_1 _24985_ (.Y(_06303_),
    .B(_00080_),
    .A_N(_05432_));
 sg13g2_buf_2 _24986_ (.A(_06303_),
    .X(_06304_));
 sg13g2_nor2_1 _24987_ (.A(_06302_),
    .B(_06304_),
    .Y(_06305_));
 sg13g2_a21oi_1 _24988_ (.A1(net832),
    .A2(_06171_),
    .Y(_06306_),
    .B1(_06305_));
 sg13g2_nand2_1 _24989_ (.Y(_06307_),
    .A(\mem.internal_data_out[0] ),
    .B(net546));
 sg13g2_o21ai_1 _24990_ (.B1(_06307_),
    .Y(_02420_),
    .A1(net546),
    .A2(_06306_));
 sg13g2_mux4_1 _24991_ (.S0(net545),
    .A0(\mem.mem_internal.data_mem[0][1] ),
    .A1(\mem.mem_internal.data_mem[1][1] ),
    .A2(\mem.mem_internal.data_mem[2][1] ),
    .A3(\mem.mem_internal.data_mem[3][1] ),
    .S1(net544),
    .X(_06308_));
 sg13g2_mux4_1 _24992_ (.S0(net545),
    .A0(\mem.mem_internal.data_mem[4][1] ),
    .A1(\mem.mem_internal.data_mem[5][1] ),
    .A2(\mem.mem_internal.data_mem[6][1] ),
    .A3(\mem.mem_internal.data_mem[7][1] ),
    .S1(net544),
    .X(_06309_));
 sg13g2_mux4_1 _24993_ (.S0(net577),
    .A0(\mem.mem_internal.data_mem[8][1] ),
    .A1(\mem.mem_internal.data_mem[9][1] ),
    .A2(\mem.mem_internal.data_mem[10][1] ),
    .A3(\mem.mem_internal.data_mem[11][1] ),
    .S1(net543),
    .X(_06310_));
 sg13g2_mux4_1 _24994_ (.S0(net542),
    .A0(\mem.mem_internal.data_mem[12][1] ),
    .A1(\mem.mem_internal.data_mem[13][1] ),
    .A2(\mem.mem_internal.data_mem[14][1] ),
    .A3(\mem.mem_internal.data_mem[15][1] ),
    .S1(net541),
    .X(_06311_));
 sg13g2_mux4_1 _24995_ (.S0(net818),
    .A0(_06308_),
    .A1(_06309_),
    .A2(_06310_),
    .A3(_06311_),
    .S1(net986),
    .X(_06312_));
 sg13g2_mux4_1 _24996_ (.S0(net540),
    .A0(\mem.mem_internal.data_mem[16][1] ),
    .A1(\mem.mem_internal.data_mem[17][1] ),
    .A2(\mem.mem_internal.data_mem[18][1] ),
    .A3(\mem.mem_internal.data_mem[19][1] ),
    .S1(net539),
    .X(_06313_));
 sg13g2_mux4_1 _24997_ (.S0(net538),
    .A0(\mem.mem_internal.data_mem[20][1] ),
    .A1(\mem.mem_internal.data_mem[21][1] ),
    .A2(\mem.mem_internal.data_mem[22][1] ),
    .A3(\mem.mem_internal.data_mem[23][1] ),
    .S1(net537),
    .X(_06314_));
 sg13g2_mux4_1 _24998_ (.S0(net576),
    .A0(\mem.mem_internal.data_mem[24][1] ),
    .A1(\mem.mem_internal.data_mem[25][1] ),
    .A2(\mem.mem_internal.data_mem[26][1] ),
    .A3(\mem.mem_internal.data_mem[27][1] ),
    .S1(net575),
    .X(_06315_));
 sg13g2_mux4_1 _24999_ (.S0(net577),
    .A0(\mem.mem_internal.data_mem[28][1] ),
    .A1(\mem.mem_internal.data_mem[29][1] ),
    .A2(\mem.mem_internal.data_mem[30][1] ),
    .A3(\mem.mem_internal.data_mem[31][1] ),
    .S1(net543),
    .X(_06316_));
 sg13g2_mux4_1 _25000_ (.S0(net818),
    .A0(_06313_),
    .A1(_06314_),
    .A2(_06315_),
    .A3(_06316_),
    .S1(net986),
    .X(_06317_));
 sg13g2_mux2_1 _25001_ (.A0(_06312_),
    .A1(_06317_),
    .S(net817),
    .X(_06318_));
 sg13g2_buf_2 _25002_ (.A(_06177_),
    .X(_06319_));
 sg13g2_mux4_1 _25003_ (.S0(net958),
    .A0(\mem.mem_internal.code_mem[0][1] ),
    .A1(\mem.mem_internal.code_mem[1][1] ),
    .A2(\mem.mem_internal.code_mem[2][1] ),
    .A3(\mem.mem_internal.code_mem[3][1] ),
    .S1(net814),
    .X(_06320_));
 sg13g2_buf_2 _25004_ (.A(_06177_),
    .X(_06321_));
 sg13g2_buf_1 _25005_ (.A(net989),
    .X(_06322_));
 sg13g2_mux4_1 _25006_ (.S0(net957),
    .A0(\mem.mem_internal.code_mem[4][1] ),
    .A1(\mem.mem_internal.code_mem[5][1] ),
    .A2(\mem.mem_internal.code_mem[6][1] ),
    .A3(\mem.mem_internal.code_mem[7][1] ),
    .S1(net813),
    .X(_06323_));
 sg13g2_buf_2 _25007_ (.A(_06237_),
    .X(_06324_));
 sg13g2_buf_1 _25008_ (.A(_06187_),
    .X(_06325_));
 sg13g2_mux4_1 _25009_ (.S0(net956),
    .A0(\mem.mem_internal.code_mem[16][1] ),
    .A1(\mem.mem_internal.code_mem[17][1] ),
    .A2(\mem.mem_internal.code_mem[18][1] ),
    .A3(\mem.mem_internal.code_mem[19][1] ),
    .S1(net955),
    .X(_06326_));
 sg13g2_buf_2 _25010_ (.A(_06237_),
    .X(_06327_));
 sg13g2_buf_2 _25011_ (.A(_06187_),
    .X(_06328_));
 sg13g2_mux4_1 _25012_ (.S0(net954),
    .A0(\mem.mem_internal.code_mem[20][1] ),
    .A1(\mem.mem_internal.code_mem[21][1] ),
    .A2(\mem.mem_internal.code_mem[22][1] ),
    .A3(\mem.mem_internal.code_mem[23][1] ),
    .S1(net953),
    .X(_06329_));
 sg13g2_buf_2 _25013_ (.A(net1236),
    .X(_06330_));
 sg13g2_buf_1 _25014_ (.A(_06153_),
    .X(_06331_));
 sg13g2_mux4_1 _25015_ (.S0(net952),
    .A0(_06320_),
    .A1(_06323_),
    .A2(_06326_),
    .A3(_06329_),
    .S1(net951),
    .X(_06332_));
 sg13g2_buf_1 _25016_ (.A(net989),
    .X(_06333_));
 sg13g2_mux4_1 _25017_ (.S0(net957),
    .A0(\mem.mem_internal.code_mem[8][1] ),
    .A1(\mem.mem_internal.code_mem[9][1] ),
    .A2(\mem.mem_internal.code_mem[10][1] ),
    .A3(\mem.mem_internal.code_mem[11][1] ),
    .S1(net812),
    .X(_06334_));
 sg13g2_buf_2 _25018_ (.A(net990),
    .X(_06335_));
 sg13g2_buf_2 _25019_ (.A(net989),
    .X(_06336_));
 sg13g2_mux4_1 _25020_ (.S0(net811),
    .A0(\mem.mem_internal.code_mem[12][1] ),
    .A1(\mem.mem_internal.code_mem[13][1] ),
    .A2(\mem.mem_internal.code_mem[14][1] ),
    .A3(\mem.mem_internal.code_mem[15][1] ),
    .S1(net810),
    .X(_06337_));
 sg13g2_buf_2 _25021_ (.A(_06172_),
    .X(_06338_));
 sg13g2_buf_2 _25022_ (.A(_06135_),
    .X(_06339_));
 sg13g2_buf_1 _25023_ (.A(_06339_),
    .X(_06340_));
 sg13g2_mux4_1 _25024_ (.S0(net950),
    .A0(\mem.mem_internal.code_mem[24][1] ),
    .A1(\mem.mem_internal.code_mem[25][1] ),
    .A2(\mem.mem_internal.code_mem[26][1] ),
    .A3(\mem.mem_internal.code_mem[27][1] ),
    .S1(net809),
    .X(_06341_));
 sg13g2_buf_2 _25025_ (.A(_06172_),
    .X(_06342_));
 sg13g2_mux4_1 _25026_ (.S0(net949),
    .A0(\mem.mem_internal.code_mem[28][1] ),
    .A1(\mem.mem_internal.code_mem[29][1] ),
    .A2(\mem.mem_internal.code_mem[30][1] ),
    .A3(\mem.mem_internal.code_mem[31][1] ),
    .S1(net816),
    .X(_06343_));
 sg13g2_buf_2 _25027_ (.A(net1236),
    .X(_06344_));
 sg13g2_buf_1 _25028_ (.A(_06153_),
    .X(_06345_));
 sg13g2_mux4_1 _25029_ (.S0(net948),
    .A0(_06334_),
    .A1(_06337_),
    .A2(_06341_),
    .A3(_06343_),
    .S1(net947),
    .X(_06346_));
 sg13g2_buf_1 _25030_ (.A(_06187_),
    .X(_06347_));
 sg13g2_mux4_1 _25031_ (.S0(net956),
    .A0(\mem.mem_internal.code_mem[128][1] ),
    .A1(\mem.mem_internal.code_mem[129][1] ),
    .A2(\mem.mem_internal.code_mem[130][1] ),
    .A3(\mem.mem_internal.code_mem[131][1] ),
    .S1(net946),
    .X(_06348_));
 sg13g2_buf_2 _25032_ (.A(_06172_),
    .X(_06349_));
 sg13g2_buf_1 _25033_ (.A(_06339_),
    .X(_06350_));
 sg13g2_mux4_1 _25034_ (.S0(net945),
    .A0(\mem.mem_internal.code_mem[132][1] ),
    .A1(\mem.mem_internal.code_mem[133][1] ),
    .A2(\mem.mem_internal.code_mem[134][1] ),
    .A3(\mem.mem_internal.code_mem[135][1] ),
    .S1(net808),
    .X(_06351_));
 sg13g2_buf_2 _25035_ (.A(_06206_),
    .X(_06352_));
 sg13g2_buf_1 _25036_ (.A(_06203_),
    .X(_06353_));
 sg13g2_mux4_1 _25037_ (.S0(net944),
    .A0(\mem.mem_internal.code_mem[144][1] ),
    .A1(\mem.mem_internal.code_mem[145][1] ),
    .A2(\mem.mem_internal.code_mem[146][1] ),
    .A3(\mem.mem_internal.code_mem[147][1] ),
    .S1(net943),
    .X(_06354_));
 sg13g2_buf_1 _25038_ (.A(_06128_),
    .X(_06355_));
 sg13g2_buf_2 _25039_ (.A(_06355_),
    .X(_06356_));
 sg13g2_buf_2 _25040_ (.A(_06134_),
    .X(_06357_));
 sg13g2_buf_2 _25041_ (.A(_06357_),
    .X(_06358_));
 sg13g2_mux4_1 _25042_ (.S0(net942),
    .A0(\mem.mem_internal.code_mem[148][1] ),
    .A1(\mem.mem_internal.code_mem[149][1] ),
    .A2(\mem.mem_internal.code_mem[150][1] ),
    .A3(\mem.mem_internal.code_mem[151][1] ),
    .S1(net941),
    .X(_06359_));
 sg13g2_buf_2 _25043_ (.A(_06210_),
    .X(_06360_));
 sg13g2_buf_1 _25044_ (.A(_06212_),
    .X(_06361_));
 sg13g2_mux4_1 _25045_ (.S0(net940),
    .A0(_06348_),
    .A1(_06351_),
    .A2(_06354_),
    .A3(_06359_),
    .S1(net939),
    .X(_06362_));
 sg13g2_buf_2 _25046_ (.A(_06237_),
    .X(_06363_));
 sg13g2_mux4_1 _25047_ (.S0(net938),
    .A0(\mem.mem_internal.code_mem[136][1] ),
    .A1(\mem.mem_internal.code_mem[137][1] ),
    .A2(\mem.mem_internal.code_mem[138][1] ),
    .A3(\mem.mem_internal.code_mem[139][1] ),
    .S1(net953),
    .X(_06364_));
 sg13g2_buf_1 _25048_ (.A(_06339_),
    .X(_06365_));
 sg13g2_mux4_1 _25049_ (.S0(_06342_),
    .A0(\mem.mem_internal.code_mem[140][1] ),
    .A1(\mem.mem_internal.code_mem[141][1] ),
    .A2(\mem.mem_internal.code_mem[142][1] ),
    .A3(\mem.mem_internal.code_mem[143][1] ),
    .S1(_06365_),
    .X(_06366_));
 sg13g2_buf_2 _25050_ (.A(_06355_),
    .X(_06367_));
 sg13g2_buf_1 _25051_ (.A(_06357_),
    .X(_06368_));
 sg13g2_mux4_1 _25052_ (.S0(net937),
    .A0(\mem.mem_internal.code_mem[152][1] ),
    .A1(\mem.mem_internal.code_mem[153][1] ),
    .A2(\mem.mem_internal.code_mem[154][1] ),
    .A3(\mem.mem_internal.code_mem[155][1] ),
    .S1(net936),
    .X(_06369_));
 sg13g2_buf_2 _25053_ (.A(_06355_),
    .X(_06370_));
 sg13g2_buf_1 _25054_ (.A(_06183_),
    .X(_06371_));
 sg13g2_mux4_1 _25055_ (.S0(net935),
    .A0(\mem.mem_internal.code_mem[156][1] ),
    .A1(\mem.mem_internal.code_mem[157][1] ),
    .A2(\mem.mem_internal.code_mem[158][1] ),
    .A3(\mem.mem_internal.code_mem[159][1] ),
    .S1(net934),
    .X(_06372_));
 sg13g2_buf_2 _25056_ (.A(_06210_),
    .X(_06373_));
 sg13g2_buf_1 _25057_ (.A(_06212_),
    .X(_06374_));
 sg13g2_mux4_1 _25058_ (.S0(net933),
    .A0(_06364_),
    .A1(_06366_),
    .A2(_06369_),
    .A3(_06372_),
    .S1(net932),
    .X(_06375_));
 sg13g2_buf_1 _25059_ (.A(_06224_),
    .X(_06376_));
 sg13g2_mux4_1 _25060_ (.S0(net1234),
    .A0(_06332_),
    .A1(_06346_),
    .A2(_06362_),
    .A3(_06375_),
    .S1(net1232),
    .X(_06377_));
 sg13g2_buf_2 _25061_ (.A(_06177_),
    .X(_06378_));
 sg13g2_mux4_1 _25062_ (.S0(net931),
    .A0(\mem.mem_internal.code_mem[32][1] ),
    .A1(\mem.mem_internal.code_mem[33][1] ),
    .A2(\mem.mem_internal.code_mem[34][1] ),
    .A3(\mem.mem_internal.code_mem[35][1] ),
    .S1(net812),
    .X(_06379_));
 sg13g2_buf_1 _25063_ (.A(net989),
    .X(_06380_));
 sg13g2_mux4_1 _25064_ (.S0(net811),
    .A0(\mem.mem_internal.code_mem[36][1] ),
    .A1(\mem.mem_internal.code_mem[37][1] ),
    .A2(\mem.mem_internal.code_mem[38][1] ),
    .A3(\mem.mem_internal.code_mem[39][1] ),
    .S1(net806),
    .X(_06381_));
 sg13g2_buf_2 _25065_ (.A(_06237_),
    .X(_06382_));
 sg13g2_buf_1 _25066_ (.A(_06339_),
    .X(_06383_));
 sg13g2_mux4_1 _25067_ (.S0(net930),
    .A0(\mem.mem_internal.code_mem[48][1] ),
    .A1(\mem.mem_internal.code_mem[49][1] ),
    .A2(\mem.mem_internal.code_mem[50][1] ),
    .A3(\mem.mem_internal.code_mem[51][1] ),
    .S1(net805),
    .X(_06384_));
 sg13g2_buf_2 _25068_ (.A(_06172_),
    .X(_06385_));
 sg13g2_buf_1 _25069_ (.A(_06174_),
    .X(_06386_));
 sg13g2_mux4_1 _25070_ (.S0(net929),
    .A0(\mem.mem_internal.code_mem[52][1] ),
    .A1(\mem.mem_internal.code_mem[53][1] ),
    .A2(\mem.mem_internal.code_mem[54][1] ),
    .A3(\mem.mem_internal.code_mem[55][1] ),
    .S1(net804),
    .X(_06387_));
 sg13g2_mux4_1 _25071_ (.S0(net952),
    .A0(_06379_),
    .A1(_06381_),
    .A2(_06384_),
    .A3(_06387_),
    .S1(net947),
    .X(_06388_));
 sg13g2_buf_2 _25072_ (.A(net990),
    .X(_06389_));
 sg13g2_mux4_1 _25073_ (.S0(net803),
    .A0(\mem.mem_internal.code_mem[40][1] ),
    .A1(\mem.mem_internal.code_mem[41][1] ),
    .A2(\mem.mem_internal.code_mem[42][1] ),
    .A3(\mem.mem_internal.code_mem[43][1] ),
    .S1(net819),
    .X(_06390_));
 sg13g2_mux4_1 _25074_ (.S0(net820),
    .A0(\mem.mem_internal.code_mem[44][1] ),
    .A1(\mem.mem_internal.code_mem[45][1] ),
    .A2(\mem.mem_internal.code_mem[46][1] ),
    .A3(\mem.mem_internal.code_mem[47][1] ),
    .S1(net819),
    .X(_06391_));
 sg13g2_buf_2 _25075_ (.A(_06177_),
    .X(_06392_));
 sg13g2_buf_2 _25076_ (.A(_06174_),
    .X(_06393_));
 sg13g2_mux4_1 _25077_ (.S0(net928),
    .A0(\mem.mem_internal.code_mem[56][1] ),
    .A1(\mem.mem_internal.code_mem[57][1] ),
    .A2(\mem.mem_internal.code_mem[58][1] ),
    .A3(\mem.mem_internal.code_mem[59][1] ),
    .S1(net802),
    .X(_06394_));
 sg13g2_buf_2 _25078_ (.A(_06177_),
    .X(_06395_));
 sg13g2_mux4_1 _25079_ (.S0(net927),
    .A0(\mem.mem_internal.code_mem[60][1] ),
    .A1(\mem.mem_internal.code_mem[61][1] ),
    .A2(\mem.mem_internal.code_mem[62][1] ),
    .A3(\mem.mem_internal.code_mem[63][1] ),
    .S1(net815),
    .X(_06396_));
 sg13g2_mux4_1 _25080_ (.S0(net988),
    .A0(_06390_),
    .A1(_06391_),
    .A2(_06394_),
    .A3(_06396_),
    .S1(net987),
    .X(_06397_));
 sg13g2_mux4_1 _25081_ (.S0(_06338_),
    .A0(\mem.mem_internal.code_mem[160][1] ),
    .A1(\mem.mem_internal.code_mem[161][1] ),
    .A2(\mem.mem_internal.code_mem[162][1] ),
    .A3(\mem.mem_internal.code_mem[163][1] ),
    .S1(net809),
    .X(_06398_));
 sg13g2_buf_2 _25082_ (.A(_06177_),
    .X(_06399_));
 sg13g2_buf_1 _25083_ (.A(_06174_),
    .X(_06400_));
 sg13g2_mux4_1 _25084_ (.S0(net926),
    .A0(\mem.mem_internal.code_mem[164][1] ),
    .A1(\mem.mem_internal.code_mem[165][1] ),
    .A2(\mem.mem_internal.code_mem[166][1] ),
    .A3(\mem.mem_internal.code_mem[167][1] ),
    .S1(net801),
    .X(_06401_));
 sg13g2_buf_2 _25085_ (.A(_06355_),
    .X(_06402_));
 sg13g2_buf_1 _25086_ (.A(_06357_),
    .X(_06403_));
 sg13g2_mux4_1 _25087_ (.S0(net925),
    .A0(\mem.mem_internal.code_mem[176][1] ),
    .A1(\mem.mem_internal.code_mem[177][1] ),
    .A2(\mem.mem_internal.code_mem[178][1] ),
    .A3(\mem.mem_internal.code_mem[179][1] ),
    .S1(net924),
    .X(_06404_));
 sg13g2_mux4_1 _25088_ (.S0(net962),
    .A0(\mem.mem_internal.code_mem[180][1] ),
    .A1(\mem.mem_internal.code_mem[181][1] ),
    .A2(\mem.mem_internal.code_mem[182][1] ),
    .A3(\mem.mem_internal.code_mem[183][1] ),
    .S1(net982),
    .X(_06405_));
 sg13g2_buf_2 _25089_ (.A(_06210_),
    .X(_06406_));
 sg13g2_buf_2 _25090_ (.A(_06153_),
    .X(_06407_));
 sg13g2_mux4_1 _25091_ (.S0(net923),
    .A0(_06398_),
    .A1(_06401_),
    .A2(_06404_),
    .A3(_06405_),
    .S1(net922),
    .X(_06408_));
 sg13g2_mux4_1 _25092_ (.S0(net949),
    .A0(\mem.mem_internal.code_mem[168][1] ),
    .A1(\mem.mem_internal.code_mem[169][1] ),
    .A2(\mem.mem_internal.code_mem[170][1] ),
    .A3(\mem.mem_internal.code_mem[171][1] ),
    .S1(net807),
    .X(_06409_));
 sg13g2_buf_2 _25093_ (.A(_06174_),
    .X(_06410_));
 sg13g2_mux4_1 _25094_ (.S0(net984),
    .A0(\mem.mem_internal.code_mem[172][1] ),
    .A1(\mem.mem_internal.code_mem[173][1] ),
    .A2(\mem.mem_internal.code_mem[174][1] ),
    .A3(\mem.mem_internal.code_mem[175][1] ),
    .S1(net800),
    .X(_06411_));
 sg13g2_buf_1 _25095_ (.A(_06183_),
    .X(_06412_));
 sg13g2_mux4_1 _25096_ (.S0(_06254_),
    .A0(\mem.mem_internal.code_mem[184][1] ),
    .A1(\mem.mem_internal.code_mem[185][1] ),
    .A2(\mem.mem_internal.code_mem[186][1] ),
    .A3(\mem.mem_internal.code_mem[187][1] ),
    .S1(net921),
    .X(_06413_));
 sg13g2_mux4_1 _25097_ (.S0(net981),
    .A0(\mem.mem_internal.code_mem[188][1] ),
    .A1(\mem.mem_internal.code_mem[189][1] ),
    .A2(\mem.mem_internal.code_mem[190][1] ),
    .A3(\mem.mem_internal.code_mem[191][1] ),
    .S1(net980),
    .X(_06414_));
 sg13g2_mux4_1 _25098_ (.S0(net979),
    .A0(_06409_),
    .A1(_06411_),
    .A2(_06413_),
    .A3(_06414_),
    .S1(net978),
    .X(_06415_));
 sg13g2_mux4_1 _25099_ (.S0(net1235),
    .A0(_06388_),
    .A1(_06397_),
    .A2(_06408_),
    .A3(_06415_),
    .S1(net1232),
    .X(_06416_));
 sg13g2_buf_2 _25100_ (.A(_06237_),
    .X(_06417_));
 sg13g2_mux4_1 _25101_ (.S0(net920),
    .A0(\mem.mem_internal.code_mem[64][1] ),
    .A1(\mem.mem_internal.code_mem[65][1] ),
    .A2(\mem.mem_internal.code_mem[66][1] ),
    .A3(\mem.mem_internal.code_mem[67][1] ),
    .S1(_06325_),
    .X(_06418_));
 sg13g2_buf_2 _25102_ (.A(_06237_),
    .X(_06419_));
 sg13g2_buf_1 _25103_ (.A(_06339_),
    .X(_06420_));
 sg13g2_mux4_1 _25104_ (.S0(net919),
    .A0(\mem.mem_internal.code_mem[68][1] ),
    .A1(\mem.mem_internal.code_mem[69][1] ),
    .A2(\mem.mem_internal.code_mem[70][1] ),
    .A3(\mem.mem_internal.code_mem[71][1] ),
    .S1(net799),
    .X(_06421_));
 sg13g2_buf_2 _25105_ (.A(_06206_),
    .X(_06422_));
 sg13g2_buf_1 _25106_ (.A(_06203_),
    .X(_06423_));
 sg13g2_mux4_1 _25107_ (.S0(net918),
    .A0(\mem.mem_internal.code_mem[80][1] ),
    .A1(\mem.mem_internal.code_mem[81][1] ),
    .A2(\mem.mem_internal.code_mem[82][1] ),
    .A3(\mem.mem_internal.code_mem[83][1] ),
    .S1(net917),
    .X(_06424_));
 sg13g2_buf_2 _25108_ (.A(_06206_),
    .X(_06425_));
 sg13g2_mux4_1 _25109_ (.S0(net916),
    .A0(\mem.mem_internal.code_mem[84][1] ),
    .A1(\mem.mem_internal.code_mem[85][1] ),
    .A2(\mem.mem_internal.code_mem[86][1] ),
    .A3(\mem.mem_internal.code_mem[87][1] ),
    .S1(net936),
    .X(_06426_));
 sg13g2_buf_1 _25110_ (.A(_06212_),
    .X(_06427_));
 sg13g2_mux4_1 _25111_ (.S0(_06360_),
    .A0(_06418_),
    .A1(_06421_),
    .A2(_06424_),
    .A3(_06426_),
    .S1(net915),
    .X(_06428_));
 sg13g2_mux4_1 _25112_ (.S0(net919),
    .A0(\mem.mem_internal.code_mem[72][1] ),
    .A1(\mem.mem_internal.code_mem[73][1] ),
    .A2(\mem.mem_internal.code_mem[74][1] ),
    .A3(\mem.mem_internal.code_mem[75][1] ),
    .S1(net808),
    .X(_06429_));
 sg13g2_mux4_1 _25113_ (.S0(net985),
    .A0(\mem.mem_internal.code_mem[76][1] ),
    .A1(\mem.mem_internal.code_mem[77][1] ),
    .A2(\mem.mem_internal.code_mem[78][1] ),
    .A3(\mem.mem_internal.code_mem[79][1] ),
    .S1(net816),
    .X(_06430_));
 sg13g2_buf_4 _25114_ (.X(_06431_),
    .A(_06355_));
 sg13g2_mux4_1 _25115_ (.S0(net914),
    .A0(\mem.mem_internal.code_mem[88][1] ),
    .A1(\mem.mem_internal.code_mem[89][1] ),
    .A2(\mem.mem_internal.code_mem[90][1] ),
    .A3(\mem.mem_internal.code_mem[91][1] ),
    .S1(_06403_),
    .X(_06432_));
 sg13g2_buf_2 _25116_ (.A(_06181_),
    .X(_06433_));
 sg13g2_buf_1 _25117_ (.A(_06183_),
    .X(_06434_));
 sg13g2_mux4_1 _25118_ (.S0(net913),
    .A0(\mem.mem_internal.code_mem[92][1] ),
    .A1(\mem.mem_internal.code_mem[93][1] ),
    .A2(\mem.mem_internal.code_mem[94][1] ),
    .A3(\mem.mem_internal.code_mem[95][1] ),
    .S1(net912),
    .X(_06435_));
 sg13g2_buf_2 _25119_ (.A(_06153_),
    .X(_06436_));
 sg13g2_mux4_1 _25120_ (.S0(net933),
    .A0(_06429_),
    .A1(_06430_),
    .A2(_06432_),
    .A3(_06435_),
    .S1(net911),
    .X(_06437_));
 sg13g2_mux4_1 _25121_ (.S0(_06422_),
    .A0(\mem.mem_internal.code_mem[192][1] ),
    .A1(\mem.mem_internal.code_mem[193][1] ),
    .A2(\mem.mem_internal.code_mem[194][1] ),
    .A3(\mem.mem_internal.code_mem[195][1] ),
    .S1(net917),
    .X(_06438_));
 sg13g2_buf_1 _25122_ (.A(_06357_),
    .X(_06439_));
 sg13g2_mux4_1 _25123_ (.S0(net914),
    .A0(\mem.mem_internal.code_mem[196][1] ),
    .A1(\mem.mem_internal.code_mem[197][1] ),
    .A2(\mem.mem_internal.code_mem[198][1] ),
    .A3(\mem.mem_internal.code_mem[199][1] ),
    .S1(net910),
    .X(_06440_));
 sg13g2_buf_1 _25124_ (.A(_06135_),
    .X(_06441_));
 sg13g2_mux4_1 _25125_ (.S0(net959),
    .A0(\mem.mem_internal.code_mem[208][1] ),
    .A1(\mem.mem_internal.code_mem[209][1] ),
    .A2(\mem.mem_internal.code_mem[210][1] ),
    .A3(\mem.mem_internal.code_mem[211][1] ),
    .S1(net909),
    .X(_06442_));
 sg13g2_buf_2 _25126_ (.A(_06129_),
    .X(_06443_));
 sg13g2_buf_1 _25127_ (.A(_06135_),
    .X(_06444_));
 sg13g2_mux4_1 _25128_ (.S0(net908),
    .A0(\mem.mem_internal.code_mem[212][1] ),
    .A1(\mem.mem_internal.code_mem[213][1] ),
    .A2(\mem.mem_internal.code_mem[214][1] ),
    .A3(\mem.mem_internal.code_mem[215][1] ),
    .S1(net907),
    .X(_06445_));
 sg13g2_buf_2 _25129_ (.A(_06148_),
    .X(_06446_));
 sg13g2_mux4_1 _25130_ (.S0(net1231),
    .A0(_06438_),
    .A1(_06440_),
    .A2(_06442_),
    .A3(_06445_),
    .S1(net960),
    .X(_06447_));
 sg13g2_buf_2 _25131_ (.A(_06206_),
    .X(_06448_));
 sg13g2_buf_1 _25132_ (.A(_06357_),
    .X(_06449_));
 sg13g2_mux4_1 _25133_ (.S0(net906),
    .A0(\mem.mem_internal.code_mem[200][1] ),
    .A1(\mem.mem_internal.code_mem[201][1] ),
    .A2(\mem.mem_internal.code_mem[202][1] ),
    .A3(\mem.mem_internal.code_mem[203][1] ),
    .S1(net905),
    .X(_06450_));
 sg13g2_buf_1 _25134_ (.A(_06183_),
    .X(_06451_));
 sg13g2_mux4_1 _25135_ (.S0(net913),
    .A0(\mem.mem_internal.code_mem[204][1] ),
    .A1(\mem.mem_internal.code_mem[205][1] ),
    .A2(\mem.mem_internal.code_mem[206][1] ),
    .A3(\mem.mem_internal.code_mem[207][1] ),
    .S1(net904),
    .X(_06452_));
 sg13g2_buf_2 _25136_ (.A(_06129_),
    .X(_06453_));
 sg13g2_mux4_1 _25137_ (.S0(net903),
    .A0(\mem.mem_internal.code_mem[216][1] ),
    .A1(\mem.mem_internal.code_mem[217][1] ),
    .A2(\mem.mem_internal.code_mem[218][1] ),
    .A3(\mem.mem_internal.code_mem[219][1] ),
    .S1(net909),
    .X(_06454_));
 sg13g2_buf_2 _25138_ (.A(_06129_),
    .X(_06455_));
 sg13g2_buf_1 _25139_ (.A(_06203_),
    .X(_06456_));
 sg13g2_mux4_1 _25140_ (.S0(net902),
    .A0(\mem.mem_internal.code_mem[220][1] ),
    .A1(\mem.mem_internal.code_mem[221][1] ),
    .A2(\mem.mem_internal.code_mem[222][1] ),
    .A3(\mem.mem_internal.code_mem[223][1] ),
    .S1(net901),
    .X(_06457_));
 sg13g2_buf_2 _25141_ (.A(_06148_),
    .X(_06458_));
 sg13g2_buf_1 _25142_ (.A(_06212_),
    .X(_06459_));
 sg13g2_mux4_1 _25143_ (.S0(net1230),
    .A0(_06450_),
    .A1(_06452_),
    .A2(_06454_),
    .A3(_06457_),
    .S1(net900),
    .X(_06460_));
 sg13g2_buf_2 _25144_ (.A(_06168_),
    .X(_06461_));
 sg13g2_buf_1 _25145_ (.A(_06224_),
    .X(_06462_));
 sg13g2_mux4_1 _25146_ (.S0(net1229),
    .A0(_06428_),
    .A1(_06437_),
    .A2(_06447_),
    .A3(_06460_),
    .S1(net1228),
    .X(_06463_));
 sg13g2_buf_1 _25147_ (.A(_06187_),
    .X(_06464_));
 sg13g2_mux4_1 _25148_ (.S0(net954),
    .A0(\mem.mem_internal.code_mem[96][1] ),
    .A1(\mem.mem_internal.code_mem[97][1] ),
    .A2(\mem.mem_internal.code_mem[98][1] ),
    .A3(\mem.mem_internal.code_mem[99][1] ),
    .S1(net899),
    .X(_06465_));
 sg13g2_buf_1 _25149_ (.A(_06339_),
    .X(_06466_));
 sg13g2_mux4_1 _25150_ (.S0(net929),
    .A0(\mem.mem_internal.code_mem[100][1] ),
    .A1(\mem.mem_internal.code_mem[101][1] ),
    .A2(\mem.mem_internal.code_mem[102][1] ),
    .A3(\mem.mem_internal.code_mem[103][1] ),
    .S1(net798),
    .X(_06467_));
 sg13g2_buf_1 _25151_ (.A(_06357_),
    .X(_06468_));
 sg13g2_mux4_1 _25152_ (.S0(_06367_),
    .A0(\mem.mem_internal.code_mem[112][1] ),
    .A1(\mem.mem_internal.code_mem[113][1] ),
    .A2(\mem.mem_internal.code_mem[114][1] ),
    .A3(\mem.mem_internal.code_mem[115][1] ),
    .S1(net898),
    .X(_06469_));
 sg13g2_buf_2 _25153_ (.A(_06355_),
    .X(_06470_));
 sg13g2_mux4_1 _25154_ (.S0(net897),
    .A0(\mem.mem_internal.code_mem[116][1] ),
    .A1(\mem.mem_internal.code_mem[117][1] ),
    .A2(\mem.mem_internal.code_mem[118][1] ),
    .A3(\mem.mem_internal.code_mem[119][1] ),
    .S1(net934),
    .X(_06471_));
 sg13g2_buf_2 _25155_ (.A(_06210_),
    .X(_06472_));
 sg13g2_mux4_1 _25156_ (.S0(net896),
    .A0(_06465_),
    .A1(_06467_),
    .A2(_06469_),
    .A3(_06471_),
    .S1(net939),
    .X(_06473_));
 sg13g2_buf_2 _25157_ (.A(_06172_),
    .X(_06474_));
 sg13g2_buf_1 _25158_ (.A(_06339_),
    .X(_06475_));
 sg13g2_mux4_1 _25159_ (.S0(net895),
    .A0(\mem.mem_internal.code_mem[104][1] ),
    .A1(\mem.mem_internal.code_mem[105][1] ),
    .A2(\mem.mem_internal.code_mem[106][1] ),
    .A3(\mem.mem_internal.code_mem[107][1] ),
    .S1(net797),
    .X(_06476_));
 sg13g2_mux4_1 _25160_ (.S0(net926),
    .A0(\mem.mem_internal.code_mem[108][1] ),
    .A1(\mem.mem_internal.code_mem[109][1] ),
    .A2(\mem.mem_internal.code_mem[110][1] ),
    .A3(\mem.mem_internal.code_mem[111][1] ),
    .S1(_06410_),
    .X(_06477_));
 sg13g2_buf_2 _25161_ (.A(_06181_),
    .X(_06478_));
 sg13g2_mux4_1 _25162_ (.S0(net894),
    .A0(\mem.mem_internal.code_mem[120][1] ),
    .A1(\mem.mem_internal.code_mem[121][1] ),
    .A2(\mem.mem_internal.code_mem[122][1] ),
    .A3(\mem.mem_internal.code_mem[123][1] ),
    .S1(net904),
    .X(_06479_));
 sg13g2_buf_2 _25163_ (.A(_06181_),
    .X(_06480_));
 sg13g2_buf_1 _25164_ (.A(_06183_),
    .X(_06481_));
 sg13g2_mux4_1 _25165_ (.S0(net893),
    .A0(\mem.mem_internal.code_mem[124][1] ),
    .A1(\mem.mem_internal.code_mem[125][1] ),
    .A2(\mem.mem_internal.code_mem[126][1] ),
    .A3(\mem.mem_internal.code_mem[127][1] ),
    .S1(net892),
    .X(_06482_));
 sg13g2_buf_2 _25166_ (.A(_06210_),
    .X(_06483_));
 sg13g2_mux4_1 _25167_ (.S0(net891),
    .A0(_06476_),
    .A1(_06477_),
    .A2(_06479_),
    .A3(_06482_),
    .S1(net922),
    .X(_06484_));
 sg13g2_mux4_1 _25168_ (.S0(net944),
    .A0(\mem.mem_internal.code_mem[224][1] ),
    .A1(\mem.mem_internal.code_mem[225][1] ),
    .A2(\mem.mem_internal.code_mem[226][1] ),
    .A3(\mem.mem_internal.code_mem[227][1] ),
    .S1(_06449_),
    .X(_06485_));
 sg13g2_buf_2 _25169_ (.A(_06355_),
    .X(_06486_));
 sg13g2_buf_1 _25170_ (.A(_06183_),
    .X(_06487_));
 sg13g2_mux4_1 _25171_ (.S0(net890),
    .A0(\mem.mem_internal.code_mem[228][1] ),
    .A1(\mem.mem_internal.code_mem[229][1] ),
    .A2(\mem.mem_internal.code_mem[230][1] ),
    .A3(\mem.mem_internal.code_mem[231][1] ),
    .S1(net889),
    .X(_06488_));
 sg13g2_buf_1 _25172_ (.A(_06135_),
    .X(_06489_));
 sg13g2_mux4_1 _25173_ (.S0(net908),
    .A0(\mem.mem_internal.code_mem[240][1] ),
    .A1(\mem.mem_internal.code_mem[241][1] ),
    .A2(\mem.mem_internal.code_mem[242][1] ),
    .A3(\mem.mem_internal.code_mem[243][1] ),
    .S1(net888),
    .X(_06490_));
 sg13g2_mux4_1 _25174_ (.S0(net975),
    .A0(\mem.mem_internal.code_mem[244][1] ),
    .A1(\mem.mem_internal.code_mem[245][1] ),
    .A2(\mem.mem_internal.code_mem[246][1] ),
    .A3(\mem.mem_internal.code_mem[247][1] ),
    .S1(net974),
    .X(_06491_));
 sg13g2_buf_1 _25175_ (.A(_06212_),
    .X(_06492_));
 sg13g2_mux4_1 _25176_ (.S0(_06458_),
    .A0(_06485_),
    .A1(_06488_),
    .A2(_06490_),
    .A3(_06491_),
    .S1(net887),
    .X(_06493_));
 sg13g2_buf_1 _25177_ (.A(_06357_),
    .X(_06494_));
 sg13g2_mux4_1 _25178_ (.S0(net897),
    .A0(\mem.mem_internal.code_mem[232][1] ),
    .A1(\mem.mem_internal.code_mem[233][1] ),
    .A2(\mem.mem_internal.code_mem[234][1] ),
    .A3(\mem.mem_internal.code_mem[235][1] ),
    .S1(net886),
    .X(_06495_));
 sg13g2_mux4_1 _25179_ (.S0(net983),
    .A0(\mem.mem_internal.code_mem[236][1] ),
    .A1(\mem.mem_internal.code_mem[237][1] ),
    .A2(\mem.mem_internal.code_mem[238][1] ),
    .A3(\mem.mem_internal.code_mem[239][1] ),
    .S1(_06481_),
    .X(_06496_));
 sg13g2_buf_2 _25180_ (.A(_06129_),
    .X(_06497_));
 sg13g2_mux4_1 _25181_ (.S0(net885),
    .A0(\mem.mem_internal.code_mem[248][1] ),
    .A1(\mem.mem_internal.code_mem[249][1] ),
    .A2(\mem.mem_internal.code_mem[250][1] ),
    .A3(\mem.mem_internal.code_mem[251][1] ),
    .S1(net907),
    .X(_06498_));
 sg13g2_mux4_1 _25182_ (.S0(_06207_),
    .A0(\mem.mem_internal.code_mem[252][1] ),
    .A1(\mem.mem_internal.code_mem[253][1] ),
    .A2(\mem.mem_internal.code_mem[254][1] ),
    .A3(\mem.mem_internal.code_mem[255][1] ),
    .S1(net972),
    .X(_06499_));
 sg13g2_mux4_1 _25183_ (.S0(net971),
    .A0(_06495_),
    .A1(_06496_),
    .A2(_06498_),
    .A3(_06499_),
    .S1(net970),
    .X(_06500_));
 sg13g2_mux4_1 _25184_ (.S0(net1234),
    .A0(_06473_),
    .A1(_06484_),
    .A2(_06493_),
    .A3(_06500_),
    .S1(net1233),
    .X(_06501_));
 sg13g2_mux4_1 _25185_ (.S0(_06300_),
    .A0(_06377_),
    .A1(_06416_),
    .A2(_06463_),
    .A3(_06501_),
    .S1(_06301_),
    .X(_06502_));
 sg13g2_nor2_1 _25186_ (.A(_06304_),
    .B(_06502_),
    .Y(_06503_));
 sg13g2_a21oi_1 _25187_ (.A1(net832),
    .A2(_06318_),
    .Y(_06504_),
    .B1(_06503_));
 sg13g2_nand2_1 _25188_ (.Y(_06505_),
    .A(\mem.internal_data_out[1] ),
    .B(net546));
 sg13g2_o21ai_1 _25189_ (.B1(_06505_),
    .Y(_02421_),
    .A1(net546),
    .A2(_06504_));
 sg13g2_mux4_1 _25190_ (.S0(net538),
    .A0(\mem.mem_internal.data_mem[0][2] ),
    .A1(\mem.mem_internal.data_mem[1][2] ),
    .A2(\mem.mem_internal.data_mem[2][2] ),
    .A3(\mem.mem_internal.data_mem[3][2] ),
    .S1(net537),
    .X(_06506_));
 sg13g2_mux4_1 _25191_ (.S0(net545),
    .A0(\mem.mem_internal.data_mem[4][2] ),
    .A1(\mem.mem_internal.data_mem[5][2] ),
    .A2(\mem.mem_internal.data_mem[6][2] ),
    .A3(\mem.mem_internal.data_mem[7][2] ),
    .S1(net544),
    .X(_06507_));
 sg13g2_mux4_1 _25192_ (.S0(net577),
    .A0(\mem.mem_internal.data_mem[8][2] ),
    .A1(\mem.mem_internal.data_mem[9][2] ),
    .A2(\mem.mem_internal.data_mem[10][2] ),
    .A3(\mem.mem_internal.data_mem[11][2] ),
    .S1(net543),
    .X(_06508_));
 sg13g2_mux4_1 _25193_ (.S0(net542),
    .A0(\mem.mem_internal.data_mem[12][2] ),
    .A1(\mem.mem_internal.data_mem[13][2] ),
    .A2(\mem.mem_internal.data_mem[14][2] ),
    .A3(\mem.mem_internal.data_mem[15][2] ),
    .S1(net541),
    .X(_06509_));
 sg13g2_mux4_1 _25194_ (.S0(_06151_),
    .A0(_06506_),
    .A1(_06507_),
    .A2(_06508_),
    .A3(_06509_),
    .S1(net986),
    .X(_06510_));
 sg13g2_mux4_1 _25195_ (.S0(_06157_),
    .A0(\mem.mem_internal.data_mem[16][2] ),
    .A1(\mem.mem_internal.data_mem[17][2] ),
    .A2(\mem.mem_internal.data_mem[18][2] ),
    .A3(\mem.mem_internal.data_mem[19][2] ),
    .S1(_06158_),
    .X(_06511_));
 sg13g2_mux4_1 _25196_ (.S0(net538),
    .A0(\mem.mem_internal.data_mem[20][2] ),
    .A1(\mem.mem_internal.data_mem[21][2] ),
    .A2(\mem.mem_internal.data_mem[22][2] ),
    .A3(\mem.mem_internal.data_mem[23][2] ),
    .S1(net537),
    .X(_06512_));
 sg13g2_mux4_1 _25197_ (.S0(net576),
    .A0(\mem.mem_internal.data_mem[24][2] ),
    .A1(\mem.mem_internal.data_mem[25][2] ),
    .A2(\mem.mem_internal.data_mem[26][2] ),
    .A3(\mem.mem_internal.data_mem[27][2] ),
    .S1(net575),
    .X(_06513_));
 sg13g2_mux4_1 _25198_ (.S0(_06163_),
    .A0(\mem.mem_internal.data_mem[28][2] ),
    .A1(\mem.mem_internal.data_mem[29][2] ),
    .A2(\mem.mem_internal.data_mem[30][2] ),
    .A3(\mem.mem_internal.data_mem[31][2] ),
    .S1(_06164_),
    .X(_06514_));
 sg13g2_mux4_1 _25199_ (.S0(net988),
    .A0(_06511_),
    .A1(_06512_),
    .A2(_06513_),
    .A3(_06514_),
    .S1(net986),
    .X(_06515_));
 sg13g2_mux2_1 _25200_ (.A0(_06510_),
    .A1(_06515_),
    .S(net817),
    .X(_06516_));
 sg13g2_mux4_1 _25201_ (.S0(net958),
    .A0(\mem.mem_internal.code_mem[0][2] ),
    .A1(\mem.mem_internal.code_mem[1][2] ),
    .A2(\mem.mem_internal.code_mem[2][2] ),
    .A3(\mem.mem_internal.code_mem[3][2] ),
    .S1(net814),
    .X(_06517_));
 sg13g2_mux4_1 _25202_ (.S0(net957),
    .A0(\mem.mem_internal.code_mem[4][2] ),
    .A1(\mem.mem_internal.code_mem[5][2] ),
    .A2(\mem.mem_internal.code_mem[6][2] ),
    .A3(\mem.mem_internal.code_mem[7][2] ),
    .S1(net813),
    .X(_06518_));
 sg13g2_mux4_1 _25203_ (.S0(net956),
    .A0(\mem.mem_internal.code_mem[16][2] ),
    .A1(\mem.mem_internal.code_mem[17][2] ),
    .A2(\mem.mem_internal.code_mem[18][2] ),
    .A3(\mem.mem_internal.code_mem[19][2] ),
    .S1(net955),
    .X(_06519_));
 sg13g2_mux4_1 _25204_ (.S0(net954),
    .A0(\mem.mem_internal.code_mem[20][2] ),
    .A1(\mem.mem_internal.code_mem[21][2] ),
    .A2(\mem.mem_internal.code_mem[22][2] ),
    .A3(\mem.mem_internal.code_mem[23][2] ),
    .S1(net953),
    .X(_06520_));
 sg13g2_mux4_1 _25205_ (.S0(_06330_),
    .A0(_06517_),
    .A1(_06518_),
    .A2(_06519_),
    .A3(_06520_),
    .S1(net951),
    .X(_06521_));
 sg13g2_mux4_1 _25206_ (.S0(net957),
    .A0(\mem.mem_internal.code_mem[8][2] ),
    .A1(\mem.mem_internal.code_mem[9][2] ),
    .A2(\mem.mem_internal.code_mem[10][2] ),
    .A3(\mem.mem_internal.code_mem[11][2] ),
    .S1(net812),
    .X(_06522_));
 sg13g2_mux4_1 _25207_ (.S0(net811),
    .A0(\mem.mem_internal.code_mem[12][2] ),
    .A1(\mem.mem_internal.code_mem[13][2] ),
    .A2(\mem.mem_internal.code_mem[14][2] ),
    .A3(\mem.mem_internal.code_mem[15][2] ),
    .S1(net810),
    .X(_06523_));
 sg13g2_mux4_1 _25208_ (.S0(net950),
    .A0(\mem.mem_internal.code_mem[24][2] ),
    .A1(\mem.mem_internal.code_mem[25][2] ),
    .A2(\mem.mem_internal.code_mem[26][2] ),
    .A3(\mem.mem_internal.code_mem[27][2] ),
    .S1(net809),
    .X(_06524_));
 sg13g2_buf_2 _25209_ (.A(_06172_),
    .X(_06525_));
 sg13g2_mux4_1 _25210_ (.S0(net884),
    .A0(\mem.mem_internal.code_mem[28][2] ),
    .A1(\mem.mem_internal.code_mem[29][2] ),
    .A2(\mem.mem_internal.code_mem[30][2] ),
    .A3(\mem.mem_internal.code_mem[31][2] ),
    .S1(net816),
    .X(_06526_));
 sg13g2_mux4_1 _25211_ (.S0(net948),
    .A0(_06522_),
    .A1(_06523_),
    .A2(_06524_),
    .A3(_06526_),
    .S1(_06345_),
    .X(_06527_));
 sg13g2_mux4_1 _25212_ (.S0(_06324_),
    .A0(\mem.mem_internal.code_mem[128][2] ),
    .A1(\mem.mem_internal.code_mem[129][2] ),
    .A2(\mem.mem_internal.code_mem[130][2] ),
    .A3(\mem.mem_internal.code_mem[131][2] ),
    .S1(net946),
    .X(_06528_));
 sg13g2_mux4_1 _25213_ (.S0(net945),
    .A0(\mem.mem_internal.code_mem[132][2] ),
    .A1(\mem.mem_internal.code_mem[133][2] ),
    .A2(\mem.mem_internal.code_mem[134][2] ),
    .A3(\mem.mem_internal.code_mem[135][2] ),
    .S1(net808),
    .X(_06529_));
 sg13g2_mux4_1 _25214_ (.S0(net944),
    .A0(\mem.mem_internal.code_mem[144][2] ),
    .A1(\mem.mem_internal.code_mem[145][2] ),
    .A2(\mem.mem_internal.code_mem[146][2] ),
    .A3(\mem.mem_internal.code_mem[147][2] ),
    .S1(net943),
    .X(_06530_));
 sg13g2_mux4_1 _25215_ (.S0(net942),
    .A0(\mem.mem_internal.code_mem[148][2] ),
    .A1(\mem.mem_internal.code_mem[149][2] ),
    .A2(\mem.mem_internal.code_mem[150][2] ),
    .A3(\mem.mem_internal.code_mem[151][2] ),
    .S1(net941),
    .X(_06531_));
 sg13g2_mux4_1 _25216_ (.S0(net940),
    .A0(_06528_),
    .A1(_06529_),
    .A2(_06530_),
    .A3(_06531_),
    .S1(net939),
    .X(_06532_));
 sg13g2_mux4_1 _25217_ (.S0(net938),
    .A0(\mem.mem_internal.code_mem[136][2] ),
    .A1(\mem.mem_internal.code_mem[137][2] ),
    .A2(\mem.mem_internal.code_mem[138][2] ),
    .A3(\mem.mem_internal.code_mem[139][2] ),
    .S1(net899),
    .X(_06533_));
 sg13g2_mux4_1 _25218_ (.S0(_06342_),
    .A0(\mem.mem_internal.code_mem[140][2] ),
    .A1(\mem.mem_internal.code_mem[141][2] ),
    .A2(\mem.mem_internal.code_mem[142][2] ),
    .A3(\mem.mem_internal.code_mem[143][2] ),
    .S1(net797),
    .X(_06534_));
 sg13g2_mux4_1 _25219_ (.S0(net937),
    .A0(\mem.mem_internal.code_mem[152][2] ),
    .A1(\mem.mem_internal.code_mem[153][2] ),
    .A2(\mem.mem_internal.code_mem[154][2] ),
    .A3(\mem.mem_internal.code_mem[155][2] ),
    .S1(net936),
    .X(_06535_));
 sg13g2_mux4_1 _25220_ (.S0(net935),
    .A0(\mem.mem_internal.code_mem[156][2] ),
    .A1(\mem.mem_internal.code_mem[157][2] ),
    .A2(\mem.mem_internal.code_mem[158][2] ),
    .A3(\mem.mem_internal.code_mem[159][2] ),
    .S1(net934),
    .X(_06536_));
 sg13g2_mux4_1 _25221_ (.S0(net933),
    .A0(_06533_),
    .A1(_06534_),
    .A2(_06535_),
    .A3(_06536_),
    .S1(net932),
    .X(_06537_));
 sg13g2_mux4_1 _25222_ (.S0(net1234),
    .A0(_06521_),
    .A1(_06527_),
    .A2(_06532_),
    .A3(_06537_),
    .S1(_06376_),
    .X(_06538_));
 sg13g2_mux4_1 _25223_ (.S0(net931),
    .A0(\mem.mem_internal.code_mem[32][2] ),
    .A1(\mem.mem_internal.code_mem[33][2] ),
    .A2(\mem.mem_internal.code_mem[34][2] ),
    .A3(\mem.mem_internal.code_mem[35][2] ),
    .S1(net812),
    .X(_06539_));
 sg13g2_mux4_1 _25224_ (.S0(net811),
    .A0(\mem.mem_internal.code_mem[36][2] ),
    .A1(\mem.mem_internal.code_mem[37][2] ),
    .A2(\mem.mem_internal.code_mem[38][2] ),
    .A3(\mem.mem_internal.code_mem[39][2] ),
    .S1(net806),
    .X(_06540_));
 sg13g2_mux4_1 _25225_ (.S0(net930),
    .A0(\mem.mem_internal.code_mem[48][2] ),
    .A1(\mem.mem_internal.code_mem[49][2] ),
    .A2(\mem.mem_internal.code_mem[50][2] ),
    .A3(\mem.mem_internal.code_mem[51][2] ),
    .S1(net805),
    .X(_06541_));
 sg13g2_mux4_1 _25226_ (.S0(net929),
    .A0(\mem.mem_internal.code_mem[52][2] ),
    .A1(\mem.mem_internal.code_mem[53][2] ),
    .A2(\mem.mem_internal.code_mem[54][2] ),
    .A3(\mem.mem_internal.code_mem[55][2] ),
    .S1(net804),
    .X(_06542_));
 sg13g2_mux4_1 _25227_ (.S0(net952),
    .A0(_06539_),
    .A1(_06540_),
    .A2(_06541_),
    .A3(_06542_),
    .S1(net947),
    .X(_06543_));
 sg13g2_mux4_1 _25228_ (.S0(net803),
    .A0(\mem.mem_internal.code_mem[40][2] ),
    .A1(\mem.mem_internal.code_mem[41][2] ),
    .A2(\mem.mem_internal.code_mem[42][2] ),
    .A3(\mem.mem_internal.code_mem[43][2] ),
    .S1(net810),
    .X(_06544_));
 sg13g2_mux4_1 _25229_ (.S0(net820),
    .A0(\mem.mem_internal.code_mem[44][2] ),
    .A1(\mem.mem_internal.code_mem[45][2] ),
    .A2(\mem.mem_internal.code_mem[46][2] ),
    .A3(\mem.mem_internal.code_mem[47][2] ),
    .S1(net819),
    .X(_06545_));
 sg13g2_mux4_1 _25230_ (.S0(net928),
    .A0(\mem.mem_internal.code_mem[56][2] ),
    .A1(\mem.mem_internal.code_mem[57][2] ),
    .A2(\mem.mem_internal.code_mem[58][2] ),
    .A3(\mem.mem_internal.code_mem[59][2] ),
    .S1(net802),
    .X(_06546_));
 sg13g2_mux4_1 _25231_ (.S0(net927),
    .A0(\mem.mem_internal.code_mem[60][2] ),
    .A1(\mem.mem_internal.code_mem[61][2] ),
    .A2(\mem.mem_internal.code_mem[62][2] ),
    .A3(\mem.mem_internal.code_mem[63][2] ),
    .S1(net815),
    .X(_06547_));
 sg13g2_mux4_1 _25232_ (.S0(_06150_),
    .A0(_06544_),
    .A1(_06545_),
    .A2(_06546_),
    .A3(_06547_),
    .S1(net987),
    .X(_06548_));
 sg13g2_mux4_1 _25233_ (.S0(net945),
    .A0(\mem.mem_internal.code_mem[160][2] ),
    .A1(\mem.mem_internal.code_mem[161][2] ),
    .A2(\mem.mem_internal.code_mem[162][2] ),
    .A3(\mem.mem_internal.code_mem[163][2] ),
    .S1(net809),
    .X(_06549_));
 sg13g2_mux4_1 _25234_ (.S0(net926),
    .A0(\mem.mem_internal.code_mem[164][2] ),
    .A1(\mem.mem_internal.code_mem[165][2] ),
    .A2(\mem.mem_internal.code_mem[166][2] ),
    .A3(\mem.mem_internal.code_mem[167][2] ),
    .S1(net801),
    .X(_06550_));
 sg13g2_mux4_1 _25235_ (.S0(net925),
    .A0(\mem.mem_internal.code_mem[176][2] ),
    .A1(\mem.mem_internal.code_mem[177][2] ),
    .A2(\mem.mem_internal.code_mem[178][2] ),
    .A3(\mem.mem_internal.code_mem[179][2] ),
    .S1(net924),
    .X(_06551_));
 sg13g2_mux4_1 _25236_ (.S0(net962),
    .A0(\mem.mem_internal.code_mem[180][2] ),
    .A1(\mem.mem_internal.code_mem[181][2] ),
    .A2(\mem.mem_internal.code_mem[182][2] ),
    .A3(\mem.mem_internal.code_mem[183][2] ),
    .S1(net912),
    .X(_06552_));
 sg13g2_mux4_1 _25237_ (.S0(net923),
    .A0(_06549_),
    .A1(_06550_),
    .A2(_06551_),
    .A3(_06552_),
    .S1(net911),
    .X(_06553_));
 sg13g2_mux4_1 _25238_ (.S0(net949),
    .A0(\mem.mem_internal.code_mem[168][2] ),
    .A1(\mem.mem_internal.code_mem[169][2] ),
    .A2(\mem.mem_internal.code_mem[170][2] ),
    .A3(\mem.mem_internal.code_mem[171][2] ),
    .S1(net807),
    .X(_06554_));
 sg13g2_mux4_1 _25239_ (.S0(net984),
    .A0(\mem.mem_internal.code_mem[172][2] ),
    .A1(\mem.mem_internal.code_mem[173][2] ),
    .A2(\mem.mem_internal.code_mem[174][2] ),
    .A3(\mem.mem_internal.code_mem[175][2] ),
    .S1(net800),
    .X(_06555_));
 sg13g2_mux4_1 _25240_ (.S0(net962),
    .A0(\mem.mem_internal.code_mem[184][2] ),
    .A1(\mem.mem_internal.code_mem[185][2] ),
    .A2(\mem.mem_internal.code_mem[186][2] ),
    .A3(\mem.mem_internal.code_mem[187][2] ),
    .S1(net921),
    .X(_06556_));
 sg13g2_mux4_1 _25241_ (.S0(net981),
    .A0(\mem.mem_internal.code_mem[188][2] ),
    .A1(\mem.mem_internal.code_mem[189][2] ),
    .A2(\mem.mem_internal.code_mem[190][2] ),
    .A3(\mem.mem_internal.code_mem[191][2] ),
    .S1(net980),
    .X(_06557_));
 sg13g2_mux4_1 _25242_ (.S0(net891),
    .A0(_06554_),
    .A1(_06555_),
    .A2(_06556_),
    .A3(_06557_),
    .S1(net978),
    .X(_06558_));
 sg13g2_mux4_1 _25243_ (.S0(net1235),
    .A0(_06543_),
    .A1(_06548_),
    .A2(_06553_),
    .A3(_06558_),
    .S1(net1232),
    .X(_06559_));
 sg13g2_mux4_1 _25244_ (.S0(net965),
    .A0(\mem.mem_internal.code_mem[64][2] ),
    .A1(\mem.mem_internal.code_mem[65][2] ),
    .A2(\mem.mem_internal.code_mem[66][2] ),
    .A3(\mem.mem_internal.code_mem[67][2] ),
    .S1(_06325_),
    .X(_06560_));
 sg13g2_mux4_1 _25245_ (.S0(net919),
    .A0(\mem.mem_internal.code_mem[68][2] ),
    .A1(\mem.mem_internal.code_mem[69][2] ),
    .A2(\mem.mem_internal.code_mem[70][2] ),
    .A3(\mem.mem_internal.code_mem[71][2] ),
    .S1(net799),
    .X(_06561_));
 sg13g2_mux4_1 _25246_ (.S0(net918),
    .A0(\mem.mem_internal.code_mem[80][2] ),
    .A1(\mem.mem_internal.code_mem[81][2] ),
    .A2(\mem.mem_internal.code_mem[82][2] ),
    .A3(\mem.mem_internal.code_mem[83][2] ),
    .S1(net964),
    .X(_06562_));
 sg13g2_mux4_1 _25247_ (.S0(net916),
    .A0(\mem.mem_internal.code_mem[84][2] ),
    .A1(\mem.mem_internal.code_mem[85][2] ),
    .A2(\mem.mem_internal.code_mem[86][2] ),
    .A3(\mem.mem_internal.code_mem[87][2] ),
    .S1(net936),
    .X(_06563_));
 sg13g2_mux4_1 _25248_ (.S0(net940),
    .A0(_06560_),
    .A1(_06561_),
    .A2(_06562_),
    .A3(_06563_),
    .S1(net915),
    .X(_06564_));
 sg13g2_mux4_1 _25249_ (.S0(net919),
    .A0(\mem.mem_internal.code_mem[72][2] ),
    .A1(\mem.mem_internal.code_mem[73][2] ),
    .A2(\mem.mem_internal.code_mem[74][2] ),
    .A3(\mem.mem_internal.code_mem[75][2] ),
    .S1(_06350_),
    .X(_06565_));
 sg13g2_mux4_1 _25250_ (.S0(net985),
    .A0(\mem.mem_internal.code_mem[76][2] ),
    .A1(\mem.mem_internal.code_mem[77][2] ),
    .A2(\mem.mem_internal.code_mem[78][2] ),
    .A3(\mem.mem_internal.code_mem[79][2] ),
    .S1(net816),
    .X(_06566_));
 sg13g2_mux4_1 _25251_ (.S0(net914),
    .A0(\mem.mem_internal.code_mem[88][2] ),
    .A1(\mem.mem_internal.code_mem[89][2] ),
    .A2(\mem.mem_internal.code_mem[90][2] ),
    .A3(\mem.mem_internal.code_mem[91][2] ),
    .S1(net910),
    .X(_06567_));
 sg13g2_mux4_1 _25252_ (.S0(net913),
    .A0(\mem.mem_internal.code_mem[92][2] ),
    .A1(\mem.mem_internal.code_mem[93][2] ),
    .A2(\mem.mem_internal.code_mem[94][2] ),
    .A3(\mem.mem_internal.code_mem[95][2] ),
    .S1(net912),
    .X(_06568_));
 sg13g2_mux4_1 _25253_ (.S0(net933),
    .A0(_06565_),
    .A1(_06566_),
    .A2(_06567_),
    .A3(_06568_),
    .S1(net911),
    .X(_06569_));
 sg13g2_mux4_1 _25254_ (.S0(net918),
    .A0(\mem.mem_internal.code_mem[192][2] ),
    .A1(\mem.mem_internal.code_mem[193][2] ),
    .A2(\mem.mem_internal.code_mem[194][2] ),
    .A3(\mem.mem_internal.code_mem[195][2] ),
    .S1(net917),
    .X(_06570_));
 sg13g2_mux4_1 _25255_ (.S0(_06431_),
    .A0(\mem.mem_internal.code_mem[196][2] ),
    .A1(\mem.mem_internal.code_mem[197][2] ),
    .A2(\mem.mem_internal.code_mem[198][2] ),
    .A3(\mem.mem_internal.code_mem[199][2] ),
    .S1(net910),
    .X(_06571_));
 sg13g2_mux4_1 _25256_ (.S0(net959),
    .A0(\mem.mem_internal.code_mem[208][2] ),
    .A1(\mem.mem_internal.code_mem[209][2] ),
    .A2(\mem.mem_internal.code_mem[210][2] ),
    .A3(\mem.mem_internal.code_mem[211][2] ),
    .S1(net961),
    .X(_06572_));
 sg13g2_mux4_1 _25257_ (.S0(net908),
    .A0(\mem.mem_internal.code_mem[212][2] ),
    .A1(\mem.mem_internal.code_mem[213][2] ),
    .A2(\mem.mem_internal.code_mem[214][2] ),
    .A3(\mem.mem_internal.code_mem[215][2] ),
    .S1(_06444_),
    .X(_06573_));
 sg13g2_mux4_1 _25258_ (.S0(net1231),
    .A0(_06570_),
    .A1(_06571_),
    .A2(_06572_),
    .A3(_06573_),
    .S1(net960),
    .X(_06574_));
 sg13g2_mux4_1 _25259_ (.S0(net906),
    .A0(\mem.mem_internal.code_mem[200][2] ),
    .A1(\mem.mem_internal.code_mem[201][2] ),
    .A2(\mem.mem_internal.code_mem[202][2] ),
    .A3(\mem.mem_internal.code_mem[203][2] ),
    .S1(net905),
    .X(_06575_));
 sg13g2_mux4_1 _25260_ (.S0(net913),
    .A0(\mem.mem_internal.code_mem[204][2] ),
    .A1(\mem.mem_internal.code_mem[205][2] ),
    .A2(\mem.mem_internal.code_mem[206][2] ),
    .A3(\mem.mem_internal.code_mem[207][2] ),
    .S1(_06451_),
    .X(_06576_));
 sg13g2_mux4_1 _25261_ (.S0(net903),
    .A0(\mem.mem_internal.code_mem[216][2] ),
    .A1(\mem.mem_internal.code_mem[217][2] ),
    .A2(\mem.mem_internal.code_mem[218][2] ),
    .A3(\mem.mem_internal.code_mem[219][2] ),
    .S1(net909),
    .X(_06577_));
 sg13g2_mux4_1 _25262_ (.S0(net902),
    .A0(\mem.mem_internal.code_mem[220][2] ),
    .A1(\mem.mem_internal.code_mem[221][2] ),
    .A2(\mem.mem_internal.code_mem[222][2] ),
    .A3(\mem.mem_internal.code_mem[223][2] ),
    .S1(net901),
    .X(_06578_));
 sg13g2_mux4_1 _25263_ (.S0(net1230),
    .A0(_06575_),
    .A1(_06576_),
    .A2(_06577_),
    .A3(_06578_),
    .S1(net900),
    .X(_06579_));
 sg13g2_mux4_1 _25264_ (.S0(net1229),
    .A0(_06564_),
    .A1(_06569_),
    .A2(_06574_),
    .A3(_06579_),
    .S1(net1228),
    .X(_06580_));
 sg13g2_mux4_1 _25265_ (.S0(net954),
    .A0(\mem.mem_internal.code_mem[96][2] ),
    .A1(\mem.mem_internal.code_mem[97][2] ),
    .A2(\mem.mem_internal.code_mem[98][2] ),
    .A3(\mem.mem_internal.code_mem[99][2] ),
    .S1(net899),
    .X(_06581_));
 sg13g2_mux4_1 _25266_ (.S0(_06385_),
    .A0(\mem.mem_internal.code_mem[100][2] ),
    .A1(\mem.mem_internal.code_mem[101][2] ),
    .A2(\mem.mem_internal.code_mem[102][2] ),
    .A3(\mem.mem_internal.code_mem[103][2] ),
    .S1(net798),
    .X(_06582_));
 sg13g2_mux4_1 _25267_ (.S0(net906),
    .A0(\mem.mem_internal.code_mem[112][2] ),
    .A1(\mem.mem_internal.code_mem[113][2] ),
    .A2(\mem.mem_internal.code_mem[114][2] ),
    .A3(\mem.mem_internal.code_mem[115][2] ),
    .S1(net898),
    .X(_06583_));
 sg13g2_mux4_1 _25268_ (.S0(net897),
    .A0(\mem.mem_internal.code_mem[116][2] ),
    .A1(\mem.mem_internal.code_mem[117][2] ),
    .A2(\mem.mem_internal.code_mem[118][2] ),
    .A3(\mem.mem_internal.code_mem[119][2] ),
    .S1(_06371_),
    .X(_06584_));
 sg13g2_mux4_1 _25269_ (.S0(net896),
    .A0(_06581_),
    .A1(_06582_),
    .A2(_06583_),
    .A3(_06584_),
    .S1(net939),
    .X(_06585_));
 sg13g2_mux4_1 _25270_ (.S0(net895),
    .A0(\mem.mem_internal.code_mem[104][2] ),
    .A1(\mem.mem_internal.code_mem[105][2] ),
    .A2(\mem.mem_internal.code_mem[106][2] ),
    .A3(\mem.mem_internal.code_mem[107][2] ),
    .S1(net797),
    .X(_06586_));
 sg13g2_mux4_1 _25271_ (.S0(net926),
    .A0(\mem.mem_internal.code_mem[108][2] ),
    .A1(\mem.mem_internal.code_mem[109][2] ),
    .A2(\mem.mem_internal.code_mem[110][2] ),
    .A3(\mem.mem_internal.code_mem[111][2] ),
    .S1(net802),
    .X(_06587_));
 sg13g2_mux4_1 _25272_ (.S0(net894),
    .A0(\mem.mem_internal.code_mem[120][2] ),
    .A1(\mem.mem_internal.code_mem[121][2] ),
    .A2(\mem.mem_internal.code_mem[122][2] ),
    .A3(\mem.mem_internal.code_mem[123][2] ),
    .S1(net904),
    .X(_06588_));
 sg13g2_mux4_1 _25273_ (.S0(net893),
    .A0(\mem.mem_internal.code_mem[124][2] ),
    .A1(\mem.mem_internal.code_mem[125][2] ),
    .A2(\mem.mem_internal.code_mem[126][2] ),
    .A3(\mem.mem_internal.code_mem[127][2] ),
    .S1(net892),
    .X(_06589_));
 sg13g2_mux4_1 _25274_ (.S0(net891),
    .A0(_06586_),
    .A1(_06587_),
    .A2(_06588_),
    .A3(_06589_),
    .S1(net922),
    .X(_06590_));
 sg13g2_mux4_1 _25275_ (.S0(net944),
    .A0(\mem.mem_internal.code_mem[224][2] ),
    .A1(\mem.mem_internal.code_mem[225][2] ),
    .A2(\mem.mem_internal.code_mem[226][2] ),
    .A3(\mem.mem_internal.code_mem[227][2] ),
    .S1(_06449_),
    .X(_06591_));
 sg13g2_mux4_1 _25276_ (.S0(net890),
    .A0(\mem.mem_internal.code_mem[228][2] ),
    .A1(\mem.mem_internal.code_mem[229][2] ),
    .A2(\mem.mem_internal.code_mem[230][2] ),
    .A3(\mem.mem_internal.code_mem[231][2] ),
    .S1(net889),
    .X(_06592_));
 sg13g2_mux4_1 _25277_ (.S0(net908),
    .A0(\mem.mem_internal.code_mem[240][2] ),
    .A1(\mem.mem_internal.code_mem[241][2] ),
    .A2(\mem.mem_internal.code_mem[242][2] ),
    .A3(\mem.mem_internal.code_mem[243][2] ),
    .S1(net888),
    .X(_06593_));
 sg13g2_mux4_1 _25278_ (.S0(net902),
    .A0(\mem.mem_internal.code_mem[244][2] ),
    .A1(\mem.mem_internal.code_mem[245][2] ),
    .A2(\mem.mem_internal.code_mem[246][2] ),
    .A3(\mem.mem_internal.code_mem[247][2] ),
    .S1(net974),
    .X(_06594_));
 sg13g2_mux4_1 _25279_ (.S0(net1230),
    .A0(_06591_),
    .A1(_06592_),
    .A2(_06593_),
    .A3(_06594_),
    .S1(net887),
    .X(_06595_));
 sg13g2_mux4_1 _25280_ (.S0(_06470_),
    .A0(\mem.mem_internal.code_mem[232][2] ),
    .A1(\mem.mem_internal.code_mem[233][2] ),
    .A2(\mem.mem_internal.code_mem[234][2] ),
    .A3(\mem.mem_internal.code_mem[235][2] ),
    .S1(net886),
    .X(_06596_));
 sg13g2_mux4_1 _25281_ (.S0(net983),
    .A0(\mem.mem_internal.code_mem[236][2] ),
    .A1(\mem.mem_internal.code_mem[237][2] ),
    .A2(\mem.mem_internal.code_mem[238][2] ),
    .A3(\mem.mem_internal.code_mem[239][2] ),
    .S1(net982),
    .X(_06597_));
 sg13g2_mux4_1 _25282_ (.S0(net885),
    .A0(\mem.mem_internal.code_mem[248][2] ),
    .A1(\mem.mem_internal.code_mem[249][2] ),
    .A2(\mem.mem_internal.code_mem[250][2] ),
    .A3(\mem.mem_internal.code_mem[251][2] ),
    .S1(net907),
    .X(_06598_));
 sg13g2_mux4_1 _25283_ (.S0(net975),
    .A0(\mem.mem_internal.code_mem[252][2] ),
    .A1(\mem.mem_internal.code_mem[253][2] ),
    .A2(\mem.mem_internal.code_mem[254][2] ),
    .A3(\mem.mem_internal.code_mem[255][2] ),
    .S1(_06208_),
    .X(_06599_));
 sg13g2_mux4_1 _25284_ (.S0(net971),
    .A0(_06596_),
    .A1(_06597_),
    .A2(_06598_),
    .A3(_06599_),
    .S1(net900),
    .X(_06600_));
 sg13g2_mux4_1 _25285_ (.S0(net1229),
    .A0(_06585_),
    .A1(_06590_),
    .A2(_06595_),
    .A3(_06600_),
    .S1(net1233),
    .X(_06601_));
 sg13g2_mux4_1 _25286_ (.S0(_06300_),
    .A0(_06538_),
    .A1(_06559_),
    .A2(_06580_),
    .A3(_06601_),
    .S1(_06301_),
    .X(_06602_));
 sg13g2_nor2_1 _25287_ (.A(_06304_),
    .B(_06602_),
    .Y(_06603_));
 sg13g2_a21oi_1 _25288_ (.A1(net832),
    .A2(_06516_),
    .Y(_06604_),
    .B1(_06603_));
 sg13g2_nand2_1 _25289_ (.Y(_06605_),
    .A(\mem.internal_data_out[2] ),
    .B(_06126_));
 sg13g2_o21ai_1 _25290_ (.B1(_06605_),
    .Y(_02422_),
    .A1(net546),
    .A2(_06604_));
 sg13g2_mux4_1 _25291_ (.S0(net538),
    .A0(\mem.mem_internal.data_mem[0][3] ),
    .A1(\mem.mem_internal.data_mem[1][3] ),
    .A2(\mem.mem_internal.data_mem[2][3] ),
    .A3(\mem.mem_internal.data_mem[3][3] ),
    .S1(net537),
    .X(_06606_));
 sg13g2_mux4_1 _25292_ (.S0(net545),
    .A0(\mem.mem_internal.data_mem[4][3] ),
    .A1(\mem.mem_internal.data_mem[5][3] ),
    .A2(\mem.mem_internal.data_mem[6][3] ),
    .A3(\mem.mem_internal.data_mem[7][3] ),
    .S1(net544),
    .X(_06607_));
 sg13g2_mux4_1 _25293_ (.S0(net577),
    .A0(\mem.mem_internal.data_mem[8][3] ),
    .A1(\mem.mem_internal.data_mem[9][3] ),
    .A2(\mem.mem_internal.data_mem[10][3] ),
    .A3(\mem.mem_internal.data_mem[11][3] ),
    .S1(net543),
    .X(_06608_));
 sg13g2_mux4_1 _25294_ (.S0(net542),
    .A0(\mem.mem_internal.data_mem[12][3] ),
    .A1(\mem.mem_internal.data_mem[13][3] ),
    .A2(\mem.mem_internal.data_mem[14][3] ),
    .A3(\mem.mem_internal.data_mem[15][3] ),
    .S1(net541),
    .X(_06609_));
 sg13g2_mux4_1 _25295_ (.S0(net818),
    .A0(_06606_),
    .A1(_06607_),
    .A2(_06608_),
    .A3(_06609_),
    .S1(_06170_),
    .X(_06610_));
 sg13g2_mux4_1 _25296_ (.S0(net540),
    .A0(\mem.mem_internal.data_mem[16][3] ),
    .A1(\mem.mem_internal.data_mem[17][3] ),
    .A2(\mem.mem_internal.data_mem[18][3] ),
    .A3(\mem.mem_internal.data_mem[19][3] ),
    .S1(net539),
    .X(_06611_));
 sg13g2_mux4_1 _25297_ (.S0(net538),
    .A0(\mem.mem_internal.data_mem[20][3] ),
    .A1(\mem.mem_internal.data_mem[21][3] ),
    .A2(\mem.mem_internal.data_mem[22][3] ),
    .A3(\mem.mem_internal.data_mem[23][3] ),
    .S1(net537),
    .X(_06612_));
 sg13g2_mux4_1 _25298_ (.S0(net576),
    .A0(\mem.mem_internal.data_mem[24][3] ),
    .A1(\mem.mem_internal.data_mem[25][3] ),
    .A2(\mem.mem_internal.data_mem[26][3] ),
    .A3(\mem.mem_internal.data_mem[27][3] ),
    .S1(net575),
    .X(_06613_));
 sg13g2_mux4_1 _25299_ (.S0(net576),
    .A0(\mem.mem_internal.data_mem[28][3] ),
    .A1(\mem.mem_internal.data_mem[29][3] ),
    .A2(\mem.mem_internal.data_mem[30][3] ),
    .A3(\mem.mem_internal.data_mem[31][3] ),
    .S1(net575),
    .X(_06614_));
 sg13g2_mux4_1 _25300_ (.S0(net988),
    .A0(_06611_),
    .A1(_06612_),
    .A2(_06613_),
    .A3(_06614_),
    .S1(net1235),
    .X(_06615_));
 sg13g2_mux2_1 _25301_ (.A0(_06610_),
    .A1(_06615_),
    .S(net817),
    .X(_06616_));
 sg13g2_mux4_1 _25302_ (.S0(net958),
    .A0(\mem.mem_internal.code_mem[0][3] ),
    .A1(\mem.mem_internal.code_mem[1][3] ),
    .A2(\mem.mem_internal.code_mem[2][3] ),
    .A3(\mem.mem_internal.code_mem[3][3] ),
    .S1(net814),
    .X(_06617_));
 sg13g2_mux4_1 _25303_ (.S0(net957),
    .A0(\mem.mem_internal.code_mem[4][3] ),
    .A1(\mem.mem_internal.code_mem[5][3] ),
    .A2(\mem.mem_internal.code_mem[6][3] ),
    .A3(\mem.mem_internal.code_mem[7][3] ),
    .S1(net813),
    .X(_06618_));
 sg13g2_mux4_1 _25304_ (.S0(net920),
    .A0(\mem.mem_internal.code_mem[16][3] ),
    .A1(\mem.mem_internal.code_mem[17][3] ),
    .A2(\mem.mem_internal.code_mem[18][3] ),
    .A3(\mem.mem_internal.code_mem[19][3] ),
    .S1(net955),
    .X(_06619_));
 sg13g2_mux4_1 _25305_ (.S0(net954),
    .A0(\mem.mem_internal.code_mem[20][3] ),
    .A1(\mem.mem_internal.code_mem[21][3] ),
    .A2(\mem.mem_internal.code_mem[22][3] ),
    .A3(\mem.mem_internal.code_mem[23][3] ),
    .S1(net953),
    .X(_06620_));
 sg13g2_mux4_1 _25306_ (.S0(net979),
    .A0(_06617_),
    .A1(_06618_),
    .A2(_06619_),
    .A3(_06620_),
    .S1(net951),
    .X(_06621_));
 sg13g2_mux4_1 _25307_ (.S0(_06321_),
    .A0(\mem.mem_internal.code_mem[8][3] ),
    .A1(\mem.mem_internal.code_mem[9][3] ),
    .A2(\mem.mem_internal.code_mem[10][3] ),
    .A3(\mem.mem_internal.code_mem[11][3] ),
    .S1(net812),
    .X(_06622_));
 sg13g2_mux4_1 _25308_ (.S0(net811),
    .A0(\mem.mem_internal.code_mem[12][3] ),
    .A1(\mem.mem_internal.code_mem[13][3] ),
    .A2(\mem.mem_internal.code_mem[14][3] ),
    .A3(\mem.mem_internal.code_mem[15][3] ),
    .S1(_06336_),
    .X(_06623_));
 sg13g2_mux4_1 _25309_ (.S0(net950),
    .A0(\mem.mem_internal.code_mem[24][3] ),
    .A1(\mem.mem_internal.code_mem[25][3] ),
    .A2(\mem.mem_internal.code_mem[26][3] ),
    .A3(\mem.mem_internal.code_mem[27][3] ),
    .S1(net809),
    .X(_06624_));
 sg13g2_mux4_1 _25310_ (.S0(net884),
    .A0(\mem.mem_internal.code_mem[28][3] ),
    .A1(\mem.mem_internal.code_mem[29][3] ),
    .A2(\mem.mem_internal.code_mem[30][3] ),
    .A3(\mem.mem_internal.code_mem[31][3] ),
    .S1(net804),
    .X(_06625_));
 sg13g2_mux4_1 _25311_ (.S0(net948),
    .A0(_06622_),
    .A1(_06623_),
    .A2(_06624_),
    .A3(_06625_),
    .S1(_06345_),
    .X(_06626_));
 sg13g2_mux4_1 _25312_ (.S0(_06324_),
    .A0(\mem.mem_internal.code_mem[128][3] ),
    .A1(\mem.mem_internal.code_mem[129][3] ),
    .A2(\mem.mem_internal.code_mem[130][3] ),
    .A3(\mem.mem_internal.code_mem[131][3] ),
    .S1(net946),
    .X(_06627_));
 sg13g2_mux4_1 _25313_ (.S0(_06349_),
    .A0(\mem.mem_internal.code_mem[132][3] ),
    .A1(\mem.mem_internal.code_mem[133][3] ),
    .A2(\mem.mem_internal.code_mem[134][3] ),
    .A3(\mem.mem_internal.code_mem[135][3] ),
    .S1(net808),
    .X(_06628_));
 sg13g2_mux4_1 _25314_ (.S0(net944),
    .A0(\mem.mem_internal.code_mem[144][3] ),
    .A1(\mem.mem_internal.code_mem[145][3] ),
    .A2(\mem.mem_internal.code_mem[146][3] ),
    .A3(\mem.mem_internal.code_mem[147][3] ),
    .S1(net943),
    .X(_06629_));
 sg13g2_mux4_1 _25315_ (.S0(net942),
    .A0(\mem.mem_internal.code_mem[148][3] ),
    .A1(\mem.mem_internal.code_mem[149][3] ),
    .A2(\mem.mem_internal.code_mem[150][3] ),
    .A3(\mem.mem_internal.code_mem[151][3] ),
    .S1(net941),
    .X(_06630_));
 sg13g2_mux4_1 _25316_ (.S0(net940),
    .A0(_06627_),
    .A1(_06628_),
    .A2(_06629_),
    .A3(_06630_),
    .S1(net939),
    .X(_06631_));
 sg13g2_mux4_1 _25317_ (.S0(net938),
    .A0(\mem.mem_internal.code_mem[136][3] ),
    .A1(\mem.mem_internal.code_mem[137][3] ),
    .A2(\mem.mem_internal.code_mem[138][3] ),
    .A3(\mem.mem_internal.code_mem[139][3] ),
    .S1(net899),
    .X(_06632_));
 sg13g2_mux4_1 _25318_ (.S0(net884),
    .A0(\mem.mem_internal.code_mem[140][3] ),
    .A1(\mem.mem_internal.code_mem[141][3] ),
    .A2(\mem.mem_internal.code_mem[142][3] ),
    .A3(\mem.mem_internal.code_mem[143][3] ),
    .S1(net797),
    .X(_06633_));
 sg13g2_mux4_1 _25319_ (.S0(net937),
    .A0(\mem.mem_internal.code_mem[152][3] ),
    .A1(\mem.mem_internal.code_mem[153][3] ),
    .A2(\mem.mem_internal.code_mem[154][3] ),
    .A3(\mem.mem_internal.code_mem[155][3] ),
    .S1(net936),
    .X(_06634_));
 sg13g2_mux4_1 _25320_ (.S0(net935),
    .A0(\mem.mem_internal.code_mem[156][3] ),
    .A1(\mem.mem_internal.code_mem[157][3] ),
    .A2(\mem.mem_internal.code_mem[158][3] ),
    .A3(\mem.mem_internal.code_mem[159][3] ),
    .S1(net934),
    .X(_06635_));
 sg13g2_mux4_1 _25321_ (.S0(net933),
    .A0(_06632_),
    .A1(_06633_),
    .A2(_06634_),
    .A3(_06635_),
    .S1(net932),
    .X(_06636_));
 sg13g2_mux4_1 _25322_ (.S0(net1234),
    .A0(_06621_),
    .A1(_06626_),
    .A2(_06631_),
    .A3(_06636_),
    .S1(_06376_),
    .X(_06637_));
 sg13g2_mux4_1 _25323_ (.S0(net931),
    .A0(\mem.mem_internal.code_mem[32][3] ),
    .A1(\mem.mem_internal.code_mem[33][3] ),
    .A2(\mem.mem_internal.code_mem[34][3] ),
    .A3(\mem.mem_internal.code_mem[35][3] ),
    .S1(net812),
    .X(_06638_));
 sg13g2_mux4_1 _25324_ (.S0(net803),
    .A0(\mem.mem_internal.code_mem[36][3] ),
    .A1(\mem.mem_internal.code_mem[37][3] ),
    .A2(\mem.mem_internal.code_mem[38][3] ),
    .A3(\mem.mem_internal.code_mem[39][3] ),
    .S1(net806),
    .X(_06639_));
 sg13g2_mux4_1 _25325_ (.S0(net930),
    .A0(\mem.mem_internal.code_mem[48][3] ),
    .A1(\mem.mem_internal.code_mem[49][3] ),
    .A2(\mem.mem_internal.code_mem[50][3] ),
    .A3(\mem.mem_internal.code_mem[51][3] ),
    .S1(net805),
    .X(_06640_));
 sg13g2_mux4_1 _25326_ (.S0(net929),
    .A0(\mem.mem_internal.code_mem[52][3] ),
    .A1(\mem.mem_internal.code_mem[53][3] ),
    .A2(\mem.mem_internal.code_mem[54][3] ),
    .A3(\mem.mem_internal.code_mem[55][3] ),
    .S1(net804),
    .X(_06641_));
 sg13g2_mux4_1 _25327_ (.S0(net952),
    .A0(_06638_),
    .A1(_06639_),
    .A2(_06640_),
    .A3(_06641_),
    .S1(net947),
    .X(_06642_));
 sg13g2_mux4_1 _25328_ (.S0(net803),
    .A0(\mem.mem_internal.code_mem[40][3] ),
    .A1(\mem.mem_internal.code_mem[41][3] ),
    .A2(\mem.mem_internal.code_mem[42][3] ),
    .A3(\mem.mem_internal.code_mem[43][3] ),
    .S1(net810),
    .X(_06643_));
 sg13g2_mux4_1 _25329_ (.S0(net820),
    .A0(\mem.mem_internal.code_mem[44][3] ),
    .A1(\mem.mem_internal.code_mem[45][3] ),
    .A2(\mem.mem_internal.code_mem[46][3] ),
    .A3(\mem.mem_internal.code_mem[47][3] ),
    .S1(net819),
    .X(_06644_));
 sg13g2_mux4_1 _25330_ (.S0(net928),
    .A0(\mem.mem_internal.code_mem[56][3] ),
    .A1(\mem.mem_internal.code_mem[57][3] ),
    .A2(\mem.mem_internal.code_mem[58][3] ),
    .A3(\mem.mem_internal.code_mem[59][3] ),
    .S1(net802),
    .X(_06645_));
 sg13g2_mux4_1 _25331_ (.S0(net927),
    .A0(\mem.mem_internal.code_mem[60][3] ),
    .A1(\mem.mem_internal.code_mem[61][3] ),
    .A2(\mem.mem_internal.code_mem[62][3] ),
    .A3(\mem.mem_internal.code_mem[63][3] ),
    .S1(net815),
    .X(_06646_));
 sg13g2_mux4_1 _25332_ (.S0(_06150_),
    .A0(_06643_),
    .A1(_06644_),
    .A2(_06645_),
    .A3(_06646_),
    .S1(net987),
    .X(_06647_));
 sg13g2_mux4_1 _25333_ (.S0(net945),
    .A0(\mem.mem_internal.code_mem[160][3] ),
    .A1(\mem.mem_internal.code_mem[161][3] ),
    .A2(\mem.mem_internal.code_mem[162][3] ),
    .A3(\mem.mem_internal.code_mem[163][3] ),
    .S1(net809),
    .X(_06648_));
 sg13g2_mux4_1 _25334_ (.S0(net928),
    .A0(\mem.mem_internal.code_mem[164][3] ),
    .A1(\mem.mem_internal.code_mem[165][3] ),
    .A2(\mem.mem_internal.code_mem[166][3] ),
    .A3(\mem.mem_internal.code_mem[167][3] ),
    .S1(net801),
    .X(_06649_));
 sg13g2_mux4_1 _25335_ (.S0(net925),
    .A0(\mem.mem_internal.code_mem[176][3] ),
    .A1(\mem.mem_internal.code_mem[177][3] ),
    .A2(\mem.mem_internal.code_mem[178][3] ),
    .A3(\mem.mem_internal.code_mem[179][3] ),
    .S1(net924),
    .X(_06650_));
 sg13g2_mux4_1 _25336_ (.S0(net962),
    .A0(\mem.mem_internal.code_mem[180][3] ),
    .A1(\mem.mem_internal.code_mem[181][3] ),
    .A2(\mem.mem_internal.code_mem[182][3] ),
    .A3(\mem.mem_internal.code_mem[183][3] ),
    .S1(net912),
    .X(_06651_));
 sg13g2_mux4_1 _25337_ (.S0(net923),
    .A0(_06648_),
    .A1(_06649_),
    .A2(_06650_),
    .A3(_06651_),
    .S1(net911),
    .X(_06652_));
 sg13g2_mux4_1 _25338_ (.S0(net949),
    .A0(\mem.mem_internal.code_mem[168][3] ),
    .A1(\mem.mem_internal.code_mem[169][3] ),
    .A2(\mem.mem_internal.code_mem[170][3] ),
    .A3(\mem.mem_internal.code_mem[171][3] ),
    .S1(net807),
    .X(_06653_));
 sg13g2_mux4_1 _25339_ (.S0(net984),
    .A0(\mem.mem_internal.code_mem[172][3] ),
    .A1(\mem.mem_internal.code_mem[173][3] ),
    .A2(\mem.mem_internal.code_mem[174][3] ),
    .A3(\mem.mem_internal.code_mem[175][3] ),
    .S1(net800),
    .X(_06654_));
 sg13g2_mux4_1 _25340_ (.S0(net894),
    .A0(\mem.mem_internal.code_mem[184][3] ),
    .A1(\mem.mem_internal.code_mem[185][3] ),
    .A2(\mem.mem_internal.code_mem[186][3] ),
    .A3(\mem.mem_internal.code_mem[187][3] ),
    .S1(net921),
    .X(_06655_));
 sg13g2_mux4_1 _25341_ (.S0(net981),
    .A0(\mem.mem_internal.code_mem[188][3] ),
    .A1(\mem.mem_internal.code_mem[189][3] ),
    .A2(\mem.mem_internal.code_mem[190][3] ),
    .A3(\mem.mem_internal.code_mem[191][3] ),
    .S1(net980),
    .X(_06656_));
 sg13g2_mux4_1 _25342_ (.S0(net891),
    .A0(_06653_),
    .A1(_06654_),
    .A2(_06655_),
    .A3(_06656_),
    .S1(net978),
    .X(_06657_));
 sg13g2_mux4_1 _25343_ (.S0(net1235),
    .A0(_06642_),
    .A1(_06647_),
    .A2(_06652_),
    .A3(_06657_),
    .S1(net1232),
    .X(_06658_));
 sg13g2_mux4_1 _25344_ (.S0(net965),
    .A0(\mem.mem_internal.code_mem[64][3] ),
    .A1(\mem.mem_internal.code_mem[65][3] ),
    .A2(\mem.mem_internal.code_mem[66][3] ),
    .A3(\mem.mem_internal.code_mem[67][3] ),
    .S1(net955),
    .X(_06659_));
 sg13g2_mux4_1 _25345_ (.S0(net919),
    .A0(\mem.mem_internal.code_mem[68][3] ),
    .A1(\mem.mem_internal.code_mem[69][3] ),
    .A2(\mem.mem_internal.code_mem[70][3] ),
    .A3(\mem.mem_internal.code_mem[71][3] ),
    .S1(net799),
    .X(_06660_));
 sg13g2_mux4_1 _25346_ (.S0(net918),
    .A0(\mem.mem_internal.code_mem[80][3] ),
    .A1(\mem.mem_internal.code_mem[81][3] ),
    .A2(\mem.mem_internal.code_mem[82][3] ),
    .A3(\mem.mem_internal.code_mem[83][3] ),
    .S1(net964),
    .X(_06661_));
 sg13g2_mux4_1 _25347_ (.S0(net916),
    .A0(\mem.mem_internal.code_mem[84][3] ),
    .A1(\mem.mem_internal.code_mem[85][3] ),
    .A2(\mem.mem_internal.code_mem[86][3] ),
    .A3(\mem.mem_internal.code_mem[87][3] ),
    .S1(net936),
    .X(_06662_));
 sg13g2_mux4_1 _25348_ (.S0(_06221_),
    .A0(_06659_),
    .A1(_06660_),
    .A2(_06661_),
    .A3(_06662_),
    .S1(net915),
    .X(_06663_));
 sg13g2_mux4_1 _25349_ (.S0(net919),
    .A0(\mem.mem_internal.code_mem[72][3] ),
    .A1(\mem.mem_internal.code_mem[73][3] ),
    .A2(\mem.mem_internal.code_mem[74][3] ),
    .A3(\mem.mem_internal.code_mem[75][3] ),
    .S1(_06420_),
    .X(_06664_));
 sg13g2_mux4_1 _25350_ (.S0(net985),
    .A0(\mem.mem_internal.code_mem[76][3] ),
    .A1(\mem.mem_internal.code_mem[77][3] ),
    .A2(\mem.mem_internal.code_mem[78][3] ),
    .A3(\mem.mem_internal.code_mem[79][3] ),
    .S1(net816),
    .X(_06665_));
 sg13g2_mux4_1 _25351_ (.S0(net914),
    .A0(\mem.mem_internal.code_mem[88][3] ),
    .A1(\mem.mem_internal.code_mem[89][3] ),
    .A2(\mem.mem_internal.code_mem[90][3] ),
    .A3(\mem.mem_internal.code_mem[91][3] ),
    .S1(net910),
    .X(_06666_));
 sg13g2_mux4_1 _25352_ (.S0(net913),
    .A0(\mem.mem_internal.code_mem[92][3] ),
    .A1(\mem.mem_internal.code_mem[93][3] ),
    .A2(\mem.mem_internal.code_mem[94][3] ),
    .A3(\mem.mem_internal.code_mem[95][3] ),
    .S1(_06434_),
    .X(_06667_));
 sg13g2_mux4_1 _25353_ (.S0(net933),
    .A0(_06664_),
    .A1(_06665_),
    .A2(_06666_),
    .A3(_06667_),
    .S1(_06436_),
    .X(_06668_));
 sg13g2_mux4_1 _25354_ (.S0(_06422_),
    .A0(\mem.mem_internal.code_mem[192][3] ),
    .A1(\mem.mem_internal.code_mem[193][3] ),
    .A2(\mem.mem_internal.code_mem[194][3] ),
    .A3(\mem.mem_internal.code_mem[195][3] ),
    .S1(net917),
    .X(_06669_));
 sg13g2_mux4_1 _25355_ (.S0(net942),
    .A0(\mem.mem_internal.code_mem[196][3] ),
    .A1(\mem.mem_internal.code_mem[197][3] ),
    .A2(\mem.mem_internal.code_mem[198][3] ),
    .A3(\mem.mem_internal.code_mem[199][3] ),
    .S1(_06439_),
    .X(_06670_));
 sg13g2_mux4_1 _25356_ (.S0(net959),
    .A0(\mem.mem_internal.code_mem[208][3] ),
    .A1(\mem.mem_internal.code_mem[209][3] ),
    .A2(\mem.mem_internal.code_mem[210][3] ),
    .A3(\mem.mem_internal.code_mem[211][3] ),
    .S1(net961),
    .X(_06671_));
 sg13g2_mux4_1 _25357_ (.S0(net908),
    .A0(\mem.mem_internal.code_mem[212][3] ),
    .A1(\mem.mem_internal.code_mem[213][3] ),
    .A2(\mem.mem_internal.code_mem[214][3] ),
    .A3(\mem.mem_internal.code_mem[215][3] ),
    .S1(net888),
    .X(_06672_));
 sg13g2_mux4_1 _25358_ (.S0(net1231),
    .A0(_06669_),
    .A1(_06670_),
    .A2(_06671_),
    .A3(_06672_),
    .S1(net960),
    .X(_06673_));
 sg13g2_mux4_1 _25359_ (.S0(_06448_),
    .A0(\mem.mem_internal.code_mem[200][3] ),
    .A1(\mem.mem_internal.code_mem[201][3] ),
    .A2(\mem.mem_internal.code_mem[202][3] ),
    .A3(\mem.mem_internal.code_mem[203][3] ),
    .S1(net905),
    .X(_06674_));
 sg13g2_mux4_1 _25360_ (.S0(_06433_),
    .A0(\mem.mem_internal.code_mem[204][3] ),
    .A1(\mem.mem_internal.code_mem[205][3] ),
    .A2(\mem.mem_internal.code_mem[206][3] ),
    .A3(\mem.mem_internal.code_mem[207][3] ),
    .S1(_06451_),
    .X(_06675_));
 sg13g2_mux4_1 _25361_ (.S0(net903),
    .A0(\mem.mem_internal.code_mem[216][3] ),
    .A1(\mem.mem_internal.code_mem[217][3] ),
    .A2(\mem.mem_internal.code_mem[218][3] ),
    .A3(\mem.mem_internal.code_mem[219][3] ),
    .S1(net909),
    .X(_06676_));
 sg13g2_mux4_1 _25362_ (.S0(_06455_),
    .A0(\mem.mem_internal.code_mem[220][3] ),
    .A1(\mem.mem_internal.code_mem[221][3] ),
    .A2(\mem.mem_internal.code_mem[222][3] ),
    .A3(\mem.mem_internal.code_mem[223][3] ),
    .S1(net901),
    .X(_06677_));
 sg13g2_mux4_1 _25363_ (.S0(net1230),
    .A0(_06674_),
    .A1(_06675_),
    .A2(_06676_),
    .A3(_06677_),
    .S1(_06459_),
    .X(_06678_));
 sg13g2_mux4_1 _25364_ (.S0(net1229),
    .A0(_06663_),
    .A1(_06668_),
    .A2(_06673_),
    .A3(_06678_),
    .S1(net1228),
    .X(_06679_));
 sg13g2_mux4_1 _25365_ (.S0(net956),
    .A0(\mem.mem_internal.code_mem[96][3] ),
    .A1(\mem.mem_internal.code_mem[97][3] ),
    .A2(\mem.mem_internal.code_mem[98][3] ),
    .A3(\mem.mem_internal.code_mem[99][3] ),
    .S1(_06464_),
    .X(_06680_));
 sg13g2_mux4_1 _25366_ (.S0(net895),
    .A0(\mem.mem_internal.code_mem[100][3] ),
    .A1(\mem.mem_internal.code_mem[101][3] ),
    .A2(\mem.mem_internal.code_mem[102][3] ),
    .A3(\mem.mem_internal.code_mem[103][3] ),
    .S1(net798),
    .X(_06681_));
 sg13g2_mux4_1 _25367_ (.S0(net906),
    .A0(\mem.mem_internal.code_mem[112][3] ),
    .A1(\mem.mem_internal.code_mem[113][3] ),
    .A2(\mem.mem_internal.code_mem[114][3] ),
    .A3(\mem.mem_internal.code_mem[115][3] ),
    .S1(net898),
    .X(_06682_));
 sg13g2_mux4_1 _25368_ (.S0(net897),
    .A0(\mem.mem_internal.code_mem[116][3] ),
    .A1(\mem.mem_internal.code_mem[117][3] ),
    .A2(\mem.mem_internal.code_mem[118][3] ),
    .A3(\mem.mem_internal.code_mem[119][3] ),
    .S1(net886),
    .X(_06683_));
 sg13g2_mux4_1 _25369_ (.S0(net896),
    .A0(_06680_),
    .A1(_06681_),
    .A2(_06682_),
    .A3(_06683_),
    .S1(net939),
    .X(_06684_));
 sg13g2_mux4_1 _25370_ (.S0(net895),
    .A0(\mem.mem_internal.code_mem[104][3] ),
    .A1(\mem.mem_internal.code_mem[105][3] ),
    .A2(\mem.mem_internal.code_mem[106][3] ),
    .A3(\mem.mem_internal.code_mem[107][3] ),
    .S1(_06475_),
    .X(_06685_));
 sg13g2_mux4_1 _25371_ (.S0(net926),
    .A0(\mem.mem_internal.code_mem[108][3] ),
    .A1(\mem.mem_internal.code_mem[109][3] ),
    .A2(\mem.mem_internal.code_mem[110][3] ),
    .A3(\mem.mem_internal.code_mem[111][3] ),
    .S1(net802),
    .X(_06686_));
 sg13g2_mux4_1 _25372_ (.S0(net894),
    .A0(\mem.mem_internal.code_mem[120][3] ),
    .A1(\mem.mem_internal.code_mem[121][3] ),
    .A2(\mem.mem_internal.code_mem[122][3] ),
    .A3(\mem.mem_internal.code_mem[123][3] ),
    .S1(net904),
    .X(_06687_));
 sg13g2_mux4_1 _25373_ (.S0(net893),
    .A0(\mem.mem_internal.code_mem[124][3] ),
    .A1(\mem.mem_internal.code_mem[125][3] ),
    .A2(\mem.mem_internal.code_mem[126][3] ),
    .A3(\mem.mem_internal.code_mem[127][3] ),
    .S1(net892),
    .X(_06688_));
 sg13g2_mux4_1 _25374_ (.S0(_06483_),
    .A0(_06685_),
    .A1(_06686_),
    .A2(_06687_),
    .A3(_06688_),
    .S1(net922),
    .X(_06689_));
 sg13g2_mux4_1 _25375_ (.S0(net944),
    .A0(\mem.mem_internal.code_mem[224][3] ),
    .A1(\mem.mem_internal.code_mem[225][3] ),
    .A2(\mem.mem_internal.code_mem[226][3] ),
    .A3(\mem.mem_internal.code_mem[227][3] ),
    .S1(net943),
    .X(_06690_));
 sg13g2_mux4_1 _25376_ (.S0(net890),
    .A0(\mem.mem_internal.code_mem[228][3] ),
    .A1(\mem.mem_internal.code_mem[229][3] ),
    .A2(\mem.mem_internal.code_mem[230][3] ),
    .A3(\mem.mem_internal.code_mem[231][3] ),
    .S1(net889),
    .X(_06691_));
 sg13g2_mux4_1 _25377_ (.S0(net908),
    .A0(\mem.mem_internal.code_mem[240][3] ),
    .A1(\mem.mem_internal.code_mem[241][3] ),
    .A2(\mem.mem_internal.code_mem[242][3] ),
    .A3(\mem.mem_internal.code_mem[243][3] ),
    .S1(net888),
    .X(_06692_));
 sg13g2_mux4_1 _25378_ (.S0(net902),
    .A0(\mem.mem_internal.code_mem[244][3] ),
    .A1(\mem.mem_internal.code_mem[245][3] ),
    .A2(\mem.mem_internal.code_mem[246][3] ),
    .A3(\mem.mem_internal.code_mem[247][3] ),
    .S1(net974),
    .X(_06693_));
 sg13g2_mux4_1 _25379_ (.S0(_06458_),
    .A0(_06690_),
    .A1(_06691_),
    .A2(_06692_),
    .A3(_06693_),
    .S1(net887),
    .X(_06694_));
 sg13g2_mux4_1 _25380_ (.S0(_06470_),
    .A0(\mem.mem_internal.code_mem[232][3] ),
    .A1(\mem.mem_internal.code_mem[233][3] ),
    .A2(\mem.mem_internal.code_mem[234][3] ),
    .A3(\mem.mem_internal.code_mem[235][3] ),
    .S1(net886),
    .X(_06695_));
 sg13g2_mux4_1 _25381_ (.S0(net983),
    .A0(\mem.mem_internal.code_mem[236][3] ),
    .A1(\mem.mem_internal.code_mem[237][3] ),
    .A2(\mem.mem_internal.code_mem[238][3] ),
    .A3(\mem.mem_internal.code_mem[239][3] ),
    .S1(net982),
    .X(_06696_));
 sg13g2_mux4_1 _25382_ (.S0(net885),
    .A0(\mem.mem_internal.code_mem[248][3] ),
    .A1(\mem.mem_internal.code_mem[249][3] ),
    .A2(\mem.mem_internal.code_mem[250][3] ),
    .A3(\mem.mem_internal.code_mem[251][3] ),
    .S1(net907),
    .X(_06697_));
 sg13g2_mux4_1 _25383_ (.S0(net975),
    .A0(\mem.mem_internal.code_mem[252][3] ),
    .A1(\mem.mem_internal.code_mem[253][3] ),
    .A2(\mem.mem_internal.code_mem[254][3] ),
    .A3(\mem.mem_internal.code_mem[255][3] ),
    .S1(_06208_),
    .X(_06698_));
 sg13g2_mux4_1 _25384_ (.S0(net971),
    .A0(_06695_),
    .A1(_06696_),
    .A2(_06697_),
    .A3(_06698_),
    .S1(net900),
    .X(_06699_));
 sg13g2_mux4_1 _25385_ (.S0(net1229),
    .A0(_06684_),
    .A1(_06689_),
    .A2(_06694_),
    .A3(_06699_),
    .S1(net1233),
    .X(_06700_));
 sg13g2_mux4_1 _25386_ (.S0(_06300_),
    .A0(_06637_),
    .A1(_06658_),
    .A2(_06679_),
    .A3(_06700_),
    .S1(_06301_),
    .X(_06701_));
 sg13g2_nor2_1 _25387_ (.A(_06304_),
    .B(_06701_),
    .Y(_06702_));
 sg13g2_a21oi_1 _25388_ (.A1(net832),
    .A2(_06616_),
    .Y(_06703_),
    .B1(_06702_));
 sg13g2_nand2_1 _25389_ (.Y(_06704_),
    .A(\mem.internal_data_out[3] ),
    .B(_06126_));
 sg13g2_o21ai_1 _25390_ (.B1(_06704_),
    .Y(_02423_),
    .A1(_06127_),
    .A2(_06703_));
 sg13g2_mux4_1 _25391_ (.S0(net538),
    .A0(\mem.mem_internal.data_mem[0][4] ),
    .A1(\mem.mem_internal.data_mem[1][4] ),
    .A2(\mem.mem_internal.data_mem[2][4] ),
    .A3(\mem.mem_internal.data_mem[3][4] ),
    .S1(net537),
    .X(_06705_));
 sg13g2_mux4_1 _25392_ (.S0(net545),
    .A0(\mem.mem_internal.data_mem[4][4] ),
    .A1(\mem.mem_internal.data_mem[5][4] ),
    .A2(\mem.mem_internal.data_mem[6][4] ),
    .A3(\mem.mem_internal.data_mem[7][4] ),
    .S1(net544),
    .X(_06706_));
 sg13g2_mux4_1 _25393_ (.S0(net577),
    .A0(\mem.mem_internal.data_mem[16][4] ),
    .A1(\mem.mem_internal.data_mem[17][4] ),
    .A2(\mem.mem_internal.data_mem[18][4] ),
    .A3(\mem.mem_internal.data_mem[19][4] ),
    .S1(net543),
    .X(_06707_));
 sg13g2_mux4_1 _25394_ (.S0(net542),
    .A0(\mem.mem_internal.data_mem[20][4] ),
    .A1(\mem.mem_internal.data_mem[21][4] ),
    .A2(\mem.mem_internal.data_mem[22][4] ),
    .A3(\mem.mem_internal.data_mem[23][4] ),
    .S1(net541),
    .X(_06708_));
 sg13g2_mux4_1 _25395_ (.S0(net818),
    .A0(_06705_),
    .A1(_06706_),
    .A2(_06707_),
    .A3(_06708_),
    .S1(net817),
    .X(_06709_));
 sg13g2_mux4_1 _25396_ (.S0(net540),
    .A0(\mem.mem_internal.data_mem[8][4] ),
    .A1(\mem.mem_internal.data_mem[9][4] ),
    .A2(\mem.mem_internal.data_mem[10][4] ),
    .A3(\mem.mem_internal.data_mem[11][4] ),
    .S1(net539),
    .X(_06710_));
 sg13g2_mux4_1 _25397_ (.S0(net540),
    .A0(\mem.mem_internal.data_mem[12][4] ),
    .A1(\mem.mem_internal.data_mem[13][4] ),
    .A2(\mem.mem_internal.data_mem[14][4] ),
    .A3(\mem.mem_internal.data_mem[15][4] ),
    .S1(net539),
    .X(_06711_));
 sg13g2_mux4_1 _25398_ (.S0(_06132_),
    .A0(\mem.mem_internal.data_mem[24][4] ),
    .A1(\mem.mem_internal.data_mem[25][4] ),
    .A2(\mem.mem_internal.data_mem[26][4] ),
    .A3(\mem.mem_internal.data_mem[27][4] ),
    .S1(net578),
    .X(_06712_));
 sg13g2_mux4_1 _25399_ (.S0(net576),
    .A0(\mem.mem_internal.data_mem[28][4] ),
    .A1(\mem.mem_internal.data_mem[29][4] ),
    .A2(\mem.mem_internal.data_mem[30][4] ),
    .A3(\mem.mem_internal.data_mem[31][4] ),
    .S1(net575),
    .X(_06713_));
 sg13g2_mux4_1 _25400_ (.S0(net988),
    .A0(_06710_),
    .A1(_06711_),
    .A2(_06712_),
    .A3(_06713_),
    .S1(net817),
    .X(_06714_));
 sg13g2_mux2_1 _25401_ (.A0(_06709_),
    .A1(_06714_),
    .S(net986),
    .X(_06715_));
 sg13g2_mux4_1 _25402_ (.S0(net958),
    .A0(\mem.mem_internal.code_mem[0][4] ),
    .A1(\mem.mem_internal.code_mem[1][4] ),
    .A2(\mem.mem_internal.code_mem[2][4] ),
    .A3(\mem.mem_internal.code_mem[3][4] ),
    .S1(net814),
    .X(_06716_));
 sg13g2_mux4_1 _25403_ (.S0(net957),
    .A0(\mem.mem_internal.code_mem[4][4] ),
    .A1(\mem.mem_internal.code_mem[5][4] ),
    .A2(\mem.mem_internal.code_mem[6][4] ),
    .A3(\mem.mem_internal.code_mem[7][4] ),
    .S1(net813),
    .X(_06717_));
 sg13g2_mux4_1 _25404_ (.S0(net920),
    .A0(\mem.mem_internal.code_mem[16][4] ),
    .A1(\mem.mem_internal.code_mem[17][4] ),
    .A2(\mem.mem_internal.code_mem[18][4] ),
    .A3(\mem.mem_internal.code_mem[19][4] ),
    .S1(net955),
    .X(_06718_));
 sg13g2_mux4_1 _25405_ (.S0(net954),
    .A0(\mem.mem_internal.code_mem[20][4] ),
    .A1(\mem.mem_internal.code_mem[21][4] ),
    .A2(\mem.mem_internal.code_mem[22][4] ),
    .A3(\mem.mem_internal.code_mem[23][4] ),
    .S1(net953),
    .X(_06719_));
 sg13g2_mux4_1 _25406_ (.S0(net979),
    .A0(_06716_),
    .A1(_06717_),
    .A2(_06718_),
    .A3(_06719_),
    .S1(net951),
    .X(_06720_));
 sg13g2_mux4_1 _25407_ (.S0(_06321_),
    .A0(\mem.mem_internal.code_mem[8][4] ),
    .A1(\mem.mem_internal.code_mem[9][4] ),
    .A2(\mem.mem_internal.code_mem[10][4] ),
    .A3(\mem.mem_internal.code_mem[11][4] ),
    .S1(net812),
    .X(_06721_));
 sg13g2_mux4_1 _25408_ (.S0(net811),
    .A0(\mem.mem_internal.code_mem[12][4] ),
    .A1(\mem.mem_internal.code_mem[13][4] ),
    .A2(\mem.mem_internal.code_mem[14][4] ),
    .A3(\mem.mem_internal.code_mem[15][4] ),
    .S1(_06336_),
    .X(_06722_));
 sg13g2_mux4_1 _25409_ (.S0(net950),
    .A0(\mem.mem_internal.code_mem[24][4] ),
    .A1(\mem.mem_internal.code_mem[25][4] ),
    .A2(\mem.mem_internal.code_mem[26][4] ),
    .A3(\mem.mem_internal.code_mem[27][4] ),
    .S1(net809),
    .X(_06723_));
 sg13g2_mux4_1 _25410_ (.S0(net884),
    .A0(\mem.mem_internal.code_mem[28][4] ),
    .A1(\mem.mem_internal.code_mem[29][4] ),
    .A2(\mem.mem_internal.code_mem[30][4] ),
    .A3(\mem.mem_internal.code_mem[31][4] ),
    .S1(net804),
    .X(_06724_));
 sg13g2_mux4_1 _25411_ (.S0(net948),
    .A0(_06721_),
    .A1(_06722_),
    .A2(_06723_),
    .A3(_06724_),
    .S1(net951),
    .X(_06725_));
 sg13g2_mux4_1 _25412_ (.S0(net920),
    .A0(\mem.mem_internal.code_mem[128][4] ),
    .A1(\mem.mem_internal.code_mem[129][4] ),
    .A2(\mem.mem_internal.code_mem[130][4] ),
    .A3(\mem.mem_internal.code_mem[131][4] ),
    .S1(net946),
    .X(_06726_));
 sg13g2_mux4_1 _25413_ (.S0(_06349_),
    .A0(\mem.mem_internal.code_mem[132][4] ),
    .A1(\mem.mem_internal.code_mem[133][4] ),
    .A2(\mem.mem_internal.code_mem[134][4] ),
    .A3(\mem.mem_internal.code_mem[135][4] ),
    .S1(net808),
    .X(_06727_));
 sg13g2_mux4_1 _25414_ (.S0(net918),
    .A0(\mem.mem_internal.code_mem[144][4] ),
    .A1(\mem.mem_internal.code_mem[145][4] ),
    .A2(\mem.mem_internal.code_mem[146][4] ),
    .A3(\mem.mem_internal.code_mem[147][4] ),
    .S1(net943),
    .X(_06728_));
 sg13g2_mux4_1 _25415_ (.S0(net942),
    .A0(\mem.mem_internal.code_mem[148][4] ),
    .A1(\mem.mem_internal.code_mem[149][4] ),
    .A2(\mem.mem_internal.code_mem[150][4] ),
    .A3(\mem.mem_internal.code_mem[151][4] ),
    .S1(net941),
    .X(_06729_));
 sg13g2_mux4_1 _25416_ (.S0(net940),
    .A0(_06726_),
    .A1(_06727_),
    .A2(_06728_),
    .A3(_06729_),
    .S1(net915),
    .X(_06730_));
 sg13g2_mux4_1 _25417_ (.S0(net938),
    .A0(\mem.mem_internal.code_mem[136][4] ),
    .A1(\mem.mem_internal.code_mem[137][4] ),
    .A2(\mem.mem_internal.code_mem[138][4] ),
    .A3(\mem.mem_internal.code_mem[139][4] ),
    .S1(net899),
    .X(_06731_));
 sg13g2_mux4_1 _25418_ (.S0(net884),
    .A0(\mem.mem_internal.code_mem[140][4] ),
    .A1(\mem.mem_internal.code_mem[141][4] ),
    .A2(\mem.mem_internal.code_mem[142][4] ),
    .A3(\mem.mem_internal.code_mem[143][4] ),
    .S1(net797),
    .X(_06732_));
 sg13g2_mux4_1 _25419_ (.S0(net937),
    .A0(\mem.mem_internal.code_mem[152][4] ),
    .A1(\mem.mem_internal.code_mem[153][4] ),
    .A2(\mem.mem_internal.code_mem[154][4] ),
    .A3(\mem.mem_internal.code_mem[155][4] ),
    .S1(net898),
    .X(_06733_));
 sg13g2_mux4_1 _25420_ (.S0(net935),
    .A0(\mem.mem_internal.code_mem[156][4] ),
    .A1(\mem.mem_internal.code_mem[157][4] ),
    .A2(\mem.mem_internal.code_mem[158][4] ),
    .A3(\mem.mem_internal.code_mem[159][4] ),
    .S1(net934),
    .X(_06734_));
 sg13g2_mux4_1 _25421_ (.S0(net896),
    .A0(_06731_),
    .A1(_06732_),
    .A2(_06733_),
    .A3(_06734_),
    .S1(net932),
    .X(_06735_));
 sg13g2_mux4_1 _25422_ (.S0(net1234),
    .A0(_06720_),
    .A1(_06725_),
    .A2(_06730_),
    .A3(_06735_),
    .S1(_06225_),
    .X(_06736_));
 sg13g2_mux4_1 _25423_ (.S0(net931),
    .A0(\mem.mem_internal.code_mem[32][4] ),
    .A1(\mem.mem_internal.code_mem[33][4] ),
    .A2(\mem.mem_internal.code_mem[34][4] ),
    .A3(\mem.mem_internal.code_mem[35][4] ),
    .S1(net813),
    .X(_06737_));
 sg13g2_mux4_1 _25424_ (.S0(net803),
    .A0(\mem.mem_internal.code_mem[36][4] ),
    .A1(\mem.mem_internal.code_mem[37][4] ),
    .A2(\mem.mem_internal.code_mem[38][4] ),
    .A3(\mem.mem_internal.code_mem[39][4] ),
    .S1(net806),
    .X(_06738_));
 sg13g2_mux4_1 _25425_ (.S0(net930),
    .A0(\mem.mem_internal.code_mem[48][4] ),
    .A1(\mem.mem_internal.code_mem[49][4] ),
    .A2(\mem.mem_internal.code_mem[50][4] ),
    .A3(\mem.mem_internal.code_mem[51][4] ),
    .S1(net805),
    .X(_06739_));
 sg13g2_mux4_1 _25426_ (.S0(net929),
    .A0(\mem.mem_internal.code_mem[52][4] ),
    .A1(\mem.mem_internal.code_mem[53][4] ),
    .A2(\mem.mem_internal.code_mem[54][4] ),
    .A3(\mem.mem_internal.code_mem[55][4] ),
    .S1(net804),
    .X(_06740_));
 sg13g2_mux4_1 _25427_ (.S0(net952),
    .A0(_06737_),
    .A1(_06738_),
    .A2(_06739_),
    .A3(_06740_),
    .S1(net947),
    .X(_06741_));
 sg13g2_mux4_1 _25428_ (.S0(_06389_),
    .A0(\mem.mem_internal.code_mem[40][4] ),
    .A1(\mem.mem_internal.code_mem[41][4] ),
    .A2(\mem.mem_internal.code_mem[42][4] ),
    .A3(\mem.mem_internal.code_mem[43][4] ),
    .S1(net810),
    .X(_06742_));
 sg13g2_mux4_1 _25429_ (.S0(net820),
    .A0(\mem.mem_internal.code_mem[44][4] ),
    .A1(\mem.mem_internal.code_mem[45][4] ),
    .A2(\mem.mem_internal.code_mem[46][4] ),
    .A3(\mem.mem_internal.code_mem[47][4] ),
    .S1(net819),
    .X(_06743_));
 sg13g2_mux4_1 _25430_ (.S0(_06392_),
    .A0(\mem.mem_internal.code_mem[56][4] ),
    .A1(\mem.mem_internal.code_mem[57][4] ),
    .A2(\mem.mem_internal.code_mem[58][4] ),
    .A3(\mem.mem_internal.code_mem[59][4] ),
    .S1(net802),
    .X(_06744_));
 sg13g2_mux4_1 _25431_ (.S0(net927),
    .A0(\mem.mem_internal.code_mem[60][4] ),
    .A1(\mem.mem_internal.code_mem[61][4] ),
    .A2(\mem.mem_internal.code_mem[62][4] ),
    .A3(\mem.mem_internal.code_mem[63][4] ),
    .S1(net815),
    .X(_06745_));
 sg13g2_mux4_1 _25432_ (.S0(net948),
    .A0(_06742_),
    .A1(_06743_),
    .A2(_06744_),
    .A3(_06745_),
    .S1(net987),
    .X(_06746_));
 sg13g2_mux4_1 _25433_ (.S0(net945),
    .A0(\mem.mem_internal.code_mem[160][4] ),
    .A1(\mem.mem_internal.code_mem[161][4] ),
    .A2(\mem.mem_internal.code_mem[162][4] ),
    .A3(\mem.mem_internal.code_mem[163][4] ),
    .S1(net805),
    .X(_06747_));
 sg13g2_mux4_1 _25434_ (.S0(net928),
    .A0(\mem.mem_internal.code_mem[164][4] ),
    .A1(\mem.mem_internal.code_mem[165][4] ),
    .A2(\mem.mem_internal.code_mem[166][4] ),
    .A3(\mem.mem_internal.code_mem[167][4] ),
    .S1(net801),
    .X(_06748_));
 sg13g2_mux4_1 _25435_ (.S0(net925),
    .A0(\mem.mem_internal.code_mem[176][4] ),
    .A1(\mem.mem_internal.code_mem[177][4] ),
    .A2(\mem.mem_internal.code_mem[178][4] ),
    .A3(\mem.mem_internal.code_mem[179][4] ),
    .S1(net924),
    .X(_06749_));
 sg13g2_mux4_1 _25436_ (.S0(net962),
    .A0(\mem.mem_internal.code_mem[180][4] ),
    .A1(\mem.mem_internal.code_mem[181][4] ),
    .A2(\mem.mem_internal.code_mem[182][4] ),
    .A3(\mem.mem_internal.code_mem[183][4] ),
    .S1(net912),
    .X(_06750_));
 sg13g2_mux4_1 _25437_ (.S0(net923),
    .A0(_06747_),
    .A1(_06748_),
    .A2(_06749_),
    .A3(_06750_),
    .S1(net911),
    .X(_06751_));
 sg13g2_mux4_1 _25438_ (.S0(net949),
    .A0(\mem.mem_internal.code_mem[168][4] ),
    .A1(\mem.mem_internal.code_mem[169][4] ),
    .A2(\mem.mem_internal.code_mem[170][4] ),
    .A3(\mem.mem_internal.code_mem[171][4] ),
    .S1(net807),
    .X(_06752_));
 sg13g2_mux4_1 _25439_ (.S0(net927),
    .A0(\mem.mem_internal.code_mem[172][4] ),
    .A1(\mem.mem_internal.code_mem[173][4] ),
    .A2(\mem.mem_internal.code_mem[174][4] ),
    .A3(\mem.mem_internal.code_mem[175][4] ),
    .S1(net800),
    .X(_06753_));
 sg13g2_mux4_1 _25440_ (.S0(net894),
    .A0(\mem.mem_internal.code_mem[184][4] ),
    .A1(\mem.mem_internal.code_mem[185][4] ),
    .A2(\mem.mem_internal.code_mem[186][4] ),
    .A3(\mem.mem_internal.code_mem[187][4] ),
    .S1(net921),
    .X(_06754_));
 sg13g2_mux4_1 _25441_ (.S0(net893),
    .A0(\mem.mem_internal.code_mem[188][4] ),
    .A1(\mem.mem_internal.code_mem[189][4] ),
    .A2(\mem.mem_internal.code_mem[190][4] ),
    .A3(\mem.mem_internal.code_mem[191][4] ),
    .S1(net980),
    .X(_06755_));
 sg13g2_mux4_1 _25442_ (.S0(net891),
    .A0(_06752_),
    .A1(_06753_),
    .A2(_06754_),
    .A3(_06755_),
    .S1(net978),
    .X(_06756_));
 sg13g2_mux4_1 _25443_ (.S0(net1235),
    .A0(_06741_),
    .A1(_06746_),
    .A2(_06751_),
    .A3(_06756_),
    .S1(net1232),
    .X(_06757_));
 sg13g2_mux4_1 _25444_ (.S0(net965),
    .A0(\mem.mem_internal.code_mem[64][4] ),
    .A1(\mem.mem_internal.code_mem[65][4] ),
    .A2(\mem.mem_internal.code_mem[66][4] ),
    .A3(\mem.mem_internal.code_mem[67][4] ),
    .S1(net966),
    .X(_06758_));
 sg13g2_mux4_1 _25445_ (.S0(_06419_),
    .A0(\mem.mem_internal.code_mem[68][4] ),
    .A1(\mem.mem_internal.code_mem[69][4] ),
    .A2(\mem.mem_internal.code_mem[70][4] ),
    .A3(\mem.mem_internal.code_mem[71][4] ),
    .S1(net799),
    .X(_06759_));
 sg13g2_mux4_1 _25446_ (.S0(net963),
    .A0(\mem.mem_internal.code_mem[80][4] ),
    .A1(\mem.mem_internal.code_mem[81][4] ),
    .A2(\mem.mem_internal.code_mem[82][4] ),
    .A3(\mem.mem_internal.code_mem[83][4] ),
    .S1(net964),
    .X(_06760_));
 sg13g2_mux4_1 _25447_ (.S0(net916),
    .A0(\mem.mem_internal.code_mem[84][4] ),
    .A1(\mem.mem_internal.code_mem[85][4] ),
    .A2(\mem.mem_internal.code_mem[86][4] ),
    .A3(\mem.mem_internal.code_mem[87][4] ),
    .S1(net936),
    .X(_06761_));
 sg13g2_mux4_1 _25448_ (.S0(net967),
    .A0(_06758_),
    .A1(_06759_),
    .A2(_06760_),
    .A3(_06761_),
    .S1(net915),
    .X(_06762_));
 sg13g2_mux4_1 _25449_ (.S0(net938),
    .A0(\mem.mem_internal.code_mem[72][4] ),
    .A1(\mem.mem_internal.code_mem[73][4] ),
    .A2(\mem.mem_internal.code_mem[74][4] ),
    .A3(\mem.mem_internal.code_mem[75][4] ),
    .S1(net799),
    .X(_06763_));
 sg13g2_mux4_1 _25450_ (.S0(net985),
    .A0(\mem.mem_internal.code_mem[76][4] ),
    .A1(\mem.mem_internal.code_mem[77][4] ),
    .A2(\mem.mem_internal.code_mem[78][4] ),
    .A3(\mem.mem_internal.code_mem[79][4] ),
    .S1(net816),
    .X(_06764_));
 sg13g2_mux4_1 _25451_ (.S0(net914),
    .A0(\mem.mem_internal.code_mem[88][4] ),
    .A1(\mem.mem_internal.code_mem[89][4] ),
    .A2(\mem.mem_internal.code_mem[90][4] ),
    .A3(\mem.mem_internal.code_mem[91][4] ),
    .S1(net910),
    .X(_06765_));
 sg13g2_mux4_1 _25452_ (.S0(net913),
    .A0(\mem.mem_internal.code_mem[92][4] ),
    .A1(\mem.mem_internal.code_mem[93][4] ),
    .A2(\mem.mem_internal.code_mem[94][4] ),
    .A3(\mem.mem_internal.code_mem[95][4] ),
    .S1(_06434_),
    .X(_06766_));
 sg13g2_mux4_1 _25453_ (.S0(net933),
    .A0(_06763_),
    .A1(_06764_),
    .A2(_06765_),
    .A3(_06766_),
    .S1(_06436_),
    .X(_06767_));
 sg13g2_mux4_1 _25454_ (.S0(net963),
    .A0(\mem.mem_internal.code_mem[192][4] ),
    .A1(\mem.mem_internal.code_mem[193][4] ),
    .A2(\mem.mem_internal.code_mem[194][4] ),
    .A3(\mem.mem_internal.code_mem[195][4] ),
    .S1(net917),
    .X(_06768_));
 sg13g2_mux4_1 _25455_ (.S0(net942),
    .A0(\mem.mem_internal.code_mem[196][4] ),
    .A1(\mem.mem_internal.code_mem[197][4] ),
    .A2(\mem.mem_internal.code_mem[198][4] ),
    .A3(\mem.mem_internal.code_mem[199][4] ),
    .S1(_06439_),
    .X(_06769_));
 sg13g2_mux4_1 _25456_ (.S0(net959),
    .A0(\mem.mem_internal.code_mem[208][4] ),
    .A1(\mem.mem_internal.code_mem[209][4] ),
    .A2(\mem.mem_internal.code_mem[210][4] ),
    .A3(\mem.mem_internal.code_mem[211][4] ),
    .S1(net961),
    .X(_06770_));
 sg13g2_mux4_1 _25457_ (.S0(net908),
    .A0(\mem.mem_internal.code_mem[212][4] ),
    .A1(\mem.mem_internal.code_mem[213][4] ),
    .A2(\mem.mem_internal.code_mem[214][4] ),
    .A3(\mem.mem_internal.code_mem[215][4] ),
    .S1(net888),
    .X(_06771_));
 sg13g2_mux4_1 _25458_ (.S0(net1231),
    .A0(_06768_),
    .A1(_06769_),
    .A2(_06770_),
    .A3(_06771_),
    .S1(net960),
    .X(_06772_));
 sg13g2_mux4_1 _25459_ (.S0(_06448_),
    .A0(\mem.mem_internal.code_mem[200][4] ),
    .A1(\mem.mem_internal.code_mem[201][4] ),
    .A2(\mem.mem_internal.code_mem[202][4] ),
    .A3(\mem.mem_internal.code_mem[203][4] ),
    .S1(net905),
    .X(_06773_));
 sg13g2_mux4_1 _25460_ (.S0(_06433_),
    .A0(\mem.mem_internal.code_mem[204][4] ),
    .A1(\mem.mem_internal.code_mem[205][4] ),
    .A2(\mem.mem_internal.code_mem[206][4] ),
    .A3(\mem.mem_internal.code_mem[207][4] ),
    .S1(net889),
    .X(_06774_));
 sg13g2_mux4_1 _25461_ (.S0(net903),
    .A0(\mem.mem_internal.code_mem[216][4] ),
    .A1(\mem.mem_internal.code_mem[217][4] ),
    .A2(\mem.mem_internal.code_mem[218][4] ),
    .A3(\mem.mem_internal.code_mem[219][4] ),
    .S1(net909),
    .X(_06775_));
 sg13g2_mux4_1 _25462_ (.S0(_06455_),
    .A0(\mem.mem_internal.code_mem[220][4] ),
    .A1(\mem.mem_internal.code_mem[221][4] ),
    .A2(\mem.mem_internal.code_mem[222][4] ),
    .A3(\mem.mem_internal.code_mem[223][4] ),
    .S1(net901),
    .X(_06776_));
 sg13g2_mux4_1 _25463_ (.S0(net1230),
    .A0(_06773_),
    .A1(_06774_),
    .A2(_06775_),
    .A3(_06776_),
    .S1(_06459_),
    .X(_06777_));
 sg13g2_mux4_1 _25464_ (.S0(net1229),
    .A0(_06762_),
    .A1(_06767_),
    .A2(_06772_),
    .A3(_06777_),
    .S1(net1228),
    .X(_06778_));
 sg13g2_mux4_1 _25465_ (.S0(net956),
    .A0(\mem.mem_internal.code_mem[96][4] ),
    .A1(\mem.mem_internal.code_mem[97][4] ),
    .A2(\mem.mem_internal.code_mem[98][4] ),
    .A3(\mem.mem_internal.code_mem[99][4] ),
    .S1(_06464_),
    .X(_06779_));
 sg13g2_mux4_1 _25466_ (.S0(net895),
    .A0(\mem.mem_internal.code_mem[100][4] ),
    .A1(\mem.mem_internal.code_mem[101][4] ),
    .A2(\mem.mem_internal.code_mem[102][4] ),
    .A3(\mem.mem_internal.code_mem[103][4] ),
    .S1(net798),
    .X(_06780_));
 sg13g2_mux4_1 _25467_ (.S0(net906),
    .A0(\mem.mem_internal.code_mem[112][4] ),
    .A1(\mem.mem_internal.code_mem[113][4] ),
    .A2(\mem.mem_internal.code_mem[114][4] ),
    .A3(\mem.mem_internal.code_mem[115][4] ),
    .S1(net898),
    .X(_06781_));
 sg13g2_mux4_1 _25468_ (.S0(net897),
    .A0(\mem.mem_internal.code_mem[116][4] ),
    .A1(\mem.mem_internal.code_mem[117][4] ),
    .A2(\mem.mem_internal.code_mem[118][4] ),
    .A3(\mem.mem_internal.code_mem[119][4] ),
    .S1(net886),
    .X(_06782_));
 sg13g2_mux4_1 _25469_ (.S0(net896),
    .A0(_06779_),
    .A1(_06780_),
    .A2(_06781_),
    .A3(_06782_),
    .S1(net939),
    .X(_06783_));
 sg13g2_mux4_1 _25470_ (.S0(net895),
    .A0(\mem.mem_internal.code_mem[104][4] ),
    .A1(\mem.mem_internal.code_mem[105][4] ),
    .A2(\mem.mem_internal.code_mem[106][4] ),
    .A3(\mem.mem_internal.code_mem[107][4] ),
    .S1(_06475_),
    .X(_06784_));
 sg13g2_mux4_1 _25471_ (.S0(net926),
    .A0(\mem.mem_internal.code_mem[108][4] ),
    .A1(\mem.mem_internal.code_mem[109][4] ),
    .A2(\mem.mem_internal.code_mem[110][4] ),
    .A3(\mem.mem_internal.code_mem[111][4] ),
    .S1(net802),
    .X(_06785_));
 sg13g2_mux4_1 _25472_ (.S0(_06478_),
    .A0(\mem.mem_internal.code_mem[120][4] ),
    .A1(\mem.mem_internal.code_mem[121][4] ),
    .A2(\mem.mem_internal.code_mem[122][4] ),
    .A3(\mem.mem_internal.code_mem[123][4] ),
    .S1(net904),
    .X(_06786_));
 sg13g2_mux4_1 _25473_ (.S0(net893),
    .A0(\mem.mem_internal.code_mem[124][4] ),
    .A1(\mem.mem_internal.code_mem[125][4] ),
    .A2(\mem.mem_internal.code_mem[126][4] ),
    .A3(\mem.mem_internal.code_mem[127][4] ),
    .S1(net892),
    .X(_06787_));
 sg13g2_mux4_1 _25474_ (.S0(_06483_),
    .A0(_06784_),
    .A1(_06785_),
    .A2(_06786_),
    .A3(_06787_),
    .S1(net922),
    .X(_06788_));
 sg13g2_mux4_1 _25475_ (.S0(net944),
    .A0(\mem.mem_internal.code_mem[224][4] ),
    .A1(\mem.mem_internal.code_mem[225][4] ),
    .A2(\mem.mem_internal.code_mem[226][4] ),
    .A3(\mem.mem_internal.code_mem[227][4] ),
    .S1(net943),
    .X(_06789_));
 sg13g2_mux4_1 _25476_ (.S0(net890),
    .A0(\mem.mem_internal.code_mem[228][4] ),
    .A1(\mem.mem_internal.code_mem[229][4] ),
    .A2(\mem.mem_internal.code_mem[230][4] ),
    .A3(\mem.mem_internal.code_mem[231][4] ),
    .S1(net889),
    .X(_06790_));
 sg13g2_mux4_1 _25477_ (.S0(net903),
    .A0(\mem.mem_internal.code_mem[240][4] ),
    .A1(\mem.mem_internal.code_mem[241][4] ),
    .A2(\mem.mem_internal.code_mem[242][4] ),
    .A3(\mem.mem_internal.code_mem[243][4] ),
    .S1(net888),
    .X(_06791_));
 sg13g2_mux4_1 _25478_ (.S0(net902),
    .A0(\mem.mem_internal.code_mem[244][4] ),
    .A1(\mem.mem_internal.code_mem[245][4] ),
    .A2(\mem.mem_internal.code_mem[246][4] ),
    .A3(\mem.mem_internal.code_mem[247][4] ),
    .S1(net901),
    .X(_06792_));
 sg13g2_mux4_1 _25479_ (.S0(net1231),
    .A0(_06789_),
    .A1(_06790_),
    .A2(_06791_),
    .A3(_06792_),
    .S1(net887),
    .X(_06793_));
 sg13g2_mux4_1 _25480_ (.S0(net925),
    .A0(\mem.mem_internal.code_mem[232][4] ),
    .A1(\mem.mem_internal.code_mem[233][4] ),
    .A2(\mem.mem_internal.code_mem[234][4] ),
    .A3(\mem.mem_internal.code_mem[235][4] ),
    .S1(_06494_),
    .X(_06794_));
 sg13g2_mux4_1 _25481_ (.S0(net983),
    .A0(\mem.mem_internal.code_mem[236][4] ),
    .A1(\mem.mem_internal.code_mem[237][4] ),
    .A2(\mem.mem_internal.code_mem[238][4] ),
    .A3(\mem.mem_internal.code_mem[239][4] ),
    .S1(net982),
    .X(_06795_));
 sg13g2_mux4_1 _25482_ (.S0(net885),
    .A0(\mem.mem_internal.code_mem[248][4] ),
    .A1(\mem.mem_internal.code_mem[249][4] ),
    .A2(\mem.mem_internal.code_mem[250][4] ),
    .A3(\mem.mem_internal.code_mem[251][4] ),
    .S1(net907),
    .X(_06796_));
 sg13g2_mux4_1 _25483_ (.S0(net975),
    .A0(\mem.mem_internal.code_mem[252][4] ),
    .A1(\mem.mem_internal.code_mem[253][4] ),
    .A2(\mem.mem_internal.code_mem[254][4] ),
    .A3(\mem.mem_internal.code_mem[255][4] ),
    .S1(net974),
    .X(_06797_));
 sg13g2_mux4_1 _25484_ (.S0(net971),
    .A0(_06794_),
    .A1(_06795_),
    .A2(_06796_),
    .A3(_06797_),
    .S1(net900),
    .X(_06798_));
 sg13g2_mux4_1 _25485_ (.S0(net1229),
    .A0(_06783_),
    .A1(_06788_),
    .A2(_06793_),
    .A3(_06798_),
    .S1(net1233),
    .X(_06799_));
 sg13g2_mux4_1 _25486_ (.S0(_06300_),
    .A0(_06736_),
    .A1(_06757_),
    .A2(_06778_),
    .A3(_06799_),
    .S1(_06301_),
    .X(_06800_));
 sg13g2_nor2_1 _25487_ (.A(_06304_),
    .B(_06800_),
    .Y(_06801_));
 sg13g2_a21oi_1 _25488_ (.A1(net832),
    .A2(_06715_),
    .Y(_06802_),
    .B1(_06801_));
 sg13g2_nand2_1 _25489_ (.Y(_06803_),
    .A(\mem.internal_data_out[4] ),
    .B(_06126_));
 sg13g2_o21ai_1 _25490_ (.B1(_06803_),
    .Y(_02424_),
    .A1(net546),
    .A2(_06802_));
 sg13g2_mux4_1 _25491_ (.S0(_06160_),
    .A0(\mem.mem_internal.data_mem[0][5] ),
    .A1(\mem.mem_internal.data_mem[1][5] ),
    .A2(\mem.mem_internal.data_mem[2][5] ),
    .A3(\mem.mem_internal.data_mem[3][5] ),
    .S1(_06161_),
    .X(_06804_));
 sg13g2_mux4_1 _25492_ (.S0(_06133_),
    .A0(\mem.mem_internal.data_mem[4][5] ),
    .A1(\mem.mem_internal.data_mem[5][5] ),
    .A2(\mem.mem_internal.data_mem[6][5] ),
    .A3(\mem.mem_internal.data_mem[7][5] ),
    .S1(_06139_),
    .X(_06805_));
 sg13g2_mux4_1 _25493_ (.S0(net577),
    .A0(\mem.mem_internal.data_mem[8][5] ),
    .A1(\mem.mem_internal.data_mem[9][5] ),
    .A2(\mem.mem_internal.data_mem[10][5] ),
    .A3(\mem.mem_internal.data_mem[11][5] ),
    .S1(net543),
    .X(_06806_));
 sg13g2_mux4_1 _25494_ (.S0(net542),
    .A0(\mem.mem_internal.data_mem[12][5] ),
    .A1(\mem.mem_internal.data_mem[13][5] ),
    .A2(\mem.mem_internal.data_mem[14][5] ),
    .A3(\mem.mem_internal.data_mem[15][5] ),
    .S1(net541),
    .X(_06807_));
 sg13g2_mux4_1 _25495_ (.S0(_06151_),
    .A0(_06804_),
    .A1(_06805_),
    .A2(_06806_),
    .A3(_06807_),
    .S1(_06170_),
    .X(_06808_));
 sg13g2_mux4_1 _25496_ (.S0(net540),
    .A0(\mem.mem_internal.data_mem[16][5] ),
    .A1(\mem.mem_internal.data_mem[17][5] ),
    .A2(\mem.mem_internal.data_mem[18][5] ),
    .A3(\mem.mem_internal.data_mem[19][5] ),
    .S1(net539),
    .X(_06809_));
 sg13g2_mux4_1 _25497_ (.S0(net540),
    .A0(\mem.mem_internal.data_mem[20][5] ),
    .A1(\mem.mem_internal.data_mem[21][5] ),
    .A2(\mem.mem_internal.data_mem[22][5] ),
    .A3(\mem.mem_internal.data_mem[23][5] ),
    .S1(net539),
    .X(_06810_));
 sg13g2_mux4_1 _25498_ (.S0(_06132_),
    .A0(\mem.mem_internal.data_mem[24][5] ),
    .A1(\mem.mem_internal.data_mem[25][5] ),
    .A2(\mem.mem_internal.data_mem[26][5] ),
    .A3(\mem.mem_internal.data_mem[27][5] ),
    .S1(net578),
    .X(_06811_));
 sg13g2_mux4_1 _25499_ (.S0(net576),
    .A0(\mem.mem_internal.data_mem[28][5] ),
    .A1(\mem.mem_internal.data_mem[29][5] ),
    .A2(\mem.mem_internal.data_mem[30][5] ),
    .A3(\mem.mem_internal.data_mem[31][5] ),
    .S1(net575),
    .X(_06812_));
 sg13g2_mux4_1 _25500_ (.S0(net988),
    .A0(_06809_),
    .A1(_06810_),
    .A2(_06811_),
    .A3(_06812_),
    .S1(net1235),
    .X(_06813_));
 sg13g2_mux2_1 _25501_ (.A0(_06808_),
    .A1(_06813_),
    .S(_06155_),
    .X(_06814_));
 sg13g2_mux4_1 _25502_ (.S0(net958),
    .A0(\mem.mem_internal.code_mem[0][5] ),
    .A1(\mem.mem_internal.code_mem[1][5] ),
    .A2(\mem.mem_internal.code_mem[2][5] ),
    .A3(\mem.mem_internal.code_mem[3][5] ),
    .S1(net814),
    .X(_06815_));
 sg13g2_mux4_1 _25503_ (.S0(net931),
    .A0(\mem.mem_internal.code_mem[4][5] ),
    .A1(\mem.mem_internal.code_mem[5][5] ),
    .A2(\mem.mem_internal.code_mem[6][5] ),
    .A3(\mem.mem_internal.code_mem[7][5] ),
    .S1(_06322_),
    .X(_06816_));
 sg13g2_mux4_1 _25504_ (.S0(net920),
    .A0(\mem.mem_internal.code_mem[16][5] ),
    .A1(\mem.mem_internal.code_mem[17][5] ),
    .A2(\mem.mem_internal.code_mem[18][5] ),
    .A3(\mem.mem_internal.code_mem[19][5] ),
    .S1(net955),
    .X(_06817_));
 sg13g2_mux4_1 _25505_ (.S0(net954),
    .A0(\mem.mem_internal.code_mem[20][5] ),
    .A1(\mem.mem_internal.code_mem[21][5] ),
    .A2(\mem.mem_internal.code_mem[22][5] ),
    .A3(\mem.mem_internal.code_mem[23][5] ),
    .S1(net953),
    .X(_06818_));
 sg13g2_mux4_1 _25506_ (.S0(net979),
    .A0(_06815_),
    .A1(_06816_),
    .A2(_06817_),
    .A3(_06818_),
    .S1(_06331_),
    .X(_06819_));
 sg13g2_mux4_1 _25507_ (.S0(net931),
    .A0(\mem.mem_internal.code_mem[8][5] ),
    .A1(\mem.mem_internal.code_mem[9][5] ),
    .A2(\mem.mem_internal.code_mem[10][5] ),
    .A3(\mem.mem_internal.code_mem[11][5] ),
    .S1(net812),
    .X(_06820_));
 sg13g2_mux4_1 _25508_ (.S0(net811),
    .A0(\mem.mem_internal.code_mem[12][5] ),
    .A1(\mem.mem_internal.code_mem[13][5] ),
    .A2(\mem.mem_internal.code_mem[14][5] ),
    .A3(\mem.mem_internal.code_mem[15][5] ),
    .S1(net806),
    .X(_06821_));
 sg13g2_mux4_1 _25509_ (.S0(net950),
    .A0(\mem.mem_internal.code_mem[24][5] ),
    .A1(\mem.mem_internal.code_mem[25][5] ),
    .A2(\mem.mem_internal.code_mem[26][5] ),
    .A3(\mem.mem_internal.code_mem[27][5] ),
    .S1(net809),
    .X(_06822_));
 sg13g2_mux4_1 _25510_ (.S0(_06525_),
    .A0(\mem.mem_internal.code_mem[28][5] ),
    .A1(\mem.mem_internal.code_mem[29][5] ),
    .A2(\mem.mem_internal.code_mem[30][5] ),
    .A3(\mem.mem_internal.code_mem[31][5] ),
    .S1(net804),
    .X(_06823_));
 sg13g2_mux4_1 _25511_ (.S0(_06344_),
    .A0(_06820_),
    .A1(_06821_),
    .A2(_06822_),
    .A3(_06823_),
    .S1(net951),
    .X(_06824_));
 sg13g2_mux4_1 _25512_ (.S0(net920),
    .A0(\mem.mem_internal.code_mem[128][5] ),
    .A1(\mem.mem_internal.code_mem[129][5] ),
    .A2(\mem.mem_internal.code_mem[130][5] ),
    .A3(\mem.mem_internal.code_mem[131][5] ),
    .S1(net946),
    .X(_06825_));
 sg13g2_mux4_1 _25513_ (.S0(net930),
    .A0(\mem.mem_internal.code_mem[132][5] ),
    .A1(\mem.mem_internal.code_mem[133][5] ),
    .A2(\mem.mem_internal.code_mem[134][5] ),
    .A3(\mem.mem_internal.code_mem[135][5] ),
    .S1(net808),
    .X(_06826_));
 sg13g2_mux4_1 _25514_ (.S0(net918),
    .A0(\mem.mem_internal.code_mem[144][5] ),
    .A1(\mem.mem_internal.code_mem[145][5] ),
    .A2(\mem.mem_internal.code_mem[146][5] ),
    .A3(\mem.mem_internal.code_mem[147][5] ),
    .S1(net943),
    .X(_06827_));
 sg13g2_mux4_1 _25515_ (.S0(net942),
    .A0(\mem.mem_internal.code_mem[148][5] ),
    .A1(\mem.mem_internal.code_mem[149][5] ),
    .A2(\mem.mem_internal.code_mem[150][5] ),
    .A3(\mem.mem_internal.code_mem[151][5] ),
    .S1(net941),
    .X(_06828_));
 sg13g2_mux4_1 _25516_ (.S0(net940),
    .A0(_06825_),
    .A1(_06826_),
    .A2(_06827_),
    .A3(_06828_),
    .S1(net915),
    .X(_06829_));
 sg13g2_mux4_1 _25517_ (.S0(net938),
    .A0(\mem.mem_internal.code_mem[136][5] ),
    .A1(\mem.mem_internal.code_mem[137][5] ),
    .A2(\mem.mem_internal.code_mem[138][5] ),
    .A3(\mem.mem_internal.code_mem[139][5] ),
    .S1(net899),
    .X(_06830_));
 sg13g2_mux4_1 _25518_ (.S0(net884),
    .A0(\mem.mem_internal.code_mem[140][5] ),
    .A1(\mem.mem_internal.code_mem[141][5] ),
    .A2(\mem.mem_internal.code_mem[142][5] ),
    .A3(\mem.mem_internal.code_mem[143][5] ),
    .S1(net797),
    .X(_06831_));
 sg13g2_mux4_1 _25519_ (.S0(net937),
    .A0(\mem.mem_internal.code_mem[152][5] ),
    .A1(\mem.mem_internal.code_mem[153][5] ),
    .A2(\mem.mem_internal.code_mem[154][5] ),
    .A3(\mem.mem_internal.code_mem[155][5] ),
    .S1(net898),
    .X(_06832_));
 sg13g2_mux4_1 _25520_ (.S0(net935),
    .A0(\mem.mem_internal.code_mem[156][5] ),
    .A1(\mem.mem_internal.code_mem[157][5] ),
    .A2(\mem.mem_internal.code_mem[158][5] ),
    .A3(\mem.mem_internal.code_mem[159][5] ),
    .S1(net934),
    .X(_06833_));
 sg13g2_mux4_1 _25521_ (.S0(net896),
    .A0(_06830_),
    .A1(_06831_),
    .A2(_06832_),
    .A3(_06833_),
    .S1(net932),
    .X(_06834_));
 sg13g2_mux4_1 _25522_ (.S0(_06223_),
    .A0(_06819_),
    .A1(_06824_),
    .A2(_06829_),
    .A3(_06834_),
    .S1(net1233),
    .X(_06835_));
 sg13g2_mux4_1 _25523_ (.S0(net958),
    .A0(\mem.mem_internal.code_mem[32][5] ),
    .A1(\mem.mem_internal.code_mem[33][5] ),
    .A2(\mem.mem_internal.code_mem[34][5] ),
    .A3(\mem.mem_internal.code_mem[35][5] ),
    .S1(net813),
    .X(_06836_));
 sg13g2_mux4_1 _25524_ (.S0(net803),
    .A0(\mem.mem_internal.code_mem[36][5] ),
    .A1(\mem.mem_internal.code_mem[37][5] ),
    .A2(\mem.mem_internal.code_mem[38][5] ),
    .A3(\mem.mem_internal.code_mem[39][5] ),
    .S1(net806),
    .X(_06837_));
 sg13g2_mux4_1 _25525_ (.S0(net930),
    .A0(\mem.mem_internal.code_mem[48][5] ),
    .A1(\mem.mem_internal.code_mem[49][5] ),
    .A2(\mem.mem_internal.code_mem[50][5] ),
    .A3(\mem.mem_internal.code_mem[51][5] ),
    .S1(net805),
    .X(_06838_));
 sg13g2_mux4_1 _25526_ (.S0(net929),
    .A0(\mem.mem_internal.code_mem[52][5] ),
    .A1(\mem.mem_internal.code_mem[53][5] ),
    .A2(\mem.mem_internal.code_mem[54][5] ),
    .A3(\mem.mem_internal.code_mem[55][5] ),
    .S1(net804),
    .X(_06839_));
 sg13g2_mux4_1 _25527_ (.S0(net952),
    .A0(_06836_),
    .A1(_06837_),
    .A2(_06838_),
    .A3(_06839_),
    .S1(net947),
    .X(_06840_));
 sg13g2_mux4_1 _25528_ (.S0(_06389_),
    .A0(\mem.mem_internal.code_mem[40][5] ),
    .A1(\mem.mem_internal.code_mem[41][5] ),
    .A2(\mem.mem_internal.code_mem[42][5] ),
    .A3(\mem.mem_internal.code_mem[43][5] ),
    .S1(net810),
    .X(_06841_));
 sg13g2_mux4_1 _25529_ (.S0(net820),
    .A0(\mem.mem_internal.code_mem[44][5] ),
    .A1(\mem.mem_internal.code_mem[45][5] ),
    .A2(\mem.mem_internal.code_mem[46][5] ),
    .A3(\mem.mem_internal.code_mem[47][5] ),
    .S1(net819),
    .X(_06842_));
 sg13g2_mux4_1 _25530_ (.S0(_06392_),
    .A0(\mem.mem_internal.code_mem[56][5] ),
    .A1(\mem.mem_internal.code_mem[57][5] ),
    .A2(\mem.mem_internal.code_mem[58][5] ),
    .A3(\mem.mem_internal.code_mem[59][5] ),
    .S1(net801),
    .X(_06843_));
 sg13g2_mux4_1 _25531_ (.S0(_06395_),
    .A0(\mem.mem_internal.code_mem[60][5] ),
    .A1(\mem.mem_internal.code_mem[61][5] ),
    .A2(\mem.mem_internal.code_mem[62][5] ),
    .A3(\mem.mem_internal.code_mem[63][5] ),
    .S1(net815),
    .X(_06844_));
 sg13g2_mux4_1 _25532_ (.S0(net948),
    .A0(_06841_),
    .A1(_06842_),
    .A2(_06843_),
    .A3(_06844_),
    .S1(net987),
    .X(_06845_));
 sg13g2_mux4_1 _25533_ (.S0(net945),
    .A0(\mem.mem_internal.code_mem[160][5] ),
    .A1(\mem.mem_internal.code_mem[161][5] ),
    .A2(\mem.mem_internal.code_mem[162][5] ),
    .A3(\mem.mem_internal.code_mem[163][5] ),
    .S1(net805),
    .X(_06846_));
 sg13g2_mux4_1 _25534_ (.S0(net928),
    .A0(\mem.mem_internal.code_mem[164][5] ),
    .A1(\mem.mem_internal.code_mem[165][5] ),
    .A2(\mem.mem_internal.code_mem[166][5] ),
    .A3(\mem.mem_internal.code_mem[167][5] ),
    .S1(net801),
    .X(_06847_));
 sg13g2_mux4_1 _25535_ (.S0(net925),
    .A0(\mem.mem_internal.code_mem[176][5] ),
    .A1(\mem.mem_internal.code_mem[177][5] ),
    .A2(\mem.mem_internal.code_mem[178][5] ),
    .A3(\mem.mem_internal.code_mem[179][5] ),
    .S1(net924),
    .X(_06848_));
 sg13g2_mux4_1 _25536_ (.S0(net962),
    .A0(\mem.mem_internal.code_mem[180][5] ),
    .A1(\mem.mem_internal.code_mem[181][5] ),
    .A2(\mem.mem_internal.code_mem[182][5] ),
    .A3(\mem.mem_internal.code_mem[183][5] ),
    .S1(net912),
    .X(_06849_));
 sg13g2_mux4_1 _25537_ (.S0(net923),
    .A0(_06846_),
    .A1(_06847_),
    .A2(_06848_),
    .A3(_06849_),
    .S1(net911),
    .X(_06850_));
 sg13g2_mux4_1 _25538_ (.S0(net949),
    .A0(\mem.mem_internal.code_mem[168][5] ),
    .A1(\mem.mem_internal.code_mem[169][5] ),
    .A2(\mem.mem_internal.code_mem[170][5] ),
    .A3(\mem.mem_internal.code_mem[171][5] ),
    .S1(net807),
    .X(_06851_));
 sg13g2_mux4_1 _25539_ (.S0(net927),
    .A0(\mem.mem_internal.code_mem[172][5] ),
    .A1(\mem.mem_internal.code_mem[173][5] ),
    .A2(\mem.mem_internal.code_mem[174][5] ),
    .A3(\mem.mem_internal.code_mem[175][5] ),
    .S1(net800),
    .X(_06852_));
 sg13g2_mux4_1 _25540_ (.S0(net894),
    .A0(\mem.mem_internal.code_mem[184][5] ),
    .A1(\mem.mem_internal.code_mem[185][5] ),
    .A2(\mem.mem_internal.code_mem[186][5] ),
    .A3(\mem.mem_internal.code_mem[187][5] ),
    .S1(net921),
    .X(_06853_));
 sg13g2_mux4_1 _25541_ (.S0(net893),
    .A0(\mem.mem_internal.code_mem[188][5] ),
    .A1(\mem.mem_internal.code_mem[189][5] ),
    .A2(\mem.mem_internal.code_mem[190][5] ),
    .A3(\mem.mem_internal.code_mem[191][5] ),
    .S1(net980),
    .X(_06854_));
 sg13g2_mux4_1 _25542_ (.S0(net891),
    .A0(_06851_),
    .A1(_06852_),
    .A2(_06853_),
    .A3(_06854_),
    .S1(net978),
    .X(_06855_));
 sg13g2_mux4_1 _25543_ (.S0(net1235),
    .A0(_06840_),
    .A1(_06845_),
    .A2(_06850_),
    .A3(_06855_),
    .S1(net1232),
    .X(_06856_));
 sg13g2_mux4_1 _25544_ (.S0(net965),
    .A0(\mem.mem_internal.code_mem[64][5] ),
    .A1(\mem.mem_internal.code_mem[65][5] ),
    .A2(\mem.mem_internal.code_mem[66][5] ),
    .A3(\mem.mem_internal.code_mem[67][5] ),
    .S1(net966),
    .X(_06857_));
 sg13g2_mux4_1 _25545_ (.S0(_06419_),
    .A0(\mem.mem_internal.code_mem[68][5] ),
    .A1(\mem.mem_internal.code_mem[69][5] ),
    .A2(\mem.mem_internal.code_mem[70][5] ),
    .A3(\mem.mem_internal.code_mem[71][5] ),
    .S1(net799),
    .X(_06858_));
 sg13g2_mux4_1 _25546_ (.S0(net963),
    .A0(\mem.mem_internal.code_mem[80][5] ),
    .A1(\mem.mem_internal.code_mem[81][5] ),
    .A2(\mem.mem_internal.code_mem[82][5] ),
    .A3(\mem.mem_internal.code_mem[83][5] ),
    .S1(net964),
    .X(_06859_));
 sg13g2_mux4_1 _25547_ (.S0(net916),
    .A0(\mem.mem_internal.code_mem[84][5] ),
    .A1(\mem.mem_internal.code_mem[85][5] ),
    .A2(\mem.mem_internal.code_mem[86][5] ),
    .A3(\mem.mem_internal.code_mem[87][5] ),
    .S1(net936),
    .X(_06860_));
 sg13g2_mux4_1 _25548_ (.S0(net967),
    .A0(_06857_),
    .A1(_06858_),
    .A2(_06859_),
    .A3(_06860_),
    .S1(_06427_),
    .X(_06861_));
 sg13g2_mux4_1 _25549_ (.S0(net938),
    .A0(\mem.mem_internal.code_mem[72][5] ),
    .A1(\mem.mem_internal.code_mem[73][5] ),
    .A2(\mem.mem_internal.code_mem[74][5] ),
    .A3(\mem.mem_internal.code_mem[75][5] ),
    .S1(net799),
    .X(_06862_));
 sg13g2_mux4_1 _25550_ (.S0(net985),
    .A0(\mem.mem_internal.code_mem[76][5] ),
    .A1(\mem.mem_internal.code_mem[77][5] ),
    .A2(\mem.mem_internal.code_mem[78][5] ),
    .A3(\mem.mem_internal.code_mem[79][5] ),
    .S1(net816),
    .X(_06863_));
 sg13g2_mux4_1 _25551_ (.S0(net914),
    .A0(\mem.mem_internal.code_mem[88][5] ),
    .A1(\mem.mem_internal.code_mem[89][5] ),
    .A2(\mem.mem_internal.code_mem[90][5] ),
    .A3(\mem.mem_internal.code_mem[91][5] ),
    .S1(net910),
    .X(_06864_));
 sg13g2_mux4_1 _25552_ (.S0(net890),
    .A0(\mem.mem_internal.code_mem[92][5] ),
    .A1(\mem.mem_internal.code_mem[93][5] ),
    .A2(\mem.mem_internal.code_mem[94][5] ),
    .A3(\mem.mem_internal.code_mem[95][5] ),
    .S1(net921),
    .X(_06865_));
 sg13g2_mux4_1 _25553_ (.S0(net933),
    .A0(_06862_),
    .A1(_06863_),
    .A2(_06864_),
    .A3(_06865_),
    .S1(net932),
    .X(_06866_));
 sg13g2_mux4_1 _25554_ (.S0(net963),
    .A0(\mem.mem_internal.code_mem[192][5] ),
    .A1(\mem.mem_internal.code_mem[193][5] ),
    .A2(\mem.mem_internal.code_mem[194][5] ),
    .A3(\mem.mem_internal.code_mem[195][5] ),
    .S1(net917),
    .X(_06867_));
 sg13g2_mux4_1 _25555_ (.S0(net942),
    .A0(\mem.mem_internal.code_mem[196][5] ),
    .A1(\mem.mem_internal.code_mem[197][5] ),
    .A2(\mem.mem_internal.code_mem[198][5] ),
    .A3(\mem.mem_internal.code_mem[199][5] ),
    .S1(net941),
    .X(_06868_));
 sg13g2_mux4_1 _25556_ (.S0(net959),
    .A0(\mem.mem_internal.code_mem[208][5] ),
    .A1(\mem.mem_internal.code_mem[209][5] ),
    .A2(\mem.mem_internal.code_mem[210][5] ),
    .A3(\mem.mem_internal.code_mem[211][5] ),
    .S1(net961),
    .X(_06869_));
 sg13g2_mux4_1 _25557_ (.S0(net908),
    .A0(\mem.mem_internal.code_mem[212][5] ),
    .A1(\mem.mem_internal.code_mem[213][5] ),
    .A2(\mem.mem_internal.code_mem[214][5] ),
    .A3(\mem.mem_internal.code_mem[215][5] ),
    .S1(net888),
    .X(_06870_));
 sg13g2_mux4_1 _25558_ (.S0(net1231),
    .A0(_06867_),
    .A1(_06868_),
    .A2(_06869_),
    .A3(_06870_),
    .S1(net960),
    .X(_06871_));
 sg13g2_mux4_1 _25559_ (.S0(net916),
    .A0(\mem.mem_internal.code_mem[200][5] ),
    .A1(\mem.mem_internal.code_mem[201][5] ),
    .A2(\mem.mem_internal.code_mem[202][5] ),
    .A3(\mem.mem_internal.code_mem[203][5] ),
    .S1(net905),
    .X(_06872_));
 sg13g2_mux4_1 _25560_ (.S0(net890),
    .A0(\mem.mem_internal.code_mem[204][5] ),
    .A1(\mem.mem_internal.code_mem[205][5] ),
    .A2(\mem.mem_internal.code_mem[206][5] ),
    .A3(\mem.mem_internal.code_mem[207][5] ),
    .S1(net889),
    .X(_06873_));
 sg13g2_mux4_1 _25561_ (.S0(_06453_),
    .A0(\mem.mem_internal.code_mem[216][5] ),
    .A1(\mem.mem_internal.code_mem[217][5] ),
    .A2(\mem.mem_internal.code_mem[218][5] ),
    .A3(\mem.mem_internal.code_mem[219][5] ),
    .S1(net909),
    .X(_06874_));
 sg13g2_mux4_1 _25562_ (.S0(net885),
    .A0(\mem.mem_internal.code_mem[220][5] ),
    .A1(\mem.mem_internal.code_mem[221][5] ),
    .A2(\mem.mem_internal.code_mem[222][5] ),
    .A3(\mem.mem_internal.code_mem[223][5] ),
    .S1(_06456_),
    .X(_06875_));
 sg13g2_mux4_1 _25563_ (.S0(net1230),
    .A0(_06872_),
    .A1(_06873_),
    .A2(_06874_),
    .A3(_06875_),
    .S1(net887),
    .X(_06876_));
 sg13g2_mux4_1 _25564_ (.S0(_06168_),
    .A0(_06861_),
    .A1(_06866_),
    .A2(_06871_),
    .A3(_06876_),
    .S1(net1228),
    .X(_06877_));
 sg13g2_mux4_1 _25565_ (.S0(net956),
    .A0(\mem.mem_internal.code_mem[96][5] ),
    .A1(\mem.mem_internal.code_mem[97][5] ),
    .A2(\mem.mem_internal.code_mem[98][5] ),
    .A3(\mem.mem_internal.code_mem[99][5] ),
    .S1(net946),
    .X(_06878_));
 sg13g2_mux4_1 _25566_ (.S0(net895),
    .A0(\mem.mem_internal.code_mem[100][5] ),
    .A1(\mem.mem_internal.code_mem[101][5] ),
    .A2(\mem.mem_internal.code_mem[102][5] ),
    .A3(\mem.mem_internal.code_mem[103][5] ),
    .S1(net798),
    .X(_06879_));
 sg13g2_mux4_1 _25567_ (.S0(net906),
    .A0(\mem.mem_internal.code_mem[112][5] ),
    .A1(\mem.mem_internal.code_mem[113][5] ),
    .A2(\mem.mem_internal.code_mem[114][5] ),
    .A3(\mem.mem_internal.code_mem[115][5] ),
    .S1(_06468_),
    .X(_06880_));
 sg13g2_mux4_1 _25568_ (.S0(net897),
    .A0(\mem.mem_internal.code_mem[116][5] ),
    .A1(\mem.mem_internal.code_mem[117][5] ),
    .A2(\mem.mem_internal.code_mem[118][5] ),
    .A3(\mem.mem_internal.code_mem[119][5] ),
    .S1(net886),
    .X(_06881_));
 sg13g2_mux4_1 _25569_ (.S0(_06472_),
    .A0(_06878_),
    .A1(_06879_),
    .A2(_06880_),
    .A3(_06881_),
    .S1(net939),
    .X(_06882_));
 sg13g2_mux4_1 _25570_ (.S0(net895),
    .A0(\mem.mem_internal.code_mem[104][5] ),
    .A1(\mem.mem_internal.code_mem[105][5] ),
    .A2(\mem.mem_internal.code_mem[106][5] ),
    .A3(\mem.mem_internal.code_mem[107][5] ),
    .S1(net798),
    .X(_06883_));
 sg13g2_mux4_1 _25571_ (.S0(net926),
    .A0(\mem.mem_internal.code_mem[108][5] ),
    .A1(\mem.mem_internal.code_mem[109][5] ),
    .A2(\mem.mem_internal.code_mem[110][5] ),
    .A3(\mem.mem_internal.code_mem[111][5] ),
    .S1(net802),
    .X(_06884_));
 sg13g2_mux4_1 _25572_ (.S0(_06478_),
    .A0(\mem.mem_internal.code_mem[120][5] ),
    .A1(\mem.mem_internal.code_mem[121][5] ),
    .A2(\mem.mem_internal.code_mem[122][5] ),
    .A3(\mem.mem_internal.code_mem[123][5] ),
    .S1(net904),
    .X(_06885_));
 sg13g2_mux4_1 _25573_ (.S0(_06480_),
    .A0(\mem.mem_internal.code_mem[124][5] ),
    .A1(\mem.mem_internal.code_mem[125][5] ),
    .A2(\mem.mem_internal.code_mem[126][5] ),
    .A3(\mem.mem_internal.code_mem[127][5] ),
    .S1(net892),
    .X(_06886_));
 sg13g2_mux4_1 _25574_ (.S0(net923),
    .A0(_06883_),
    .A1(_06884_),
    .A2(_06885_),
    .A3(_06886_),
    .S1(net922),
    .X(_06887_));
 sg13g2_mux4_1 _25575_ (.S0(net944),
    .A0(\mem.mem_internal.code_mem[224][5] ),
    .A1(\mem.mem_internal.code_mem[225][5] ),
    .A2(\mem.mem_internal.code_mem[226][5] ),
    .A3(\mem.mem_internal.code_mem[227][5] ),
    .S1(net943),
    .X(_06888_));
 sg13g2_mux4_1 _25576_ (.S0(net935),
    .A0(\mem.mem_internal.code_mem[228][5] ),
    .A1(\mem.mem_internal.code_mem[229][5] ),
    .A2(\mem.mem_internal.code_mem[230][5] ),
    .A3(\mem.mem_internal.code_mem[231][5] ),
    .S1(_06487_),
    .X(_06889_));
 sg13g2_mux4_1 _25577_ (.S0(net903),
    .A0(\mem.mem_internal.code_mem[240][5] ),
    .A1(\mem.mem_internal.code_mem[241][5] ),
    .A2(\mem.mem_internal.code_mem[242][5] ),
    .A3(\mem.mem_internal.code_mem[243][5] ),
    .S1(net888),
    .X(_06890_));
 sg13g2_mux4_1 _25578_ (.S0(net902),
    .A0(\mem.mem_internal.code_mem[244][5] ),
    .A1(\mem.mem_internal.code_mem[245][5] ),
    .A2(\mem.mem_internal.code_mem[246][5] ),
    .A3(\mem.mem_internal.code_mem[247][5] ),
    .S1(net901),
    .X(_06891_));
 sg13g2_mux4_1 _25579_ (.S0(net1231),
    .A0(_06888_),
    .A1(_06889_),
    .A2(_06890_),
    .A3(_06891_),
    .S1(net887),
    .X(_06892_));
 sg13g2_mux4_1 _25580_ (.S0(net925),
    .A0(\mem.mem_internal.code_mem[232][5] ),
    .A1(\mem.mem_internal.code_mem[233][5] ),
    .A2(\mem.mem_internal.code_mem[234][5] ),
    .A3(\mem.mem_internal.code_mem[235][5] ),
    .S1(_06494_),
    .X(_06893_));
 sg13g2_mux4_1 _25581_ (.S0(net983),
    .A0(\mem.mem_internal.code_mem[236][5] ),
    .A1(\mem.mem_internal.code_mem[237][5] ),
    .A2(\mem.mem_internal.code_mem[238][5] ),
    .A3(\mem.mem_internal.code_mem[239][5] ),
    .S1(net982),
    .X(_06894_));
 sg13g2_mux4_1 _25582_ (.S0(net885),
    .A0(\mem.mem_internal.code_mem[248][5] ),
    .A1(\mem.mem_internal.code_mem[249][5] ),
    .A2(\mem.mem_internal.code_mem[250][5] ),
    .A3(\mem.mem_internal.code_mem[251][5] ),
    .S1(net907),
    .X(_06895_));
 sg13g2_mux4_1 _25583_ (.S0(net975),
    .A0(\mem.mem_internal.code_mem[252][5] ),
    .A1(\mem.mem_internal.code_mem[253][5] ),
    .A2(\mem.mem_internal.code_mem[254][5] ),
    .A3(\mem.mem_internal.code_mem[255][5] ),
    .S1(net974),
    .X(_06896_));
 sg13g2_mux4_1 _25584_ (.S0(net971),
    .A0(_06893_),
    .A1(_06894_),
    .A2(_06895_),
    .A3(_06896_),
    .S1(net900),
    .X(_06897_));
 sg13g2_mux4_1 _25585_ (.S0(net1229),
    .A0(_06882_),
    .A1(_06887_),
    .A2(_06892_),
    .A3(_06897_),
    .S1(net1228),
    .X(_06898_));
 sg13g2_mux4_1 _25586_ (.S0(_06300_),
    .A0(_06835_),
    .A1(_06856_),
    .A2(_06877_),
    .A3(_06898_),
    .S1(_06301_),
    .X(_06899_));
 sg13g2_nor2_1 _25587_ (.A(_06304_),
    .B(_06899_),
    .Y(_06900_));
 sg13g2_a21oi_1 _25588_ (.A1(net832),
    .A2(_06814_),
    .Y(_06901_),
    .B1(_06900_));
 sg13g2_nand2_1 _25589_ (.Y(_06902_),
    .A(\mem.internal_data_out[5] ),
    .B(_06126_));
 sg13g2_o21ai_1 _25590_ (.B1(_06902_),
    .Y(_02425_),
    .A1(net546),
    .A2(_06901_));
 sg13g2_mux4_1 _25591_ (.S0(net538),
    .A0(\mem.mem_internal.data_mem[0][6] ),
    .A1(\mem.mem_internal.data_mem[1][6] ),
    .A2(\mem.mem_internal.data_mem[2][6] ),
    .A3(\mem.mem_internal.data_mem[3][6] ),
    .S1(net537),
    .X(_06903_));
 sg13g2_mux4_1 _25592_ (.S0(_06133_),
    .A0(\mem.mem_internal.data_mem[4][6] ),
    .A1(\mem.mem_internal.data_mem[5][6] ),
    .A2(\mem.mem_internal.data_mem[6][6] ),
    .A3(\mem.mem_internal.data_mem[7][6] ),
    .S1(_06139_),
    .X(_06904_));
 sg13g2_mux4_1 _25593_ (.S0(_06142_),
    .A0(\mem.mem_internal.data_mem[16][6] ),
    .A1(\mem.mem_internal.data_mem[17][6] ),
    .A2(\mem.mem_internal.data_mem[18][6] ),
    .A3(\mem.mem_internal.data_mem[19][6] ),
    .S1(_06143_),
    .X(_06905_));
 sg13g2_mux4_1 _25594_ (.S0(net542),
    .A0(\mem.mem_internal.data_mem[20][6] ),
    .A1(\mem.mem_internal.data_mem[21][6] ),
    .A2(\mem.mem_internal.data_mem[22][6] ),
    .A3(\mem.mem_internal.data_mem[23][6] ),
    .S1(net541),
    .X(_06906_));
 sg13g2_mux4_1 _25595_ (.S0(net818),
    .A0(_06903_),
    .A1(_06904_),
    .A2(_06905_),
    .A3(_06906_),
    .S1(net817),
    .X(_06907_));
 sg13g2_mux4_1 _25596_ (.S0(_06145_),
    .A0(\mem.mem_internal.data_mem[8][6] ),
    .A1(\mem.mem_internal.data_mem[9][6] ),
    .A2(\mem.mem_internal.data_mem[10][6] ),
    .A3(\mem.mem_internal.data_mem[11][6] ),
    .S1(_06146_),
    .X(_06908_));
 sg13g2_mux4_1 _25597_ (.S0(_06157_),
    .A0(\mem.mem_internal.data_mem[12][6] ),
    .A1(\mem.mem_internal.data_mem[13][6] ),
    .A2(\mem.mem_internal.data_mem[14][6] ),
    .A3(\mem.mem_internal.data_mem[15][6] ),
    .S1(_06158_),
    .X(_06909_));
 sg13g2_mux4_1 _25598_ (.S0(_06132_),
    .A0(\mem.mem_internal.data_mem[24][6] ),
    .A1(\mem.mem_internal.data_mem[25][6] ),
    .A2(\mem.mem_internal.data_mem[26][6] ),
    .A3(\mem.mem_internal.data_mem[27][6] ),
    .S1(net578),
    .X(_06910_));
 sg13g2_mux4_1 _25599_ (.S0(net576),
    .A0(\mem.mem_internal.data_mem[28][6] ),
    .A1(\mem.mem_internal.data_mem[29][6] ),
    .A2(\mem.mem_internal.data_mem[30][6] ),
    .A3(\mem.mem_internal.data_mem[31][6] ),
    .S1(net575),
    .X(_06911_));
 sg13g2_mux4_1 _25600_ (.S0(net988),
    .A0(_06908_),
    .A1(_06909_),
    .A2(_06910_),
    .A3(_06911_),
    .S1(net987),
    .X(_06912_));
 sg13g2_mux2_1 _25601_ (.A0(_06907_),
    .A1(_06912_),
    .S(net986),
    .X(_06913_));
 sg13g2_mux4_1 _25602_ (.S0(_06319_),
    .A0(\mem.mem_internal.code_mem[0][6] ),
    .A1(\mem.mem_internal.code_mem[1][6] ),
    .A2(\mem.mem_internal.code_mem[2][6] ),
    .A3(\mem.mem_internal.code_mem[3][6] ),
    .S1(_06232_),
    .X(_06914_));
 sg13g2_mux4_1 _25603_ (.S0(net931),
    .A0(\mem.mem_internal.code_mem[4][6] ),
    .A1(\mem.mem_internal.code_mem[5][6] ),
    .A2(\mem.mem_internal.code_mem[6][6] ),
    .A3(\mem.mem_internal.code_mem[7][6] ),
    .S1(_06322_),
    .X(_06915_));
 sg13g2_mux4_1 _25604_ (.S0(net920),
    .A0(\mem.mem_internal.code_mem[16][6] ),
    .A1(\mem.mem_internal.code_mem[17][6] ),
    .A2(\mem.mem_internal.code_mem[18][6] ),
    .A3(\mem.mem_internal.code_mem[19][6] ),
    .S1(net955),
    .X(_06916_));
 sg13g2_mux4_1 _25605_ (.S0(net954),
    .A0(\mem.mem_internal.code_mem[20][6] ),
    .A1(\mem.mem_internal.code_mem[21][6] ),
    .A2(\mem.mem_internal.code_mem[22][6] ),
    .A3(\mem.mem_internal.code_mem[23][6] ),
    .S1(_06328_),
    .X(_06917_));
 sg13g2_mux4_1 _25606_ (.S0(_06190_),
    .A0(_06914_),
    .A1(_06915_),
    .A2(_06916_),
    .A3(_06917_),
    .S1(_06331_),
    .X(_06918_));
 sg13g2_mux4_1 _25607_ (.S0(_06378_),
    .A0(\mem.mem_internal.code_mem[8][6] ),
    .A1(\mem.mem_internal.code_mem[9][6] ),
    .A2(\mem.mem_internal.code_mem[10][6] ),
    .A3(\mem.mem_internal.code_mem[11][6] ),
    .S1(_06333_),
    .X(_06919_));
 sg13g2_mux4_1 _25608_ (.S0(_06335_),
    .A0(\mem.mem_internal.code_mem[12][6] ),
    .A1(\mem.mem_internal.code_mem[13][6] ),
    .A2(\mem.mem_internal.code_mem[14][6] ),
    .A3(\mem.mem_internal.code_mem[15][6] ),
    .S1(_06380_),
    .X(_06920_));
 sg13g2_mux4_1 _25609_ (.S0(net950),
    .A0(\mem.mem_internal.code_mem[24][6] ),
    .A1(\mem.mem_internal.code_mem[25][6] ),
    .A2(\mem.mem_internal.code_mem[26][6] ),
    .A3(\mem.mem_internal.code_mem[27][6] ),
    .S1(_06340_),
    .X(_06921_));
 sg13g2_mux4_1 _25610_ (.S0(_06525_),
    .A0(\mem.mem_internal.code_mem[28][6] ),
    .A1(\mem.mem_internal.code_mem[29][6] ),
    .A2(\mem.mem_internal.code_mem[30][6] ),
    .A3(\mem.mem_internal.code_mem[31][6] ),
    .S1(_06386_),
    .X(_06922_));
 sg13g2_mux4_1 _25611_ (.S0(_06344_),
    .A0(_06919_),
    .A1(_06920_),
    .A2(_06921_),
    .A3(_06922_),
    .S1(net951),
    .X(_06923_));
 sg13g2_mux4_1 _25612_ (.S0(_06417_),
    .A0(\mem.mem_internal.code_mem[128][6] ),
    .A1(\mem.mem_internal.code_mem[129][6] ),
    .A2(\mem.mem_internal.code_mem[130][6] ),
    .A3(\mem.mem_internal.code_mem[131][6] ),
    .S1(net946),
    .X(_06924_));
 sg13g2_mux4_1 _25613_ (.S0(_06382_),
    .A0(\mem.mem_internal.code_mem[132][6] ),
    .A1(\mem.mem_internal.code_mem[133][6] ),
    .A2(\mem.mem_internal.code_mem[134][6] ),
    .A3(\mem.mem_internal.code_mem[135][6] ),
    .S1(net808),
    .X(_06925_));
 sg13g2_mux4_1 _25614_ (.S0(net918),
    .A0(\mem.mem_internal.code_mem[144][6] ),
    .A1(\mem.mem_internal.code_mem[145][6] ),
    .A2(\mem.mem_internal.code_mem[146][6] ),
    .A3(\mem.mem_internal.code_mem[147][6] ),
    .S1(net917),
    .X(_06926_));
 sg13g2_mux4_1 _25615_ (.S0(_06367_),
    .A0(\mem.mem_internal.code_mem[148][6] ),
    .A1(\mem.mem_internal.code_mem[149][6] ),
    .A2(\mem.mem_internal.code_mem[150][6] ),
    .A3(\mem.mem_internal.code_mem[151][6] ),
    .S1(net941),
    .X(_06927_));
 sg13g2_mux4_1 _25616_ (.S0(net940),
    .A0(_06924_),
    .A1(_06925_),
    .A2(_06926_),
    .A3(_06927_),
    .S1(net915),
    .X(_06928_));
 sg13g2_mux4_1 _25617_ (.S0(net938),
    .A0(\mem.mem_internal.code_mem[136][6] ),
    .A1(\mem.mem_internal.code_mem[137][6] ),
    .A2(\mem.mem_internal.code_mem[138][6] ),
    .A3(\mem.mem_internal.code_mem[139][6] ),
    .S1(net899),
    .X(_06929_));
 sg13g2_mux4_1 _25618_ (.S0(net884),
    .A0(\mem.mem_internal.code_mem[140][6] ),
    .A1(\mem.mem_internal.code_mem[141][6] ),
    .A2(\mem.mem_internal.code_mem[142][6] ),
    .A3(\mem.mem_internal.code_mem[143][6] ),
    .S1(net797),
    .X(_06930_));
 sg13g2_mux4_1 _25619_ (.S0(net937),
    .A0(\mem.mem_internal.code_mem[152][6] ),
    .A1(\mem.mem_internal.code_mem[153][6] ),
    .A2(\mem.mem_internal.code_mem[154][6] ),
    .A3(\mem.mem_internal.code_mem[155][6] ),
    .S1(net898),
    .X(_06931_));
 sg13g2_mux4_1 _25620_ (.S0(net935),
    .A0(\mem.mem_internal.code_mem[156][6] ),
    .A1(\mem.mem_internal.code_mem[157][6] ),
    .A2(\mem.mem_internal.code_mem[158][6] ),
    .A3(\mem.mem_internal.code_mem[159][6] ),
    .S1(net934),
    .X(_06932_));
 sg13g2_mux4_1 _25621_ (.S0(net896),
    .A0(_06929_),
    .A1(_06930_),
    .A2(_06931_),
    .A3(_06932_),
    .S1(net932),
    .X(_06933_));
 sg13g2_mux4_1 _25622_ (.S0(_06223_),
    .A0(_06918_),
    .A1(_06923_),
    .A2(_06928_),
    .A3(_06933_),
    .S1(_06225_),
    .X(_06934_));
 sg13g2_mux4_1 _25623_ (.S0(net958),
    .A0(\mem.mem_internal.code_mem[32][6] ),
    .A1(\mem.mem_internal.code_mem[33][6] ),
    .A2(\mem.mem_internal.code_mem[34][6] ),
    .A3(\mem.mem_internal.code_mem[35][6] ),
    .S1(net813),
    .X(_06935_));
 sg13g2_mux4_1 _25624_ (.S0(net803),
    .A0(\mem.mem_internal.code_mem[36][6] ),
    .A1(\mem.mem_internal.code_mem[37][6] ),
    .A2(\mem.mem_internal.code_mem[38][6] ),
    .A3(\mem.mem_internal.code_mem[39][6] ),
    .S1(net806),
    .X(_06936_));
 sg13g2_mux4_1 _25625_ (.S0(net930),
    .A0(\mem.mem_internal.code_mem[48][6] ),
    .A1(\mem.mem_internal.code_mem[49][6] ),
    .A2(\mem.mem_internal.code_mem[50][6] ),
    .A3(\mem.mem_internal.code_mem[51][6] ),
    .S1(net805),
    .X(_06937_));
 sg13g2_mux4_1 _25626_ (.S0(net929),
    .A0(\mem.mem_internal.code_mem[52][6] ),
    .A1(\mem.mem_internal.code_mem[53][6] ),
    .A2(\mem.mem_internal.code_mem[54][6] ),
    .A3(\mem.mem_internal.code_mem[55][6] ),
    .S1(net807),
    .X(_06938_));
 sg13g2_mux4_1 _25627_ (.S0(net952),
    .A0(_06935_),
    .A1(_06936_),
    .A2(_06937_),
    .A3(_06938_),
    .S1(net947),
    .X(_06939_));
 sg13g2_mux4_1 _25628_ (.S0(net957),
    .A0(\mem.mem_internal.code_mem[40][6] ),
    .A1(\mem.mem_internal.code_mem[41][6] ),
    .A2(\mem.mem_internal.code_mem[42][6] ),
    .A3(\mem.mem_internal.code_mem[43][6] ),
    .S1(net810),
    .X(_06940_));
 sg13g2_mux4_1 _25629_ (.S0(_06131_),
    .A0(\mem.mem_internal.code_mem[44][6] ),
    .A1(\mem.mem_internal.code_mem[45][6] ),
    .A2(\mem.mem_internal.code_mem[46][6] ),
    .A3(\mem.mem_internal.code_mem[47][6] ),
    .S1(_06137_),
    .X(_06941_));
 sg13g2_mux4_1 _25630_ (.S0(net985),
    .A0(\mem.mem_internal.code_mem[56][6] ),
    .A1(\mem.mem_internal.code_mem[57][6] ),
    .A2(\mem.mem_internal.code_mem[58][6] ),
    .A3(\mem.mem_internal.code_mem[59][6] ),
    .S1(_06400_),
    .X(_06942_));
 sg13g2_mux4_1 _25631_ (.S0(_06395_),
    .A0(\mem.mem_internal.code_mem[60][6] ),
    .A1(\mem.mem_internal.code_mem[61][6] ),
    .A2(\mem.mem_internal.code_mem[62][6] ),
    .A3(\mem.mem_internal.code_mem[63][6] ),
    .S1(net800),
    .X(_06943_));
 sg13g2_mux4_1 _25632_ (.S0(net948),
    .A0(_06940_),
    .A1(_06941_),
    .A2(_06942_),
    .A3(_06943_),
    .S1(_06154_),
    .X(_06944_));
 sg13g2_mux4_1 _25633_ (.S0(net945),
    .A0(\mem.mem_internal.code_mem[160][6] ),
    .A1(\mem.mem_internal.code_mem[161][6] ),
    .A2(\mem.mem_internal.code_mem[162][6] ),
    .A3(\mem.mem_internal.code_mem[163][6] ),
    .S1(_06383_),
    .X(_06945_));
 sg13g2_mux4_1 _25634_ (.S0(net928),
    .A0(\mem.mem_internal.code_mem[164][6] ),
    .A1(\mem.mem_internal.code_mem[165][6] ),
    .A2(\mem.mem_internal.code_mem[166][6] ),
    .A3(\mem.mem_internal.code_mem[167][6] ),
    .S1(net801),
    .X(_06946_));
 sg13g2_mux4_1 _25635_ (.S0(net925),
    .A0(\mem.mem_internal.code_mem[176][6] ),
    .A1(\mem.mem_internal.code_mem[177][6] ),
    .A2(\mem.mem_internal.code_mem[178][6] ),
    .A3(\mem.mem_internal.code_mem[179][6] ),
    .S1(net924),
    .X(_06947_));
 sg13g2_mux4_1 _25636_ (.S0(net962),
    .A0(\mem.mem_internal.code_mem[180][6] ),
    .A1(\mem.mem_internal.code_mem[181][6] ),
    .A2(\mem.mem_internal.code_mem[182][6] ),
    .A3(\mem.mem_internal.code_mem[183][6] ),
    .S1(net912),
    .X(_06948_));
 sg13g2_mux4_1 _25637_ (.S0(net923),
    .A0(_06945_),
    .A1(_06946_),
    .A2(_06947_),
    .A3(_06948_),
    .S1(net911),
    .X(_06949_));
 sg13g2_mux4_1 _25638_ (.S0(net949),
    .A0(\mem.mem_internal.code_mem[168][6] ),
    .A1(\mem.mem_internal.code_mem[169][6] ),
    .A2(\mem.mem_internal.code_mem[170][6] ),
    .A3(\mem.mem_internal.code_mem[171][6] ),
    .S1(net807),
    .X(_06950_));
 sg13g2_mux4_1 _25639_ (.S0(net927),
    .A0(\mem.mem_internal.code_mem[172][6] ),
    .A1(\mem.mem_internal.code_mem[173][6] ),
    .A2(\mem.mem_internal.code_mem[174][6] ),
    .A3(\mem.mem_internal.code_mem[175][6] ),
    .S1(net800),
    .X(_06951_));
 sg13g2_mux4_1 _25640_ (.S0(net894),
    .A0(\mem.mem_internal.code_mem[184][6] ),
    .A1(\mem.mem_internal.code_mem[185][6] ),
    .A2(\mem.mem_internal.code_mem[186][6] ),
    .A3(\mem.mem_internal.code_mem[187][6] ),
    .S1(net921),
    .X(_06952_));
 sg13g2_mux4_1 _25641_ (.S0(net893),
    .A0(\mem.mem_internal.code_mem[188][6] ),
    .A1(\mem.mem_internal.code_mem[189][6] ),
    .A2(\mem.mem_internal.code_mem[190][6] ),
    .A3(\mem.mem_internal.code_mem[191][6] ),
    .S1(net892),
    .X(_06953_));
 sg13g2_mux4_1 _25642_ (.S0(net891),
    .A0(_06950_),
    .A1(_06951_),
    .A2(_06952_),
    .A3(_06953_),
    .S1(net922),
    .X(_06954_));
 sg13g2_mux4_1 _25643_ (.S0(_06169_),
    .A0(_06939_),
    .A1(_06944_),
    .A2(_06949_),
    .A3(_06954_),
    .S1(net1232),
    .X(_06955_));
 sg13g2_mux4_1 _25644_ (.S0(net965),
    .A0(\mem.mem_internal.code_mem[64][6] ),
    .A1(\mem.mem_internal.code_mem[65][6] ),
    .A2(\mem.mem_internal.code_mem[66][6] ),
    .A3(\mem.mem_internal.code_mem[67][6] ),
    .S1(net966),
    .X(_06956_));
 sg13g2_mux4_1 _25645_ (.S0(net919),
    .A0(\mem.mem_internal.code_mem[68][6] ),
    .A1(\mem.mem_internal.code_mem[69][6] ),
    .A2(\mem.mem_internal.code_mem[70][6] ),
    .A3(\mem.mem_internal.code_mem[71][6] ),
    .S1(net953),
    .X(_06957_));
 sg13g2_mux4_1 _25646_ (.S0(net963),
    .A0(\mem.mem_internal.code_mem[80][6] ),
    .A1(\mem.mem_internal.code_mem[81][6] ),
    .A2(\mem.mem_internal.code_mem[82][6] ),
    .A3(\mem.mem_internal.code_mem[83][6] ),
    .S1(net964),
    .X(_06958_));
 sg13g2_mux4_1 _25647_ (.S0(net916),
    .A0(\mem.mem_internal.code_mem[84][6] ),
    .A1(\mem.mem_internal.code_mem[85][6] ),
    .A2(\mem.mem_internal.code_mem[86][6] ),
    .A3(\mem.mem_internal.code_mem[87][6] ),
    .S1(_06368_),
    .X(_06959_));
 sg13g2_mux4_1 _25648_ (.S0(net967),
    .A0(_06956_),
    .A1(_06957_),
    .A2(_06958_),
    .A3(_06959_),
    .S1(_06427_),
    .X(_06960_));
 sg13g2_mux4_1 _25649_ (.S0(_06363_),
    .A0(\mem.mem_internal.code_mem[72][6] ),
    .A1(\mem.mem_internal.code_mem[73][6] ),
    .A2(\mem.mem_internal.code_mem[74][6] ),
    .A3(\mem.mem_internal.code_mem[75][6] ),
    .S1(_06420_),
    .X(_06961_));
 sg13g2_mux4_1 _25650_ (.S0(_06173_),
    .A0(\mem.mem_internal.code_mem[76][6] ),
    .A1(\mem.mem_internal.code_mem[77][6] ),
    .A2(\mem.mem_internal.code_mem[78][6] ),
    .A3(\mem.mem_internal.code_mem[79][6] ),
    .S1(_06175_),
    .X(_06962_));
 sg13g2_mux4_1 _25651_ (.S0(net914),
    .A0(\mem.mem_internal.code_mem[88][6] ),
    .A1(\mem.mem_internal.code_mem[89][6] ),
    .A2(\mem.mem_internal.code_mem[90][6] ),
    .A3(\mem.mem_internal.code_mem[91][6] ),
    .S1(net910),
    .X(_06963_));
 sg13g2_mux4_1 _25652_ (.S0(net890),
    .A0(\mem.mem_internal.code_mem[92][6] ),
    .A1(\mem.mem_internal.code_mem[93][6] ),
    .A2(\mem.mem_internal.code_mem[94][6] ),
    .A3(\mem.mem_internal.code_mem[95][6] ),
    .S1(_06412_),
    .X(_06964_));
 sg13g2_mux4_1 _25653_ (.S0(_06373_),
    .A0(_06961_),
    .A1(_06962_),
    .A2(_06963_),
    .A3(_06964_),
    .S1(_06374_),
    .X(_06965_));
 sg13g2_mux4_1 _25654_ (.S0(_06250_),
    .A0(\mem.mem_internal.code_mem[192][6] ),
    .A1(\mem.mem_internal.code_mem[193][6] ),
    .A2(\mem.mem_internal.code_mem[194][6] ),
    .A3(\mem.mem_internal.code_mem[195][6] ),
    .S1(_06423_),
    .X(_06966_));
 sg13g2_mux4_1 _25655_ (.S0(_06356_),
    .A0(\mem.mem_internal.code_mem[196][6] ),
    .A1(\mem.mem_internal.code_mem[197][6] ),
    .A2(\mem.mem_internal.code_mem[198][6] ),
    .A3(\mem.mem_internal.code_mem[199][6] ),
    .S1(_06358_),
    .X(_06967_));
 sg13g2_mux4_1 _25656_ (.S0(net959),
    .A0(\mem.mem_internal.code_mem[208][6] ),
    .A1(\mem.mem_internal.code_mem[209][6] ),
    .A2(\mem.mem_internal.code_mem[210][6] ),
    .A3(\mem.mem_internal.code_mem[211][6] ),
    .S1(net961),
    .X(_06968_));
 sg13g2_mux4_1 _25657_ (.S0(_06443_),
    .A0(\mem.mem_internal.code_mem[212][6] ),
    .A1(\mem.mem_internal.code_mem[213][6] ),
    .A2(\mem.mem_internal.code_mem[214][6] ),
    .A3(\mem.mem_internal.code_mem[215][6] ),
    .S1(_06489_),
    .X(_06969_));
 sg13g2_mux4_1 _25658_ (.S0(net1231),
    .A0(_06966_),
    .A1(_06967_),
    .A2(_06968_),
    .A3(_06969_),
    .S1(_06275_),
    .X(_06970_));
 sg13g2_mux4_1 _25659_ (.S0(_06425_),
    .A0(\mem.mem_internal.code_mem[200][6] ),
    .A1(\mem.mem_internal.code_mem[201][6] ),
    .A2(\mem.mem_internal.code_mem[202][6] ),
    .A3(\mem.mem_internal.code_mem[203][6] ),
    .S1(net905),
    .X(_06971_));
 sg13g2_mux4_1 _25660_ (.S0(_06486_),
    .A0(\mem.mem_internal.code_mem[204][6] ),
    .A1(\mem.mem_internal.code_mem[205][6] ),
    .A2(\mem.mem_internal.code_mem[206][6] ),
    .A3(\mem.mem_internal.code_mem[207][6] ),
    .S1(net889),
    .X(_06972_));
 sg13g2_mux4_1 _25661_ (.S0(_06453_),
    .A0(\mem.mem_internal.code_mem[216][6] ),
    .A1(\mem.mem_internal.code_mem[217][6] ),
    .A2(\mem.mem_internal.code_mem[218][6] ),
    .A3(\mem.mem_internal.code_mem[219][6] ),
    .S1(_06441_),
    .X(_06973_));
 sg13g2_mux4_1 _25662_ (.S0(_06497_),
    .A0(\mem.mem_internal.code_mem[220][6] ),
    .A1(\mem.mem_internal.code_mem[221][6] ),
    .A2(\mem.mem_internal.code_mem[222][6] ),
    .A3(\mem.mem_internal.code_mem[223][6] ),
    .S1(_06456_),
    .X(_06974_));
 sg13g2_mux4_1 _25663_ (.S0(net1230),
    .A0(_06971_),
    .A1(_06972_),
    .A2(_06973_),
    .A3(_06974_),
    .S1(net887),
    .X(_06975_));
 sg13g2_mux4_1 _25664_ (.S0(_06168_),
    .A0(_06960_),
    .A1(_06965_),
    .A2(_06970_),
    .A3(_06975_),
    .S1(net1228),
    .X(_06976_));
 sg13g2_mux4_1 _25665_ (.S0(net956),
    .A0(\mem.mem_internal.code_mem[96][6] ),
    .A1(\mem.mem_internal.code_mem[97][6] ),
    .A2(\mem.mem_internal.code_mem[98][6] ),
    .A3(\mem.mem_internal.code_mem[99][6] ),
    .S1(_06347_),
    .X(_06977_));
 sg13g2_mux4_1 _25666_ (.S0(_06474_),
    .A0(\mem.mem_internal.code_mem[100][6] ),
    .A1(\mem.mem_internal.code_mem[101][6] ),
    .A2(\mem.mem_internal.code_mem[102][6] ),
    .A3(\mem.mem_internal.code_mem[103][6] ),
    .S1(_06466_),
    .X(_06978_));
 sg13g2_mux4_1 _25667_ (.S0(net906),
    .A0(\mem.mem_internal.code_mem[112][6] ),
    .A1(\mem.mem_internal.code_mem[113][6] ),
    .A2(\mem.mem_internal.code_mem[114][6] ),
    .A3(\mem.mem_internal.code_mem[115][6] ),
    .S1(_06468_),
    .X(_06979_));
 sg13g2_mux4_1 _25668_ (.S0(net897),
    .A0(\mem.mem_internal.code_mem[116][6] ),
    .A1(\mem.mem_internal.code_mem[117][6] ),
    .A2(\mem.mem_internal.code_mem[118][6] ),
    .A3(\mem.mem_internal.code_mem[119][6] ),
    .S1(net886),
    .X(_06980_));
 sg13g2_mux4_1 _25669_ (.S0(_06472_),
    .A0(_06977_),
    .A1(_06978_),
    .A2(_06979_),
    .A3(_06980_),
    .S1(_06361_),
    .X(_06981_));
 sg13g2_mux4_1 _25670_ (.S0(net950),
    .A0(\mem.mem_internal.code_mem[104][6] ),
    .A1(\mem.mem_internal.code_mem[105][6] ),
    .A2(\mem.mem_internal.code_mem[106][6] ),
    .A3(\mem.mem_internal.code_mem[107][6] ),
    .S1(net798),
    .X(_06982_));
 sg13g2_mux4_1 _25671_ (.S0(_06399_),
    .A0(\mem.mem_internal.code_mem[108][6] ),
    .A1(\mem.mem_internal.code_mem[109][6] ),
    .A2(\mem.mem_internal.code_mem[110][6] ),
    .A3(\mem.mem_internal.code_mem[111][6] ),
    .S1(_06393_),
    .X(_06983_));
 sg13g2_mux4_1 _25672_ (.S0(net913),
    .A0(\mem.mem_internal.code_mem[120][6] ),
    .A1(\mem.mem_internal.code_mem[121][6] ),
    .A2(\mem.mem_internal.code_mem[122][6] ),
    .A3(\mem.mem_internal.code_mem[123][6] ),
    .S1(net904),
    .X(_06984_));
 sg13g2_mux4_1 _25673_ (.S0(_06480_),
    .A0(\mem.mem_internal.code_mem[124][6] ),
    .A1(\mem.mem_internal.code_mem[125][6] ),
    .A2(\mem.mem_internal.code_mem[126][6] ),
    .A3(\mem.mem_internal.code_mem[127][6] ),
    .S1(net892),
    .X(_06985_));
 sg13g2_mux4_1 _25674_ (.S0(_06406_),
    .A0(_06982_),
    .A1(_06983_),
    .A2(_06984_),
    .A3(_06985_),
    .S1(_06407_),
    .X(_06986_));
 sg13g2_mux4_1 _25675_ (.S0(_06352_),
    .A0(\mem.mem_internal.code_mem[224][6] ),
    .A1(\mem.mem_internal.code_mem[225][6] ),
    .A2(\mem.mem_internal.code_mem[226][6] ),
    .A3(\mem.mem_internal.code_mem[227][6] ),
    .S1(_06353_),
    .X(_06987_));
 sg13g2_mux4_1 _25676_ (.S0(_06370_),
    .A0(\mem.mem_internal.code_mem[228][6] ),
    .A1(\mem.mem_internal.code_mem[229][6] ),
    .A2(\mem.mem_internal.code_mem[230][6] ),
    .A3(\mem.mem_internal.code_mem[231][6] ),
    .S1(_06487_),
    .X(_06988_));
 sg13g2_mux4_1 _25677_ (.S0(net903),
    .A0(\mem.mem_internal.code_mem[240][6] ),
    .A1(\mem.mem_internal.code_mem[241][6] ),
    .A2(\mem.mem_internal.code_mem[242][6] ),
    .A3(\mem.mem_internal.code_mem[243][6] ),
    .S1(net909),
    .X(_06989_));
 sg13g2_mux4_1 _25678_ (.S0(net902),
    .A0(\mem.mem_internal.code_mem[244][6] ),
    .A1(\mem.mem_internal.code_mem[245][6] ),
    .A2(\mem.mem_internal.code_mem[246][6] ),
    .A3(\mem.mem_internal.code_mem[247][6] ),
    .S1(net901),
    .X(_06990_));
 sg13g2_mux4_1 _25679_ (.S0(_06446_),
    .A0(_06987_),
    .A1(_06988_),
    .A2(_06989_),
    .A3(_06990_),
    .S1(_06492_),
    .X(_06991_));
 sg13g2_mux4_1 _25680_ (.S0(_06402_),
    .A0(\mem.mem_internal.code_mem[232][6] ),
    .A1(\mem.mem_internal.code_mem[233][6] ),
    .A2(\mem.mem_internal.code_mem[234][6] ),
    .A3(\mem.mem_internal.code_mem[235][6] ),
    .S1(net924),
    .X(_06992_));
 sg13g2_mux4_1 _25681_ (.S0(_06182_),
    .A0(\mem.mem_internal.code_mem[236][6] ),
    .A1(\mem.mem_internal.code_mem[237][6] ),
    .A2(\mem.mem_internal.code_mem[238][6] ),
    .A3(\mem.mem_internal.code_mem[239][6] ),
    .S1(net982),
    .X(_06993_));
 sg13g2_mux4_1 _25682_ (.S0(net885),
    .A0(\mem.mem_internal.code_mem[248][6] ),
    .A1(\mem.mem_internal.code_mem[249][6] ),
    .A2(\mem.mem_internal.code_mem[250][6] ),
    .A3(\mem.mem_internal.code_mem[251][6] ),
    .S1(net907),
    .X(_06994_));
 sg13g2_mux4_1 _25683_ (.S0(_06202_),
    .A0(\mem.mem_internal.code_mem[252][6] ),
    .A1(\mem.mem_internal.code_mem[253][6] ),
    .A2(\mem.mem_internal.code_mem[254][6] ),
    .A3(\mem.mem_internal.code_mem[255][6] ),
    .S1(_06204_),
    .X(_06995_));
 sg13g2_mux4_1 _25684_ (.S0(_06211_),
    .A0(_06992_),
    .A1(_06993_),
    .A2(_06994_),
    .A3(_06995_),
    .S1(net900),
    .X(_06996_));
 sg13g2_mux4_1 _25685_ (.S0(_06461_),
    .A0(_06981_),
    .A1(_06986_),
    .A2(_06991_),
    .A3(_06996_),
    .S1(_06462_),
    .X(_06997_));
 sg13g2_mux4_1 _25686_ (.S0(_06300_),
    .A0(_06934_),
    .A1(_06955_),
    .A2(_06976_),
    .A3(_06997_),
    .S1(_06301_),
    .X(_06998_));
 sg13g2_nor2_1 _25687_ (.A(_06304_),
    .B(_06998_),
    .Y(_06999_));
 sg13g2_a21oi_1 _25688_ (.A1(net832),
    .A2(_06913_),
    .Y(_07000_),
    .B1(_06999_));
 sg13g2_nand2_1 _25689_ (.Y(_07001_),
    .A(\mem.internal_data_out[6] ),
    .B(_06126_));
 sg13g2_o21ai_1 _25690_ (.B1(_07001_),
    .Y(_02426_),
    .A1(_06127_),
    .A2(_07000_));
 sg13g2_mux4_1 _25691_ (.S0(net538),
    .A0(\mem.mem_internal.data_mem[0][7] ),
    .A1(\mem.mem_internal.data_mem[1][7] ),
    .A2(\mem.mem_internal.data_mem[2][7] ),
    .A3(\mem.mem_internal.data_mem[3][7] ),
    .S1(net537),
    .X(_07002_));
 sg13g2_mux4_1 _25692_ (.S0(net545),
    .A0(\mem.mem_internal.data_mem[4][7] ),
    .A1(\mem.mem_internal.data_mem[5][7] ),
    .A2(\mem.mem_internal.data_mem[6][7] ),
    .A3(\mem.mem_internal.data_mem[7][7] ),
    .S1(net544),
    .X(_07003_));
 sg13g2_mux4_1 _25693_ (.S0(_06142_),
    .A0(\mem.mem_internal.data_mem[16][7] ),
    .A1(\mem.mem_internal.data_mem[17][7] ),
    .A2(\mem.mem_internal.data_mem[18][7] ),
    .A3(\mem.mem_internal.data_mem[19][7] ),
    .S1(_06143_),
    .X(_07004_));
 sg13g2_mux4_1 _25694_ (.S0(net542),
    .A0(\mem.mem_internal.data_mem[20][7] ),
    .A1(\mem.mem_internal.data_mem[21][7] ),
    .A2(\mem.mem_internal.data_mem[22][7] ),
    .A3(\mem.mem_internal.data_mem[23][7] ),
    .S1(net541),
    .X(_07005_));
 sg13g2_mux4_1 _25695_ (.S0(net818),
    .A0(_07002_),
    .A1(_07003_),
    .A2(_07004_),
    .A3(_07005_),
    .S1(_06155_),
    .X(_07006_));
 sg13g2_mux4_1 _25696_ (.S0(_06145_),
    .A0(\mem.mem_internal.data_mem[8][7] ),
    .A1(\mem.mem_internal.data_mem[9][7] ),
    .A2(\mem.mem_internal.data_mem[10][7] ),
    .A3(\mem.mem_internal.data_mem[11][7] ),
    .S1(_06146_),
    .X(_07007_));
 sg13g2_mux4_1 _25697_ (.S0(net540),
    .A0(\mem.mem_internal.data_mem[12][7] ),
    .A1(\mem.mem_internal.data_mem[13][7] ),
    .A2(\mem.mem_internal.data_mem[14][7] ),
    .A3(\mem.mem_internal.data_mem[15][7] ),
    .S1(net539),
    .X(_07008_));
 sg13g2_mux4_1 _25698_ (.S0(_06132_),
    .A0(\mem.mem_internal.data_mem[24][7] ),
    .A1(\mem.mem_internal.data_mem[25][7] ),
    .A2(\mem.mem_internal.data_mem[26][7] ),
    .A3(\mem.mem_internal.data_mem[27][7] ),
    .S1(net578),
    .X(_07009_));
 sg13g2_mux4_1 _25699_ (.S0(_06163_),
    .A0(\mem.mem_internal.data_mem[28][7] ),
    .A1(\mem.mem_internal.data_mem[29][7] ),
    .A2(\mem.mem_internal.data_mem[30][7] ),
    .A3(\mem.mem_internal.data_mem[31][7] ),
    .S1(_06164_),
    .X(_07010_));
 sg13g2_mux4_1 _25700_ (.S0(net988),
    .A0(_07007_),
    .A1(_07008_),
    .A2(_07009_),
    .A3(_07010_),
    .S1(net987),
    .X(_07011_));
 sg13g2_mux2_1 _25701_ (.A0(_07006_),
    .A1(_07011_),
    .S(net986),
    .X(_07012_));
 sg13g2_mux4_1 _25702_ (.S0(_06319_),
    .A0(\mem.mem_internal.code_mem[0][7] ),
    .A1(\mem.mem_internal.code_mem[1][7] ),
    .A2(\mem.mem_internal.code_mem[2][7] ),
    .A3(\mem.mem_internal.code_mem[3][7] ),
    .S1(_06232_),
    .X(_07013_));
 sg13g2_mux4_1 _25703_ (.S0(net931),
    .A0(\mem.mem_internal.code_mem[4][7] ),
    .A1(\mem.mem_internal.code_mem[5][7] ),
    .A2(\mem.mem_internal.code_mem[6][7] ),
    .A3(\mem.mem_internal.code_mem[7][7] ),
    .S1(net814),
    .X(_07014_));
 sg13g2_mux4_1 _25704_ (.S0(net920),
    .A0(\mem.mem_internal.code_mem[16][7] ),
    .A1(\mem.mem_internal.code_mem[17][7] ),
    .A2(\mem.mem_internal.code_mem[18][7] ),
    .A3(\mem.mem_internal.code_mem[19][7] ),
    .S1(net955),
    .X(_07015_));
 sg13g2_mux4_1 _25705_ (.S0(_06327_),
    .A0(\mem.mem_internal.code_mem[20][7] ),
    .A1(\mem.mem_internal.code_mem[21][7] ),
    .A2(\mem.mem_internal.code_mem[22][7] ),
    .A3(\mem.mem_internal.code_mem[23][7] ),
    .S1(_06328_),
    .X(_07016_));
 sg13g2_mux4_1 _25706_ (.S0(_06190_),
    .A0(_07013_),
    .A1(_07014_),
    .A2(_07015_),
    .A3(_07016_),
    .S1(_06191_),
    .X(_07017_));
 sg13g2_mux4_1 _25707_ (.S0(_06378_),
    .A0(\mem.mem_internal.code_mem[8][7] ),
    .A1(\mem.mem_internal.code_mem[9][7] ),
    .A2(\mem.mem_internal.code_mem[10][7] ),
    .A3(\mem.mem_internal.code_mem[11][7] ),
    .S1(_06333_),
    .X(_07018_));
 sg13g2_mux4_1 _25708_ (.S0(_06335_),
    .A0(\mem.mem_internal.code_mem[12][7] ),
    .A1(\mem.mem_internal.code_mem[13][7] ),
    .A2(\mem.mem_internal.code_mem[14][7] ),
    .A3(\mem.mem_internal.code_mem[15][7] ),
    .S1(_06380_),
    .X(_07019_));
 sg13g2_mux4_1 _25709_ (.S0(net950),
    .A0(\mem.mem_internal.code_mem[24][7] ),
    .A1(\mem.mem_internal.code_mem[25][7] ),
    .A2(\mem.mem_internal.code_mem[26][7] ),
    .A3(\mem.mem_internal.code_mem[27][7] ),
    .S1(_06340_),
    .X(_07020_));
 sg13g2_mux4_1 _25710_ (.S0(_06385_),
    .A0(\mem.mem_internal.code_mem[28][7] ),
    .A1(\mem.mem_internal.code_mem[29][7] ),
    .A2(\mem.mem_internal.code_mem[30][7] ),
    .A3(\mem.mem_internal.code_mem[31][7] ),
    .S1(_06386_),
    .X(_07021_));
 sg13g2_mux4_1 _25711_ (.S0(_06330_),
    .A0(_07018_),
    .A1(_07019_),
    .A2(_07020_),
    .A3(_07021_),
    .S1(net951),
    .X(_07022_));
 sg13g2_mux4_1 _25712_ (.S0(_06417_),
    .A0(\mem.mem_internal.code_mem[128][7] ),
    .A1(\mem.mem_internal.code_mem[129][7] ),
    .A2(\mem.mem_internal.code_mem[130][7] ),
    .A3(\mem.mem_internal.code_mem[131][7] ),
    .S1(net946),
    .X(_07023_));
 sg13g2_mux4_1 _25713_ (.S0(_06382_),
    .A0(\mem.mem_internal.code_mem[132][7] ),
    .A1(\mem.mem_internal.code_mem[133][7] ),
    .A2(\mem.mem_internal.code_mem[134][7] ),
    .A3(\mem.mem_internal.code_mem[135][7] ),
    .S1(net808),
    .X(_07024_));
 sg13g2_mux4_1 _25714_ (.S0(net918),
    .A0(\mem.mem_internal.code_mem[144][7] ),
    .A1(\mem.mem_internal.code_mem[145][7] ),
    .A2(\mem.mem_internal.code_mem[146][7] ),
    .A3(\mem.mem_internal.code_mem[147][7] ),
    .S1(net917),
    .X(_07025_));
 sg13g2_mux4_1 _25715_ (.S0(net937),
    .A0(\mem.mem_internal.code_mem[148][7] ),
    .A1(\mem.mem_internal.code_mem[149][7] ),
    .A2(\mem.mem_internal.code_mem[150][7] ),
    .A3(\mem.mem_internal.code_mem[151][7] ),
    .S1(net941),
    .X(_07026_));
 sg13g2_mux4_1 _25716_ (.S0(net940),
    .A0(_07023_),
    .A1(_07024_),
    .A2(_07025_),
    .A3(_07026_),
    .S1(net915),
    .X(_07027_));
 sg13g2_mux4_1 _25717_ (.S0(_06327_),
    .A0(\mem.mem_internal.code_mem[136][7] ),
    .A1(\mem.mem_internal.code_mem[137][7] ),
    .A2(\mem.mem_internal.code_mem[138][7] ),
    .A3(\mem.mem_internal.code_mem[139][7] ),
    .S1(net899),
    .X(_07028_));
 sg13g2_mux4_1 _25718_ (.S0(net884),
    .A0(\mem.mem_internal.code_mem[140][7] ),
    .A1(\mem.mem_internal.code_mem[141][7] ),
    .A2(\mem.mem_internal.code_mem[142][7] ),
    .A3(\mem.mem_internal.code_mem[143][7] ),
    .S1(net797),
    .X(_07029_));
 sg13g2_mux4_1 _25719_ (.S0(net937),
    .A0(\mem.mem_internal.code_mem[152][7] ),
    .A1(\mem.mem_internal.code_mem[153][7] ),
    .A2(\mem.mem_internal.code_mem[154][7] ),
    .A3(\mem.mem_internal.code_mem[155][7] ),
    .S1(net898),
    .X(_07030_));
 sg13g2_mux4_1 _25720_ (.S0(net935),
    .A0(\mem.mem_internal.code_mem[156][7] ),
    .A1(\mem.mem_internal.code_mem[157][7] ),
    .A2(\mem.mem_internal.code_mem[158][7] ),
    .A3(\mem.mem_internal.code_mem[159][7] ),
    .S1(net934),
    .X(_07031_));
 sg13g2_mux4_1 _25721_ (.S0(net896),
    .A0(_07028_),
    .A1(_07029_),
    .A2(_07030_),
    .A3(_07031_),
    .S1(net932),
    .X(_07032_));
 sg13g2_mux4_1 _25722_ (.S0(net1234),
    .A0(_07017_),
    .A1(_07022_),
    .A2(_07027_),
    .A3(_07032_),
    .S1(net1233),
    .X(_07033_));
 sg13g2_mux4_1 _25723_ (.S0(net958),
    .A0(\mem.mem_internal.code_mem[32][7] ),
    .A1(\mem.mem_internal.code_mem[33][7] ),
    .A2(\mem.mem_internal.code_mem[34][7] ),
    .A3(\mem.mem_internal.code_mem[35][7] ),
    .S1(net813),
    .X(_07034_));
 sg13g2_mux4_1 _25724_ (.S0(net803),
    .A0(\mem.mem_internal.code_mem[36][7] ),
    .A1(\mem.mem_internal.code_mem[37][7] ),
    .A2(\mem.mem_internal.code_mem[38][7] ),
    .A3(\mem.mem_internal.code_mem[39][7] ),
    .S1(net806),
    .X(_07035_));
 sg13g2_mux4_1 _25725_ (.S0(net930),
    .A0(\mem.mem_internal.code_mem[48][7] ),
    .A1(\mem.mem_internal.code_mem[49][7] ),
    .A2(\mem.mem_internal.code_mem[50][7] ),
    .A3(\mem.mem_internal.code_mem[51][7] ),
    .S1(_06350_),
    .X(_07036_));
 sg13g2_mux4_1 _25726_ (.S0(net929),
    .A0(\mem.mem_internal.code_mem[52][7] ),
    .A1(\mem.mem_internal.code_mem[53][7] ),
    .A2(\mem.mem_internal.code_mem[54][7] ),
    .A3(\mem.mem_internal.code_mem[55][7] ),
    .S1(_06365_),
    .X(_07037_));
 sg13g2_mux4_1 _25727_ (.S0(net952),
    .A0(_07034_),
    .A1(_07035_),
    .A2(_07036_),
    .A3(_07037_),
    .S1(net947),
    .X(_07038_));
 sg13g2_mux4_1 _25728_ (.S0(net957),
    .A0(\mem.mem_internal.code_mem[40][7] ),
    .A1(\mem.mem_internal.code_mem[41][7] ),
    .A2(\mem.mem_internal.code_mem[42][7] ),
    .A3(\mem.mem_internal.code_mem[43][7] ),
    .S1(net810),
    .X(_07039_));
 sg13g2_mux4_1 _25729_ (.S0(net811),
    .A0(\mem.mem_internal.code_mem[44][7] ),
    .A1(\mem.mem_internal.code_mem[45][7] ),
    .A2(\mem.mem_internal.code_mem[46][7] ),
    .A3(\mem.mem_internal.code_mem[47][7] ),
    .S1(_06137_),
    .X(_07040_));
 sg13g2_mux4_1 _25730_ (.S0(net985),
    .A0(\mem.mem_internal.code_mem[56][7] ),
    .A1(\mem.mem_internal.code_mem[57][7] ),
    .A2(\mem.mem_internal.code_mem[58][7] ),
    .A3(\mem.mem_internal.code_mem[59][7] ),
    .S1(_06400_),
    .X(_07041_));
 sg13g2_mux4_1 _25731_ (.S0(net926),
    .A0(\mem.mem_internal.code_mem[60][7] ),
    .A1(\mem.mem_internal.code_mem[61][7] ),
    .A2(\mem.mem_internal.code_mem[62][7] ),
    .A3(\mem.mem_internal.code_mem[63][7] ),
    .S1(_06410_),
    .X(_07042_));
 sg13g2_mux4_1 _25732_ (.S0(net948),
    .A0(_07039_),
    .A1(_07040_),
    .A2(_07041_),
    .A3(_07042_),
    .S1(_06154_),
    .X(_07043_));
 sg13g2_mux4_1 _25733_ (.S0(net945),
    .A0(\mem.mem_internal.code_mem[160][7] ),
    .A1(\mem.mem_internal.code_mem[161][7] ),
    .A2(\mem.mem_internal.code_mem[162][7] ),
    .A3(\mem.mem_internal.code_mem[163][7] ),
    .S1(_06383_),
    .X(_07044_));
 sg13g2_mux4_1 _25734_ (.S0(net928),
    .A0(\mem.mem_internal.code_mem[164][7] ),
    .A1(\mem.mem_internal.code_mem[165][7] ),
    .A2(\mem.mem_internal.code_mem[166][7] ),
    .A3(\mem.mem_internal.code_mem[167][7] ),
    .S1(net801),
    .X(_07045_));
 sg13g2_mux4_1 _25735_ (.S0(_06431_),
    .A0(\mem.mem_internal.code_mem[176][7] ),
    .A1(\mem.mem_internal.code_mem[177][7] ),
    .A2(\mem.mem_internal.code_mem[178][7] ),
    .A3(\mem.mem_internal.code_mem[179][7] ),
    .S1(net924),
    .X(_07046_));
 sg13g2_mux4_1 _25736_ (.S0(net962),
    .A0(\mem.mem_internal.code_mem[180][7] ),
    .A1(\mem.mem_internal.code_mem[181][7] ),
    .A2(\mem.mem_internal.code_mem[182][7] ),
    .A3(\mem.mem_internal.code_mem[183][7] ),
    .S1(net912),
    .X(_07047_));
 sg13g2_mux4_1 _25737_ (.S0(net923),
    .A0(_07044_),
    .A1(_07045_),
    .A2(_07046_),
    .A3(_07047_),
    .S1(net911),
    .X(_07048_));
 sg13g2_mux4_1 _25738_ (.S0(net949),
    .A0(\mem.mem_internal.code_mem[168][7] ),
    .A1(\mem.mem_internal.code_mem[169][7] ),
    .A2(\mem.mem_internal.code_mem[170][7] ),
    .A3(\mem.mem_internal.code_mem[171][7] ),
    .S1(net807),
    .X(_07049_));
 sg13g2_mux4_1 _25739_ (.S0(net927),
    .A0(\mem.mem_internal.code_mem[172][7] ),
    .A1(\mem.mem_internal.code_mem[173][7] ),
    .A2(\mem.mem_internal.code_mem[174][7] ),
    .A3(\mem.mem_internal.code_mem[175][7] ),
    .S1(net800),
    .X(_07050_));
 sg13g2_mux4_1 _25740_ (.S0(net894),
    .A0(\mem.mem_internal.code_mem[184][7] ),
    .A1(\mem.mem_internal.code_mem[185][7] ),
    .A2(\mem.mem_internal.code_mem[186][7] ),
    .A3(\mem.mem_internal.code_mem[187][7] ),
    .S1(net921),
    .X(_07051_));
 sg13g2_mux4_1 _25741_ (.S0(net893),
    .A0(\mem.mem_internal.code_mem[188][7] ),
    .A1(\mem.mem_internal.code_mem[189][7] ),
    .A2(\mem.mem_internal.code_mem[190][7] ),
    .A3(\mem.mem_internal.code_mem[191][7] ),
    .S1(net892),
    .X(_07052_));
 sg13g2_mux4_1 _25742_ (.S0(net891),
    .A0(_07049_),
    .A1(_07050_),
    .A2(_07051_),
    .A3(_07052_),
    .S1(net922),
    .X(_07053_));
 sg13g2_mux4_1 _25743_ (.S0(_06169_),
    .A0(_07038_),
    .A1(_07043_),
    .A2(_07048_),
    .A3(_07053_),
    .S1(net1232),
    .X(_07054_));
 sg13g2_mux4_1 _25744_ (.S0(_06238_),
    .A0(\mem.mem_internal.code_mem[64][7] ),
    .A1(\mem.mem_internal.code_mem[65][7] ),
    .A2(\mem.mem_internal.code_mem[66][7] ),
    .A3(\mem.mem_internal.code_mem[67][7] ),
    .S1(net966),
    .X(_07055_));
 sg13g2_mux4_1 _25745_ (.S0(net919),
    .A0(\mem.mem_internal.code_mem[68][7] ),
    .A1(\mem.mem_internal.code_mem[69][7] ),
    .A2(\mem.mem_internal.code_mem[70][7] ),
    .A3(\mem.mem_internal.code_mem[71][7] ),
    .S1(net953),
    .X(_07056_));
 sg13g2_mux4_1 _25746_ (.S0(net963),
    .A0(\mem.mem_internal.code_mem[80][7] ),
    .A1(\mem.mem_internal.code_mem[81][7] ),
    .A2(\mem.mem_internal.code_mem[82][7] ),
    .A3(\mem.mem_internal.code_mem[83][7] ),
    .S1(net964),
    .X(_07057_));
 sg13g2_mux4_1 _25747_ (.S0(net916),
    .A0(\mem.mem_internal.code_mem[84][7] ),
    .A1(\mem.mem_internal.code_mem[85][7] ),
    .A2(\mem.mem_internal.code_mem[86][7] ),
    .A3(\mem.mem_internal.code_mem[87][7] ),
    .S1(_06368_),
    .X(_07058_));
 sg13g2_mux4_1 _25748_ (.S0(_06221_),
    .A0(_07055_),
    .A1(_07056_),
    .A2(_07057_),
    .A3(_07058_),
    .S1(net970),
    .X(_07059_));
 sg13g2_mux4_1 _25749_ (.S0(_06363_),
    .A0(\mem.mem_internal.code_mem[72][7] ),
    .A1(\mem.mem_internal.code_mem[73][7] ),
    .A2(\mem.mem_internal.code_mem[74][7] ),
    .A3(\mem.mem_internal.code_mem[75][7] ),
    .S1(net799),
    .X(_07060_));
 sg13g2_mux4_1 _25750_ (.S0(_06173_),
    .A0(\mem.mem_internal.code_mem[76][7] ),
    .A1(\mem.mem_internal.code_mem[77][7] ),
    .A2(\mem.mem_internal.code_mem[78][7] ),
    .A3(\mem.mem_internal.code_mem[79][7] ),
    .S1(_06175_),
    .X(_07061_));
 sg13g2_mux4_1 _25751_ (.S0(net914),
    .A0(\mem.mem_internal.code_mem[88][7] ),
    .A1(\mem.mem_internal.code_mem[89][7] ),
    .A2(\mem.mem_internal.code_mem[90][7] ),
    .A3(\mem.mem_internal.code_mem[91][7] ),
    .S1(net910),
    .X(_07062_));
 sg13g2_mux4_1 _25752_ (.S0(net890),
    .A0(\mem.mem_internal.code_mem[92][7] ),
    .A1(\mem.mem_internal.code_mem[93][7] ),
    .A2(\mem.mem_internal.code_mem[94][7] ),
    .A3(\mem.mem_internal.code_mem[95][7] ),
    .S1(_06412_),
    .X(_07063_));
 sg13g2_mux4_1 _25753_ (.S0(_06373_),
    .A0(_07060_),
    .A1(_07061_),
    .A2(_07062_),
    .A3(_07063_),
    .S1(_06374_),
    .X(_07064_));
 sg13g2_mux4_1 _25754_ (.S0(_06250_),
    .A0(\mem.mem_internal.code_mem[192][7] ),
    .A1(\mem.mem_internal.code_mem[193][7] ),
    .A2(\mem.mem_internal.code_mem[194][7] ),
    .A3(\mem.mem_internal.code_mem[195][7] ),
    .S1(_06423_),
    .X(_07065_));
 sg13g2_mux4_1 _25755_ (.S0(_06356_),
    .A0(\mem.mem_internal.code_mem[196][7] ),
    .A1(\mem.mem_internal.code_mem[197][7] ),
    .A2(\mem.mem_internal.code_mem[198][7] ),
    .A3(\mem.mem_internal.code_mem[199][7] ),
    .S1(_06358_),
    .X(_07066_));
 sg13g2_mux4_1 _25756_ (.S0(_06291_),
    .A0(\mem.mem_internal.code_mem[208][7] ),
    .A1(\mem.mem_internal.code_mem[209][7] ),
    .A2(\mem.mem_internal.code_mem[210][7] ),
    .A3(\mem.mem_internal.code_mem[211][7] ),
    .S1(_06273_),
    .X(_07067_));
 sg13g2_mux4_1 _25757_ (.S0(_06443_),
    .A0(\mem.mem_internal.code_mem[212][7] ),
    .A1(\mem.mem_internal.code_mem[213][7] ),
    .A2(\mem.mem_internal.code_mem[214][7] ),
    .A3(\mem.mem_internal.code_mem[215][7] ),
    .S1(_06489_),
    .X(_07068_));
 sg13g2_mux4_1 _25758_ (.S0(_06149_),
    .A0(_07065_),
    .A1(_07066_),
    .A2(_07067_),
    .A3(_07068_),
    .S1(_06275_),
    .X(_07069_));
 sg13g2_mux4_1 _25759_ (.S0(_06425_),
    .A0(\mem.mem_internal.code_mem[200][7] ),
    .A1(\mem.mem_internal.code_mem[201][7] ),
    .A2(\mem.mem_internal.code_mem[202][7] ),
    .A3(\mem.mem_internal.code_mem[203][7] ),
    .S1(net905),
    .X(_07070_));
 sg13g2_mux4_1 _25760_ (.S0(_06486_),
    .A0(\mem.mem_internal.code_mem[204][7] ),
    .A1(\mem.mem_internal.code_mem[205][7] ),
    .A2(\mem.mem_internal.code_mem[206][7] ),
    .A3(\mem.mem_internal.code_mem[207][7] ),
    .S1(net889),
    .X(_07071_));
 sg13g2_mux4_1 _25761_ (.S0(_06291_),
    .A0(\mem.mem_internal.code_mem[216][7] ),
    .A1(\mem.mem_internal.code_mem[217][7] ),
    .A2(\mem.mem_internal.code_mem[218][7] ),
    .A3(\mem.mem_internal.code_mem[219][7] ),
    .S1(_06441_),
    .X(_07072_));
 sg13g2_mux4_1 _25762_ (.S0(_06497_),
    .A0(\mem.mem_internal.code_mem[220][7] ),
    .A1(\mem.mem_internal.code_mem[221][7] ),
    .A2(\mem.mem_internal.code_mem[222][7] ),
    .A3(\mem.mem_internal.code_mem[223][7] ),
    .S1(_06444_),
    .X(_07073_));
 sg13g2_mux4_1 _25763_ (.S0(net1230),
    .A0(_07070_),
    .A1(_07071_),
    .A2(_07072_),
    .A3(_07073_),
    .S1(net887),
    .X(_07074_));
 sg13g2_mux4_1 _25764_ (.S0(_06168_),
    .A0(_07059_),
    .A1(_07064_),
    .A2(_07069_),
    .A3(_07074_),
    .S1(net1228),
    .X(_07075_));
 sg13g2_mux4_1 _25765_ (.S0(net956),
    .A0(\mem.mem_internal.code_mem[96][7] ),
    .A1(\mem.mem_internal.code_mem[97][7] ),
    .A2(\mem.mem_internal.code_mem[98][7] ),
    .A3(\mem.mem_internal.code_mem[99][7] ),
    .S1(_06347_),
    .X(_07076_));
 sg13g2_mux4_1 _25766_ (.S0(_06474_),
    .A0(\mem.mem_internal.code_mem[100][7] ),
    .A1(\mem.mem_internal.code_mem[101][7] ),
    .A2(\mem.mem_internal.code_mem[102][7] ),
    .A3(\mem.mem_internal.code_mem[103][7] ),
    .S1(_06466_),
    .X(_07077_));
 sg13g2_mux4_1 _25767_ (.S0(net906),
    .A0(\mem.mem_internal.code_mem[112][7] ),
    .A1(\mem.mem_internal.code_mem[113][7] ),
    .A2(\mem.mem_internal.code_mem[114][7] ),
    .A3(\mem.mem_internal.code_mem[115][7] ),
    .S1(net905),
    .X(_07078_));
 sg13g2_mux4_1 _25768_ (.S0(net897),
    .A0(\mem.mem_internal.code_mem[116][7] ),
    .A1(\mem.mem_internal.code_mem[117][7] ),
    .A2(\mem.mem_internal.code_mem[118][7] ),
    .A3(\mem.mem_internal.code_mem[119][7] ),
    .S1(net886),
    .X(_07079_));
 sg13g2_mux4_1 _25769_ (.S0(_06360_),
    .A0(_07076_),
    .A1(_07077_),
    .A2(_07078_),
    .A3(_07079_),
    .S1(_06361_),
    .X(_07080_));
 sg13g2_mux4_1 _25770_ (.S0(_06338_),
    .A0(\mem.mem_internal.code_mem[104][7] ),
    .A1(\mem.mem_internal.code_mem[105][7] ),
    .A2(\mem.mem_internal.code_mem[106][7] ),
    .A3(\mem.mem_internal.code_mem[107][7] ),
    .S1(net798),
    .X(_07081_));
 sg13g2_mux4_1 _25771_ (.S0(_06399_),
    .A0(\mem.mem_internal.code_mem[108][7] ),
    .A1(\mem.mem_internal.code_mem[109][7] ),
    .A2(\mem.mem_internal.code_mem[110][7] ),
    .A3(\mem.mem_internal.code_mem[111][7] ),
    .S1(_06393_),
    .X(_07082_));
 sg13g2_mux4_1 _25772_ (.S0(net913),
    .A0(\mem.mem_internal.code_mem[120][7] ),
    .A1(\mem.mem_internal.code_mem[121][7] ),
    .A2(\mem.mem_internal.code_mem[122][7] ),
    .A3(\mem.mem_internal.code_mem[123][7] ),
    .S1(net904),
    .X(_07083_));
 sg13g2_mux4_1 _25773_ (.S0(net983),
    .A0(\mem.mem_internal.code_mem[124][7] ),
    .A1(\mem.mem_internal.code_mem[125][7] ),
    .A2(\mem.mem_internal.code_mem[126][7] ),
    .A3(\mem.mem_internal.code_mem[127][7] ),
    .S1(_06481_),
    .X(_07084_));
 sg13g2_mux4_1 _25774_ (.S0(_06406_),
    .A0(_07081_),
    .A1(_07082_),
    .A2(_07083_),
    .A3(_07084_),
    .S1(_06407_),
    .X(_07085_));
 sg13g2_mux4_1 _25775_ (.S0(_06352_),
    .A0(\mem.mem_internal.code_mem[224][7] ),
    .A1(\mem.mem_internal.code_mem[225][7] ),
    .A2(\mem.mem_internal.code_mem[226][7] ),
    .A3(\mem.mem_internal.code_mem[227][7] ),
    .S1(_06353_),
    .X(_07086_));
 sg13g2_mux4_1 _25776_ (.S0(_06370_),
    .A0(\mem.mem_internal.code_mem[228][7] ),
    .A1(\mem.mem_internal.code_mem[229][7] ),
    .A2(\mem.mem_internal.code_mem[230][7] ),
    .A3(\mem.mem_internal.code_mem[231][7] ),
    .S1(_06371_),
    .X(_07087_));
 sg13g2_mux4_1 _25777_ (.S0(net903),
    .A0(\mem.mem_internal.code_mem[240][7] ),
    .A1(\mem.mem_internal.code_mem[241][7] ),
    .A2(\mem.mem_internal.code_mem[242][7] ),
    .A3(\mem.mem_internal.code_mem[243][7] ),
    .S1(net909),
    .X(_07088_));
 sg13g2_mux4_1 _25778_ (.S0(net902),
    .A0(\mem.mem_internal.code_mem[244][7] ),
    .A1(\mem.mem_internal.code_mem[245][7] ),
    .A2(\mem.mem_internal.code_mem[246][7] ),
    .A3(\mem.mem_internal.code_mem[247][7] ),
    .S1(net901),
    .X(_07089_));
 sg13g2_mux4_1 _25779_ (.S0(_06446_),
    .A0(_07086_),
    .A1(_07087_),
    .A2(_07088_),
    .A3(_07089_),
    .S1(_06492_),
    .X(_07090_));
 sg13g2_mux4_1 _25780_ (.S0(_06402_),
    .A0(\mem.mem_internal.code_mem[232][7] ),
    .A1(\mem.mem_internal.code_mem[233][7] ),
    .A2(\mem.mem_internal.code_mem[234][7] ),
    .A3(\mem.mem_internal.code_mem[235][7] ),
    .S1(_06403_),
    .X(_07091_));
 sg13g2_mux4_1 _25781_ (.S0(_06182_),
    .A0(\mem.mem_internal.code_mem[236][7] ),
    .A1(\mem.mem_internal.code_mem[237][7] ),
    .A2(\mem.mem_internal.code_mem[238][7] ),
    .A3(\mem.mem_internal.code_mem[239][7] ),
    .S1(_06184_),
    .X(_07092_));
 sg13g2_mux4_1 _25782_ (.S0(net885),
    .A0(\mem.mem_internal.code_mem[248][7] ),
    .A1(\mem.mem_internal.code_mem[249][7] ),
    .A2(\mem.mem_internal.code_mem[250][7] ),
    .A3(\mem.mem_internal.code_mem[251][7] ),
    .S1(net907),
    .X(_07093_));
 sg13g2_mux4_1 _25783_ (.S0(_06202_),
    .A0(\mem.mem_internal.code_mem[252][7] ),
    .A1(\mem.mem_internal.code_mem[253][7] ),
    .A2(\mem.mem_internal.code_mem[254][7] ),
    .A3(\mem.mem_internal.code_mem[255][7] ),
    .S1(_06204_),
    .X(_07094_));
 sg13g2_mux4_1 _25784_ (.S0(_06211_),
    .A0(_07091_),
    .A1(_07092_),
    .A2(_07093_),
    .A3(_07094_),
    .S1(net900),
    .X(_07095_));
 sg13g2_mux4_1 _25785_ (.S0(_06461_),
    .A0(_07080_),
    .A1(_07085_),
    .A2(_07090_),
    .A3(_07095_),
    .S1(_06462_),
    .X(_07096_));
 sg13g2_mux4_1 _25786_ (.S0(_06300_),
    .A0(_07033_),
    .A1(_07054_),
    .A2(_07075_),
    .A3(_07096_),
    .S1(_06301_),
    .X(_07097_));
 sg13g2_nor2_1 _25787_ (.A(_06304_),
    .B(_07097_),
    .Y(_07098_));
 sg13g2_a21oi_1 _25788_ (.A1(net832),
    .A2(_07012_),
    .Y(_07099_),
    .B1(_07098_));
 sg13g2_nand2_1 _25789_ (.Y(_07100_),
    .A(\mem.internal_data_out[7] ),
    .B(_06126_));
 sg13g2_o21ai_1 _25790_ (.B1(_07100_),
    .Y(_02427_),
    .A1(net546),
    .A2(_07099_));
 sg13g2_buf_1 _25791_ (.A(_09881_),
    .X(_07101_));
 sg13g2_or3_1 _25792_ (.A(net1275),
    .B(net1227),
    .C(_10088_),
    .X(_07102_));
 sg13g2_nand3_1 _25793_ (.B(net1227),
    .C(net1272),
    .A(net1275),
    .Y(_07103_));
 sg13g2_o21ai_1 _25794_ (.B1(_07103_),
    .Y(_07104_),
    .A1(_00072_),
    .A2(_07102_));
 sg13g2_nand4_1 _25795_ (.B(_09890_),
    .C(_09919_),
    .A(net1278),
    .Y(_07105_),
    .D(_07104_));
 sg13g2_nand2_1 _25796_ (.Y(_07106_),
    .A(\mem.mem_internal.memory_type_data ),
    .B(_10084_));
 sg13g2_o21ai_1 _25797_ (.B1(_07106_),
    .Y(_02472_),
    .A1(net780),
    .A2(_07105_));
 sg13g2_mux2_1 _25798_ (.A0(\stack[22][0] ),
    .A1(\stack[23][0] ),
    .S(_09617_),
    .X(_07107_));
 sg13g2_and2_1 _25799_ (.A(net1280),
    .B(net1279),
    .X(_07108_));
 sg13g2_buf_2 _25800_ (.A(_07108_),
    .X(_07109_));
 sg13g2_nand2_1 _25801_ (.Y(_07110_),
    .A(net874),
    .B(\stack[21][0] ));
 sg13g2_nand2b_1 _25802_ (.Y(_07111_),
    .B(\stack[20][0] ),
    .A_N(net867));
 sg13g2_nand3_1 _25803_ (.B(_07110_),
    .C(_07111_),
    .A(_07109_),
    .Y(_07112_));
 sg13g2_o21ai_1 _25804_ (.B1(_07112_),
    .Y(_07113_),
    .A1(net863),
    .A2(_07107_));
 sg13g2_buf_1 _25805_ (.A(_09686_),
    .X(_07114_));
 sg13g2_nor2b_1 _25806_ (.A(net1281),
    .B_N(net1279),
    .Y(_07115_));
 sg13g2_buf_2 _25807_ (.A(_07115_),
    .X(_07116_));
 sg13g2_nand2_1 _25808_ (.Y(_07117_),
    .A(_09734_),
    .B(\stack[19][0] ));
 sg13g2_nand2b_1 _25809_ (.Y(_07118_),
    .B(\stack[16][0] ),
    .A_N(_09713_));
 sg13g2_a22oi_1 _25810_ (.Y(_07119_),
    .B1(_07118_),
    .B2(_09694_),
    .A2(_07117_),
    .A1(_07116_));
 sg13g2_a221oi_1 _25811_ (.B2(\stack[17][0] ),
    .C1(_07119_),
    .B1(net574),
    .A1(\stack[18][0] ),
    .Y(_07120_),
    .A2(net865));
 sg13g2_nor2_1 _25812_ (.A(net1311),
    .B(net1310),
    .Y(_07121_));
 sg13g2_buf_2 _25813_ (.A(_07121_),
    .X(_07122_));
 sg13g2_xnor2_1 _25814_ (.Y(_07123_),
    .A(_09632_),
    .B(_07122_));
 sg13g2_buf_2 _25815_ (.A(_07123_),
    .X(_07124_));
 sg13g2_nor3_1 _25816_ (.A(_09622_),
    .B(_09677_),
    .C(_09654_),
    .Y(_07125_));
 sg13g2_xnor2_1 _25817_ (.Y(_07126_),
    .A(_09653_),
    .B(_07125_));
 sg13g2_buf_2 _25818_ (.A(_07126_),
    .X(_07127_));
 sg13g2_nor2_1 _25819_ (.A(_07124_),
    .B(_07127_),
    .Y(_07128_));
 sg13g2_o21ai_1 _25820_ (.B1(_07128_),
    .Y(_07129_),
    .A1(_07113_),
    .A2(_07120_));
 sg13g2_buf_1 _25821_ (.A(_09689_),
    .X(_07130_));
 sg13g2_nand2b_1 _25822_ (.Y(_07131_),
    .B(\stack[26][0] ),
    .A_N(net1195));
 sg13g2_nand2_1 _25823_ (.Y(_07132_),
    .A(net864),
    .B(\stack[25][0] ));
 sg13g2_a22oi_1 _25824_ (.Y(_07133_),
    .B1(_07132_),
    .B2(_09694_),
    .A2(_07131_),
    .A1(_07116_));
 sg13g2_a221oi_1 _25825_ (.B2(\stack[24][0] ),
    .C1(_07133_),
    .B1(net1197),
    .A1(\stack[27][0] ),
    .Y(_07134_),
    .A2(net796));
 sg13g2_nand2b_1 _25826_ (.Y(_07135_),
    .B(\stack[28][0] ),
    .A_N(net867));
 sg13g2_nand2_1 _25827_ (.Y(_07136_),
    .A(net874),
    .B(\stack[31][0] ));
 sg13g2_a22oi_1 _25828_ (.Y(_07137_),
    .B1(_07136_),
    .B2(_07122_),
    .A2(_07135_),
    .A1(_07109_));
 sg13g2_a221oi_1 _25829_ (.B2(\stack[29][0] ),
    .C1(_07137_),
    .B1(net574),
    .A1(\stack[30][0] ),
    .Y(_07138_),
    .A2(net865));
 sg13g2_xnor2_1 _25830_ (.Y(_07139_),
    .A(_09633_),
    .B(_07122_));
 sg13g2_buf_2 _25831_ (.A(_07139_),
    .X(_07140_));
 sg13g2_nor2_1 _25832_ (.A(_07140_),
    .B(_07127_),
    .Y(_07141_));
 sg13g2_o21ai_1 _25833_ (.B1(_07141_),
    .Y(_07142_),
    .A1(_07134_),
    .A2(_07138_));
 sg13g2_nand2b_1 _25834_ (.Y(_07143_),
    .B(\stack[10][0] ),
    .A_N(net1195));
 sg13g2_nand2_1 _25835_ (.Y(_07144_),
    .A(net867),
    .B(\stack[9][0] ));
 sg13g2_a22oi_1 _25836_ (.Y(_07145_),
    .B1(_07144_),
    .B2(_09694_),
    .A2(_07143_),
    .A1(_07116_));
 sg13g2_a221oi_1 _25837_ (.B2(\stack[8][0] ),
    .C1(_07145_),
    .B1(net1197),
    .A1(\stack[11][0] ),
    .Y(_07146_),
    .A2(net796));
 sg13g2_nand2b_1 _25838_ (.Y(_07147_),
    .B(\stack[12][0] ),
    .A_N(net1195));
 sg13g2_nand2_1 _25839_ (.Y(_07148_),
    .A(net864),
    .B(\stack[15][0] ));
 sg13g2_a22oi_1 _25840_ (.Y(_07149_),
    .B1(_07148_),
    .B2(_07122_),
    .A2(_07147_),
    .A1(_07109_));
 sg13g2_a221oi_1 _25841_ (.B2(\stack[13][0] ),
    .C1(_07149_),
    .B1(net574),
    .A1(\stack[14][0] ),
    .Y(_07150_),
    .A2(net865));
 sg13g2_xnor2_1 _25842_ (.Y(_07151_),
    .A(_09652_),
    .B(_07125_));
 sg13g2_buf_2 _25843_ (.A(_07151_),
    .X(_07152_));
 sg13g2_nor2_1 _25844_ (.A(_07140_),
    .B(_07152_),
    .Y(_07153_));
 sg13g2_o21ai_1 _25845_ (.B1(_07153_),
    .Y(_07154_),
    .A1(_07146_),
    .A2(_07150_));
 sg13g2_buf_8 _25846_ (.A(_07140_),
    .X(_07155_));
 sg13g2_mux4_1 _25847_ (.S0(net1199),
    .A0(\stack[7][0] ),
    .A1(\stack[1][0] ),
    .A2(\stack[3][0] ),
    .A3(\stack[5][0] ),
    .S1(net861),
    .X(_07156_));
 sg13g2_nand2_1 _25848_ (.Y(_07157_),
    .A(net788),
    .B(_07156_));
 sg13g2_mux4_1 _25849_ (.S0(_09702_),
    .A0(\stack[6][0] ),
    .A1(\stack[0][0] ),
    .A2(\stack[2][0] ),
    .A3(\stack[4][0] ),
    .S1(_09746_),
    .X(_07158_));
 sg13g2_nand2_1 _25850_ (.Y(_07159_),
    .A(net785),
    .B(_07158_));
 sg13g2_nand4_1 _25851_ (.B(_07127_),
    .C(_07157_),
    .A(net536),
    .Y(_07160_),
    .D(_07159_));
 sg13g2_nand4_1 _25852_ (.B(_07142_),
    .C(_07154_),
    .A(_07129_),
    .Y(_07161_),
    .D(_07160_));
 sg13g2_buf_1 _25853_ (.A(_07161_),
    .X(_07162_));
 sg13g2_buf_2 _25854_ (.A(_07162_),
    .X(_07163_));
 sg13g2_nand2_1 _25855_ (.Y(_07164_),
    .A(_05441_),
    .B(net781));
 sg13g2_o21ai_1 _25856_ (.B1(_07164_),
    .Y(_02474_),
    .A1(net781),
    .A2(_07163_));
 sg13g2_nor3_1 _25857_ (.A(_09632_),
    .B(_09670_),
    .C(_09743_),
    .Y(_07165_));
 sg13g2_inv_1 _25858_ (.Y(_07166_),
    .A(_09623_));
 sg13g2_o21ai_1 _25859_ (.B1(net861),
    .Y(_07167_),
    .A1(net864),
    .A2(\stack[2][1] ));
 sg13g2_nand2b_1 _25860_ (.Y(_07168_),
    .B(net1311),
    .A_N(_09634_));
 sg13g2_buf_2 _25861_ (.A(_07168_),
    .X(_07169_));
 sg13g2_or2_1 _25862_ (.X(_07170_),
    .B(\stack[3][1] ),
    .A(_09661_));
 sg13g2_o21ai_1 _25863_ (.B1(_07170_),
    .Y(_07171_),
    .A1(\stack[1][1] ),
    .A2(_07169_));
 sg13g2_or3_1 _25864_ (.A(net1200),
    .B(net1201),
    .C(\stack[0][1] ),
    .X(_07172_));
 sg13g2_nand3_1 _25865_ (.B(_09652_),
    .C(_07172_),
    .A(_09632_),
    .Y(_07173_));
 sg13g2_a221oi_1 _25866_ (.B2(_09735_),
    .C1(_07173_),
    .B1(_07171_),
    .A1(_07166_),
    .Y(_07174_),
    .A2(_07167_));
 sg13g2_or2_1 _25867_ (.X(_07175_),
    .B(_07174_),
    .A(_07165_));
 sg13g2_buf_1 _25868_ (.A(net796),
    .X(_07176_));
 sg13g2_inv_1 _25869_ (.Y(_07177_),
    .A(\stack[6][1] ));
 sg13g2_buf_1 _25870_ (.A(_07122_),
    .X(_07178_));
 sg13g2_buf_1 _25871_ (.A(_09681_),
    .X(_07179_));
 sg13g2_o21ai_1 _25872_ (.B1(_09742_),
    .Y(_07180_),
    .A1(\stack[5][1] ),
    .A2(net794));
 sg13g2_nand3b_1 _25873_ (.B(_09675_),
    .C(net1279),
    .Y(_07181_),
    .A_N(net1282));
 sg13g2_buf_2 _25874_ (.A(_07181_),
    .X(_07182_));
 sg13g2_nor2_1 _25875_ (.A(\stack[4][1] ),
    .B(_07182_),
    .Y(_07183_));
 sg13g2_a221oi_1 _25876_ (.B2(net784),
    .C1(_07183_),
    .B1(_07180_),
    .A1(_07177_),
    .Y(_07184_),
    .A2(net795));
 sg13g2_a21o_1 _25877_ (.A2(net573),
    .A1(\stack[7][1] ),
    .B1(_07184_),
    .X(_07185_));
 sg13g2_xnor2_1 _25878_ (.Y(_07186_),
    .A(_09622_),
    .B(_09677_));
 sg13g2_buf_1 _25879_ (.A(_07186_),
    .X(_07187_));
 sg13g2_buf_1 _25880_ (.A(_07187_),
    .X(_07188_));
 sg13g2_mux4_1 _25881_ (.S0(_09617_),
    .A0(\stack[18][1] ),
    .A1(\stack[19][1] ),
    .A2(\stack[16][1] ),
    .A3(\stack[17][1] ),
    .S1(_09624_),
    .X(_07189_));
 sg13g2_nor2_1 _25882_ (.A(net572),
    .B(_07189_),
    .Y(_07190_));
 sg13g2_nor3_1 _25883_ (.A(_07124_),
    .B(_07127_),
    .C(_07190_),
    .Y(_07191_));
 sg13g2_inv_1 _25884_ (.Y(_07192_),
    .A(\stack[22][1] ));
 sg13g2_o21ai_1 _25885_ (.B1(net863),
    .Y(_07193_),
    .A1(\stack[21][1] ),
    .A2(net794));
 sg13g2_nor2_1 _25886_ (.A(\stack[20][1] ),
    .B(_07182_),
    .Y(_07194_));
 sg13g2_a221oi_1 _25887_ (.B2(_09618_),
    .C1(_07194_),
    .B1(_07193_),
    .A1(_07192_),
    .Y(_07195_),
    .A2(net795));
 sg13g2_a21o_1 _25888_ (.A2(net573),
    .A1(\stack[23][1] ),
    .B1(_07195_),
    .X(_07196_));
 sg13g2_a22oi_1 _25889_ (.Y(_07197_),
    .B1(_07191_),
    .B2(_07196_),
    .A2(_07185_),
    .A1(_07175_));
 sg13g2_buf_1 _25890_ (.A(_07197_),
    .X(_07198_));
 sg13g2_a21oi_1 _25891_ (.A1(net870),
    .A2(\stack[12][1] ),
    .Y(_07199_),
    .B1(net794));
 sg13g2_a21oi_1 _25892_ (.A1(net874),
    .A2(\stack[15][1] ),
    .Y(_07200_),
    .B1(_09742_));
 sg13g2_or2_1 _25893_ (.X(_07201_),
    .B(_07200_),
    .A(_07199_));
 sg13g2_a22oi_1 _25894_ (.Y(_07202_),
    .B1(_09686_),
    .B2(\stack[13][1] ),
    .A2(net865),
    .A1(\stack[14][1] ));
 sg13g2_inv_1 _25895_ (.Y(_07203_),
    .A(\stack[9][1] ));
 sg13g2_a21oi_1 _25896_ (.A1(_07203_),
    .A2(_09694_),
    .Y(_07204_),
    .B1(_07116_));
 sg13g2_inv_1 _25897_ (.Y(_07205_),
    .A(_09687_));
 sg13g2_nor2_1 _25898_ (.A(net1198),
    .B(\stack[8][1] ),
    .Y(_07206_));
 sg13g2_a22oi_1 _25899_ (.Y(_07207_),
    .B1(_07206_),
    .B2(net1197),
    .A2(_07116_),
    .A1(_07205_));
 sg13g2_o21ai_1 _25900_ (.B1(_07207_),
    .Y(_07208_),
    .A1(net870),
    .A2(_07204_));
 sg13g2_nand2_1 _25901_ (.Y(_07209_),
    .A(\stack[11][1] ),
    .B(net796));
 sg13g2_a221oi_1 _25902_ (.B2(_07209_),
    .C1(_07152_),
    .B1(_07208_),
    .A1(_07201_),
    .Y(_07210_),
    .A2(_07202_));
 sg13g2_xor2_1 _25903_ (.B(net1201),
    .A(net1280),
    .X(_07211_));
 sg13g2_buf_4 _25904_ (.X(_07212_),
    .A(_07211_));
 sg13g2_mux4_1 _25905_ (.S0(net867),
    .A0(\stack[30][1] ),
    .A1(\stack[31][1] ),
    .A2(\stack[28][1] ),
    .A3(\stack[29][1] ),
    .S1(net862),
    .X(_07213_));
 sg13g2_nor2_1 _25906_ (.A(_07212_),
    .B(_07213_),
    .Y(_07214_));
 sg13g2_and2_1 _25907_ (.A(net862),
    .B(\stack[25][1] ),
    .X(_07215_));
 sg13g2_nand2_1 _25908_ (.Y(_07216_),
    .A(net867),
    .B(\stack[27][1] ));
 sg13g2_nand2b_1 _25909_ (.Y(_07217_),
    .B(\stack[24][1] ),
    .A_N(net867));
 sg13g2_a22oi_1 _25910_ (.Y(_07218_),
    .B1(_07217_),
    .B2(_09694_),
    .A2(_07216_),
    .A1(_07116_));
 sg13g2_a221oi_1 _25911_ (.B2(net788),
    .C1(_07218_),
    .B1(_07215_),
    .A1(\stack[26][1] ),
    .Y(_07219_),
    .A2(net865));
 sg13g2_nor3_1 _25912_ (.A(_07127_),
    .B(_07214_),
    .C(_07219_),
    .Y(_07220_));
 sg13g2_o21ai_1 _25913_ (.B1(_07124_),
    .Y(_07221_),
    .A1(_07210_),
    .A2(_07220_));
 sg13g2_buf_1 _25914_ (.A(_07221_),
    .X(_07222_));
 sg13g2_nand2_1 _25915_ (.Y(_07223_),
    .A(_07198_),
    .B(_07222_));
 sg13g2_buf_2 _25916_ (.A(_07223_),
    .X(_07224_));
 sg13g2_mux2_1 _25917_ (.A0(_07224_),
    .A1(_05446_),
    .S(net781),
    .X(_02475_));
 sg13g2_buf_1 _25918_ (.A(_07127_),
    .X(_07225_));
 sg13g2_and2_1 _25919_ (.A(\stack[7][2] ),
    .B(net796),
    .X(_07226_));
 sg13g2_inv_1 _25920_ (.Y(_07227_),
    .A(\stack[6][2] ));
 sg13g2_o21ai_1 _25921_ (.B1(_09742_),
    .Y(_07228_),
    .A1(\stack[5][2] ),
    .A2(net794));
 sg13g2_nor2_1 _25922_ (.A(\stack[4][2] ),
    .B(_07182_),
    .Y(_07229_));
 sg13g2_a221oi_1 _25923_ (.B2(net786),
    .C1(_07229_),
    .B1(_07228_),
    .A1(_07227_),
    .Y(_07230_),
    .A2(_07178_));
 sg13g2_inv_1 _25924_ (.Y(_07231_),
    .A(\stack[2][2] ));
 sg13g2_and2_1 _25925_ (.A(net1198),
    .B(_09719_),
    .X(_07232_));
 sg13g2_buf_2 _25926_ (.A(_07232_),
    .X(_07233_));
 sg13g2_buf_1 _25927_ (.A(_07169_),
    .X(_07234_));
 sg13g2_o21ai_1 _25928_ (.B1(net793),
    .Y(_07235_),
    .A1(\stack[3][2] ),
    .A2(net866));
 sg13g2_nor2_1 _25929_ (.A(\stack[0][2] ),
    .B(net793),
    .Y(_07236_));
 sg13g2_a221oi_1 _25930_ (.B2(net788),
    .C1(_07236_),
    .B1(_07235_),
    .A1(_07231_),
    .Y(_07237_),
    .A2(_07233_));
 sg13g2_o21ai_1 _25931_ (.B1(_07237_),
    .Y(_07238_),
    .A1(_07226_),
    .A2(_07230_));
 sg13g2_nand3_1 _25932_ (.B(net574),
    .C(_07230_),
    .A(\stack[1][2] ),
    .Y(_07239_));
 sg13g2_nand4_1 _25933_ (.B(_07225_),
    .C(_07238_),
    .A(net536),
    .Y(_07240_),
    .D(_07239_));
 sg13g2_mux4_1 _25934_ (.S0(net874),
    .A0(\stack[30][2] ),
    .A1(\stack[31][2] ),
    .A2(\stack[28][2] ),
    .A3(\stack[29][2] ),
    .S1(net873),
    .X(_07241_));
 sg13g2_nand2_1 _25935_ (.Y(_07242_),
    .A(net572),
    .B(_07241_));
 sg13g2_mux4_1 _25936_ (.S0(net864),
    .A0(\stack[26][2] ),
    .A1(\stack[27][2] ),
    .A2(\stack[24][2] ),
    .A3(\stack[25][2] ),
    .S1(net873),
    .X(_07243_));
 sg13g2_nand2_1 _25937_ (.Y(_07244_),
    .A(_07212_),
    .B(_07243_));
 sg13g2_a21oi_1 _25938_ (.A1(_07242_),
    .A2(_07244_),
    .Y(_07245_),
    .B1(net535));
 sg13g2_inv_1 _25939_ (.Y(_07246_),
    .A(\stack[15][2] ));
 sg13g2_a21oi_1 _25940_ (.A1(_07246_),
    .A2(net795),
    .Y(_07247_),
    .B1(_07109_));
 sg13g2_inv_1 _25941_ (.Y(_07248_),
    .A(\stack[14][2] ));
 sg13g2_inv_1 _25942_ (.Y(_07249_),
    .A(\stack[12][2] ));
 sg13g2_a22oi_1 _25943_ (.Y(_07250_),
    .B1(_07109_),
    .B2(_07249_),
    .A2(_09635_),
    .A1(_07248_));
 sg13g2_o21ai_1 _25944_ (.B1(_07250_),
    .Y(_07251_),
    .A1(net785),
    .A2(_07247_));
 sg13g2_nand2_1 _25945_ (.Y(_07252_),
    .A(\stack[13][2] ),
    .B(net574));
 sg13g2_mux4_1 _25946_ (.S0(net864),
    .A0(\stack[10][2] ),
    .A1(\stack[11][2] ),
    .A2(\stack[8][2] ),
    .A3(\stack[9][2] ),
    .S1(net873),
    .X(_07253_));
 sg13g2_o21ai_1 _25947_ (.B1(_07127_),
    .Y(_07254_),
    .A1(net572),
    .A2(_07253_));
 sg13g2_a21oi_1 _25948_ (.A1(_07251_),
    .A2(_07252_),
    .Y(_07255_),
    .B1(_07254_));
 sg13g2_or3_1 _25949_ (.A(net536),
    .B(_07245_),
    .C(_07255_),
    .X(_07256_));
 sg13g2_mux4_1 _25950_ (.S0(_09714_),
    .A0(\stack[22][2] ),
    .A1(\stack[23][2] ),
    .A2(\stack[20][2] ),
    .A3(\stack[21][2] ),
    .S1(net860),
    .X(_07257_));
 sg13g2_nor2_1 _25951_ (.A(_07212_),
    .B(_07257_),
    .Y(_07258_));
 sg13g2_inv_1 _25952_ (.Y(_07259_),
    .A(\stack[16][2] ));
 sg13g2_nor2b_1 _25953_ (.A(net1279),
    .B_N(net1197),
    .Y(_07260_));
 sg13g2_buf_8 _25954_ (.A(_07260_),
    .X(_07261_));
 sg13g2_o21ai_1 _25955_ (.B1(net866),
    .Y(_07262_),
    .A1(\stack[17][2] ),
    .A2(_07169_));
 sg13g2_buf_8 _25956_ (.A(net866),
    .X(_07263_));
 sg13g2_nor2_1 _25957_ (.A(\stack[18][2] ),
    .B(net571),
    .Y(_07264_));
 sg13g2_a221oi_1 _25958_ (.B2(net788),
    .C1(_07264_),
    .B1(_07262_),
    .A1(_07259_),
    .Y(_07265_),
    .A2(_07261_));
 sg13g2_a21oi_1 _25959_ (.A1(\stack[19][2] ),
    .A2(net573),
    .Y(_07266_),
    .B1(_07265_));
 sg13g2_o21ai_1 _25960_ (.B1(_07128_),
    .Y(_07267_),
    .A1(_07258_),
    .A2(_07266_));
 sg13g2_nand3_1 _25961_ (.B(_07256_),
    .C(_07267_),
    .A(_07240_),
    .Y(_07268_));
 sg13g2_buf_2 _25962_ (.A(_07268_),
    .X(_07269_));
 sg13g2_nand2_1 _25963_ (.Y(_07270_),
    .A(_05449_),
    .B(net859));
 sg13g2_o21ai_1 _25964_ (.B1(_07270_),
    .Y(_02476_),
    .A1(net781),
    .A2(_07269_));
 sg13g2_inv_1 _25965_ (.Y(_07271_),
    .A(\stack[16][3] ));
 sg13g2_o21ai_1 _25966_ (.B1(_07263_),
    .Y(_07272_),
    .A1(\stack[17][3] ),
    .A2(_07234_));
 sg13g2_nor2_1 _25967_ (.A(\stack[18][3] ),
    .B(_07263_),
    .Y(_07273_));
 sg13g2_a221oi_1 _25968_ (.B2(net560),
    .C1(_07273_),
    .B1(_07272_),
    .A1(_07271_),
    .Y(_07274_),
    .A2(_07261_));
 sg13g2_a21oi_1 _25969_ (.A1(\stack[19][3] ),
    .A2(net573),
    .Y(_07275_),
    .B1(_07274_));
 sg13g2_mux4_1 _25970_ (.S0(net784),
    .A0(\stack[22][3] ),
    .A1(\stack[23][3] ),
    .A2(\stack[20][3] ),
    .A3(\stack[21][3] ),
    .S1(net787),
    .X(_07276_));
 sg13g2_o21ai_1 _25971_ (.B1(_07152_),
    .Y(_07277_),
    .A1(_07212_),
    .A2(_07276_));
 sg13g2_nor2_1 _25972_ (.A(_07275_),
    .B(_07277_),
    .Y(_07278_));
 sg13g2_inv_1 _25973_ (.Y(_07279_),
    .A(\stack[6][3] ));
 sg13g2_o21ai_1 _25974_ (.B1(net863),
    .Y(_07280_),
    .A1(\stack[5][3] ),
    .A2(_07179_));
 sg13g2_nor2_1 _25975_ (.A(\stack[4][3] ),
    .B(_07182_),
    .Y(_07281_));
 sg13g2_a221oi_1 _25976_ (.B2(net560),
    .C1(_07281_),
    .B1(_07280_),
    .A1(_07279_),
    .Y(_07282_),
    .A2(net795));
 sg13g2_a21oi_1 _25977_ (.A1(\stack[7][3] ),
    .A2(net573),
    .Y(_07283_),
    .B1(_07282_));
 sg13g2_mux4_1 _25978_ (.S0(_09735_),
    .A0(\stack[2][3] ),
    .A1(\stack[3][3] ),
    .A2(\stack[0][3] ),
    .A3(\stack[1][3] ),
    .S1(_09853_),
    .X(_07284_));
 sg13g2_o21ai_1 _25979_ (.B1(_07225_),
    .Y(_07285_),
    .A1(net572),
    .A2(_07284_));
 sg13g2_o21ai_1 _25980_ (.B1(net536),
    .Y(_07286_),
    .A1(_07283_),
    .A2(_07285_));
 sg13g2_inv_1 _25981_ (.Y(_07287_),
    .A(\stack[24][3] ));
 sg13g2_o21ai_1 _25982_ (.B1(net571),
    .Y(_07288_),
    .A1(\stack[25][3] ),
    .A2(net793));
 sg13g2_nor2_1 _25983_ (.A(\stack[26][3] ),
    .B(net571),
    .Y(_07289_));
 sg13g2_a221oi_1 _25984_ (.B2(net560),
    .C1(_07289_),
    .B1(_07288_),
    .A1(_07287_),
    .Y(_07290_),
    .A2(_07261_));
 sg13g2_and2_1 _25985_ (.A(\stack[27][3] ),
    .B(net796),
    .X(_07291_));
 sg13g2_mux4_1 _25986_ (.S0(net869),
    .A0(\stack[30][3] ),
    .A1(\stack[31][3] ),
    .A2(\stack[28][3] ),
    .A3(\stack[29][3] ),
    .S1(net860),
    .X(_07292_));
 sg13g2_nand2b_1 _25987_ (.Y(_07293_),
    .B(net572),
    .A_N(_07292_));
 sg13g2_o21ai_1 _25988_ (.B1(_07293_),
    .Y(_07294_),
    .A1(_07290_),
    .A2(_07291_));
 sg13g2_o21ai_1 _25989_ (.B1(net863),
    .Y(_07295_),
    .A1(\stack[12][3] ),
    .A2(net794));
 sg13g2_nand3_1 _25990_ (.B(net1280),
    .C(net1201),
    .A(net1206),
    .Y(_07296_));
 sg13g2_buf_2 _25991_ (.A(_07296_),
    .X(_07297_));
 sg13g2_or3_1 _25992_ (.A(net1202),
    .B(net861),
    .C(\stack[15][3] ),
    .X(_07298_));
 sg13g2_o21ai_1 _25993_ (.B1(_07298_),
    .Y(_07299_),
    .A1(\stack[13][3] ),
    .A2(_07297_));
 sg13g2_a21oi_1 _25994_ (.A1(net785),
    .A2(_07295_),
    .Y(_07300_),
    .B1(_07299_));
 sg13g2_and2_1 _25995_ (.A(\stack[14][3] ),
    .B(net865),
    .X(_07301_));
 sg13g2_inv_1 _25996_ (.Y(_07302_),
    .A(\stack[10][3] ));
 sg13g2_o21ai_1 _25997_ (.B1(net793),
    .Y(_07303_),
    .A1(\stack[11][3] ),
    .A2(net571));
 sg13g2_nor2_1 _25998_ (.A(\stack[8][3] ),
    .B(net793),
    .Y(_07304_));
 sg13g2_a221oi_1 _25999_ (.B2(net561),
    .C1(_07304_),
    .B1(_07303_),
    .A1(_07302_),
    .Y(_07305_),
    .A2(_07233_));
 sg13g2_o21ai_1 _26000_ (.B1(_07305_),
    .Y(_07306_),
    .A1(_07300_),
    .A2(_07301_));
 sg13g2_inv_1 _26001_ (.Y(_07307_),
    .A(\stack[9][3] ));
 sg13g2_nor4_1 _26002_ (.A(net785),
    .B(_07166_),
    .C(_07307_),
    .D(_07299_),
    .Y(_07308_));
 sg13g2_nor2b_1 _26003_ (.A(_07308_),
    .B_N(_07153_),
    .Y(_07309_));
 sg13g2_a22oi_1 _26004_ (.Y(_07310_),
    .B1(_07306_),
    .B2(_07309_),
    .A2(_07294_),
    .A1(_07141_));
 sg13g2_o21ai_1 _26005_ (.B1(_07310_),
    .Y(_07311_),
    .A1(_07278_),
    .A2(_07286_));
 sg13g2_buf_1 _26006_ (.A(_07311_),
    .X(_07312_));
 sg13g2_buf_1 _26007_ (.A(_07312_),
    .X(_07313_));
 sg13g2_nand2_1 _26008_ (.Y(_07314_),
    .A(_05453_),
    .B(net859));
 sg13g2_o21ai_1 _26009_ (.B1(_07314_),
    .Y(_02477_),
    .A1(net781),
    .A2(_07313_));
 sg13g2_inv_1 _26010_ (.Y(_07315_),
    .A(\stack[26][4] ));
 sg13g2_mux2_1 _26011_ (.A0(\stack[24][4] ),
    .A1(\stack[28][4] ),
    .S(_09678_),
    .X(_07316_));
 sg13g2_or3_1 _26012_ (.A(net1204),
    .B(net1198),
    .C(\stack[30][4] ),
    .X(_07317_));
 sg13g2_o21ai_1 _26013_ (.B1(_07317_),
    .Y(_07318_),
    .A1(_07166_),
    .A2(_07316_));
 sg13g2_mux2_1 _26014_ (.A0(\stack[25][4] ),
    .A1(\stack[29][4] ),
    .S(_09678_),
    .X(_07319_));
 sg13g2_a221oi_1 _26015_ (.B2(net862),
    .C1(net870),
    .B1(_07319_),
    .A1(_09858_),
    .Y(_07320_),
    .A2(_07122_));
 sg13g2_a221oi_1 _26016_ (.B2(_09683_),
    .C1(_07320_),
    .B1(_07318_),
    .A1(_07315_),
    .Y(_07321_),
    .A2(_07116_));
 sg13g2_nor2_1 _26017_ (.A(_09633_),
    .B(_09858_),
    .Y(_07322_));
 sg13g2_nor2_1 _26018_ (.A(net1198),
    .B(_09632_),
    .Y(_07323_));
 sg13g2_a221oi_1 _26019_ (.B2(_09632_),
    .C1(_07323_),
    .B1(_09742_),
    .A1(_09696_),
    .Y(_07324_),
    .A2(\stack[27][4] ));
 sg13g2_a221oi_1 _26020_ (.B2(_07322_),
    .C1(_07324_),
    .B1(net795),
    .A1(net860),
    .Y(_07325_),
    .A2(_09633_));
 sg13g2_mux4_1 _26021_ (.S0(net1200),
    .A0(\stack[22][4] ),
    .A1(\stack[23][4] ),
    .A2(\stack[20][4] ),
    .A3(\stack[21][4] ),
    .S1(net1202),
    .X(_07326_));
 sg13g2_nand2_1 _26022_ (.Y(_07327_),
    .A(_07187_),
    .B(_07326_));
 sg13g2_mux4_1 _26023_ (.S0(_09695_),
    .A0(\stack[18][4] ),
    .A1(\stack[19][4] ),
    .A2(\stack[16][4] ),
    .A3(\stack[17][4] ),
    .S1(net1202),
    .X(_07328_));
 sg13g2_nand2_1 _26024_ (.Y(_07329_),
    .A(_07212_),
    .B(_07328_));
 sg13g2_nand3_1 _26025_ (.B(_07327_),
    .C(_07329_),
    .A(_07155_),
    .Y(_07330_));
 sg13g2_o21ai_1 _26026_ (.B1(_07330_),
    .Y(_07331_),
    .A1(_07321_),
    .A2(_07325_));
 sg13g2_mux4_1 _26027_ (.S0(net1195),
    .A0(\stack[14][4] ),
    .A1(\stack[15][4] ),
    .A2(\stack[12][4] ),
    .A3(\stack[13][4] ),
    .S1(net862),
    .X(_07332_));
 sg13g2_mux4_1 _26028_ (.S0(net1195),
    .A0(\stack[10][4] ),
    .A1(\stack[11][4] ),
    .A2(\stack[8][4] ),
    .A3(\stack[9][4] ),
    .S1(net862),
    .X(_07333_));
 sg13g2_mux4_1 _26029_ (.S0(net1195),
    .A0(\stack[6][4] ),
    .A1(\stack[7][4] ),
    .A2(\stack[4][4] ),
    .A3(\stack[5][4] ),
    .S1(net1202),
    .X(_07334_));
 sg13g2_mux4_1 _26030_ (.S0(_09783_),
    .A0(\stack[2][4] ),
    .A1(\stack[3][4] ),
    .A2(\stack[0][4] ),
    .A3(\stack[1][4] ),
    .S1(net1202),
    .X(_07335_));
 sg13g2_mux4_1 _26031_ (.S0(_07212_),
    .A0(_07332_),
    .A1(_07333_),
    .A2(_07334_),
    .A3(_07335_),
    .S1(_07140_),
    .X(_07336_));
 sg13g2_nand2_1 _26032_ (.Y(_07337_),
    .A(net535),
    .B(_07336_));
 sg13g2_o21ai_1 _26033_ (.B1(_07337_),
    .Y(_07338_),
    .A1(net535),
    .A2(_07331_));
 sg13g2_buf_2 _26034_ (.A(_07338_),
    .X(_07339_));
 sg13g2_inv_1 _26035_ (.Y(_07340_),
    .A(_07339_));
 sg13g2_nand2_1 _26036_ (.Y(_07341_),
    .A(_05457_),
    .B(net859));
 sg13g2_o21ai_1 _26037_ (.B1(_07341_),
    .Y(_02478_),
    .A1(net781),
    .A2(_07340_));
 sg13g2_inv_1 _26038_ (.Y(_07342_),
    .A(\stack[24][5] ));
 sg13g2_o21ai_1 _26039_ (.B1(net866),
    .Y(_07343_),
    .A1(\stack[25][5] ),
    .A2(_07169_));
 sg13g2_nor2_1 _26040_ (.A(\stack[26][5] ),
    .B(net571),
    .Y(_07344_));
 sg13g2_a221oi_1 _26041_ (.B2(net560),
    .C1(_07344_),
    .B1(_07343_),
    .A1(_07342_),
    .Y(_07345_),
    .A2(_07261_));
 sg13g2_and2_1 _26042_ (.A(\stack[27][5] ),
    .B(_07176_),
    .X(_07346_));
 sg13g2_inv_1 _26043_ (.Y(_07347_),
    .A(\stack[28][5] ));
 sg13g2_o21ai_1 _26044_ (.B1(net794),
    .Y(_07348_),
    .A1(\stack[31][5] ),
    .A2(net863));
 sg13g2_nor2_1 _26045_ (.A(\stack[30][5] ),
    .B(net871),
    .Y(_07349_));
 sg13g2_a221oi_1 _26046_ (.B2(net561),
    .C1(_07349_),
    .B1(_07348_),
    .A1(_07347_),
    .Y(_07350_),
    .A2(_07109_));
 sg13g2_o21ai_1 _26047_ (.B1(_07350_),
    .Y(_07351_),
    .A1(_07345_),
    .A2(_07346_));
 sg13g2_nand3_1 _26048_ (.B(net574),
    .C(_07345_),
    .A(\stack[29][5] ),
    .Y(_07352_));
 sg13g2_a21o_1 _26049_ (.A2(_07352_),
    .A1(_07351_),
    .B1(net535),
    .X(_07353_));
 sg13g2_inv_1 _26050_ (.Y(_07354_),
    .A(\stack[14][5] ));
 sg13g2_o21ai_1 _26051_ (.B1(net863),
    .Y(_07355_),
    .A1(\stack[13][5] ),
    .A2(net794));
 sg13g2_nor2_1 _26052_ (.A(\stack[12][5] ),
    .B(_07182_),
    .Y(_07356_));
 sg13g2_a221oi_1 _26053_ (.B2(net561),
    .C1(_07356_),
    .B1(_07355_),
    .A1(_07354_),
    .Y(_07357_),
    .A2(net795));
 sg13g2_a21o_1 _26054_ (.A2(net573),
    .A1(\stack[15][5] ),
    .B1(_07357_),
    .X(_07358_));
 sg13g2_mux4_1 _26055_ (.S0(net784),
    .A0(\stack[10][5] ),
    .A1(\stack[11][5] ),
    .A2(\stack[8][5] ),
    .A3(\stack[9][5] ),
    .S1(net860),
    .X(_07359_));
 sg13g2_nor2_1 _26056_ (.A(net572),
    .B(_07359_),
    .Y(_07360_));
 sg13g2_nor2_1 _26057_ (.A(_07152_),
    .B(_07360_),
    .Y(_07361_));
 sg13g2_a21oi_1 _26058_ (.A1(_07358_),
    .A2(_07361_),
    .Y(_07362_),
    .B1(net536));
 sg13g2_nand2_1 _26059_ (.Y(_07363_),
    .A(_07353_),
    .B(_07362_));
 sg13g2_inv_1 _26060_ (.Y(_07364_),
    .A(\stack[16][5] ));
 sg13g2_o21ai_1 _26061_ (.B1(net571),
    .Y(_07365_),
    .A1(\stack[17][5] ),
    .A2(_07234_));
 sg13g2_nor2_1 _26062_ (.A(\stack[18][5] ),
    .B(net571),
    .Y(_07366_));
 sg13g2_a221oi_1 _26063_ (.B2(_09823_),
    .C1(_07366_),
    .B1(_07365_),
    .A1(_07364_),
    .Y(_07367_),
    .A2(_07261_));
 sg13g2_inv_1 _26064_ (.Y(_07368_),
    .A(\stack[22][5] ));
 sg13g2_o21ai_1 _26065_ (.B1(_09743_),
    .Y(_07369_),
    .A1(\stack[21][5] ),
    .A2(_07179_));
 sg13g2_nor2_1 _26066_ (.A(\stack[20][5] ),
    .B(_07182_),
    .Y(_07370_));
 sg13g2_a221oi_1 _26067_ (.B2(_09823_),
    .C1(_07370_),
    .B1(_07369_),
    .A1(_07368_),
    .Y(_07371_),
    .A2(_07178_));
 sg13g2_a21oi_1 _26068_ (.A1(_07367_),
    .A2(_07371_),
    .Y(_07372_),
    .B1(_07176_));
 sg13g2_nor2_1 _26069_ (.A(\stack[19][5] ),
    .B(_07367_),
    .Y(_07373_));
 sg13g2_o21ai_1 _26070_ (.B1(_07152_),
    .Y(_07374_),
    .A1(\stack[23][5] ),
    .A2(_07371_));
 sg13g2_or3_1 _26071_ (.A(_07372_),
    .B(_07373_),
    .C(_07374_),
    .X(_07375_));
 sg13g2_inv_1 _26072_ (.Y(_07376_),
    .A(\stack[2][5] ));
 sg13g2_o21ai_1 _26073_ (.B1(net793),
    .Y(_07377_),
    .A1(\stack[3][5] ),
    .A2(net571));
 sg13g2_nor2_1 _26074_ (.A(\stack[0][5] ),
    .B(net793),
    .Y(_07378_));
 sg13g2_a221oi_1 _26075_ (.B2(_09812_),
    .C1(_07378_),
    .B1(_07377_),
    .A1(_07376_),
    .Y(_07379_),
    .A2(_07233_));
 sg13g2_a21o_1 _26076_ (.A2(net574),
    .A1(\stack[1][5] ),
    .B1(_07379_),
    .X(_07380_));
 sg13g2_mux4_1 _26077_ (.S0(net784),
    .A0(\stack[6][5] ),
    .A1(\stack[7][5] ),
    .A2(\stack[4][5] ),
    .A3(\stack[5][5] ),
    .S1(_09853_),
    .X(_07381_));
 sg13g2_inv_1 _26078_ (.Y(_07382_),
    .A(_07381_));
 sg13g2_a21oi_1 _26079_ (.A1(_07188_),
    .A2(_07382_),
    .Y(_07383_),
    .B1(_07152_));
 sg13g2_a21oi_1 _26080_ (.A1(_07380_),
    .A2(_07383_),
    .Y(_07384_),
    .B1(_07124_));
 sg13g2_nand2_1 _26081_ (.Y(_07385_),
    .A(_07375_),
    .B(_07384_));
 sg13g2_nand2_1 _26082_ (.Y(_07386_),
    .A(_07363_),
    .B(_07385_));
 sg13g2_buf_2 _26083_ (.A(_07386_),
    .X(_07387_));
 sg13g2_nand2_1 _26084_ (.Y(_07388_),
    .A(_05463_),
    .B(net859));
 sg13g2_o21ai_1 _26085_ (.B1(_07388_),
    .Y(_02479_),
    .A1(net781),
    .A2(_07387_));
 sg13g2_mux4_1 _26086_ (.S0(net864),
    .A0(\stack[30][6] ),
    .A1(\stack[31][6] ),
    .A2(\stack[28][6] ),
    .A3(\stack[29][6] ),
    .S1(net862),
    .X(_07389_));
 sg13g2_mux4_1 _26087_ (.S0(_09734_),
    .A0(\stack[26][6] ),
    .A1(\stack[27][6] ),
    .A2(\stack[24][6] ),
    .A3(\stack[25][6] ),
    .S1(net873),
    .X(_07390_));
 sg13g2_mux4_1 _26088_ (.S0(_09713_),
    .A0(\stack[22][6] ),
    .A1(\stack[23][6] ),
    .A2(\stack[20][6] ),
    .A3(\stack[21][6] ),
    .S1(_09745_),
    .X(_07391_));
 sg13g2_mux4_1 _26089_ (.S0(net867),
    .A0(\stack[18][6] ),
    .A1(\stack[19][6] ),
    .A2(\stack[16][6] ),
    .A3(\stack[17][6] ),
    .S1(_09745_),
    .X(_07392_));
 sg13g2_mux4_1 _26090_ (.S0(_07212_),
    .A0(_07389_),
    .A1(_07390_),
    .A2(_07391_),
    .A3(_07392_),
    .S1(_07155_),
    .X(_07393_));
 sg13g2_or2_1 _26091_ (.X(_07394_),
    .B(_07393_),
    .A(net535));
 sg13g2_buf_1 _26092_ (.A(_07394_),
    .X(_07395_));
 sg13g2_inv_1 _26093_ (.Y(_07396_),
    .A(\stack[14][6] ));
 sg13g2_o21ai_1 _26094_ (.B1(net863),
    .Y(_07397_),
    .A1(\stack[13][6] ),
    .A2(net794));
 sg13g2_nor2_1 _26095_ (.A(\stack[12][6] ),
    .B(_07182_),
    .Y(_07398_));
 sg13g2_a221oi_1 _26096_ (.B2(net788),
    .C1(_07398_),
    .B1(_07397_),
    .A1(_07396_),
    .Y(_07399_),
    .A2(net795));
 sg13g2_and2_1 _26097_ (.A(\stack[15][6] ),
    .B(net796),
    .X(_07400_));
 sg13g2_mux4_1 _26098_ (.S0(net1195),
    .A0(\stack[10][6] ),
    .A1(\stack[11][6] ),
    .A2(\stack[8][6] ),
    .A3(\stack[9][6] ),
    .S1(net862),
    .X(_07401_));
 sg13g2_nor2_1 _26099_ (.A(net572),
    .B(_07401_),
    .Y(_07402_));
 sg13g2_nor2_1 _26100_ (.A(net536),
    .B(_07402_),
    .Y(_07403_));
 sg13g2_o21ai_1 _26101_ (.B1(_07403_),
    .Y(_07404_),
    .A1(_07399_),
    .A2(_07400_));
 sg13g2_inv_1 _26102_ (.Y(_07405_),
    .A(\stack[2][6] ));
 sg13g2_o21ai_1 _26103_ (.B1(_07169_),
    .Y(_07406_),
    .A1(\stack[3][6] ),
    .A2(_09727_));
 sg13g2_nor2_1 _26104_ (.A(\stack[0][6] ),
    .B(net793),
    .Y(_07407_));
 sg13g2_a221oi_1 _26105_ (.B2(_09618_),
    .C1(_07407_),
    .B1(_07406_),
    .A1(_07405_),
    .Y(_07408_),
    .A2(_07233_));
 sg13g2_and2_1 _26106_ (.A(\stack[1][6] ),
    .B(net574),
    .X(_07409_));
 sg13g2_mux4_1 _26107_ (.S0(_09783_),
    .A0(\stack[6][6] ),
    .A1(\stack[7][6] ),
    .A2(\stack[4][6] ),
    .A3(\stack[5][6] ),
    .S1(_09676_),
    .X(_07410_));
 sg13g2_inv_1 _26108_ (.Y(_07411_),
    .A(_07410_));
 sg13g2_a21oi_1 _26109_ (.A1(_07188_),
    .A2(_07411_),
    .Y(_07412_),
    .B1(_07124_));
 sg13g2_o21ai_1 _26110_ (.B1(_07412_),
    .Y(_07413_),
    .A1(_07408_),
    .A2(_07409_));
 sg13g2_nand3_1 _26111_ (.B(_07404_),
    .C(_07413_),
    .A(net535),
    .Y(_07414_));
 sg13g2_buf_1 _26112_ (.A(_07414_),
    .X(_07415_));
 sg13g2_nand2_2 _26113_ (.Y(_07416_),
    .A(_07395_),
    .B(_07415_));
 sg13g2_nand2_1 _26114_ (.Y(_07417_),
    .A(_05467_),
    .B(net859));
 sg13g2_o21ai_1 _26115_ (.B1(_07417_),
    .Y(_02480_),
    .A1(net781),
    .A2(_07416_));
 sg13g2_inv_1 _26116_ (.Y(_07418_),
    .A(\stack[8][7] ));
 sg13g2_o21ai_1 _26117_ (.B1(_09726_),
    .Y(_07419_),
    .A1(\stack[9][7] ),
    .A2(_07169_));
 sg13g2_nor2_1 _26118_ (.A(\stack[10][7] ),
    .B(net866),
    .Y(_07420_));
 sg13g2_a221oi_1 _26119_ (.B2(net869),
    .C1(_07420_),
    .B1(_07419_),
    .A1(_07418_),
    .Y(_07421_),
    .A2(_07261_));
 sg13g2_and2_1 _26120_ (.A(\stack[11][7] ),
    .B(_07130_),
    .X(_07422_));
 sg13g2_mux4_1 _26121_ (.S0(net1200),
    .A0(\stack[14][7] ),
    .A1(\stack[15][7] ),
    .A2(\stack[12][7] ),
    .A3(\stack[13][7] ),
    .S1(net1199),
    .X(_07423_));
 sg13g2_nand2b_1 _26122_ (.Y(_07424_),
    .B(_07187_),
    .A_N(_07423_));
 sg13g2_o21ai_1 _26123_ (.B1(_07424_),
    .Y(_07425_),
    .A1(_07421_),
    .A2(_07422_));
 sg13g2_inv_1 _26124_ (.Y(_07426_),
    .A(\stack[24][7] ));
 sg13g2_o21ai_1 _26125_ (.B1(_09726_),
    .Y(_07427_),
    .A1(\stack[25][7] ),
    .A2(_07169_));
 sg13g2_nor2_1 _26126_ (.A(\stack[26][7] ),
    .B(net866),
    .Y(_07428_));
 sg13g2_a221oi_1 _26127_ (.B2(net869),
    .C1(_07428_),
    .B1(_07427_),
    .A1(_07426_),
    .Y(_07429_),
    .A2(_07261_));
 sg13g2_and2_1 _26128_ (.A(\stack[27][7] ),
    .B(net796),
    .X(_07430_));
 sg13g2_mux4_1 _26129_ (.S0(net1200),
    .A0(\stack[30][7] ),
    .A1(\stack[31][7] ),
    .A2(\stack[28][7] ),
    .A3(\stack[29][7] ),
    .S1(net1199),
    .X(_07431_));
 sg13g2_nand2b_1 _26130_ (.Y(_07432_),
    .B(net572),
    .A_N(_07431_));
 sg13g2_o21ai_1 _26131_ (.B1(_07432_),
    .Y(_07433_),
    .A1(_07429_),
    .A2(_07430_));
 sg13g2_mux4_1 _26132_ (.S0(_09676_),
    .A0(\stack[6][7] ),
    .A1(\stack[0][7] ),
    .A2(\stack[2][7] ),
    .A3(\stack[4][7] ),
    .S1(_09746_),
    .X(_07434_));
 sg13g2_mux4_1 _26133_ (.S0(_09675_),
    .A0(\stack[7][7] ),
    .A1(\stack[1][7] ),
    .A2(\stack[3][7] ),
    .A3(\stack[5][7] ),
    .S1(_09711_),
    .X(_07435_));
 sg13g2_and2_1 _26134_ (.A(_09714_),
    .B(_07435_),
    .X(_07436_));
 sg13g2_a21oi_1 _26135_ (.A1(net785),
    .A2(_07434_),
    .Y(_07437_),
    .B1(_07436_));
 sg13g2_inv_1 _26136_ (.Y(_07438_),
    .A(\stack[16][7] ));
 sg13g2_o21ai_1 _26137_ (.B1(_09726_),
    .Y(_07439_),
    .A1(\stack[17][7] ),
    .A2(_07169_));
 sg13g2_nor2_1 _26138_ (.A(\stack[18][7] ),
    .B(net866),
    .Y(_07440_));
 sg13g2_a221oi_1 _26139_ (.B2(net869),
    .C1(_07440_),
    .B1(_07439_),
    .A1(_07438_),
    .Y(_07441_),
    .A2(_07261_));
 sg13g2_and2_1 _26140_ (.A(\stack[19][7] ),
    .B(_07130_),
    .X(_07442_));
 sg13g2_mux4_1 _26141_ (.S0(_09695_),
    .A0(\stack[22][7] ),
    .A1(\stack[23][7] ),
    .A2(\stack[20][7] ),
    .A3(\stack[21][7] ),
    .S1(_09702_),
    .X(_07443_));
 sg13g2_nand2b_1 _26142_ (.Y(_07444_),
    .B(_07187_),
    .A_N(_07443_));
 sg13g2_o21ai_1 _26143_ (.B1(_07444_),
    .Y(_07445_),
    .A1(_07441_),
    .A2(_07442_));
 sg13g2_mux4_1 _26144_ (.S0(_07152_),
    .A0(_07425_),
    .A1(_07433_),
    .A2(_07437_),
    .A3(_07445_),
    .S1(net536),
    .X(_07446_));
 sg13g2_buf_2 _26145_ (.A(_07446_),
    .X(_07447_));
 sg13g2_nand2_1 _26146_ (.Y(_07448_),
    .A(_05471_),
    .B(_09911_));
 sg13g2_o21ai_1 _26147_ (.B1(_07448_),
    .Y(_02481_),
    .A1(_10080_),
    .A2(_07447_));
 sg13g2_mux2_1 _26148_ (.A0(\exec.memory_input[0] ),
    .A1(_10047_),
    .S(_10030_),
    .X(_02482_));
 sg13g2_mux2_1 _26149_ (.A0(\exec.memory_input[1] ),
    .A1(_10041_),
    .S(net783),
    .X(_02483_));
 sg13g2_mux2_1 _26150_ (.A0(\exec.memory_input[2] ),
    .A1(_10052_),
    .S(net783),
    .X(_02484_));
 sg13g2_mux2_1 _26151_ (.A0(\exec.memory_input[3] ),
    .A1(_10049_),
    .S(net783),
    .X(_02485_));
 sg13g2_mux2_1 _26152_ (.A0(\exec.memory_input[4] ),
    .A1(_10040_),
    .S(net783),
    .X(_02486_));
 sg13g2_mux2_1 _26153_ (.A0(\exec.memory_input[5] ),
    .A1(_10044_),
    .S(net783),
    .X(_02487_));
 sg13g2_mux2_1 _26154_ (.A0(\exec.memory_input[6] ),
    .A1(_10054_),
    .S(net783),
    .X(_02488_));
 sg13g2_nor2_1 _26155_ (.A(\exec.memory_input[7] ),
    .B(net783),
    .Y(_07449_));
 sg13g2_a21oi_1 _26156_ (.A1(net783),
    .A2(_10043_),
    .Y(_02489_),
    .B1(_07449_));
 sg13g2_and4_1 _26157_ (.A(_07162_),
    .B(_07198_),
    .C(_07222_),
    .D(_07447_),
    .X(_07450_));
 sg13g2_a21oi_1 _26158_ (.A1(_07395_),
    .A2(_07415_),
    .Y(_07451_),
    .B1(_07339_));
 sg13g2_and4_1 _26159_ (.A(_07269_),
    .B(_07312_),
    .C(_07450_),
    .D(_07451_),
    .X(_07452_));
 sg13g2_buf_8 _26160_ (.A(_07452_),
    .X(_07453_));
 sg13g2_a22oi_1 _26161_ (.Y(_07454_),
    .B1(_07375_),
    .B2(_07384_),
    .A2(_07362_),
    .A1(_07353_));
 sg13g2_buf_1 _26162_ (.A(_07454_),
    .X(_07455_));
 sg13g2_nand2b_1 _26163_ (.Y(_07456_),
    .B(net1305),
    .A_N(\exec.opcode[0] ));
 sg13g2_and2_1 _26164_ (.A(_09883_),
    .B(_07456_),
    .X(_07457_));
 sg13g2_nor3_1 _26165_ (.A(net1278),
    .B(net1307),
    .C(_09870_),
    .Y(_07458_));
 sg13g2_nand2b_1 _26166_ (.Y(_07459_),
    .B(net1227),
    .A_N(net1277));
 sg13g2_nand3b_1 _26167_ (.B(net1277),
    .C(_09878_),
    .Y(_07460_),
    .A_N(net1227));
 sg13g2_o21ai_1 _26168_ (.B1(_07460_),
    .Y(_07461_),
    .A1(net1306),
    .A2(_07459_));
 sg13g2_nor3_1 _26169_ (.A(_09913_),
    .B(_09870_),
    .C(_09873_),
    .Y(_07462_));
 sg13g2_nand2_1 _26170_ (.Y(_07463_),
    .A(_09880_),
    .B(_09881_));
 sg13g2_xnor2_1 _26171_ (.Y(_07464_),
    .A(_09876_),
    .B(net1308));
 sg13g2_nor4_1 _26172_ (.A(_07463_),
    .B(_09918_),
    .C(_07456_),
    .D(_07464_),
    .Y(_07465_));
 sg13g2_buf_2 _26173_ (.A(_07465_),
    .X(_07466_));
 sg13g2_a221oi_1 _26174_ (.B2(_07462_),
    .C1(_07466_),
    .B1(_07461_),
    .A1(_07457_),
    .Y(_07467_),
    .A2(_07458_));
 sg13g2_buf_2 _26175_ (.A(_07467_),
    .X(_07468_));
 sg13g2_inv_1 _26176_ (.Y(_07469_),
    .A(_07468_));
 sg13g2_or4_1 _26177_ (.A(_09876_),
    .B(net1306),
    .C(_09880_),
    .D(_09881_),
    .X(_07470_));
 sg13g2_or4_1 _26178_ (.A(net1305),
    .B(_09869_),
    .C(_09918_),
    .D(_07470_),
    .X(_07471_));
 sg13g2_buf_1 _26179_ (.A(_07471_),
    .X(_07472_));
 sg13g2_nand3_1 _26180_ (.B(_07472_),
    .C(_07468_),
    .A(net559),
    .Y(_07473_));
 sg13g2_buf_1 _26181_ (.A(_07473_),
    .X(_07474_));
 sg13g2_buf_2 _26182_ (.A(\exec.sp[4] ),
    .X(_07475_));
 sg13g2_inv_2 _26183_ (.Y(_07476_),
    .A(_07475_));
 sg13g2_nor4_1 _26184_ (.A(net1307),
    .B(net1309),
    .C(_07463_),
    .D(_09901_),
    .Y(_07477_));
 sg13g2_buf_2 _26185_ (.A(_07477_),
    .X(_07478_));
 sg13g2_or2_1 _26186_ (.X(_07479_),
    .B(_09881_),
    .A(_09880_));
 sg13g2_nor4_1 _26187_ (.A(net1306),
    .B(_09901_),
    .C(_09918_),
    .D(_07479_),
    .Y(_07480_));
 sg13g2_o21ai_1 _26188_ (.B1(net1278),
    .Y(_07481_),
    .A1(_07478_),
    .A2(_07480_));
 sg13g2_inv_1 _26189_ (.Y(_07482_),
    .A(_09878_));
 sg13g2_nand2_1 _26190_ (.Y(_07483_),
    .A(_07482_),
    .B(_07478_));
 sg13g2_nor4_1 _26191_ (.A(_09912_),
    .B(_09898_),
    .C(_09899_),
    .D(_09901_),
    .Y(_07484_));
 sg13g2_nor4_1 _26192_ (.A(net1306),
    .B(net1227),
    .C(_09901_),
    .D(_09918_),
    .Y(_07485_));
 sg13g2_o21ai_1 _26193_ (.B1(net1277),
    .Y(_07486_),
    .A1(_07484_),
    .A2(_07485_));
 sg13g2_inv_1 _26194_ (.Y(_07487_),
    .A(_09654_));
 sg13g2_nor2_2 _26195_ (.A(_07487_),
    .B(_07297_),
    .Y(_07488_));
 sg13g2_nand4_1 _26196_ (.B(_07483_),
    .C(_07486_),
    .A(_07481_),
    .Y(_07489_),
    .D(_07488_));
 sg13g2_xnor2_1 _26197_ (.Y(_07490_),
    .A(_07476_),
    .B(_07489_));
 sg13g2_nor2_1 _26198_ (.A(_07474_),
    .B(_07490_),
    .Y(_07491_));
 sg13g2_nor3_1 _26199_ (.A(_07455_),
    .B(_07469_),
    .C(_07491_),
    .Y(_07492_));
 sg13g2_nand2_1 _26200_ (.Y(_07493_),
    .A(_07472_),
    .B(_07468_));
 sg13g2_a21oi_1 _26201_ (.A1(_09730_),
    .A2(_07493_),
    .Y(_07494_),
    .B1(_07491_));
 sg13g2_a21o_1 _26202_ (.A2(_07492_),
    .A1(net406),
    .B1(_07494_),
    .X(_07495_));
 sg13g2_buf_1 _26203_ (.A(_07495_),
    .X(_07496_));
 sg13g2_buf_8 _26204_ (.A(_07455_),
    .X(_07497_));
 sg13g2_buf_1 _26205_ (.A(_07472_),
    .X(_07498_));
 sg13g2_nor3_1 _26206_ (.A(net535),
    .B(net454),
    .C(_07498_),
    .Y(_07499_));
 sg13g2_nor2_1 _26207_ (.A(net559),
    .B(net535),
    .Y(_07500_));
 sg13g2_a21oi_2 _26208_ (.B1(_07500_),
    .Y(_07501_),
    .A2(_07499_),
    .A1(net406));
 sg13g2_nand2_1 _26209_ (.Y(_07502_),
    .A(_07496_),
    .B(_07501_));
 sg13g2_buf_8 _26210_ (.A(_07502_),
    .X(_07503_));
 sg13g2_nand3_1 _26211_ (.B(_07483_),
    .C(_07486_),
    .A(_07481_),
    .Y(_07504_));
 sg13g2_buf_8 _26212_ (.A(_07504_),
    .X(_07505_));
 sg13g2_nand2_1 _26213_ (.Y(_07506_),
    .A(_07166_),
    .B(_07468_));
 sg13g2_buf_1 _26214_ (.A(net564),
    .X(_07507_));
 sg13g2_nand2_1 _26215_ (.Y(_07508_),
    .A(net525),
    .B(_07469_));
 sg13g2_o21ai_1 _26216_ (.B1(_07508_),
    .Y(_07509_),
    .A1(_07505_),
    .A2(_07506_));
 sg13g2_mux2_1 _26217_ (.A0(_07468_),
    .A1(_07474_),
    .S(net530),
    .X(_07510_));
 sg13g2_a21oi_1 _26218_ (.A1(net559),
    .A2(_07472_),
    .Y(_07511_),
    .B1(_07507_));
 sg13g2_a21oi_1 _26219_ (.A1(net525),
    .A2(_07505_),
    .Y(_07512_),
    .B1(_07511_));
 sg13g2_o21ai_1 _26220_ (.B1(_07512_),
    .Y(_07513_),
    .A1(net531),
    .A2(_07510_));
 sg13g2_a21oi_1 _26221_ (.A1(net531),
    .A2(_07509_),
    .Y(_07514_),
    .B1(_07513_));
 sg13g2_nand3_1 _26222_ (.B(_07514_),
    .C(_07453_),
    .A(_07387_),
    .Y(_07515_));
 sg13g2_buf_1 _26223_ (.A(_07515_),
    .X(_07516_));
 sg13g2_nand4_1 _26224_ (.B(_07312_),
    .C(_07450_),
    .A(_07269_),
    .Y(_07517_),
    .D(_07451_));
 sg13g2_buf_2 _26225_ (.A(_07517_),
    .X(_07518_));
 sg13g2_nor3_1 _26226_ (.A(net525),
    .B(_07505_),
    .C(_07493_),
    .Y(_07519_));
 sg13g2_a21o_1 _26227_ (.A2(_07493_),
    .A1(net525),
    .B1(_07519_),
    .X(_07520_));
 sg13g2_nand2_1 _26228_ (.Y(_07521_),
    .A(net530),
    .B(net559));
 sg13g2_mux2_1 _26229_ (.A0(_07521_),
    .A1(net525),
    .S(_07493_),
    .X(_07522_));
 sg13g2_nor2_1 _26230_ (.A(net525),
    .B(net559),
    .Y(_07523_));
 sg13g2_a21oi_1 _26231_ (.A1(net525),
    .A2(_07505_),
    .Y(_07524_),
    .B1(_07523_));
 sg13g2_o21ai_1 _26232_ (.B1(_07524_),
    .Y(_07525_),
    .A1(net531),
    .A2(_07522_));
 sg13g2_a21oi_1 _26233_ (.A1(net531),
    .A2(_07520_),
    .Y(_07526_),
    .B1(_07525_));
 sg13g2_o21ai_1 _26234_ (.B1(_07526_),
    .Y(_07527_),
    .A1(net454),
    .A2(_07518_));
 sg13g2_buf_1 _26235_ (.A(_07527_),
    .X(_07528_));
 sg13g2_nand2_1 _26236_ (.Y(_07529_),
    .A(_07516_),
    .B(_07528_));
 sg13g2_buf_1 _26237_ (.A(_07529_),
    .X(_07530_));
 sg13g2_nand2b_1 _26238_ (.Y(_07531_),
    .B(net140),
    .A_N(_07503_));
 sg13g2_buf_1 _26239_ (.A(_00067_),
    .X(_07532_));
 sg13g2_xnor2_1 _26240_ (.Y(_07533_),
    .A(_07532_),
    .B(_07114_));
 sg13g2_nor2_1 _26241_ (.A(_07505_),
    .B(_07474_),
    .Y(_07534_));
 sg13g2_nand2_1 _26242_ (.Y(_07535_),
    .A(_07533_),
    .B(_07534_));
 sg13g2_o21ai_1 _26243_ (.B1(net559),
    .Y(_07536_),
    .A1(net531),
    .A2(_07468_));
 sg13g2_nand2_1 _26244_ (.Y(_07537_),
    .A(net795),
    .B(_07536_));
 sg13g2_nand2_1 _26245_ (.Y(_07538_),
    .A(net525),
    .B(_10002_));
 sg13g2_o21ai_1 _26246_ (.B1(_07538_),
    .Y(_07539_),
    .A1(_09732_),
    .A2(_07468_));
 sg13g2_o21ai_1 _26247_ (.B1(net868),
    .Y(_07540_),
    .A1(_07505_),
    .A2(_07539_));
 sg13g2_nand3_1 _26248_ (.B(_07537_),
    .C(_07540_),
    .A(_07535_),
    .Y(_07541_));
 sg13g2_buf_1 _26249_ (.A(net534),
    .X(_07542_));
 sg13g2_a221oi_1 _26250_ (.B2(_07453_),
    .C1(net524),
    .B1(_07387_),
    .A1(_09669_),
    .Y(_07543_),
    .A2(_09642_));
 sg13g2_nor4_2 _26251_ (.A(_07212_),
    .B(net454),
    .C(_07498_),
    .Y(_07544_),
    .D(_07518_));
 sg13g2_nor3_2 _26252_ (.A(_07541_),
    .B(_07543_),
    .C(_07544_),
    .Y(_07545_));
 sg13g2_buf_8 _26253_ (.A(_07545_),
    .X(_07546_));
 sg13g2_buf_8 _26254_ (.A(net143),
    .X(_07547_));
 sg13g2_xnor2_1 _26255_ (.Y(_07548_),
    .A(_07487_),
    .B(_07297_));
 sg13g2_a21oi_1 _26256_ (.A1(_09654_),
    .A2(_07505_),
    .Y(_07549_),
    .B1(_07534_));
 sg13g2_a22oi_1 _26257_ (.Y(_07550_),
    .B1(_07469_),
    .B2(_09710_),
    .A2(_07124_),
    .A1(_10002_));
 sg13g2_a22oi_1 _26258_ (.Y(_07551_),
    .B1(_07549_),
    .B2(_07550_),
    .A2(_07548_),
    .A1(_07534_));
 sg13g2_nor4_1 _26259_ (.A(_09893_),
    .B(net1308),
    .C(_09918_),
    .D(_07470_),
    .Y(_07552_));
 sg13g2_buf_1 _26260_ (.A(_07552_),
    .X(_07553_));
 sg13g2_nand2_1 _26261_ (.Y(_07554_),
    .A(_09710_),
    .B(_07553_));
 sg13g2_a21oi_1 _26262_ (.A1(_07387_),
    .A2(net406),
    .Y(_07555_),
    .B1(_07554_));
 sg13g2_nor4_1 _26263_ (.A(net536),
    .B(_07497_),
    .C(_07542_),
    .D(_07518_),
    .Y(_07556_));
 sg13g2_nor3_1 _26264_ (.A(_07551_),
    .B(_07555_),
    .C(_07556_),
    .Y(_07557_));
 sg13g2_buf_1 _26265_ (.A(_07557_),
    .X(_07558_));
 sg13g2_buf_8 _26266_ (.A(net142),
    .X(_07559_));
 sg13g2_buf_1 _26267_ (.A(_00065_),
    .X(_07560_));
 sg13g2_buf_1 _26268_ (.A(_07553_),
    .X(_07561_));
 sg13g2_o21ai_1 _26269_ (.B1(_07561_),
    .Y(_07562_),
    .A1(_07560_),
    .A2(_07387_));
 sg13g2_nor2_1 _26270_ (.A(_09877_),
    .B(_07482_),
    .Y(_07563_));
 sg13g2_nand2_1 _26271_ (.Y(_07564_),
    .A(_07478_),
    .B(_07563_));
 sg13g2_and4_1 _26272_ (.A(_10152_),
    .B(_09897_),
    .C(net534),
    .D(_07564_),
    .X(_07565_));
 sg13g2_and4_1 _26273_ (.A(net1277),
    .B(_09912_),
    .C(_09879_),
    .D(_09919_),
    .X(_07566_));
 sg13g2_buf_1 _26274_ (.A(_07566_),
    .X(_07567_));
 sg13g2_buf_1 _26275_ (.A(_07567_),
    .X(_07568_));
 sg13g2_a21oi_1 _26276_ (.A1(_07486_),
    .A2(_07565_),
    .Y(_07569_),
    .B1(net523));
 sg13g2_inv_1 _26277_ (.Y(_07570_),
    .A(_07569_));
 sg13g2_nand2_1 _26278_ (.Y(_07571_),
    .A(_07560_),
    .B(net534));
 sg13g2_nor2_1 _26279_ (.A(_10002_),
    .B(_07505_),
    .Y(_07572_));
 sg13g2_mux2_1 _26280_ (.A0(_09723_),
    .A1(_07571_),
    .S(_07572_),
    .X(_07573_));
 sg13g2_buf_2 _26281_ (.A(_07573_),
    .X(_07574_));
 sg13g2_inv_1 _26282_ (.Y(_07575_),
    .A(_07574_));
 sg13g2_o21ai_1 _26283_ (.B1(_07575_),
    .Y(_07576_),
    .A1(net533),
    .A2(_07570_));
 sg13g2_inv_1 _26284_ (.Y(_07577_),
    .A(_07560_));
 sg13g2_o21ai_1 _26285_ (.B1(_07570_),
    .Y(_07578_),
    .A1(_07577_),
    .A2(_07575_));
 sg13g2_nor2_2 _26286_ (.A(_07497_),
    .B(_07518_),
    .Y(_07579_));
 sg13g2_nand2_1 _26287_ (.Y(_07580_),
    .A(_07577_),
    .B(_07574_));
 sg13g2_nor2_1 _26288_ (.A(_10143_),
    .B(_00068_),
    .Y(_07581_));
 sg13g2_o21ai_1 _26289_ (.B1(_07581_),
    .Y(_07582_),
    .A1(net406),
    .A2(_07580_));
 sg13g2_a221oi_1 _26290_ (.B2(_07579_),
    .C1(_07582_),
    .B1(_07578_),
    .A1(_07562_),
    .Y(_07583_),
    .A2(_07576_));
 sg13g2_buf_1 _26291_ (.A(_07583_),
    .X(_07584_));
 sg13g2_buf_1 _26292_ (.A(_07584_),
    .X(_07585_));
 sg13g2_nand3_1 _26293_ (.B(net138),
    .C(net137),
    .A(net139),
    .Y(_07586_));
 sg13g2_buf_1 _26294_ (.A(_07586_),
    .X(_07587_));
 sg13g2_nor2_1 _26295_ (.A(_07531_),
    .B(_07587_),
    .Y(_07588_));
 sg13g2_buf_2 _26296_ (.A(_07588_),
    .X(_07589_));
 sg13g2_buf_1 _26297_ (.A(_07589_),
    .X(_07590_));
 sg13g2_buf_1 _26298_ (.A(net1302),
    .X(_07591_));
 sg13g2_nor2_1 _26299_ (.A(net868),
    .B(_09654_),
    .Y(_07592_));
 sg13g2_nand2_1 _26300_ (.Y(_07593_),
    .A(_07476_),
    .B(_07592_));
 sg13g2_buf_1 _26301_ (.A(_07593_),
    .X(_07594_));
 sg13g2_and2_1 _26302_ (.A(_09924_),
    .B(net3),
    .X(_07595_));
 sg13g2_buf_1 _26303_ (.A(_07595_),
    .X(_07596_));
 sg13g2_and3_1 _26304_ (.X(_07597_),
    .A(_09906_),
    .B(_09922_),
    .C(_07596_));
 sg13g2_buf_1 _26305_ (.A(_07597_),
    .X(_07598_));
 sg13g2_nand2_1 _26306_ (.Y(_07599_),
    .A(_09732_),
    .B(_07598_));
 sg13g2_buf_2 _26307_ (.A(_07599_),
    .X(_07600_));
 sg13g2_nor2_1 _26308_ (.A(_07594_),
    .B(_07600_),
    .Y(_07601_));
 sg13g2_buf_1 _26309_ (.A(_07601_),
    .X(_07602_));
 sg13g2_nand4_1 _26310_ (.B(_07528_),
    .C(_07496_),
    .A(_07516_),
    .Y(_07603_),
    .D(_07501_));
 sg13g2_buf_2 _26311_ (.A(_07603_),
    .X(_07604_));
 sg13g2_or3_1 _26312_ (.A(_07541_),
    .B(_07543_),
    .C(_07544_),
    .X(_07605_));
 sg13g2_buf_1 _26313_ (.A(_07605_),
    .X(_07606_));
 sg13g2_buf_8 _26314_ (.A(_07606_),
    .X(_07607_));
 sg13g2_or3_1 _26315_ (.A(_07551_),
    .B(_07555_),
    .C(_07556_),
    .X(_07608_));
 sg13g2_buf_2 _26316_ (.A(_07608_),
    .X(_07609_));
 sg13g2_buf_8 _26317_ (.A(_07609_),
    .X(_07610_));
 sg13g2_nand3_1 _26318_ (.B(_07581_),
    .C(_07568_),
    .A(_07574_),
    .Y(_07611_));
 sg13g2_buf_1 _26319_ (.A(_07611_),
    .X(_07612_));
 sg13g2_or4_1 _26320_ (.A(_07604_),
    .B(_07607_),
    .C(net135),
    .D(_07612_),
    .X(_07613_));
 sg13g2_buf_1 _26321_ (.A(_07613_),
    .X(_07614_));
 sg13g2_nor2_1 _26322_ (.A(net1270),
    .B(net509),
    .Y(_07615_));
 sg13g2_and2_1 _26323_ (.A(_07614_),
    .B(_07615_),
    .X(_07616_));
 sg13g2_buf_2 _26324_ (.A(_07616_),
    .X(_07617_));
 sg13g2_a22oi_1 _26325_ (.Y(_07618_),
    .B1(_07617_),
    .B2(\stack[0][0] ),
    .A2(net509),
    .A1(net1226));
 sg13g2_buf_1 _26326_ (.A(net495),
    .X(_07619_));
 sg13g2_buf_1 _26327_ (.A(net480),
    .X(_07620_));
 sg13g2_nor2_2 _26328_ (.A(net140),
    .B(_07503_),
    .Y(_07621_));
 sg13g2_nor3_1 _26329_ (.A(net136),
    .B(net135),
    .C(_07612_),
    .Y(_07622_));
 sg13g2_and2_1 _26330_ (.A(_07621_),
    .B(_07622_),
    .X(_07623_));
 sg13g2_buf_1 _26331_ (.A(_07623_),
    .X(_07624_));
 sg13g2_nand2_1 _26332_ (.Y(_07625_),
    .A(_07481_),
    .B(_07483_));
 sg13g2_xor2_1 _26333_ (.B(_07101_),
    .A(_09877_),
    .X(_07626_));
 sg13g2_nand4_1 _26334_ (.B(net1277),
    .C(_09875_),
    .A(net1275),
    .Y(_07627_),
    .D(_07626_));
 sg13g2_nand2_1 _26335_ (.Y(_07628_),
    .A(net534),
    .B(_07627_));
 sg13g2_buf_1 _26336_ (.A(_07628_),
    .X(_07629_));
 sg13g2_nor3_1 _26337_ (.A(net1307),
    .B(net1309),
    .C(_09901_),
    .Y(_07630_));
 sg13g2_nand4_1 _26338_ (.B(_09912_),
    .C(_09916_),
    .A(_09890_),
    .Y(_07631_),
    .D(_07630_));
 sg13g2_buf_1 _26339_ (.A(_07631_),
    .X(_07632_));
 sg13g2_nand4_1 _26340_ (.B(net1227),
    .C(_09875_),
    .A(_09890_),
    .Y(_07633_),
    .D(_09916_));
 sg13g2_buf_1 _26341_ (.A(_07633_),
    .X(_07634_));
 sg13g2_nand2_1 _26342_ (.Y(_07635_),
    .A(_07632_),
    .B(_07634_));
 sg13g2_or2_1 _26343_ (.X(_07636_),
    .B(_07567_),
    .A(_07466_));
 sg13g2_buf_1 _26344_ (.A(_07636_),
    .X(_07637_));
 sg13g2_nor4_1 _26345_ (.A(_07625_),
    .B(net518),
    .C(_07635_),
    .D(_07637_),
    .Y(_07638_));
 sg13g2_buf_1 _26346_ (.A(_07638_),
    .X(_07639_));
 sg13g2_buf_1 _26347_ (.A(_07639_),
    .X(_07640_));
 sg13g2_nor2_1 _26348_ (.A(net1308),
    .B(_09918_),
    .Y(_07641_));
 sg13g2_and4_1 _26349_ (.A(net1305),
    .B(_09883_),
    .C(_09916_),
    .D(_07641_),
    .X(_07642_));
 sg13g2_buf_1 _26350_ (.A(_07642_),
    .X(_07643_));
 sg13g2_nand2_1 _26351_ (.Y(_07644_),
    .A(_09885_),
    .B(_09919_));
 sg13g2_nand2_1 _26352_ (.Y(_07645_),
    .A(_07632_),
    .B(_07644_));
 sg13g2_a21oi_1 _26353_ (.A1(net481),
    .A2(_07643_),
    .Y(_07646_),
    .B1(_07645_));
 sg13g2_and2_1 _26354_ (.A(_09916_),
    .B(_07478_),
    .X(_07647_));
 sg13g2_buf_2 _26355_ (.A(_07647_),
    .X(_07648_));
 sg13g2_a21oi_1 _26356_ (.A1(net1275),
    .A2(_07478_),
    .Y(_07649_),
    .B1(_07480_));
 sg13g2_nor2_1 _26357_ (.A(_09913_),
    .B(_07649_),
    .Y(_07650_));
 sg13g2_buf_2 _26358_ (.A(_07650_),
    .X(_07651_));
 sg13g2_a221oi_1 _26359_ (.B2(\exec.memory_input[0] ),
    .C1(_07639_),
    .B1(_07651_),
    .A1(net486),
    .Y(_07652_),
    .A2(_07648_));
 sg13g2_o21ai_1 _26360_ (.B1(_07652_),
    .Y(_07653_),
    .A1(_09772_),
    .A2(_07646_));
 sg13g2_inv_1 _26361_ (.Y(_07654_),
    .A(_07653_));
 sg13g2_and4_1 _26362_ (.A(net1275),
    .B(_09889_),
    .C(_09875_),
    .D(_07626_),
    .X(_07655_));
 sg13g2_buf_1 _26363_ (.A(_07655_),
    .X(_07656_));
 sg13g2_a21oi_1 _26364_ (.A1(net495),
    .A2(_07656_),
    .Y(_07657_),
    .B1(net533));
 sg13g2_nor3_1 _26365_ (.A(net495),
    .B(_07466_),
    .C(_07656_),
    .Y(_07658_));
 sg13g2_a21oi_1 _26366_ (.A1(net495),
    .A2(_07634_),
    .Y(_07659_),
    .B1(_07658_));
 sg13g2_nor3_1 _26367_ (.A(net481),
    .B(net523),
    .C(_07659_),
    .Y(_07660_));
 sg13g2_a21o_1 _26368_ (.A2(_07657_),
    .A1(net481),
    .B1(_07660_),
    .X(_07661_));
 sg13g2_a22oi_1 _26369_ (.Y(_07662_),
    .B1(_07654_),
    .B2(_07661_),
    .A2(net479),
    .A1(_07482_));
 sg13g2_buf_1 _26370_ (.A(_07662_),
    .X(_07663_));
 sg13g2_buf_1 _26371_ (.A(_07663_),
    .X(_07664_));
 sg13g2_buf_1 _26372_ (.A(_07664_),
    .X(_07665_));
 sg13g2_a22oi_1 _26373_ (.Y(_07666_),
    .B1(_07589_),
    .B2(net131),
    .A2(_07624_),
    .A1(net453));
 sg13g2_o21ai_1 _26374_ (.B1(_07666_),
    .Y(_02523_),
    .A1(net65),
    .A2(_07618_));
 sg13g2_buf_1 _26375_ (.A(net1299),
    .X(_07667_));
 sg13g2_buf_1 _26376_ (.A(net1225),
    .X(_07668_));
 sg13g2_a22oi_1 _26377_ (.Y(_07669_),
    .B1(_07617_),
    .B2(\stack[0][1] ),
    .A2(net509),
    .A1(net883));
 sg13g2_nand3_1 _26378_ (.B(_09883_),
    .C(_07563_),
    .A(_09875_),
    .Y(_07670_));
 sg13g2_buf_1 _26379_ (.A(_07670_),
    .X(_07671_));
 sg13g2_xnor2_1 _26380_ (.Y(_07672_),
    .A(net481),
    .B(_07671_));
 sg13g2_a21oi_1 _26381_ (.A1(_09772_),
    .A2(net524),
    .Y(_07673_),
    .B1(_07672_));
 sg13g2_and3_1 _26382_ (.X(_07674_),
    .A(_09875_),
    .B(_09883_),
    .C(_07563_));
 sg13g2_buf_1 _26383_ (.A(_07674_),
    .X(_07675_));
 sg13g2_nor2_2 _26384_ (.A(_07553_),
    .B(_07675_),
    .Y(_07676_));
 sg13g2_buf_1 _26385_ (.A(_07675_),
    .X(_07677_));
 sg13g2_mux2_1 _26386_ (.A0(_07676_),
    .A1(net517),
    .S(net481),
    .X(_07678_));
 sg13g2_a221oi_1 _26387_ (.B2(net495),
    .C1(net486),
    .B1(_07678_),
    .A1(_07163_),
    .Y(_07679_),
    .A2(_07561_));
 sg13g2_a21oi_1 _26388_ (.A1(_10096_),
    .A2(_07673_),
    .Y(_07680_),
    .B1(_07679_));
 sg13g2_xor2_1 _26389_ (.B(_07680_),
    .A(_07224_),
    .X(_07681_));
 sg13g2_or4_1 _26390_ (.A(_07463_),
    .B(_09918_),
    .C(_07456_),
    .D(_07464_),
    .X(_07682_));
 sg13g2_buf_1 _26391_ (.A(_07682_),
    .X(_07683_));
 sg13g2_and4_1 _26392_ (.A(_09890_),
    .B(net1227),
    .C(_09875_),
    .D(_09916_),
    .X(_07684_));
 sg13g2_buf_1 _26393_ (.A(_07684_),
    .X(_07685_));
 sg13g2_nand2_1 _26394_ (.Y(_07686_),
    .A(net486),
    .B(_07685_));
 sg13g2_o21ai_1 _26395_ (.B1(_07686_),
    .Y(_07687_),
    .A1(net486),
    .A2(_07683_));
 sg13g2_o21ai_1 _26396_ (.B1(_07224_),
    .Y(_07688_),
    .A1(net523),
    .A2(_07687_));
 sg13g2_nand4_1 _26397_ (.B(_09883_),
    .C(_09916_),
    .A(net1305),
    .Y(_07689_),
    .D(_07641_));
 sg13g2_buf_1 _26398_ (.A(_07689_),
    .X(_07690_));
 sg13g2_nor2_1 _26399_ (.A(_07224_),
    .B(_07690_),
    .Y(_07691_));
 sg13g2_o21ai_1 _26400_ (.B1(net486),
    .Y(_07692_),
    .A1(_07645_),
    .A2(_07691_));
 sg13g2_nand2_1 _26401_ (.Y(_07693_),
    .A(net485),
    .B(_07648_));
 sg13g2_and2_1 _26402_ (.A(_09885_),
    .B(_07630_),
    .X(_07694_));
 sg13g2_buf_2 _26403_ (.A(_07694_),
    .X(_07695_));
 sg13g2_a221oi_1 _26404_ (.B2(net495),
    .C1(_07639_),
    .B1(_07695_),
    .A1(\exec.memory_input[1] ),
    .Y(_07696_),
    .A2(_07651_));
 sg13g2_nand4_1 _26405_ (.B(_07692_),
    .C(_07693_),
    .A(_07688_),
    .Y(_07697_),
    .D(_07696_));
 sg13g2_a21oi_1 _26406_ (.A1(net518),
    .A2(_07681_),
    .Y(_07698_),
    .B1(_07697_));
 sg13g2_a21oi_1 _26407_ (.A1(_09913_),
    .A2(_07640_),
    .Y(_07699_),
    .B1(_07698_));
 sg13g2_buf_1 _26408_ (.A(_07699_),
    .X(_07700_));
 sg13g2_buf_1 _26409_ (.A(_07700_),
    .X(_07701_));
 sg13g2_buf_1 _26410_ (.A(net119),
    .X(_07702_));
 sg13g2_a22oi_1 _26411_ (.Y(_07703_),
    .B1(_07589_),
    .B2(net105),
    .A2(_07624_),
    .A1(net447));
 sg13g2_o21ai_1 _26412_ (.B1(_07703_),
    .Y(_02524_),
    .A1(net65),
    .A2(_07669_));
 sg13g2_buf_1 _26413_ (.A(net1301),
    .X(_07704_));
 sg13g2_buf_1 _26414_ (.A(net1224),
    .X(_07705_));
 sg13g2_a22oi_1 _26415_ (.Y(_07706_),
    .B1(_07617_),
    .B2(\stack[0][2] ),
    .A2(net509),
    .A1(net882));
 sg13g2_buf_1 _26416_ (.A(net485),
    .X(_07707_));
 sg13g2_nand2_1 _26417_ (.Y(_07708_),
    .A(_10182_),
    .B(_07644_));
 sg13g2_o21ai_1 _26418_ (.B1(_07466_),
    .Y(_07709_),
    .A1(_07269_),
    .A2(_07708_));
 sg13g2_nand2_1 _26419_ (.Y(_07710_),
    .A(_07632_),
    .B(_07709_));
 sg13g2_o21ai_1 _26420_ (.B1(_09807_),
    .Y(_07711_),
    .A1(_07269_),
    .A2(_07683_));
 sg13g2_a21oi_1 _26421_ (.A1(net485),
    .A2(_07685_),
    .Y(_07712_),
    .B1(net523));
 sg13g2_a221oi_1 _26422_ (.B2(\exec.memory_input[2] ),
    .C1(net479),
    .B1(_07651_),
    .A1(_10176_),
    .Y(_07713_),
    .A2(_07648_));
 sg13g2_o21ai_1 _26423_ (.B1(_07713_),
    .Y(_07714_),
    .A1(_07269_),
    .A2(_07712_));
 sg13g2_a221oi_1 _26424_ (.B2(_07711_),
    .C1(_07714_),
    .B1(_07710_),
    .A1(net473),
    .Y(_07715_),
    .A2(_07695_));
 sg13g2_and4_1 _26425_ (.A(_09668_),
    .B(_09700_),
    .C(_09706_),
    .D(_07676_),
    .X(_07716_));
 sg13g2_a221oi_1 _26426_ (.B2(net486),
    .C1(_07716_),
    .B1(_07677_),
    .A1(_07198_),
    .Y(_07717_),
    .A2(_07222_));
 sg13g2_nor2_1 _26427_ (.A(net481),
    .B(_07716_),
    .Y(_07718_));
 sg13g2_a21oi_1 _26428_ (.A1(_07198_),
    .A2(_07222_),
    .Y(_07719_),
    .B1(net481));
 sg13g2_nor4_2 _26429_ (.A(_09771_),
    .B(_07717_),
    .C(_07718_),
    .Y(_07720_),
    .D(_07719_));
 sg13g2_nand2_1 _26430_ (.Y(_07721_),
    .A(net563),
    .B(_07472_));
 sg13g2_a221oi_1 _26431_ (.B2(_09768_),
    .C1(_07721_),
    .B1(_09764_),
    .A1(_09755_),
    .Y(_07722_),
    .A2(_09759_));
 sg13g2_nand2_1 _26432_ (.Y(_07723_),
    .A(_09710_),
    .B(_07472_));
 sg13g2_a221oi_1 _26433_ (.B2(_09749_),
    .C1(_07723_),
    .B1(_09739_),
    .A1(_09722_),
    .Y(_07724_),
    .A2(_09731_));
 sg13g2_or3_1 _26434_ (.A(_07677_),
    .B(_07722_),
    .C(_07724_),
    .X(_07725_));
 sg13g2_a22oi_1 _26435_ (.Y(_07726_),
    .B1(_07725_),
    .B2(net486),
    .A2(_07553_),
    .A1(net481));
 sg13g2_nor2_1 _26436_ (.A(_07224_),
    .B(_07726_),
    .Y(_07727_));
 sg13g2_nor2_1 _26437_ (.A(_07720_),
    .B(_07727_),
    .Y(_07728_));
 sg13g2_nand2_1 _26438_ (.Y(_07729_),
    .A(_10182_),
    .B(net517));
 sg13g2_nand4_1 _26439_ (.B(_09771_),
    .C(_10182_),
    .A(_09708_),
    .Y(_07730_),
    .D(net534));
 sg13g2_and2_1 _26440_ (.A(_09807_),
    .B(_07676_),
    .X(_07731_));
 sg13g2_o21ai_1 _26441_ (.B1(_07731_),
    .Y(_07732_),
    .A1(_10096_),
    .A2(_10164_));
 sg13g2_nand3_1 _26442_ (.B(_07730_),
    .C(_07732_),
    .A(_07729_),
    .Y(_07733_));
 sg13g2_xnor2_1 _26443_ (.Y(_07734_),
    .A(_07269_),
    .B(_07733_));
 sg13g2_xnor2_1 _26444_ (.Y(_07735_),
    .A(_07728_),
    .B(_07734_));
 sg13g2_nand2_1 _26445_ (.Y(_07736_),
    .A(net518),
    .B(_07735_));
 sg13g2_a22oi_1 _26446_ (.Y(_07737_),
    .B1(_07715_),
    .B2(_07736_),
    .A2(_07640_),
    .A1(_09912_));
 sg13g2_buf_2 _26447_ (.A(_07737_),
    .X(_07738_));
 sg13g2_buf_1 _26448_ (.A(_07738_),
    .X(_07739_));
 sg13g2_buf_2 _26449_ (.A(net118),
    .X(_07740_));
 sg13g2_a22oi_1 _26450_ (.Y(_07741_),
    .B1(_07589_),
    .B2(net104),
    .A2(_07624_),
    .A1(net452));
 sg13g2_o21ai_1 _26451_ (.B1(_07741_),
    .Y(_02525_),
    .A1(net65),
    .A2(_07706_));
 sg13g2_buf_1 _26452_ (.A(net1300),
    .X(_07742_));
 sg13g2_buf_1 _26453_ (.A(net1223),
    .X(_07743_));
 sg13g2_a22oi_1 _26454_ (.Y(_07744_),
    .B1(_07617_),
    .B2(\stack[0][3] ),
    .A2(_07602_),
    .A1(net881));
 sg13g2_buf_1 _26455_ (.A(net510),
    .X(_07745_));
 sg13g2_buf_1 _26456_ (.A(_07604_),
    .X(_07746_));
 sg13g2_nand2_1 _26457_ (.Y(_07747_),
    .A(net143),
    .B(net142));
 sg13g2_buf_2 _26458_ (.A(_07747_),
    .X(_07748_));
 sg13g2_nand2_1 _26459_ (.Y(_07749_),
    .A(_07581_),
    .B(_07568_));
 sg13g2_buf_1 _26460_ (.A(_07749_),
    .X(_07750_));
 sg13g2_buf_1 _26461_ (.A(_07750_),
    .X(_07751_));
 sg13g2_xnor2_1 _26462_ (.Y(_07752_),
    .A(_07560_),
    .B(_07579_));
 sg13g2_o21ai_1 _26463_ (.B1(_07574_),
    .Y(_07753_),
    .A1(net524),
    .A2(_07752_));
 sg13g2_buf_2 _26464_ (.A(_07753_),
    .X(_07754_));
 sg13g2_buf_1 _26465_ (.A(_07754_),
    .X(_07755_));
 sg13g2_nor4_1 _26466_ (.A(net130),
    .B(_07748_),
    .C(net491),
    .D(net129),
    .Y(_07756_));
 sg13g2_nand2b_1 _26467_ (.Y(_07757_),
    .B(_07644_),
    .A_N(net455));
 sg13g2_o21ai_1 _26468_ (.B1(_07632_),
    .Y(_07758_),
    .A1(net455),
    .A2(_07634_));
 sg13g2_a21o_1 _26469_ (.A2(_07757_),
    .A1(_07466_),
    .B1(_07758_),
    .X(_07759_));
 sg13g2_a21oi_1 _26470_ (.A1(_09788_),
    .A2(_07466_),
    .Y(_07760_),
    .B1(net523));
 sg13g2_a21o_1 _26471_ (.A2(_07651_),
    .A1(\exec.memory_input[3] ),
    .B1(_07639_),
    .X(_07761_));
 sg13g2_a221oi_1 _26472_ (.B2(_10182_),
    .C1(_07761_),
    .B1(_07695_),
    .A1(_09864_),
    .Y(_07762_),
    .A2(_07648_));
 sg13g2_o21ai_1 _26473_ (.B1(_07762_),
    .Y(_07763_),
    .A1(net455),
    .A2(_07760_));
 sg13g2_a21oi_1 _26474_ (.A1(net510),
    .A2(_07759_),
    .Y(_07764_),
    .B1(_07763_));
 sg13g2_nor3_1 _26475_ (.A(_07720_),
    .B(_07727_),
    .C(_07733_),
    .Y(_07765_));
 sg13g2_and3_1 _26476_ (.X(_07766_),
    .A(_07240_),
    .B(_07256_),
    .C(_07267_));
 sg13g2_o21ai_1 _26477_ (.B1(_07766_),
    .Y(_07767_),
    .A1(_07224_),
    .A2(_07726_));
 sg13g2_nand4_1 _26478_ (.B(_07729_),
    .C(_07730_),
    .A(_07766_),
    .Y(_07768_),
    .D(_07732_));
 sg13g2_o21ai_1 _26479_ (.B1(_07768_),
    .Y(_07769_),
    .A1(_07720_),
    .A2(_07767_));
 sg13g2_or2_1 _26480_ (.X(_07770_),
    .B(_07769_),
    .A(_07765_));
 sg13g2_buf_1 _26481_ (.A(_07770_),
    .X(_07771_));
 sg13g2_inv_1 _26482_ (.Y(_07772_),
    .A(_07676_));
 sg13g2_nand4_1 _26483_ (.B(_09771_),
    .C(_09807_),
    .A(_09708_),
    .Y(_07773_),
    .D(net534));
 sg13g2_nor2_1 _26484_ (.A(_09788_),
    .B(net517),
    .Y(_07774_));
 sg13g2_a221oi_1 _26485_ (.B2(_07774_),
    .C1(_10189_),
    .B1(_07773_),
    .A1(_09788_),
    .Y(_07775_),
    .A2(_07772_));
 sg13g2_buf_2 _26486_ (.A(_07775_),
    .X(_07776_));
 sg13g2_xor2_1 _26487_ (.B(_07776_),
    .A(net455),
    .X(_07777_));
 sg13g2_xnor2_1 _26488_ (.Y(_07778_),
    .A(_07771_),
    .B(_07777_));
 sg13g2_nor2_1 _26489_ (.A(net533),
    .B(_07656_),
    .Y(_07779_));
 sg13g2_buf_1 _26490_ (.A(_07779_),
    .X(_07780_));
 sg13g2_and2_1 _26491_ (.A(_07780_),
    .B(_07764_),
    .X(_07781_));
 sg13g2_a221oi_1 _26492_ (.B2(_07778_),
    .C1(_07781_),
    .B1(_07764_),
    .A1(_09890_),
    .Y(_07782_),
    .A2(net479));
 sg13g2_buf_2 _26493_ (.A(_07782_),
    .X(_07783_));
 sg13g2_buf_1 _26494_ (.A(_07783_),
    .X(_07784_));
 sg13g2_buf_8 _26495_ (.A(_07784_),
    .X(_07785_));
 sg13g2_a22oi_1 _26496_ (.Y(_07786_),
    .B1(net91),
    .B2(_07590_),
    .A2(_07756_),
    .A1(net492));
 sg13g2_o21ai_1 _26497_ (.B1(_07786_),
    .Y(_02526_),
    .A1(_07590_),
    .A2(_07744_));
 sg13g2_buf_1 _26498_ (.A(_10022_),
    .X(_07787_));
 sg13g2_nand2_1 _26499_ (.Y(_07788_),
    .A(net1222),
    .B(net509));
 sg13g2_nand3_1 _26500_ (.B(_07621_),
    .C(_07622_),
    .A(_10190_),
    .Y(_07789_));
 sg13g2_nand2_1 _26501_ (.Y(_07790_),
    .A(\stack[0][4] ),
    .B(_07617_));
 sg13g2_nand3_1 _26502_ (.B(_07789_),
    .C(_07790_),
    .A(_07788_),
    .Y(_07791_));
 sg13g2_nand2_1 _26503_ (.Y(_07792_),
    .A(net496),
    .B(_07676_));
 sg13g2_nand2_1 _26504_ (.Y(_07793_),
    .A(_09864_),
    .B(net534));
 sg13g2_mux2_1 _26505_ (.A0(_07792_),
    .A1(_07793_),
    .S(_10189_),
    .X(_07794_));
 sg13g2_a21oi_1 _26506_ (.A1(_09864_),
    .A2(net517),
    .Y(_07795_),
    .B1(_07340_));
 sg13g2_nand2_1 _26507_ (.Y(_07796_),
    .A(_07794_),
    .B(_07795_));
 sg13g2_nand3_1 _26508_ (.B(net487),
    .C(_09809_),
    .A(_09708_),
    .Y(_07797_));
 sg13g2_or2_1 _26509_ (.X(_07798_),
    .B(_07793_),
    .A(_07339_));
 sg13g2_a21oi_1 _26510_ (.A1(_07797_),
    .A2(_07671_),
    .Y(_07799_),
    .B1(_07798_));
 sg13g2_nand2_1 _26511_ (.Y(_07800_),
    .A(_10117_),
    .B(net534));
 sg13g2_nor4_2 _26512_ (.A(_10189_),
    .B(_07339_),
    .C(net517),
    .Y(_07801_),
    .D(_07800_));
 sg13g2_nor2_1 _26513_ (.A(_07799_),
    .B(_07801_),
    .Y(_07802_));
 sg13g2_nand3_1 _26514_ (.B(_07796_),
    .C(_07802_),
    .A(net518),
    .Y(_07803_));
 sg13g2_a21o_1 _26515_ (.A2(_07802_),
    .A1(_07796_),
    .B1(_07780_),
    .X(_07804_));
 sg13g2_or2_1 _26516_ (.X(_07805_),
    .B(_07776_),
    .A(net455));
 sg13g2_nand2_1 _26517_ (.Y(_07806_),
    .A(net455),
    .B(_07776_));
 sg13g2_o21ai_1 _26518_ (.B1(_07806_),
    .Y(_07807_),
    .A1(_07765_),
    .A2(_07769_));
 sg13g2_nand2_1 _26519_ (.Y(_07808_),
    .A(_07805_),
    .B(_07807_));
 sg13g2_mux2_1 _26520_ (.A0(_07803_),
    .A1(_07804_),
    .S(_07808_),
    .X(_07809_));
 sg13g2_inv_1 _26521_ (.Y(_07810_),
    .A(_07632_));
 sg13g2_a221oi_1 _26522_ (.B2(\exec.memory_input[4] ),
    .C1(net479),
    .B1(_07651_),
    .A1(_09864_),
    .Y(_07811_),
    .A2(_07810_));
 sg13g2_a22oi_1 _26523_ (.Y(_07812_),
    .B1(_07695_),
    .B2(net510),
    .A2(_07648_),
    .A1(net471));
 sg13g2_nand3b_1 _26524_ (.B(_07634_),
    .C(_07644_),
    .Y(_07813_),
    .A_N(net523));
 sg13g2_a21oi_1 _26525_ (.A1(_09864_),
    .A2(_07339_),
    .Y(_07814_),
    .B1(_07690_));
 sg13g2_nand2_1 _26526_ (.Y(_07815_),
    .A(_07339_),
    .B(_07637_));
 sg13g2_a22oi_1 _26527_ (.Y(_07816_),
    .B1(_07815_),
    .B2(net496),
    .A2(_07683_),
    .A1(_07340_));
 sg13g2_o21ai_1 _26528_ (.B1(_07816_),
    .Y(_07817_),
    .A1(_07813_),
    .A2(_07814_));
 sg13g2_and3_1 _26529_ (.X(_07818_),
    .A(_07811_),
    .B(_07812_),
    .C(_07817_));
 sg13g2_or4_1 _26530_ (.A(_07625_),
    .B(net518),
    .C(_07635_),
    .D(_07637_),
    .X(_07819_));
 sg13g2_buf_1 _26531_ (.A(_07819_),
    .X(_07820_));
 sg13g2_nor2_1 _26532_ (.A(_09893_),
    .B(_07820_),
    .Y(_07821_));
 sg13g2_a21o_1 _26533_ (.A2(_07818_),
    .A1(_07809_),
    .B1(_07821_),
    .X(_07822_));
 sg13g2_buf_1 _26534_ (.A(_07822_),
    .X(_07823_));
 sg13g2_buf_1 _26535_ (.A(_07823_),
    .X(_07824_));
 sg13g2_nand2_1 _26536_ (.Y(_07825_),
    .A(_07789_),
    .B(net102));
 sg13g2_mux2_1 _26537_ (.A0(_07791_),
    .A1(_07825_),
    .S(net65),
    .X(_02527_));
 sg13g2_nand2_1 _26538_ (.Y(_07826_),
    .A(_07797_),
    .B(_07671_));
 sg13g2_nor2_1 _26539_ (.A(_07339_),
    .B(_07793_),
    .Y(_07827_));
 sg13g2_a221oi_1 _26540_ (.B2(_07827_),
    .C1(_07801_),
    .B1(_07826_),
    .A1(net455),
    .Y(_07828_),
    .A2(_07776_));
 sg13g2_o21ai_1 _26541_ (.B1(_07828_),
    .Y(_07829_),
    .A1(_07765_),
    .A2(_07769_));
 sg13g2_or4_1 _26542_ (.A(net455),
    .B(_07776_),
    .C(_07799_),
    .D(_07801_),
    .X(_07830_));
 sg13g2_and2_1 _26543_ (.A(_07796_),
    .B(_07830_),
    .X(_07831_));
 sg13g2_o21ai_1 _26544_ (.B1(_10199_),
    .Y(_07832_),
    .A1(_10197_),
    .A2(net517));
 sg13g2_nand3_1 _26545_ (.B(_10201_),
    .C(_07671_),
    .A(net472),
    .Y(_07833_));
 sg13g2_a21oi_2 _26546_ (.B1(_07553_),
    .Y(_07834_),
    .A2(_07833_),
    .A1(_07832_));
 sg13g2_xnor2_1 _26547_ (.Y(_07835_),
    .A(net454),
    .B(_07834_));
 sg13g2_a221oi_1 _26548_ (.B2(_07831_),
    .C1(_07835_),
    .B1(_07829_),
    .A1(net524),
    .Y(_07836_),
    .A2(_07627_));
 sg13g2_nand4_1 _26549_ (.B(_07829_),
    .C(_07831_),
    .A(_07629_),
    .Y(_07837_),
    .D(_07835_));
 sg13g2_mux2_1 _26550_ (.A0(_07643_),
    .A1(_07685_),
    .S(net454),
    .X(_07838_));
 sg13g2_a21oi_1 _26551_ (.A1(net472),
    .A2(_07643_),
    .Y(_07839_),
    .B1(_07838_));
 sg13g2_nand2b_1 _26552_ (.Y(_07840_),
    .B(_07839_),
    .A_N(_07645_));
 sg13g2_o21ai_1 _26553_ (.B1(net472),
    .Y(_07841_),
    .A1(_07387_),
    .A2(_07683_));
 sg13g2_inv_1 _26554_ (.Y(_07842_),
    .A(_07695_));
 sg13g2_a221oi_1 _26555_ (.B2(\exec.memory_input[5] ),
    .C1(_07639_),
    .B1(_07651_),
    .A1(net483),
    .Y(_07843_),
    .A2(_07648_));
 sg13g2_o21ai_1 _26556_ (.B1(_07843_),
    .Y(_07844_),
    .A1(net496),
    .A2(_07842_));
 sg13g2_a221oi_1 _26557_ (.B2(_07841_),
    .C1(_07844_),
    .B1(_07840_),
    .A1(net454),
    .Y(_07845_),
    .A2(net523));
 sg13g2_nand3b_1 _26558_ (.B(_07837_),
    .C(_07845_),
    .Y(_07846_),
    .A_N(_07836_));
 sg13g2_o21ai_1 _26559_ (.B1(_07846_),
    .Y(_07847_),
    .A1(_09869_),
    .A2(_07820_));
 sg13g2_buf_2 _26560_ (.A(_07847_),
    .X(_07848_));
 sg13g2_buf_1 _26561_ (.A(_07848_),
    .X(_07849_));
 sg13g2_buf_1 _26562_ (.A(net1298),
    .X(_07850_));
 sg13g2_a221oi_1 _26563_ (.B2(\stack[0][5] ),
    .C1(_07589_),
    .B1(_07617_),
    .A1(net1221),
    .Y(_07851_),
    .A2(net509));
 sg13g2_a21o_1 _26564_ (.A2(net90),
    .A1(_07589_),
    .B1(_07851_),
    .X(_07852_));
 sg13g2_o21ai_1 _26565_ (.B1(_07852_),
    .Y(_02528_),
    .A1(net446),
    .A2(_07614_));
 sg13g2_buf_1 _26566_ (.A(_10017_),
    .X(_07853_));
 sg13g2_buf_1 _26567_ (.A(net1220),
    .X(_07854_));
 sg13g2_a22oi_1 _26568_ (.Y(_07855_),
    .B1(_07617_),
    .B2(\stack[0][6] ),
    .A2(net509),
    .A1(net880));
 sg13g2_buf_1 _26569_ (.A(net483),
    .X(_07856_));
 sg13g2_buf_1 _26570_ (.A(net451),
    .X(_07857_));
 sg13g2_a221oi_1 _26571_ (.B2(\exec.memory_input[6] ),
    .C1(net479),
    .B1(_07651_),
    .A1(net483),
    .Y(_07858_),
    .A2(_07810_));
 sg13g2_a22oi_1 _26572_ (.Y(_07859_),
    .B1(_07695_),
    .B2(net471),
    .A2(_07648_),
    .A1(net474));
 sg13g2_and2_1 _26573_ (.A(_07395_),
    .B(_07415_),
    .X(_07860_));
 sg13g2_buf_1 _26574_ (.A(_07860_),
    .X(_07861_));
 sg13g2_a21oi_1 _26575_ (.A1(net497),
    .A2(_07861_),
    .Y(_07862_),
    .B1(_07690_));
 sg13g2_nand2_1 _26576_ (.Y(_07863_),
    .A(_07861_),
    .B(_07637_));
 sg13g2_a22oi_1 _26577_ (.Y(_07864_),
    .B1(_07863_),
    .B2(_10134_),
    .A2(_07683_),
    .A1(_07416_));
 sg13g2_o21ai_1 _26578_ (.B1(_07864_),
    .Y(_07865_),
    .A1(_07813_),
    .A2(_07862_));
 sg13g2_nand3_1 _26579_ (.B(_07859_),
    .C(_07865_),
    .A(_07858_),
    .Y(_07866_));
 sg13g2_nand2b_1 _26580_ (.Y(_07867_),
    .B(net479),
    .A_N(_09871_));
 sg13g2_nand2_1 _26581_ (.Y(_07868_),
    .A(_07866_),
    .B(_07867_));
 sg13g2_nor2b_1 _26582_ (.A(_07834_),
    .B_N(_07828_),
    .Y(_07869_));
 sg13g2_a21oi_1 _26583_ (.A1(_07796_),
    .A2(_07830_),
    .Y(_07870_),
    .B1(_07834_));
 sg13g2_a221oi_1 _26584_ (.B2(_07869_),
    .C1(_07870_),
    .B1(_07771_),
    .A1(_07363_),
    .Y(_07871_),
    .A2(_07385_));
 sg13g2_buf_1 _26585_ (.A(_07871_),
    .X(_07872_));
 sg13g2_nand3_1 _26586_ (.B(_07796_),
    .C(_07834_),
    .A(_07805_),
    .Y(_07873_));
 sg13g2_or2_1 _26587_ (.X(_07874_),
    .B(_07801_),
    .A(_07799_));
 sg13g2_a221oi_1 _26588_ (.B2(_07833_),
    .C1(net533),
    .B1(_07832_),
    .A1(_07794_),
    .Y(_07875_),
    .A2(_07795_));
 sg13g2_and2_1 _26589_ (.A(_07313_),
    .B(_07776_),
    .X(_07876_));
 sg13g2_a22oi_1 _26590_ (.Y(_07877_),
    .B1(_07875_),
    .B2(_07876_),
    .A2(_07834_),
    .A1(_07874_));
 sg13g2_o21ai_1 _26591_ (.B1(_07877_),
    .Y(_07878_),
    .A1(_07771_),
    .A2(_07873_));
 sg13g2_buf_1 _26592_ (.A(_07878_),
    .X(_07879_));
 sg13g2_nand3_1 _26593_ (.B(_07416_),
    .C(net524),
    .A(_09822_),
    .Y(_07880_));
 sg13g2_nand3_1 _26594_ (.B(_07416_),
    .C(net524),
    .A(_10134_),
    .Y(_07881_));
 sg13g2_a21oi_1 _26595_ (.A1(net472),
    .A2(_10197_),
    .Y(_07882_),
    .B1(net517));
 sg13g2_mux2_1 _26596_ (.A0(_07880_),
    .A1(_07881_),
    .S(_07882_),
    .X(_07883_));
 sg13g2_nor2_1 _26597_ (.A(net497),
    .B(_07772_),
    .Y(_07884_));
 sg13g2_o21ai_1 _26598_ (.B1(_07884_),
    .Y(_07885_),
    .A1(net471),
    .A2(_10201_));
 sg13g2_nand4_1 _26599_ (.B(net472),
    .C(_10197_),
    .A(net497),
    .Y(_07886_),
    .D(net524));
 sg13g2_nand2_1 _26600_ (.Y(_07887_),
    .A(net497),
    .B(net517));
 sg13g2_nand4_1 _26601_ (.B(_07885_),
    .C(_07886_),
    .A(_07861_),
    .Y(_07888_),
    .D(_07887_));
 sg13g2_buf_1 _26602_ (.A(_07888_),
    .X(_07889_));
 sg13g2_nand2_1 _26603_ (.Y(_07890_),
    .A(_07883_),
    .B(_07889_));
 sg13g2_nand2_1 _26604_ (.Y(_07891_),
    .A(net518),
    .B(_07890_));
 sg13g2_or3_1 _26605_ (.A(_07872_),
    .B(_07879_),
    .C(_07891_),
    .X(_07892_));
 sg13g2_buf_2 _26606_ (.A(_07892_),
    .X(_07893_));
 sg13g2_nor2_1 _26607_ (.A(_07780_),
    .B(_07890_),
    .Y(_07894_));
 sg13g2_nor3_1 _26608_ (.A(net454),
    .B(_07780_),
    .C(_07890_),
    .Y(_07895_));
 sg13g2_a21oi_1 _26609_ (.A1(_07771_),
    .A2(_07869_),
    .Y(_07896_),
    .B1(_07870_));
 sg13g2_a22oi_1 _26610_ (.Y(_07897_),
    .B1(_07895_),
    .B2(_07896_),
    .A2(_07894_),
    .A1(_07879_));
 sg13g2_nand3_1 _26611_ (.B(_07893_),
    .C(_07897_),
    .A(_07868_),
    .Y(_07898_));
 sg13g2_buf_8 _26612_ (.A(_07898_),
    .X(_07899_));
 sg13g2_buf_8 _26613_ (.A(_07899_),
    .X(_07900_));
 sg13g2_a22oi_1 _26614_ (.Y(_07901_),
    .B1(net46),
    .B2(net65),
    .A2(_07756_),
    .A1(net405));
 sg13g2_o21ai_1 _26615_ (.B1(_07901_),
    .Y(_02529_),
    .A1(net65),
    .A2(_07855_));
 sg13g2_inv_1 _26616_ (.Y(_07902_),
    .A(_07447_));
 sg13g2_and3_1 _26617_ (.X(_07903_),
    .A(_09659_),
    .B(_09867_),
    .C(_07671_));
 sg13g2_a21oi_1 _26618_ (.A1(_09867_),
    .A2(_07671_),
    .Y(_07904_),
    .B1(net474));
 sg13g2_nor3_1 _26619_ (.A(net533),
    .B(_07903_),
    .C(_07904_),
    .Y(_07905_));
 sg13g2_xnor2_1 _26620_ (.Y(_07906_),
    .A(_07902_),
    .B(_07905_));
 sg13g2_nor2_1 _26621_ (.A(_07780_),
    .B(_07906_),
    .Y(_07907_));
 sg13g2_xnor2_1 _26622_ (.Y(_07908_),
    .A(net497),
    .B(_07882_));
 sg13g2_nor2_1 _26623_ (.A(net533),
    .B(_07908_),
    .Y(_07909_));
 sg13g2_nor3_1 _26624_ (.A(_07909_),
    .B(_07872_),
    .C(_07879_),
    .Y(_07910_));
 sg13g2_nor3_1 _26625_ (.A(net454),
    .B(net533),
    .C(_07908_),
    .Y(_07911_));
 sg13g2_a221oi_1 _26626_ (.B2(_07896_),
    .C1(_07416_),
    .B1(_07911_),
    .A1(_07909_),
    .Y(_07912_),
    .A2(_07879_));
 sg13g2_or2_1 _26627_ (.X(_07913_),
    .B(_07912_),
    .A(_07910_));
 sg13g2_nor2_1 _26628_ (.A(_07872_),
    .B(_07879_),
    .Y(_07914_));
 sg13g2_nand3_1 _26629_ (.B(_07889_),
    .C(_07906_),
    .A(net518),
    .Y(_07915_));
 sg13g2_nor4_1 _26630_ (.A(_07861_),
    .B(net533),
    .C(_07780_),
    .D(_07908_),
    .Y(_07916_));
 sg13g2_a221oi_1 _26631_ (.B2(net483),
    .C1(net479),
    .B1(_07695_),
    .A1(\exec.memory_input[7] ),
    .Y(_07917_),
    .A2(_07651_));
 sg13g2_a21oi_1 _26632_ (.A1(_07447_),
    .A2(_07643_),
    .Y(_07918_),
    .B1(_07645_));
 sg13g2_or2_1 _26633_ (.X(_07919_),
    .B(_07918_),
    .A(_10138_));
 sg13g2_nand2_1 _26634_ (.Y(_07920_),
    .A(net474),
    .B(_07685_));
 sg13g2_o21ai_1 _26635_ (.B1(_07920_),
    .Y(_07921_),
    .A1(net474),
    .A2(_07683_));
 sg13g2_o21ai_1 _26636_ (.B1(_07902_),
    .Y(_07922_),
    .A1(net523),
    .A2(_07921_));
 sg13g2_nand3_1 _26637_ (.B(_07919_),
    .C(_07922_),
    .A(_07917_),
    .Y(_07923_));
 sg13g2_nand2b_1 _26638_ (.Y(_07924_),
    .B(net479),
    .A_N(net1309));
 sg13g2_a22oi_1 _26639_ (.Y(_07925_),
    .B1(_07923_),
    .B2(_07924_),
    .A2(_07916_),
    .A1(_07906_));
 sg13g2_o21ai_1 _26640_ (.B1(_07925_),
    .Y(_07926_),
    .A1(_07914_),
    .A2(_07915_));
 sg13g2_a21oi_1 _26641_ (.A1(_07907_),
    .A2(_07913_),
    .Y(_07927_),
    .B1(_07926_));
 sg13g2_buf_2 _26642_ (.A(_07927_),
    .X(_07928_));
 sg13g2_buf_8 _26643_ (.A(_07928_),
    .X(_07929_));
 sg13g2_buf_1 _26644_ (.A(_10024_),
    .X(_07930_));
 sg13g2_nor2_1 _26645_ (.A(_10138_),
    .B(_07614_),
    .Y(_07931_));
 sg13g2_a221oi_1 _26646_ (.B2(\stack[0][7] ),
    .C1(_07931_),
    .B1(_07617_),
    .A1(net1219),
    .Y(_07932_),
    .A2(net509));
 sg13g2_nor2b_1 _26647_ (.A(net65),
    .B_N(_07932_),
    .Y(_07933_));
 sg13g2_a21oi_1 _26648_ (.A1(net65),
    .A2(net45),
    .Y(_02530_),
    .B1(_07933_));
 sg13g2_buf_8 _26649_ (.A(net136),
    .X(_07934_));
 sg13g2_nor2_1 _26650_ (.A(net128),
    .B(_07559_),
    .Y(_07935_));
 sg13g2_buf_2 _26651_ (.A(_07935_),
    .X(_07936_));
 sg13g2_nor2b_1 _26652_ (.A(_07604_),
    .B_N(net137),
    .Y(_07937_));
 sg13g2_buf_2 _26653_ (.A(_07937_),
    .X(_07938_));
 sg13g2_nand2_1 _26654_ (.Y(_07939_),
    .A(_07936_),
    .B(_07938_));
 sg13g2_nor2_1 _26655_ (.A(_09712_),
    .B(_07487_),
    .Y(_07940_));
 sg13g2_nand2_1 _26656_ (.Y(_07941_),
    .A(_07476_),
    .B(_07940_));
 sg13g2_buf_2 _26657_ (.A(_07941_),
    .X(_07942_));
 sg13g2_nand2_1 _26658_ (.Y(_07943_),
    .A(_09717_),
    .B(_07598_));
 sg13g2_nor2_1 _26659_ (.A(_07942_),
    .B(_07943_),
    .Y(_07944_));
 sg13g2_buf_1 _26660_ (.A(_07944_),
    .X(_07945_));
 sg13g2_nor2_1 _26661_ (.A(_07575_),
    .B(_07750_),
    .Y(_07946_));
 sg13g2_buf_1 _26662_ (.A(_07946_),
    .X(_07947_));
 sg13g2_inv_1 _26663_ (.Y(_07948_),
    .A(_07494_));
 sg13g2_nand2_1 _26664_ (.Y(_07949_),
    .A(net406),
    .B(_07492_));
 sg13g2_a21o_1 _26665_ (.A2(_07499_),
    .A1(net406),
    .B1(_07500_),
    .X(_07950_));
 sg13g2_a221oi_1 _26666_ (.B2(_07949_),
    .C1(_07950_),
    .B1(_07948_),
    .A1(_07516_),
    .Y(_07951_),
    .A2(_07528_));
 sg13g2_buf_2 _26667_ (.A(_07951_),
    .X(_07952_));
 sg13g2_and4_1 _26668_ (.A(net128),
    .B(net135),
    .C(net299),
    .D(_07952_),
    .X(_07953_));
 sg13g2_nor3_1 _26669_ (.A(net1270),
    .B(_07945_),
    .C(_07953_),
    .Y(_07954_));
 sg13g2_buf_2 _26670_ (.A(_07954_),
    .X(_07955_));
 sg13g2_nand2_1 _26671_ (.Y(_07956_),
    .A(_07939_),
    .B(_07955_));
 sg13g2_buf_2 _26672_ (.A(_07956_),
    .X(_07957_));
 sg13g2_and2_1 _26673_ (.A(_07936_),
    .B(_07938_),
    .X(_07958_));
 sg13g2_buf_2 _26674_ (.A(_07958_),
    .X(_07959_));
 sg13g2_buf_1 _26675_ (.A(_10165_),
    .X(_07960_));
 sg13g2_buf_1 _26676_ (.A(net1302),
    .X(_07961_));
 sg13g2_and3_1 _26677_ (.X(_07962_),
    .A(net1218),
    .B(_07939_),
    .C(net508));
 sg13g2_a221oi_1 _26678_ (.B2(net478),
    .C1(_07962_),
    .B1(_07953_),
    .A1(net134),
    .Y(_07963_),
    .A2(_07959_));
 sg13g2_nor2_1 _26679_ (.A(\stack[10][0] ),
    .B(_07957_),
    .Y(_07964_));
 sg13g2_a21oi_1 _26680_ (.A1(_07957_),
    .A2(_07963_),
    .Y(_02531_),
    .B1(_07964_));
 sg13g2_buf_8 _26681_ (.A(_07959_),
    .X(_07965_));
 sg13g2_nand2_1 _26682_ (.Y(_07966_),
    .A(net1225),
    .B(net508));
 sg13g2_nand2_1 _26683_ (.Y(_07967_),
    .A(_07606_),
    .B(_07609_));
 sg13g2_buf_2 _26684_ (.A(_07967_),
    .X(_07968_));
 sg13g2_buf_8 _26685_ (.A(_07968_),
    .X(_07969_));
 sg13g2_nand2b_1 _26686_ (.Y(_07970_),
    .B(_07952_),
    .A_N(_07750_));
 sg13g2_buf_1 _26687_ (.A(_07970_),
    .X(_07971_));
 sg13g2_nor3_1 _26688_ (.A(_07754_),
    .B(net117),
    .C(_07971_),
    .Y(_07972_));
 sg13g2_buf_2 _26689_ (.A(_07972_),
    .X(_07973_));
 sg13g2_a22oi_1 _26690_ (.Y(_07974_),
    .B1(_07973_),
    .B2(net473),
    .A2(_07959_),
    .A1(net119));
 sg13g2_o21ai_1 _26691_ (.B1(_07974_),
    .Y(_07975_),
    .A1(net44),
    .A2(_07966_));
 sg13g2_mux2_1 _26692_ (.A0(_09687_),
    .A1(_07975_),
    .S(_07957_),
    .X(_02532_));
 sg13g2_buf_1 _26693_ (.A(net1301),
    .X(_07976_));
 sg13g2_nand2_1 _26694_ (.Y(_07977_),
    .A(net1217),
    .B(net508));
 sg13g2_buf_1 _26695_ (.A(net485),
    .X(_07978_));
 sg13g2_a22oi_1 _26696_ (.Y(_07979_),
    .B1(_07973_),
    .B2(net450),
    .A2(_07959_),
    .A1(net118));
 sg13g2_o21ai_1 _26697_ (.B1(_07979_),
    .Y(_07980_),
    .A1(net44),
    .A2(_07977_));
 sg13g2_mux2_1 _26698_ (.A0(\stack[10][2] ),
    .A1(_07980_),
    .S(_07957_),
    .X(_02533_));
 sg13g2_buf_2 _26699_ (.A(_07783_),
    .X(_07981_));
 sg13g2_and3_1 _26700_ (.X(_07982_),
    .A(net1223),
    .B(_07939_),
    .C(net508));
 sg13g2_a221oi_1 _26701_ (.B2(net492),
    .C1(_07982_),
    .B1(_07973_),
    .A1(net101),
    .Y(_07983_),
    .A2(_07959_));
 sg13g2_nor2_1 _26702_ (.A(\stack[10][3] ),
    .B(_07957_),
    .Y(_07984_));
 sg13g2_a21oi_1 _26703_ (.A1(_07957_),
    .A2(_07983_),
    .Y(_02534_),
    .B1(_07984_));
 sg13g2_buf_1 _26704_ (.A(_07823_),
    .X(_07985_));
 sg13g2_a21oi_1 _26705_ (.A1(net484),
    .A2(_07973_),
    .Y(_07986_),
    .B1(_07955_));
 sg13g2_a21oi_1 _26706_ (.A1(net1222),
    .A2(net508),
    .Y(_07987_),
    .B1(net44));
 sg13g2_inv_1 _26707_ (.Y(_07988_),
    .A(_07955_));
 sg13g2_nor3_1 _26708_ (.A(\stack[10][4] ),
    .B(net44),
    .C(_07988_),
    .Y(_07989_));
 sg13g2_a221oi_1 _26709_ (.B2(_07987_),
    .C1(_07989_),
    .B1(_07986_),
    .A1(_07985_),
    .Y(_02535_),
    .A2(net44));
 sg13g2_buf_1 _26710_ (.A(_07848_),
    .X(_07990_));
 sg13g2_buf_1 _26711_ (.A(net1298),
    .X(_07991_));
 sg13g2_a21oi_1 _26712_ (.A1(net1216),
    .A2(net508),
    .Y(_07992_),
    .B1(_07955_));
 sg13g2_a21o_1 _26713_ (.A2(_07973_),
    .A1(net471),
    .B1(_07959_),
    .X(_07993_));
 sg13g2_inv_1 _26714_ (.Y(_07994_),
    .A(_07993_));
 sg13g2_nor2_1 _26715_ (.A(\stack[10][5] ),
    .B(_07957_),
    .Y(_07995_));
 sg13g2_a221oi_1 _26716_ (.B2(_07994_),
    .C1(_07995_),
    .B1(_07992_),
    .A1(_07990_),
    .Y(_02536_),
    .A2(net44));
 sg13g2_and3_1 _26717_ (.X(_07996_),
    .A(_07868_),
    .B(_07893_),
    .C(_07897_));
 sg13g2_buf_2 _26718_ (.A(_07996_),
    .X(_07997_));
 sg13g2_buf_1 _26719_ (.A(net1220),
    .X(_07998_));
 sg13g2_a21oi_1 _26720_ (.A1(net879),
    .A2(net508),
    .Y(_07999_),
    .B1(_07955_));
 sg13g2_buf_1 _26721_ (.A(net483),
    .X(_08000_));
 sg13g2_a21oi_1 _26722_ (.A1(net449),
    .A2(_07973_),
    .Y(_08001_),
    .B1(_07965_));
 sg13g2_nor2_1 _26723_ (.A(\stack[10][6] ),
    .B(_07957_),
    .Y(_08002_));
 sg13g2_a221oi_1 _26724_ (.B2(_08001_),
    .C1(_08002_),
    .B1(_07999_),
    .A1(_07997_),
    .Y(_02537_),
    .A2(net44));
 sg13g2_buf_8 _26725_ (.A(_07928_),
    .X(_08003_));
 sg13g2_nand2_1 _26726_ (.Y(_08004_),
    .A(\stack[10][7] ),
    .B(_07955_));
 sg13g2_buf_1 _26727_ (.A(_10024_),
    .X(_08005_));
 sg13g2_buf_1 _26728_ (.A(net445),
    .X(_08006_));
 sg13g2_a221oi_1 _26729_ (.B2(net298),
    .C1(_07965_),
    .B1(_07973_),
    .A1(net1215),
    .Y(_08007_),
    .A2(net508));
 sg13g2_a22oi_1 _26730_ (.Y(_02538_),
    .B1(_08004_),
    .B2(_08007_),
    .A2(net44),
    .A1(net43));
 sg13g2_buf_8 _26731_ (.A(_07952_),
    .X(_08008_));
 sg13g2_nor2_1 _26732_ (.A(net143),
    .B(net138),
    .Y(_08009_));
 sg13g2_buf_2 _26733_ (.A(_08009_),
    .X(_08010_));
 sg13g2_nor2_1 _26734_ (.A(_07574_),
    .B(_07750_),
    .Y(_08011_));
 sg13g2_buf_1 _26735_ (.A(_08011_),
    .X(_08012_));
 sg13g2_nand3_1 _26736_ (.B(_08010_),
    .C(net404),
    .A(net127),
    .Y(_08013_));
 sg13g2_buf_1 _26737_ (.A(_08013_),
    .X(_08014_));
 sg13g2_nand2_1 _26738_ (.Y(_08015_),
    .A(_07114_),
    .B(_07598_));
 sg13g2_buf_1 _26739_ (.A(_08015_),
    .X(_08016_));
 sg13g2_buf_1 _26740_ (.A(_08016_),
    .X(_08017_));
 sg13g2_nor2_1 _26741_ (.A(_07942_),
    .B(net516),
    .Y(_08018_));
 sg13g2_buf_2 _26742_ (.A(_08018_),
    .X(_08019_));
 sg13g2_nand2_1 _26743_ (.Y(_08020_),
    .A(net1302),
    .B(_08019_));
 sg13g2_nand2_1 _26744_ (.Y(_08021_),
    .A(_07654_),
    .B(_07661_));
 sg13g2_o21ai_1 _26745_ (.B1(_08021_),
    .Y(_08022_),
    .A1(net1275),
    .A2(_07820_));
 sg13g2_buf_1 _26746_ (.A(_08022_),
    .X(_08023_));
 sg13g2_a21oi_1 _26747_ (.A1(_07387_),
    .A2(net406),
    .Y(_08024_),
    .B1(_07542_));
 sg13g2_a21oi_1 _26748_ (.A1(_07577_),
    .A2(_08024_),
    .Y(_08025_),
    .B1(_07570_));
 sg13g2_nand2_1 _26749_ (.Y(_08026_),
    .A(_07574_),
    .B(_07581_));
 sg13g2_or2_1 _26750_ (.X(_08027_),
    .B(_08026_),
    .A(_08025_));
 sg13g2_buf_2 _26751_ (.A(_08027_),
    .X(_08028_));
 sg13g2_buf_1 _26752_ (.A(_08028_),
    .X(_08029_));
 sg13g2_nor3_1 _26753_ (.A(_07531_),
    .B(net117),
    .C(net126),
    .Y(_08030_));
 sg13g2_buf_2 _26754_ (.A(_08030_),
    .X(_08031_));
 sg13g2_mux2_1 _26755_ (.A0(_08020_),
    .A1(_08023_),
    .S(_08031_),
    .X(_08032_));
 sg13g2_o21ai_1 _26756_ (.B1(_08032_),
    .Y(_08033_),
    .A1(net487),
    .A2(_08014_));
 sg13g2_or2_1 _26757_ (.X(_08034_),
    .B(_07750_),
    .A(_07574_));
 sg13g2_buf_1 _26758_ (.A(_08034_),
    .X(_08035_));
 sg13g2_buf_1 _26759_ (.A(_08035_),
    .X(_08036_));
 sg13g2_a21oi_1 _26760_ (.A1(net297),
    .A2(net126),
    .Y(_08037_),
    .B1(net117));
 sg13g2_o21ai_1 _26761_ (.B1(net1304),
    .Y(_08038_),
    .A1(_07942_),
    .A2(net516));
 sg13g2_a21oi_1 _26762_ (.A1(net127),
    .A2(_08037_),
    .Y(_08039_),
    .B1(_08038_));
 sg13g2_buf_1 _26763_ (.A(_08039_),
    .X(_08040_));
 sg13g2_mux2_1 _26764_ (.A0(_08033_),
    .A1(\stack[11][0] ),
    .S(net64),
    .X(_02539_));
 sg13g2_inv_1 _26765_ (.Y(_08041_),
    .A(\stack[11][1] ));
 sg13g2_inv_1 _26766_ (.Y(_08042_),
    .A(_08014_));
 sg13g2_buf_8 _26767_ (.A(_08031_),
    .X(_08043_));
 sg13g2_nand2b_1 _26768_ (.Y(_08044_),
    .B(net63),
    .A_N(_07700_));
 sg13g2_a21o_1 _26769_ (.A2(_08019_),
    .A1(net1299),
    .B1(_08031_),
    .X(_08045_));
 sg13g2_a221oi_1 _26770_ (.B2(_08045_),
    .C1(net64),
    .B1(_08044_),
    .A1(net447),
    .Y(_08046_),
    .A2(_08042_));
 sg13g2_a21oi_1 _26771_ (.A1(_08041_),
    .A2(net64),
    .Y(_02540_),
    .B1(_08046_));
 sg13g2_inv_1 _26772_ (.Y(_08047_),
    .A(\stack[11][2] ));
 sg13g2_nand2b_1 _26773_ (.Y(_08048_),
    .B(net63),
    .A_N(_07738_));
 sg13g2_a21o_1 _26774_ (.A2(_08019_),
    .A1(net1301),
    .B1(_08031_),
    .X(_08049_));
 sg13g2_a221oi_1 _26775_ (.B2(_08049_),
    .C1(net64),
    .B1(_08048_),
    .A1(net452),
    .Y(_08050_),
    .A2(_08042_));
 sg13g2_a21oi_1 _26776_ (.A1(_08047_),
    .A2(net64),
    .Y(_02541_),
    .B1(_08050_));
 sg13g2_inv_1 _26777_ (.Y(_08051_),
    .A(\stack[11][3] ));
 sg13g2_nand2b_1 _26778_ (.Y(_08052_),
    .B(net63),
    .A_N(_07783_));
 sg13g2_a21o_1 _26779_ (.A2(_08019_),
    .A1(net1300),
    .B1(_08031_),
    .X(_08053_));
 sg13g2_a221oi_1 _26780_ (.B2(_08053_),
    .C1(_08039_),
    .B1(_08052_),
    .A1(net492),
    .Y(_08054_),
    .A2(_08042_));
 sg13g2_a21oi_1 _26781_ (.A1(_08051_),
    .A2(net64),
    .Y(_02542_),
    .B1(_08054_));
 sg13g2_inv_1 _26782_ (.Y(_08055_),
    .A(\stack[11][4] ));
 sg13g2_nor2b_1 _26783_ (.A(_08031_),
    .B_N(_08019_),
    .Y(_08056_));
 sg13g2_a221oi_1 _26784_ (.B2(net1222),
    .C1(_08039_),
    .B1(_08056_),
    .A1(net484),
    .Y(_08057_),
    .A2(_08042_));
 sg13g2_a21oi_2 _26785_ (.B1(_07821_),
    .Y(_08058_),
    .A2(_07818_),
    .A1(_07809_));
 sg13g2_nand2_1 _26786_ (.Y(_08059_),
    .A(_08058_),
    .B(net63));
 sg13g2_a22oi_1 _26787_ (.Y(_02543_),
    .B1(_08057_),
    .B2(_08059_),
    .A2(net64),
    .A1(_08055_));
 sg13g2_buf_1 _26788_ (.A(net471),
    .X(_08060_));
 sg13g2_buf_1 _26789_ (.A(_07848_),
    .X(_08061_));
 sg13g2_buf_1 _26790_ (.A(net1298),
    .X(_08062_));
 sg13g2_inv_1 _26791_ (.Y(_08063_),
    .A(\stack[11][5] ));
 sg13g2_nor2_1 _26792_ (.A(_08063_),
    .B(_08038_),
    .Y(_08064_));
 sg13g2_a221oi_1 _26793_ (.B2(_08064_),
    .C1(net63),
    .B1(_08014_),
    .A1(net1214),
    .Y(_08065_),
    .A2(_08019_));
 sg13g2_a21oi_1 _26794_ (.A1(net88),
    .A2(net63),
    .Y(_08066_),
    .B1(_08065_));
 sg13g2_a21o_1 _26795_ (.A2(_08042_),
    .A1(net403),
    .B1(_08066_),
    .X(_02544_));
 sg13g2_inv_1 _26796_ (.Y(_08067_),
    .A(\stack[11][6] ));
 sg13g2_buf_8 _26797_ (.A(_07899_),
    .X(_08068_));
 sg13g2_nand2_1 _26798_ (.Y(_08069_),
    .A(net42),
    .B(net63));
 sg13g2_nand2_1 _26799_ (.Y(_08070_),
    .A(net1220),
    .B(_08019_));
 sg13g2_nand4_1 _26800_ (.B(net127),
    .C(_08010_),
    .A(net483),
    .Y(_08071_),
    .D(net404));
 sg13g2_o21ai_1 _26801_ (.B1(_08071_),
    .Y(_08072_),
    .A1(_08043_),
    .A2(_08070_));
 sg13g2_nor2_1 _26802_ (.A(_08040_),
    .B(_08072_),
    .Y(_08073_));
 sg13g2_a22oi_1 _26803_ (.Y(_02545_),
    .B1(_08069_),
    .B2(_08073_),
    .A2(net64),
    .A1(_08067_));
 sg13g2_inv_1 _26804_ (.Y(_08074_),
    .A(\stack[11][7] ));
 sg13g2_buf_8 _26805_ (.A(_07928_),
    .X(_08075_));
 sg13g2_buf_1 _26806_ (.A(_10024_),
    .X(_08076_));
 sg13g2_nand2_1 _26807_ (.Y(_08077_),
    .A(net1213),
    .B(_08019_));
 sg13g2_o21ai_1 _26808_ (.B1(_08077_),
    .Y(_08078_),
    .A1(_10138_),
    .A2(_08014_));
 sg13g2_nor3_1 _26809_ (.A(_08039_),
    .B(_08043_),
    .C(_08078_),
    .Y(_08079_));
 sg13g2_a221oi_1 _26810_ (.B2(net41),
    .C1(_08079_),
    .B1(net63),
    .A1(_08074_),
    .Y(_02546_),
    .A2(_08040_));
 sg13g2_inv_1 _26811_ (.Y(_08080_),
    .A(\stack[12][0] ));
 sg13g2_buf_8 _26812_ (.A(net135),
    .X(_08081_));
 sg13g2_and4_1 _26813_ (.A(net128),
    .B(net125),
    .C(net127),
    .D(net137),
    .X(_08082_));
 sg13g2_buf_8 _26814_ (.A(_08082_),
    .X(_08083_));
 sg13g2_nor2_1 _26815_ (.A(_07487_),
    .B(_07532_),
    .Y(_08084_));
 sg13g2_nand2_1 _26816_ (.Y(_08085_),
    .A(_07476_),
    .B(_08084_));
 sg13g2_buf_2 _26817_ (.A(_08085_),
    .X(_08086_));
 sg13g2_nor2_1 _26818_ (.A(_07600_),
    .B(_08086_),
    .Y(_08087_));
 sg13g2_buf_1 _26819_ (.A(_08087_),
    .X(_08088_));
 sg13g2_buf_1 _26820_ (.A(_07612_),
    .X(_08089_));
 sg13g2_or4_1 _26821_ (.A(net130),
    .B(net139),
    .C(net138),
    .D(net296),
    .X(_08090_));
 sg13g2_nand3b_1 _26822_ (.B(net1304),
    .C(_08090_),
    .Y(_08091_),
    .A_N(_08088_));
 sg13g2_nor2_1 _26823_ (.A(net99),
    .B(_08091_),
    .Y(_08092_));
 sg13g2_buf_1 _26824_ (.A(_08092_),
    .X(_08093_));
 sg13g2_nor3_1 _26825_ (.A(net130),
    .B(net296),
    .C(net117),
    .Y(_08094_));
 sg13g2_buf_2 _26826_ (.A(_08094_),
    .X(_08095_));
 sg13g2_nand2_1 _26827_ (.Y(_08096_),
    .A(net1302),
    .B(_08088_));
 sg13g2_nor2_1 _26828_ (.A(net99),
    .B(_08096_),
    .Y(_08097_));
 sg13g2_a221oi_1 _26829_ (.B2(net480),
    .C1(_08097_),
    .B1(_08095_),
    .A1(_07663_),
    .Y(_08098_),
    .A2(net99));
 sg13g2_nor2b_1 _26830_ (.A(net62),
    .B_N(_08098_),
    .Y(_08099_));
 sg13g2_a21oi_1 _26831_ (.A1(_08080_),
    .A2(net62),
    .Y(_02547_),
    .B1(_08099_));
 sg13g2_buf_1 _26832_ (.A(net1299),
    .X(_08100_));
 sg13g2_and2_1 _26833_ (.A(_07952_),
    .B(_07584_),
    .X(_08101_));
 sg13g2_buf_2 _26834_ (.A(_08101_),
    .X(_08102_));
 sg13g2_nand2_2 _26835_ (.Y(_08103_),
    .A(_08010_),
    .B(_08102_));
 sg13g2_nand3_1 _26836_ (.B(_08103_),
    .C(_08088_),
    .A(net1212),
    .Y(_08104_));
 sg13g2_buf_1 _26837_ (.A(net473),
    .X(_08105_));
 sg13g2_a22oi_1 _26838_ (.Y(_08106_),
    .B1(_08095_),
    .B2(net402),
    .A2(net99),
    .A1(net119));
 sg13g2_nand2_1 _26839_ (.Y(_08107_),
    .A(_08104_),
    .B(_08106_));
 sg13g2_mux2_1 _26840_ (.A0(_08107_),
    .A1(\stack[12][1] ),
    .S(net62),
    .X(_02548_));
 sg13g2_nand3_1 _26841_ (.B(_08103_),
    .C(_08088_),
    .A(net1217),
    .Y(_08108_));
 sg13g2_a22oi_1 _26842_ (.Y(_08109_),
    .B1(_08095_),
    .B2(net450),
    .A2(net99),
    .A1(net118));
 sg13g2_nand2_1 _26843_ (.Y(_08110_),
    .A(_08108_),
    .B(_08109_));
 sg13g2_mux2_1 _26844_ (.A0(_08110_),
    .A1(\stack[12][2] ),
    .S(net62),
    .X(_02549_));
 sg13g2_buf_1 _26845_ (.A(net1300),
    .X(_08111_));
 sg13g2_nand3_1 _26846_ (.B(_08103_),
    .C(_08088_),
    .A(net1211),
    .Y(_08112_));
 sg13g2_a22oi_1 _26847_ (.Y(_08113_),
    .B1(_08095_),
    .B2(net510),
    .A2(net99),
    .A1(net103));
 sg13g2_nand2_1 _26848_ (.Y(_08114_),
    .A(_08112_),
    .B(_08113_));
 sg13g2_mux2_1 _26849_ (.A0(_08114_),
    .A1(\stack[12][3] ),
    .S(net62),
    .X(_02550_));
 sg13g2_buf_1 _26850_ (.A(_07823_),
    .X(_08115_));
 sg13g2_nor2b_1 _26851_ (.A(_08083_),
    .B_N(_08088_),
    .Y(_08116_));
 sg13g2_buf_1 _26852_ (.A(_10022_),
    .X(_08117_));
 sg13g2_a22oi_1 _26853_ (.Y(_08118_),
    .B1(_08116_),
    .B2(net1210),
    .A2(_08095_),
    .A1(net493));
 sg13g2_o21ai_1 _26854_ (.B1(_08118_),
    .Y(_08119_),
    .A1(net98),
    .A2(_08103_));
 sg13g2_mux2_1 _26855_ (.A0(_08119_),
    .A1(\stack[12][4] ),
    .S(_08093_),
    .X(_02551_));
 sg13g2_inv_1 _26856_ (.Y(_08120_),
    .A(\stack[12][5] ));
 sg13g2_buf_1 _26857_ (.A(net471),
    .X(_08121_));
 sg13g2_a21oi_1 _26858_ (.A1(net1298),
    .A2(_08088_),
    .Y(_08122_),
    .B1(net99));
 sg13g2_nand2_1 _26859_ (.Y(_08123_),
    .A(_08091_),
    .B(_08122_));
 sg13g2_a21oi_1 _26860_ (.A1(net401),
    .A2(_08095_),
    .Y(_08124_),
    .B1(_08123_));
 sg13g2_a221oi_1 _26861_ (.B2(_08120_),
    .C1(_08124_),
    .B1(net62),
    .A1(net89),
    .Y(_02552_),
    .A2(_08083_));
 sg13g2_inv_1 _26862_ (.Y(_08125_),
    .A(\stack[12][6] ));
 sg13g2_nand2_1 _26863_ (.Y(_08126_),
    .A(net42),
    .B(net99));
 sg13g2_a221oi_1 _26864_ (.B2(net879),
    .C1(net62),
    .B1(_08116_),
    .A1(net449),
    .Y(_08127_),
    .A2(_08095_));
 sg13g2_a22oi_1 _26865_ (.Y(_02553_),
    .B1(_08126_),
    .B2(_08127_),
    .A2(net62),
    .A1(_08125_));
 sg13g2_and2_1 _26866_ (.A(net1219),
    .B(_08116_),
    .X(_08128_));
 sg13g2_a221oi_1 _26867_ (.B2(\stack[12][7] ),
    .C1(_08128_),
    .B1(_08093_),
    .A1(net298),
    .Y(_08129_),
    .A2(_08095_));
 sg13g2_o21ai_1 _26868_ (.B1(_08129_),
    .Y(_02554_),
    .A1(net45),
    .A2(_08103_));
 sg13g2_or4_1 _26869_ (.A(_07604_),
    .B(net143),
    .C(net142),
    .D(net297),
    .X(_08130_));
 sg13g2_buf_2 _26870_ (.A(_08130_),
    .X(_08131_));
 sg13g2_nand2_1 _26871_ (.Y(_08132_),
    .A(net573),
    .B(_07598_));
 sg13g2_buf_1 _26872_ (.A(_08132_),
    .X(_08133_));
 sg13g2_nor2_1 _26873_ (.A(_08086_),
    .B(net522),
    .Y(_08134_));
 sg13g2_buf_1 _26874_ (.A(_08134_),
    .X(_08135_));
 sg13g2_nand2_1 _26875_ (.Y(_08136_),
    .A(net1302),
    .B(net507));
 sg13g2_nor3_1 _26876_ (.A(net130),
    .B(_07968_),
    .C(net126),
    .Y(_08137_));
 sg13g2_buf_2 _26877_ (.A(_08137_),
    .X(_08138_));
 sg13g2_mux2_1 _26878_ (.A0(_08136_),
    .A1(_08023_),
    .S(_08138_),
    .X(_08139_));
 sg13g2_o21ai_1 _26879_ (.B1(_08139_),
    .Y(_08140_),
    .A1(net487),
    .A2(_08131_));
 sg13g2_buf_8 _26880_ (.A(_08138_),
    .X(_08141_));
 sg13g2_nand3b_1 _26881_ (.B(_08131_),
    .C(net1276),
    .Y(_08142_),
    .A_N(_08134_));
 sg13g2_buf_1 _26882_ (.A(_08142_),
    .X(_08143_));
 sg13g2_nor2_2 _26883_ (.A(net87),
    .B(_08143_),
    .Y(_08144_));
 sg13g2_mux2_1 _26884_ (.A0(_08140_),
    .A1(\stack[13][0] ),
    .S(_08144_),
    .X(_02555_));
 sg13g2_nor2b_1 _26885_ (.A(net119),
    .B_N(_08138_),
    .Y(_08145_));
 sg13g2_a21oi_1 _26886_ (.A1(net1225),
    .A2(net507),
    .Y(_08146_),
    .B1(net87));
 sg13g2_inv_1 _26887_ (.Y(_08147_),
    .A(_08131_));
 sg13g2_nand2_1 _26888_ (.Y(_08148_),
    .A(net402),
    .B(_08147_));
 sg13g2_o21ai_1 _26889_ (.B1(_08148_),
    .Y(_08149_),
    .A1(_08145_),
    .A2(_08146_));
 sg13g2_mux2_1 _26890_ (.A0(_08149_),
    .A1(\stack[13][1] ),
    .S(_08144_),
    .X(_02556_));
 sg13g2_nor2b_1 _26891_ (.A(net118),
    .B_N(_08138_),
    .Y(_08150_));
 sg13g2_a21oi_1 _26892_ (.A1(net1224),
    .A2(net507),
    .Y(_08151_),
    .B1(net87));
 sg13g2_nand2_1 _26893_ (.Y(_08152_),
    .A(net450),
    .B(_08147_));
 sg13g2_o21ai_1 _26894_ (.B1(_08152_),
    .Y(_08153_),
    .A1(_08150_),
    .A2(_08151_));
 sg13g2_mux2_1 _26895_ (.A0(_08153_),
    .A1(\stack[13][2] ),
    .S(_08144_),
    .X(_02557_));
 sg13g2_nor2b_1 _26896_ (.A(net103),
    .B_N(_08138_),
    .Y(_08154_));
 sg13g2_a21oi_1 _26897_ (.A1(net1223),
    .A2(net507),
    .Y(_08155_),
    .B1(_08138_));
 sg13g2_nand2_1 _26898_ (.Y(_08156_),
    .A(net494),
    .B(_08147_));
 sg13g2_o21ai_1 _26899_ (.B1(_08156_),
    .Y(_08157_),
    .A1(_08154_),
    .A2(_08155_));
 sg13g2_mux2_1 _26900_ (.A0(_08157_),
    .A1(\stack[13][3] ),
    .S(_08144_),
    .X(_02558_));
 sg13g2_buf_1 _26901_ (.A(_10022_),
    .X(_08158_));
 sg13g2_and2_1 _26902_ (.A(net1273),
    .B(_08131_),
    .X(_08159_));
 sg13g2_nor2b_1 _26903_ (.A(_08135_),
    .B_N(\stack[13][4] ),
    .Y(_08160_));
 sg13g2_a221oi_1 _26904_ (.B2(_08160_),
    .C1(net87),
    .B1(_08159_),
    .A1(net1209),
    .Y(_08161_),
    .A2(net507));
 sg13g2_a21o_1 _26905_ (.A2(net87),
    .A1(net98),
    .B1(_08161_),
    .X(_08162_));
 sg13g2_o21ai_1 _26906_ (.B1(_08162_),
    .Y(_02559_),
    .A1(net496),
    .A2(_08131_));
 sg13g2_nand2_1 _26907_ (.Y(_08163_),
    .A(net1221),
    .B(net507));
 sg13g2_o21ai_1 _26908_ (.B1(_08163_),
    .Y(_08164_),
    .A1(net446),
    .A2(_08131_));
 sg13g2_inv_1 _26909_ (.Y(_08165_),
    .A(\stack[13][5] ));
 sg13g2_nor2_1 _26910_ (.A(_08165_),
    .B(_08143_),
    .Y(_08166_));
 sg13g2_nor3_1 _26911_ (.A(_08141_),
    .B(_08164_),
    .C(_08166_),
    .Y(_08167_));
 sg13g2_a21oi_1 _26912_ (.A1(net89),
    .A2(net87),
    .Y(_02560_),
    .B1(_08167_));
 sg13g2_and2_1 _26913_ (.A(_07893_),
    .B(_07897_),
    .X(_08168_));
 sg13g2_buf_1 _26914_ (.A(_08168_),
    .X(_08169_));
 sg13g2_nand3_1 _26915_ (.B(_08169_),
    .C(net87),
    .A(_07868_),
    .Y(_08170_));
 sg13g2_inv_1 _26916_ (.Y(_08171_),
    .A(_08138_));
 sg13g2_nand2_1 _26917_ (.Y(_08172_),
    .A(net451),
    .B(_08147_));
 sg13g2_nand2_1 _26918_ (.Y(_08173_),
    .A(net1220),
    .B(net507));
 sg13g2_nand4_1 _26919_ (.B(_08143_),
    .C(_08172_),
    .A(_08171_),
    .Y(_08174_),
    .D(_08173_));
 sg13g2_or3_1 _26920_ (.A(\stack[13][6] ),
    .B(_08141_),
    .C(_08143_),
    .X(_08175_));
 sg13g2_and3_1 _26921_ (.X(_02561_),
    .A(_08170_),
    .B(_08174_),
    .C(_08175_));
 sg13g2_a22oi_1 _26922_ (.Y(_08176_),
    .B1(_08147_),
    .B2(net445),
    .A2(_08135_),
    .A1(net1219));
 sg13g2_nand3b_1 _26923_ (.B(_08159_),
    .C(\stack[13][7] ),
    .Y(_08177_),
    .A_N(net507));
 sg13g2_a21o_1 _26924_ (.A2(_08177_),
    .A1(_08176_),
    .B1(net87),
    .X(_08178_));
 sg13g2_o21ai_1 _26925_ (.B1(_08178_),
    .Y(_02562_),
    .A1(net45),
    .A2(_08171_));
 sg13g2_nand2_1 _26926_ (.Y(_08179_),
    .A(_07938_),
    .B(_08010_));
 sg13g2_a22oi_1 _26927_ (.Y(_08180_),
    .B1(_07496_),
    .B2(_07501_),
    .A2(_07528_),
    .A1(_07516_));
 sg13g2_buf_2 _26928_ (.A(_08180_),
    .X(_08181_));
 sg13g2_buf_8 _26929_ (.A(_08181_),
    .X(_08182_));
 sg13g2_buf_1 _26930_ (.A(_07943_),
    .X(_08183_));
 sg13g2_o21ai_1 _26931_ (.B1(_09906_),
    .Y(_08184_),
    .A1(net532),
    .A2(_08086_));
 sg13g2_a21oi_1 _26932_ (.A1(_07622_),
    .A2(net124),
    .Y(_08185_),
    .B1(_08184_));
 sg13g2_buf_2 _26933_ (.A(_08185_),
    .X(_08186_));
 sg13g2_nand2_1 _26934_ (.Y(_08187_),
    .A(_08179_),
    .B(_08186_));
 sg13g2_buf_2 _26935_ (.A(_08187_),
    .X(_08188_));
 sg13g2_and2_1 _26936_ (.A(_07938_),
    .B(_08010_),
    .X(_08189_));
 sg13g2_buf_1 _26937_ (.A(_08189_),
    .X(_08190_));
 sg13g2_nand2_1 _26938_ (.Y(_08191_),
    .A(net140),
    .B(_07502_));
 sg13g2_buf_1 _26939_ (.A(_08191_),
    .X(_08192_));
 sg13g2_nor4_1 _26940_ (.A(_07748_),
    .B(net491),
    .C(_07754_),
    .D(net116),
    .Y(_08193_));
 sg13g2_buf_2 _26941_ (.A(_08193_),
    .X(_08194_));
 sg13g2_nor2_1 _26942_ (.A(net532),
    .B(_08086_),
    .Y(_08195_));
 sg13g2_buf_2 _26943_ (.A(_08195_),
    .X(_08196_));
 sg13g2_and3_1 _26944_ (.X(_08197_),
    .A(net1218),
    .B(_08179_),
    .C(_08196_));
 sg13g2_a221oi_1 _26945_ (.B2(net478),
    .C1(_08197_),
    .B1(_08194_),
    .A1(net134),
    .Y(_08198_),
    .A2(_08190_));
 sg13g2_nor2_1 _26946_ (.A(\stack[14][0] ),
    .B(_08188_),
    .Y(_08199_));
 sg13g2_a21oi_1 _26947_ (.A1(_08188_),
    .A2(_08198_),
    .Y(_02563_),
    .B1(_08199_));
 sg13g2_buf_1 _26948_ (.A(_08190_),
    .X(_08200_));
 sg13g2_nand2_1 _26949_ (.Y(_08201_),
    .A(net1225),
    .B(_08196_));
 sg13g2_a22oi_1 _26950_ (.Y(_08202_),
    .B1(_08194_),
    .B2(net473),
    .A2(_08190_),
    .A1(net119));
 sg13g2_o21ai_1 _26951_ (.B1(_08202_),
    .Y(_08203_),
    .A1(net61),
    .A2(_08201_));
 sg13g2_mux2_1 _26952_ (.A0(\stack[14][1] ),
    .A1(_08203_),
    .S(_08188_),
    .X(_02564_));
 sg13g2_nand2_1 _26953_ (.Y(_08204_),
    .A(net1224),
    .B(_08196_));
 sg13g2_a22oi_1 _26954_ (.Y(_08205_),
    .B1(_08194_),
    .B2(net450),
    .A2(_08190_),
    .A1(net118));
 sg13g2_o21ai_1 _26955_ (.B1(_08205_),
    .Y(_08206_),
    .A1(net61),
    .A2(_08204_));
 sg13g2_mux2_1 _26956_ (.A0(\stack[14][2] ),
    .A1(_08206_),
    .S(_08188_),
    .X(_02565_));
 sg13g2_nand2_1 _26957_ (.Y(_08207_),
    .A(net1211),
    .B(_08196_));
 sg13g2_a22oi_1 _26958_ (.Y(_08208_),
    .B1(_08194_),
    .B2(net510),
    .A2(_08190_),
    .A1(net103));
 sg13g2_o21ai_1 _26959_ (.B1(_08208_),
    .Y(_08209_),
    .A1(_08190_),
    .A2(_08207_));
 sg13g2_mux2_1 _26960_ (.A0(\stack[14][3] ),
    .A1(_08209_),
    .S(_08188_),
    .X(_02566_));
 sg13g2_nor2_1 _26961_ (.A(\stack[14][4] ),
    .B(net61),
    .Y(_08210_));
 sg13g2_a21o_1 _26962_ (.A2(_08194_),
    .A1(net493),
    .B1(_08186_),
    .X(_08211_));
 sg13g2_a221oi_1 _26963_ (.B2(net1222),
    .C1(_08211_),
    .B1(_08196_),
    .A1(_07938_),
    .Y(_08212_),
    .A2(_08010_));
 sg13g2_a221oi_1 _26964_ (.B2(_08210_),
    .C1(_08212_),
    .B1(_08186_),
    .A1(net100),
    .Y(_02567_),
    .A2(net61));
 sg13g2_a21oi_1 _26965_ (.A1(net1216),
    .A2(_08196_),
    .Y(_08213_),
    .B1(_08186_));
 sg13g2_a21oi_1 _26966_ (.A1(net401),
    .A2(_08194_),
    .Y(_08214_),
    .B1(_08200_));
 sg13g2_nor2_1 _26967_ (.A(\stack[14][5] ),
    .B(_08188_),
    .Y(_08215_));
 sg13g2_a221oi_1 _26968_ (.B2(_08214_),
    .C1(_08215_),
    .B1(_08213_),
    .A1(net88),
    .Y(_02568_),
    .A2(net61));
 sg13g2_a21oi_1 _26969_ (.A1(net879),
    .A2(_08196_),
    .Y(_08216_),
    .B1(_08186_));
 sg13g2_a21oi_1 _26970_ (.A1(net449),
    .A2(_08194_),
    .Y(_08217_),
    .B1(_08200_));
 sg13g2_nor2_1 _26971_ (.A(\stack[14][6] ),
    .B(_08188_),
    .Y(_08218_));
 sg13g2_a221oi_1 _26972_ (.B2(_08217_),
    .C1(_08218_),
    .B1(_08216_),
    .A1(_07997_),
    .Y(_02569_),
    .A2(net61));
 sg13g2_nand2_1 _26973_ (.Y(_08219_),
    .A(\stack[14][7] ),
    .B(_08186_));
 sg13g2_a221oi_1 _26974_ (.B2(net298),
    .C1(net61),
    .B1(_08194_),
    .A1(net1215),
    .Y(_08220_),
    .A2(_08196_));
 sg13g2_a22oi_1 _26975_ (.Y(_02570_),
    .B1(_08219_),
    .B2(_08220_),
    .A2(net61),
    .A1(net45));
 sg13g2_inv_1 _26976_ (.Y(_08221_),
    .A(\stack[15][0] ));
 sg13g2_nor4_1 _26977_ (.A(_07606_),
    .B(_07609_),
    .C(_08025_),
    .D(_08026_),
    .Y(_08222_));
 sg13g2_buf_2 _26978_ (.A(_08222_),
    .X(_08223_));
 sg13g2_and2_1 _26979_ (.A(net124),
    .B(_08223_),
    .X(_08224_));
 sg13g2_buf_2 _26980_ (.A(_08224_),
    .X(_08225_));
 sg13g2_nor2_1 _26981_ (.A(_08016_),
    .B(_08086_),
    .Y(_08226_));
 sg13g2_buf_2 _26982_ (.A(_08226_),
    .X(_08227_));
 sg13g2_nand4_1 _26983_ (.B(net142),
    .C(net404),
    .A(net143),
    .Y(_08228_),
    .D(net124));
 sg13g2_nand3b_1 _26984_ (.B(_08228_),
    .C(net1304),
    .Y(_08229_),
    .A_N(_08227_));
 sg13g2_buf_1 _26985_ (.A(_08229_),
    .X(_08230_));
 sg13g2_nor2_1 _26986_ (.A(_08225_),
    .B(_08230_),
    .Y(_08231_));
 sg13g2_buf_2 _26987_ (.A(_08231_),
    .X(_08232_));
 sg13g2_nor3_1 _26988_ (.A(_07748_),
    .B(net297),
    .C(net116),
    .Y(_08233_));
 sg13g2_buf_2 _26989_ (.A(_08233_),
    .X(_08234_));
 sg13g2_buf_1 _26990_ (.A(_08023_),
    .X(_08235_));
 sg13g2_buf_8 _26991_ (.A(_08225_),
    .X(_08236_));
 sg13g2_nand2_1 _26992_ (.Y(_08237_),
    .A(net123),
    .B(net86));
 sg13g2_buf_1 _26993_ (.A(net1302),
    .X(_08238_));
 sg13g2_a21o_1 _26994_ (.A2(_08227_),
    .A1(net1208),
    .B1(_08225_),
    .X(_08239_));
 sg13g2_a221oi_1 _26995_ (.B2(_08239_),
    .C1(_08232_),
    .B1(_08237_),
    .A1(net478),
    .Y(_08240_),
    .A2(_08234_));
 sg13g2_a21oi_1 _26996_ (.A1(_08221_),
    .A2(_08232_),
    .Y(_02571_),
    .B1(_08240_));
 sg13g2_inv_1 _26997_ (.Y(_08241_),
    .A(\stack[15][1] ));
 sg13g2_nand2b_1 _26998_ (.Y(_08242_),
    .B(net86),
    .A_N(_07700_));
 sg13g2_a21o_1 _26999_ (.A2(_08227_),
    .A1(net1299),
    .B1(_08225_),
    .X(_08243_));
 sg13g2_a221oi_1 _27000_ (.B2(_08243_),
    .C1(_08232_),
    .B1(_08242_),
    .A1(net447),
    .Y(_08244_),
    .A2(_08234_));
 sg13g2_a21oi_1 _27001_ (.A1(_08241_),
    .A2(_08232_),
    .Y(_02572_),
    .B1(_08244_));
 sg13g2_nand2b_1 _27002_ (.Y(_08245_),
    .B(net86),
    .A_N(_07738_));
 sg13g2_a21o_1 _27003_ (.A2(_08227_),
    .A1(net1301),
    .B1(_08225_),
    .X(_08246_));
 sg13g2_a221oi_1 _27004_ (.B2(_08246_),
    .C1(_08232_),
    .B1(_08245_),
    .A1(net452),
    .Y(_08247_),
    .A2(_08234_));
 sg13g2_a21oi_1 _27005_ (.A1(_07246_),
    .A2(_08232_),
    .Y(_02573_),
    .B1(_08247_));
 sg13g2_inv_1 _27006_ (.Y(_08248_),
    .A(\stack[15][3] ));
 sg13g2_nand2b_1 _27007_ (.Y(_08249_),
    .B(_08225_),
    .A_N(_07783_));
 sg13g2_a21o_1 _27008_ (.A2(_08227_),
    .A1(net1300),
    .B1(_08225_),
    .X(_08250_));
 sg13g2_a221oi_1 _27009_ (.B2(_08250_),
    .C1(_08232_),
    .B1(_08249_),
    .A1(net492),
    .Y(_08251_),
    .A2(_08234_));
 sg13g2_a21oi_1 _27010_ (.A1(_08248_),
    .A2(_08232_),
    .Y(_02574_),
    .B1(_08251_));
 sg13g2_inv_2 _27011_ (.Y(_08252_),
    .A(_10022_));
 sg13g2_nor3_1 _27012_ (.A(_08252_),
    .B(net516),
    .C(_08086_),
    .Y(_08253_));
 sg13g2_nand2_2 _27013_ (.Y(_08254_),
    .A(net124),
    .B(_08223_));
 sg13g2_a22oi_1 _27014_ (.Y(_08255_),
    .B1(_08253_),
    .B2(_08254_),
    .A2(_08234_),
    .A1(net484));
 sg13g2_inv_1 _27015_ (.Y(_08256_),
    .A(_08230_));
 sg13g2_nor2_1 _27016_ (.A(net86),
    .B(_08256_),
    .Y(_08257_));
 sg13g2_nor3_1 _27017_ (.A(\stack[15][4] ),
    .B(_08236_),
    .C(_08230_),
    .Y(_08258_));
 sg13g2_a221oi_1 _27018_ (.B2(_08257_),
    .C1(_08258_),
    .B1(_08255_),
    .A1(net100),
    .Y(_02575_),
    .A2(net86));
 sg13g2_and2_1 _27019_ (.A(net90),
    .B(net86),
    .X(_08259_));
 sg13g2_a221oi_1 _27020_ (.B2(\stack[15][5] ),
    .C1(net86),
    .B1(_08256_),
    .A1(net1216),
    .Y(_08260_),
    .A2(_08227_));
 sg13g2_nand2_1 _27021_ (.Y(_08261_),
    .A(net403),
    .B(_08234_));
 sg13g2_o21ai_1 _27022_ (.B1(_08261_),
    .Y(_02576_),
    .A1(_08259_),
    .A2(_08260_));
 sg13g2_and2_1 _27023_ (.A(_07866_),
    .B(_07867_),
    .X(_08262_));
 sg13g2_buf_1 _27024_ (.A(_08262_),
    .X(_08263_));
 sg13g2_nor2_1 _27025_ (.A(_08263_),
    .B(_08254_),
    .Y(_08264_));
 sg13g2_nor4_1 _27026_ (.A(_10018_),
    .B(net516),
    .C(_08086_),
    .D(_08225_),
    .Y(_08265_));
 sg13g2_a221oi_1 _27027_ (.B2(net451),
    .C1(_08265_),
    .B1(_08234_),
    .A1(_08263_),
    .Y(_08266_),
    .A2(net86));
 sg13g2_nor3_1 _27028_ (.A(\stack[15][6] ),
    .B(_08236_),
    .C(_08230_),
    .Y(_08267_));
 sg13g2_a221oi_1 _27029_ (.B2(_08257_),
    .C1(_08267_),
    .B1(_08266_),
    .A1(_08169_),
    .Y(_02577_),
    .A2(_08264_));
 sg13g2_nand3_1 _27030_ (.B(\stack[15][7] ),
    .C(_08228_),
    .A(net1192),
    .Y(_08268_));
 sg13g2_nand2_1 _27031_ (.Y(_08269_),
    .A(net1213),
    .B(_08227_));
 sg13g2_o21ai_1 _27032_ (.B1(_08269_),
    .Y(_08270_),
    .A1(_08227_),
    .A2(_08268_));
 sg13g2_a22oi_1 _27033_ (.Y(_08271_),
    .B1(_08270_),
    .B2(_08254_),
    .A2(_08234_),
    .A1(net298));
 sg13g2_o21ai_1 _27034_ (.B1(_08271_),
    .Y(_02578_),
    .A1(net41),
    .A2(_08254_));
 sg13g2_nor2_1 _27035_ (.A(_07587_),
    .B(net116),
    .Y(_08272_));
 sg13g2_buf_2 _27036_ (.A(_08272_),
    .X(_08273_));
 sg13g2_buf_1 _27037_ (.A(_08273_),
    .X(_08274_));
 sg13g2_nand2_2 _27038_ (.Y(_08275_),
    .A(_07475_),
    .B(_07592_));
 sg13g2_nor2_1 _27039_ (.A(_07600_),
    .B(_08275_),
    .Y(_08276_));
 sg13g2_buf_2 _27040_ (.A(_08276_),
    .X(_08277_));
 sg13g2_nor2_1 _27041_ (.A(_10144_),
    .B(_08277_),
    .Y(_08278_));
 sg13g2_a221oi_1 _27042_ (.B2(net531),
    .C1(_07525_),
    .B1(_07520_),
    .A1(_07387_),
    .Y(_08279_),
    .A2(net406));
 sg13g2_a221oi_1 _27043_ (.B2(_07501_),
    .C1(_08279_),
    .B1(_07496_),
    .A1(_07514_),
    .Y(_08280_),
    .A2(_07579_));
 sg13g2_buf_1 _27044_ (.A(_08280_),
    .X(_08281_));
 sg13g2_nand4_1 _27045_ (.B(net138),
    .C(net299),
    .A(net139),
    .Y(_08282_),
    .D(net133));
 sg13g2_buf_1 _27046_ (.A(_08282_),
    .X(_08283_));
 sg13g2_and2_1 _27047_ (.A(_08278_),
    .B(_08283_),
    .X(_08284_));
 sg13g2_buf_2 _27048_ (.A(_08284_),
    .X(_08285_));
 sg13g2_a22oi_1 _27049_ (.Y(_08286_),
    .B1(_08285_),
    .B2(\stack[16][0] ),
    .A2(_08277_),
    .A1(net1226));
 sg13g2_nand2b_1 _27050_ (.Y(_08287_),
    .B(net141),
    .A_N(net140));
 sg13g2_buf_2 _27051_ (.A(_08287_),
    .X(_08288_));
 sg13g2_buf_8 _27052_ (.A(_08288_),
    .X(_08289_));
 sg13g2_nor4_1 _27053_ (.A(_07748_),
    .B(net491),
    .C(net129),
    .D(net97),
    .Y(_08290_));
 sg13g2_buf_2 _27054_ (.A(_08290_),
    .X(_08291_));
 sg13g2_a22oi_1 _27055_ (.Y(_08292_),
    .B1(_08291_),
    .B2(net453),
    .A2(net60),
    .A1(net131));
 sg13g2_o21ai_1 _27056_ (.B1(_08292_),
    .Y(_02579_),
    .A1(net60),
    .A2(_08286_));
 sg13g2_a22oi_1 _27057_ (.Y(_08293_),
    .B1(_08285_),
    .B2(\stack[16][1] ),
    .A2(_08277_),
    .A1(net883));
 sg13g2_buf_1 _27058_ (.A(_08105_),
    .X(_08294_));
 sg13g2_a22oi_1 _27059_ (.Y(_08295_),
    .B1(_08291_),
    .B2(_08294_),
    .A2(net60),
    .A1(net105));
 sg13g2_o21ai_1 _27060_ (.B1(_08295_),
    .Y(_02580_),
    .A1(net60),
    .A2(_08293_));
 sg13g2_a22oi_1 _27061_ (.Y(_08296_),
    .B1(_08285_),
    .B2(\stack[16][2] ),
    .A2(_08277_),
    .A1(net882));
 sg13g2_buf_1 _27062_ (.A(net450),
    .X(_08297_));
 sg13g2_a22oi_1 _27063_ (.Y(_08298_),
    .B1(_08291_),
    .B2(_08297_),
    .A2(_08273_),
    .A1(net104));
 sg13g2_o21ai_1 _27064_ (.B1(_08298_),
    .Y(_02581_),
    .A1(net60),
    .A2(_08296_));
 sg13g2_a22oi_1 _27065_ (.Y(_08299_),
    .B1(_08285_),
    .B2(\stack[16][3] ),
    .A2(_08277_),
    .A1(net881));
 sg13g2_buf_1 _27066_ (.A(_10178_),
    .X(_08300_));
 sg13g2_a22oi_1 _27067_ (.Y(_08301_),
    .B1(_08291_),
    .B2(net477),
    .A2(_08273_),
    .A1(net91));
 sg13g2_o21ai_1 _27068_ (.B1(_08301_),
    .Y(_02582_),
    .A1(net60),
    .A2(_08299_));
 sg13g2_buf_1 _27069_ (.A(_07600_),
    .X(_08302_));
 sg13g2_nor3_1 _27070_ (.A(_08252_),
    .B(net521),
    .C(_08275_),
    .Y(_08303_));
 sg13g2_nor4_1 _27071_ (.A(net496),
    .B(_07748_),
    .C(net296),
    .D(net97),
    .Y(_08304_));
 sg13g2_and2_1 _27072_ (.A(\stack[16][4] ),
    .B(_08285_),
    .X(_08305_));
 sg13g2_nor4_1 _27073_ (.A(_08273_),
    .B(_08303_),
    .C(_08304_),
    .D(_08305_),
    .Y(_08306_));
 sg13g2_a21oi_1 _27074_ (.A1(_07985_),
    .A2(net60),
    .Y(_02583_),
    .B1(_08306_));
 sg13g2_a221oi_1 _27075_ (.B2(\stack[16][5] ),
    .C1(_08273_),
    .B1(_08285_),
    .A1(_07850_),
    .Y(_08307_),
    .A2(_08277_));
 sg13g2_a21o_1 _27076_ (.A2(_08273_),
    .A1(net90),
    .B1(_08307_),
    .X(_08308_));
 sg13g2_o21ai_1 _27077_ (.B1(_08308_),
    .Y(_02584_),
    .A1(net446),
    .A2(_08283_));
 sg13g2_a22oi_1 _27078_ (.Y(_08309_),
    .B1(_08285_),
    .B2(\stack[16][6] ),
    .A2(_08277_),
    .A1(net880));
 sg13g2_a22oi_1 _27079_ (.Y(_08310_),
    .B1(_08291_),
    .B2(net405),
    .A2(_08273_),
    .A1(net46));
 sg13g2_o21ai_1 _27080_ (.B1(_08310_),
    .Y(_02585_),
    .A1(net60),
    .A2(_08309_));
 sg13g2_nor2_1 _27081_ (.A(_10138_),
    .B(_08283_),
    .Y(_08311_));
 sg13g2_a221oi_1 _27082_ (.B2(\stack[16][7] ),
    .C1(_08311_),
    .B1(_08285_),
    .A1(_07930_),
    .Y(_08312_),
    .A2(_08277_));
 sg13g2_nor2b_1 _27083_ (.A(_08274_),
    .B_N(_08312_),
    .Y(_08313_));
 sg13g2_a21oi_1 _27084_ (.A1(net43),
    .A2(_08274_),
    .Y(_02586_),
    .B1(_08313_));
 sg13g2_and2_1 _27085_ (.A(_08223_),
    .B(net133),
    .X(_08314_));
 sg13g2_buf_2 _27086_ (.A(_08314_),
    .X(_08315_));
 sg13g2_buf_1 _27087_ (.A(_08315_),
    .X(_08316_));
 sg13g2_nor2_1 _27088_ (.A(net522),
    .B(_08275_),
    .Y(_08317_));
 sg13g2_buf_1 _27089_ (.A(_08317_),
    .X(_08318_));
 sg13g2_buf_1 _27090_ (.A(_08318_),
    .X(_08319_));
 sg13g2_nand4_1 _27091_ (.B(net138),
    .C(net404),
    .A(net139),
    .Y(_08320_),
    .D(net133));
 sg13g2_and2_1 _27092_ (.A(_09908_),
    .B(_08320_),
    .X(_08321_));
 sg13g2_buf_2 _27093_ (.A(_08321_),
    .X(_08322_));
 sg13g2_nand3b_1 _27094_ (.B(_08322_),
    .C(\stack[17][0] ),
    .Y(_08323_),
    .A_N(net490));
 sg13g2_nor3_1 _27095_ (.A(_07748_),
    .B(_08036_),
    .C(net97),
    .Y(_08324_));
 sg13g2_buf_2 _27096_ (.A(_08324_),
    .X(_08325_));
 sg13g2_a221oi_1 _27097_ (.B2(net1226),
    .C1(_08315_),
    .B1(net490),
    .A1(_07960_),
    .Y(_08326_),
    .A2(_08325_));
 sg13g2_a22oi_1 _27098_ (.Y(_02587_),
    .B1(_08323_),
    .B2(_08326_),
    .A2(_08316_),
    .A1(net123));
 sg13g2_nor2b_1 _27099_ (.A(net490),
    .B_N(\stack[17][1] ),
    .Y(_08327_));
 sg13g2_a22oi_1 _27100_ (.Y(_08328_),
    .B1(_08327_),
    .B2(_08322_),
    .A2(net490),
    .A1(net883));
 sg13g2_a22oi_1 _27101_ (.Y(_08329_),
    .B1(net85),
    .B2(net105),
    .A2(_08325_),
    .A1(net447));
 sg13g2_o21ai_1 _27102_ (.B1(_08329_),
    .Y(_02588_),
    .A1(net85),
    .A2(_08328_));
 sg13g2_nor2b_1 _27103_ (.A(net490),
    .B_N(\stack[17][2] ),
    .Y(_08330_));
 sg13g2_a22oi_1 _27104_ (.Y(_08331_),
    .B1(_08330_),
    .B2(_08322_),
    .A2(net490),
    .A1(net882));
 sg13g2_a22oi_1 _27105_ (.Y(_08332_),
    .B1(net85),
    .B2(net104),
    .A2(_08325_),
    .A1(net452));
 sg13g2_o21ai_1 _27106_ (.B1(_08332_),
    .Y(_02589_),
    .A1(_08316_),
    .A2(_08331_));
 sg13g2_nor2b_1 _27107_ (.A(_08318_),
    .B_N(\stack[17][3] ),
    .Y(_08333_));
 sg13g2_a22oi_1 _27108_ (.Y(_08334_),
    .B1(_08333_),
    .B2(_08322_),
    .A2(net490),
    .A1(net881));
 sg13g2_a22oi_1 _27109_ (.Y(_08335_),
    .B1(net85),
    .B2(net91),
    .A2(_08325_),
    .A1(net492));
 sg13g2_o21ai_1 _27110_ (.B1(_08335_),
    .Y(_02590_),
    .A1(net85),
    .A2(_08334_));
 sg13g2_buf_1 _27111_ (.A(_10190_),
    .X(_08336_));
 sg13g2_nor2b_1 _27112_ (.A(_08318_),
    .B_N(\stack[17][4] ),
    .Y(_08337_));
 sg13g2_a221oi_1 _27113_ (.B2(_08322_),
    .C1(_08315_),
    .B1(_08337_),
    .A1(net1210),
    .Y(_08338_),
    .A2(_08318_));
 sg13g2_a21oi_1 _27114_ (.A1(net102),
    .A2(_08315_),
    .Y(_08339_),
    .B1(_08338_));
 sg13g2_a21o_1 _27115_ (.A2(_08325_),
    .A1(net476),
    .B1(_08339_),
    .X(_02591_));
 sg13g2_nor2b_1 _27116_ (.A(_08318_),
    .B_N(\stack[17][5] ),
    .Y(_08340_));
 sg13g2_a221oi_1 _27117_ (.B2(_08322_),
    .C1(_08315_),
    .B1(_08340_),
    .A1(net1214),
    .Y(_08341_),
    .A2(_08318_));
 sg13g2_a21oi_1 _27118_ (.A1(net88),
    .A2(_08315_),
    .Y(_08342_),
    .B1(_08341_));
 sg13g2_a21o_1 _27119_ (.A2(_08325_),
    .A1(net403),
    .B1(_08342_),
    .X(_02592_));
 sg13g2_nor2b_1 _27120_ (.A(_08318_),
    .B_N(\stack[17][6] ),
    .Y(_08343_));
 sg13g2_a22oi_1 _27121_ (.Y(_08344_),
    .B1(_08343_),
    .B2(_08322_),
    .A2(_08319_),
    .A1(net880));
 sg13g2_a22oi_1 _27122_ (.Y(_08345_),
    .B1(net85),
    .B2(net42),
    .A2(_08325_),
    .A1(net405));
 sg13g2_o21ai_1 _27123_ (.B1(_08345_),
    .Y(_02593_),
    .A1(net85),
    .A2(_08344_));
 sg13g2_nand3b_1 _27124_ (.B(_08322_),
    .C(\stack[17][7] ),
    .Y(_08346_),
    .A_N(net490));
 sg13g2_buf_1 _27125_ (.A(net445),
    .X(_08347_));
 sg13g2_a221oi_1 _27126_ (.B2(net1215),
    .C1(_08315_),
    .B1(_08319_),
    .A1(net294),
    .Y(_08348_),
    .A2(_08325_));
 sg13g2_a22oi_1 _27127_ (.Y(_02594_),
    .B1(_08346_),
    .B2(_08348_),
    .A2(net85),
    .A1(net45));
 sg13g2_nand4_1 _27128_ (.B(_07559_),
    .C(net299),
    .A(net128),
    .Y(_08349_),
    .D(net124));
 sg13g2_nor2_1 _27129_ (.A(_07587_),
    .B(_08289_),
    .Y(_08350_));
 sg13g2_buf_1 _27130_ (.A(_08350_),
    .X(_08351_));
 sg13g2_nor2_1 _27131_ (.A(net532),
    .B(_08275_),
    .Y(_08352_));
 sg13g2_buf_1 _27132_ (.A(_08352_),
    .X(_08353_));
 sg13g2_nor2_1 _27133_ (.A(_10143_),
    .B(net515),
    .Y(_08354_));
 sg13g2_and2_1 _27134_ (.A(_08349_),
    .B(_08354_),
    .X(_08355_));
 sg13g2_buf_2 _27135_ (.A(_08355_),
    .X(_08356_));
 sg13g2_a221oi_1 _27136_ (.B2(\stack[18][0] ),
    .C1(_08350_),
    .B1(_08356_),
    .A1(net1208),
    .Y(_08357_),
    .A2(net515));
 sg13g2_a21o_1 _27137_ (.A2(net59),
    .A1(net123),
    .B1(_08357_),
    .X(_08358_));
 sg13g2_o21ai_1 _27138_ (.B1(_08358_),
    .Y(_02595_),
    .A1(net487),
    .A2(_08349_));
 sg13g2_nand2_1 _27139_ (.Y(_08359_),
    .A(_07606_),
    .B(net142));
 sg13g2_buf_1 _27140_ (.A(_08359_),
    .X(_08360_));
 sg13g2_nor3_1 _27141_ (.A(_08089_),
    .B(net116),
    .C(net122),
    .Y(_08361_));
 sg13g2_buf_2 _27142_ (.A(_08361_),
    .X(_08362_));
 sg13g2_a22oi_1 _27143_ (.Y(_08363_),
    .B1(_08362_),
    .B2(net402),
    .A2(net515),
    .A1(net1212));
 sg13g2_nand2_1 _27144_ (.Y(_08364_),
    .A(\stack[18][1] ),
    .B(_08356_));
 sg13g2_nand2_1 _27145_ (.Y(_08365_),
    .A(_08363_),
    .B(_08364_));
 sg13g2_mux2_1 _27146_ (.A0(_08365_),
    .A1(net105),
    .S(net59),
    .X(_02596_));
 sg13g2_a22oi_1 _27147_ (.Y(_08366_),
    .B1(_08362_),
    .B2(_07978_),
    .A2(net515),
    .A1(net1217));
 sg13g2_nand2_1 _27148_ (.Y(_08367_),
    .A(\stack[18][2] ),
    .B(_08356_));
 sg13g2_nand2_1 _27149_ (.Y(_08368_),
    .A(_08366_),
    .B(_08367_));
 sg13g2_mux2_1 _27150_ (.A0(_08368_),
    .A1(net104),
    .S(net59),
    .X(_02597_));
 sg13g2_a22oi_1 _27151_ (.Y(_08369_),
    .B1(_08362_),
    .B2(net494),
    .A2(net515),
    .A1(net1211));
 sg13g2_nand2_1 _27152_ (.Y(_08370_),
    .A(\stack[18][3] ),
    .B(_08356_));
 sg13g2_nand2_1 _27153_ (.Y(_08371_),
    .A(_08369_),
    .B(_08370_));
 sg13g2_mux2_1 _27154_ (.A0(_08371_),
    .A1(net91),
    .S(net59),
    .X(_02598_));
 sg13g2_a221oi_1 _27155_ (.B2(\stack[18][4] ),
    .C1(_08350_),
    .B1(_08356_),
    .A1(_08158_),
    .Y(_08372_),
    .A2(net515));
 sg13g2_a21oi_1 _27156_ (.A1(net102),
    .A2(net59),
    .Y(_08373_),
    .B1(_08372_));
 sg13g2_a21o_1 _27157_ (.A2(_08362_),
    .A1(net476),
    .B1(_08373_),
    .X(_02599_));
 sg13g2_a221oi_1 _27158_ (.B2(\stack[18][5] ),
    .C1(_08350_),
    .B1(_08356_),
    .A1(net1214),
    .Y(_08374_),
    .A2(net515));
 sg13g2_a21oi_1 _27159_ (.A1(net88),
    .A2(net59),
    .Y(_08375_),
    .B1(_08374_));
 sg13g2_a21o_1 _27160_ (.A2(_08362_),
    .A1(net403),
    .B1(_08375_),
    .X(_02600_));
 sg13g2_and2_1 _27161_ (.A(_07997_),
    .B(net59),
    .X(_08376_));
 sg13g2_a221oi_1 _27162_ (.B2(\stack[18][6] ),
    .C1(_08351_),
    .B1(_08356_),
    .A1(net879),
    .Y(_08377_),
    .A2(net515));
 sg13g2_nand2_1 _27163_ (.Y(_08378_),
    .A(net405),
    .B(_08362_));
 sg13g2_o21ai_1 _27164_ (.B1(_08378_),
    .Y(_02601_),
    .A1(_08376_),
    .A2(_08377_));
 sg13g2_a221oi_1 _27165_ (.B2(net294),
    .C1(net59),
    .B1(_08362_),
    .A1(net1215),
    .Y(_08379_),
    .A2(_08353_));
 sg13g2_nand2_1 _27166_ (.Y(_08380_),
    .A(\stack[18][7] ),
    .B(_08356_));
 sg13g2_a22oi_1 _27167_ (.Y(_02602_),
    .B1(_08379_),
    .B2(_08380_),
    .A2(_08351_),
    .A1(net45));
 sg13g2_inv_1 _27168_ (.Y(_08381_),
    .A(net141));
 sg13g2_nor2_2 _27169_ (.A(_07545_),
    .B(_07609_),
    .Y(_08382_));
 sg13g2_nand2_1 _27170_ (.Y(_08383_),
    .A(net140),
    .B(_08382_));
 sg13g2_nor3_1 _27171_ (.A(_08381_),
    .B(net126),
    .C(_08383_),
    .Y(_08384_));
 sg13g2_buf_2 _27172_ (.A(_08384_),
    .X(_08385_));
 sg13g2_buf_1 _27173_ (.A(_08385_),
    .X(_08386_));
 sg13g2_nor2_1 _27174_ (.A(net516),
    .B(_08275_),
    .Y(_08387_));
 sg13g2_buf_1 _27175_ (.A(_08387_),
    .X(_08388_));
 sg13g2_buf_1 _27176_ (.A(_08388_),
    .X(_08389_));
 sg13g2_buf_1 _27177_ (.A(net1270),
    .X(_08390_));
 sg13g2_nor3_1 _27178_ (.A(net297),
    .B(_08192_),
    .C(net122),
    .Y(_08391_));
 sg13g2_buf_1 _27179_ (.A(_08391_),
    .X(_08392_));
 sg13g2_nor2_1 _27180_ (.A(net878),
    .B(net83),
    .Y(_08393_));
 sg13g2_buf_2 _27181_ (.A(_08393_),
    .X(_08394_));
 sg13g2_nor2b_1 _27182_ (.A(net475),
    .B_N(\stack[19][0] ),
    .Y(_08395_));
 sg13g2_a22oi_1 _27183_ (.Y(_08396_),
    .B1(_08394_),
    .B2(_08395_),
    .A2(net475),
    .A1(net1226));
 sg13g2_a22oi_1 _27184_ (.Y(_08397_),
    .B1(net84),
    .B2(net131),
    .A2(net83),
    .A1(net453));
 sg13g2_o21ai_1 _27185_ (.B1(_08397_),
    .Y(_02603_),
    .A1(net84),
    .A2(_08396_));
 sg13g2_nor2b_1 _27186_ (.A(_08388_),
    .B_N(\stack[19][1] ),
    .Y(_08398_));
 sg13g2_a22oi_1 _27187_ (.Y(_08399_),
    .B1(_08394_),
    .B2(_08398_),
    .A2(net475),
    .A1(net883));
 sg13g2_a22oi_1 _27188_ (.Y(_08400_),
    .B1(net84),
    .B2(_07702_),
    .A2(net83),
    .A1(net447));
 sg13g2_o21ai_1 _27189_ (.B1(_08400_),
    .Y(_02604_),
    .A1(net84),
    .A2(_08399_));
 sg13g2_nor2b_1 _27190_ (.A(_08388_),
    .B_N(\stack[19][2] ),
    .Y(_08401_));
 sg13g2_a22oi_1 _27191_ (.Y(_08402_),
    .B1(_08394_),
    .B2(_08401_),
    .A2(net475),
    .A1(net882));
 sg13g2_a22oi_1 _27192_ (.Y(_08403_),
    .B1(_08385_),
    .B2(net104),
    .A2(net83),
    .A1(_07707_));
 sg13g2_o21ai_1 _27193_ (.B1(_08403_),
    .Y(_02605_),
    .A1(net84),
    .A2(_08402_));
 sg13g2_nor2b_1 _27194_ (.A(_08388_),
    .B_N(\stack[19][3] ),
    .Y(_08404_));
 sg13g2_a22oi_1 _27195_ (.Y(_08405_),
    .B1(_08394_),
    .B2(_08404_),
    .A2(net475),
    .A1(net881));
 sg13g2_a22oi_1 _27196_ (.Y(_08406_),
    .B1(_08385_),
    .B2(_07785_),
    .A2(net83),
    .A1(_07745_));
 sg13g2_o21ai_1 _27197_ (.B1(_08406_),
    .Y(_02606_),
    .A1(net84),
    .A2(_08405_));
 sg13g2_nor2b_1 _27198_ (.A(_08388_),
    .B_N(\stack[19][4] ),
    .Y(_08407_));
 sg13g2_a22oi_1 _27199_ (.Y(_08408_),
    .B1(_08394_),
    .B2(_08407_),
    .A2(net475),
    .A1(net1222));
 sg13g2_a22oi_1 _27200_ (.Y(_08409_),
    .B1(_08385_),
    .B2(_08058_),
    .A2(net83),
    .A1(_10191_));
 sg13g2_o21ai_1 _27201_ (.B1(_08409_),
    .Y(_02607_),
    .A1(net84),
    .A2(_08408_));
 sg13g2_and2_1 _27202_ (.A(_07848_),
    .B(_08385_),
    .X(_08410_));
 sg13g2_nor2b_1 _27203_ (.A(_08388_),
    .B_N(\stack[19][5] ),
    .Y(_08411_));
 sg13g2_a221oi_1 _27204_ (.B2(_08411_),
    .C1(_08385_),
    .B1(_08394_),
    .A1(net1216),
    .Y(_08412_),
    .A2(net475));
 sg13g2_nand2_1 _27205_ (.Y(_08413_),
    .A(net401),
    .B(net83));
 sg13g2_o21ai_1 _27206_ (.B1(_08413_),
    .Y(_02608_),
    .A1(_08410_),
    .A2(_08412_));
 sg13g2_nor2b_1 _27207_ (.A(_08388_),
    .B_N(\stack[19][6] ),
    .Y(_08414_));
 sg13g2_a22oi_1 _27208_ (.Y(_08415_),
    .B1(_08394_),
    .B2(_08414_),
    .A2(net475),
    .A1(net880));
 sg13g2_a22oi_1 _27209_ (.Y(_08416_),
    .B1(_08385_),
    .B2(_07900_),
    .A2(net83),
    .A1(_08000_));
 sg13g2_o21ai_1 _27210_ (.B1(_08416_),
    .Y(_02609_),
    .A1(net84),
    .A2(_08415_));
 sg13g2_nor2b_1 _27211_ (.A(_08389_),
    .B_N(\stack[19][7] ),
    .Y(_08417_));
 sg13g2_a22oi_1 _27212_ (.Y(_08418_),
    .B1(_08394_),
    .B2(_08417_),
    .A2(_08389_),
    .A1(net1215));
 sg13g2_a21oi_1 _27213_ (.A1(_08006_),
    .A2(_08392_),
    .Y(_08419_),
    .B1(_08386_));
 sg13g2_a22oi_1 _27214_ (.Y(_02610_),
    .B1(_08418_),
    .B2(_08419_),
    .A2(_08386_),
    .A1(net45));
 sg13g2_nor4_1 _27215_ (.A(_07604_),
    .B(net136),
    .C(net135),
    .D(_08035_),
    .Y(_08420_));
 sg13g2_buf_1 _27216_ (.A(_08420_),
    .X(_08421_));
 sg13g2_nor2_1 _27217_ (.A(_07594_),
    .B(net522),
    .Y(_08422_));
 sg13g2_buf_1 _27218_ (.A(_08422_),
    .X(_08423_));
 sg13g2_a22oi_1 _27219_ (.Y(_08424_),
    .B1(net506),
    .B2(net1226),
    .A2(net115),
    .A1(_07619_));
 sg13g2_nor3_1 _27220_ (.A(net878),
    .B(_08421_),
    .C(_08422_),
    .Y(_08425_));
 sg13g2_buf_2 _27221_ (.A(_08425_),
    .X(_08426_));
 sg13g2_nand2_1 _27222_ (.Y(_08427_),
    .A(\stack[1][0] ),
    .B(_08426_));
 sg13g2_nand2_1 _27223_ (.Y(_08428_),
    .A(_08424_),
    .B(_08427_));
 sg13g2_and2_1 _27224_ (.A(_07621_),
    .B(_08223_),
    .X(_08429_));
 sg13g2_buf_2 _27225_ (.A(_08429_),
    .X(_08430_));
 sg13g2_buf_1 _27226_ (.A(_08430_),
    .X(_08431_));
 sg13g2_mux2_1 _27227_ (.A0(_08428_),
    .A1(net131),
    .S(net82),
    .X(_02611_));
 sg13g2_a22oi_1 _27228_ (.Y(_08432_),
    .B1(_08426_),
    .B2(\stack[1][1] ),
    .A2(_08423_),
    .A1(net883));
 sg13g2_a22oi_1 _27229_ (.Y(_08433_),
    .B1(net115),
    .B2(net295),
    .A2(net82),
    .A1(net105));
 sg13g2_o21ai_1 _27230_ (.B1(_08433_),
    .Y(_02612_),
    .A1(net82),
    .A2(_08432_));
 sg13g2_a22oi_1 _27231_ (.Y(_08434_),
    .B1(_08426_),
    .B2(\stack[1][2] ),
    .A2(_08423_),
    .A1(net882));
 sg13g2_a22oi_1 _27232_ (.Y(_08435_),
    .B1(net115),
    .B2(net400),
    .A2(net82),
    .A1(net104));
 sg13g2_o21ai_1 _27233_ (.B1(_08435_),
    .Y(_02613_),
    .A1(net82),
    .A2(_08434_));
 sg13g2_a22oi_1 _27234_ (.Y(_08436_),
    .B1(_08426_),
    .B2(\stack[1][3] ),
    .A2(net506),
    .A1(net881));
 sg13g2_a22oi_1 _27235_ (.Y(_08437_),
    .B1(net115),
    .B2(net477),
    .A2(_08431_),
    .A1(net91));
 sg13g2_o21ai_1 _27236_ (.B1(_08437_),
    .Y(_02614_),
    .A1(_08431_),
    .A2(_08436_));
 sg13g2_a221oi_1 _27237_ (.B2(\stack[1][4] ),
    .C1(_08430_),
    .B1(_08426_),
    .A1(net1209),
    .Y(_08438_),
    .A2(net506));
 sg13g2_a21oi_1 _27238_ (.A1(net102),
    .A2(_08430_),
    .Y(_08439_),
    .B1(_08438_));
 sg13g2_a21o_1 _27239_ (.A2(net115),
    .A1(net476),
    .B1(_08439_),
    .X(_02615_));
 sg13g2_nor2_1 _27240_ (.A(net878),
    .B(_08421_),
    .Y(_08440_));
 sg13g2_nor2b_1 _27241_ (.A(net506),
    .B_N(\stack[1][5] ),
    .Y(_08441_));
 sg13g2_a221oi_1 _27242_ (.B2(_08441_),
    .C1(_08430_),
    .B1(_08440_),
    .A1(net1214),
    .Y(_08442_),
    .A2(net506));
 sg13g2_a21oi_1 _27243_ (.A1(_08061_),
    .A2(_08430_),
    .Y(_08443_),
    .B1(_08442_));
 sg13g2_a21o_1 _27244_ (.A2(net115),
    .A1(net403),
    .B1(_08443_),
    .X(_02616_));
 sg13g2_nor2b_1 _27245_ (.A(net506),
    .B_N(\stack[1][6] ),
    .Y(_08444_));
 sg13g2_a22oi_1 _27246_ (.Y(_08445_),
    .B1(_08440_),
    .B2(_08444_),
    .A2(net506),
    .A1(_07854_));
 sg13g2_a22oi_1 _27247_ (.Y(_08446_),
    .B1(net115),
    .B2(net405),
    .A2(_08430_),
    .A1(net46));
 sg13g2_o21ai_1 _27248_ (.B1(_08446_),
    .Y(_02617_),
    .A1(net82),
    .A2(_08445_));
 sg13g2_nand2_1 _27249_ (.Y(_08447_),
    .A(\stack[1][7] ),
    .B(_08426_));
 sg13g2_a221oi_1 _27250_ (.B2(_08005_),
    .C1(net82),
    .B1(net506),
    .A1(net294),
    .Y(_08448_),
    .A2(net115));
 sg13g2_a22oi_1 _27251_ (.Y(_02618_),
    .B1(_08447_),
    .B2(_08448_),
    .A2(net82),
    .A1(_07929_));
 sg13g2_nor2_1 _27252_ (.A(_09654_),
    .B(_07532_),
    .Y(_08449_));
 sg13g2_nand2_1 _27253_ (.Y(_08450_),
    .A(_07475_),
    .B(_08449_));
 sg13g2_buf_2 _27254_ (.A(_08450_),
    .X(_08451_));
 sg13g2_nor2_1 _27255_ (.A(_07600_),
    .B(_08451_),
    .Y(_08452_));
 sg13g2_buf_2 _27256_ (.A(_08452_),
    .X(_08453_));
 sg13g2_nor2_1 _27257_ (.A(net1191),
    .B(_08453_),
    .Y(_08454_));
 sg13g2_nand4_1 _27258_ (.B(net138),
    .C(net299),
    .A(net128),
    .Y(_08455_),
    .D(_08281_));
 sg13g2_buf_1 _27259_ (.A(_08455_),
    .X(_08456_));
 sg13g2_and2_1 _27260_ (.A(_08454_),
    .B(_08456_),
    .X(_08457_));
 sg13g2_buf_1 _27261_ (.A(_08457_),
    .X(_08458_));
 sg13g2_a21oi_1 _27262_ (.A1(net1218),
    .A2(_08453_),
    .Y(_08459_),
    .B1(net58));
 sg13g2_and2_1 _27263_ (.A(_07530_),
    .B(_08382_),
    .X(_08460_));
 sg13g2_buf_2 _27264_ (.A(_08460_),
    .X(_08461_));
 sg13g2_and3_1 _27265_ (.X(_08462_),
    .A(net141),
    .B(_07585_),
    .C(_08461_));
 sg13g2_buf_2 _27266_ (.A(_08462_),
    .X(_08463_));
 sg13g2_mux2_1 _27267_ (.A0(_08459_),
    .A1(net123),
    .S(_08463_),
    .X(_08464_));
 sg13g2_nand2b_1 _27268_ (.Y(_08465_),
    .B(_07620_),
    .A_N(_08456_));
 sg13g2_buf_8 _27269_ (.A(_08463_),
    .X(_08466_));
 sg13g2_nor2_1 _27270_ (.A(\stack[20][0] ),
    .B(net57),
    .Y(_08467_));
 sg13g2_a22oi_1 _27271_ (.Y(_02619_),
    .B1(_08467_),
    .B2(net58),
    .A2(_08465_),
    .A1(_08464_));
 sg13g2_a22oi_1 _27272_ (.Y(_08468_),
    .B1(net58),
    .B2(\stack[20][1] ),
    .A2(_08453_),
    .A1(net883));
 sg13g2_nor4_2 _27273_ (.A(net491),
    .B(_07755_),
    .C(_08289_),
    .Y(_08469_),
    .D(net122));
 sg13g2_a22oi_1 _27274_ (.Y(_08470_),
    .B1(_08469_),
    .B2(net295),
    .A2(net57),
    .A1(_07702_));
 sg13g2_o21ai_1 _27275_ (.B1(_08470_),
    .Y(_02620_),
    .A1(net57),
    .A2(_08468_));
 sg13g2_a22oi_1 _27276_ (.Y(_08471_),
    .B1(net58),
    .B2(\stack[20][2] ),
    .A2(_08453_),
    .A1(net882));
 sg13g2_a22oi_1 _27277_ (.Y(_08472_),
    .B1(_08469_),
    .B2(net400),
    .A2(net57),
    .A1(_07740_));
 sg13g2_o21ai_1 _27278_ (.B1(_08472_),
    .Y(_02621_),
    .A1(net57),
    .A2(_08471_));
 sg13g2_a22oi_1 _27279_ (.Y(_08473_),
    .B1(net58),
    .B2(\stack[20][3] ),
    .A2(_08453_),
    .A1(net881));
 sg13g2_a22oi_1 _27280_ (.Y(_08474_),
    .B1(_08469_),
    .B2(net477),
    .A2(_08463_),
    .A1(net91));
 sg13g2_o21ai_1 _27281_ (.B1(_08474_),
    .Y(_02622_),
    .A1(net57),
    .A2(_08473_));
 sg13g2_a22oi_1 _27282_ (.Y(_08475_),
    .B1(net58),
    .B2(\stack[20][4] ),
    .A2(_08453_),
    .A1(_08117_));
 sg13g2_mux2_1 _27283_ (.A0(_08475_),
    .A1(net98),
    .S(_08463_),
    .X(_08476_));
 sg13g2_o21ai_1 _27284_ (.B1(_08476_),
    .Y(_02623_),
    .A1(net496),
    .A2(_08456_));
 sg13g2_nand2_1 _27285_ (.Y(_08477_),
    .A(_10023_),
    .B(_08453_));
 sg13g2_o21ai_1 _27286_ (.B1(_08477_),
    .Y(_08478_),
    .A1(net472),
    .A2(_08456_));
 sg13g2_and2_1 _27287_ (.A(\stack[20][5] ),
    .B(net58),
    .X(_08479_));
 sg13g2_nor3_1 _27288_ (.A(net57),
    .B(_08478_),
    .C(_08479_),
    .Y(_08480_));
 sg13g2_a21oi_1 _27289_ (.A1(net89),
    .A2(net57),
    .Y(_02624_),
    .B1(_08480_));
 sg13g2_a22oi_1 _27290_ (.Y(_08481_),
    .B1(_08458_),
    .B2(\stack[20][6] ),
    .A2(_08453_),
    .A1(net880));
 sg13g2_a22oi_1 _27291_ (.Y(_08482_),
    .B1(_08469_),
    .B2(net405),
    .A2(_08463_),
    .A1(net46));
 sg13g2_o21ai_1 _27292_ (.B1(_08482_),
    .Y(_02625_),
    .A1(_08466_),
    .A2(_08481_));
 sg13g2_nor2_1 _27293_ (.A(\stack[20][7] ),
    .B(_08463_),
    .Y(_08483_));
 sg13g2_nor3_1 _27294_ (.A(_10025_),
    .B(_08302_),
    .C(_08451_),
    .Y(_08484_));
 sg13g2_and2_1 _27295_ (.A(net445),
    .B(_08469_),
    .X(_08485_));
 sg13g2_nor4_1 _27296_ (.A(_08463_),
    .B(_08458_),
    .C(_08484_),
    .D(_08485_),
    .Y(_08486_));
 sg13g2_a221oi_1 _27297_ (.B2(_08483_),
    .C1(_08486_),
    .B1(net58),
    .A1(_08075_),
    .Y(_02626_),
    .A2(_08466_));
 sg13g2_nor2_1 _27298_ (.A(net522),
    .B(_08451_),
    .Y(_08487_));
 sg13g2_buf_1 _27299_ (.A(_08487_),
    .X(_08488_));
 sg13g2_and4_1 _27300_ (.A(net136),
    .B(net142),
    .C(net404),
    .D(_08281_),
    .X(_08489_));
 sg13g2_buf_1 _27301_ (.A(_08489_),
    .X(_08490_));
 sg13g2_nor3_1 _27302_ (.A(net1191),
    .B(net505),
    .C(net114),
    .Y(_08491_));
 sg13g2_buf_1 _27303_ (.A(_08491_),
    .X(_08492_));
 sg13g2_a21oi_1 _27304_ (.A1(net1218),
    .A2(net505),
    .Y(_08493_),
    .B1(net81));
 sg13g2_nor4_1 _27305_ (.A(net140),
    .B(_08381_),
    .C(net126),
    .D(net122),
    .Y(_08494_));
 sg13g2_buf_2 _27306_ (.A(_08494_),
    .X(_08495_));
 sg13g2_mux2_1 _27307_ (.A0(_08493_),
    .A1(_08235_),
    .S(_08495_),
    .X(_08496_));
 sg13g2_nand2_1 _27308_ (.Y(_08497_),
    .A(net453),
    .B(net114));
 sg13g2_buf_1 _27309_ (.A(_08495_),
    .X(_08498_));
 sg13g2_nor2_1 _27310_ (.A(\stack[21][0] ),
    .B(net80),
    .Y(_08499_));
 sg13g2_a22oi_1 _27311_ (.Y(_02627_),
    .B1(_08499_),
    .B2(net81),
    .A2(_08497_),
    .A1(_08496_));
 sg13g2_a22oi_1 _27312_ (.Y(_08500_),
    .B1(net81),
    .B2(\stack[21][1] ),
    .A2(net505),
    .A1(net883));
 sg13g2_a22oi_1 _27313_ (.Y(_08501_),
    .B1(net114),
    .B2(net295),
    .A2(net80),
    .A1(net105));
 sg13g2_o21ai_1 _27314_ (.B1(_08501_),
    .Y(_02628_),
    .A1(net80),
    .A2(_08500_));
 sg13g2_a22oi_1 _27315_ (.Y(_08502_),
    .B1(net81),
    .B2(\stack[21][2] ),
    .A2(net505),
    .A1(net882));
 sg13g2_a22oi_1 _27316_ (.Y(_08503_),
    .B1(net114),
    .B2(net400),
    .A2(_08498_),
    .A1(_07740_));
 sg13g2_o21ai_1 _27317_ (.B1(_08503_),
    .Y(_02629_),
    .A1(net80),
    .A2(_08502_));
 sg13g2_a22oi_1 _27318_ (.Y(_08504_),
    .B1(net81),
    .B2(\stack[21][3] ),
    .A2(net505),
    .A1(net881));
 sg13g2_a22oi_1 _27319_ (.Y(_08505_),
    .B1(net114),
    .B2(net477),
    .A2(net80),
    .A1(_07785_));
 sg13g2_o21ai_1 _27320_ (.B1(_08505_),
    .Y(_02630_),
    .A1(net80),
    .A2(_08504_));
 sg13g2_a221oi_1 _27321_ (.B2(\stack[21][4] ),
    .C1(_08495_),
    .B1(net81),
    .A1(net1209),
    .Y(_08506_),
    .A2(net505));
 sg13g2_a21oi_1 _27322_ (.A1(_07824_),
    .A2(_08495_),
    .Y(_08507_),
    .B1(_08506_));
 sg13g2_a21o_1 _27323_ (.A2(net114),
    .A1(net476),
    .B1(_08507_),
    .X(_02631_));
 sg13g2_a221oi_1 _27324_ (.B2(\stack[21][5] ),
    .C1(_08495_),
    .B1(net81),
    .A1(net1214),
    .Y(_08508_),
    .A2(net505));
 sg13g2_a21oi_1 _27325_ (.A1(_08061_),
    .A2(_08495_),
    .Y(_08509_),
    .B1(_08508_));
 sg13g2_a21o_1 _27326_ (.A2(net114),
    .A1(net403),
    .B1(_08509_),
    .X(_02632_));
 sg13g2_a22oi_1 _27327_ (.Y(_08510_),
    .B1(net81),
    .B2(\stack[21][6] ),
    .A2(_08488_),
    .A1(net880));
 sg13g2_a22oi_1 _27328_ (.Y(_08511_),
    .B1(net114),
    .B2(net405),
    .A2(_08495_),
    .A1(net46));
 sg13g2_o21ai_1 _27329_ (.B1(_08511_),
    .Y(_02633_),
    .A1(net80),
    .A2(_08510_));
 sg13g2_and2_1 _27330_ (.A(net445),
    .B(_08490_),
    .X(_08512_));
 sg13g2_a221oi_1 _27331_ (.B2(\stack[21][7] ),
    .C1(_08512_),
    .B1(_08492_),
    .A1(net1219),
    .Y(_08513_),
    .A2(net505));
 sg13g2_nor2b_1 _27332_ (.A(_08498_),
    .B_N(_08513_),
    .Y(_08514_));
 sg13g2_a21oi_1 _27333_ (.A1(net43),
    .A2(net80),
    .Y(_02634_),
    .B1(_08514_));
 sg13g2_nor3_1 _27334_ (.A(_07934_),
    .B(net138),
    .C(_08089_),
    .Y(_08515_));
 sg13g2_o21ai_1 _27335_ (.B1(net1304),
    .Y(_08516_),
    .A1(_08183_),
    .A2(_08451_));
 sg13g2_a21oi_1 _27336_ (.A1(net124),
    .A2(_08515_),
    .Y(_08517_),
    .B1(_08516_));
 sg13g2_buf_2 _27337_ (.A(_08517_),
    .X(_08518_));
 sg13g2_nand2_1 _27338_ (.Y(_08519_),
    .A(\stack[22][0] ),
    .B(_08518_));
 sg13g2_and2_1 _27339_ (.A(net124),
    .B(_08515_),
    .X(_08520_));
 sg13g2_buf_1 _27340_ (.A(_08520_),
    .X(_08521_));
 sg13g2_nor2_1 _27341_ (.A(net532),
    .B(_08451_),
    .Y(_08522_));
 sg13g2_buf_2 _27342_ (.A(_08522_),
    .X(_08523_));
 sg13g2_a22oi_1 _27343_ (.Y(_08524_),
    .B1(_08523_),
    .B2(net1218),
    .A2(_08521_),
    .A1(_07619_));
 sg13g2_nand2_1 _27344_ (.Y(_08525_),
    .A(_08519_),
    .B(_08524_));
 sg13g2_nand2_1 _27345_ (.Y(_08526_),
    .A(net137),
    .B(net133));
 sg13g2_nor2_1 _27346_ (.A(net122),
    .B(_08526_),
    .Y(_08527_));
 sg13g2_buf_2 _27347_ (.A(_08527_),
    .X(_08528_));
 sg13g2_buf_1 _27348_ (.A(_08528_),
    .X(_08529_));
 sg13g2_mux2_1 _27349_ (.A0(_08525_),
    .A1(net131),
    .S(net79),
    .X(_02635_));
 sg13g2_a22oi_1 _27350_ (.Y(_08530_),
    .B1(_08518_),
    .B2(\stack[22][1] ),
    .A2(_08523_),
    .A1(_07668_));
 sg13g2_buf_1 _27351_ (.A(_07700_),
    .X(_08531_));
 sg13g2_nand2_1 _27352_ (.Y(_08532_),
    .A(_07545_),
    .B(_07609_));
 sg13g2_buf_1 _27353_ (.A(_08532_),
    .X(_08533_));
 sg13g2_nor4_2 _27354_ (.A(_07751_),
    .B(net129),
    .C(_08533_),
    .Y(_08534_),
    .D(_08192_));
 sg13g2_a22oi_1 _27355_ (.Y(_08535_),
    .B1(_08534_),
    .B2(net295),
    .A2(net79),
    .A1(net113));
 sg13g2_o21ai_1 _27356_ (.B1(_08535_),
    .Y(_02636_),
    .A1(net79),
    .A2(_08530_));
 sg13g2_a22oi_1 _27357_ (.Y(_08536_),
    .B1(_08518_),
    .B2(\stack[22][2] ),
    .A2(_08523_),
    .A1(_07705_));
 sg13g2_buf_1 _27358_ (.A(_07738_),
    .X(_08537_));
 sg13g2_a22oi_1 _27359_ (.Y(_08538_),
    .B1(_08534_),
    .B2(_08297_),
    .A2(net79),
    .A1(net112));
 sg13g2_o21ai_1 _27360_ (.B1(_08538_),
    .Y(_02637_),
    .A1(net79),
    .A2(_08536_));
 sg13g2_a22oi_1 _27361_ (.Y(_08539_),
    .B1(_08518_),
    .B2(\stack[22][3] ),
    .A2(_08523_),
    .A1(_07743_));
 sg13g2_a22oi_1 _27362_ (.Y(_08540_),
    .B1(_08534_),
    .B2(net477),
    .A2(net79),
    .A1(net101));
 sg13g2_o21ai_1 _27363_ (.B1(_08540_),
    .Y(_02638_),
    .A1(net79),
    .A2(_08539_));
 sg13g2_a221oi_1 _27364_ (.B2(\stack[22][4] ),
    .C1(_08528_),
    .B1(_08518_),
    .A1(net1209),
    .Y(_08541_),
    .A2(_08523_));
 sg13g2_a21oi_1 _27365_ (.A1(net102),
    .A2(_08528_),
    .Y(_08542_),
    .B1(_08541_));
 sg13g2_a21o_1 _27366_ (.A2(_08521_),
    .A1(net476),
    .B1(_08542_),
    .X(_02639_));
 sg13g2_a221oi_1 _27367_ (.B2(net1216),
    .C1(_08528_),
    .B1(_08523_),
    .A1(_08121_),
    .Y(_08543_),
    .A2(_08521_));
 sg13g2_nand2_1 _27368_ (.Y(_08544_),
    .A(\stack[22][5] ),
    .B(_08518_));
 sg13g2_a22oi_1 _27369_ (.Y(_02640_),
    .B1(_08543_),
    .B2(_08544_),
    .A2(net79),
    .A1(net89));
 sg13g2_a22oi_1 _27370_ (.Y(_08545_),
    .B1(_08518_),
    .B2(\stack[22][6] ),
    .A2(_08523_),
    .A1(net880));
 sg13g2_a22oi_1 _27371_ (.Y(_08546_),
    .B1(_08534_),
    .B2(_07857_),
    .A2(_08528_),
    .A1(_07900_));
 sg13g2_o21ai_1 _27372_ (.B1(_08546_),
    .Y(_02641_),
    .A1(_08529_),
    .A2(_08545_));
 sg13g2_a221oi_1 _27373_ (.B2(_08005_),
    .C1(_08528_),
    .B1(_08523_),
    .A1(_08347_),
    .Y(_08547_),
    .A2(_08521_));
 sg13g2_nand2_1 _27374_ (.Y(_08548_),
    .A(\stack[22][7] ),
    .B(_08518_));
 sg13g2_a22oi_1 _27375_ (.Y(_02642_),
    .B1(_08547_),
    .B2(_08548_),
    .A2(_08529_),
    .A1(_07929_));
 sg13g2_nor2_1 _27376_ (.A(_08016_),
    .B(_08451_),
    .Y(_08549_));
 sg13g2_buf_1 _27377_ (.A(_08549_),
    .X(_08550_));
 sg13g2_and4_1 _27378_ (.A(net143),
    .B(_07610_),
    .C(_08012_),
    .D(_08181_),
    .X(_08551_));
 sg13g2_buf_1 _27379_ (.A(_08551_),
    .X(_08552_));
 sg13g2_nor3_1 _27380_ (.A(net1191),
    .B(net504),
    .C(net111),
    .Y(_08553_));
 sg13g2_buf_1 _27381_ (.A(_08553_),
    .X(_08554_));
 sg13g2_a21oi_1 _27382_ (.A1(_07961_),
    .A2(net504),
    .Y(_08555_),
    .B1(net78));
 sg13g2_nand3_1 _27383_ (.B(net139),
    .C(net125),
    .A(net140),
    .Y(_08556_));
 sg13g2_nor3_1 _27384_ (.A(_08381_),
    .B(net126),
    .C(_08556_),
    .Y(_08557_));
 sg13g2_buf_2 _27385_ (.A(_08557_),
    .X(_08558_));
 sg13g2_mux2_1 _27386_ (.A0(_08555_),
    .A1(_08235_),
    .S(_08558_),
    .X(_08559_));
 sg13g2_nand2_1 _27387_ (.Y(_08560_),
    .A(net453),
    .B(net111));
 sg13g2_buf_8 _27388_ (.A(_08558_),
    .X(_08561_));
 sg13g2_nor2_1 _27389_ (.A(\stack[23][0] ),
    .B(net56),
    .Y(_08562_));
 sg13g2_a22oi_1 _27390_ (.Y(_02643_),
    .B1(_08562_),
    .B2(net78),
    .A2(_08560_),
    .A1(_08559_));
 sg13g2_a22oi_1 _27391_ (.Y(_08563_),
    .B1(net78),
    .B2(\stack[23][1] ),
    .A2(net504),
    .A1(_07668_));
 sg13g2_a22oi_1 _27392_ (.Y(_08564_),
    .B1(net111),
    .B2(_08294_),
    .A2(net56),
    .A1(net113));
 sg13g2_o21ai_1 _27393_ (.B1(_08564_),
    .Y(_02644_),
    .A1(net56),
    .A2(_08563_));
 sg13g2_a22oi_1 _27394_ (.Y(_08565_),
    .B1(net78),
    .B2(\stack[23][2] ),
    .A2(net504),
    .A1(_07705_));
 sg13g2_a22oi_1 _27395_ (.Y(_08566_),
    .B1(net111),
    .B2(net400),
    .A2(net56),
    .A1(net112));
 sg13g2_o21ai_1 _27396_ (.B1(_08566_),
    .Y(_02645_),
    .A1(net56),
    .A2(_08565_));
 sg13g2_a22oi_1 _27397_ (.Y(_08567_),
    .B1(net78),
    .B2(\stack[23][3] ),
    .A2(net504),
    .A1(_07743_));
 sg13g2_a22oi_1 _27398_ (.Y(_08568_),
    .B1(net111),
    .B2(net477),
    .A2(_08561_),
    .A1(net101));
 sg13g2_o21ai_1 _27399_ (.B1(_08568_),
    .Y(_02646_),
    .A1(_08561_),
    .A2(_08567_));
 sg13g2_a221oi_1 _27400_ (.B2(\stack[23][4] ),
    .C1(_08558_),
    .B1(_08554_),
    .A1(net1209),
    .Y(_08569_),
    .A2(_08550_));
 sg13g2_a21oi_1 _27401_ (.A1(net102),
    .A2(_08558_),
    .Y(_08570_),
    .B1(_08569_));
 sg13g2_a21o_1 _27402_ (.A2(_08552_),
    .A1(net476),
    .B1(_08570_),
    .X(_02647_));
 sg13g2_a221oi_1 _27403_ (.B2(\stack[23][5] ),
    .C1(_08558_),
    .B1(net78),
    .A1(net1214),
    .Y(_08571_),
    .A2(net504));
 sg13g2_a21oi_1 _27404_ (.A1(_07849_),
    .A2(_08558_),
    .Y(_08572_),
    .B1(_08571_));
 sg13g2_a21o_1 _27405_ (.A2(net111),
    .A1(_08060_),
    .B1(_08572_),
    .X(_02648_));
 sg13g2_a22oi_1 _27406_ (.Y(_08573_),
    .B1(net78),
    .B2(\stack[23][6] ),
    .A2(net504),
    .A1(net880));
 sg13g2_a22oi_1 _27407_ (.Y(_08574_),
    .B1(net111),
    .B2(_07857_),
    .A2(_08558_),
    .A1(_07899_));
 sg13g2_o21ai_1 _27408_ (.B1(_08574_),
    .Y(_02649_),
    .A1(net56),
    .A2(_08573_));
 sg13g2_and2_1 _27409_ (.A(_09660_),
    .B(net111),
    .X(_08575_));
 sg13g2_a221oi_1 _27410_ (.B2(\stack[23][7] ),
    .C1(_08575_),
    .B1(net78),
    .A1(net1213),
    .Y(_08576_),
    .A2(net504));
 sg13g2_nor2b_1 _27411_ (.A(net56),
    .B_N(_08576_),
    .Y(_08577_));
 sg13g2_a21oi_1 _27412_ (.A1(net43),
    .A2(net56),
    .Y(_02650_),
    .B1(_08577_));
 sg13g2_nand2_1 _27413_ (.Y(_08578_),
    .A(net137),
    .B(_08182_));
 sg13g2_o21ai_1 _27414_ (.B1(_08578_),
    .Y(_08579_),
    .A1(net296),
    .A2(_08288_));
 sg13g2_nand2_1 _27415_ (.Y(_08580_),
    .A(_07475_),
    .B(_07940_));
 sg13g2_buf_2 _27416_ (.A(_08580_),
    .X(_08581_));
 sg13g2_o21ai_1 _27417_ (.B1(net1304),
    .Y(_08582_),
    .A1(_07600_),
    .A2(_08581_));
 sg13g2_buf_1 _27418_ (.A(_08582_),
    .X(_08583_));
 sg13g2_a21o_1 _27419_ (.A2(_08579_),
    .A1(_07936_),
    .B1(_08583_),
    .X(_08584_));
 sg13g2_buf_2 _27420_ (.A(_08584_),
    .X(_08585_));
 sg13g2_nor2_1 _27421_ (.A(net121),
    .B(_08578_),
    .Y(_08586_));
 sg13g2_buf_2 _27422_ (.A(_08586_),
    .X(_08587_));
 sg13g2_buf_1 _27423_ (.A(_08587_),
    .X(_08588_));
 sg13g2_nor4_1 _27424_ (.A(net491),
    .B(_07754_),
    .C(net121),
    .D(net97),
    .Y(_08589_));
 sg13g2_buf_2 _27425_ (.A(_08589_),
    .X(_08590_));
 sg13g2_nor2_1 _27426_ (.A(net521),
    .B(_08581_),
    .Y(_08591_));
 sg13g2_buf_2 _27427_ (.A(_08591_),
    .X(_08592_));
 sg13g2_nand2_1 _27428_ (.Y(_08593_),
    .A(net1208),
    .B(_08592_));
 sg13g2_nor2_1 _27429_ (.A(_08587_),
    .B(_08593_),
    .Y(_08594_));
 sg13g2_a221oi_1 _27430_ (.B2(net478),
    .C1(_08594_),
    .B1(_08590_),
    .A1(net134),
    .Y(_08595_),
    .A2(net55));
 sg13g2_nor2_1 _27431_ (.A(\stack[24][0] ),
    .B(_08585_),
    .Y(_08596_));
 sg13g2_a21oi_1 _27432_ (.A1(_08585_),
    .A2(_08595_),
    .Y(_02651_),
    .B1(_08596_));
 sg13g2_nand2_1 _27433_ (.Y(_08597_),
    .A(net1225),
    .B(_08592_));
 sg13g2_a22oi_1 _27434_ (.Y(_08598_),
    .B1(_08590_),
    .B2(net473),
    .A2(_08587_),
    .A1(_07701_));
 sg13g2_o21ai_1 _27435_ (.B1(_08598_),
    .Y(_08599_),
    .A1(net55),
    .A2(_08597_));
 sg13g2_mux2_1 _27436_ (.A0(\stack[24][1] ),
    .A1(_08599_),
    .S(_08585_),
    .X(_02652_));
 sg13g2_nand2_1 _27437_ (.Y(_08600_),
    .A(net1224),
    .B(_08592_));
 sg13g2_a22oi_1 _27438_ (.Y(_08601_),
    .B1(_08590_),
    .B2(_10183_),
    .A2(_08587_),
    .A1(net118));
 sg13g2_o21ai_1 _27439_ (.B1(_08601_),
    .Y(_08602_),
    .A1(net55),
    .A2(_08600_));
 sg13g2_mux2_1 _27440_ (.A0(\stack[24][2] ),
    .A1(_08602_),
    .S(_08585_),
    .X(_02653_));
 sg13g2_nand2_1 _27441_ (.Y(_08603_),
    .A(net1223),
    .B(_08592_));
 sg13g2_a22oi_1 _27442_ (.Y(_08604_),
    .B1(_08590_),
    .B2(_10177_),
    .A2(_08587_),
    .A1(_07783_));
 sg13g2_o21ai_1 _27443_ (.B1(_08604_),
    .Y(_08605_),
    .A1(net55),
    .A2(_08603_));
 sg13g2_mux2_1 _27444_ (.A0(\stack[24][3] ),
    .A1(_08605_),
    .S(_08585_),
    .X(_02654_));
 sg13g2_a21oi_1 _27445_ (.A1(net1222),
    .A2(_08592_),
    .Y(_08606_),
    .B1(net55));
 sg13g2_a21oi_1 _27446_ (.A1(net102),
    .A2(net55),
    .Y(_08607_),
    .B1(_08606_));
 sg13g2_a21oi_1 _27447_ (.A1(_07936_),
    .A2(_08579_),
    .Y(_08608_),
    .B1(_08583_));
 sg13g2_a22oi_1 _27448_ (.Y(_08609_),
    .B1(_08590_),
    .B2(net484),
    .A2(_08608_),
    .A1(\stack[24][4] ));
 sg13g2_nand2b_1 _27449_ (.Y(_02655_),
    .B(_08609_),
    .A_N(_08607_));
 sg13g2_a21oi_1 _27450_ (.A1(_07991_),
    .A2(_08592_),
    .Y(_08610_),
    .B1(net55));
 sg13g2_nor3_1 _27451_ (.A(net296),
    .B(net121),
    .C(net97),
    .Y(_08611_));
 sg13g2_nor2_1 _27452_ (.A(_08583_),
    .B(_08590_),
    .Y(_08612_));
 sg13g2_a21oi_1 _27453_ (.A1(net401),
    .A2(_08611_),
    .Y(_08613_),
    .B1(_08612_));
 sg13g2_nor2_1 _27454_ (.A(\stack[24][5] ),
    .B(_08585_),
    .Y(_08614_));
 sg13g2_a221oi_1 _27455_ (.B2(_08613_),
    .C1(_08614_),
    .B1(_08610_),
    .A1(net88),
    .Y(_02656_),
    .A2(net55));
 sg13g2_nor4_1 _27456_ (.A(_10018_),
    .B(net521),
    .C(_08581_),
    .D(_08587_),
    .Y(_08615_));
 sg13g2_a221oi_1 _27457_ (.B2(net451),
    .C1(_08615_),
    .B1(_08611_),
    .A1(_07899_),
    .Y(_08616_),
    .A2(_08588_));
 sg13g2_nor2_1 _27458_ (.A(\stack[24][6] ),
    .B(_08585_),
    .Y(_08617_));
 sg13g2_a21oi_1 _27459_ (.A1(_08585_),
    .A2(_08616_),
    .Y(_02657_),
    .B1(_08617_));
 sg13g2_nand2_1 _27460_ (.Y(_08618_),
    .A(_07889_),
    .B(_07906_));
 sg13g2_or2_1 _27461_ (.X(_08619_),
    .B(_08618_),
    .A(_07914_));
 sg13g2_xnor2_1 _27462_ (.Y(_08620_),
    .A(_07447_),
    .B(_07905_));
 sg13g2_o21ai_1 _27463_ (.B1(_08620_),
    .Y(_08621_),
    .A1(_07910_),
    .A2(_07912_));
 sg13g2_nand2_1 _27464_ (.Y(_08622_),
    .A(net518),
    .B(_08588_));
 sg13g2_a21o_1 _27465_ (.A2(_08621_),
    .A1(_08619_),
    .B1(_08622_),
    .X(_08623_));
 sg13g2_nand2_1 _27466_ (.Y(_08624_),
    .A(_07925_),
    .B(_08587_));
 sg13g2_a21o_1 _27467_ (.A2(_08592_),
    .A1(_08076_),
    .B1(_08587_),
    .X(_08625_));
 sg13g2_a221oi_1 _27468_ (.B2(_08625_),
    .C1(_08608_),
    .B1(_08624_),
    .A1(net294),
    .Y(_08626_),
    .A2(_08590_));
 sg13g2_a22oi_1 _27469_ (.Y(_02658_),
    .B1(_08623_),
    .B2(_08626_),
    .A2(_08608_),
    .A1(_07426_));
 sg13g2_nor3_1 _27470_ (.A(_08532_),
    .B(_08028_),
    .C(_08288_),
    .Y(_08627_));
 sg13g2_buf_2 _27471_ (.A(_08627_),
    .X(_08628_));
 sg13g2_nand4_1 _27472_ (.B(net125),
    .C(net404),
    .A(_07547_),
    .Y(_08629_),
    .D(net133));
 sg13g2_nor2_1 _27473_ (.A(net522),
    .B(_08581_),
    .Y(_08630_));
 sg13g2_buf_1 _27474_ (.A(_08630_),
    .X(_08631_));
 sg13g2_nor2_1 _27475_ (.A(net1270),
    .B(net503),
    .Y(_08632_));
 sg13g2_and2_1 _27476_ (.A(_08629_),
    .B(_08632_),
    .X(_08633_));
 sg13g2_buf_1 _27477_ (.A(_08633_),
    .X(_08634_));
 sg13g2_nand2b_1 _27478_ (.Y(_08635_),
    .B(_08634_),
    .A_N(_08628_));
 sg13g2_buf_8 _27479_ (.A(_08635_),
    .X(_08636_));
 sg13g2_buf_1 _27480_ (.A(_08628_),
    .X(_08637_));
 sg13g2_nor3_1 _27481_ (.A(net121),
    .B(net297),
    .C(net97),
    .Y(_08638_));
 sg13g2_buf_1 _27482_ (.A(_08638_),
    .X(_08639_));
 sg13g2_nand2_1 _27483_ (.Y(_08640_),
    .A(net1208),
    .B(net503));
 sg13g2_nor2_1 _27484_ (.A(_08628_),
    .B(_08640_),
    .Y(_08641_));
 sg13g2_a221oi_1 _27485_ (.B2(net480),
    .C1(_08641_),
    .B1(_08639_),
    .A1(net134),
    .Y(_08642_),
    .A2(net54));
 sg13g2_nor2_1 _27486_ (.A(\stack[25][0] ),
    .B(net40),
    .Y(_08643_));
 sg13g2_a21oi_1 _27487_ (.A1(net40),
    .A2(_08642_),
    .Y(_02659_),
    .B1(_08643_));
 sg13g2_nand2_1 _27488_ (.Y(_08644_),
    .A(_10021_),
    .B(net503));
 sg13g2_nor2_1 _27489_ (.A(_08628_),
    .B(_08644_),
    .Y(_08645_));
 sg13g2_a221oi_1 _27490_ (.B2(net447),
    .C1(_08645_),
    .B1(_08639_),
    .A1(net113),
    .Y(_08646_),
    .A2(net54));
 sg13g2_nor2_1 _27491_ (.A(\stack[25][1] ),
    .B(net40),
    .Y(_08647_));
 sg13g2_a21oi_1 _27492_ (.A1(net40),
    .A2(_08646_),
    .Y(_02660_),
    .B1(_08647_));
 sg13g2_nand2_1 _27493_ (.Y(_08648_),
    .A(net1301),
    .B(_08631_));
 sg13g2_nor2_1 _27494_ (.A(_08628_),
    .B(_08648_),
    .Y(_08649_));
 sg13g2_a221oi_1 _27495_ (.B2(net452),
    .C1(_08649_),
    .B1(_08639_),
    .A1(net112),
    .Y(_08650_),
    .A2(_08628_));
 sg13g2_nor2_1 _27496_ (.A(\stack[25][2] ),
    .B(net40),
    .Y(_08651_));
 sg13g2_a21oi_1 _27497_ (.A1(net40),
    .A2(_08650_),
    .Y(_02661_),
    .B1(_08651_));
 sg13g2_nand2_1 _27498_ (.Y(_08652_),
    .A(net1300),
    .B(net503));
 sg13g2_nor2_1 _27499_ (.A(_08628_),
    .B(_08652_),
    .Y(_08653_));
 sg13g2_a221oi_1 _27500_ (.B2(net492),
    .C1(_08653_),
    .B1(_08639_),
    .A1(net101),
    .Y(_08654_),
    .A2(_08628_));
 sg13g2_nor2_1 _27501_ (.A(\stack[25][3] ),
    .B(_08636_),
    .Y(_08655_));
 sg13g2_a21oi_1 _27502_ (.A1(_08636_),
    .A2(_08654_),
    .Y(_02662_),
    .B1(_08655_));
 sg13g2_nand2_1 _27503_ (.Y(_08656_),
    .A(\stack[25][4] ),
    .B(_08634_));
 sg13g2_a221oi_1 _27504_ (.B2(net1222),
    .C1(net54),
    .B1(net503),
    .A1(net484),
    .Y(_08657_),
    .A2(_08639_));
 sg13g2_a22oi_1 _27505_ (.Y(_02663_),
    .B1(_08656_),
    .B2(_08657_),
    .A2(net54),
    .A1(net100));
 sg13g2_and2_1 _27506_ (.A(_07850_),
    .B(net503),
    .X(_08658_));
 sg13g2_nor2_1 _27507_ (.A(net446),
    .B(_08629_),
    .Y(_08659_));
 sg13g2_and2_1 _27508_ (.A(\stack[25][5] ),
    .B(_08634_),
    .X(_08660_));
 sg13g2_nor4_1 _27509_ (.A(net54),
    .B(_08658_),
    .C(_08659_),
    .D(_08660_),
    .Y(_08661_));
 sg13g2_a21oi_1 _27510_ (.A1(net89),
    .A2(net54),
    .Y(_02664_),
    .B1(_08661_));
 sg13g2_a21oi_1 _27511_ (.A1(net879),
    .A2(net503),
    .Y(_08662_),
    .B1(_08634_));
 sg13g2_a21oi_1 _27512_ (.A1(net449),
    .A2(_08639_),
    .Y(_08663_),
    .B1(_08637_));
 sg13g2_nor2_1 _27513_ (.A(\stack[25][6] ),
    .B(net40),
    .Y(_08664_));
 sg13g2_a221oi_1 _27514_ (.B2(_08663_),
    .C1(_08664_),
    .B1(_08662_),
    .A1(_07997_),
    .Y(_02665_),
    .A2(net54));
 sg13g2_a221oi_1 _27515_ (.B2(net1215),
    .C1(net54),
    .B1(net503),
    .A1(net294),
    .Y(_08665_),
    .A2(_08639_));
 sg13g2_nor2_1 _27516_ (.A(\stack[25][7] ),
    .B(_08635_),
    .Y(_08666_));
 sg13g2_a221oi_1 _27517_ (.B2(_08665_),
    .C1(_08666_),
    .B1(net40),
    .A1(net41),
    .Y(_02666_),
    .A2(_08637_));
 sg13g2_nor2_1 _27518_ (.A(net532),
    .B(_08581_),
    .Y(_08667_));
 sg13g2_buf_1 _27519_ (.A(_08667_),
    .X(_08668_));
 sg13g2_nand4_1 _27520_ (.B(net135),
    .C(_07946_),
    .A(net136),
    .Y(_08669_),
    .D(_08181_));
 sg13g2_buf_1 _27521_ (.A(_08669_),
    .X(_08670_));
 sg13g2_nand3b_1 _27522_ (.B(_08670_),
    .C(_09907_),
    .Y(_08671_),
    .A_N(_08668_));
 sg13g2_nand4_1 _27523_ (.B(_08081_),
    .C(net137),
    .A(_07547_),
    .Y(_08672_),
    .D(net133));
 sg13g2_buf_1 _27524_ (.A(_08672_),
    .X(_08673_));
 sg13g2_nand2b_1 _27525_ (.Y(_08674_),
    .B(_08673_),
    .A_N(_08671_));
 sg13g2_buf_1 _27526_ (.A(_08674_),
    .X(_08675_));
 sg13g2_buf_1 _27527_ (.A(_08675_),
    .X(_08676_));
 sg13g2_nor3_2 _27528_ (.A(net296),
    .B(net117),
    .C(net116),
    .Y(_08677_));
 sg13g2_buf_1 _27529_ (.A(_08673_),
    .X(_08678_));
 sg13g2_nand3_1 _27530_ (.B(net77),
    .C(_08668_),
    .A(net1302),
    .Y(_08679_));
 sg13g2_o21ai_1 _27531_ (.B1(_08679_),
    .Y(_08680_),
    .A1(net123),
    .A2(net77));
 sg13g2_a21oi_1 _27532_ (.A1(net478),
    .A2(_08677_),
    .Y(_08681_),
    .B1(_08680_));
 sg13g2_nor2_1 _27533_ (.A(\stack[26][0] ),
    .B(net39),
    .Y(_08682_));
 sg13g2_a21oi_1 _27534_ (.A1(net39),
    .A2(_08681_),
    .Y(_02667_),
    .B1(_08682_));
 sg13g2_nor2_1 _27535_ (.A(net121),
    .B(_08526_),
    .Y(_08683_));
 sg13g2_buf_1 _27536_ (.A(_08683_),
    .X(_08684_));
 sg13g2_and3_1 _27537_ (.X(_08685_),
    .A(net1225),
    .B(net77),
    .C(_08668_));
 sg13g2_a221oi_1 _27538_ (.B2(net447),
    .C1(_08685_),
    .B1(_08677_),
    .A1(net113),
    .Y(_08686_),
    .A2(_08684_));
 sg13g2_nor2_1 _27539_ (.A(\stack[26][1] ),
    .B(net39),
    .Y(_08687_));
 sg13g2_a21oi_1 _27540_ (.A1(net39),
    .A2(_08686_),
    .Y(_02668_),
    .B1(_08687_));
 sg13g2_and3_1 _27541_ (.X(_08688_),
    .A(net1224),
    .B(net77),
    .C(_08668_));
 sg13g2_a221oi_1 _27542_ (.B2(net452),
    .C1(_08688_),
    .B1(_08677_),
    .A1(net112),
    .Y(_08689_),
    .A2(_08684_));
 sg13g2_nor2_1 _27543_ (.A(\stack[26][2] ),
    .B(net39),
    .Y(_08690_));
 sg13g2_a21oi_1 _27544_ (.A1(net39),
    .A2(_08689_),
    .Y(_02669_),
    .B1(_08690_));
 sg13g2_nor4_1 _27545_ (.A(net491),
    .B(net129),
    .C(net117),
    .D(net116),
    .Y(_08691_));
 sg13g2_and3_1 _27546_ (.X(_08692_),
    .A(net1223),
    .B(net77),
    .C(_08668_));
 sg13g2_a221oi_1 _27547_ (.B2(net492),
    .C1(_08692_),
    .B1(_08691_),
    .A1(net101),
    .Y(_08693_),
    .A2(_08684_));
 sg13g2_nor2_1 _27548_ (.A(\stack[26][3] ),
    .B(net39),
    .Y(_08694_));
 sg13g2_a21oi_1 _27549_ (.A1(net39),
    .A2(_08693_),
    .Y(_02670_),
    .B1(_08694_));
 sg13g2_and2_1 _27550_ (.A(_08678_),
    .B(_08668_),
    .X(_08695_));
 sg13g2_a22oi_1 _27551_ (.Y(_08696_),
    .B1(_08695_),
    .B2(net1210),
    .A2(_08677_),
    .A1(net493));
 sg13g2_o21ai_1 _27552_ (.B1(_08696_),
    .Y(_08697_),
    .A1(net98),
    .A2(_08678_));
 sg13g2_mux2_1 _27553_ (.A0(\stack[26][4] ),
    .A1(_08697_),
    .S(_08676_),
    .X(_02671_));
 sg13g2_or2_1 _27554_ (.X(_08698_),
    .B(_08670_),
    .A(_10127_));
 sg13g2_nand2_1 _27555_ (.Y(_08699_),
    .A(net1298),
    .B(_08668_));
 sg13g2_nand4_1 _27556_ (.B(_08671_),
    .C(_08698_),
    .A(net77),
    .Y(_08700_),
    .D(_08699_));
 sg13g2_o21ai_1 _27557_ (.B1(_08700_),
    .Y(_08701_),
    .A1(\stack[26][5] ),
    .A2(_08675_));
 sg13g2_a21oi_1 _27558_ (.A1(net89),
    .A2(_08684_),
    .Y(_02672_),
    .B1(_08701_));
 sg13g2_nor2_1 _27559_ (.A(_10134_),
    .B(_08670_),
    .Y(_08702_));
 sg13g2_a221oi_1 _27560_ (.B2(net879),
    .C1(_08702_),
    .B1(_08695_),
    .A1(_07899_),
    .Y(_08703_),
    .A2(_08684_));
 sg13g2_nor2_1 _27561_ (.A(\stack[26][6] ),
    .B(_08675_),
    .Y(_08704_));
 sg13g2_a21oi_1 _27562_ (.A1(_08676_),
    .A2(_08703_),
    .Y(_02673_),
    .B1(_08704_));
 sg13g2_a21oi_1 _27563_ (.A1(_08619_),
    .A2(_08621_),
    .Y(_08705_),
    .B1(_07780_));
 sg13g2_inv_1 _27564_ (.Y(_08706_),
    .A(\stack[26][7] ));
 sg13g2_nor3_1 _27565_ (.A(_10025_),
    .B(net532),
    .C(_08581_),
    .Y(_08707_));
 sg13g2_nor2_1 _27566_ (.A(_07925_),
    .B(net77),
    .Y(_08708_));
 sg13g2_a221oi_1 _27567_ (.B2(net77),
    .C1(_08708_),
    .B1(_08707_),
    .A1(net445),
    .Y(_08709_),
    .A2(_08691_));
 sg13g2_o21ai_1 _27568_ (.B1(_08709_),
    .Y(_08710_),
    .A1(_08706_),
    .A2(_08675_));
 sg13g2_a21o_1 _27569_ (.A2(_08684_),
    .A1(_08705_),
    .B1(_08710_),
    .X(_02674_));
 sg13g2_nor3_1 _27570_ (.A(_07968_),
    .B(_08028_),
    .C(net116),
    .Y(_08711_));
 sg13g2_buf_2 _27571_ (.A(_08711_),
    .X(_08712_));
 sg13g2_and4_1 _27572_ (.A(net136),
    .B(net135),
    .C(net404),
    .D(_08182_),
    .X(_08713_));
 sg13g2_buf_2 _27573_ (.A(_08713_),
    .X(_08714_));
 sg13g2_nor2_1 _27574_ (.A(net516),
    .B(_08581_),
    .Y(_08715_));
 sg13g2_buf_2 _27575_ (.A(_08715_),
    .X(_08716_));
 sg13g2_nor3_2 _27576_ (.A(net878),
    .B(_08714_),
    .C(_08716_),
    .Y(_08717_));
 sg13g2_nand2b_1 _27577_ (.Y(_08718_),
    .B(_08717_),
    .A_N(_08712_));
 sg13g2_buf_1 _27578_ (.A(_08718_),
    .X(_08719_));
 sg13g2_buf_1 _27579_ (.A(_08712_),
    .X(_08720_));
 sg13g2_nand2_1 _27580_ (.Y(_08721_),
    .A(net1208),
    .B(_08716_));
 sg13g2_nor2_1 _27581_ (.A(net53),
    .B(_08721_),
    .Y(_08722_));
 sg13g2_a221oi_1 _27582_ (.B2(net480),
    .C1(_08722_),
    .B1(_08714_),
    .A1(_07664_),
    .Y(_08723_),
    .A2(net53));
 sg13g2_nor2_1 _27583_ (.A(\stack[27][0] ),
    .B(net38),
    .Y(_08724_));
 sg13g2_a21oi_1 _27584_ (.A1(net38),
    .A2(_08723_),
    .Y(_02675_),
    .B1(_08724_));
 sg13g2_nand2_1 _27585_ (.Y(_08725_),
    .A(_10021_),
    .B(_08716_));
 sg13g2_nor2_1 _27586_ (.A(_08712_),
    .B(_08725_),
    .Y(_08726_));
 sg13g2_a221oi_1 _27587_ (.B2(_08105_),
    .C1(_08726_),
    .B1(_08714_),
    .A1(net113),
    .Y(_08727_),
    .A2(net53));
 sg13g2_nor2_1 _27588_ (.A(\stack[27][1] ),
    .B(net38),
    .Y(_08728_));
 sg13g2_a21oi_1 _27589_ (.A1(net38),
    .A2(_08727_),
    .Y(_02676_),
    .B1(_08728_));
 sg13g2_nand2_1 _27590_ (.Y(_08729_),
    .A(_10015_),
    .B(_08716_));
 sg13g2_nor2_1 _27591_ (.A(_08712_),
    .B(_08729_),
    .Y(_08730_));
 sg13g2_a221oi_1 _27592_ (.B2(net452),
    .C1(_08730_),
    .B1(_08714_),
    .A1(net112),
    .Y(_08731_),
    .A2(net53));
 sg13g2_nor2_1 _27593_ (.A(\stack[27][2] ),
    .B(net38),
    .Y(_08732_));
 sg13g2_a21oi_1 _27594_ (.A1(net38),
    .A2(_08731_),
    .Y(_02677_),
    .B1(_08732_));
 sg13g2_nand2_1 _27595_ (.Y(_08733_),
    .A(net1300),
    .B(_08716_));
 sg13g2_nor2_1 _27596_ (.A(_08712_),
    .B(_08733_),
    .Y(_08734_));
 sg13g2_a221oi_1 _27597_ (.B2(net494),
    .C1(_08734_),
    .B1(_08714_),
    .A1(net101),
    .Y(_08735_),
    .A2(net53));
 sg13g2_nor2_1 _27598_ (.A(\stack[27][3] ),
    .B(net38),
    .Y(_08736_));
 sg13g2_a21oi_1 _27599_ (.A1(net38),
    .A2(_08735_),
    .Y(_02678_),
    .B1(_08736_));
 sg13g2_inv_1 _27600_ (.Y(_08737_),
    .A(\stack[27][4] ));
 sg13g2_nor2b_1 _27601_ (.A(_08712_),
    .B_N(_08717_),
    .Y(_08738_));
 sg13g2_nand2_1 _27602_ (.Y(_08739_),
    .A(_10191_),
    .B(_08714_));
 sg13g2_a21oi_1 _27603_ (.A1(net1210),
    .A2(_08716_),
    .Y(_08740_),
    .B1(_08717_));
 sg13g2_inv_1 _27604_ (.Y(_08741_),
    .A(_08712_));
 sg13g2_mux2_1 _27605_ (.A0(net98),
    .A1(_08740_),
    .S(_08741_),
    .X(_08742_));
 sg13g2_a22oi_1 _27606_ (.Y(_02679_),
    .B1(_08739_),
    .B2(_08742_),
    .A2(_08738_),
    .A1(_08737_));
 sg13g2_a21oi_1 _27607_ (.A1(_07991_),
    .A2(_08716_),
    .Y(_08743_),
    .B1(_08717_));
 sg13g2_nor3_1 _27608_ (.A(net117),
    .B(net297),
    .C(net116),
    .Y(_08744_));
 sg13g2_a21oi_1 _27609_ (.A1(net401),
    .A2(_08744_),
    .Y(_08745_),
    .B1(net53));
 sg13g2_nor2_1 _27610_ (.A(\stack[27][5] ),
    .B(_08719_),
    .Y(_08746_));
 sg13g2_a221oi_1 _27611_ (.B2(_08745_),
    .C1(_08746_),
    .B1(_08743_),
    .A1(net88),
    .Y(_02680_),
    .A2(_08720_));
 sg13g2_inv_1 _27612_ (.Y(_08747_),
    .A(\stack[27][6] ));
 sg13g2_nand2_1 _27613_ (.Y(_08748_),
    .A(net42),
    .B(net53));
 sg13g2_nor3_1 _27614_ (.A(_10018_),
    .B(_08017_),
    .C(_08581_),
    .Y(_08749_));
 sg13g2_a221oi_1 _27615_ (.B2(_08741_),
    .C1(_08738_),
    .B1(_08749_),
    .A1(net449),
    .Y(_08750_),
    .A2(_08744_));
 sg13g2_a22oi_1 _27616_ (.Y(_02681_),
    .B1(_08748_),
    .B2(_08750_),
    .A2(_08738_),
    .A1(_08747_));
 sg13g2_a221oi_1 _27617_ (.B2(net1215),
    .C1(net53),
    .B1(_08716_),
    .A1(net294),
    .Y(_08751_),
    .A2(_08714_));
 sg13g2_nor2_1 _27618_ (.A(\stack[27][7] ),
    .B(_08718_),
    .Y(_08752_));
 sg13g2_a221oi_1 _27619_ (.B2(_08751_),
    .C1(_08752_),
    .B1(_08719_),
    .A1(_08075_),
    .Y(_02682_),
    .A2(_08720_));
 sg13g2_nand2_1 _27620_ (.Y(_08753_),
    .A(_07475_),
    .B(_08084_));
 sg13g2_buf_2 _27621_ (.A(_08753_),
    .X(_08754_));
 sg13g2_nor2_1 _27622_ (.A(_07600_),
    .B(_08754_),
    .Y(_08755_));
 sg13g2_buf_2 _27623_ (.A(_08755_),
    .X(_08756_));
 sg13g2_nand4_1 _27624_ (.B(net125),
    .C(_07947_),
    .A(_07934_),
    .Y(_08757_),
    .D(net133));
 sg13g2_nand3b_1 _27625_ (.B(_08757_),
    .C(_09907_),
    .Y(_08758_),
    .A_N(_08756_));
 sg13g2_buf_1 _27626_ (.A(_08758_),
    .X(_08759_));
 sg13g2_or2_1 _27627_ (.X(_08760_),
    .B(_08578_),
    .A(_07968_));
 sg13g2_buf_2 _27628_ (.A(_08760_),
    .X(_08761_));
 sg13g2_nand2b_1 _27629_ (.Y(_08762_),
    .B(_08761_),
    .A_N(_08759_));
 sg13g2_buf_2 _27630_ (.A(_08762_),
    .X(_08763_));
 sg13g2_nor3_2 _27631_ (.A(net296),
    .B(_07969_),
    .C(net97),
    .Y(_08764_));
 sg13g2_and4_1 _27632_ (.A(net128),
    .B(_08081_),
    .C(net137),
    .D(net124),
    .X(_08765_));
 sg13g2_buf_1 _27633_ (.A(_08765_),
    .X(_08766_));
 sg13g2_buf_1 _27634_ (.A(_08766_),
    .X(_08767_));
 sg13g2_a21oi_1 _27635_ (.A1(net1302),
    .A2(_08756_),
    .Y(_08768_),
    .B1(net76));
 sg13g2_a21oi_1 _27636_ (.A1(net123),
    .A2(net76),
    .Y(_08769_),
    .B1(_08768_));
 sg13g2_a21oi_1 _27637_ (.A1(net478),
    .A2(_08764_),
    .Y(_08770_),
    .B1(_08769_));
 sg13g2_nor2_1 _27638_ (.A(\stack[28][0] ),
    .B(_08763_),
    .Y(_08771_));
 sg13g2_a21oi_1 _27639_ (.A1(_08763_),
    .A2(_08770_),
    .Y(_02683_),
    .B1(_08771_));
 sg13g2_nand3_1 _27640_ (.B(_08761_),
    .C(_08756_),
    .A(net1212),
    .Y(_08772_));
 sg13g2_nor4_2 _27641_ (.A(net491),
    .B(net129),
    .C(_07969_),
    .Y(_08773_),
    .D(net97));
 sg13g2_a22oi_1 _27642_ (.Y(_08774_),
    .B1(_08773_),
    .B2(net402),
    .A2(net76),
    .A1(net119));
 sg13g2_nand2_1 _27643_ (.Y(_08775_),
    .A(_08772_),
    .B(_08774_));
 sg13g2_mux2_1 _27644_ (.A0(\stack[28][1] ),
    .A1(_08775_),
    .S(_08763_),
    .X(_02684_));
 sg13g2_nand3_1 _27645_ (.B(_08761_),
    .C(_08756_),
    .A(net1224),
    .Y(_08776_));
 sg13g2_a22oi_1 _27646_ (.Y(_08777_),
    .B1(_08773_),
    .B2(net485),
    .A2(net76),
    .A1(_07738_));
 sg13g2_and2_1 _27647_ (.A(_08776_),
    .B(_08777_),
    .X(_08778_));
 sg13g2_nor2_1 _27648_ (.A(\stack[28][2] ),
    .B(_08763_),
    .Y(_08779_));
 sg13g2_a21oi_1 _27649_ (.A1(_08763_),
    .A2(_08778_),
    .Y(_02685_),
    .B1(_08779_));
 sg13g2_and3_1 _27650_ (.X(_08780_),
    .A(_07742_),
    .B(_08761_),
    .C(_08756_));
 sg13g2_a221oi_1 _27651_ (.B2(net494),
    .C1(_08780_),
    .B1(_08773_),
    .A1(net103),
    .Y(_08781_),
    .A2(net76));
 sg13g2_nor2_1 _27652_ (.A(\stack[28][3] ),
    .B(_08763_),
    .Y(_08782_));
 sg13g2_a21oi_1 _27653_ (.A1(_08763_),
    .A2(_08781_),
    .Y(_02686_),
    .B1(_08782_));
 sg13g2_nor2b_1 _27654_ (.A(_08766_),
    .B_N(_08756_),
    .Y(_08783_));
 sg13g2_a22oi_1 _27655_ (.Y(_08784_),
    .B1(_08783_),
    .B2(net1210),
    .A2(_08764_),
    .A1(net493));
 sg13g2_o21ai_1 _27656_ (.B1(_08784_),
    .Y(_08785_),
    .A1(net98),
    .A2(_08761_));
 sg13g2_mux2_1 _27657_ (.A0(\stack[28][4] ),
    .A1(_08785_),
    .S(_08763_),
    .X(_02687_));
 sg13g2_nor2_1 _27658_ (.A(_08767_),
    .B(_08759_),
    .Y(_08786_));
 sg13g2_a21oi_1 _27659_ (.A1(net1298),
    .A2(_08756_),
    .Y(_08787_),
    .B1(net76));
 sg13g2_nand2_1 _27660_ (.Y(_08788_),
    .A(_08759_),
    .B(_08787_));
 sg13g2_a21oi_1 _27661_ (.A1(net401),
    .A2(_08764_),
    .Y(_08789_),
    .B1(_08788_));
 sg13g2_a221oi_1 _27662_ (.B2(_07347_),
    .C1(_08789_),
    .B1(_08786_),
    .A1(net88),
    .Y(_02688_),
    .A2(_08767_));
 sg13g2_inv_1 _27663_ (.Y(_08790_),
    .A(\stack[28][6] ));
 sg13g2_nand2_1 _27664_ (.Y(_08791_),
    .A(net42),
    .B(net76));
 sg13g2_nor3_1 _27665_ (.A(_10018_),
    .B(net521),
    .C(_08754_),
    .Y(_08792_));
 sg13g2_a221oi_1 _27666_ (.B2(_08761_),
    .C1(_08786_),
    .B1(_08792_),
    .A1(_08000_),
    .Y(_08793_),
    .A2(_08773_));
 sg13g2_a22oi_1 _27667_ (.Y(_02689_),
    .B1(_08791_),
    .B2(_08793_),
    .A2(_08786_),
    .A1(_08790_));
 sg13g2_inv_1 _27668_ (.Y(_08794_),
    .A(\stack[28][7] ));
 sg13g2_or2_1 _27669_ (.X(_08795_),
    .B(_08759_),
    .A(_08794_));
 sg13g2_a22oi_1 _27670_ (.Y(_08796_),
    .B1(_08764_),
    .B2(net294),
    .A2(_08756_),
    .A1(net1219));
 sg13g2_and3_1 _27671_ (.X(_08797_),
    .A(_08761_),
    .B(_08795_),
    .C(_08796_));
 sg13g2_a21oi_1 _27672_ (.A1(net43),
    .A2(net76),
    .Y(_02690_),
    .B1(_08797_));
 sg13g2_or3_1 _27673_ (.A(_07968_),
    .B(_08028_),
    .C(_08288_),
    .X(_08798_));
 sg13g2_buf_2 _27674_ (.A(_08798_),
    .X(_08799_));
 sg13g2_nor2_1 _27675_ (.A(net134),
    .B(_08799_),
    .Y(_08800_));
 sg13g2_nor2_1 _27676_ (.A(net522),
    .B(_08754_),
    .Y(_08801_));
 sg13g2_buf_2 _27677_ (.A(_08801_),
    .X(_08802_));
 sg13g2_nor3_1 _27678_ (.A(net117),
    .B(net126),
    .C(_08288_),
    .Y(_08803_));
 sg13g2_buf_1 _27679_ (.A(_08803_),
    .X(_08804_));
 sg13g2_a21oi_1 _27680_ (.A1(net1208),
    .A2(_08802_),
    .Y(_08805_),
    .B1(net75));
 sg13g2_and4_1 _27681_ (.A(net136),
    .B(_07609_),
    .C(_08011_),
    .D(net133),
    .X(_08806_));
 sg13g2_buf_8 _27682_ (.A(_08806_),
    .X(_08807_));
 sg13g2_nand2_1 _27683_ (.Y(_08808_),
    .A(net480),
    .B(net110));
 sg13g2_o21ai_1 _27684_ (.B1(_08808_),
    .Y(_08809_),
    .A1(_08800_),
    .A2(_08805_));
 sg13g2_nor3_1 _27685_ (.A(net1270),
    .B(_08802_),
    .C(net110),
    .Y(_08810_));
 sg13g2_nand2_1 _27686_ (.Y(_08811_),
    .A(_08799_),
    .B(_08810_));
 sg13g2_buf_1 _27687_ (.A(_08811_),
    .X(_08812_));
 sg13g2_mux2_1 _27688_ (.A0(\stack[29][0] ),
    .A1(_08809_),
    .S(net37),
    .X(_02691_));
 sg13g2_and3_1 _27689_ (.X(_08813_),
    .A(_07667_),
    .B(_08799_),
    .C(_08802_));
 sg13g2_a221oi_1 _27690_ (.B2(net402),
    .C1(_08813_),
    .B1(net110),
    .A1(net113),
    .Y(_08814_),
    .A2(net75));
 sg13g2_nor2_1 _27691_ (.A(\stack[29][1] ),
    .B(net37),
    .Y(_08815_));
 sg13g2_a21oi_1 _27692_ (.A1(net37),
    .A2(_08814_),
    .Y(_02692_),
    .B1(_08815_));
 sg13g2_and3_1 _27693_ (.X(_08816_),
    .A(_07704_),
    .B(_08799_),
    .C(_08802_));
 sg13g2_a221oi_1 _27694_ (.B2(net450),
    .C1(_08816_),
    .B1(net110),
    .A1(net112),
    .Y(_08817_),
    .A2(net75));
 sg13g2_nor2_1 _27695_ (.A(\stack[29][2] ),
    .B(net37),
    .Y(_08818_));
 sg13g2_a21oi_1 _27696_ (.A1(net37),
    .A2(_08817_),
    .Y(_02693_),
    .B1(_08818_));
 sg13g2_and3_1 _27697_ (.X(_08819_),
    .A(_07742_),
    .B(_08799_),
    .C(_08802_));
 sg13g2_a221oi_1 _27698_ (.B2(net494),
    .C1(_08819_),
    .B1(net110),
    .A1(net103),
    .Y(_08820_),
    .A2(net75));
 sg13g2_nor2_1 _27699_ (.A(\stack[29][3] ),
    .B(net37),
    .Y(_08821_));
 sg13g2_a21oi_1 _27700_ (.A1(net37),
    .A2(_08820_),
    .Y(_02694_),
    .B1(_08821_));
 sg13g2_or2_1 _27701_ (.X(_08822_),
    .B(_08754_),
    .A(net522));
 sg13g2_nor2_1 _27702_ (.A(_08252_),
    .B(_08822_),
    .Y(_08823_));
 sg13g2_and2_1 _27703_ (.A(_09864_),
    .B(net110),
    .X(_08824_));
 sg13g2_or4_1 _27704_ (.A(net75),
    .B(_08810_),
    .C(_08823_),
    .D(_08824_),
    .X(_08825_));
 sg13g2_o21ai_1 _27705_ (.B1(_08825_),
    .Y(_08826_),
    .A1(\stack[29][4] ),
    .A2(_08812_));
 sg13g2_a21oi_1 _27706_ (.A1(net100),
    .A2(_08804_),
    .Y(_02695_),
    .B1(_08826_));
 sg13g2_a21o_1 _27707_ (.A2(net110),
    .A1(net471),
    .B1(net75),
    .X(_08827_));
 sg13g2_a221oi_1 _27708_ (.B2(\stack[29][5] ),
    .C1(_08827_),
    .B1(_08810_),
    .A1(net1216),
    .Y(_08828_),
    .A2(_08802_));
 sg13g2_a21oi_1 _27709_ (.A1(net89),
    .A2(net75),
    .Y(_02696_),
    .B1(_08828_));
 sg13g2_nand2_1 _27710_ (.Y(_08829_),
    .A(net451),
    .B(net110));
 sg13g2_nand3_1 _27711_ (.B(_08799_),
    .C(_08802_),
    .A(net1220),
    .Y(_08830_));
 sg13g2_and3_1 _27712_ (.X(_08831_),
    .A(net37),
    .B(_08829_),
    .C(_08830_));
 sg13g2_nand2_1 _27713_ (.Y(_08832_),
    .A(net46),
    .B(net75));
 sg13g2_nor2_1 _27714_ (.A(\stack[29][6] ),
    .B(_08812_),
    .Y(_08833_));
 sg13g2_a21oi_1 _27715_ (.A1(_08831_),
    .A2(_08832_),
    .Y(_02697_),
    .B1(_08833_));
 sg13g2_nand3_1 _27716_ (.B(\stack[29][7] ),
    .C(_08822_),
    .A(net1192),
    .Y(_08834_));
 sg13g2_nand2_1 _27717_ (.Y(_08835_),
    .A(_08076_),
    .B(_08802_));
 sg13g2_o21ai_1 _27718_ (.B1(_08835_),
    .Y(_08836_),
    .A1(_08807_),
    .A2(_08834_));
 sg13g2_a22oi_1 _27719_ (.Y(_08837_),
    .B1(_08836_),
    .B2(_08799_),
    .A2(_08807_),
    .A1(net298));
 sg13g2_o21ai_1 _27720_ (.B1(_08837_),
    .Y(_02698_),
    .A1(net41),
    .A2(_08799_));
 sg13g2_nor2_1 _27721_ (.A(net130),
    .B(_07587_),
    .Y(_08838_));
 sg13g2_buf_2 _27722_ (.A(_08838_),
    .X(_08839_));
 sg13g2_buf_1 _27723_ (.A(_08839_),
    .X(_08840_));
 sg13g2_nor2_1 _27724_ (.A(_07594_),
    .B(net532),
    .Y(_08841_));
 sg13g2_buf_1 _27725_ (.A(_08841_),
    .X(_08842_));
 sg13g2_nor3_1 _27726_ (.A(_07754_),
    .B(_07971_),
    .C(net122),
    .Y(_08843_));
 sg13g2_buf_1 _27727_ (.A(_08843_),
    .X(_08844_));
 sg13g2_nor2_1 _27728_ (.A(net878),
    .B(net74),
    .Y(_08845_));
 sg13g2_nor2b_1 _27729_ (.A(net502),
    .B_N(\stack[2][0] ),
    .Y(_08846_));
 sg13g2_a22oi_1 _27730_ (.Y(_08847_),
    .B1(_08845_),
    .B2(_08846_),
    .A2(net502),
    .A1(net1226));
 sg13g2_a22oi_1 _27731_ (.Y(_08848_),
    .B1(net74),
    .B2(net453),
    .A2(net52),
    .A1(net131));
 sg13g2_o21ai_1 _27732_ (.B1(_08848_),
    .Y(_02699_),
    .A1(net52),
    .A2(_08847_));
 sg13g2_nand4_1 _27733_ (.B(net138),
    .C(net299),
    .A(net128),
    .Y(_08849_),
    .D(_08008_));
 sg13g2_nor2_1 _27734_ (.A(net1191),
    .B(net502),
    .Y(_08850_));
 sg13g2_and2_1 _27735_ (.A(_08849_),
    .B(_08850_),
    .X(_08851_));
 sg13g2_buf_2 _27736_ (.A(_08851_),
    .X(_08852_));
 sg13g2_a22oi_1 _27737_ (.Y(_08853_),
    .B1(_08852_),
    .B2(\stack[2][1] ),
    .A2(net502),
    .A1(net883));
 sg13g2_a22oi_1 _27738_ (.Y(_08854_),
    .B1(net74),
    .B2(net295),
    .A2(net52),
    .A1(net113));
 sg13g2_o21ai_1 _27739_ (.B1(_08854_),
    .Y(_02700_),
    .A1(net52),
    .A2(_08853_));
 sg13g2_a22oi_1 _27740_ (.Y(_08855_),
    .B1(_08852_),
    .B2(\stack[2][2] ),
    .A2(net502),
    .A1(net882));
 sg13g2_a22oi_1 _27741_ (.Y(_08856_),
    .B1(net74),
    .B2(net400),
    .A2(net52),
    .A1(net112));
 sg13g2_o21ai_1 _27742_ (.B1(_08856_),
    .Y(_02701_),
    .A1(_08840_),
    .A2(_08855_));
 sg13g2_nor2b_1 _27743_ (.A(_08842_),
    .B_N(\stack[2][3] ),
    .Y(_08857_));
 sg13g2_a22oi_1 _27744_ (.Y(_08858_),
    .B1(_08845_),
    .B2(_08857_),
    .A2(_08842_),
    .A1(net881));
 sg13g2_a22oi_1 _27745_ (.Y(_08859_),
    .B1(_08844_),
    .B2(net477),
    .A2(_08839_),
    .A1(net101));
 sg13g2_o21ai_1 _27746_ (.B1(_08859_),
    .Y(_02702_),
    .A1(_08840_),
    .A2(_08858_));
 sg13g2_a221oi_1 _27747_ (.B2(\stack[2][4] ),
    .C1(_08839_),
    .B1(_08852_),
    .A1(net1209),
    .Y(_08860_),
    .A2(net502));
 sg13g2_a21oi_1 _27748_ (.A1(_07824_),
    .A2(_08839_),
    .Y(_08861_),
    .B1(_08860_));
 sg13g2_a21o_1 _27749_ (.A2(net74),
    .A1(net476),
    .B1(_08861_),
    .X(_02703_));
 sg13g2_a221oi_1 _27750_ (.B2(\stack[2][5] ),
    .C1(_08839_),
    .B1(_08852_),
    .A1(net1221),
    .Y(_08862_),
    .A2(net502));
 sg13g2_a21oi_1 _27751_ (.A1(_07849_),
    .A2(_08839_),
    .Y(_08863_),
    .B1(_08862_));
 sg13g2_a21o_1 _27752_ (.A2(net74),
    .A1(net403),
    .B1(_08863_),
    .X(_02704_));
 sg13g2_nand2_1 _27753_ (.Y(_08864_),
    .A(net1220),
    .B(net502));
 sg13g2_a22oi_1 _27754_ (.Y(_08865_),
    .B1(_08852_),
    .B2(\stack[2][6] ),
    .A2(net74),
    .A1(_07856_));
 sg13g2_nand2_1 _27755_ (.Y(_08866_),
    .A(_08864_),
    .B(_08865_));
 sg13g2_mux2_1 _27756_ (.A0(_08866_),
    .A1(net42),
    .S(net52),
    .X(_02705_));
 sg13g2_nor3_1 _27757_ (.A(_10025_),
    .B(_07594_),
    .C(_08183_),
    .Y(_08867_));
 sg13g2_a221oi_1 _27758_ (.B2(\stack[2][7] ),
    .C1(_08867_),
    .B1(_08852_),
    .A1(net445),
    .Y(_08868_),
    .A2(net74));
 sg13g2_nor2b_1 _27759_ (.A(net52),
    .B_N(_08868_),
    .Y(_08869_));
 sg13g2_a21oi_1 _27760_ (.A1(net43),
    .A2(net52),
    .Y(_02706_),
    .B1(_08869_));
 sg13g2_nor2_1 _27761_ (.A(_07968_),
    .B(_08526_),
    .Y(_08870_));
 sg13g2_buf_1 _27762_ (.A(_08870_),
    .X(_08871_));
 sg13g2_nor2_1 _27763_ (.A(_07943_),
    .B(_08754_),
    .Y(_08872_));
 sg13g2_buf_1 _27764_ (.A(_08872_),
    .X(_08873_));
 sg13g2_and4_1 _27765_ (.A(net143),
    .B(net142),
    .C(_07947_),
    .D(_07952_),
    .X(_08874_));
 sg13g2_nor3_1 _27766_ (.A(net1270),
    .B(net520),
    .C(_08874_),
    .Y(_08875_));
 sg13g2_buf_1 _27767_ (.A(_08875_),
    .X(_08876_));
 sg13g2_nand2b_1 _27768_ (.Y(_08877_),
    .B(_08876_),
    .A_N(net96));
 sg13g2_buf_2 _27769_ (.A(_08877_),
    .X(_08878_));
 sg13g2_nor3_1 _27770_ (.A(_07748_),
    .B(net129),
    .C(_07971_),
    .Y(_08879_));
 sg13g2_buf_2 _27771_ (.A(_08879_),
    .X(_08880_));
 sg13g2_nand2_1 _27772_ (.Y(_08881_),
    .A(_08238_),
    .B(net520));
 sg13g2_nor2_1 _27773_ (.A(net96),
    .B(_08881_),
    .Y(_08882_));
 sg13g2_a221oi_1 _27774_ (.B2(net480),
    .C1(_08882_),
    .B1(_08880_),
    .A1(net134),
    .Y(_08883_),
    .A2(net96));
 sg13g2_nor2_1 _27775_ (.A(\stack[30][0] ),
    .B(_08878_),
    .Y(_08884_));
 sg13g2_a21oi_1 _27776_ (.A1(_08878_),
    .A2(_08883_),
    .Y(_02707_),
    .B1(_08884_));
 sg13g2_buf_1 _27777_ (.A(net96),
    .X(_08885_));
 sg13g2_nand2_1 _27778_ (.Y(_08886_),
    .A(_07667_),
    .B(net520));
 sg13g2_a22oi_1 _27779_ (.Y(_08887_),
    .B1(_08880_),
    .B2(net473),
    .A2(net96),
    .A1(_07700_));
 sg13g2_o21ai_1 _27780_ (.B1(_08887_),
    .Y(_08888_),
    .A1(net73),
    .A2(_08886_));
 sg13g2_mux2_1 _27781_ (.A0(\stack[30][1] ),
    .A1(_08888_),
    .S(_08878_),
    .X(_02708_));
 sg13g2_nand2_1 _27782_ (.Y(_08889_),
    .A(_07704_),
    .B(net520));
 sg13g2_a22oi_1 _27783_ (.Y(_08890_),
    .B1(_08880_),
    .B2(_10183_),
    .A2(net96),
    .A1(_07739_));
 sg13g2_o21ai_1 _27784_ (.B1(_08890_),
    .Y(_08891_),
    .A1(net73),
    .A2(_08889_));
 sg13g2_mux2_1 _27785_ (.A0(\stack[30][2] ),
    .A1(_08891_),
    .S(_08878_),
    .X(_02709_));
 sg13g2_nand2_1 _27786_ (.Y(_08892_),
    .A(net1300),
    .B(net520));
 sg13g2_nor2_1 _27787_ (.A(net96),
    .B(_08892_),
    .Y(_08893_));
 sg13g2_a221oi_1 _27788_ (.B2(_10178_),
    .C1(_08893_),
    .B1(_08874_),
    .A1(net103),
    .Y(_08894_),
    .A2(net96));
 sg13g2_nor2_1 _27789_ (.A(\stack[30][3] ),
    .B(_08878_),
    .Y(_08895_));
 sg13g2_a21oi_1 _27790_ (.A1(_08878_),
    .A2(_08894_),
    .Y(_02710_),
    .B1(_08895_));
 sg13g2_nor2_1 _27791_ (.A(\stack[30][4] ),
    .B(_08885_),
    .Y(_08896_));
 sg13g2_a21oi_1 _27792_ (.A1(net493),
    .A2(_08880_),
    .Y(_08897_),
    .B1(_08876_));
 sg13g2_a21oi_1 _27793_ (.A1(net1210),
    .A2(_08873_),
    .Y(_08898_),
    .B1(_08871_));
 sg13g2_and2_1 _27794_ (.A(_08897_),
    .B(_08898_),
    .X(_08899_));
 sg13g2_a221oi_1 _27795_ (.B2(_08896_),
    .C1(_08899_),
    .B1(_08876_),
    .A1(net100),
    .Y(_02711_),
    .A2(_08885_));
 sg13g2_a21oi_1 _27796_ (.A1(net1216),
    .A2(net520),
    .Y(_08900_),
    .B1(_08876_));
 sg13g2_a21oi_1 _27797_ (.A1(net401),
    .A2(_08880_),
    .Y(_08901_),
    .B1(net73));
 sg13g2_nor2_1 _27798_ (.A(\stack[30][5] ),
    .B(_08878_),
    .Y(_08902_));
 sg13g2_a221oi_1 _27799_ (.B2(_08901_),
    .C1(_08902_),
    .B1(_08900_),
    .A1(net88),
    .Y(_02712_),
    .A2(net73));
 sg13g2_a21oi_1 _27800_ (.A1(net879),
    .A2(net520),
    .Y(_08903_),
    .B1(_08876_));
 sg13g2_a21oi_1 _27801_ (.A1(net451),
    .A2(_08880_),
    .Y(_08904_),
    .B1(net73));
 sg13g2_nor2_1 _27802_ (.A(\stack[30][6] ),
    .B(_08878_),
    .Y(_08905_));
 sg13g2_a221oi_1 _27803_ (.B2(_08904_),
    .C1(_08905_),
    .B1(_08903_),
    .A1(_07997_),
    .Y(_02713_),
    .A2(net73));
 sg13g2_nand2_1 _27804_ (.Y(_08906_),
    .A(\stack[30][7] ),
    .B(_08876_));
 sg13g2_a221oi_1 _27805_ (.B2(_08006_),
    .C1(net73),
    .B1(_08880_),
    .A1(net1215),
    .Y(_08907_),
    .A2(net520));
 sg13g2_a22oi_1 _27806_ (.Y(_02714_),
    .B1(_08906_),
    .B2(_08907_),
    .A2(net73),
    .A1(net45));
 sg13g2_nand2_1 _27807_ (.Y(_08908_),
    .A(net127),
    .B(_08223_));
 sg13g2_buf_2 _27808_ (.A(_08908_),
    .X(_08909_));
 sg13g2_nor2_1 _27809_ (.A(net516),
    .B(_08754_),
    .Y(_08910_));
 sg13g2_buf_1 _27810_ (.A(_08910_),
    .X(_08911_));
 sg13g2_and4_1 _27811_ (.A(net143),
    .B(net142),
    .C(_07952_),
    .D(net404),
    .X(_08912_));
 sg13g2_buf_1 _27812_ (.A(_08912_),
    .X(_08913_));
 sg13g2_nor3_2 _27813_ (.A(net1191),
    .B(net489),
    .C(net109),
    .Y(_08914_));
 sg13g2_nand2_1 _27814_ (.Y(_08915_),
    .A(_08909_),
    .B(_08914_));
 sg13g2_buf_2 _27815_ (.A(_08915_),
    .X(_08916_));
 sg13g2_and2_1 _27816_ (.A(net127),
    .B(_08223_),
    .X(_08917_));
 sg13g2_buf_1 _27817_ (.A(_08917_),
    .X(_08918_));
 sg13g2_buf_1 _27818_ (.A(_08918_),
    .X(_08919_));
 sg13g2_and3_1 _27819_ (.X(_08920_),
    .A(net1218),
    .B(_08909_),
    .C(net489));
 sg13g2_a221oi_1 _27820_ (.B2(net480),
    .C1(_08920_),
    .B1(net109),
    .A1(net134),
    .Y(_08921_),
    .A2(net72));
 sg13g2_nor2_1 _27821_ (.A(\stack[31][0] ),
    .B(_08916_),
    .Y(_08922_));
 sg13g2_a21oi_1 _27822_ (.A1(_08916_),
    .A2(_08921_),
    .Y(_02715_),
    .B1(_08922_));
 sg13g2_and3_1 _27823_ (.X(_08923_),
    .A(net1225),
    .B(_08909_),
    .C(net489));
 sg13g2_a221oi_1 _27824_ (.B2(net402),
    .C1(_08923_),
    .B1(net109),
    .A1(net119),
    .Y(_08924_),
    .A2(net72));
 sg13g2_nor2_1 _27825_ (.A(\stack[31][1] ),
    .B(_08916_),
    .Y(_08925_));
 sg13g2_a21oi_1 _27826_ (.A1(_08916_),
    .A2(_08924_),
    .Y(_02716_),
    .B1(_08925_));
 sg13g2_and3_1 _27827_ (.X(_08926_),
    .A(net1224),
    .B(_08909_),
    .C(net489));
 sg13g2_a221oi_1 _27828_ (.B2(net450),
    .C1(_08926_),
    .B1(net109),
    .A1(net118),
    .Y(_08927_),
    .A2(net72));
 sg13g2_nor2_1 _27829_ (.A(\stack[31][2] ),
    .B(_08916_),
    .Y(_08928_));
 sg13g2_a21oi_1 _27830_ (.A1(_08916_),
    .A2(_08927_),
    .Y(_02717_),
    .B1(_08928_));
 sg13g2_and3_1 _27831_ (.X(_08929_),
    .A(net1223),
    .B(_08909_),
    .C(net489));
 sg13g2_a221oi_1 _27832_ (.B2(net494),
    .C1(_08929_),
    .B1(net109),
    .A1(net103),
    .Y(_08930_),
    .A2(net72));
 sg13g2_nor2_1 _27833_ (.A(\stack[31][3] ),
    .B(_08916_),
    .Y(_08931_));
 sg13g2_a21oi_1 _27834_ (.A1(_08916_),
    .A2(_08930_),
    .Y(_02718_),
    .B1(_08931_));
 sg13g2_nor2_1 _27835_ (.A(_09858_),
    .B(net72),
    .Y(_08932_));
 sg13g2_inv_1 _27836_ (.Y(_08933_),
    .A(_08913_));
 sg13g2_nor2_1 _27837_ (.A(net496),
    .B(_08933_),
    .Y(_08934_));
 sg13g2_nor3_1 _27838_ (.A(_08252_),
    .B(net516),
    .C(_08754_),
    .Y(_08935_));
 sg13g2_nor4_1 _27839_ (.A(net72),
    .B(_08914_),
    .C(_08934_),
    .D(_08935_),
    .Y(_08936_));
 sg13g2_a221oi_1 _27840_ (.B2(_08932_),
    .C1(_08936_),
    .B1(_08914_),
    .A1(net100),
    .Y(_02719_),
    .A2(net72));
 sg13g2_a221oi_1 _27841_ (.B2(\stack[31][5] ),
    .C1(net72),
    .B1(_08914_),
    .A1(net1221),
    .Y(_08937_),
    .A2(net489));
 sg13g2_a21o_1 _27842_ (.A2(_08919_),
    .A1(net90),
    .B1(_08937_),
    .X(_08938_));
 sg13g2_o21ai_1 _27843_ (.B1(_08938_),
    .Y(_02720_),
    .A1(net446),
    .A2(_08933_));
 sg13g2_nand2_1 _27844_ (.Y(_08939_),
    .A(_10017_),
    .B(_08911_));
 sg13g2_a21oi_1 _27845_ (.A1(net127),
    .A2(_08223_),
    .Y(_08940_),
    .B1(_08939_));
 sg13g2_a221oi_1 _27846_ (.B2(net483),
    .C1(_08940_),
    .B1(net109),
    .A1(_08263_),
    .Y(_08941_),
    .A2(_08918_));
 sg13g2_inv_1 _27847_ (.Y(_08942_),
    .A(\stack[31][6] ));
 sg13g2_mux2_1 _27848_ (.A0(_08941_),
    .A1(_08942_),
    .S(_08914_),
    .X(_08943_));
 sg13g2_and2_1 _27849_ (.A(_08919_),
    .B(_08941_),
    .X(_08944_));
 sg13g2_a22oi_1 _27850_ (.Y(_02721_),
    .B1(_08944_),
    .B2(_08169_),
    .A2(_08943_),
    .A1(_08909_));
 sg13g2_nand3b_1 _27851_ (.B(\stack[31][7] ),
    .C(_10415_),
    .Y(_08945_),
    .A_N(net489));
 sg13g2_nand2_1 _27852_ (.Y(_08946_),
    .A(net1213),
    .B(net489));
 sg13g2_o21ai_1 _27853_ (.B1(_08946_),
    .Y(_08947_),
    .A1(net109),
    .A2(_08945_));
 sg13g2_a22oi_1 _27854_ (.Y(_08948_),
    .B1(_08947_),
    .B2(_08909_),
    .A2(net109),
    .A1(net298));
 sg13g2_o21ai_1 _27855_ (.B1(_08948_),
    .Y(_02722_),
    .A1(net41),
    .A2(_08909_));
 sg13g2_nor2_1 _27856_ (.A(net141),
    .B(net126),
    .Y(_08949_));
 sg13g2_and2_1 _27857_ (.A(_08461_),
    .B(_08949_),
    .X(_08950_));
 sg13g2_buf_2 _27858_ (.A(_08950_),
    .X(_08951_));
 sg13g2_buf_1 _27859_ (.A(_08951_),
    .X(_08952_));
 sg13g2_nor2_1 _27860_ (.A(_07594_),
    .B(_08017_),
    .Y(_08953_));
 sg13g2_buf_1 _27861_ (.A(_08953_),
    .X(_08954_));
 sg13g2_nand4_1 _27862_ (.B(_07558_),
    .C(_07952_),
    .A(_07607_),
    .Y(_08955_),
    .D(_08011_));
 sg13g2_buf_1 _27863_ (.A(_08955_),
    .X(_08956_));
 sg13g2_and2_1 _27864_ (.A(_09906_),
    .B(_08956_),
    .X(_08957_));
 sg13g2_buf_1 _27865_ (.A(_08957_),
    .X(_08958_));
 sg13g2_nor2b_1 _27866_ (.A(_08953_),
    .B_N(_08958_),
    .Y(_08959_));
 sg13g2_buf_2 _27867_ (.A(_08959_),
    .X(_08960_));
 sg13g2_a22oi_1 _27868_ (.Y(_08961_),
    .B1(_08960_),
    .B2(\stack[3][0] ),
    .A2(net488),
    .A1(net1226));
 sg13g2_nor3_1 _27869_ (.A(_07531_),
    .B(_08036_),
    .C(_08360_),
    .Y(_08962_));
 sg13g2_buf_1 _27870_ (.A(_08962_),
    .X(_08963_));
 sg13g2_a22oi_1 _27871_ (.Y(_08964_),
    .B1(net51),
    .B2(net131),
    .A2(_08963_),
    .A1(net478));
 sg13g2_o21ai_1 _27872_ (.B1(_08964_),
    .Y(_02723_),
    .A1(net51),
    .A2(_08961_));
 sg13g2_a22oi_1 _27873_ (.Y(_08965_),
    .B1(_08960_),
    .B2(\stack[3][1] ),
    .A2(net488),
    .A1(net1212));
 sg13g2_a22oi_1 _27874_ (.Y(_08966_),
    .B1(net51),
    .B2(net105),
    .A2(_08963_),
    .A1(_10098_));
 sg13g2_o21ai_1 _27875_ (.B1(_08966_),
    .Y(_02724_),
    .A1(net51),
    .A2(_08965_));
 sg13g2_a22oi_1 _27876_ (.Y(_08967_),
    .B1(_08960_),
    .B2(\stack[3][2] ),
    .A2(net488),
    .A1(net1217));
 sg13g2_a22oi_1 _27877_ (.Y(_08968_),
    .B1(_08952_),
    .B2(net104),
    .A2(_08963_),
    .A1(net452));
 sg13g2_o21ai_1 _27878_ (.B1(_08968_),
    .Y(_02725_),
    .A1(net51),
    .A2(_08967_));
 sg13g2_a22oi_1 _27879_ (.Y(_08969_),
    .B1(_08960_),
    .B2(\stack[3][3] ),
    .A2(_08954_),
    .A1(net1211));
 sg13g2_a22oi_1 _27880_ (.Y(_08970_),
    .B1(_08952_),
    .B2(net91),
    .A2(_08963_),
    .A1(_07745_));
 sg13g2_o21ai_1 _27881_ (.B1(_08970_),
    .Y(_02726_),
    .A1(net51),
    .A2(_08969_));
 sg13g2_and2_1 _27882_ (.A(net98),
    .B(_08951_),
    .X(_08971_));
 sg13g2_a221oi_1 _27883_ (.B2(\stack[3][4] ),
    .C1(_08951_),
    .B1(_08960_),
    .A1(_07787_),
    .Y(_08972_),
    .A2(_08954_));
 sg13g2_nand2_1 _27884_ (.Y(_08973_),
    .A(_08336_),
    .B(_08963_));
 sg13g2_o21ai_1 _27885_ (.B1(_08973_),
    .Y(_02727_),
    .A1(_08971_),
    .A2(_08972_));
 sg13g2_nor2b_1 _27886_ (.A(net488),
    .B_N(\stack[3][5] ),
    .Y(_08974_));
 sg13g2_a22oi_1 _27887_ (.Y(_08975_),
    .B1(_08974_),
    .B2(_08958_),
    .A2(net488),
    .A1(net1214));
 sg13g2_mux2_1 _27888_ (.A0(_08975_),
    .A1(net90),
    .S(_08951_),
    .X(_08976_));
 sg13g2_o21ai_1 _27889_ (.B1(_08976_),
    .Y(_02728_),
    .A1(net446),
    .A2(_08956_));
 sg13g2_nor2b_1 _27890_ (.A(net488),
    .B_N(\stack[3][6] ),
    .Y(_08977_));
 sg13g2_a22oi_1 _27891_ (.Y(_08978_),
    .B1(_08977_),
    .B2(_08958_),
    .A2(net488),
    .A1(net879));
 sg13g2_a22oi_1 _27892_ (.Y(_08979_),
    .B1(_08951_),
    .B2(net46),
    .A2(_08963_),
    .A1(net449));
 sg13g2_o21ai_1 _27893_ (.B1(_08979_),
    .Y(_02729_),
    .A1(net51),
    .A2(_08978_));
 sg13g2_nand2_1 _27894_ (.Y(_08980_),
    .A(net1213),
    .B(net488));
 sg13g2_o21ai_1 _27895_ (.B1(_08980_),
    .Y(_08981_),
    .A1(_10138_),
    .A2(_08956_));
 sg13g2_a221oi_1 _27896_ (.B2(\stack[3][7] ),
    .C1(_08981_),
    .B1(_08960_),
    .A1(_08461_),
    .Y(_08982_),
    .A2(_08949_));
 sg13g2_a21oi_1 _27897_ (.A1(net43),
    .A2(net51),
    .Y(_02730_),
    .B1(_08982_));
 sg13g2_nor2b_1 _27898_ (.A(net141),
    .B_N(_07585_),
    .Y(_08983_));
 sg13g2_and2_1 _27899_ (.A(_08461_),
    .B(_08983_),
    .X(_08984_));
 sg13g2_buf_1 _27900_ (.A(_08984_),
    .X(_08985_));
 sg13g2_nand2_2 _27901_ (.Y(_08986_),
    .A(_07476_),
    .B(_08449_));
 sg13g2_nor2_1 _27902_ (.A(_08302_),
    .B(_08986_),
    .Y(_08987_));
 sg13g2_buf_2 _27903_ (.A(_08987_),
    .X(_08988_));
 sg13g2_nor4_2 _27904_ (.A(_07746_),
    .B(net139),
    .C(net125),
    .Y(_08989_),
    .D(net296));
 sg13g2_nor2_1 _27905_ (.A(_08390_),
    .B(_08989_),
    .Y(_08990_));
 sg13g2_buf_2 _27906_ (.A(_08990_),
    .X(_08991_));
 sg13g2_or2_1 _27907_ (.X(_08992_),
    .B(_08986_),
    .A(net521));
 sg13g2_buf_2 _27908_ (.A(_08992_),
    .X(_08993_));
 sg13g2_and2_1 _27909_ (.A(\stack[4][0] ),
    .B(_08993_),
    .X(_08994_));
 sg13g2_a22oi_1 _27910_ (.Y(_08995_),
    .B1(_08991_),
    .B2(_08994_),
    .A2(_08988_),
    .A1(_07591_));
 sg13g2_nor4_2 _27911_ (.A(_07746_),
    .B(_07751_),
    .C(net129),
    .Y(_08996_),
    .D(net122));
 sg13g2_a22oi_1 _27912_ (.Y(_08997_),
    .B1(_08996_),
    .B2(net453),
    .A2(net71),
    .A1(_07665_));
 sg13g2_o21ai_1 _27913_ (.B1(_08997_),
    .Y(_02731_),
    .A1(net71),
    .A2(_08995_));
 sg13g2_and2_1 _27914_ (.A(\stack[4][1] ),
    .B(_08993_),
    .X(_08998_));
 sg13g2_a22oi_1 _27915_ (.Y(_08999_),
    .B1(_08991_),
    .B2(_08998_),
    .A2(_08988_),
    .A1(net1212));
 sg13g2_a22oi_1 _27916_ (.Y(_09000_),
    .B1(_08996_),
    .B2(net295),
    .A2(net71),
    .A1(net113));
 sg13g2_o21ai_1 _27917_ (.B1(_09000_),
    .Y(_02732_),
    .A1(_08985_),
    .A2(_08999_));
 sg13g2_and2_1 _27918_ (.A(\stack[4][2] ),
    .B(_08993_),
    .X(_09001_));
 sg13g2_a22oi_1 _27919_ (.Y(_09002_),
    .B1(_08991_),
    .B2(_09001_),
    .A2(_08988_),
    .A1(net1217));
 sg13g2_a22oi_1 _27920_ (.Y(_09003_),
    .B1(_08996_),
    .B2(net400),
    .A2(net71),
    .A1(net112));
 sg13g2_o21ai_1 _27921_ (.B1(_09003_),
    .Y(_02733_),
    .A1(net71),
    .A2(_09002_));
 sg13g2_and2_1 _27922_ (.A(\stack[4][3] ),
    .B(_08993_),
    .X(_09004_));
 sg13g2_a22oi_1 _27923_ (.Y(_09005_),
    .B1(_08991_),
    .B2(_09004_),
    .A2(_08988_),
    .A1(net1211));
 sg13g2_a22oi_1 _27924_ (.Y(_09006_),
    .B1(_08996_),
    .B2(net477),
    .A2(net71),
    .A1(net101));
 sg13g2_o21ai_1 _27925_ (.B1(_09006_),
    .Y(_02734_),
    .A1(net71),
    .A2(_09005_));
 sg13g2_nand3_1 _27926_ (.B(net299),
    .C(_08382_),
    .A(_07621_),
    .Y(_09007_));
 sg13g2_buf_1 _27927_ (.A(_09007_),
    .X(_09008_));
 sg13g2_and2_1 _27928_ (.A(\stack[4][4] ),
    .B(_08993_),
    .X(_09009_));
 sg13g2_a22oi_1 _27929_ (.Y(_09010_),
    .B1(_08991_),
    .B2(_09009_),
    .A2(_08988_),
    .A1(_08117_));
 sg13g2_nand2_2 _27930_ (.Y(_09011_),
    .A(_08461_),
    .B(_08983_));
 sg13g2_mux2_1 _27931_ (.A0(_08115_),
    .A1(_09010_),
    .S(_09011_),
    .X(_09012_));
 sg13g2_o21ai_1 _27932_ (.B1(_09012_),
    .Y(_02735_),
    .A1(net496),
    .A2(_09008_));
 sg13g2_and2_1 _27933_ (.A(\stack[4][5] ),
    .B(_08993_),
    .X(_09013_));
 sg13g2_a22oi_1 _27934_ (.Y(_09014_),
    .B1(_08991_),
    .B2(_09013_),
    .A2(_08988_),
    .A1(_08062_));
 sg13g2_mux2_1 _27935_ (.A0(net90),
    .A1(_09014_),
    .S(_09011_),
    .X(_09015_));
 sg13g2_o21ai_1 _27936_ (.B1(_09015_),
    .Y(_02736_),
    .A1(_10128_),
    .A2(_09008_));
 sg13g2_nor2_1 _27937_ (.A(_08068_),
    .B(_09011_),
    .Y(_09016_));
 sg13g2_nand4_1 _27938_ (.B(\stack[4][6] ),
    .C(_08993_),
    .A(_09995_),
    .Y(_09017_),
    .D(_09008_));
 sg13g2_a22oi_1 _27939_ (.Y(_09018_),
    .B1(_08989_),
    .B2(_07856_),
    .A2(_08988_),
    .A1(net1220));
 sg13g2_nand3_1 _27940_ (.B(_09017_),
    .C(_09018_),
    .A(_09011_),
    .Y(_09019_));
 sg13g2_nor2b_1 _27941_ (.A(_09016_),
    .B_N(_09019_),
    .Y(_02737_));
 sg13g2_nand4_1 _27942_ (.B(\stack[4][7] ),
    .C(_08993_),
    .A(_09995_),
    .Y(_09020_),
    .D(_09008_));
 sg13g2_a22oi_1 _27943_ (.Y(_09021_),
    .B1(_08989_),
    .B2(_08347_),
    .A2(_08988_),
    .A1(_07930_));
 sg13g2_and3_1 _27944_ (.X(_09022_),
    .A(_09011_),
    .B(_09020_),
    .C(_09021_));
 sg13g2_a21oi_1 _27945_ (.A1(net43),
    .A2(net71),
    .Y(_02738_),
    .B1(_09022_));
 sg13g2_nor4_1 _27946_ (.A(net140),
    .B(net141),
    .C(_08029_),
    .D(net122),
    .Y(_09023_));
 sg13g2_buf_2 _27947_ (.A(_09023_),
    .X(_09024_));
 sg13g2_buf_1 _27948_ (.A(_09024_),
    .X(_09025_));
 sg13g2_nor2_1 _27949_ (.A(_08133_),
    .B(_08986_),
    .Y(_09026_));
 sg13g2_buf_1 _27950_ (.A(_09026_),
    .X(_09027_));
 sg13g2_nor4_1 _27951_ (.A(_07604_),
    .B(_07546_),
    .C(_07610_),
    .D(_08035_),
    .Y(_09028_));
 sg13g2_buf_1 _27952_ (.A(_09028_),
    .X(_09029_));
 sg13g2_nor2_1 _27953_ (.A(_08390_),
    .B(_09029_),
    .Y(_09030_));
 sg13g2_nor2b_1 _27954_ (.A(net501),
    .B_N(\stack[5][0] ),
    .Y(_09031_));
 sg13g2_a22oi_1 _27955_ (.Y(_09032_),
    .B1(_09030_),
    .B2(_09031_),
    .A2(net501),
    .A1(_07591_));
 sg13g2_a22oi_1 _27956_ (.Y(_09033_),
    .B1(net70),
    .B2(net131),
    .A2(net108),
    .A1(_07960_));
 sg13g2_o21ai_1 _27957_ (.B1(_09033_),
    .Y(_02739_),
    .A1(net70),
    .A2(_09032_));
 sg13g2_nor3_1 _27958_ (.A(net1191),
    .B(net108),
    .C(_09026_),
    .Y(_09034_));
 sg13g2_buf_2 _27959_ (.A(_09034_),
    .X(_09035_));
 sg13g2_a22oi_1 _27960_ (.Y(_09036_),
    .B1(_09035_),
    .B2(\stack[5][1] ),
    .A2(_09027_),
    .A1(net1212));
 sg13g2_a22oi_1 _27961_ (.Y(_09037_),
    .B1(net70),
    .B2(net105),
    .A2(net108),
    .A1(_10098_));
 sg13g2_o21ai_1 _27962_ (.B1(_09037_),
    .Y(_02740_),
    .A1(_09025_),
    .A2(_09036_));
 sg13g2_a22oi_1 _27963_ (.Y(_09038_),
    .B1(_09035_),
    .B2(\stack[5][2] ),
    .A2(_09027_),
    .A1(net1217));
 sg13g2_a22oi_1 _27964_ (.Y(_09039_),
    .B1(_09025_),
    .B2(net104),
    .A2(net108),
    .A1(_07707_));
 sg13g2_o21ai_1 _27965_ (.B1(_09039_),
    .Y(_02741_),
    .A1(net70),
    .A2(_09038_));
 sg13g2_a22oi_1 _27966_ (.Y(_09040_),
    .B1(_09035_),
    .B2(\stack[5][3] ),
    .A2(net501),
    .A1(net1211));
 sg13g2_a22oi_1 _27967_ (.Y(_09041_),
    .B1(_09024_),
    .B2(net91),
    .A2(net108),
    .A1(net492));
 sg13g2_o21ai_1 _27968_ (.B1(_09041_),
    .Y(_02742_),
    .A1(net70),
    .A2(_09040_));
 sg13g2_and2_1 _27969_ (.A(_08115_),
    .B(_09024_),
    .X(_09042_));
 sg13g2_a221oi_1 _27970_ (.B2(\stack[5][4] ),
    .C1(_09024_),
    .B1(_09035_),
    .A1(_07787_),
    .Y(_09043_),
    .A2(net501));
 sg13g2_nand2_1 _27971_ (.Y(_09044_),
    .A(net476),
    .B(net108));
 sg13g2_o21ai_1 _27972_ (.B1(_09044_),
    .Y(_02743_),
    .A1(_09042_),
    .A2(_09043_));
 sg13g2_and2_1 _27973_ (.A(_07848_),
    .B(_09024_),
    .X(_09045_));
 sg13g2_a221oi_1 _27974_ (.B2(\stack[5][5] ),
    .C1(_09024_),
    .B1(_09035_),
    .A1(_08062_),
    .Y(_09046_),
    .A2(net501));
 sg13g2_nand2_1 _27975_ (.Y(_09047_),
    .A(_08121_),
    .B(net108));
 sg13g2_o21ai_1 _27976_ (.B1(_09047_),
    .Y(_02744_),
    .A1(_09045_),
    .A2(_09046_));
 sg13g2_nor2b_1 _27977_ (.A(net501),
    .B_N(\stack[5][6] ),
    .Y(_09048_));
 sg13g2_a22oi_1 _27978_ (.Y(_09049_),
    .B1(_09030_),
    .B2(_09048_),
    .A2(net501),
    .A1(_07998_));
 sg13g2_a22oi_1 _27979_ (.Y(_09050_),
    .B1(_09024_),
    .B2(net46),
    .A2(_09029_),
    .A1(net449));
 sg13g2_o21ai_1 _27980_ (.B1(_09050_),
    .Y(_02745_),
    .A1(net70),
    .A2(_09049_));
 sg13g2_and2_1 _27981_ (.A(net474),
    .B(net108),
    .X(_09051_));
 sg13g2_a221oi_1 _27982_ (.B2(\stack[5][7] ),
    .C1(_09051_),
    .B1(_09035_),
    .A1(net1213),
    .Y(_09052_),
    .A2(net501));
 sg13g2_nor2b_1 _27983_ (.A(net70),
    .B_N(_09052_),
    .Y(_09053_));
 sg13g2_a21oi_1 _27984_ (.A1(_08003_),
    .A2(net70),
    .Y(_02746_),
    .B1(_09053_));
 sg13g2_and2_1 _27985_ (.A(_07938_),
    .B(_08382_),
    .X(_09054_));
 sg13g2_buf_1 _27986_ (.A(_09054_),
    .X(_09055_));
 sg13g2_buf_1 _27987_ (.A(_09055_),
    .X(_09056_));
 sg13g2_nor2_1 _27988_ (.A(net532),
    .B(_08986_),
    .Y(_09057_));
 sg13g2_buf_1 _27989_ (.A(_09057_),
    .X(_09058_));
 sg13g2_nand4_1 _27990_ (.B(net125),
    .C(net299),
    .A(net139),
    .Y(_09059_),
    .D(_08008_));
 sg13g2_buf_1 _27991_ (.A(_09059_),
    .X(_09060_));
 sg13g2_and2_1 _27992_ (.A(_09984_),
    .B(_09060_),
    .X(_09061_));
 sg13g2_nor2b_1 _27993_ (.A(net514),
    .B_N(\stack[6][0] ),
    .Y(_09062_));
 sg13g2_a22oi_1 _27994_ (.Y(_09063_),
    .B1(_09061_),
    .B2(_09062_),
    .A2(net514),
    .A1(net1226));
 sg13g2_nor3_1 _27995_ (.A(_07755_),
    .B(_08533_),
    .C(_07971_),
    .Y(_09064_));
 sg13g2_buf_2 _27996_ (.A(_09064_),
    .X(_09065_));
 sg13g2_a22oi_1 _27997_ (.Y(_09066_),
    .B1(_09065_),
    .B2(net453),
    .A2(net50),
    .A1(_07665_));
 sg13g2_o21ai_1 _27998_ (.B1(_09066_),
    .Y(_02747_),
    .A1(net50),
    .A2(_09063_));
 sg13g2_inv_1 _27999_ (.Y(_09067_),
    .A(net514));
 sg13g2_and3_1 _28000_ (.X(_09068_),
    .A(_09908_),
    .B(_09067_),
    .C(_09060_));
 sg13g2_buf_2 _28001_ (.A(_09068_),
    .X(_09069_));
 sg13g2_a22oi_1 _28002_ (.Y(_09070_),
    .B1(_09069_),
    .B2(\stack[6][1] ),
    .A2(net514),
    .A1(_08100_));
 sg13g2_a22oi_1 _28003_ (.Y(_09071_),
    .B1(_09065_),
    .B2(net295),
    .A2(net50),
    .A1(_08531_));
 sg13g2_o21ai_1 _28004_ (.B1(_09071_),
    .Y(_02748_),
    .A1(_09056_),
    .A2(_09070_));
 sg13g2_a22oi_1 _28005_ (.Y(_09072_),
    .B1(_09069_),
    .B2(\stack[6][2] ),
    .A2(net514),
    .A1(_07976_));
 sg13g2_a22oi_1 _28006_ (.Y(_09073_),
    .B1(_09065_),
    .B2(net400),
    .A2(net50),
    .A1(_08537_));
 sg13g2_o21ai_1 _28007_ (.B1(_09073_),
    .Y(_02749_),
    .A1(net50),
    .A2(_09072_));
 sg13g2_a22oi_1 _28008_ (.Y(_09074_),
    .B1(_09069_),
    .B2(\stack[6][3] ),
    .A2(_09058_),
    .A1(_08111_));
 sg13g2_a22oi_1 _28009_ (.Y(_09075_),
    .B1(_09065_),
    .B2(_08300_),
    .A2(_09056_),
    .A1(_07981_));
 sg13g2_o21ai_1 _28010_ (.B1(_09075_),
    .Y(_02750_),
    .A1(net50),
    .A2(_09074_));
 sg13g2_nor2b_1 _28011_ (.A(net514),
    .B_N(\stack[6][4] ),
    .Y(_09076_));
 sg13g2_a221oi_1 _28012_ (.B2(_09076_),
    .C1(_09055_),
    .B1(_09061_),
    .A1(net1209),
    .Y(_09077_),
    .A2(net514));
 sg13g2_a21o_1 _28013_ (.A2(net50),
    .A1(net98),
    .B1(_09077_),
    .X(_09078_));
 sg13g2_o21ai_1 _28014_ (.B1(_09078_),
    .Y(_02751_),
    .A1(_10118_),
    .A2(_09060_));
 sg13g2_a221oi_1 _28015_ (.B2(\stack[6][5] ),
    .C1(_09055_),
    .B1(_09069_),
    .A1(net1221),
    .Y(_09079_),
    .A2(net514));
 sg13g2_a21oi_1 _28016_ (.A1(net90),
    .A2(net50),
    .Y(_09080_),
    .B1(_09079_));
 sg13g2_a21o_1 _28017_ (.A2(_09065_),
    .A1(_08060_),
    .B1(_09080_),
    .X(_02752_));
 sg13g2_a22oi_1 _28018_ (.Y(_09081_),
    .B1(_09069_),
    .B2(\stack[6][6] ),
    .A2(_09065_),
    .A1(net451));
 sg13g2_o21ai_1 _28019_ (.B1(_09081_),
    .Y(_09082_),
    .A1(_10018_),
    .A2(_09067_));
 sg13g2_nand2_1 _28020_ (.Y(_09083_),
    .A(_07938_),
    .B(_08382_));
 sg13g2_mux2_1 _28021_ (.A0(_08068_),
    .A1(_09082_),
    .S(_09083_),
    .X(_02753_));
 sg13g2_nor2_1 _28022_ (.A(_10025_),
    .B(_09067_),
    .Y(_09084_));
 sg13g2_a21o_1 _28023_ (.A2(_09069_),
    .A1(\stack[6][7] ),
    .B1(_09084_),
    .X(_09085_));
 sg13g2_a22oi_1 _28024_ (.Y(_09086_),
    .B1(_09085_),
    .B2(_09083_),
    .A2(_09065_),
    .A1(net298));
 sg13g2_o21ai_1 _28025_ (.B1(_09086_),
    .Y(_02754_),
    .A1(net41),
    .A2(_09083_));
 sg13g2_nor2_1 _28026_ (.A(_08016_),
    .B(_08986_),
    .Y(_09087_));
 sg13g2_buf_1 _28027_ (.A(_09087_),
    .X(_09088_));
 sg13g2_and4_1 _28028_ (.A(_07546_),
    .B(net135),
    .C(_07952_),
    .D(_08012_),
    .X(_09089_));
 sg13g2_buf_1 _28029_ (.A(_09089_),
    .X(_09090_));
 sg13g2_nor3_1 _28030_ (.A(_10144_),
    .B(net500),
    .C(net107),
    .Y(_09091_));
 sg13g2_buf_1 _28031_ (.A(_09091_),
    .X(_09092_));
 sg13g2_a21oi_1 _28032_ (.A1(_07961_),
    .A2(net500),
    .Y(_09093_),
    .B1(net69));
 sg13g2_nor3_1 _28033_ (.A(net141),
    .B(_08029_),
    .C(_08556_),
    .Y(_09094_));
 sg13g2_buf_2 _28034_ (.A(_09094_),
    .X(_09095_));
 sg13g2_mux2_1 _28035_ (.A0(_09093_),
    .A1(net123),
    .S(_09095_),
    .X(_09096_));
 sg13g2_nand2_1 _28036_ (.Y(_09097_),
    .A(_07620_),
    .B(net107));
 sg13g2_buf_8 _28037_ (.A(_09095_),
    .X(_09098_));
 sg13g2_nor2_1 _28038_ (.A(\stack[7][0] ),
    .B(net49),
    .Y(_09099_));
 sg13g2_a22oi_1 _28039_ (.Y(_02755_),
    .B1(_09099_),
    .B2(_09092_),
    .A2(_09097_),
    .A1(_09096_));
 sg13g2_a22oi_1 _28040_ (.Y(_09100_),
    .B1(net69),
    .B2(\stack[7][1] ),
    .A2(net500),
    .A1(_08100_));
 sg13g2_a22oi_1 _28041_ (.Y(_09101_),
    .B1(net107),
    .B2(net295),
    .A2(net49),
    .A1(_08531_));
 sg13g2_o21ai_1 _28042_ (.B1(_09101_),
    .Y(_02756_),
    .A1(_09098_),
    .A2(_09100_));
 sg13g2_a22oi_1 _28043_ (.Y(_09102_),
    .B1(net69),
    .B2(\stack[7][2] ),
    .A2(net500),
    .A1(_07976_));
 sg13g2_a22oi_1 _28044_ (.Y(_09103_),
    .B1(net107),
    .B2(net400),
    .A2(net49),
    .A1(_08537_));
 sg13g2_o21ai_1 _28045_ (.B1(_09103_),
    .Y(_02757_),
    .A1(net49),
    .A2(_09102_));
 sg13g2_a22oi_1 _28046_ (.Y(_09104_),
    .B1(net69),
    .B2(\stack[7][3] ),
    .A2(_09088_),
    .A1(_08111_));
 sg13g2_a22oi_1 _28047_ (.Y(_09105_),
    .B1(_09090_),
    .B2(_08300_),
    .A2(net49),
    .A1(_07981_));
 sg13g2_o21ai_1 _28048_ (.B1(_09105_),
    .Y(_02758_),
    .A1(_09098_),
    .A2(_09104_));
 sg13g2_a221oi_1 _28049_ (.B2(\stack[7][4] ),
    .C1(_09095_),
    .B1(net69),
    .A1(_08158_),
    .Y(_09106_),
    .A2(net500));
 sg13g2_a21oi_1 _28050_ (.A1(net102),
    .A2(_09095_),
    .Y(_09107_),
    .B1(_09106_));
 sg13g2_a21o_1 _28051_ (.A2(net107),
    .A1(_08336_),
    .B1(_09107_),
    .X(_02759_));
 sg13g2_a221oi_1 _28052_ (.B2(\stack[7][5] ),
    .C1(_09095_),
    .B1(net69),
    .A1(net1221),
    .Y(_09108_),
    .A2(net500));
 sg13g2_a21oi_1 _28053_ (.A1(net90),
    .A2(_09095_),
    .Y(_09109_),
    .B1(_09108_));
 sg13g2_a21o_1 _28054_ (.A2(net107),
    .A1(net403),
    .B1(_09109_),
    .X(_02760_));
 sg13g2_a22oi_1 _28055_ (.Y(_09110_),
    .B1(net69),
    .B2(\stack[7][6] ),
    .A2(net500),
    .A1(_07998_));
 sg13g2_a22oi_1 _28056_ (.Y(_09111_),
    .B1(net107),
    .B2(net405),
    .A2(_09095_),
    .A1(_07899_));
 sg13g2_o21ai_1 _28057_ (.B1(_09111_),
    .Y(_02761_),
    .A1(net49),
    .A2(_09110_));
 sg13g2_and2_1 _28058_ (.A(_09660_),
    .B(net107),
    .X(_09112_));
 sg13g2_a221oi_1 _28059_ (.B2(\stack[7][7] ),
    .C1(_09112_),
    .B1(net69),
    .A1(net1213),
    .Y(_09113_),
    .A2(net500));
 sg13g2_nor2b_1 _28060_ (.A(net49),
    .B_N(_09113_),
    .Y(_09114_));
 sg13g2_a21oi_1 _28061_ (.A1(_08003_),
    .A2(net49),
    .Y(_02762_),
    .B1(_09114_));
 sg13g2_inv_1 _28062_ (.Y(_09115_),
    .A(\stack[8][0] ));
 sg13g2_a21o_1 _28063_ (.A2(net299),
    .A1(_07621_),
    .B1(_08102_),
    .X(_09116_));
 sg13g2_o21ai_1 _28064_ (.B1(net1304),
    .Y(_09117_),
    .A1(net521),
    .A2(_07942_));
 sg13g2_a21oi_1 _28065_ (.A1(_07936_),
    .A2(_09116_),
    .Y(_09118_),
    .B1(_09117_));
 sg13g2_buf_1 _28066_ (.A(_09118_),
    .X(_09119_));
 sg13g2_and4_1 _28067_ (.A(net139),
    .B(net125),
    .C(net127),
    .D(net137),
    .X(_09120_));
 sg13g2_buf_1 _28068_ (.A(_09120_),
    .X(_09121_));
 sg13g2_nand2_1 _28069_ (.Y(_09122_),
    .A(net123),
    .B(net95));
 sg13g2_nor2_1 _28070_ (.A(net521),
    .B(_07942_),
    .Y(_09123_));
 sg13g2_buf_1 _28071_ (.A(_09123_),
    .X(_09124_));
 sg13g2_a21o_1 _28072_ (.A2(_09124_),
    .A1(net1208),
    .B1(net95),
    .X(_09125_));
 sg13g2_nor4_1 _28073_ (.A(net130),
    .B(net491),
    .C(_07754_),
    .D(net121),
    .Y(_09126_));
 sg13g2_buf_1 _28074_ (.A(_09126_),
    .X(_09127_));
 sg13g2_a221oi_1 _28075_ (.B2(net478),
    .C1(net48),
    .B1(net94),
    .A1(_09122_),
    .Y(_09128_),
    .A2(_09125_));
 sg13g2_a21oi_1 _28076_ (.A1(_09115_),
    .A2(net48),
    .Y(_02763_),
    .B1(_09128_));
 sg13g2_nand2_2 _28077_ (.Y(_09129_),
    .A(_07936_),
    .B(_08102_));
 sg13g2_nand3_1 _28078_ (.B(_09124_),
    .C(_09129_),
    .A(net1212),
    .Y(_09130_));
 sg13g2_a22oi_1 _28079_ (.Y(_09131_),
    .B1(net94),
    .B2(net402),
    .A2(net95),
    .A1(net119));
 sg13g2_nand2_1 _28080_ (.Y(_09132_),
    .A(_09130_),
    .B(_09131_));
 sg13g2_mux2_1 _28081_ (.A0(_09132_),
    .A1(\stack[8][1] ),
    .S(net48),
    .X(_02764_));
 sg13g2_nand3_1 _28082_ (.B(_09124_),
    .C(_09129_),
    .A(net1217),
    .Y(_09133_));
 sg13g2_a22oi_1 _28083_ (.Y(_09134_),
    .B1(net94),
    .B2(net450),
    .A2(net95),
    .A1(net118));
 sg13g2_nand2_1 _28084_ (.Y(_09135_),
    .A(_09133_),
    .B(_09134_));
 sg13g2_mux2_1 _28085_ (.A0(_09135_),
    .A1(\stack[8][2] ),
    .S(net48),
    .X(_02765_));
 sg13g2_nand2_1 _28086_ (.Y(_09136_),
    .A(net1211),
    .B(_09124_));
 sg13g2_a22oi_1 _28087_ (.Y(_09137_),
    .B1(net94),
    .B2(net510),
    .A2(net95),
    .A1(net103));
 sg13g2_o21ai_1 _28088_ (.B1(_09137_),
    .Y(_09138_),
    .A1(net95),
    .A2(_09136_));
 sg13g2_mux2_1 _28089_ (.A0(_09138_),
    .A1(\stack[8][3] ),
    .S(net48),
    .X(_02766_));
 sg13g2_nor2b_1 _28090_ (.A(net95),
    .B_N(_09124_),
    .Y(_09139_));
 sg13g2_and2_1 _28091_ (.A(net1210),
    .B(_09139_),
    .X(_09140_));
 sg13g2_a221oi_1 _28092_ (.B2(net484),
    .C1(_09140_),
    .B1(net94),
    .A1(\stack[8][4] ),
    .Y(_09141_),
    .A2(net48));
 sg13g2_o21ai_1 _28093_ (.B1(_09141_),
    .Y(_02767_),
    .A1(net100),
    .A2(_09129_));
 sg13g2_inv_1 _28094_ (.Y(_09142_),
    .A(\stack[8][5] ));
 sg13g2_nand2_1 _28095_ (.Y(_09143_),
    .A(net1298),
    .B(_09124_));
 sg13g2_o21ai_1 _28096_ (.B1(_09143_),
    .Y(_09144_),
    .A1(_09117_),
    .A2(net94));
 sg13g2_a221oi_1 _28097_ (.B2(net401),
    .C1(_09144_),
    .B1(_09127_),
    .A1(_07936_),
    .Y(_09145_),
    .A2(_08102_));
 sg13g2_a221oi_1 _28098_ (.B2(net89),
    .C1(_09145_),
    .B1(net95),
    .A1(_09142_),
    .Y(_02768_),
    .A2(net48));
 sg13g2_inv_1 _28099_ (.Y(_09146_),
    .A(\stack[8][6] ));
 sg13g2_nand2_1 _28100_ (.Y(_09147_),
    .A(net42),
    .B(_09121_));
 sg13g2_nor3_1 _28101_ (.A(_10018_),
    .B(net521),
    .C(_07942_),
    .Y(_09148_));
 sg13g2_a221oi_1 _28102_ (.B2(_09129_),
    .C1(_09119_),
    .B1(_09148_),
    .A1(net449),
    .Y(_09149_),
    .A2(net94));
 sg13g2_a22oi_1 _28103_ (.Y(_02769_),
    .B1(_09147_),
    .B2(_09149_),
    .A2(net48),
    .A1(_09146_));
 sg13g2_and2_1 _28104_ (.A(net1219),
    .B(_09139_),
    .X(_09150_));
 sg13g2_a221oi_1 _28105_ (.B2(net298),
    .C1(_09150_),
    .B1(net94),
    .A1(\stack[8][7] ),
    .Y(_09151_),
    .A2(_09119_));
 sg13g2_o21ai_1 _28106_ (.B1(_09151_),
    .Y(_02770_),
    .A1(net41),
    .A2(_09129_));
 sg13g2_nor3_1 _28107_ (.A(net130),
    .B(net121),
    .C(_08028_),
    .Y(_09152_));
 sg13g2_buf_2 _28108_ (.A(_09152_),
    .X(_09153_));
 sg13g2_or4_1 _28109_ (.A(_07604_),
    .B(net136),
    .C(_07558_),
    .D(net297),
    .X(_09154_));
 sg13g2_nor2_1 _28110_ (.A(_07942_),
    .B(net522),
    .Y(_09155_));
 sg13g2_buf_1 _28111_ (.A(_09155_),
    .X(_09156_));
 sg13g2_nor2_1 _28112_ (.A(net1270),
    .B(net499),
    .Y(_09157_));
 sg13g2_and2_1 _28113_ (.A(_09154_),
    .B(_09157_),
    .X(_09158_));
 sg13g2_buf_1 _28114_ (.A(_09158_),
    .X(_09159_));
 sg13g2_nand2b_1 _28115_ (.Y(_09160_),
    .B(_09159_),
    .A_N(_09153_));
 sg13g2_buf_1 _28116_ (.A(_09160_),
    .X(_09161_));
 sg13g2_buf_1 _28117_ (.A(_09153_),
    .X(_09162_));
 sg13g2_nor3_1 _28118_ (.A(net130),
    .B(net121),
    .C(net297),
    .Y(_09163_));
 sg13g2_buf_2 _28119_ (.A(_09163_),
    .X(_09164_));
 sg13g2_nand2_1 _28120_ (.Y(_09165_),
    .A(_08238_),
    .B(net499));
 sg13g2_nor2_1 _28121_ (.A(_09153_),
    .B(_09165_),
    .Y(_09166_));
 sg13g2_a221oi_1 _28122_ (.B2(net480),
    .C1(_09166_),
    .B1(_09164_),
    .A1(net134),
    .Y(_09167_),
    .A2(net68));
 sg13g2_nor2_1 _28123_ (.A(\stack[9][0] ),
    .B(net47),
    .Y(_09168_));
 sg13g2_a21oi_1 _28124_ (.A1(net47),
    .A2(_09167_),
    .Y(_02771_),
    .B1(_09168_));
 sg13g2_nand2_1 _28125_ (.Y(_09169_),
    .A(net1299),
    .B(net499));
 sg13g2_nor2_1 _28126_ (.A(_09153_),
    .B(_09169_),
    .Y(_09170_));
 sg13g2_a221oi_1 _28127_ (.B2(net402),
    .C1(_09170_),
    .B1(_09164_),
    .A1(_07701_),
    .Y(_09171_),
    .A2(net68));
 sg13g2_nor2_1 _28128_ (.A(\stack[9][1] ),
    .B(net47),
    .Y(_09172_));
 sg13g2_a21oi_1 _28129_ (.A1(net47),
    .A2(_09171_),
    .Y(_02772_),
    .B1(_09172_));
 sg13g2_nand2_1 _28130_ (.Y(_09173_),
    .A(_10015_),
    .B(net499));
 sg13g2_nor2_1 _28131_ (.A(_09153_),
    .B(_09173_),
    .Y(_09174_));
 sg13g2_a221oi_1 _28132_ (.B2(_07978_),
    .C1(_09174_),
    .B1(_09164_),
    .A1(_07739_),
    .Y(_09175_),
    .A2(net68));
 sg13g2_nor2_1 _28133_ (.A(\stack[9][2] ),
    .B(net47),
    .Y(_09176_));
 sg13g2_a21oi_1 _28134_ (.A1(net47),
    .A2(_09175_),
    .Y(_02773_),
    .B1(_09176_));
 sg13g2_nand2_1 _28135_ (.Y(_09177_),
    .A(net1300),
    .B(net499));
 sg13g2_nor2_1 _28136_ (.A(_09153_),
    .B(_09177_),
    .Y(_09178_));
 sg13g2_a221oi_1 _28137_ (.B2(net494),
    .C1(_09178_),
    .B1(_09164_),
    .A1(_07784_),
    .Y(_09179_),
    .A2(_09153_));
 sg13g2_nor2_1 _28138_ (.A(\stack[9][3] ),
    .B(_09161_),
    .Y(_09180_));
 sg13g2_a21oi_1 _28139_ (.A1(net47),
    .A2(_09179_),
    .Y(_02774_),
    .B1(_09180_));
 sg13g2_nand2_1 _28140_ (.Y(_09181_),
    .A(\stack[9][4] ),
    .B(_09159_));
 sg13g2_a221oi_1 _28141_ (.B2(net1222),
    .C1(net68),
    .B1(net499),
    .A1(net484),
    .Y(_09182_),
    .A2(_09164_));
 sg13g2_a22oi_1 _28142_ (.Y(_02775_),
    .B1(_09181_),
    .B2(_09182_),
    .A2(net68),
    .A1(net100));
 sg13g2_and2_1 _28143_ (.A(net1221),
    .B(net499),
    .X(_09183_));
 sg13g2_nor2_1 _28144_ (.A(net446),
    .B(_09154_),
    .Y(_09184_));
 sg13g2_and2_1 _28145_ (.A(\stack[9][5] ),
    .B(_09159_),
    .X(_09185_));
 sg13g2_nor4_1 _28146_ (.A(_09162_),
    .B(_09183_),
    .C(_09184_),
    .D(_09185_),
    .Y(_09186_));
 sg13g2_a21oi_1 _28147_ (.A1(_07990_),
    .A2(net68),
    .Y(_02776_),
    .B1(_09186_));
 sg13g2_a22oi_1 _28148_ (.Y(_09187_),
    .B1(net499),
    .B2(net1220),
    .A2(_09164_),
    .A1(net451));
 sg13g2_nand2_1 _28149_ (.Y(_09188_),
    .A(\stack[9][6] ),
    .B(_09159_));
 sg13g2_nand2_1 _28150_ (.Y(_09189_),
    .A(_09187_),
    .B(_09188_));
 sg13g2_mux2_1 _28151_ (.A0(_09189_),
    .A1(net42),
    .S(net68),
    .X(_02777_));
 sg13g2_a221oi_1 _28152_ (.B2(net1219),
    .C1(_09162_),
    .B1(_09156_),
    .A1(net294),
    .Y(_09190_),
    .A2(_09164_));
 sg13g2_nor2_1 _28153_ (.A(\stack[9][7] ),
    .B(_09161_),
    .Y(_09191_));
 sg13g2_a221oi_1 _28154_ (.B2(_09190_),
    .C1(_09191_),
    .B1(net47),
    .A1(net41),
    .Y(_02778_),
    .A2(net68));
 sg13g2_buf_1 _28155_ (.A(\exec.out_of_order_exec ),
    .X(_09192_));
 sg13g2_inv_1 _28156_ (.Y(_09193_),
    .A(_09192_));
 sg13g2_a21oi_1 _28157_ (.A1(_09193_),
    .A2(_09927_),
    .Y(_02499_),
    .B1(_09933_));
 sg13g2_buf_2 _28158_ (.A(net878),
    .X(_09194_));
 sg13g2_buf_1 _28159_ (.A(net792),
    .X(_09195_));
 sg13g2_buf_1 _28160_ (.A(net120),
    .X(_09196_));
 sg13g2_nor2_1 _28161_ (.A(_09944_),
    .B(_09964_),
    .Y(_09197_));
 sg13g2_nor2b_1 _28162_ (.A(net93),
    .B_N(_09197_),
    .Y(_09198_));
 sg13g2_a21oi_1 _28163_ (.A1(_09944_),
    .A2(net93),
    .Y(_09199_),
    .B1(_09198_));
 sg13g2_nor2_1 _28164_ (.A(_09195_),
    .B(_09199_),
    .Y(_00090_));
 sg13g2_buf_1 _28165_ (.A(_10066_),
    .X(_09200_));
 sg13g2_nor2_1 _28166_ (.A(_09942_),
    .B(_09947_),
    .Y(_09201_));
 sg13g2_and2_1 _28167_ (.A(_09950_),
    .B(_09201_),
    .X(_09202_));
 sg13g2_and2_1 _28168_ (.A(_09951_),
    .B(_09202_),
    .X(_09203_));
 sg13g2_and2_1 _28169_ (.A(_09952_),
    .B(_09203_),
    .X(_09204_));
 sg13g2_and2_1 _28170_ (.A(_09953_),
    .B(_09204_),
    .X(_09205_));
 sg13g2_nand3_1 _28171_ (.B(_09956_),
    .C(_09205_),
    .A(_09955_),
    .Y(_09206_));
 sg13g2_buf_1 _28172_ (.A(_09206_),
    .X(_09207_));
 sg13g2_a21o_1 _28173_ (.A2(_09207_),
    .A1(net448),
    .B1(net93),
    .X(_09208_));
 sg13g2_or2_1 _28174_ (.X(_09209_),
    .B(_10149_),
    .A(_09964_));
 sg13g2_buf_1 _28175_ (.A(_09209_),
    .X(_09210_));
 sg13g2_buf_1 _28176_ (.A(_09210_),
    .X(_09211_));
 sg13g2_nor3_1 _28177_ (.A(_09957_),
    .B(_09207_),
    .C(_09211_),
    .Y(_09212_));
 sg13g2_a21oi_1 _28178_ (.A1(_09957_),
    .A2(_09208_),
    .Y(_09213_),
    .B1(_09212_));
 sg13g2_nor2_1 _28179_ (.A(net570),
    .B(_09213_),
    .Y(_00091_));
 sg13g2_buf_1 _28180_ (.A(net1193),
    .X(_09214_));
 sg13g2_inv_1 _28181_ (.Y(_09215_),
    .A(_09957_));
 sg13g2_nor2_1 _28182_ (.A(_09215_),
    .B(_09207_),
    .Y(_09216_));
 sg13g2_nand2b_1 _28183_ (.Y(_09217_),
    .B(_09216_),
    .A_N(_09939_));
 sg13g2_nor2_1 _28184_ (.A(_09964_),
    .B(_09216_),
    .Y(_09218_));
 sg13g2_o21ai_1 _28185_ (.B1(_09939_),
    .Y(_09219_),
    .A1(_10157_),
    .A2(_09218_));
 sg13g2_o21ai_1 _28186_ (.B1(_09219_),
    .Y(_09220_),
    .A1(net67),
    .A2(_09217_));
 sg13g2_and2_1 _28187_ (.A(net791),
    .B(_09220_),
    .X(_00092_));
 sg13g2_nand2_1 _28188_ (.Y(_09221_),
    .A(_09939_),
    .B(_09216_));
 sg13g2_a21o_1 _28189_ (.A2(_09221_),
    .A1(_09200_),
    .B1(net93),
    .X(_09222_));
 sg13g2_nor3_1 _28190_ (.A(_09940_),
    .B(_09210_),
    .C(_09221_),
    .Y(_09223_));
 sg13g2_a21oi_1 _28191_ (.A1(_09940_),
    .A2(_09222_),
    .Y(_09224_),
    .B1(_09223_));
 sg13g2_nor2_1 _28192_ (.A(net570),
    .B(_09224_),
    .Y(_00093_));
 sg13g2_inv_1 _28193_ (.Y(_09225_),
    .A(_09940_));
 sg13g2_nor3_1 _28194_ (.A(_09225_),
    .B(net93),
    .C(_09221_),
    .Y(_09226_));
 sg13g2_nor2_1 _28195_ (.A(\delay_cycles[13] ),
    .B(_09226_),
    .Y(_09227_));
 sg13g2_o21ai_1 _28196_ (.B1(net791),
    .Y(_09228_),
    .A1(net448),
    .A2(net93));
 sg13g2_nor2_1 _28197_ (.A(_09227_),
    .B(_09228_),
    .Y(_00094_));
 sg13g2_and2_1 _28198_ (.A(net1192),
    .B(_10157_),
    .X(_09229_));
 sg13g2_buf_1 _28199_ (.A(_09229_),
    .X(_09230_));
 sg13g2_and2_1 _28200_ (.A(\delay_cycles[14] ),
    .B(net66),
    .X(_00095_));
 sg13g2_and2_1 _28201_ (.A(\delay_cycles[15] ),
    .B(net66),
    .X(_00096_));
 sg13g2_and2_1 _28202_ (.A(\delay_cycles[16] ),
    .B(net66),
    .X(_00097_));
 sg13g2_and2_1 _28203_ (.A(\delay_cycles[17] ),
    .B(net66),
    .X(_00098_));
 sg13g2_and2_1 _28204_ (.A(\delay_cycles[18] ),
    .B(net66),
    .X(_00099_));
 sg13g2_and2_1 _28205_ (.A(\delay_cycles[19] ),
    .B(net66),
    .X(_00100_));
 sg13g2_nand2b_1 _28206_ (.Y(_09231_),
    .B(_09944_),
    .A_N(_09943_));
 sg13g2_o21ai_1 _28207_ (.B1(_09943_),
    .Y(_09232_),
    .A1(net120),
    .A2(_09197_));
 sg13g2_o21ai_1 _28208_ (.B1(_09232_),
    .Y(_09233_),
    .A1(net67),
    .A2(_09231_));
 sg13g2_and2_1 _28209_ (.A(_09214_),
    .B(_09233_),
    .X(_00101_));
 sg13g2_and2_1 _28210_ (.A(\delay_cycles[20] ),
    .B(_09230_),
    .X(_00102_));
 sg13g2_and2_1 _28211_ (.A(\delay_cycles[21] ),
    .B(_09230_),
    .X(_00103_));
 sg13g2_and2_1 _28212_ (.A(\delay_cycles[22] ),
    .B(net66),
    .X(_00104_));
 sg13g2_and2_1 _28213_ (.A(\delay_cycles[23] ),
    .B(net66),
    .X(_00105_));
 sg13g2_nand2_1 _28214_ (.Y(_09234_),
    .A(_09943_),
    .B(_09944_));
 sg13g2_nor3_1 _28215_ (.A(_09945_),
    .B(_09234_),
    .C(net120),
    .Y(_09235_));
 sg13g2_a21o_1 _28216_ (.A2(_09234_),
    .A1(_09945_),
    .B1(_09235_),
    .X(_09236_));
 sg13g2_a22oi_1 _28217_ (.Y(_09237_),
    .B1(_09236_),
    .B2(net448),
    .A2(_09196_),
    .A1(_09945_));
 sg13g2_nor2_1 _28218_ (.A(net570),
    .B(_09237_),
    .Y(_00106_));
 sg13g2_a21o_1 _28219_ (.A2(_09200_),
    .A1(_09947_),
    .B1(_09196_),
    .X(_09238_));
 sg13g2_nor3_1 _28220_ (.A(\delay_cycles[3] ),
    .B(_09947_),
    .C(_09211_),
    .Y(_09239_));
 sg13g2_a21oi_1 _28221_ (.A1(\delay_cycles[3] ),
    .A2(_09238_),
    .Y(_09240_),
    .B1(_09239_));
 sg13g2_nor2_1 _28222_ (.A(_09195_),
    .B(_09240_),
    .Y(_00107_));
 sg13g2_a21o_1 _28223_ (.A2(_10066_),
    .A1(_09949_),
    .B1(net93),
    .X(_09241_));
 sg13g2_nor3_1 _28224_ (.A(_09950_),
    .B(_09949_),
    .C(net67),
    .Y(_09242_));
 sg13g2_a21oi_1 _28225_ (.A1(_09950_),
    .A2(_09241_),
    .Y(_09243_),
    .B1(_09242_));
 sg13g2_nor2_1 _28226_ (.A(net570),
    .B(_09243_),
    .Y(_00108_));
 sg13g2_nand2_1 _28227_ (.Y(_09244_),
    .A(_09950_),
    .B(_09201_));
 sg13g2_a21o_1 _28228_ (.A2(_09244_),
    .A1(net448),
    .B1(net93),
    .X(_09245_));
 sg13g2_nor3_1 _28229_ (.A(_09951_),
    .B(_09244_),
    .C(net67),
    .Y(_09246_));
 sg13g2_a21oi_1 _28230_ (.A1(_09951_),
    .A2(_09245_),
    .Y(_09247_),
    .B1(_09246_));
 sg13g2_nor2_1 _28231_ (.A(net570),
    .B(_09247_),
    .Y(_00109_));
 sg13g2_nand2_1 _28232_ (.Y(_09248_),
    .A(_09951_),
    .B(_09202_));
 sg13g2_a21o_1 _28233_ (.A2(_09248_),
    .A1(net448),
    .B1(net120),
    .X(_09249_));
 sg13g2_nor3_1 _28234_ (.A(_09952_),
    .B(_09248_),
    .C(net67),
    .Y(_09250_));
 sg13g2_a21oi_1 _28235_ (.A1(_09952_),
    .A2(_09249_),
    .Y(_09251_),
    .B1(_09250_));
 sg13g2_nor2_1 _28236_ (.A(net570),
    .B(_09251_),
    .Y(_00110_));
 sg13g2_nand2_1 _28237_ (.Y(_09252_),
    .A(_09952_),
    .B(_09203_));
 sg13g2_a21o_1 _28238_ (.A2(_09252_),
    .A1(net448),
    .B1(net120),
    .X(_09253_));
 sg13g2_nor3_1 _28239_ (.A(_09953_),
    .B(_09252_),
    .C(net67),
    .Y(_09254_));
 sg13g2_a21oi_1 _28240_ (.A1(_09953_),
    .A2(_09253_),
    .Y(_09255_),
    .B1(_09254_));
 sg13g2_nor2_1 _28241_ (.A(net570),
    .B(_09255_),
    .Y(_00111_));
 sg13g2_nand2_1 _28242_ (.Y(_09256_),
    .A(_09953_),
    .B(_09204_));
 sg13g2_a21o_1 _28243_ (.A2(_09256_),
    .A1(net448),
    .B1(net120),
    .X(_09257_));
 sg13g2_nor3_1 _28244_ (.A(_09955_),
    .B(_09256_),
    .C(net67),
    .Y(_09258_));
 sg13g2_a21oi_1 _28245_ (.A1(_09955_),
    .A2(_09257_),
    .Y(_09259_),
    .B1(_09258_));
 sg13g2_nor2_1 _28246_ (.A(net570),
    .B(_09259_),
    .Y(_00112_));
 sg13g2_buf_2 _28247_ (.A(net792),
    .X(_09260_));
 sg13g2_nand2_1 _28248_ (.Y(_09261_),
    .A(_09955_),
    .B(_09205_));
 sg13g2_a21o_1 _28249_ (.A2(_09261_),
    .A1(net448),
    .B1(net120),
    .X(_09262_));
 sg13g2_nor3_1 _28250_ (.A(_09956_),
    .B(_09261_),
    .C(net67),
    .Y(_09263_));
 sg13g2_a21oi_1 _28251_ (.A1(_09956_),
    .A2(_09262_),
    .Y(_09264_),
    .B1(_09263_));
 sg13g2_nor2_1 _28252_ (.A(_09260_),
    .B(_09264_),
    .Y(_00113_));
 sg13g2_o21ai_1 _28253_ (.B1(net791),
    .Y(_09265_),
    .A1(_00081_),
    .A2(_06123_));
 sg13g2_a21oi_1 _28254_ (.A1(_10237_),
    .A2(_10239_),
    .Y(_09266_),
    .B1(_10238_));
 sg13g2_nor2_1 _28255_ (.A(_09265_),
    .B(_09266_),
    .Y(_02162_));
 sg13g2_inv_1 _28256_ (.Y(_09267_),
    .A(_10238_));
 sg13g2_nand2_1 _28257_ (.Y(_09268_),
    .A(net791),
    .B(_10237_));
 sg13g2_a21oi_1 _28258_ (.A1(_09267_),
    .A2(_10239_),
    .Y(_02163_),
    .B1(_09268_));
 sg13g2_inv_1 _28259_ (.Y(_09269_),
    .A(_10237_));
 sg13g2_a21oi_1 _28260_ (.A1(_09269_),
    .A2(_09267_),
    .Y(_09270_),
    .B1(_09986_));
 sg13g2_nor2_1 _28261_ (.A(_10240_),
    .B(_09270_),
    .Y(_02428_));
 sg13g2_nor3_1 _28262_ (.A(_10236_),
    .B(net775),
    .C(_04224_),
    .Y(_09271_));
 sg13g2_buf_2 _28263_ (.A(_09271_),
    .X(_09272_));
 sg13g2_buf_2 _28264_ (.A(_10236_),
    .X(_09273_));
 sg13g2_nor3_1 _28265_ (.A(_09273_),
    .B(net554),
    .C(_04224_),
    .Y(_09274_));
 sg13g2_buf_2 _28266_ (.A(_09274_),
    .X(_09275_));
 sg13g2_nor3_1 _28267_ (.A(_10236_),
    .B(net778),
    .C(_04224_),
    .Y(_09276_));
 sg13g2_buf_2 _28268_ (.A(_09276_),
    .X(_09277_));
 sg13g2_and2_1 _28269_ (.A(net21),
    .B(_09277_),
    .X(_09278_));
 sg13g2_a221oi_1 _28270_ (.B2(net5),
    .C1(_09278_),
    .B1(_09275_),
    .A1(\mem.mem_io.porta_out[0] ),
    .Y(_09279_),
    .A2(_09272_));
 sg13g2_buf_1 _28271_ (.A(net558),
    .X(_09280_));
 sg13g2_a21oi_1 _28272_ (.A1(net1294),
    .A2(_10293_),
    .Y(_09281_),
    .B1(_10395_));
 sg13g2_o21ai_1 _28273_ (.B1(_00070_),
    .Y(_09282_),
    .A1(_04224_),
    .A2(_09281_));
 sg13g2_nand2_1 _28274_ (.Y(_09283_),
    .A(_09280_),
    .B(_09282_));
 sg13g2_buf_2 _28275_ (.A(_09283_),
    .X(_09284_));
 sg13g2_nor2_1 _28276_ (.A(_10372_),
    .B(_04224_),
    .Y(_09285_));
 sg13g2_buf_2 _28277_ (.A(_09285_),
    .X(_09286_));
 sg13g2_buf_1 _28278_ (.A(_09286_),
    .X(_09287_));
 sg13g2_nor2_1 _28279_ (.A(_10444_),
    .B(_04224_),
    .Y(_09288_));
 sg13g2_buf_2 _28280_ (.A(_09288_),
    .X(_09289_));
 sg13g2_buf_1 _28281_ (.A(_09289_),
    .X(_09290_));
 sg13g2_a22oi_1 _28282_ (.Y(_09291_),
    .B1(net512),
    .B2(\mem.mem_io.porta_oe[0] ),
    .A2(_09287_),
    .A1(net13));
 sg13g2_nor2_1 _28283_ (.A(net1207),
    .B(_09291_),
    .Y(_09292_));
 sg13g2_nor2_1 _28284_ (.A(_09284_),
    .B(_09292_),
    .Y(_09293_));
 sg13g2_o21ai_1 _28285_ (.B1(net791),
    .Y(_09294_),
    .A1(\mem.io_data_out[0] ),
    .A2(net519));
 sg13g2_a21oi_1 _28286_ (.A1(_09279_),
    .A2(_09293_),
    .Y(_02429_),
    .B1(_09294_));
 sg13g2_and2_1 _28287_ (.A(net22),
    .B(_09277_),
    .X(_09295_));
 sg13g2_a221oi_1 _28288_ (.B2(net6),
    .C1(_09295_),
    .B1(_09275_),
    .A1(\mem.mem_io.porta_out[1] ),
    .Y(_09296_),
    .A2(_09272_));
 sg13g2_a22oi_1 _28289_ (.Y(_09297_),
    .B1(net512),
    .B2(\mem.mem_io.porta_oe[1] ),
    .A2(_09287_),
    .A1(net14));
 sg13g2_nor2_1 _28290_ (.A(net1207),
    .B(_09297_),
    .Y(_09298_));
 sg13g2_nor2_1 _28291_ (.A(_09284_),
    .B(_09298_),
    .Y(_09299_));
 sg13g2_o21ai_1 _28292_ (.B1(net857),
    .Y(_09300_),
    .A1(\mem.io_data_out[1] ),
    .A2(net519));
 sg13g2_a21oi_1 _28293_ (.A1(_09296_),
    .A2(_09299_),
    .Y(_02430_),
    .B1(_09300_));
 sg13g2_and2_1 _28294_ (.A(net23),
    .B(_09277_),
    .X(_09301_));
 sg13g2_a221oi_1 _28295_ (.B2(net7),
    .C1(_09301_),
    .B1(_09275_),
    .A1(\mem.mem_io.porta_out[2] ),
    .Y(_09302_),
    .A2(_09272_));
 sg13g2_buf_1 _28296_ (.A(\mem.mem_io.porta_oe[2] ),
    .X(_09303_));
 sg13g2_a22oi_1 _28297_ (.Y(_09304_),
    .B1(_09289_),
    .B2(_09303_),
    .A2(_09286_),
    .A1(net15));
 sg13g2_nor2_1 _28298_ (.A(net1207),
    .B(_09304_),
    .Y(_09305_));
 sg13g2_nor2_1 _28299_ (.A(_09284_),
    .B(_09305_),
    .Y(_09306_));
 sg13g2_o21ai_1 _28300_ (.B1(net857),
    .Y(_09307_),
    .A1(\mem.io_data_out[2] ),
    .A2(net519));
 sg13g2_a21oi_1 _28301_ (.A1(_09302_),
    .A2(_09306_),
    .Y(_02431_),
    .B1(_09307_));
 sg13g2_and2_1 _28302_ (.A(net24),
    .B(_09277_),
    .X(_09308_));
 sg13g2_a221oi_1 _28303_ (.B2(net8),
    .C1(_09308_),
    .B1(_09275_),
    .A1(\mem.mem_io.porta_out[3] ),
    .Y(_09309_),
    .A2(_09272_));
 sg13g2_a22oi_1 _28304_ (.Y(_09310_),
    .B1(_09289_),
    .B2(\mem.mem_io.porta_oe[3] ),
    .A2(_09286_),
    .A1(net16));
 sg13g2_nor2_1 _28305_ (.A(net1207),
    .B(_09310_),
    .Y(_09311_));
 sg13g2_nor2_1 _28306_ (.A(_09284_),
    .B(_09311_),
    .Y(_09312_));
 sg13g2_o21ai_1 _28307_ (.B1(net857),
    .Y(_09313_),
    .A1(\mem.io_data_out[3] ),
    .A2(net519));
 sg13g2_a21oi_1 _28308_ (.A1(_09309_),
    .A2(_09312_),
    .Y(_02432_),
    .B1(_09313_));
 sg13g2_and2_1 _28309_ (.A(net25),
    .B(_09277_),
    .X(_09314_));
 sg13g2_a221oi_1 _28310_ (.B2(net9),
    .C1(_09314_),
    .B1(_09275_),
    .A1(\mem.mem_io.porta_out[4] ),
    .Y(_09315_),
    .A2(_09272_));
 sg13g2_a22oi_1 _28311_ (.Y(_09316_),
    .B1(_09289_),
    .B2(\mem.mem_io.porta_oe[4] ),
    .A2(_09286_),
    .A1(net17));
 sg13g2_nor2_1 _28312_ (.A(net1207),
    .B(_09316_),
    .Y(_09317_));
 sg13g2_nor2_1 _28313_ (.A(_09284_),
    .B(_09317_),
    .Y(_09318_));
 sg13g2_o21ai_1 _28314_ (.B1(net857),
    .Y(_09319_),
    .A1(\mem.io_data_out[4] ),
    .A2(net519));
 sg13g2_a21oi_1 _28315_ (.A1(_09315_),
    .A2(_09318_),
    .Y(_02433_),
    .B1(_09319_));
 sg13g2_and2_1 _28316_ (.A(net26),
    .B(_09277_),
    .X(_09320_));
 sg13g2_a221oi_1 _28317_ (.B2(net10),
    .C1(_09320_),
    .B1(_09275_),
    .A1(\mem.mem_io.porta_out[5] ),
    .Y(_09321_),
    .A2(_09272_));
 sg13g2_a22oi_1 _28318_ (.Y(_09322_),
    .B1(_09289_),
    .B2(\mem.mem_io.porta_oe[5] ),
    .A2(_09286_),
    .A1(net18));
 sg13g2_nor2_1 _28319_ (.A(net1207),
    .B(_09322_),
    .Y(_09323_));
 sg13g2_nor2_1 _28320_ (.A(_09284_),
    .B(_09323_),
    .Y(_09324_));
 sg13g2_o21ai_1 _28321_ (.B1(net857),
    .Y(_09325_),
    .A1(\mem.io_data_out[5] ),
    .A2(net519));
 sg13g2_a21oi_1 _28322_ (.A1(_09321_),
    .A2(_09324_),
    .Y(_02434_),
    .B1(_09325_));
 sg13g2_and2_1 _28323_ (.A(net27),
    .B(_09277_),
    .X(_09326_));
 sg13g2_a221oi_1 _28324_ (.B2(net11),
    .C1(_09326_),
    .B1(_09275_),
    .A1(\mem.mem_io.porta_out[6] ),
    .Y(_09327_),
    .A2(_09272_));
 sg13g2_a22oi_1 _28325_ (.Y(_09328_),
    .B1(_09289_),
    .B2(\mem.mem_io.porta_oe[6] ),
    .A2(_09286_),
    .A1(net19));
 sg13g2_nor2_1 _28326_ (.A(net1207),
    .B(_09328_),
    .Y(_09329_));
 sg13g2_nor2_1 _28327_ (.A(_09284_),
    .B(_09329_),
    .Y(_09330_));
 sg13g2_o21ai_1 _28328_ (.B1(net857),
    .Y(_09331_),
    .A1(\mem.io_data_out[6] ),
    .A2(net519));
 sg13g2_a21oi_1 _28329_ (.A1(_09327_),
    .A2(_09330_),
    .Y(_02435_),
    .B1(_09331_));
 sg13g2_and2_1 _28330_ (.A(net28),
    .B(_09277_),
    .X(_09332_));
 sg13g2_a221oi_1 _28331_ (.B2(net12),
    .C1(_09332_),
    .B1(_09275_),
    .A1(\mem.mem_io.porta_out[7] ),
    .Y(_09333_),
    .A2(_09272_));
 sg13g2_a22oi_1 _28332_ (.Y(_09334_),
    .B1(_09289_),
    .B2(\mem.mem_io.porta_oe[7] ),
    .A2(_09286_),
    .A1(net20));
 sg13g2_nor2_1 _28333_ (.A(net1207),
    .B(_09334_),
    .Y(_09335_));
 sg13g2_nor2_1 _28334_ (.A(_09284_),
    .B(_09335_),
    .Y(_09336_));
 sg13g2_o21ai_1 _28335_ (.B1(net857),
    .Y(_09337_),
    .A1(\mem.io_data_out[7] ),
    .A2(net519));
 sg13g2_a21oi_1 _28336_ (.A1(_09333_),
    .A2(_09336_),
    .Y(_02436_),
    .B1(_09337_));
 sg13g2_and2_1 _28337_ (.A(net791),
    .B(_09280_),
    .X(_02437_));
 sg13g2_and2_1 _28338_ (.A(_05430_),
    .B(net558),
    .X(_09338_));
 sg13g2_buf_1 _28339_ (.A(_09338_),
    .X(_09339_));
 sg13g2_buf_1 _28340_ (.A(net511),
    .X(_09340_));
 sg13g2_and2_1 _28341_ (.A(net791),
    .B(_09340_),
    .X(_02438_));
 sg13g2_nand3_1 _28342_ (.B(net512),
    .C(net498),
    .A(net1292),
    .Y(_09341_));
 sg13g2_nand2_1 _28343_ (.Y(_09342_),
    .A(_09289_),
    .B(_09339_));
 sg13g2_buf_2 _28344_ (.A(_09342_),
    .X(_09343_));
 sg13g2_nand2_1 _28345_ (.Y(_09344_),
    .A(\mem.mem_io.porta_oe[0] ),
    .B(_09343_));
 sg13g2_buf_2 _28346_ (.A(net878),
    .X(_09345_));
 sg13g2_a21oi_1 _28347_ (.A1(_09341_),
    .A2(_09344_),
    .Y(_02439_),
    .B1(net790));
 sg13g2_nand3_1 _28348_ (.B(_09290_),
    .C(_09340_),
    .A(_05445_),
    .Y(_09346_));
 sg13g2_nand2_1 _28349_ (.Y(_09347_),
    .A(\mem.mem_io.porta_oe[1] ),
    .B(_09343_));
 sg13g2_a21oi_1 _28350_ (.A1(_09346_),
    .A2(_09347_),
    .Y(_02440_),
    .B1(net790));
 sg13g2_nand3_1 _28351_ (.B(_09290_),
    .C(net498),
    .A(net1290),
    .Y(_09348_));
 sg13g2_nand2_1 _28352_ (.Y(_09349_),
    .A(_09303_),
    .B(_09343_));
 sg13g2_a21oi_1 _28353_ (.A1(_09348_),
    .A2(_09349_),
    .Y(_02441_),
    .B1(net790));
 sg13g2_nand3_1 _28354_ (.B(net512),
    .C(net498),
    .A(net1289),
    .Y(_09350_));
 sg13g2_nand2_1 _28355_ (.Y(_09351_),
    .A(\mem.mem_io.porta_oe[3] ),
    .B(_09343_));
 sg13g2_buf_1 _28356_ (.A(net878),
    .X(_09352_));
 sg13g2_a21oi_1 _28357_ (.A1(_09350_),
    .A2(_09351_),
    .Y(_02442_),
    .B1(net789));
 sg13g2_nand3_1 _28358_ (.B(net512),
    .C(net498),
    .A(net1288),
    .Y(_09353_));
 sg13g2_nand2_1 _28359_ (.Y(_09354_),
    .A(\mem.mem_io.porta_oe[4] ),
    .B(_09343_));
 sg13g2_a21oi_1 _28360_ (.A1(_09353_),
    .A2(_09354_),
    .Y(_02443_),
    .B1(net789));
 sg13g2_nand3_1 _28361_ (.B(net512),
    .C(net498),
    .A(net1287),
    .Y(_09355_));
 sg13g2_nand2_1 _28362_ (.Y(_09356_),
    .A(\mem.mem_io.porta_oe[5] ),
    .B(_09343_));
 sg13g2_a21oi_1 _28363_ (.A1(_09355_),
    .A2(_09356_),
    .Y(_02444_),
    .B1(_09352_));
 sg13g2_nand3_1 _28364_ (.B(net512),
    .C(net498),
    .A(net1286),
    .Y(_09357_));
 sg13g2_nand2_1 _28365_ (.Y(_09358_),
    .A(\mem.mem_io.porta_oe[6] ),
    .B(_09343_));
 sg13g2_a21oi_1 _28366_ (.A1(_09357_),
    .A2(_09358_),
    .Y(_02445_),
    .B1(_09352_));
 sg13g2_nand3_1 _28367_ (.B(net512),
    .C(net498),
    .A(net1285),
    .Y(_09359_));
 sg13g2_nand2_1 _28368_ (.Y(_09360_),
    .A(\mem.mem_io.porta_oe[7] ),
    .B(_09343_));
 sg13g2_a21oi_1 _28369_ (.A1(_09359_),
    .A2(_09360_),
    .Y(_02446_),
    .B1(net789));
 sg13g2_nand3_1 _28370_ (.B(net558),
    .C(_04225_),
    .A(_10236_),
    .Y(_09361_));
 sg13g2_buf_1 _28371_ (.A(_09361_),
    .X(_09362_));
 sg13g2_or2_1 _28372_ (.X(_09363_),
    .B(_09362_),
    .A(net775));
 sg13g2_buf_2 _28373_ (.A(_09363_),
    .X(_09364_));
 sg13g2_nand2_1 _28374_ (.Y(_09365_),
    .A(\mem.mem_io.porta_out[0] ),
    .B(_09364_));
 sg13g2_o21ai_1 _28375_ (.B1(net775),
    .Y(_09366_),
    .A1(\mem.mem_io.past_write ),
    .A2(_10422_));
 sg13g2_nor2b_1 _28376_ (.A(_09362_),
    .B_N(_09366_),
    .Y(_09367_));
 sg13g2_buf_2 _28377_ (.A(_09367_),
    .X(_09368_));
 sg13g2_nand2_1 _28378_ (.Y(_09369_),
    .A(_05441_),
    .B(_09368_));
 sg13g2_xnor2_1 _28379_ (.Y(_09370_),
    .A(_09365_),
    .B(_09369_));
 sg13g2_nor2_1 _28380_ (.A(_09260_),
    .B(_09370_),
    .Y(_02447_));
 sg13g2_nand2_1 _28381_ (.Y(_09371_),
    .A(\mem.mem_io.porta_out[1] ),
    .B(_09364_));
 sg13g2_nand2_1 _28382_ (.Y(_09372_),
    .A(net1291),
    .B(_09368_));
 sg13g2_xnor2_1 _28383_ (.Y(_09373_),
    .A(_09371_),
    .B(_09372_));
 sg13g2_nor2_1 _28384_ (.A(net569),
    .B(_09373_),
    .Y(_02448_));
 sg13g2_nand2_1 _28385_ (.Y(_09374_),
    .A(\mem.mem_io.porta_out[2] ),
    .B(_09364_));
 sg13g2_nand2_1 _28386_ (.Y(_09375_),
    .A(_05449_),
    .B(_09368_));
 sg13g2_xnor2_1 _28387_ (.Y(_09376_),
    .A(_09374_),
    .B(_09375_));
 sg13g2_nor2_1 _28388_ (.A(net569),
    .B(_09376_),
    .Y(_02449_));
 sg13g2_nand2_1 _28389_ (.Y(_09377_),
    .A(\mem.mem_io.porta_out[3] ),
    .B(_09364_));
 sg13g2_nand2_1 _28390_ (.Y(_09378_),
    .A(_05453_),
    .B(_09368_));
 sg13g2_xnor2_1 _28391_ (.Y(_09379_),
    .A(_09377_),
    .B(_09378_));
 sg13g2_nor2_1 _28392_ (.A(net569),
    .B(_09379_),
    .Y(_02450_));
 sg13g2_nand2_1 _28393_ (.Y(_09380_),
    .A(\mem.mem_io.porta_out[4] ),
    .B(_09364_));
 sg13g2_nand2_1 _28394_ (.Y(_09381_),
    .A(_05457_),
    .B(_09368_));
 sg13g2_xnor2_1 _28395_ (.Y(_09382_),
    .A(_09380_),
    .B(_09381_));
 sg13g2_nor2_1 _28396_ (.A(net569),
    .B(_09382_),
    .Y(_02451_));
 sg13g2_nand2_1 _28397_ (.Y(_09383_),
    .A(\mem.mem_io.porta_out[5] ),
    .B(_09364_));
 sg13g2_nand2_1 _28398_ (.Y(_09384_),
    .A(_05463_),
    .B(_09368_));
 sg13g2_xnor2_1 _28399_ (.Y(_09385_),
    .A(_09383_),
    .B(_09384_));
 sg13g2_nor2_1 _28400_ (.A(net569),
    .B(_09385_),
    .Y(_02452_));
 sg13g2_nand2_1 _28401_ (.Y(_09386_),
    .A(\mem.mem_io.porta_out[6] ),
    .B(_09364_));
 sg13g2_nand2_1 _28402_ (.Y(_09387_),
    .A(_05467_),
    .B(_09368_));
 sg13g2_xnor2_1 _28403_ (.Y(_09388_),
    .A(_09386_),
    .B(_09387_));
 sg13g2_nor2_1 _28404_ (.A(net569),
    .B(_09388_),
    .Y(_02453_));
 sg13g2_nand2_1 _28405_ (.Y(_09389_),
    .A(\mem.mem_io.porta_out[7] ),
    .B(_09364_));
 sg13g2_nand2_1 _28406_ (.Y(_09390_),
    .A(net1285),
    .B(_09368_));
 sg13g2_xnor2_1 _28407_ (.Y(_09391_),
    .A(_09389_),
    .B(_09390_));
 sg13g2_nor2_1 _28408_ (.A(net569),
    .B(_09391_),
    .Y(_02454_));
 sg13g2_nand3_1 _28409_ (.B(net513),
    .C(net498),
    .A(net1292),
    .Y(_09392_));
 sg13g2_nand2_1 _28410_ (.Y(_09393_),
    .A(_09286_),
    .B(_09339_));
 sg13g2_buf_2 _28411_ (.A(_09393_),
    .X(_09394_));
 sg13g2_nand2_1 _28412_ (.Y(_09395_),
    .A(net13),
    .B(_09394_));
 sg13g2_a21oi_1 _28413_ (.A1(_09392_),
    .A2(_09395_),
    .Y(_02455_),
    .B1(net789));
 sg13g2_nand3_1 _28414_ (.B(net513),
    .C(net511),
    .A(net1291),
    .Y(_09396_));
 sg13g2_nand2_1 _28415_ (.Y(_09397_),
    .A(net14),
    .B(_09394_));
 sg13g2_a21oi_1 _28416_ (.A1(_09396_),
    .A2(_09397_),
    .Y(_02456_),
    .B1(net789));
 sg13g2_nand3_1 _28417_ (.B(net513),
    .C(net511),
    .A(net1290),
    .Y(_09398_));
 sg13g2_nand2_1 _28418_ (.Y(_09399_),
    .A(net15),
    .B(_09394_));
 sg13g2_a21oi_1 _28419_ (.A1(_09398_),
    .A2(_09399_),
    .Y(_02457_),
    .B1(net789));
 sg13g2_nand3_1 _28420_ (.B(net513),
    .C(net511),
    .A(net1289),
    .Y(_09400_));
 sg13g2_nand2_1 _28421_ (.Y(_09401_),
    .A(net16),
    .B(_09394_));
 sg13g2_a21oi_1 _28422_ (.A1(_09400_),
    .A2(_09401_),
    .Y(_02458_),
    .B1(net789));
 sg13g2_nand3_1 _28423_ (.B(net513),
    .C(net511),
    .A(net1288),
    .Y(_09402_));
 sg13g2_nand2_1 _28424_ (.Y(_09403_),
    .A(net17),
    .B(_09394_));
 sg13g2_a21oi_1 _28425_ (.A1(_09402_),
    .A2(_09403_),
    .Y(_02459_),
    .B1(net789));
 sg13g2_nand3_1 _28426_ (.B(net513),
    .C(net511),
    .A(net1287),
    .Y(_09404_));
 sg13g2_nand2_1 _28427_ (.Y(_09405_),
    .A(net18),
    .B(_09394_));
 sg13g2_a21oi_1 _28428_ (.A1(_09404_),
    .A2(_09405_),
    .Y(_02460_),
    .B1(net792));
 sg13g2_nand3_1 _28429_ (.B(net513),
    .C(net511),
    .A(net1286),
    .Y(_09406_));
 sg13g2_nand2_1 _28430_ (.Y(_09407_),
    .A(net19),
    .B(_09394_));
 sg13g2_a21oi_1 _28431_ (.A1(_09406_),
    .A2(_09407_),
    .Y(_02461_),
    .B1(net792));
 sg13g2_nand3_1 _28432_ (.B(net513),
    .C(net511),
    .A(net1285),
    .Y(_09408_));
 sg13g2_nand2_1 _28433_ (.Y(_09409_),
    .A(net20),
    .B(_09394_));
 sg13g2_a21oi_1 _28434_ (.A1(_09408_),
    .A2(_09409_),
    .Y(_02462_),
    .B1(net792));
 sg13g2_o21ai_1 _28435_ (.B1(net778),
    .Y(_09410_),
    .A1(\mem.mem_io.past_write ),
    .A2(net779));
 sg13g2_nor2b_1 _28436_ (.A(_09362_),
    .B_N(_09410_),
    .Y(_09411_));
 sg13g2_buf_2 _28437_ (.A(_09411_),
    .X(_09412_));
 sg13g2_nand2_1 _28438_ (.Y(_09413_),
    .A(net1292),
    .B(_09412_));
 sg13g2_or2_1 _28439_ (.X(_09414_),
    .B(_09362_),
    .A(net778));
 sg13g2_buf_2 _28440_ (.A(_09414_),
    .X(_09415_));
 sg13g2_nand2_1 _28441_ (.Y(_09416_),
    .A(net21),
    .B(_09415_));
 sg13g2_xnor2_1 _28442_ (.Y(_09417_),
    .A(_09413_),
    .B(_09416_));
 sg13g2_nor2_1 _28443_ (.A(net569),
    .B(_09417_),
    .Y(_02463_));
 sg13g2_buf_2 _28444_ (.A(net792),
    .X(_09418_));
 sg13g2_nand2_1 _28445_ (.Y(_09419_),
    .A(net1291),
    .B(_09412_));
 sg13g2_nand2_1 _28446_ (.Y(_09420_),
    .A(net22),
    .B(_09415_));
 sg13g2_xnor2_1 _28447_ (.Y(_09421_),
    .A(_09419_),
    .B(_09420_));
 sg13g2_nor2_1 _28448_ (.A(net568),
    .B(_09421_),
    .Y(_02464_));
 sg13g2_nand2_1 _28449_ (.Y(_09422_),
    .A(net1290),
    .B(_09412_));
 sg13g2_nand2_1 _28450_ (.Y(_09423_),
    .A(net23),
    .B(_09415_));
 sg13g2_xnor2_1 _28451_ (.Y(_09424_),
    .A(_09422_),
    .B(_09423_));
 sg13g2_nor2_1 _28452_ (.A(net568),
    .B(_09424_),
    .Y(_02465_));
 sg13g2_nand2_1 _28453_ (.Y(_09425_),
    .A(net1289),
    .B(_09412_));
 sg13g2_nand2_1 _28454_ (.Y(_09426_),
    .A(net24),
    .B(_09415_));
 sg13g2_xnor2_1 _28455_ (.Y(_09427_),
    .A(_09425_),
    .B(_09426_));
 sg13g2_nor2_1 _28456_ (.A(net568),
    .B(_09427_),
    .Y(_02466_));
 sg13g2_nand2_1 _28457_ (.Y(_09428_),
    .A(net1288),
    .B(_09412_));
 sg13g2_nand2_1 _28458_ (.Y(_09429_),
    .A(net25),
    .B(_09415_));
 sg13g2_xnor2_1 _28459_ (.Y(_09430_),
    .A(_09428_),
    .B(_09429_));
 sg13g2_nor2_1 _28460_ (.A(net568),
    .B(_09430_),
    .Y(_02467_));
 sg13g2_nand2_1 _28461_ (.Y(_09431_),
    .A(net1287),
    .B(_09412_));
 sg13g2_nand2_1 _28462_ (.Y(_09432_),
    .A(net26),
    .B(_09415_));
 sg13g2_xnor2_1 _28463_ (.Y(_09433_),
    .A(_09431_),
    .B(_09432_));
 sg13g2_nor2_1 _28464_ (.A(net568),
    .B(_09433_),
    .Y(_02468_));
 sg13g2_nand2_1 _28465_ (.Y(_09434_),
    .A(net1286),
    .B(_09412_));
 sg13g2_nand2_1 _28466_ (.Y(_09435_),
    .A(net27),
    .B(_09415_));
 sg13g2_xnor2_1 _28467_ (.Y(_09436_),
    .A(_09434_),
    .B(_09435_));
 sg13g2_nor2_1 _28468_ (.A(net568),
    .B(_09436_),
    .Y(_02469_));
 sg13g2_nand2_1 _28469_ (.Y(_09437_),
    .A(_05471_),
    .B(_09412_));
 sg13g2_nand2_1 _28470_ (.Y(_09438_),
    .A(net28),
    .B(_09415_));
 sg13g2_xnor2_1 _28471_ (.Y(_09439_),
    .A(_09437_),
    .B(_09438_));
 sg13g2_nor2_1 _28472_ (.A(net568),
    .B(_09439_),
    .Y(_02470_));
 sg13g2_nor3_1 _28473_ (.A(_09991_),
    .B(_09987_),
    .C(_10008_),
    .Y(_09440_));
 sg13g2_a21oi_1 _28474_ (.A1(_09991_),
    .A2(_10008_),
    .Y(_09441_),
    .B1(_09987_));
 sg13g2_nor2_1 _28475_ (.A(_10004_),
    .B(_09441_),
    .Y(_09442_));
 sg13g2_nor3_1 _28476_ (.A(net792),
    .B(_09440_),
    .C(_09442_),
    .Y(_02471_));
 sg13g2_nor2_1 _28477_ (.A(_09987_),
    .B(_10008_),
    .Y(_09443_));
 sg13g2_a22oi_1 _28478_ (.Y(_09444_),
    .B1(_09443_),
    .B2(_09273_),
    .A2(_10004_),
    .A1(_09987_));
 sg13g2_nor2_1 _28479_ (.A(net568),
    .B(_09444_),
    .Y(_02473_));
 sg13g2_nor2_2 _28480_ (.A(_09418_),
    .B(_10025_),
    .Y(_02490_));
 sg13g2_nand2_1 _28481_ (.Y(_09445_),
    .A(net1208),
    .B(net858));
 sg13g2_nand2_1 _28482_ (.Y(_09446_),
    .A(net1275),
    .B(net1194));
 sg13g2_a21oi_1 _28483_ (.A1(_09445_),
    .A2(_09446_),
    .Y(_09447_),
    .B1(net557));
 sg13g2_a21oi_1 _28484_ (.A1(_10047_),
    .A2(net557),
    .Y(_09448_),
    .B1(_09447_));
 sg13g2_nor2_1 _28485_ (.A(_09418_),
    .B(_09448_),
    .Y(_02491_));
 sg13g2_buf_1 _28486_ (.A(net792),
    .X(_09449_));
 sg13g2_nand2_1 _28487_ (.Y(_09450_),
    .A(net1299),
    .B(net858));
 sg13g2_nand2_1 _28488_ (.Y(_09451_),
    .A(net1278),
    .B(net1194));
 sg13g2_a21oi_1 _28489_ (.A1(_09450_),
    .A2(_09451_),
    .Y(_09452_),
    .B1(net782));
 sg13g2_a21oi_1 _28490_ (.A1(_10041_),
    .A2(net557),
    .Y(_09453_),
    .B1(_09452_));
 sg13g2_nor2_1 _28491_ (.A(net567),
    .B(_09453_),
    .Y(_02492_));
 sg13g2_nand2_1 _28492_ (.Y(_09454_),
    .A(net1301),
    .B(net858));
 sg13g2_nand2_1 _28493_ (.Y(_09455_),
    .A(net1227),
    .B(net1194));
 sg13g2_a21oi_1 _28494_ (.A1(_09454_),
    .A2(_09455_),
    .Y(_09456_),
    .B1(net782));
 sg13g2_a21oi_1 _28495_ (.A1(_10052_),
    .A2(net557),
    .Y(_09457_),
    .B1(_09456_));
 sg13g2_nor2_1 _28496_ (.A(net567),
    .B(_09457_),
    .Y(_02493_));
 sg13g2_nand2_1 _28497_ (.Y(_09458_),
    .A(net1223),
    .B(net858));
 sg13g2_nand2_1 _28498_ (.Y(_09459_),
    .A(net1277),
    .B(net1194));
 sg13g2_a21oi_1 _28499_ (.A1(_09458_),
    .A2(_09459_),
    .Y(_09460_),
    .B1(net782));
 sg13g2_a21oi_1 _28500_ (.A1(_10049_),
    .A2(net557),
    .Y(_09461_),
    .B1(_09460_));
 sg13g2_nor2_1 _28501_ (.A(net567),
    .B(_09461_),
    .Y(_02494_));
 sg13g2_nand2_1 _28502_ (.Y(_09462_),
    .A(net1209),
    .B(net858));
 sg13g2_nand2_1 _28503_ (.Y(_09463_),
    .A(net1305),
    .B(net1194));
 sg13g2_a21oi_1 _28504_ (.A1(_09462_),
    .A2(_09463_),
    .Y(_09464_),
    .B1(net782));
 sg13g2_a21oi_1 _28505_ (.A1(_10040_),
    .A2(_10072_),
    .Y(_09465_),
    .B1(_09464_));
 sg13g2_nor2_1 _28506_ (.A(net567),
    .B(_09465_),
    .Y(_02495_));
 sg13g2_nand2_1 _28507_ (.Y(_09466_),
    .A(net1221),
    .B(net858));
 sg13g2_nand2_1 _28508_ (.Y(_09467_),
    .A(net1308),
    .B(net1194));
 sg13g2_a21oi_1 _28509_ (.A1(_09466_),
    .A2(_09467_),
    .Y(_09468_),
    .B1(net782));
 sg13g2_a21oi_1 _28510_ (.A1(_10044_),
    .A2(net557),
    .Y(_09469_),
    .B1(_09468_));
 sg13g2_nor2_1 _28511_ (.A(net567),
    .B(_09469_),
    .Y(_02496_));
 sg13g2_nand2_1 _28512_ (.Y(_09470_),
    .A(_07853_),
    .B(net858));
 sg13g2_nand2_1 _28513_ (.Y(_09471_),
    .A(net1307),
    .B(net1194));
 sg13g2_a21oi_1 _28514_ (.A1(_09470_),
    .A2(_09471_),
    .Y(_09472_),
    .B1(net782));
 sg13g2_a21oi_1 _28515_ (.A1(_10054_),
    .A2(net557),
    .Y(_09473_),
    .B1(_09472_));
 sg13g2_nor2_1 _28516_ (.A(net567),
    .B(_09473_),
    .Y(_02497_));
 sg13g2_nand2_1 _28517_ (.Y(_09474_),
    .A(net1213),
    .B(_10064_));
 sg13g2_nand2_1 _28518_ (.Y(_09475_),
    .A(net1309),
    .B(_09926_));
 sg13g2_a21oi_1 _28519_ (.A1(_09474_),
    .A2(_09475_),
    .Y(_09476_),
    .B1(net782));
 sg13g2_a21oi_1 _28520_ (.A1(_10042_),
    .A2(net557),
    .Y(_09477_),
    .B1(_09476_));
 sg13g2_nor2_1 _28521_ (.A(net567),
    .B(_09477_),
    .Y(_02498_));
 sg13g2_and2_1 _28522_ (.A(net791),
    .B(net1),
    .X(_02500_));
 sg13g2_buf_1 _28523_ (.A(net1272),
    .X(_09478_));
 sg13g2_inv_1 _28524_ (.Y(_09479_),
    .A(_09922_));
 sg13g2_buf_4 _28525_ (.X(_09480_),
    .A(_09479_));
 sg13g2_and2_1 _28526_ (.A(_09480_),
    .B(_09925_),
    .X(_09481_));
 sg13g2_buf_4 _28527_ (.X(_09482_),
    .A(_09481_));
 sg13g2_mux2_1 _28528_ (.A0(_10086_),
    .A1(net1218),
    .S(_09482_),
    .X(_09483_));
 sg13g2_buf_1 _28529_ (.A(net1272),
    .X(_09484_));
 sg13g2_o21ai_1 _28530_ (.B1(_07564_),
    .Y(_09485_),
    .A1(net524),
    .A2(_07579_));
 sg13g2_buf_2 _28531_ (.A(_09485_),
    .X(_09486_));
 sg13g2_buf_1 _28532_ (.A(_09486_),
    .X(_09487_));
 sg13g2_xor2_1 _28533_ (.B(_09192_),
    .A(_10086_),
    .X(_09488_));
 sg13g2_nor2_1 _28534_ (.A(_09487_),
    .B(_09488_),
    .Y(_09489_));
 sg13g2_a21oi_1 _28535_ (.A1(net495),
    .A2(_09487_),
    .Y(_09490_),
    .B1(_09489_));
 sg13g2_nand2_1 _28536_ (.Y(_09491_),
    .A(net876),
    .B(_09490_));
 sg13g2_o21ai_1 _28537_ (.B1(_09491_),
    .Y(_09492_),
    .A1(net877),
    .A2(_09483_));
 sg13g2_nor2_1 _28538_ (.A(_09449_),
    .B(_09492_),
    .Y(_02501_));
 sg13g2_mux2_1 _28539_ (.A0(_10099_),
    .A1(net1225),
    .S(_09482_),
    .X(_09493_));
 sg13g2_xor2_1 _28540_ (.B(_10099_),
    .A(_10086_),
    .X(_09494_));
 sg13g2_nand2_1 _28541_ (.Y(_09495_),
    .A(_09192_),
    .B(_00073_));
 sg13g2_o21ai_1 _28542_ (.B1(_09495_),
    .Y(_09496_),
    .A1(_09192_),
    .A2(_09494_));
 sg13g2_nor2_1 _28543_ (.A(net132),
    .B(_09496_),
    .Y(_09497_));
 sg13g2_a21oi_1 _28544_ (.A1(_10097_),
    .A2(net132),
    .Y(_09498_),
    .B1(_09497_));
 sg13g2_nand2_1 _28545_ (.Y(_09499_),
    .A(net876),
    .B(_09498_));
 sg13g2_o21ai_1 _28546_ (.B1(_09499_),
    .Y(_09500_),
    .A1(net877),
    .A2(_09493_));
 sg13g2_nor2_1 _28547_ (.A(_09449_),
    .B(_09500_),
    .Y(_02502_));
 sg13g2_mux2_1 _28548_ (.A0(_10104_),
    .A1(net1224),
    .S(_09482_),
    .X(_09501_));
 sg13g2_and3_1 _28549_ (.X(_09502_),
    .A(_10086_),
    .B(_10099_),
    .C(_09193_));
 sg13g2_buf_1 _28550_ (.A(_09502_),
    .X(_09503_));
 sg13g2_xor2_1 _28551_ (.B(_09503_),
    .A(_00074_),
    .X(_09504_));
 sg13g2_nor2_1 _28552_ (.A(_09486_),
    .B(_09504_),
    .Y(_09505_));
 sg13g2_a21oi_1 _28553_ (.A1(net485),
    .A2(net132),
    .Y(_09506_),
    .B1(_09505_));
 sg13g2_nand2_1 _28554_ (.Y(_09507_),
    .A(net876),
    .B(_09506_));
 sg13g2_o21ai_1 _28555_ (.B1(_09507_),
    .Y(_09508_),
    .A1(net877),
    .A2(_09501_));
 sg13g2_nor2_1 _28556_ (.A(net567),
    .B(_09508_),
    .Y(_02503_));
 sg13g2_buf_1 _28557_ (.A(_09194_),
    .X(_09509_));
 sg13g2_mux2_1 _28558_ (.A0(_10108_),
    .A1(net1223),
    .S(_09482_),
    .X(_09510_));
 sg13g2_nand2_1 _28559_ (.Y(_09511_),
    .A(_10104_),
    .B(_09503_));
 sg13g2_xnor2_1 _28560_ (.Y(_09512_),
    .A(_00075_),
    .B(_09511_));
 sg13g2_nor2_1 _28561_ (.A(_09486_),
    .B(_09512_),
    .Y(_09513_));
 sg13g2_a21oi_1 _28562_ (.A1(_10177_),
    .A2(net132),
    .Y(_09514_),
    .B1(_09513_));
 sg13g2_nand2_1 _28563_ (.Y(_09515_),
    .A(net876),
    .B(_09514_));
 sg13g2_o21ai_1 _28564_ (.B1(_09515_),
    .Y(_09516_),
    .A1(net877),
    .A2(_09510_));
 sg13g2_nor2_1 _28565_ (.A(net566),
    .B(_09516_),
    .Y(_02504_));
 sg13g2_mux2_1 _28566_ (.A0(_10119_),
    .A1(net1210),
    .S(_09482_),
    .X(_09517_));
 sg13g2_and3_1 _28567_ (.X(_09518_),
    .A(_10104_),
    .B(_10108_),
    .C(_09503_));
 sg13g2_buf_1 _28568_ (.A(_09518_),
    .X(_09519_));
 sg13g2_xor2_1 _28569_ (.B(_09519_),
    .A(_00076_),
    .X(_09520_));
 sg13g2_nor2_1 _28570_ (.A(_09486_),
    .B(_09520_),
    .Y(_09521_));
 sg13g2_a21oi_1 _28571_ (.A1(net493),
    .A2(net132),
    .Y(_09522_),
    .B1(_09521_));
 sg13g2_nand2_1 _28572_ (.Y(_09523_),
    .A(net876),
    .B(_09522_));
 sg13g2_o21ai_1 _28573_ (.B1(_09523_),
    .Y(_09524_),
    .A1(net877),
    .A2(_09517_));
 sg13g2_nor2_1 _28574_ (.A(net566),
    .B(_09524_),
    .Y(_02505_));
 sg13g2_mux2_1 _28575_ (.A0(_10129_),
    .A1(net1214),
    .S(_09482_),
    .X(_09525_));
 sg13g2_nand2_1 _28576_ (.Y(_09526_),
    .A(_10119_),
    .B(_09519_));
 sg13g2_xnor2_1 _28577_ (.Y(_09527_),
    .A(_00077_),
    .B(_09526_));
 sg13g2_nor2_1 _28578_ (.A(_09486_),
    .B(_09527_),
    .Y(_09528_));
 sg13g2_a21oi_1 _28579_ (.A1(_10199_),
    .A2(net132),
    .Y(_09529_),
    .B1(_09528_));
 sg13g2_nand2_1 _28580_ (.Y(_09530_),
    .A(_09484_),
    .B(_09529_));
 sg13g2_o21ai_1 _28581_ (.B1(_09530_),
    .Y(_09531_),
    .A1(net877),
    .A2(_09525_));
 sg13g2_nor2_1 _28582_ (.A(_09509_),
    .B(_09531_),
    .Y(_02506_));
 sg13g2_mux2_1 _28583_ (.A0(_10133_),
    .A1(_07853_),
    .S(_09482_),
    .X(_09532_));
 sg13g2_nand3_1 _28584_ (.B(_10129_),
    .C(_09519_),
    .A(_10119_),
    .Y(_09533_));
 sg13g2_xnor2_1 _28585_ (.Y(_09534_),
    .A(_00078_),
    .B(_09533_));
 sg13g2_nor2_1 _28586_ (.A(_09486_),
    .B(_09534_),
    .Y(_09535_));
 sg13g2_a21oi_1 _28587_ (.A1(_10211_),
    .A2(net132),
    .Y(_09536_),
    .B1(_09535_));
 sg13g2_nand2_1 _28588_ (.Y(_09537_),
    .A(net876),
    .B(_09536_));
 sg13g2_o21ai_1 _28589_ (.B1(_09537_),
    .Y(_09538_),
    .A1(net876),
    .A2(_09532_));
 sg13g2_nor2_1 _28590_ (.A(net566),
    .B(_09538_),
    .Y(_02507_));
 sg13g2_mux2_1 _28591_ (.A0(\exec.pc[7] ),
    .A1(net1219),
    .S(_09482_),
    .X(_09539_));
 sg13g2_nand4_1 _28592_ (.B(_10129_),
    .C(_10133_),
    .A(_10119_),
    .Y(_09540_),
    .D(_09519_));
 sg13g2_xnor2_1 _28593_ (.Y(_09541_),
    .A(_00079_),
    .B(_09540_));
 sg13g2_nor2_1 _28594_ (.A(_09486_),
    .B(_09541_),
    .Y(_09542_));
 sg13g2_a21oi_1 _28595_ (.A1(_10222_),
    .A2(net132),
    .Y(_09543_),
    .B1(_09542_));
 sg13g2_nand2_1 _28596_ (.Y(_09544_),
    .A(net1272),
    .B(_09543_));
 sg13g2_o21ai_1 _28597_ (.B1(_09544_),
    .Y(_09545_),
    .A1(net876),
    .A2(_09539_));
 sg13g2_nor2_1 _28598_ (.A(net566),
    .B(_09545_),
    .Y(_02508_));
 sg13g2_buf_2 _28599_ (.A(ui_in[3]),
    .X(_09546_));
 sg13g2_buf_1 _28600_ (.A(_09546_),
    .X(_09547_));
 sg13g2_buf_1 _28601_ (.A(_09924_),
    .X(_09548_));
 sg13g2_mux4_1 _28602_ (.S0(_09480_),
    .A0(_09914_),
    .A1(_10086_),
    .A2(_10165_),
    .A3(_07577_),
    .S1(net1283),
    .X(_09549_));
 sg13g2_nor2b_1 _28603_ (.A(net1284),
    .B_N(net4),
    .Y(_09550_));
 sg13g2_a21oi_1 _28604_ (.A1(net1284),
    .A2(_09549_),
    .Y(_09551_),
    .B1(_09550_));
 sg13g2_nor2_1 _28605_ (.A(net566),
    .B(_09551_),
    .Y(_02509_));
 sg13g2_inv_1 _28606_ (.Y(_09552_),
    .A(_00066_));
 sg13g2_mux4_1 _28607_ (.S0(_09480_),
    .A0(net1278),
    .A1(_10099_),
    .A2(_10097_),
    .A3(_09552_),
    .S1(net1283),
    .X(_09553_));
 sg13g2_nor2b_1 _28608_ (.A(_09546_),
    .B_N(net1218),
    .Y(_09554_));
 sg13g2_a21oi_1 _28609_ (.A1(net1284),
    .A2(_09553_),
    .Y(_09555_),
    .B1(_09554_));
 sg13g2_nor2_1 _28610_ (.A(net566),
    .B(_09555_),
    .Y(_02510_));
 sg13g2_inv_1 _28611_ (.Y(_09556_),
    .A(_07532_));
 sg13g2_mux4_1 _28612_ (.S0(_09480_),
    .A0(_07101_),
    .A1(_10104_),
    .A2(net485),
    .A3(_09556_),
    .S1(net1283),
    .X(_09557_));
 sg13g2_nor2b_1 _28613_ (.A(_09546_),
    .B_N(net1212),
    .Y(_09558_));
 sg13g2_a21oi_1 _28614_ (.A1(net1284),
    .A2(_09557_),
    .Y(_09559_),
    .B1(_09558_));
 sg13g2_nor2_1 _28615_ (.A(net566),
    .B(_09559_),
    .Y(_02511_));
 sg13g2_mux4_1 _28616_ (.S0(_09480_),
    .A0(_09889_),
    .A1(_10108_),
    .A2(net510),
    .A3(_09633_),
    .S1(net1283),
    .X(_09560_));
 sg13g2_nor2b_1 _28617_ (.A(_09546_),
    .B_N(net1217),
    .Y(_09561_));
 sg13g2_a21oi_1 _28618_ (.A1(net1284),
    .A2(_09560_),
    .Y(_09562_),
    .B1(_09561_));
 sg13g2_nor2_1 _28619_ (.A(net566),
    .B(_09562_),
    .Y(_02512_));
 sg13g2_mux4_1 _28620_ (.S0(_09480_),
    .A0(net1305),
    .A1(_10119_),
    .A2(net493),
    .A3(_09653_),
    .S1(net1283),
    .X(_09563_));
 sg13g2_nor2b_1 _28621_ (.A(_09546_),
    .B_N(net1211),
    .Y(_09564_));
 sg13g2_a21oi_1 _28622_ (.A1(net1284),
    .A2(_09563_),
    .Y(_09565_),
    .B1(_09564_));
 sg13g2_nor2_1 _28623_ (.A(_09509_),
    .B(_09565_),
    .Y(_02513_));
 sg13g2_nand2_1 _28624_ (.Y(_09566_),
    .A(_09548_),
    .B(_09922_));
 sg13g2_buf_2 _28625_ (.A(_09566_),
    .X(_09567_));
 sg13g2_mux2_1 _28626_ (.A0(_10129_),
    .A1(net1308),
    .S(_09923_),
    .X(_09568_));
 sg13g2_nand2b_1 _28627_ (.Y(_09569_),
    .B(_09568_),
    .A_N(net1283));
 sg13g2_o21ai_1 _28628_ (.B1(_09569_),
    .Y(_09570_),
    .A1(net446),
    .A2(_09567_));
 sg13g2_nor2_1 _28629_ (.A(_08252_),
    .B(_09547_),
    .Y(_09571_));
 sg13g2_a21oi_1 _28630_ (.A1(net1284),
    .A2(_09570_),
    .Y(_09572_),
    .B1(_09571_));
 sg13g2_nor2_1 _28631_ (.A(net790),
    .B(_09572_),
    .Y(_02514_));
 sg13g2_mux2_1 _28632_ (.A0(_10133_),
    .A1(net1307),
    .S(net1303),
    .X(_09573_));
 sg13g2_nand2b_1 _28633_ (.Y(_09574_),
    .B(_09573_),
    .A_N(net1283));
 sg13g2_nand2b_1 _28634_ (.Y(_09575_),
    .B(_10211_),
    .A_N(_09567_));
 sg13g2_nand3_1 _28635_ (.B(_09574_),
    .C(_09575_),
    .A(_09546_),
    .Y(_09576_));
 sg13g2_o21ai_1 _28636_ (.B1(_09576_),
    .Y(_09577_),
    .A1(net1216),
    .A2(net1284));
 sg13g2_nor2_1 _28637_ (.A(net790),
    .B(_09577_),
    .Y(_02515_));
 sg13g2_mux2_1 _28638_ (.A0(\exec.pc[7] ),
    .A1(net1309),
    .S(net1303),
    .X(_09578_));
 sg13g2_nand2b_1 _28639_ (.Y(_09579_),
    .B(_09578_),
    .A_N(_09548_));
 sg13g2_nand2b_1 _28640_ (.Y(_09580_),
    .B(_10222_),
    .A_N(_09567_));
 sg13g2_nand3_1 _28641_ (.B(_09579_),
    .C(_09580_),
    .A(_09546_),
    .Y(_09581_));
 sg13g2_o21ai_1 _28642_ (.B1(_09581_),
    .Y(_09582_),
    .A1(_07854_),
    .A2(_09547_));
 sg13g2_nor2_1 _28643_ (.A(net790),
    .B(_09582_),
    .Y(_02516_));
 sg13g2_nor2_1 _28644_ (.A(_09903_),
    .B(_10064_),
    .Y(_09583_));
 sg13g2_o21ai_1 _28645_ (.B1(net857),
    .Y(_09584_),
    .A1(net2),
    .A2(_09931_));
 sg13g2_a21oi_1 _28646_ (.A1(_09931_),
    .A2(_09583_),
    .Y(_02517_),
    .B1(_09584_));
 sg13g2_buf_1 _28647_ (.A(_07596_),
    .X(_09585_));
 sg13g2_mux2_1 _28648_ (.A0(_10014_),
    .A1(_07560_),
    .S(net1303),
    .X(_09586_));
 sg13g2_nor2_1 _28649_ (.A(_09723_),
    .B(net875),
    .Y(_09587_));
 sg13g2_a21oi_1 _28650_ (.A1(net875),
    .A2(_09586_),
    .Y(_09588_),
    .B1(_09587_));
 sg13g2_nor2_1 _28651_ (.A(net1272),
    .B(_09588_),
    .Y(_09589_));
 sg13g2_a21oi_1 _28652_ (.A1(net877),
    .A2(net129),
    .Y(_09590_),
    .B1(_09589_));
 sg13g2_nor2_1 _28653_ (.A(net790),
    .B(_09590_),
    .Y(_02518_));
 sg13g2_o21ai_1 _28654_ (.B1(net875),
    .Y(_09591_),
    .A1(net531),
    .A2(_09480_));
 sg13g2_mux2_1 _28655_ (.A0(net1299),
    .A1(net573),
    .S(net1303),
    .X(_09592_));
 sg13g2_a221oi_1 _28656_ (.B2(net875),
    .C1(net1272),
    .B1(_09592_),
    .A1(_07507_),
    .Y(_09593_),
    .A2(_09591_));
 sg13g2_a21oi_1 _28657_ (.A1(_09484_),
    .A2(_07530_),
    .Y(_09594_),
    .B1(_09593_));
 sg13g2_and2_1 _28658_ (.A(_09214_),
    .B(_09594_),
    .X(_02519_));
 sg13g2_nand3_1 _28659_ (.B(net1303),
    .C(_07533_),
    .A(net1283),
    .Y(_09595_));
 sg13g2_nand2_1 _28660_ (.Y(_09596_),
    .A(net1301),
    .B(_09567_));
 sg13g2_nand3_1 _28661_ (.B(_09595_),
    .C(_09596_),
    .A(net875),
    .Y(_09597_));
 sg13g2_o21ai_1 _28662_ (.B1(_09597_),
    .Y(_09598_),
    .A1(_09712_),
    .A2(net875));
 sg13g2_nor2_1 _28663_ (.A(net1272),
    .B(_09598_),
    .Y(_09599_));
 sg13g2_a21oi_1 _28664_ (.A1(net877),
    .A2(net128),
    .Y(_09600_),
    .B1(_09599_));
 sg13g2_nor2_1 _28665_ (.A(net790),
    .B(_09600_),
    .Y(_02520_));
 sg13g2_nand2_1 _28666_ (.Y(_09601_),
    .A(_10016_),
    .B(_09567_));
 sg13g2_o21ai_1 _28667_ (.B1(_09601_),
    .Y(_09602_),
    .A1(_07488_),
    .A2(_09567_));
 sg13g2_nor2b_1 _28668_ (.A(_09602_),
    .B_N(net875),
    .Y(_09603_));
 sg13g2_nand2b_1 _28669_ (.Y(_09604_),
    .B(_07297_),
    .A_N(_09567_));
 sg13g2_a21oi_1 _28670_ (.A1(net875),
    .A2(_09604_),
    .Y(_09605_),
    .B1(_09654_));
 sg13g2_nor3_1 _28671_ (.A(_10075_),
    .B(_09603_),
    .C(_09605_),
    .Y(_09606_));
 sg13g2_a21oi_1 _28672_ (.A1(_09478_),
    .A2(net125),
    .Y(_09607_),
    .B1(_09606_));
 sg13g2_nor2_1 _28673_ (.A(_09345_),
    .B(_09607_),
    .Y(_02521_));
 sg13g2_nand3_1 _28674_ (.B(_09923_),
    .C(_07488_),
    .A(_07475_),
    .Y(_09608_));
 sg13g2_o21ai_1 _28675_ (.B1(_09608_),
    .Y(_09609_),
    .A1(net1303),
    .A2(_10022_));
 sg13g2_o21ai_1 _28676_ (.B1(_09585_),
    .Y(_09610_),
    .A1(_09480_),
    .A2(_07488_));
 sg13g2_a221oi_1 _28677_ (.B2(_07476_),
    .C1(_10075_),
    .B1(_09610_),
    .A1(_09585_),
    .Y(_09611_),
    .A2(_09609_));
 sg13g2_a21oi_1 _28678_ (.A1(_09478_),
    .A2(net141),
    .Y(_09612_),
    .B1(_09611_));
 sg13g2_nor2_1 _28679_ (.A(_09345_),
    .B(_09612_),
    .Y(_02522_));
 sg13g2_mux2_1 _28680_ (.A0(_09928_),
    .A1(\mem.mem_io.porta_out[0] ),
    .S(\mem.mem_io.porta_oe[0] ),
    .X(net29));
 sg13g2_mux2_1 _28681_ (.A0(_09929_),
    .A1(\mem.mem_io.porta_out[1] ),
    .S(\mem.mem_io.porta_oe[1] ),
    .X(net30));
 sg13g2_nand2_1 _28682_ (.Y(_09613_),
    .A(\mem.mem_io.porta_out[2] ),
    .B(_09303_));
 sg13g2_o21ai_1 _28683_ (.B1(_09613_),
    .Y(net31),
    .A1(_09935_),
    .A2(_09303_));
 sg13g2_mux2_1 _28684_ (.A0(o_shift_out),
    .A1(\mem.mem_io.porta_out[3] ),
    .S(\mem.mem_io.porta_oe[3] ),
    .X(net32));
 sg13g2_and2_1 _28685_ (.A(\mem.mem_io.porta_out[4] ),
    .B(\mem.mem_io.porta_oe[4] ),
    .X(net33));
 sg13g2_and2_1 _28686_ (.A(\mem.mem_io.porta_out[5] ),
    .B(\mem.mem_io.porta_oe[5] ),
    .X(net34));
 sg13g2_and2_1 _28687_ (.A(\mem.mem_io.porta_out[6] ),
    .B(\mem.mem_io.porta_oe[6] ),
    .X(net35));
 sg13g2_and2_1 _28688_ (.A(\mem.mem_io.porta_out[7] ),
    .B(\mem.mem_io.porta_oe[7] ),
    .X(net36));
 sg13g2_dfrbp_1 _28689_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1312),
    .D(_00015_),
    .Q_N(_15692_),
    .Q(_00000_));
 sg13g2_dfrbp_1 _28690_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1313),
    .D(_00016_),
    .Q_N(_15693_),
    .Q(_00001_));
 sg13g2_dfrbp_1 _28691_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1314),
    .D(_00017_),
    .Q_N(_15694_),
    .Q(_00002_));
 sg13g2_dfrbp_1 _28692_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1315),
    .D(_00018_),
    .Q_N(_15695_),
    .Q(_00003_));
 sg13g2_dfrbp_1 _28693_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1316),
    .D(_00019_),
    .Q_N(_15696_),
    .Q(_00004_));
 sg13g2_dfrbp_1 _28694_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1317),
    .D(_00020_),
    .Q_N(_15697_),
    .Q(_00005_));
 sg13g2_dfrbp_1 _28695_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1318),
    .D(_00021_),
    .Q_N(_15698_),
    .Q(_00006_));
 sg13g2_dfrbp_1 _28696_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1319),
    .D(_00022_),
    .Q_N(_15691_),
    .Q(_00007_));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_dfrbp_1 \delay_counter[0]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1320),
    .D(_00082_),
    .Q_N(_15690_),
    .Q(\delay_counter[0] ));
 sg13g2_dfrbp_1 \delay_counter[1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1321),
    .D(_00083_),
    .Q_N(_15689_),
    .Q(\delay_counter[1] ));
 sg13g2_dfrbp_1 \delay_counter[2]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1322),
    .D(_00084_),
    .Q_N(_15688_),
    .Q(\delay_counter[2] ));
 sg13g2_dfrbp_1 \delay_counter[3]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1323),
    .D(_00085_),
    .Q_N(_15687_),
    .Q(\delay_counter[3] ));
 sg13g2_dfrbp_1 \delay_counter[4]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1324),
    .D(_00086_),
    .Q_N(_15686_),
    .Q(\delay_counter[4] ));
 sg13g2_dfrbp_1 \delay_counter[5]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1325),
    .D(_00087_),
    .Q_N(_15685_),
    .Q(\delay_counter[5] ));
 sg13g2_dfrbp_1 \delay_counter[6]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1326),
    .D(_00088_),
    .Q_N(_15684_),
    .Q(\delay_counter[6] ));
 sg13g2_dfrbp_1 \delay_counter[7]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1327),
    .D(_00089_),
    .Q_N(_15683_),
    .Q(\delay_counter[7] ));
 sg13g2_dfrbp_1 \delay_cycles[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1328),
    .D(_00090_),
    .Q_N(_15682_),
    .Q(\delay_cycles[0] ));
 sg13g2_dfrbp_1 \delay_cycles[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1329),
    .D(_00091_),
    .Q_N(_15681_),
    .Q(\delay_cycles[10] ));
 sg13g2_dfrbp_1 \delay_cycles[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1330),
    .D(_00092_),
    .Q_N(_15680_),
    .Q(\delay_cycles[11] ));
 sg13g2_dfrbp_1 \delay_cycles[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1331),
    .D(_00093_),
    .Q_N(_15679_),
    .Q(\delay_cycles[12] ));
 sg13g2_dfrbp_1 \delay_cycles[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1332),
    .D(_00094_),
    .Q_N(_15678_),
    .Q(\delay_cycles[13] ));
 sg13g2_dfrbp_1 \delay_cycles[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1333),
    .D(_00095_),
    .Q_N(_15677_),
    .Q(\delay_cycles[14] ));
 sg13g2_dfrbp_1 \delay_cycles[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1334),
    .D(_00096_),
    .Q_N(_15676_),
    .Q(\delay_cycles[15] ));
 sg13g2_dfrbp_1 \delay_cycles[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1335),
    .D(_00097_),
    .Q_N(_15675_),
    .Q(\delay_cycles[16] ));
 sg13g2_dfrbp_1 \delay_cycles[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1336),
    .D(_00098_),
    .Q_N(_15674_),
    .Q(\delay_cycles[17] ));
 sg13g2_dfrbp_1 \delay_cycles[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1337),
    .D(_00099_),
    .Q_N(_15673_),
    .Q(\delay_cycles[18] ));
 sg13g2_dfrbp_1 \delay_cycles[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1338),
    .D(_00100_),
    .Q_N(_15672_),
    .Q(\delay_cycles[19] ));
 sg13g2_dfrbp_1 \delay_cycles[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1339),
    .D(_00101_),
    .Q_N(_15671_),
    .Q(\delay_cycles[1] ));
 sg13g2_dfrbp_1 \delay_cycles[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1340),
    .D(_00102_),
    .Q_N(_15670_),
    .Q(\delay_cycles[20] ));
 sg13g2_dfrbp_1 \delay_cycles[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1341),
    .D(_00103_),
    .Q_N(_15669_),
    .Q(\delay_cycles[21] ));
 sg13g2_dfrbp_1 \delay_cycles[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1342),
    .D(_00104_),
    .Q_N(_15668_),
    .Q(\delay_cycles[22] ));
 sg13g2_dfrbp_1 \delay_cycles[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1343),
    .D(_00105_),
    .Q_N(_15667_),
    .Q(\delay_cycles[23] ));
 sg13g2_dfrbp_1 \delay_cycles[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1344),
    .D(_00106_),
    .Q_N(_15666_),
    .Q(\delay_cycles[2] ));
 sg13g2_dfrbp_1 \delay_cycles[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1345),
    .D(_00107_),
    .Q_N(_15665_),
    .Q(\delay_cycles[3] ));
 sg13g2_dfrbp_1 \delay_cycles[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1346),
    .D(_00108_),
    .Q_N(_15664_),
    .Q(\delay_cycles[4] ));
 sg13g2_dfrbp_1 \delay_cycles[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1347),
    .D(_00109_),
    .Q_N(_15663_),
    .Q(\delay_cycles[5] ));
 sg13g2_dfrbp_1 \delay_cycles[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1348),
    .D(_00110_),
    .Q_N(_15662_),
    .Q(\delay_cycles[6] ));
 sg13g2_dfrbp_1 \delay_cycles[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1349),
    .D(_00111_),
    .Q_N(_15661_),
    .Q(\delay_cycles[7] ));
 sg13g2_dfrbp_1 \delay_cycles[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1350),
    .D(_00112_),
    .Q_N(_15660_),
    .Q(\delay_cycles[8] ));
 sg13g2_dfrbp_1 \delay_cycles[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1351),
    .D(_00113_),
    .Q_N(_15659_),
    .Q(\delay_cycles[9] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1352),
    .D(_00114_),
    .Q_N(_15658_),
    .Q(\mem.mem_internal.code_mem[0][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1353),
    .D(_00115_),
    .Q_N(_15657_),
    .Q(\mem.mem_internal.code_mem[0][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[0][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1354),
    .D(_00116_),
    .Q_N(_15656_),
    .Q(\mem.mem_internal.code_mem[0][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1355),
    .D(_00117_),
    .Q_N(_15655_),
    .Q(\mem.mem_internal.code_mem[0][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[0][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1356),
    .D(_00118_),
    .Q_N(_15654_),
    .Q(\mem.mem_internal.code_mem[0][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[0][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1357),
    .D(_00119_),
    .Q_N(_15653_),
    .Q(\mem.mem_internal.code_mem[0][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[0][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1358),
    .D(_00120_),
    .Q_N(_15652_),
    .Q(\mem.mem_internal.code_mem[0][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[0][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1359),
    .D(_00121_),
    .Q_N(_15651_),
    .Q(\mem.mem_internal.code_mem[0][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[100][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1360),
    .D(_00122_),
    .Q_N(_15650_),
    .Q(\mem.mem_internal.code_mem[100][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[100][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1361),
    .D(_00123_),
    .Q_N(_15649_),
    .Q(\mem.mem_internal.code_mem[100][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[100][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1362),
    .D(_00124_),
    .Q_N(_15648_),
    .Q(\mem.mem_internal.code_mem[100][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[100][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1363),
    .D(_00125_),
    .Q_N(_15647_),
    .Q(\mem.mem_internal.code_mem[100][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[100][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1364),
    .D(_00126_),
    .Q_N(_15646_),
    .Q(\mem.mem_internal.code_mem[100][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[100][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1365),
    .D(_00127_),
    .Q_N(_15645_),
    .Q(\mem.mem_internal.code_mem[100][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[100][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1366),
    .D(_00128_),
    .Q_N(_15644_),
    .Q(\mem.mem_internal.code_mem[100][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[100][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1367),
    .D(_00129_),
    .Q_N(_15643_),
    .Q(\mem.mem_internal.code_mem[100][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[101][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1368),
    .D(_00130_),
    .Q_N(_15642_),
    .Q(\mem.mem_internal.code_mem[101][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[101][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1369),
    .D(_00131_),
    .Q_N(_15641_),
    .Q(\mem.mem_internal.code_mem[101][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[101][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1370),
    .D(_00132_),
    .Q_N(_15640_),
    .Q(\mem.mem_internal.code_mem[101][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[101][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1371),
    .D(_00133_),
    .Q_N(_15639_),
    .Q(\mem.mem_internal.code_mem[101][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[101][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1372),
    .D(_00134_),
    .Q_N(_15638_),
    .Q(\mem.mem_internal.code_mem[101][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[101][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1373),
    .D(_00135_),
    .Q_N(_15637_),
    .Q(\mem.mem_internal.code_mem[101][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[101][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1374),
    .D(_00136_),
    .Q_N(_15636_),
    .Q(\mem.mem_internal.code_mem[101][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[101][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1375),
    .D(_00137_),
    .Q_N(_15635_),
    .Q(\mem.mem_internal.code_mem[101][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[102][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1376),
    .D(_00138_),
    .Q_N(_15634_),
    .Q(\mem.mem_internal.code_mem[102][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[102][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1377),
    .D(_00139_),
    .Q_N(_15633_),
    .Q(\mem.mem_internal.code_mem[102][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[102][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1378),
    .D(_00140_),
    .Q_N(_15632_),
    .Q(\mem.mem_internal.code_mem[102][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[102][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1379),
    .D(_00141_),
    .Q_N(_15631_),
    .Q(\mem.mem_internal.code_mem[102][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[102][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1380),
    .D(_00142_),
    .Q_N(_15630_),
    .Q(\mem.mem_internal.code_mem[102][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[102][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1381),
    .D(_00143_),
    .Q_N(_15629_),
    .Q(\mem.mem_internal.code_mem[102][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[102][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1382),
    .D(_00144_),
    .Q_N(_15628_),
    .Q(\mem.mem_internal.code_mem[102][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[102][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1383),
    .D(_00145_),
    .Q_N(_15627_),
    .Q(\mem.mem_internal.code_mem[102][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[103][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1384),
    .D(_00146_),
    .Q_N(_15626_),
    .Q(\mem.mem_internal.code_mem[103][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[103][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1385),
    .D(_00147_),
    .Q_N(_15625_),
    .Q(\mem.mem_internal.code_mem[103][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[103][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1386),
    .D(_00148_),
    .Q_N(_15624_),
    .Q(\mem.mem_internal.code_mem[103][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[103][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1387),
    .D(_00149_),
    .Q_N(_15623_),
    .Q(\mem.mem_internal.code_mem[103][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[103][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1388),
    .D(_00150_),
    .Q_N(_15622_),
    .Q(\mem.mem_internal.code_mem[103][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[103][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1389),
    .D(_00151_),
    .Q_N(_15621_),
    .Q(\mem.mem_internal.code_mem[103][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[103][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1390),
    .D(_00152_),
    .Q_N(_15620_),
    .Q(\mem.mem_internal.code_mem[103][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[103][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1391),
    .D(_00153_),
    .Q_N(_15619_),
    .Q(\mem.mem_internal.code_mem[103][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[104][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1392),
    .D(_00154_),
    .Q_N(_15618_),
    .Q(\mem.mem_internal.code_mem[104][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[104][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1393),
    .D(_00155_),
    .Q_N(_15617_),
    .Q(\mem.mem_internal.code_mem[104][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[104][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1394),
    .D(_00156_),
    .Q_N(_15616_),
    .Q(\mem.mem_internal.code_mem[104][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[104][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1395),
    .D(_00157_),
    .Q_N(_15615_),
    .Q(\mem.mem_internal.code_mem[104][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[104][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1396),
    .D(_00158_),
    .Q_N(_15614_),
    .Q(\mem.mem_internal.code_mem[104][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[104][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1397),
    .D(_00159_),
    .Q_N(_15613_),
    .Q(\mem.mem_internal.code_mem[104][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[104][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1398),
    .D(_00160_),
    .Q_N(_15612_),
    .Q(\mem.mem_internal.code_mem[104][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[104][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1399),
    .D(_00161_),
    .Q_N(_15611_),
    .Q(\mem.mem_internal.code_mem[104][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[105][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1400),
    .D(_00162_),
    .Q_N(_15610_),
    .Q(\mem.mem_internal.code_mem[105][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[105][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1401),
    .D(_00163_),
    .Q_N(_15609_),
    .Q(\mem.mem_internal.code_mem[105][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[105][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1402),
    .D(_00164_),
    .Q_N(_15608_),
    .Q(\mem.mem_internal.code_mem[105][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[105][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1403),
    .D(_00165_),
    .Q_N(_15607_),
    .Q(\mem.mem_internal.code_mem[105][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[105][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1404),
    .D(_00166_),
    .Q_N(_15606_),
    .Q(\mem.mem_internal.code_mem[105][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[105][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1405),
    .D(_00167_),
    .Q_N(_15605_),
    .Q(\mem.mem_internal.code_mem[105][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[105][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1406),
    .D(_00168_),
    .Q_N(_15604_),
    .Q(\mem.mem_internal.code_mem[105][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[105][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1407),
    .D(_00169_),
    .Q_N(_15603_),
    .Q(\mem.mem_internal.code_mem[105][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[106][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1408),
    .D(_00170_),
    .Q_N(_15602_),
    .Q(\mem.mem_internal.code_mem[106][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[106][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1409),
    .D(_00171_),
    .Q_N(_15601_),
    .Q(\mem.mem_internal.code_mem[106][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[106][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1410),
    .D(_00172_),
    .Q_N(_15600_),
    .Q(\mem.mem_internal.code_mem[106][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[106][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1411),
    .D(_00173_),
    .Q_N(_15599_),
    .Q(\mem.mem_internal.code_mem[106][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[106][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1412),
    .D(_00174_),
    .Q_N(_15598_),
    .Q(\mem.mem_internal.code_mem[106][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[106][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1413),
    .D(_00175_),
    .Q_N(_15597_),
    .Q(\mem.mem_internal.code_mem[106][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[106][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1414),
    .D(_00176_),
    .Q_N(_15596_),
    .Q(\mem.mem_internal.code_mem[106][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[106][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1415),
    .D(_00177_),
    .Q_N(_15595_),
    .Q(\mem.mem_internal.code_mem[106][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[107][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1416),
    .D(_00178_),
    .Q_N(_15594_),
    .Q(\mem.mem_internal.code_mem[107][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[107][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1417),
    .D(_00179_),
    .Q_N(_15593_),
    .Q(\mem.mem_internal.code_mem[107][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[107][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1418),
    .D(_00180_),
    .Q_N(_15592_),
    .Q(\mem.mem_internal.code_mem[107][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[107][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1419),
    .D(_00181_),
    .Q_N(_15591_),
    .Q(\mem.mem_internal.code_mem[107][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[107][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1420),
    .D(_00182_),
    .Q_N(_15590_),
    .Q(\mem.mem_internal.code_mem[107][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[107][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1421),
    .D(_00183_),
    .Q_N(_15589_),
    .Q(\mem.mem_internal.code_mem[107][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[107][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1422),
    .D(_00184_),
    .Q_N(_15588_),
    .Q(\mem.mem_internal.code_mem[107][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[107][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1423),
    .D(_00185_),
    .Q_N(_15587_),
    .Q(\mem.mem_internal.code_mem[107][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[108][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1424),
    .D(_00186_),
    .Q_N(_15586_),
    .Q(\mem.mem_internal.code_mem[108][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[108][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1425),
    .D(_00187_),
    .Q_N(_15585_),
    .Q(\mem.mem_internal.code_mem[108][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[108][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1426),
    .D(_00188_),
    .Q_N(_15584_),
    .Q(\mem.mem_internal.code_mem[108][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[108][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1427),
    .D(_00189_),
    .Q_N(_15583_),
    .Q(\mem.mem_internal.code_mem[108][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[108][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1428),
    .D(_00190_),
    .Q_N(_15582_),
    .Q(\mem.mem_internal.code_mem[108][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[108][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1429),
    .D(_00191_),
    .Q_N(_15581_),
    .Q(\mem.mem_internal.code_mem[108][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[108][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1430),
    .D(_00192_),
    .Q_N(_15580_),
    .Q(\mem.mem_internal.code_mem[108][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[108][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1431),
    .D(_00193_),
    .Q_N(_15579_),
    .Q(\mem.mem_internal.code_mem[108][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[109][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1432),
    .D(_00194_),
    .Q_N(_15578_),
    .Q(\mem.mem_internal.code_mem[109][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[109][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1433),
    .D(_00195_),
    .Q_N(_15577_),
    .Q(\mem.mem_internal.code_mem[109][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[109][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1434),
    .D(_00196_),
    .Q_N(_15576_),
    .Q(\mem.mem_internal.code_mem[109][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[109][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1435),
    .D(_00197_),
    .Q_N(_15575_),
    .Q(\mem.mem_internal.code_mem[109][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[109][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1436),
    .D(_00198_),
    .Q_N(_15574_),
    .Q(\mem.mem_internal.code_mem[109][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[109][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1437),
    .D(_00199_),
    .Q_N(_15573_),
    .Q(\mem.mem_internal.code_mem[109][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[109][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1438),
    .D(_00200_),
    .Q_N(_15572_),
    .Q(\mem.mem_internal.code_mem[109][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[109][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1439),
    .D(_00201_),
    .Q_N(_15571_),
    .Q(\mem.mem_internal.code_mem[109][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[10][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1440),
    .D(_00202_),
    .Q_N(_15570_),
    .Q(\mem.mem_internal.code_mem[10][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[10][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1441),
    .D(_00203_),
    .Q_N(_15569_),
    .Q(\mem.mem_internal.code_mem[10][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[10][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1442),
    .D(_00204_),
    .Q_N(_15568_),
    .Q(\mem.mem_internal.code_mem[10][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[10][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1443),
    .D(_00205_),
    .Q_N(_15567_),
    .Q(\mem.mem_internal.code_mem[10][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[10][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1444),
    .D(_00206_),
    .Q_N(_15566_),
    .Q(\mem.mem_internal.code_mem[10][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[10][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1445),
    .D(_00207_),
    .Q_N(_15565_),
    .Q(\mem.mem_internal.code_mem[10][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[10][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1446),
    .D(_00208_),
    .Q_N(_15564_),
    .Q(\mem.mem_internal.code_mem[10][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[10][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1447),
    .D(_00209_),
    .Q_N(_15563_),
    .Q(\mem.mem_internal.code_mem[10][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[110][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1448),
    .D(_00210_),
    .Q_N(_15562_),
    .Q(\mem.mem_internal.code_mem[110][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[110][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1449),
    .D(_00211_),
    .Q_N(_15561_),
    .Q(\mem.mem_internal.code_mem[110][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[110][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1450),
    .D(_00212_),
    .Q_N(_15560_),
    .Q(\mem.mem_internal.code_mem[110][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[110][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1451),
    .D(_00213_),
    .Q_N(_15559_),
    .Q(\mem.mem_internal.code_mem[110][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[110][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1452),
    .D(_00214_),
    .Q_N(_15558_),
    .Q(\mem.mem_internal.code_mem[110][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[110][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1453),
    .D(_00215_),
    .Q_N(_15557_),
    .Q(\mem.mem_internal.code_mem[110][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[110][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1454),
    .D(_00216_),
    .Q_N(_15556_),
    .Q(\mem.mem_internal.code_mem[110][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[110][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1455),
    .D(_00217_),
    .Q_N(_15555_),
    .Q(\mem.mem_internal.code_mem[110][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[111][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1456),
    .D(_00218_),
    .Q_N(_15554_),
    .Q(\mem.mem_internal.code_mem[111][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[111][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1457),
    .D(_00219_),
    .Q_N(_15553_),
    .Q(\mem.mem_internal.code_mem[111][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[111][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1458),
    .D(_00220_),
    .Q_N(_15552_),
    .Q(\mem.mem_internal.code_mem[111][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[111][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1459),
    .D(_00221_),
    .Q_N(_15551_),
    .Q(\mem.mem_internal.code_mem[111][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[111][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1460),
    .D(_00222_),
    .Q_N(_15550_),
    .Q(\mem.mem_internal.code_mem[111][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[111][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1461),
    .D(_00223_),
    .Q_N(_15549_),
    .Q(\mem.mem_internal.code_mem[111][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[111][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1462),
    .D(_00224_),
    .Q_N(_15548_),
    .Q(\mem.mem_internal.code_mem[111][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[111][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1463),
    .D(_00225_),
    .Q_N(_15547_),
    .Q(\mem.mem_internal.code_mem[111][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[112][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1464),
    .D(_00226_),
    .Q_N(_15546_),
    .Q(\mem.mem_internal.code_mem[112][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[112][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1465),
    .D(_00227_),
    .Q_N(_15545_),
    .Q(\mem.mem_internal.code_mem[112][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[112][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1466),
    .D(_00228_),
    .Q_N(_15544_),
    .Q(\mem.mem_internal.code_mem[112][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[112][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1467),
    .D(_00229_),
    .Q_N(_15543_),
    .Q(\mem.mem_internal.code_mem[112][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[112][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1468),
    .D(_00230_),
    .Q_N(_15542_),
    .Q(\mem.mem_internal.code_mem[112][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[112][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1469),
    .D(_00231_),
    .Q_N(_15541_),
    .Q(\mem.mem_internal.code_mem[112][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[112][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1470),
    .D(_00232_),
    .Q_N(_15540_),
    .Q(\mem.mem_internal.code_mem[112][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[112][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1471),
    .D(_00233_),
    .Q_N(_15539_),
    .Q(\mem.mem_internal.code_mem[112][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[113][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1472),
    .D(_00234_),
    .Q_N(_15538_),
    .Q(\mem.mem_internal.code_mem[113][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[113][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1473),
    .D(_00235_),
    .Q_N(_15537_),
    .Q(\mem.mem_internal.code_mem[113][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[113][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1474),
    .D(_00236_),
    .Q_N(_15536_),
    .Q(\mem.mem_internal.code_mem[113][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[113][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1475),
    .D(_00237_),
    .Q_N(_15535_),
    .Q(\mem.mem_internal.code_mem[113][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[113][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1476),
    .D(_00238_),
    .Q_N(_15534_),
    .Q(\mem.mem_internal.code_mem[113][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[113][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1477),
    .D(_00239_),
    .Q_N(_15533_),
    .Q(\mem.mem_internal.code_mem[113][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[113][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1478),
    .D(_00240_),
    .Q_N(_15532_),
    .Q(\mem.mem_internal.code_mem[113][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[113][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1479),
    .D(_00241_),
    .Q_N(_15531_),
    .Q(\mem.mem_internal.code_mem[113][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[114][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1480),
    .D(_00242_),
    .Q_N(_15530_),
    .Q(\mem.mem_internal.code_mem[114][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[114][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1481),
    .D(_00243_),
    .Q_N(_15529_),
    .Q(\mem.mem_internal.code_mem[114][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[114][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1482),
    .D(_00244_),
    .Q_N(_15528_),
    .Q(\mem.mem_internal.code_mem[114][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[114][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1483),
    .D(_00245_),
    .Q_N(_15527_),
    .Q(\mem.mem_internal.code_mem[114][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[114][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1484),
    .D(_00246_),
    .Q_N(_15526_),
    .Q(\mem.mem_internal.code_mem[114][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[114][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1485),
    .D(_00247_),
    .Q_N(_15525_),
    .Q(\mem.mem_internal.code_mem[114][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[114][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1486),
    .D(_00248_),
    .Q_N(_15524_),
    .Q(\mem.mem_internal.code_mem[114][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[114][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1487),
    .D(_00249_),
    .Q_N(_15523_),
    .Q(\mem.mem_internal.code_mem[114][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[115][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1488),
    .D(_00250_),
    .Q_N(_15522_),
    .Q(\mem.mem_internal.code_mem[115][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[115][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1489),
    .D(_00251_),
    .Q_N(_15521_),
    .Q(\mem.mem_internal.code_mem[115][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[115][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1490),
    .D(_00252_),
    .Q_N(_15520_),
    .Q(\mem.mem_internal.code_mem[115][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[115][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1491),
    .D(_00253_),
    .Q_N(_15519_),
    .Q(\mem.mem_internal.code_mem[115][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[115][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1492),
    .D(_00254_),
    .Q_N(_15518_),
    .Q(\mem.mem_internal.code_mem[115][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[115][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1493),
    .D(_00255_),
    .Q_N(_15517_),
    .Q(\mem.mem_internal.code_mem[115][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[115][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1494),
    .D(_00256_),
    .Q_N(_15516_),
    .Q(\mem.mem_internal.code_mem[115][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[115][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1495),
    .D(_00257_),
    .Q_N(_15515_),
    .Q(\mem.mem_internal.code_mem[115][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[116][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1496),
    .D(_00258_),
    .Q_N(_15514_),
    .Q(\mem.mem_internal.code_mem[116][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[116][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1497),
    .D(_00259_),
    .Q_N(_15513_),
    .Q(\mem.mem_internal.code_mem[116][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[116][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1498),
    .D(_00260_),
    .Q_N(_15512_),
    .Q(\mem.mem_internal.code_mem[116][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[116][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1499),
    .D(_00261_),
    .Q_N(_15511_),
    .Q(\mem.mem_internal.code_mem[116][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[116][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1500),
    .D(_00262_),
    .Q_N(_15510_),
    .Q(\mem.mem_internal.code_mem[116][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[116][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1501),
    .D(_00263_),
    .Q_N(_15509_),
    .Q(\mem.mem_internal.code_mem[116][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[116][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1502),
    .D(_00264_),
    .Q_N(_15508_),
    .Q(\mem.mem_internal.code_mem[116][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[116][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1503),
    .D(_00265_),
    .Q_N(_15507_),
    .Q(\mem.mem_internal.code_mem[116][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[117][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1504),
    .D(_00266_),
    .Q_N(_15506_),
    .Q(\mem.mem_internal.code_mem[117][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[117][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1505),
    .D(_00267_),
    .Q_N(_15505_),
    .Q(\mem.mem_internal.code_mem[117][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[117][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1506),
    .D(_00268_),
    .Q_N(_15504_),
    .Q(\mem.mem_internal.code_mem[117][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[117][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1507),
    .D(_00269_),
    .Q_N(_15503_),
    .Q(\mem.mem_internal.code_mem[117][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[117][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1508),
    .D(_00270_),
    .Q_N(_15502_),
    .Q(\mem.mem_internal.code_mem[117][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[117][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1509),
    .D(_00271_),
    .Q_N(_15501_),
    .Q(\mem.mem_internal.code_mem[117][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[117][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1510),
    .D(_00272_),
    .Q_N(_15500_),
    .Q(\mem.mem_internal.code_mem[117][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[117][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1511),
    .D(_00273_),
    .Q_N(_15499_),
    .Q(\mem.mem_internal.code_mem[117][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[118][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1512),
    .D(_00274_),
    .Q_N(_15498_),
    .Q(\mem.mem_internal.code_mem[118][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[118][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1513),
    .D(_00275_),
    .Q_N(_15497_),
    .Q(\mem.mem_internal.code_mem[118][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[118][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1514),
    .D(_00276_),
    .Q_N(_15496_),
    .Q(\mem.mem_internal.code_mem[118][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[118][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1515),
    .D(_00277_),
    .Q_N(_15495_),
    .Q(\mem.mem_internal.code_mem[118][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[118][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1516),
    .D(_00278_),
    .Q_N(_15494_),
    .Q(\mem.mem_internal.code_mem[118][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[118][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1517),
    .D(_00279_),
    .Q_N(_15493_),
    .Q(\mem.mem_internal.code_mem[118][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[118][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1518),
    .D(_00280_),
    .Q_N(_15492_),
    .Q(\mem.mem_internal.code_mem[118][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[118][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1519),
    .D(_00281_),
    .Q_N(_15491_),
    .Q(\mem.mem_internal.code_mem[118][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[119][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1520),
    .D(_00282_),
    .Q_N(_15490_),
    .Q(\mem.mem_internal.code_mem[119][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[119][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1521),
    .D(_00283_),
    .Q_N(_15489_),
    .Q(\mem.mem_internal.code_mem[119][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[119][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1522),
    .D(_00284_),
    .Q_N(_15488_),
    .Q(\mem.mem_internal.code_mem[119][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[119][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1523),
    .D(_00285_),
    .Q_N(_15487_),
    .Q(\mem.mem_internal.code_mem[119][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[119][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1524),
    .D(_00286_),
    .Q_N(_15486_),
    .Q(\mem.mem_internal.code_mem[119][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[119][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1525),
    .D(_00287_),
    .Q_N(_15485_),
    .Q(\mem.mem_internal.code_mem[119][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[119][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1526),
    .D(_00288_),
    .Q_N(_15484_),
    .Q(\mem.mem_internal.code_mem[119][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[119][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1527),
    .D(_00289_),
    .Q_N(_15483_),
    .Q(\mem.mem_internal.code_mem[119][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[11][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1528),
    .D(_00290_),
    .Q_N(_15482_),
    .Q(\mem.mem_internal.code_mem[11][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[11][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1529),
    .D(_00291_),
    .Q_N(_15481_),
    .Q(\mem.mem_internal.code_mem[11][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[11][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1530),
    .D(_00292_),
    .Q_N(_15480_),
    .Q(\mem.mem_internal.code_mem[11][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[11][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1531),
    .D(_00293_),
    .Q_N(_15479_),
    .Q(\mem.mem_internal.code_mem[11][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[11][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1532),
    .D(_00294_),
    .Q_N(_15478_),
    .Q(\mem.mem_internal.code_mem[11][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[11][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1533),
    .D(_00295_),
    .Q_N(_15477_),
    .Q(\mem.mem_internal.code_mem[11][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[11][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1534),
    .D(_00296_),
    .Q_N(_15476_),
    .Q(\mem.mem_internal.code_mem[11][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[11][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1535),
    .D(_00297_),
    .Q_N(_15475_),
    .Q(\mem.mem_internal.code_mem[11][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[120][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1536),
    .D(_00298_),
    .Q_N(_15474_),
    .Q(\mem.mem_internal.code_mem[120][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[120][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1537),
    .D(_00299_),
    .Q_N(_15473_),
    .Q(\mem.mem_internal.code_mem[120][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[120][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1538),
    .D(_00300_),
    .Q_N(_15472_),
    .Q(\mem.mem_internal.code_mem[120][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[120][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1539),
    .D(_00301_),
    .Q_N(_15471_),
    .Q(\mem.mem_internal.code_mem[120][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[120][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1540),
    .D(_00302_),
    .Q_N(_15470_),
    .Q(\mem.mem_internal.code_mem[120][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[120][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1541),
    .D(_00303_),
    .Q_N(_15469_),
    .Q(\mem.mem_internal.code_mem[120][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[120][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1542),
    .D(_00304_),
    .Q_N(_15468_),
    .Q(\mem.mem_internal.code_mem[120][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[120][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1543),
    .D(_00305_),
    .Q_N(_15467_),
    .Q(\mem.mem_internal.code_mem[120][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[121][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1544),
    .D(_00306_),
    .Q_N(_15466_),
    .Q(\mem.mem_internal.code_mem[121][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[121][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1545),
    .D(_00307_),
    .Q_N(_15465_),
    .Q(\mem.mem_internal.code_mem[121][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[121][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1546),
    .D(_00308_),
    .Q_N(_15464_),
    .Q(\mem.mem_internal.code_mem[121][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[121][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1547),
    .D(_00309_),
    .Q_N(_15463_),
    .Q(\mem.mem_internal.code_mem[121][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[121][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1548),
    .D(_00310_),
    .Q_N(_15462_),
    .Q(\mem.mem_internal.code_mem[121][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[121][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1549),
    .D(_00311_),
    .Q_N(_15461_),
    .Q(\mem.mem_internal.code_mem[121][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[121][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1550),
    .D(_00312_),
    .Q_N(_15460_),
    .Q(\mem.mem_internal.code_mem[121][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[121][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1551),
    .D(_00313_),
    .Q_N(_15459_),
    .Q(\mem.mem_internal.code_mem[121][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[122][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1552),
    .D(_00314_),
    .Q_N(_15458_),
    .Q(\mem.mem_internal.code_mem[122][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[122][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1553),
    .D(_00315_),
    .Q_N(_15457_),
    .Q(\mem.mem_internal.code_mem[122][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[122][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1554),
    .D(_00316_),
    .Q_N(_15456_),
    .Q(\mem.mem_internal.code_mem[122][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[122][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1555),
    .D(_00317_),
    .Q_N(_15455_),
    .Q(\mem.mem_internal.code_mem[122][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[122][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1556),
    .D(_00318_),
    .Q_N(_15454_),
    .Q(\mem.mem_internal.code_mem[122][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[122][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1557),
    .D(_00319_),
    .Q_N(_15453_),
    .Q(\mem.mem_internal.code_mem[122][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[122][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1558),
    .D(_00320_),
    .Q_N(_15452_),
    .Q(\mem.mem_internal.code_mem[122][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[122][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1559),
    .D(_00321_),
    .Q_N(_15451_),
    .Q(\mem.mem_internal.code_mem[122][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[123][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1560),
    .D(_00322_),
    .Q_N(_15450_),
    .Q(\mem.mem_internal.code_mem[123][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[123][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1561),
    .D(_00323_),
    .Q_N(_15449_),
    .Q(\mem.mem_internal.code_mem[123][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[123][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1562),
    .D(_00324_),
    .Q_N(_15448_),
    .Q(\mem.mem_internal.code_mem[123][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[123][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1563),
    .D(_00325_),
    .Q_N(_15447_),
    .Q(\mem.mem_internal.code_mem[123][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[123][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1564),
    .D(_00326_),
    .Q_N(_15446_),
    .Q(\mem.mem_internal.code_mem[123][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[123][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1565),
    .D(_00327_),
    .Q_N(_15445_),
    .Q(\mem.mem_internal.code_mem[123][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[123][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1566),
    .D(_00328_),
    .Q_N(_15444_),
    .Q(\mem.mem_internal.code_mem[123][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[123][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1567),
    .D(_00329_),
    .Q_N(_15443_),
    .Q(\mem.mem_internal.code_mem[123][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[124][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1568),
    .D(_00330_),
    .Q_N(_15442_),
    .Q(\mem.mem_internal.code_mem[124][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[124][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1569),
    .D(_00331_),
    .Q_N(_15441_),
    .Q(\mem.mem_internal.code_mem[124][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[124][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1570),
    .D(_00332_),
    .Q_N(_15440_),
    .Q(\mem.mem_internal.code_mem[124][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[124][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1571),
    .D(_00333_),
    .Q_N(_15439_),
    .Q(\mem.mem_internal.code_mem[124][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[124][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1572),
    .D(_00334_),
    .Q_N(_15438_),
    .Q(\mem.mem_internal.code_mem[124][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[124][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1573),
    .D(_00335_),
    .Q_N(_15437_),
    .Q(\mem.mem_internal.code_mem[124][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[124][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1574),
    .D(_00336_),
    .Q_N(_15436_),
    .Q(\mem.mem_internal.code_mem[124][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[124][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1575),
    .D(_00337_),
    .Q_N(_15435_),
    .Q(\mem.mem_internal.code_mem[124][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[125][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1576),
    .D(_00338_),
    .Q_N(_15434_),
    .Q(\mem.mem_internal.code_mem[125][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[125][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1577),
    .D(_00339_),
    .Q_N(_15433_),
    .Q(\mem.mem_internal.code_mem[125][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[125][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1578),
    .D(_00340_),
    .Q_N(_15432_),
    .Q(\mem.mem_internal.code_mem[125][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[125][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1579),
    .D(_00341_),
    .Q_N(_15431_),
    .Q(\mem.mem_internal.code_mem[125][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[125][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1580),
    .D(_00342_),
    .Q_N(_15430_),
    .Q(\mem.mem_internal.code_mem[125][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[125][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1581),
    .D(_00343_),
    .Q_N(_15429_),
    .Q(\mem.mem_internal.code_mem[125][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[125][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1582),
    .D(_00344_),
    .Q_N(_15428_),
    .Q(\mem.mem_internal.code_mem[125][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[125][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1583),
    .D(_00345_),
    .Q_N(_15427_),
    .Q(\mem.mem_internal.code_mem[125][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[126][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1584),
    .D(_00346_),
    .Q_N(_15426_),
    .Q(\mem.mem_internal.code_mem[126][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[126][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1585),
    .D(_00347_),
    .Q_N(_15425_),
    .Q(\mem.mem_internal.code_mem[126][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[126][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1586),
    .D(_00348_),
    .Q_N(_15424_),
    .Q(\mem.mem_internal.code_mem[126][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[126][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1587),
    .D(_00349_),
    .Q_N(_15423_),
    .Q(\mem.mem_internal.code_mem[126][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[126][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1588),
    .D(_00350_),
    .Q_N(_15422_),
    .Q(\mem.mem_internal.code_mem[126][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[126][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1589),
    .D(_00351_),
    .Q_N(_15421_),
    .Q(\mem.mem_internal.code_mem[126][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[126][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1590),
    .D(_00352_),
    .Q_N(_15420_),
    .Q(\mem.mem_internal.code_mem[126][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[126][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1591),
    .D(_00353_),
    .Q_N(_15419_),
    .Q(\mem.mem_internal.code_mem[126][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[127][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1592),
    .D(_00354_),
    .Q_N(_15418_),
    .Q(\mem.mem_internal.code_mem[127][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[127][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1593),
    .D(_00355_),
    .Q_N(_15417_),
    .Q(\mem.mem_internal.code_mem[127][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[127][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1594),
    .D(_00356_),
    .Q_N(_15416_),
    .Q(\mem.mem_internal.code_mem[127][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[127][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1595),
    .D(_00357_),
    .Q_N(_15415_),
    .Q(\mem.mem_internal.code_mem[127][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[127][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1596),
    .D(_00358_),
    .Q_N(_15414_),
    .Q(\mem.mem_internal.code_mem[127][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[127][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1597),
    .D(_00359_),
    .Q_N(_15413_),
    .Q(\mem.mem_internal.code_mem[127][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[127][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1598),
    .D(_00360_),
    .Q_N(_15412_),
    .Q(\mem.mem_internal.code_mem[127][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[127][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1599),
    .D(_00361_),
    .Q_N(_15411_),
    .Q(\mem.mem_internal.code_mem[127][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[128][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1600),
    .D(_00362_),
    .Q_N(_15410_),
    .Q(\mem.mem_internal.code_mem[128][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[128][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1601),
    .D(_00363_),
    .Q_N(_15409_),
    .Q(\mem.mem_internal.code_mem[128][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[128][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1602),
    .D(_00364_),
    .Q_N(_15408_),
    .Q(\mem.mem_internal.code_mem[128][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[128][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1603),
    .D(_00365_),
    .Q_N(_15407_),
    .Q(\mem.mem_internal.code_mem[128][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[128][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1604),
    .D(_00366_),
    .Q_N(_15406_),
    .Q(\mem.mem_internal.code_mem[128][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[128][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1605),
    .D(_00367_),
    .Q_N(_15405_),
    .Q(\mem.mem_internal.code_mem[128][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[128][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1606),
    .D(_00368_),
    .Q_N(_15404_),
    .Q(\mem.mem_internal.code_mem[128][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[128][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1607),
    .D(_00369_),
    .Q_N(_15403_),
    .Q(\mem.mem_internal.code_mem[128][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[129][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1608),
    .D(_00370_),
    .Q_N(_15402_),
    .Q(\mem.mem_internal.code_mem[129][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[129][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1609),
    .D(_00371_),
    .Q_N(_15401_),
    .Q(\mem.mem_internal.code_mem[129][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[129][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1610),
    .D(_00372_),
    .Q_N(_15400_),
    .Q(\mem.mem_internal.code_mem[129][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[129][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1611),
    .D(_00373_),
    .Q_N(_15399_),
    .Q(\mem.mem_internal.code_mem[129][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[129][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1612),
    .D(_00374_),
    .Q_N(_15398_),
    .Q(\mem.mem_internal.code_mem[129][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[129][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1613),
    .D(_00375_),
    .Q_N(_15397_),
    .Q(\mem.mem_internal.code_mem[129][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[129][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1614),
    .D(_00376_),
    .Q_N(_15396_),
    .Q(\mem.mem_internal.code_mem[129][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[129][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1615),
    .D(_00377_),
    .Q_N(_15395_),
    .Q(\mem.mem_internal.code_mem[129][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[12][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1616),
    .D(_00378_),
    .Q_N(_15394_),
    .Q(\mem.mem_internal.code_mem[12][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[12][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1617),
    .D(_00379_),
    .Q_N(_15393_),
    .Q(\mem.mem_internal.code_mem[12][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[12][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1618),
    .D(_00380_),
    .Q_N(_15392_),
    .Q(\mem.mem_internal.code_mem[12][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[12][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1619),
    .D(_00381_),
    .Q_N(_15391_),
    .Q(\mem.mem_internal.code_mem[12][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[12][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1620),
    .D(_00382_),
    .Q_N(_15390_),
    .Q(\mem.mem_internal.code_mem[12][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[12][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1621),
    .D(_00383_),
    .Q_N(_15389_),
    .Q(\mem.mem_internal.code_mem[12][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[12][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1622),
    .D(_00384_),
    .Q_N(_15388_),
    .Q(\mem.mem_internal.code_mem[12][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[12][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1623),
    .D(_00385_),
    .Q_N(_15387_),
    .Q(\mem.mem_internal.code_mem[12][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[130][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1624),
    .D(_00386_),
    .Q_N(_15386_),
    .Q(\mem.mem_internal.code_mem[130][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[130][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1625),
    .D(_00387_),
    .Q_N(_15385_),
    .Q(\mem.mem_internal.code_mem[130][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[130][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1626),
    .D(_00388_),
    .Q_N(_15384_),
    .Q(\mem.mem_internal.code_mem[130][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[130][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1627),
    .D(_00389_),
    .Q_N(_15383_),
    .Q(\mem.mem_internal.code_mem[130][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[130][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1628),
    .D(_00390_),
    .Q_N(_15382_),
    .Q(\mem.mem_internal.code_mem[130][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[130][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1629),
    .D(_00391_),
    .Q_N(_15381_),
    .Q(\mem.mem_internal.code_mem[130][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[130][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1630),
    .D(_00392_),
    .Q_N(_15380_),
    .Q(\mem.mem_internal.code_mem[130][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[130][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1631),
    .D(_00393_),
    .Q_N(_15379_),
    .Q(\mem.mem_internal.code_mem[130][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[131][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1632),
    .D(_00394_),
    .Q_N(_15378_),
    .Q(\mem.mem_internal.code_mem[131][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[131][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1633),
    .D(_00395_),
    .Q_N(_15377_),
    .Q(\mem.mem_internal.code_mem[131][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[131][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1634),
    .D(_00396_),
    .Q_N(_15376_),
    .Q(\mem.mem_internal.code_mem[131][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[131][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1635),
    .D(_00397_),
    .Q_N(_15375_),
    .Q(\mem.mem_internal.code_mem[131][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[131][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1636),
    .D(_00398_),
    .Q_N(_15374_),
    .Q(\mem.mem_internal.code_mem[131][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[131][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1637),
    .D(_00399_),
    .Q_N(_15373_),
    .Q(\mem.mem_internal.code_mem[131][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[131][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1638),
    .D(_00400_),
    .Q_N(_15372_),
    .Q(\mem.mem_internal.code_mem[131][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[131][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1639),
    .D(_00401_),
    .Q_N(_15371_),
    .Q(\mem.mem_internal.code_mem[131][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[132][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1640),
    .D(_00402_),
    .Q_N(_15370_),
    .Q(\mem.mem_internal.code_mem[132][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[132][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1641),
    .D(_00403_),
    .Q_N(_15369_),
    .Q(\mem.mem_internal.code_mem[132][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[132][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1642),
    .D(_00404_),
    .Q_N(_15368_),
    .Q(\mem.mem_internal.code_mem[132][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[132][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1643),
    .D(_00405_),
    .Q_N(_15367_),
    .Q(\mem.mem_internal.code_mem[132][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[132][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1644),
    .D(_00406_),
    .Q_N(_15366_),
    .Q(\mem.mem_internal.code_mem[132][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[132][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1645),
    .D(_00407_),
    .Q_N(_15365_),
    .Q(\mem.mem_internal.code_mem[132][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[132][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1646),
    .D(_00408_),
    .Q_N(_15364_),
    .Q(\mem.mem_internal.code_mem[132][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[132][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1647),
    .D(_00409_),
    .Q_N(_15363_),
    .Q(\mem.mem_internal.code_mem[132][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[133][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1648),
    .D(_00410_),
    .Q_N(_15362_),
    .Q(\mem.mem_internal.code_mem[133][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[133][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1649),
    .D(_00411_),
    .Q_N(_15361_),
    .Q(\mem.mem_internal.code_mem[133][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[133][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1650),
    .D(_00412_),
    .Q_N(_15360_),
    .Q(\mem.mem_internal.code_mem[133][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[133][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1651),
    .D(_00413_),
    .Q_N(_15359_),
    .Q(\mem.mem_internal.code_mem[133][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[133][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1652),
    .D(_00414_),
    .Q_N(_15358_),
    .Q(\mem.mem_internal.code_mem[133][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[133][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1653),
    .D(_00415_),
    .Q_N(_15357_),
    .Q(\mem.mem_internal.code_mem[133][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[133][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1654),
    .D(_00416_),
    .Q_N(_15356_),
    .Q(\mem.mem_internal.code_mem[133][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[133][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1655),
    .D(_00417_),
    .Q_N(_15355_),
    .Q(\mem.mem_internal.code_mem[133][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[134][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1656),
    .D(_00418_),
    .Q_N(_15354_),
    .Q(\mem.mem_internal.code_mem[134][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[134][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1657),
    .D(_00419_),
    .Q_N(_15353_),
    .Q(\mem.mem_internal.code_mem[134][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[134][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1658),
    .D(_00420_),
    .Q_N(_15352_),
    .Q(\mem.mem_internal.code_mem[134][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[134][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1659),
    .D(_00421_),
    .Q_N(_15351_),
    .Q(\mem.mem_internal.code_mem[134][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[134][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1660),
    .D(_00422_),
    .Q_N(_15350_),
    .Q(\mem.mem_internal.code_mem[134][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[134][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1661),
    .D(_00423_),
    .Q_N(_15349_),
    .Q(\mem.mem_internal.code_mem[134][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[134][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1662),
    .D(_00424_),
    .Q_N(_15348_),
    .Q(\mem.mem_internal.code_mem[134][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[134][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1663),
    .D(_00425_),
    .Q_N(_15347_),
    .Q(\mem.mem_internal.code_mem[134][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[135][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1664),
    .D(_00426_),
    .Q_N(_15346_),
    .Q(\mem.mem_internal.code_mem[135][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[135][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1665),
    .D(_00427_),
    .Q_N(_15345_),
    .Q(\mem.mem_internal.code_mem[135][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[135][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1666),
    .D(_00428_),
    .Q_N(_15344_),
    .Q(\mem.mem_internal.code_mem[135][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[135][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1667),
    .D(_00429_),
    .Q_N(_15343_),
    .Q(\mem.mem_internal.code_mem[135][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[135][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1668),
    .D(_00430_),
    .Q_N(_15342_),
    .Q(\mem.mem_internal.code_mem[135][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[135][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1669),
    .D(_00431_),
    .Q_N(_15341_),
    .Q(\mem.mem_internal.code_mem[135][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[135][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1670),
    .D(_00432_),
    .Q_N(_15340_),
    .Q(\mem.mem_internal.code_mem[135][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[135][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1671),
    .D(_00433_),
    .Q_N(_15339_),
    .Q(\mem.mem_internal.code_mem[135][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[136][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1672),
    .D(_00434_),
    .Q_N(_15338_),
    .Q(\mem.mem_internal.code_mem[136][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[136][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1673),
    .D(_00435_),
    .Q_N(_15337_),
    .Q(\mem.mem_internal.code_mem[136][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[136][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1674),
    .D(_00436_),
    .Q_N(_15336_),
    .Q(\mem.mem_internal.code_mem[136][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[136][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1675),
    .D(_00437_),
    .Q_N(_15335_),
    .Q(\mem.mem_internal.code_mem[136][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[136][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1676),
    .D(_00438_),
    .Q_N(_15334_),
    .Q(\mem.mem_internal.code_mem[136][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[136][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1677),
    .D(_00439_),
    .Q_N(_15333_),
    .Q(\mem.mem_internal.code_mem[136][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[136][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1678),
    .D(_00440_),
    .Q_N(_15332_),
    .Q(\mem.mem_internal.code_mem[136][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[136][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1679),
    .D(_00441_),
    .Q_N(_15331_),
    .Q(\mem.mem_internal.code_mem[136][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[137][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1680),
    .D(_00442_),
    .Q_N(_15330_),
    .Q(\mem.mem_internal.code_mem[137][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[137][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1681),
    .D(_00443_),
    .Q_N(_15329_),
    .Q(\mem.mem_internal.code_mem[137][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[137][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1682),
    .D(_00444_),
    .Q_N(_15328_),
    .Q(\mem.mem_internal.code_mem[137][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[137][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1683),
    .D(_00445_),
    .Q_N(_15327_),
    .Q(\mem.mem_internal.code_mem[137][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[137][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1684),
    .D(_00446_),
    .Q_N(_15326_),
    .Q(\mem.mem_internal.code_mem[137][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[137][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1685),
    .D(_00447_),
    .Q_N(_15325_),
    .Q(\mem.mem_internal.code_mem[137][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[137][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1686),
    .D(_00448_),
    .Q_N(_15324_),
    .Q(\mem.mem_internal.code_mem[137][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[137][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1687),
    .D(_00449_),
    .Q_N(_15323_),
    .Q(\mem.mem_internal.code_mem[137][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[138][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1688),
    .D(_00450_),
    .Q_N(_15322_),
    .Q(\mem.mem_internal.code_mem[138][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[138][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1689),
    .D(_00451_),
    .Q_N(_15321_),
    .Q(\mem.mem_internal.code_mem[138][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[138][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1690),
    .D(_00452_),
    .Q_N(_15320_),
    .Q(\mem.mem_internal.code_mem[138][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[138][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1691),
    .D(_00453_),
    .Q_N(_15319_),
    .Q(\mem.mem_internal.code_mem[138][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[138][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1692),
    .D(_00454_),
    .Q_N(_15318_),
    .Q(\mem.mem_internal.code_mem[138][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[138][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1693),
    .D(_00455_),
    .Q_N(_15317_),
    .Q(\mem.mem_internal.code_mem[138][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[138][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1694),
    .D(_00456_),
    .Q_N(_15316_),
    .Q(\mem.mem_internal.code_mem[138][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[138][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1695),
    .D(_00457_),
    .Q_N(_15315_),
    .Q(\mem.mem_internal.code_mem[138][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[139][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1696),
    .D(_00458_),
    .Q_N(_15314_),
    .Q(\mem.mem_internal.code_mem[139][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[139][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1697),
    .D(_00459_),
    .Q_N(_15313_),
    .Q(\mem.mem_internal.code_mem[139][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[139][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1698),
    .D(_00460_),
    .Q_N(_15312_),
    .Q(\mem.mem_internal.code_mem[139][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[139][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1699),
    .D(_00461_),
    .Q_N(_15311_),
    .Q(\mem.mem_internal.code_mem[139][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[139][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1700),
    .D(_00462_),
    .Q_N(_15310_),
    .Q(\mem.mem_internal.code_mem[139][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[139][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1701),
    .D(_00463_),
    .Q_N(_15309_),
    .Q(\mem.mem_internal.code_mem[139][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[139][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1702),
    .D(_00464_),
    .Q_N(_15308_),
    .Q(\mem.mem_internal.code_mem[139][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[139][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1703),
    .D(_00465_),
    .Q_N(_15307_),
    .Q(\mem.mem_internal.code_mem[139][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[13][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1704),
    .D(_00466_),
    .Q_N(_15306_),
    .Q(\mem.mem_internal.code_mem[13][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[13][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1705),
    .D(_00467_),
    .Q_N(_15305_),
    .Q(\mem.mem_internal.code_mem[13][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[13][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1706),
    .D(_00468_),
    .Q_N(_15304_),
    .Q(\mem.mem_internal.code_mem[13][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[13][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1707),
    .D(_00469_),
    .Q_N(_15303_),
    .Q(\mem.mem_internal.code_mem[13][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[13][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1708),
    .D(_00470_),
    .Q_N(_15302_),
    .Q(\mem.mem_internal.code_mem[13][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[13][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1709),
    .D(_00471_),
    .Q_N(_15301_),
    .Q(\mem.mem_internal.code_mem[13][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[13][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1710),
    .D(_00472_),
    .Q_N(_15300_),
    .Q(\mem.mem_internal.code_mem[13][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[13][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1711),
    .D(_00473_),
    .Q_N(_15299_),
    .Q(\mem.mem_internal.code_mem[13][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[140][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1712),
    .D(_00474_),
    .Q_N(_15298_),
    .Q(\mem.mem_internal.code_mem[140][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[140][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1713),
    .D(_00475_),
    .Q_N(_15297_),
    .Q(\mem.mem_internal.code_mem[140][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[140][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1714),
    .D(_00476_),
    .Q_N(_15296_),
    .Q(\mem.mem_internal.code_mem[140][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[140][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1715),
    .D(_00477_),
    .Q_N(_15295_),
    .Q(\mem.mem_internal.code_mem[140][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[140][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1716),
    .D(_00478_),
    .Q_N(_15294_),
    .Q(\mem.mem_internal.code_mem[140][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[140][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1717),
    .D(_00479_),
    .Q_N(_15293_),
    .Q(\mem.mem_internal.code_mem[140][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[140][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1718),
    .D(_00480_),
    .Q_N(_15292_),
    .Q(\mem.mem_internal.code_mem[140][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[140][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1719),
    .D(_00481_),
    .Q_N(_15291_),
    .Q(\mem.mem_internal.code_mem[140][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[141][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1720),
    .D(_00482_),
    .Q_N(_15290_),
    .Q(\mem.mem_internal.code_mem[141][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[141][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1721),
    .D(_00483_),
    .Q_N(_15289_),
    .Q(\mem.mem_internal.code_mem[141][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[141][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1722),
    .D(_00484_),
    .Q_N(_15288_),
    .Q(\mem.mem_internal.code_mem[141][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[141][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1723),
    .D(_00485_),
    .Q_N(_15287_),
    .Q(\mem.mem_internal.code_mem[141][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[141][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1724),
    .D(_00486_),
    .Q_N(_15286_),
    .Q(\mem.mem_internal.code_mem[141][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[141][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1725),
    .D(_00487_),
    .Q_N(_15285_),
    .Q(\mem.mem_internal.code_mem[141][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[141][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1726),
    .D(_00488_),
    .Q_N(_15284_),
    .Q(\mem.mem_internal.code_mem[141][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[141][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1727),
    .D(_00489_),
    .Q_N(_15283_),
    .Q(\mem.mem_internal.code_mem[141][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[142][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1728),
    .D(_00490_),
    .Q_N(_15282_),
    .Q(\mem.mem_internal.code_mem[142][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[142][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1729),
    .D(_00491_),
    .Q_N(_15281_),
    .Q(\mem.mem_internal.code_mem[142][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[142][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1730),
    .D(_00492_),
    .Q_N(_15280_),
    .Q(\mem.mem_internal.code_mem[142][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[142][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1731),
    .D(_00493_),
    .Q_N(_15279_),
    .Q(\mem.mem_internal.code_mem[142][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[142][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1732),
    .D(_00494_),
    .Q_N(_15278_),
    .Q(\mem.mem_internal.code_mem[142][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[142][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1733),
    .D(_00495_),
    .Q_N(_15277_),
    .Q(\mem.mem_internal.code_mem[142][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[142][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1734),
    .D(_00496_),
    .Q_N(_15276_),
    .Q(\mem.mem_internal.code_mem[142][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[142][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1735),
    .D(_00497_),
    .Q_N(_15275_),
    .Q(\mem.mem_internal.code_mem[142][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[143][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1736),
    .D(_00498_),
    .Q_N(_15274_),
    .Q(\mem.mem_internal.code_mem[143][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[143][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1737),
    .D(_00499_),
    .Q_N(_15273_),
    .Q(\mem.mem_internal.code_mem[143][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[143][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1738),
    .D(_00500_),
    .Q_N(_15272_),
    .Q(\mem.mem_internal.code_mem[143][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[143][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1739),
    .D(_00501_),
    .Q_N(_15271_),
    .Q(\mem.mem_internal.code_mem[143][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[143][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1740),
    .D(_00502_),
    .Q_N(_15270_),
    .Q(\mem.mem_internal.code_mem[143][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[143][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1741),
    .D(_00503_),
    .Q_N(_15269_),
    .Q(\mem.mem_internal.code_mem[143][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[143][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1742),
    .D(_00504_),
    .Q_N(_15268_),
    .Q(\mem.mem_internal.code_mem[143][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[143][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1743),
    .D(_00505_),
    .Q_N(_15267_),
    .Q(\mem.mem_internal.code_mem[143][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[144][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1744),
    .D(_00506_),
    .Q_N(_15266_),
    .Q(\mem.mem_internal.code_mem[144][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[144][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1745),
    .D(_00507_),
    .Q_N(_15265_),
    .Q(\mem.mem_internal.code_mem[144][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[144][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1746),
    .D(_00508_),
    .Q_N(_15264_),
    .Q(\mem.mem_internal.code_mem[144][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[144][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1747),
    .D(_00509_),
    .Q_N(_15263_),
    .Q(\mem.mem_internal.code_mem[144][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[144][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1748),
    .D(_00510_),
    .Q_N(_15262_),
    .Q(\mem.mem_internal.code_mem[144][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[144][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1749),
    .D(_00511_),
    .Q_N(_15261_),
    .Q(\mem.mem_internal.code_mem[144][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[144][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1750),
    .D(_00512_),
    .Q_N(_15260_),
    .Q(\mem.mem_internal.code_mem[144][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[144][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1751),
    .D(_00513_),
    .Q_N(_15259_),
    .Q(\mem.mem_internal.code_mem[144][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[145][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1752),
    .D(_00514_),
    .Q_N(_15258_),
    .Q(\mem.mem_internal.code_mem[145][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[145][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1753),
    .D(_00515_),
    .Q_N(_15257_),
    .Q(\mem.mem_internal.code_mem[145][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[145][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1754),
    .D(_00516_),
    .Q_N(_15256_),
    .Q(\mem.mem_internal.code_mem[145][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[145][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1755),
    .D(_00517_),
    .Q_N(_15255_),
    .Q(\mem.mem_internal.code_mem[145][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[145][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1756),
    .D(_00518_),
    .Q_N(_15254_),
    .Q(\mem.mem_internal.code_mem[145][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[145][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1757),
    .D(_00519_),
    .Q_N(_15253_),
    .Q(\mem.mem_internal.code_mem[145][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[145][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1758),
    .D(_00520_),
    .Q_N(_15252_),
    .Q(\mem.mem_internal.code_mem[145][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[145][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1759),
    .D(_00521_),
    .Q_N(_15251_),
    .Q(\mem.mem_internal.code_mem[145][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[146][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1760),
    .D(_00522_),
    .Q_N(_15250_),
    .Q(\mem.mem_internal.code_mem[146][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[146][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1761),
    .D(_00523_),
    .Q_N(_15249_),
    .Q(\mem.mem_internal.code_mem[146][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[146][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1762),
    .D(_00524_),
    .Q_N(_15248_),
    .Q(\mem.mem_internal.code_mem[146][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[146][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1763),
    .D(_00525_),
    .Q_N(_15247_),
    .Q(\mem.mem_internal.code_mem[146][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[146][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1764),
    .D(_00526_),
    .Q_N(_15246_),
    .Q(\mem.mem_internal.code_mem[146][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[146][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1765),
    .D(_00527_),
    .Q_N(_15245_),
    .Q(\mem.mem_internal.code_mem[146][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[146][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1766),
    .D(_00528_),
    .Q_N(_15244_),
    .Q(\mem.mem_internal.code_mem[146][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[146][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1767),
    .D(_00529_),
    .Q_N(_15243_),
    .Q(\mem.mem_internal.code_mem[146][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[147][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1768),
    .D(_00530_),
    .Q_N(_15242_),
    .Q(\mem.mem_internal.code_mem[147][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[147][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1769),
    .D(_00531_),
    .Q_N(_15241_),
    .Q(\mem.mem_internal.code_mem[147][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[147][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1770),
    .D(_00532_),
    .Q_N(_15240_),
    .Q(\mem.mem_internal.code_mem[147][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[147][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1771),
    .D(_00533_),
    .Q_N(_15239_),
    .Q(\mem.mem_internal.code_mem[147][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[147][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1772),
    .D(_00534_),
    .Q_N(_15238_),
    .Q(\mem.mem_internal.code_mem[147][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[147][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1773),
    .D(_00535_),
    .Q_N(_15237_),
    .Q(\mem.mem_internal.code_mem[147][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[147][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1774),
    .D(_00536_),
    .Q_N(_15236_),
    .Q(\mem.mem_internal.code_mem[147][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[147][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1775),
    .D(_00537_),
    .Q_N(_15235_),
    .Q(\mem.mem_internal.code_mem[147][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[148][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1776),
    .D(_00538_),
    .Q_N(_15234_),
    .Q(\mem.mem_internal.code_mem[148][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[148][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1777),
    .D(_00539_),
    .Q_N(_15233_),
    .Q(\mem.mem_internal.code_mem[148][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[148][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1778),
    .D(_00540_),
    .Q_N(_15232_),
    .Q(\mem.mem_internal.code_mem[148][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[148][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1779),
    .D(_00541_),
    .Q_N(_15231_),
    .Q(\mem.mem_internal.code_mem[148][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[148][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1780),
    .D(_00542_),
    .Q_N(_15230_),
    .Q(\mem.mem_internal.code_mem[148][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[148][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1781),
    .D(_00543_),
    .Q_N(_15229_),
    .Q(\mem.mem_internal.code_mem[148][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[148][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1782),
    .D(_00544_),
    .Q_N(_15228_),
    .Q(\mem.mem_internal.code_mem[148][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[148][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1783),
    .D(_00545_),
    .Q_N(_15227_),
    .Q(\mem.mem_internal.code_mem[148][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[149][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1784),
    .D(_00546_),
    .Q_N(_15226_),
    .Q(\mem.mem_internal.code_mem[149][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[149][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1785),
    .D(_00547_),
    .Q_N(_15225_),
    .Q(\mem.mem_internal.code_mem[149][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[149][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1786),
    .D(_00548_),
    .Q_N(_15224_),
    .Q(\mem.mem_internal.code_mem[149][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[149][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1787),
    .D(_00549_),
    .Q_N(_15223_),
    .Q(\mem.mem_internal.code_mem[149][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[149][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1788),
    .D(_00550_),
    .Q_N(_15222_),
    .Q(\mem.mem_internal.code_mem[149][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[149][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1789),
    .D(_00551_),
    .Q_N(_15221_),
    .Q(\mem.mem_internal.code_mem[149][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[149][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1790),
    .D(_00552_),
    .Q_N(_15220_),
    .Q(\mem.mem_internal.code_mem[149][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[149][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1791),
    .D(_00553_),
    .Q_N(_15219_),
    .Q(\mem.mem_internal.code_mem[149][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[14][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1792),
    .D(_00554_),
    .Q_N(_15218_),
    .Q(\mem.mem_internal.code_mem[14][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[14][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1793),
    .D(_00555_),
    .Q_N(_15217_),
    .Q(\mem.mem_internal.code_mem[14][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[14][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1794),
    .D(_00556_),
    .Q_N(_15216_),
    .Q(\mem.mem_internal.code_mem[14][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[14][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1795),
    .D(_00557_),
    .Q_N(_15215_),
    .Q(\mem.mem_internal.code_mem[14][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[14][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1796),
    .D(_00558_),
    .Q_N(_15214_),
    .Q(\mem.mem_internal.code_mem[14][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[14][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1797),
    .D(_00559_),
    .Q_N(_15213_),
    .Q(\mem.mem_internal.code_mem[14][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[14][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1798),
    .D(_00560_),
    .Q_N(_15212_),
    .Q(\mem.mem_internal.code_mem[14][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[14][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1799),
    .D(_00561_),
    .Q_N(_15211_),
    .Q(\mem.mem_internal.code_mem[14][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[150][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1800),
    .D(_00562_),
    .Q_N(_15210_),
    .Q(\mem.mem_internal.code_mem[150][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[150][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1801),
    .D(_00563_),
    .Q_N(_15209_),
    .Q(\mem.mem_internal.code_mem[150][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[150][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1802),
    .D(_00564_),
    .Q_N(_15208_),
    .Q(\mem.mem_internal.code_mem[150][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[150][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1803),
    .D(_00565_),
    .Q_N(_15207_),
    .Q(\mem.mem_internal.code_mem[150][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[150][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1804),
    .D(_00566_),
    .Q_N(_15206_),
    .Q(\mem.mem_internal.code_mem[150][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[150][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1805),
    .D(_00567_),
    .Q_N(_15205_),
    .Q(\mem.mem_internal.code_mem[150][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[150][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1806),
    .D(_00568_),
    .Q_N(_15204_),
    .Q(\mem.mem_internal.code_mem[150][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[150][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1807),
    .D(_00569_),
    .Q_N(_15203_),
    .Q(\mem.mem_internal.code_mem[150][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[151][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1808),
    .D(_00570_),
    .Q_N(_15202_),
    .Q(\mem.mem_internal.code_mem[151][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[151][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1809),
    .D(_00571_),
    .Q_N(_15201_),
    .Q(\mem.mem_internal.code_mem[151][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[151][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1810),
    .D(_00572_),
    .Q_N(_15200_),
    .Q(\mem.mem_internal.code_mem[151][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[151][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1811),
    .D(_00573_),
    .Q_N(_15199_),
    .Q(\mem.mem_internal.code_mem[151][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[151][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1812),
    .D(_00574_),
    .Q_N(_15198_),
    .Q(\mem.mem_internal.code_mem[151][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[151][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1813),
    .D(_00575_),
    .Q_N(_15197_),
    .Q(\mem.mem_internal.code_mem[151][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[151][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1814),
    .D(_00576_),
    .Q_N(_15196_),
    .Q(\mem.mem_internal.code_mem[151][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[151][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1815),
    .D(_00577_),
    .Q_N(_15195_),
    .Q(\mem.mem_internal.code_mem[151][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[152][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1816),
    .D(_00578_),
    .Q_N(_15194_),
    .Q(\mem.mem_internal.code_mem[152][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[152][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1817),
    .D(_00579_),
    .Q_N(_15193_),
    .Q(\mem.mem_internal.code_mem[152][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[152][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1818),
    .D(_00580_),
    .Q_N(_15192_),
    .Q(\mem.mem_internal.code_mem[152][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[152][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1819),
    .D(_00581_),
    .Q_N(_15191_),
    .Q(\mem.mem_internal.code_mem[152][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[152][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1820),
    .D(_00582_),
    .Q_N(_15190_),
    .Q(\mem.mem_internal.code_mem[152][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[152][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1821),
    .D(_00583_),
    .Q_N(_15189_),
    .Q(\mem.mem_internal.code_mem[152][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[152][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1822),
    .D(_00584_),
    .Q_N(_15188_),
    .Q(\mem.mem_internal.code_mem[152][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[152][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1823),
    .D(_00585_),
    .Q_N(_15187_),
    .Q(\mem.mem_internal.code_mem[152][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[153][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1824),
    .D(_00586_),
    .Q_N(_15186_),
    .Q(\mem.mem_internal.code_mem[153][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[153][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1825),
    .D(_00587_),
    .Q_N(_15185_),
    .Q(\mem.mem_internal.code_mem[153][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[153][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1826),
    .D(_00588_),
    .Q_N(_15184_),
    .Q(\mem.mem_internal.code_mem[153][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[153][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1827),
    .D(_00589_),
    .Q_N(_15183_),
    .Q(\mem.mem_internal.code_mem[153][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[153][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1828),
    .D(_00590_),
    .Q_N(_15182_),
    .Q(\mem.mem_internal.code_mem[153][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[153][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1829),
    .D(_00591_),
    .Q_N(_15181_),
    .Q(\mem.mem_internal.code_mem[153][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[153][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1830),
    .D(_00592_),
    .Q_N(_15180_),
    .Q(\mem.mem_internal.code_mem[153][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[153][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1831),
    .D(_00593_),
    .Q_N(_15179_),
    .Q(\mem.mem_internal.code_mem[153][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[154][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1832),
    .D(_00594_),
    .Q_N(_15178_),
    .Q(\mem.mem_internal.code_mem[154][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[154][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1833),
    .D(_00595_),
    .Q_N(_15177_),
    .Q(\mem.mem_internal.code_mem[154][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[154][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1834),
    .D(_00596_),
    .Q_N(_15176_),
    .Q(\mem.mem_internal.code_mem[154][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[154][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1835),
    .D(_00597_),
    .Q_N(_15175_),
    .Q(\mem.mem_internal.code_mem[154][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[154][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1836),
    .D(_00598_),
    .Q_N(_15174_),
    .Q(\mem.mem_internal.code_mem[154][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[154][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1837),
    .D(_00599_),
    .Q_N(_15173_),
    .Q(\mem.mem_internal.code_mem[154][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[154][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1838),
    .D(_00600_),
    .Q_N(_15172_),
    .Q(\mem.mem_internal.code_mem[154][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[154][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1839),
    .D(_00601_),
    .Q_N(_15171_),
    .Q(\mem.mem_internal.code_mem[154][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[155][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1840),
    .D(_00602_),
    .Q_N(_15170_),
    .Q(\mem.mem_internal.code_mem[155][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[155][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1841),
    .D(_00603_),
    .Q_N(_15169_),
    .Q(\mem.mem_internal.code_mem[155][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[155][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1842),
    .D(_00604_),
    .Q_N(_15168_),
    .Q(\mem.mem_internal.code_mem[155][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[155][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1843),
    .D(_00605_),
    .Q_N(_15167_),
    .Q(\mem.mem_internal.code_mem[155][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[155][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1844),
    .D(_00606_),
    .Q_N(_15166_),
    .Q(\mem.mem_internal.code_mem[155][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[155][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1845),
    .D(_00607_),
    .Q_N(_15165_),
    .Q(\mem.mem_internal.code_mem[155][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[155][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1846),
    .D(_00608_),
    .Q_N(_15164_),
    .Q(\mem.mem_internal.code_mem[155][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[155][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1847),
    .D(_00609_),
    .Q_N(_15163_),
    .Q(\mem.mem_internal.code_mem[155][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[156][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1848),
    .D(_00610_),
    .Q_N(_15162_),
    .Q(\mem.mem_internal.code_mem[156][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[156][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1849),
    .D(_00611_),
    .Q_N(_15161_),
    .Q(\mem.mem_internal.code_mem[156][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[156][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1850),
    .D(_00612_),
    .Q_N(_15160_),
    .Q(\mem.mem_internal.code_mem[156][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[156][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1851),
    .D(_00613_),
    .Q_N(_15159_),
    .Q(\mem.mem_internal.code_mem[156][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[156][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1852),
    .D(_00614_),
    .Q_N(_15158_),
    .Q(\mem.mem_internal.code_mem[156][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[156][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1853),
    .D(_00615_),
    .Q_N(_15157_),
    .Q(\mem.mem_internal.code_mem[156][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[156][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1854),
    .D(_00616_),
    .Q_N(_15156_),
    .Q(\mem.mem_internal.code_mem[156][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[156][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1855),
    .D(_00617_),
    .Q_N(_15155_),
    .Q(\mem.mem_internal.code_mem[156][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[157][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1856),
    .D(_00618_),
    .Q_N(_15154_),
    .Q(\mem.mem_internal.code_mem[157][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[157][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1857),
    .D(_00619_),
    .Q_N(_15153_),
    .Q(\mem.mem_internal.code_mem[157][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[157][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1858),
    .D(_00620_),
    .Q_N(_15152_),
    .Q(\mem.mem_internal.code_mem[157][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[157][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1859),
    .D(_00621_),
    .Q_N(_15151_),
    .Q(\mem.mem_internal.code_mem[157][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[157][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1860),
    .D(_00622_),
    .Q_N(_15150_),
    .Q(\mem.mem_internal.code_mem[157][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[157][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1861),
    .D(_00623_),
    .Q_N(_15149_),
    .Q(\mem.mem_internal.code_mem[157][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[157][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1862),
    .D(_00624_),
    .Q_N(_15148_),
    .Q(\mem.mem_internal.code_mem[157][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[157][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1863),
    .D(_00625_),
    .Q_N(_15147_),
    .Q(\mem.mem_internal.code_mem[157][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[158][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1864),
    .D(_00626_),
    .Q_N(_15146_),
    .Q(\mem.mem_internal.code_mem[158][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[158][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1865),
    .D(_00627_),
    .Q_N(_15145_),
    .Q(\mem.mem_internal.code_mem[158][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[158][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1866),
    .D(_00628_),
    .Q_N(_15144_),
    .Q(\mem.mem_internal.code_mem[158][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[158][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1867),
    .D(_00629_),
    .Q_N(_15143_),
    .Q(\mem.mem_internal.code_mem[158][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[158][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1868),
    .D(_00630_),
    .Q_N(_15142_),
    .Q(\mem.mem_internal.code_mem[158][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[158][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1869),
    .D(_00631_),
    .Q_N(_15141_),
    .Q(\mem.mem_internal.code_mem[158][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[158][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1870),
    .D(_00632_),
    .Q_N(_15140_),
    .Q(\mem.mem_internal.code_mem[158][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[158][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1871),
    .D(_00633_),
    .Q_N(_15139_),
    .Q(\mem.mem_internal.code_mem[158][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[159][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1872),
    .D(_00634_),
    .Q_N(_15138_),
    .Q(\mem.mem_internal.code_mem[159][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[159][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1873),
    .D(_00635_),
    .Q_N(_15137_),
    .Q(\mem.mem_internal.code_mem[159][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[159][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1874),
    .D(_00636_),
    .Q_N(_15136_),
    .Q(\mem.mem_internal.code_mem[159][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[159][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1875),
    .D(_00637_),
    .Q_N(_15135_),
    .Q(\mem.mem_internal.code_mem[159][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[159][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1876),
    .D(_00638_),
    .Q_N(_15134_),
    .Q(\mem.mem_internal.code_mem[159][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[159][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1877),
    .D(_00639_),
    .Q_N(_15133_),
    .Q(\mem.mem_internal.code_mem[159][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[159][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1878),
    .D(_00640_),
    .Q_N(_15132_),
    .Q(\mem.mem_internal.code_mem[159][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[159][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1879),
    .D(_00641_),
    .Q_N(_15131_),
    .Q(\mem.mem_internal.code_mem[159][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[15][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1880),
    .D(_00642_),
    .Q_N(_15130_),
    .Q(\mem.mem_internal.code_mem[15][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[15][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1881),
    .D(_00643_),
    .Q_N(_15129_),
    .Q(\mem.mem_internal.code_mem[15][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[15][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1882),
    .D(_00644_),
    .Q_N(_15128_),
    .Q(\mem.mem_internal.code_mem[15][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[15][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1883),
    .D(_00645_),
    .Q_N(_15127_),
    .Q(\mem.mem_internal.code_mem[15][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[15][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1884),
    .D(_00646_),
    .Q_N(_15126_),
    .Q(\mem.mem_internal.code_mem[15][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[15][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1885),
    .D(_00647_),
    .Q_N(_15125_),
    .Q(\mem.mem_internal.code_mem[15][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[15][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1886),
    .D(_00648_),
    .Q_N(_15124_),
    .Q(\mem.mem_internal.code_mem[15][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[15][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1887),
    .D(_00649_),
    .Q_N(_15123_),
    .Q(\mem.mem_internal.code_mem[15][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[160][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1888),
    .D(_00650_),
    .Q_N(_15122_),
    .Q(\mem.mem_internal.code_mem[160][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[160][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1889),
    .D(_00651_),
    .Q_N(_15121_),
    .Q(\mem.mem_internal.code_mem[160][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[160][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1890),
    .D(_00652_),
    .Q_N(_15120_),
    .Q(\mem.mem_internal.code_mem[160][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[160][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1891),
    .D(_00653_),
    .Q_N(_15119_),
    .Q(\mem.mem_internal.code_mem[160][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[160][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1892),
    .D(_00654_),
    .Q_N(_15118_),
    .Q(\mem.mem_internal.code_mem[160][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[160][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1893),
    .D(_00655_),
    .Q_N(_15117_),
    .Q(\mem.mem_internal.code_mem[160][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[160][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net1894),
    .D(_00656_),
    .Q_N(_15116_),
    .Q(\mem.mem_internal.code_mem[160][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[160][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1895),
    .D(_00657_),
    .Q_N(_15115_),
    .Q(\mem.mem_internal.code_mem[160][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[161][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1896),
    .D(_00658_),
    .Q_N(_15114_),
    .Q(\mem.mem_internal.code_mem[161][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[161][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1897),
    .D(_00659_),
    .Q_N(_15113_),
    .Q(\mem.mem_internal.code_mem[161][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[161][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1898),
    .D(_00660_),
    .Q_N(_15112_),
    .Q(\mem.mem_internal.code_mem[161][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[161][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1899),
    .D(_00661_),
    .Q_N(_15111_),
    .Q(\mem.mem_internal.code_mem[161][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[161][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1900),
    .D(_00662_),
    .Q_N(_15110_),
    .Q(\mem.mem_internal.code_mem[161][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[161][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1901),
    .D(_00663_),
    .Q_N(_15109_),
    .Q(\mem.mem_internal.code_mem[161][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[161][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1902),
    .D(_00664_),
    .Q_N(_15108_),
    .Q(\mem.mem_internal.code_mem[161][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[161][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1903),
    .D(_00665_),
    .Q_N(_15107_),
    .Q(\mem.mem_internal.code_mem[161][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[162][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1904),
    .D(_00666_),
    .Q_N(_15106_),
    .Q(\mem.mem_internal.code_mem[162][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[162][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1905),
    .D(_00667_),
    .Q_N(_15105_),
    .Q(\mem.mem_internal.code_mem[162][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[162][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1906),
    .D(_00668_),
    .Q_N(_15104_),
    .Q(\mem.mem_internal.code_mem[162][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[162][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1907),
    .D(_00669_),
    .Q_N(_15103_),
    .Q(\mem.mem_internal.code_mem[162][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[162][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1908),
    .D(_00670_),
    .Q_N(_15102_),
    .Q(\mem.mem_internal.code_mem[162][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[162][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1909),
    .D(_00671_),
    .Q_N(_15101_),
    .Q(\mem.mem_internal.code_mem[162][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[162][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1910),
    .D(_00672_),
    .Q_N(_15100_),
    .Q(\mem.mem_internal.code_mem[162][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[162][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1911),
    .D(_00673_),
    .Q_N(_15099_),
    .Q(\mem.mem_internal.code_mem[162][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[163][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1912),
    .D(_00674_),
    .Q_N(_15098_),
    .Q(\mem.mem_internal.code_mem[163][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[163][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1913),
    .D(_00675_),
    .Q_N(_15097_),
    .Q(\mem.mem_internal.code_mem[163][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[163][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1914),
    .D(_00676_),
    .Q_N(_15096_),
    .Q(\mem.mem_internal.code_mem[163][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[163][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1915),
    .D(_00677_),
    .Q_N(_15095_),
    .Q(\mem.mem_internal.code_mem[163][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[163][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1916),
    .D(_00678_),
    .Q_N(_15094_),
    .Q(\mem.mem_internal.code_mem[163][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[163][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1917),
    .D(_00679_),
    .Q_N(_15093_),
    .Q(\mem.mem_internal.code_mem[163][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[163][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1918),
    .D(_00680_),
    .Q_N(_15092_),
    .Q(\mem.mem_internal.code_mem[163][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[163][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1919),
    .D(_00681_),
    .Q_N(_15091_),
    .Q(\mem.mem_internal.code_mem[163][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[164][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1920),
    .D(_00682_),
    .Q_N(_15090_),
    .Q(\mem.mem_internal.code_mem[164][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[164][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1921),
    .D(_00683_),
    .Q_N(_15089_),
    .Q(\mem.mem_internal.code_mem[164][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[164][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1922),
    .D(_00684_),
    .Q_N(_15088_),
    .Q(\mem.mem_internal.code_mem[164][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[164][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1923),
    .D(_00685_),
    .Q_N(_15087_),
    .Q(\mem.mem_internal.code_mem[164][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[164][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1924),
    .D(_00686_),
    .Q_N(_15086_),
    .Q(\mem.mem_internal.code_mem[164][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[164][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1925),
    .D(_00687_),
    .Q_N(_15085_),
    .Q(\mem.mem_internal.code_mem[164][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[164][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1926),
    .D(_00688_),
    .Q_N(_15084_),
    .Q(\mem.mem_internal.code_mem[164][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[164][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1927),
    .D(_00689_),
    .Q_N(_15083_),
    .Q(\mem.mem_internal.code_mem[164][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[165][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1928),
    .D(_00690_),
    .Q_N(_15082_),
    .Q(\mem.mem_internal.code_mem[165][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[165][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1929),
    .D(_00691_),
    .Q_N(_15081_),
    .Q(\mem.mem_internal.code_mem[165][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[165][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1930),
    .D(_00692_),
    .Q_N(_15080_),
    .Q(\mem.mem_internal.code_mem[165][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[165][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1931),
    .D(_00693_),
    .Q_N(_15079_),
    .Q(\mem.mem_internal.code_mem[165][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[165][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1932),
    .D(_00694_),
    .Q_N(_15078_),
    .Q(\mem.mem_internal.code_mem[165][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[165][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1933),
    .D(_00695_),
    .Q_N(_15077_),
    .Q(\mem.mem_internal.code_mem[165][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[165][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1934),
    .D(_00696_),
    .Q_N(_15076_),
    .Q(\mem.mem_internal.code_mem[165][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[165][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1935),
    .D(_00697_),
    .Q_N(_15075_),
    .Q(\mem.mem_internal.code_mem[165][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[166][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1936),
    .D(_00698_),
    .Q_N(_15074_),
    .Q(\mem.mem_internal.code_mem[166][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[166][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1937),
    .D(_00699_),
    .Q_N(_15073_),
    .Q(\mem.mem_internal.code_mem[166][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[166][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1938),
    .D(_00700_),
    .Q_N(_15072_),
    .Q(\mem.mem_internal.code_mem[166][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[166][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1939),
    .D(_00701_),
    .Q_N(_15071_),
    .Q(\mem.mem_internal.code_mem[166][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[166][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1940),
    .D(_00702_),
    .Q_N(_15070_),
    .Q(\mem.mem_internal.code_mem[166][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[166][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1941),
    .D(_00703_),
    .Q_N(_15069_),
    .Q(\mem.mem_internal.code_mem[166][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[166][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1942),
    .D(_00704_),
    .Q_N(_15068_),
    .Q(\mem.mem_internal.code_mem[166][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[166][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1943),
    .D(_00705_),
    .Q_N(_15067_),
    .Q(\mem.mem_internal.code_mem[166][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[167][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1944),
    .D(_00706_),
    .Q_N(_15066_),
    .Q(\mem.mem_internal.code_mem[167][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[167][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1945),
    .D(_00707_),
    .Q_N(_15065_),
    .Q(\mem.mem_internal.code_mem[167][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[167][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1946),
    .D(_00708_),
    .Q_N(_15064_),
    .Q(\mem.mem_internal.code_mem[167][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[167][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1947),
    .D(_00709_),
    .Q_N(_15063_),
    .Q(\mem.mem_internal.code_mem[167][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[167][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1948),
    .D(_00710_),
    .Q_N(_15062_),
    .Q(\mem.mem_internal.code_mem[167][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[167][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1949),
    .D(_00711_),
    .Q_N(_15061_),
    .Q(\mem.mem_internal.code_mem[167][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[167][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1950),
    .D(_00712_),
    .Q_N(_15060_),
    .Q(\mem.mem_internal.code_mem[167][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[167][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1951),
    .D(_00713_),
    .Q_N(_15059_),
    .Q(\mem.mem_internal.code_mem[167][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[168][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1952),
    .D(_00714_),
    .Q_N(_15058_),
    .Q(\mem.mem_internal.code_mem[168][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[168][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1953),
    .D(_00715_),
    .Q_N(_15057_),
    .Q(\mem.mem_internal.code_mem[168][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[168][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1954),
    .D(_00716_),
    .Q_N(_15056_),
    .Q(\mem.mem_internal.code_mem[168][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[168][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1955),
    .D(_00717_),
    .Q_N(_15055_),
    .Q(\mem.mem_internal.code_mem[168][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[168][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1956),
    .D(_00718_),
    .Q_N(_15054_),
    .Q(\mem.mem_internal.code_mem[168][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[168][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1957),
    .D(_00719_),
    .Q_N(_15053_),
    .Q(\mem.mem_internal.code_mem[168][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[168][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1958),
    .D(_00720_),
    .Q_N(_15052_),
    .Q(\mem.mem_internal.code_mem[168][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[168][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1959),
    .D(_00721_),
    .Q_N(_15051_),
    .Q(\mem.mem_internal.code_mem[168][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[169][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1960),
    .D(_00722_),
    .Q_N(_15050_),
    .Q(\mem.mem_internal.code_mem[169][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[169][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1961),
    .D(_00723_),
    .Q_N(_15049_),
    .Q(\mem.mem_internal.code_mem[169][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[169][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1962),
    .D(_00724_),
    .Q_N(_15048_),
    .Q(\mem.mem_internal.code_mem[169][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[169][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1963),
    .D(_00725_),
    .Q_N(_15047_),
    .Q(\mem.mem_internal.code_mem[169][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[169][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1964),
    .D(_00726_),
    .Q_N(_15046_),
    .Q(\mem.mem_internal.code_mem[169][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[169][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1965),
    .D(_00727_),
    .Q_N(_15045_),
    .Q(\mem.mem_internal.code_mem[169][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[169][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1966),
    .D(_00728_),
    .Q_N(_15044_),
    .Q(\mem.mem_internal.code_mem[169][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[169][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1967),
    .D(_00729_),
    .Q_N(_15043_),
    .Q(\mem.mem_internal.code_mem[169][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[16][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1968),
    .D(_00730_),
    .Q_N(_15042_),
    .Q(\mem.mem_internal.code_mem[16][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[16][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1969),
    .D(_00731_),
    .Q_N(_15041_),
    .Q(\mem.mem_internal.code_mem[16][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[16][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1970),
    .D(_00732_),
    .Q_N(_15040_),
    .Q(\mem.mem_internal.code_mem[16][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[16][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1971),
    .D(_00733_),
    .Q_N(_15039_),
    .Q(\mem.mem_internal.code_mem[16][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[16][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1972),
    .D(_00734_),
    .Q_N(_15038_),
    .Q(\mem.mem_internal.code_mem[16][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[16][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1973),
    .D(_00735_),
    .Q_N(_15037_),
    .Q(\mem.mem_internal.code_mem[16][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[16][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1974),
    .D(_00736_),
    .Q_N(_15036_),
    .Q(\mem.mem_internal.code_mem[16][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[16][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1975),
    .D(_00737_),
    .Q_N(_15035_),
    .Q(\mem.mem_internal.code_mem[16][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[170][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1976),
    .D(_00738_),
    .Q_N(_15034_),
    .Q(\mem.mem_internal.code_mem[170][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[170][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1977),
    .D(_00739_),
    .Q_N(_15033_),
    .Q(\mem.mem_internal.code_mem[170][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[170][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1978),
    .D(_00740_),
    .Q_N(_15032_),
    .Q(\mem.mem_internal.code_mem[170][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[170][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1979),
    .D(_00741_),
    .Q_N(_15031_),
    .Q(\mem.mem_internal.code_mem[170][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[170][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1980),
    .D(_00742_),
    .Q_N(_15030_),
    .Q(\mem.mem_internal.code_mem[170][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[170][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1981),
    .D(_00743_),
    .Q_N(_15029_),
    .Q(\mem.mem_internal.code_mem[170][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[170][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1982),
    .D(_00744_),
    .Q_N(_15028_),
    .Q(\mem.mem_internal.code_mem[170][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[170][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1983),
    .D(_00745_),
    .Q_N(_15027_),
    .Q(\mem.mem_internal.code_mem[170][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[171][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1984),
    .D(_00746_),
    .Q_N(_15026_),
    .Q(\mem.mem_internal.code_mem[171][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[171][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1985),
    .D(_00747_),
    .Q_N(_15025_),
    .Q(\mem.mem_internal.code_mem[171][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[171][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1986),
    .D(_00748_),
    .Q_N(_15024_),
    .Q(\mem.mem_internal.code_mem[171][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[171][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1987),
    .D(_00749_),
    .Q_N(_15023_),
    .Q(\mem.mem_internal.code_mem[171][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[171][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1988),
    .D(_00750_),
    .Q_N(_15022_),
    .Q(\mem.mem_internal.code_mem[171][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[171][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1989),
    .D(_00751_),
    .Q_N(_15021_),
    .Q(\mem.mem_internal.code_mem[171][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[171][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1990),
    .D(_00752_),
    .Q_N(_15020_),
    .Q(\mem.mem_internal.code_mem[171][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[171][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1991),
    .D(_00753_),
    .Q_N(_15019_),
    .Q(\mem.mem_internal.code_mem[171][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[172][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1992),
    .D(_00754_),
    .Q_N(_15018_),
    .Q(\mem.mem_internal.code_mem[172][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[172][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1993),
    .D(_00755_),
    .Q_N(_15017_),
    .Q(\mem.mem_internal.code_mem[172][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[172][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1994),
    .D(_00756_),
    .Q_N(_15016_),
    .Q(\mem.mem_internal.code_mem[172][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[172][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1995),
    .D(_00757_),
    .Q_N(_15015_),
    .Q(\mem.mem_internal.code_mem[172][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[172][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1996),
    .D(_00758_),
    .Q_N(_15014_),
    .Q(\mem.mem_internal.code_mem[172][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[172][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1997),
    .D(_00759_),
    .Q_N(_15013_),
    .Q(\mem.mem_internal.code_mem[172][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[172][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1998),
    .D(_00760_),
    .Q_N(_15012_),
    .Q(\mem.mem_internal.code_mem[172][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[172][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1999),
    .D(_00761_),
    .Q_N(_15011_),
    .Q(\mem.mem_internal.code_mem[172][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[173][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2000),
    .D(_00762_),
    .Q_N(_15010_),
    .Q(\mem.mem_internal.code_mem[173][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[173][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2001),
    .D(_00763_),
    .Q_N(_15009_),
    .Q(\mem.mem_internal.code_mem[173][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[173][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2002),
    .D(_00764_),
    .Q_N(_15008_),
    .Q(\mem.mem_internal.code_mem[173][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[173][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2003),
    .D(_00765_),
    .Q_N(_15007_),
    .Q(\mem.mem_internal.code_mem[173][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[173][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2004),
    .D(_00766_),
    .Q_N(_15006_),
    .Q(\mem.mem_internal.code_mem[173][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[173][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2005),
    .D(_00767_),
    .Q_N(_15005_),
    .Q(\mem.mem_internal.code_mem[173][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[173][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2006),
    .D(_00768_),
    .Q_N(_15004_),
    .Q(\mem.mem_internal.code_mem[173][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[173][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2007),
    .D(_00769_),
    .Q_N(_15003_),
    .Q(\mem.mem_internal.code_mem[173][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[174][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2008),
    .D(_00770_),
    .Q_N(_15002_),
    .Q(\mem.mem_internal.code_mem[174][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[174][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2009),
    .D(_00771_),
    .Q_N(_15001_),
    .Q(\mem.mem_internal.code_mem[174][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[174][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2010),
    .D(_00772_),
    .Q_N(_15000_),
    .Q(\mem.mem_internal.code_mem[174][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[174][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2011),
    .D(_00773_),
    .Q_N(_14999_),
    .Q(\mem.mem_internal.code_mem[174][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[174][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2012),
    .D(_00774_),
    .Q_N(_14998_),
    .Q(\mem.mem_internal.code_mem[174][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[174][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2013),
    .D(_00775_),
    .Q_N(_14997_),
    .Q(\mem.mem_internal.code_mem[174][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[174][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2014),
    .D(_00776_),
    .Q_N(_14996_),
    .Q(\mem.mem_internal.code_mem[174][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[174][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2015),
    .D(_00777_),
    .Q_N(_14995_),
    .Q(\mem.mem_internal.code_mem[174][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[175][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2016),
    .D(_00778_),
    .Q_N(_14994_),
    .Q(\mem.mem_internal.code_mem[175][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[175][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2017),
    .D(_00779_),
    .Q_N(_14993_),
    .Q(\mem.mem_internal.code_mem[175][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[175][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2018),
    .D(_00780_),
    .Q_N(_14992_),
    .Q(\mem.mem_internal.code_mem[175][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[175][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2019),
    .D(_00781_),
    .Q_N(_14991_),
    .Q(\mem.mem_internal.code_mem[175][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[175][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2020),
    .D(_00782_),
    .Q_N(_14990_),
    .Q(\mem.mem_internal.code_mem[175][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[175][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2021),
    .D(_00783_),
    .Q_N(_14989_),
    .Q(\mem.mem_internal.code_mem[175][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[175][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2022),
    .D(_00784_),
    .Q_N(_14988_),
    .Q(\mem.mem_internal.code_mem[175][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[175][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2023),
    .D(_00785_),
    .Q_N(_14987_),
    .Q(\mem.mem_internal.code_mem[175][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[176][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2024),
    .D(_00786_),
    .Q_N(_14986_),
    .Q(\mem.mem_internal.code_mem[176][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[176][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2025),
    .D(_00787_),
    .Q_N(_14985_),
    .Q(\mem.mem_internal.code_mem[176][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[176][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net2026),
    .D(_00788_),
    .Q_N(_14984_),
    .Q(\mem.mem_internal.code_mem[176][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[176][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net2027),
    .D(_00789_),
    .Q_N(_14983_),
    .Q(\mem.mem_internal.code_mem[176][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[176][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net2028),
    .D(_00790_),
    .Q_N(_14982_),
    .Q(\mem.mem_internal.code_mem[176][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[176][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net2029),
    .D(_00791_),
    .Q_N(_14981_),
    .Q(\mem.mem_internal.code_mem[176][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[176][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net2030),
    .D(_00792_),
    .Q_N(_14980_),
    .Q(\mem.mem_internal.code_mem[176][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[176][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net2031),
    .D(_00793_),
    .Q_N(_14979_),
    .Q(\mem.mem_internal.code_mem[176][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[177][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2032),
    .D(_00794_),
    .Q_N(_14978_),
    .Q(\mem.mem_internal.code_mem[177][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[177][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2033),
    .D(_00795_),
    .Q_N(_14977_),
    .Q(\mem.mem_internal.code_mem[177][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[177][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net2034),
    .D(_00796_),
    .Q_N(_14976_),
    .Q(\mem.mem_internal.code_mem[177][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[177][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net2035),
    .D(_00797_),
    .Q_N(_14975_),
    .Q(\mem.mem_internal.code_mem[177][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[177][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net2036),
    .D(_00798_),
    .Q_N(_14974_),
    .Q(\mem.mem_internal.code_mem[177][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[177][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net2037),
    .D(_00799_),
    .Q_N(_14973_),
    .Q(\mem.mem_internal.code_mem[177][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[177][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net2038),
    .D(_00800_),
    .Q_N(_14972_),
    .Q(\mem.mem_internal.code_mem[177][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[177][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net2039),
    .D(_00801_),
    .Q_N(_14971_),
    .Q(\mem.mem_internal.code_mem[177][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[178][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2040),
    .D(_00802_),
    .Q_N(_14970_),
    .Q(\mem.mem_internal.code_mem[178][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[178][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2041),
    .D(_00803_),
    .Q_N(_14969_),
    .Q(\mem.mem_internal.code_mem[178][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[178][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net2042),
    .D(_00804_),
    .Q_N(_14968_),
    .Q(\mem.mem_internal.code_mem[178][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[178][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net2043),
    .D(_00805_),
    .Q_N(_14967_),
    .Q(\mem.mem_internal.code_mem[178][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[178][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net2044),
    .D(_00806_),
    .Q_N(_14966_),
    .Q(\mem.mem_internal.code_mem[178][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[178][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net2045),
    .D(_00807_),
    .Q_N(_14965_),
    .Q(\mem.mem_internal.code_mem[178][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[178][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2046),
    .D(_00808_),
    .Q_N(_14964_),
    .Q(\mem.mem_internal.code_mem[178][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[178][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net2047),
    .D(_00809_),
    .Q_N(_14963_),
    .Q(\mem.mem_internal.code_mem[178][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[179][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2048),
    .D(_00810_),
    .Q_N(_14962_),
    .Q(\mem.mem_internal.code_mem[179][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[179][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2049),
    .D(_00811_),
    .Q_N(_14961_),
    .Q(\mem.mem_internal.code_mem[179][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[179][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net2050),
    .D(_00812_),
    .Q_N(_14960_),
    .Q(\mem.mem_internal.code_mem[179][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[179][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net2051),
    .D(_00813_),
    .Q_N(_14959_),
    .Q(\mem.mem_internal.code_mem[179][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[179][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net2052),
    .D(_00814_),
    .Q_N(_14958_),
    .Q(\mem.mem_internal.code_mem[179][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[179][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net2053),
    .D(_00815_),
    .Q_N(_14957_),
    .Q(\mem.mem_internal.code_mem[179][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[179][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net2054),
    .D(_00816_),
    .Q_N(_14956_),
    .Q(\mem.mem_internal.code_mem[179][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[179][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net2055),
    .D(_00817_),
    .Q_N(_14955_),
    .Q(\mem.mem_internal.code_mem[179][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[17][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2056),
    .D(_00818_),
    .Q_N(_14954_),
    .Q(\mem.mem_internal.code_mem[17][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[17][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2057),
    .D(_00819_),
    .Q_N(_14953_),
    .Q(\mem.mem_internal.code_mem[17][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[17][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2058),
    .D(_00820_),
    .Q_N(_14952_),
    .Q(\mem.mem_internal.code_mem[17][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[17][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2059),
    .D(_00821_),
    .Q_N(_14951_),
    .Q(\mem.mem_internal.code_mem[17][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[17][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2060),
    .D(_00822_),
    .Q_N(_14950_),
    .Q(\mem.mem_internal.code_mem[17][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[17][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2061),
    .D(_00823_),
    .Q_N(_14949_),
    .Q(\mem.mem_internal.code_mem[17][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[17][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2062),
    .D(_00824_),
    .Q_N(_14948_),
    .Q(\mem.mem_internal.code_mem[17][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[17][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2063),
    .D(_00825_),
    .Q_N(_14947_),
    .Q(\mem.mem_internal.code_mem[17][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[180][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2064),
    .D(_00826_),
    .Q_N(_14946_),
    .Q(\mem.mem_internal.code_mem[180][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[180][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2065),
    .D(_00827_),
    .Q_N(_14945_),
    .Q(\mem.mem_internal.code_mem[180][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[180][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net2066),
    .D(_00828_),
    .Q_N(_14944_),
    .Q(\mem.mem_internal.code_mem[180][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[180][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2067),
    .D(_00829_),
    .Q_N(_14943_),
    .Q(\mem.mem_internal.code_mem[180][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[180][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net2068),
    .D(_00830_),
    .Q_N(_14942_),
    .Q(\mem.mem_internal.code_mem[180][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[180][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2069),
    .D(_00831_),
    .Q_N(_14941_),
    .Q(\mem.mem_internal.code_mem[180][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[180][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2070),
    .D(_00832_),
    .Q_N(_14940_),
    .Q(\mem.mem_internal.code_mem[180][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[180][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net2071),
    .D(_00833_),
    .Q_N(_14939_),
    .Q(\mem.mem_internal.code_mem[180][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[181][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2072),
    .D(_00834_),
    .Q_N(_14938_),
    .Q(\mem.mem_internal.code_mem[181][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[181][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2073),
    .D(_00835_),
    .Q_N(_14937_),
    .Q(\mem.mem_internal.code_mem[181][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[181][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net2074),
    .D(_00836_),
    .Q_N(_14936_),
    .Q(\mem.mem_internal.code_mem[181][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[181][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2075),
    .D(_00837_),
    .Q_N(_14935_),
    .Q(\mem.mem_internal.code_mem[181][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[181][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net2076),
    .D(_00838_),
    .Q_N(_14934_),
    .Q(\mem.mem_internal.code_mem[181][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[181][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2077),
    .D(_00839_),
    .Q_N(_14933_),
    .Q(\mem.mem_internal.code_mem[181][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[181][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2078),
    .D(_00840_),
    .Q_N(_14932_),
    .Q(\mem.mem_internal.code_mem[181][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[181][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2079),
    .D(_00841_),
    .Q_N(_14931_),
    .Q(\mem.mem_internal.code_mem[181][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[182][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2080),
    .D(_00842_),
    .Q_N(_14930_),
    .Q(\mem.mem_internal.code_mem[182][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[182][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2081),
    .D(_00843_),
    .Q_N(_14929_),
    .Q(\mem.mem_internal.code_mem[182][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[182][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net2082),
    .D(_00844_),
    .Q_N(_14928_),
    .Q(\mem.mem_internal.code_mem[182][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[182][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2083),
    .D(_00845_),
    .Q_N(_14927_),
    .Q(\mem.mem_internal.code_mem[182][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[182][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2084),
    .D(_00846_),
    .Q_N(_14926_),
    .Q(\mem.mem_internal.code_mem[182][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[182][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2085),
    .D(_00847_),
    .Q_N(_14925_),
    .Q(\mem.mem_internal.code_mem[182][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[182][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2086),
    .D(_00848_),
    .Q_N(_14924_),
    .Q(\mem.mem_internal.code_mem[182][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[182][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net2087),
    .D(_00849_),
    .Q_N(_14923_),
    .Q(\mem.mem_internal.code_mem[182][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[183][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2088),
    .D(_00850_),
    .Q_N(_14922_),
    .Q(\mem.mem_internal.code_mem[183][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[183][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2089),
    .D(_00851_),
    .Q_N(_14921_),
    .Q(\mem.mem_internal.code_mem[183][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[183][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net2090),
    .D(_00852_),
    .Q_N(_14920_),
    .Q(\mem.mem_internal.code_mem[183][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[183][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2091),
    .D(_00853_),
    .Q_N(_14919_),
    .Q(\mem.mem_internal.code_mem[183][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[183][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2092),
    .D(_00854_),
    .Q_N(_14918_),
    .Q(\mem.mem_internal.code_mem[183][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[183][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2093),
    .D(_00855_),
    .Q_N(_14917_),
    .Q(\mem.mem_internal.code_mem[183][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[183][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2094),
    .D(_00856_),
    .Q_N(_14916_),
    .Q(\mem.mem_internal.code_mem[183][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[183][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2095),
    .D(_00857_),
    .Q_N(_14915_),
    .Q(\mem.mem_internal.code_mem[183][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[184][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2096),
    .D(_00858_),
    .Q_N(_14914_),
    .Q(\mem.mem_internal.code_mem[184][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[184][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2097),
    .D(_00859_),
    .Q_N(_14913_),
    .Q(\mem.mem_internal.code_mem[184][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[184][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2098),
    .D(_00860_),
    .Q_N(_14912_),
    .Q(\mem.mem_internal.code_mem[184][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[184][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2099),
    .D(_00861_),
    .Q_N(_14911_),
    .Q(\mem.mem_internal.code_mem[184][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[184][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2100),
    .D(_00862_),
    .Q_N(_14910_),
    .Q(\mem.mem_internal.code_mem[184][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[184][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2101),
    .D(_00863_),
    .Q_N(_14909_),
    .Q(\mem.mem_internal.code_mem[184][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[184][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2102),
    .D(_00864_),
    .Q_N(_14908_),
    .Q(\mem.mem_internal.code_mem[184][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[184][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2103),
    .D(_00865_),
    .Q_N(_14907_),
    .Q(\mem.mem_internal.code_mem[184][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[185][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2104),
    .D(_00866_),
    .Q_N(_14906_),
    .Q(\mem.mem_internal.code_mem[185][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[185][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2105),
    .D(_00867_),
    .Q_N(_14905_),
    .Q(\mem.mem_internal.code_mem[185][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[185][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2106),
    .D(_00868_),
    .Q_N(_14904_),
    .Q(\mem.mem_internal.code_mem[185][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[185][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2107),
    .D(_00869_),
    .Q_N(_14903_),
    .Q(\mem.mem_internal.code_mem[185][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[185][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2108),
    .D(_00870_),
    .Q_N(_14902_),
    .Q(\mem.mem_internal.code_mem[185][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[185][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2109),
    .D(_00871_),
    .Q_N(_14901_),
    .Q(\mem.mem_internal.code_mem[185][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[185][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2110),
    .D(_00872_),
    .Q_N(_14900_),
    .Q(\mem.mem_internal.code_mem[185][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[185][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2111),
    .D(_00873_),
    .Q_N(_14899_),
    .Q(\mem.mem_internal.code_mem[185][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[186][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2112),
    .D(_00874_),
    .Q_N(_14898_),
    .Q(\mem.mem_internal.code_mem[186][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[186][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2113),
    .D(_00875_),
    .Q_N(_14897_),
    .Q(\mem.mem_internal.code_mem[186][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[186][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2114),
    .D(_00876_),
    .Q_N(_14896_),
    .Q(\mem.mem_internal.code_mem[186][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[186][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2115),
    .D(_00877_),
    .Q_N(_14895_),
    .Q(\mem.mem_internal.code_mem[186][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[186][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2116),
    .D(_00878_),
    .Q_N(_14894_),
    .Q(\mem.mem_internal.code_mem[186][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[186][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2117),
    .D(_00879_),
    .Q_N(_14893_),
    .Q(\mem.mem_internal.code_mem[186][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[186][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2118),
    .D(_00880_),
    .Q_N(_14892_),
    .Q(\mem.mem_internal.code_mem[186][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[186][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2119),
    .D(_00881_),
    .Q_N(_14891_),
    .Q(\mem.mem_internal.code_mem[186][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[187][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2120),
    .D(_00882_),
    .Q_N(_14890_),
    .Q(\mem.mem_internal.code_mem[187][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[187][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2121),
    .D(_00883_),
    .Q_N(_14889_),
    .Q(\mem.mem_internal.code_mem[187][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[187][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2122),
    .D(_00884_),
    .Q_N(_14888_),
    .Q(\mem.mem_internal.code_mem[187][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[187][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2123),
    .D(_00885_),
    .Q_N(_14887_),
    .Q(\mem.mem_internal.code_mem[187][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[187][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2124),
    .D(_00886_),
    .Q_N(_14886_),
    .Q(\mem.mem_internal.code_mem[187][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[187][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2125),
    .D(_00887_),
    .Q_N(_14885_),
    .Q(\mem.mem_internal.code_mem[187][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[187][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2126),
    .D(_00888_),
    .Q_N(_14884_),
    .Q(\mem.mem_internal.code_mem[187][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[187][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2127),
    .D(_00889_),
    .Q_N(_14883_),
    .Q(\mem.mem_internal.code_mem[187][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[188][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2128),
    .D(_00890_),
    .Q_N(_14882_),
    .Q(\mem.mem_internal.code_mem[188][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[188][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2129),
    .D(_00891_),
    .Q_N(_14881_),
    .Q(\mem.mem_internal.code_mem[188][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[188][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2130),
    .D(_00892_),
    .Q_N(_14880_),
    .Q(\mem.mem_internal.code_mem[188][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[188][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2131),
    .D(_00893_),
    .Q_N(_14879_),
    .Q(\mem.mem_internal.code_mem[188][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[188][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2132),
    .D(_00894_),
    .Q_N(_14878_),
    .Q(\mem.mem_internal.code_mem[188][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[188][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2133),
    .D(_00895_),
    .Q_N(_14877_),
    .Q(\mem.mem_internal.code_mem[188][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[188][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2134),
    .D(_00896_),
    .Q_N(_14876_),
    .Q(\mem.mem_internal.code_mem[188][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[188][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2135),
    .D(_00897_),
    .Q_N(_14875_),
    .Q(\mem.mem_internal.code_mem[188][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[189][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2136),
    .D(_00898_),
    .Q_N(_14874_),
    .Q(\mem.mem_internal.code_mem[189][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[189][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2137),
    .D(_00899_),
    .Q_N(_14873_),
    .Q(\mem.mem_internal.code_mem[189][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[189][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2138),
    .D(_00900_),
    .Q_N(_14872_),
    .Q(\mem.mem_internal.code_mem[189][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[189][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2139),
    .D(_00901_),
    .Q_N(_14871_),
    .Q(\mem.mem_internal.code_mem[189][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[189][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2140),
    .D(_00902_),
    .Q_N(_14870_),
    .Q(\mem.mem_internal.code_mem[189][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[189][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2141),
    .D(_00903_),
    .Q_N(_14869_),
    .Q(\mem.mem_internal.code_mem[189][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[189][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2142),
    .D(_00904_),
    .Q_N(_14868_),
    .Q(\mem.mem_internal.code_mem[189][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[189][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2143),
    .D(_00905_),
    .Q_N(_14867_),
    .Q(\mem.mem_internal.code_mem[189][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[18][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2144),
    .D(_00906_),
    .Q_N(_14866_),
    .Q(\mem.mem_internal.code_mem[18][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[18][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2145),
    .D(_00907_),
    .Q_N(_14865_),
    .Q(\mem.mem_internal.code_mem[18][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[18][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2146),
    .D(_00908_),
    .Q_N(_14864_),
    .Q(\mem.mem_internal.code_mem[18][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[18][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2147),
    .D(_00909_),
    .Q_N(_14863_),
    .Q(\mem.mem_internal.code_mem[18][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[18][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2148),
    .D(_00910_),
    .Q_N(_14862_),
    .Q(\mem.mem_internal.code_mem[18][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[18][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2149),
    .D(_00911_),
    .Q_N(_14861_),
    .Q(\mem.mem_internal.code_mem[18][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[18][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2150),
    .D(_00912_),
    .Q_N(_14860_),
    .Q(\mem.mem_internal.code_mem[18][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[18][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2151),
    .D(_00913_),
    .Q_N(_14859_),
    .Q(\mem.mem_internal.code_mem[18][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[190][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2152),
    .D(_00914_),
    .Q_N(_14858_),
    .Q(\mem.mem_internal.code_mem[190][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[190][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2153),
    .D(_00915_),
    .Q_N(_14857_),
    .Q(\mem.mem_internal.code_mem[190][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[190][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2154),
    .D(_00916_),
    .Q_N(_14856_),
    .Q(\mem.mem_internal.code_mem[190][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[190][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2155),
    .D(_00917_),
    .Q_N(_14855_),
    .Q(\mem.mem_internal.code_mem[190][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[190][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2156),
    .D(_00918_),
    .Q_N(_14854_),
    .Q(\mem.mem_internal.code_mem[190][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[190][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2157),
    .D(_00919_),
    .Q_N(_14853_),
    .Q(\mem.mem_internal.code_mem[190][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[190][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2158),
    .D(_00920_),
    .Q_N(_14852_),
    .Q(\mem.mem_internal.code_mem[190][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[190][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2159),
    .D(_00921_),
    .Q_N(_14851_),
    .Q(\mem.mem_internal.code_mem[190][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[191][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2160),
    .D(_00922_),
    .Q_N(_14850_),
    .Q(\mem.mem_internal.code_mem[191][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[191][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2161),
    .D(_00923_),
    .Q_N(_14849_),
    .Q(\mem.mem_internal.code_mem[191][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[191][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2162),
    .D(_00924_),
    .Q_N(_14848_),
    .Q(\mem.mem_internal.code_mem[191][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[191][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2163),
    .D(_00925_),
    .Q_N(_14847_),
    .Q(\mem.mem_internal.code_mem[191][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[191][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2164),
    .D(_00926_),
    .Q_N(_14846_),
    .Q(\mem.mem_internal.code_mem[191][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[191][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2165),
    .D(_00927_),
    .Q_N(_14845_),
    .Q(\mem.mem_internal.code_mem[191][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[191][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2166),
    .D(_00928_),
    .Q_N(_14844_),
    .Q(\mem.mem_internal.code_mem[191][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[191][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2167),
    .D(_00929_),
    .Q_N(_14843_),
    .Q(\mem.mem_internal.code_mem[191][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[192][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2168),
    .D(_00930_),
    .Q_N(_14842_),
    .Q(\mem.mem_internal.code_mem[192][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[192][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2169),
    .D(_00931_),
    .Q_N(_14841_),
    .Q(\mem.mem_internal.code_mem[192][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[192][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2170),
    .D(_00932_),
    .Q_N(_14840_),
    .Q(\mem.mem_internal.code_mem[192][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[192][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2171),
    .D(_00933_),
    .Q_N(_14839_),
    .Q(\mem.mem_internal.code_mem[192][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[192][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2172),
    .D(_00934_),
    .Q_N(_14838_),
    .Q(\mem.mem_internal.code_mem[192][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[192][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2173),
    .D(_00935_),
    .Q_N(_14837_),
    .Q(\mem.mem_internal.code_mem[192][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[192][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2174),
    .D(_00936_),
    .Q_N(_14836_),
    .Q(\mem.mem_internal.code_mem[192][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[192][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2175),
    .D(_00937_),
    .Q_N(_14835_),
    .Q(\mem.mem_internal.code_mem[192][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[193][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2176),
    .D(_00938_),
    .Q_N(_14834_),
    .Q(\mem.mem_internal.code_mem[193][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[193][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2177),
    .D(_00939_),
    .Q_N(_14833_),
    .Q(\mem.mem_internal.code_mem[193][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[193][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2178),
    .D(_00940_),
    .Q_N(_14832_),
    .Q(\mem.mem_internal.code_mem[193][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[193][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2179),
    .D(_00941_),
    .Q_N(_14831_),
    .Q(\mem.mem_internal.code_mem[193][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[193][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2180),
    .D(_00942_),
    .Q_N(_14830_),
    .Q(\mem.mem_internal.code_mem[193][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[193][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2181),
    .D(_00943_),
    .Q_N(_14829_),
    .Q(\mem.mem_internal.code_mem[193][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[193][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2182),
    .D(_00944_),
    .Q_N(_14828_),
    .Q(\mem.mem_internal.code_mem[193][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[193][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2183),
    .D(_00945_),
    .Q_N(_14827_),
    .Q(\mem.mem_internal.code_mem[193][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[194][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2184),
    .D(_00946_),
    .Q_N(_14826_),
    .Q(\mem.mem_internal.code_mem[194][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[194][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2185),
    .D(_00947_),
    .Q_N(_14825_),
    .Q(\mem.mem_internal.code_mem[194][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[194][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2186),
    .D(_00948_),
    .Q_N(_14824_),
    .Q(\mem.mem_internal.code_mem[194][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[194][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2187),
    .D(_00949_),
    .Q_N(_14823_),
    .Q(\mem.mem_internal.code_mem[194][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[194][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2188),
    .D(_00950_),
    .Q_N(_14822_),
    .Q(\mem.mem_internal.code_mem[194][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[194][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2189),
    .D(_00951_),
    .Q_N(_14821_),
    .Q(\mem.mem_internal.code_mem[194][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[194][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2190),
    .D(_00952_),
    .Q_N(_14820_),
    .Q(\mem.mem_internal.code_mem[194][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[194][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2191),
    .D(_00953_),
    .Q_N(_14819_),
    .Q(\mem.mem_internal.code_mem[194][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[195][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2192),
    .D(_00954_),
    .Q_N(_14818_),
    .Q(\mem.mem_internal.code_mem[195][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[195][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2193),
    .D(_00955_),
    .Q_N(_14817_),
    .Q(\mem.mem_internal.code_mem[195][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[195][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2194),
    .D(_00956_),
    .Q_N(_14816_),
    .Q(\mem.mem_internal.code_mem[195][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[195][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2195),
    .D(_00957_),
    .Q_N(_14815_),
    .Q(\mem.mem_internal.code_mem[195][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[195][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2196),
    .D(_00958_),
    .Q_N(_14814_),
    .Q(\mem.mem_internal.code_mem[195][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[195][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2197),
    .D(_00959_),
    .Q_N(_14813_),
    .Q(\mem.mem_internal.code_mem[195][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[195][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2198),
    .D(_00960_),
    .Q_N(_14812_),
    .Q(\mem.mem_internal.code_mem[195][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[195][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2199),
    .D(_00961_),
    .Q_N(_14811_),
    .Q(\mem.mem_internal.code_mem[195][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[196][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2200),
    .D(_00962_),
    .Q_N(_14810_),
    .Q(\mem.mem_internal.code_mem[196][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[196][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2201),
    .D(_00963_),
    .Q_N(_14809_),
    .Q(\mem.mem_internal.code_mem[196][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[196][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2202),
    .D(_00964_),
    .Q_N(_14808_),
    .Q(\mem.mem_internal.code_mem[196][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[196][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2203),
    .D(_00965_),
    .Q_N(_14807_),
    .Q(\mem.mem_internal.code_mem[196][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[196][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2204),
    .D(_00966_),
    .Q_N(_14806_),
    .Q(\mem.mem_internal.code_mem[196][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[196][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2205),
    .D(_00967_),
    .Q_N(_14805_),
    .Q(\mem.mem_internal.code_mem[196][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[196][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2206),
    .D(_00968_),
    .Q_N(_14804_),
    .Q(\mem.mem_internal.code_mem[196][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[196][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2207),
    .D(_00969_),
    .Q_N(_14803_),
    .Q(\mem.mem_internal.code_mem[196][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[197][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2208),
    .D(_00970_),
    .Q_N(_14802_),
    .Q(\mem.mem_internal.code_mem[197][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[197][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2209),
    .D(_00971_),
    .Q_N(_14801_),
    .Q(\mem.mem_internal.code_mem[197][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[197][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2210),
    .D(_00972_),
    .Q_N(_14800_),
    .Q(\mem.mem_internal.code_mem[197][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[197][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2211),
    .D(_00973_),
    .Q_N(_14799_),
    .Q(\mem.mem_internal.code_mem[197][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[197][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2212),
    .D(_00974_),
    .Q_N(_14798_),
    .Q(\mem.mem_internal.code_mem[197][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[197][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2213),
    .D(_00975_),
    .Q_N(_14797_),
    .Q(\mem.mem_internal.code_mem[197][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[197][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2214),
    .D(_00976_),
    .Q_N(_14796_),
    .Q(\mem.mem_internal.code_mem[197][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[197][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2215),
    .D(_00977_),
    .Q_N(_14795_),
    .Q(\mem.mem_internal.code_mem[197][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[198][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2216),
    .D(_00978_),
    .Q_N(_14794_),
    .Q(\mem.mem_internal.code_mem[198][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[198][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2217),
    .D(_00979_),
    .Q_N(_14793_),
    .Q(\mem.mem_internal.code_mem[198][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[198][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2218),
    .D(_00980_),
    .Q_N(_14792_),
    .Q(\mem.mem_internal.code_mem[198][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[198][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2219),
    .D(_00981_),
    .Q_N(_14791_),
    .Q(\mem.mem_internal.code_mem[198][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[198][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2220),
    .D(_00982_),
    .Q_N(_14790_),
    .Q(\mem.mem_internal.code_mem[198][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[198][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2221),
    .D(_00983_),
    .Q_N(_14789_),
    .Q(\mem.mem_internal.code_mem[198][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[198][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2222),
    .D(_00984_),
    .Q_N(_14788_),
    .Q(\mem.mem_internal.code_mem[198][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[198][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2223),
    .D(_00985_),
    .Q_N(_14787_),
    .Q(\mem.mem_internal.code_mem[198][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[199][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2224),
    .D(_00986_),
    .Q_N(_14786_),
    .Q(\mem.mem_internal.code_mem[199][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[199][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2225),
    .D(_00987_),
    .Q_N(_14785_),
    .Q(\mem.mem_internal.code_mem[199][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[199][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2226),
    .D(_00988_),
    .Q_N(_14784_),
    .Q(\mem.mem_internal.code_mem[199][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[199][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2227),
    .D(_00989_),
    .Q_N(_14783_),
    .Q(\mem.mem_internal.code_mem[199][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[199][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2228),
    .D(_00990_),
    .Q_N(_14782_),
    .Q(\mem.mem_internal.code_mem[199][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[199][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2229),
    .D(_00991_),
    .Q_N(_14781_),
    .Q(\mem.mem_internal.code_mem[199][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[199][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2230),
    .D(_00992_),
    .Q_N(_14780_),
    .Q(\mem.mem_internal.code_mem[199][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[199][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2231),
    .D(_00993_),
    .Q_N(_14779_),
    .Q(\mem.mem_internal.code_mem[199][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[19][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2232),
    .D(_00994_),
    .Q_N(_14778_),
    .Q(\mem.mem_internal.code_mem[19][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[19][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2233),
    .D(_00995_),
    .Q_N(_14777_),
    .Q(\mem.mem_internal.code_mem[19][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[19][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2234),
    .D(_00996_),
    .Q_N(_14776_),
    .Q(\mem.mem_internal.code_mem[19][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[19][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2235),
    .D(_00997_),
    .Q_N(_14775_),
    .Q(\mem.mem_internal.code_mem[19][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[19][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2236),
    .D(_00998_),
    .Q_N(_14774_),
    .Q(\mem.mem_internal.code_mem[19][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[19][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2237),
    .D(_00999_),
    .Q_N(_14773_),
    .Q(\mem.mem_internal.code_mem[19][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[19][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2238),
    .D(_01000_),
    .Q_N(_14772_),
    .Q(\mem.mem_internal.code_mem[19][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[19][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2239),
    .D(_01001_),
    .Q_N(_14771_),
    .Q(\mem.mem_internal.code_mem[19][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2240),
    .D(_01002_),
    .Q_N(_14770_),
    .Q(\mem.mem_internal.code_mem[1][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2241),
    .D(_01003_),
    .Q_N(_14769_),
    .Q(\mem.mem_internal.code_mem[1][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[1][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2242),
    .D(_01004_),
    .Q_N(_14768_),
    .Q(\mem.mem_internal.code_mem[1][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2243),
    .D(_01005_),
    .Q_N(_14767_),
    .Q(\mem.mem_internal.code_mem[1][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[1][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2244),
    .D(_01006_),
    .Q_N(_14766_),
    .Q(\mem.mem_internal.code_mem[1][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[1][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2245),
    .D(_01007_),
    .Q_N(_14765_),
    .Q(\mem.mem_internal.code_mem[1][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[1][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2246),
    .D(_01008_),
    .Q_N(_14764_),
    .Q(\mem.mem_internal.code_mem[1][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[1][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2247),
    .D(_01009_),
    .Q_N(_14763_),
    .Q(\mem.mem_internal.code_mem[1][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[200][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2248),
    .D(_01010_),
    .Q_N(_14762_),
    .Q(\mem.mem_internal.code_mem[200][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[200][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2249),
    .D(_01011_),
    .Q_N(_14761_),
    .Q(\mem.mem_internal.code_mem[200][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[200][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2250),
    .D(_01012_),
    .Q_N(_14760_),
    .Q(\mem.mem_internal.code_mem[200][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[200][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2251),
    .D(_01013_),
    .Q_N(_14759_),
    .Q(\mem.mem_internal.code_mem[200][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[200][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2252),
    .D(_01014_),
    .Q_N(_14758_),
    .Q(\mem.mem_internal.code_mem[200][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[200][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2253),
    .D(_01015_),
    .Q_N(_14757_),
    .Q(\mem.mem_internal.code_mem[200][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[200][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2254),
    .D(_01016_),
    .Q_N(_14756_),
    .Q(\mem.mem_internal.code_mem[200][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[200][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2255),
    .D(_01017_),
    .Q_N(_14755_),
    .Q(\mem.mem_internal.code_mem[200][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[201][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2256),
    .D(_01018_),
    .Q_N(_14754_),
    .Q(\mem.mem_internal.code_mem[201][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[201][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2257),
    .D(_01019_),
    .Q_N(_14753_),
    .Q(\mem.mem_internal.code_mem[201][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[201][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2258),
    .D(_01020_),
    .Q_N(_14752_),
    .Q(\mem.mem_internal.code_mem[201][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[201][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2259),
    .D(_01021_),
    .Q_N(_14751_),
    .Q(\mem.mem_internal.code_mem[201][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[201][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2260),
    .D(_01022_),
    .Q_N(_14750_),
    .Q(\mem.mem_internal.code_mem[201][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[201][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2261),
    .D(_01023_),
    .Q_N(_14749_),
    .Q(\mem.mem_internal.code_mem[201][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[201][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2262),
    .D(_01024_),
    .Q_N(_14748_),
    .Q(\mem.mem_internal.code_mem[201][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[201][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2263),
    .D(_01025_),
    .Q_N(_14747_),
    .Q(\mem.mem_internal.code_mem[201][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[202][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2264),
    .D(_01026_),
    .Q_N(_14746_),
    .Q(\mem.mem_internal.code_mem[202][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[202][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2265),
    .D(_01027_),
    .Q_N(_14745_),
    .Q(\mem.mem_internal.code_mem[202][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[202][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2266),
    .D(_01028_),
    .Q_N(_14744_),
    .Q(\mem.mem_internal.code_mem[202][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[202][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2267),
    .D(_01029_),
    .Q_N(_14743_),
    .Q(\mem.mem_internal.code_mem[202][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[202][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2268),
    .D(_01030_),
    .Q_N(_14742_),
    .Q(\mem.mem_internal.code_mem[202][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[202][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2269),
    .D(_01031_),
    .Q_N(_14741_),
    .Q(\mem.mem_internal.code_mem[202][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[202][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2270),
    .D(_01032_),
    .Q_N(_14740_),
    .Q(\mem.mem_internal.code_mem[202][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[202][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2271),
    .D(_01033_),
    .Q_N(_14739_),
    .Q(\mem.mem_internal.code_mem[202][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[203][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2272),
    .D(_01034_),
    .Q_N(_14738_),
    .Q(\mem.mem_internal.code_mem[203][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[203][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2273),
    .D(_01035_),
    .Q_N(_14737_),
    .Q(\mem.mem_internal.code_mem[203][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[203][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2274),
    .D(_01036_),
    .Q_N(_14736_),
    .Q(\mem.mem_internal.code_mem[203][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[203][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2275),
    .D(_01037_),
    .Q_N(_14735_),
    .Q(\mem.mem_internal.code_mem[203][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[203][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2276),
    .D(_01038_),
    .Q_N(_14734_),
    .Q(\mem.mem_internal.code_mem[203][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[203][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2277),
    .D(_01039_),
    .Q_N(_14733_),
    .Q(\mem.mem_internal.code_mem[203][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[203][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2278),
    .D(_01040_),
    .Q_N(_14732_),
    .Q(\mem.mem_internal.code_mem[203][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[203][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2279),
    .D(_01041_),
    .Q_N(_14731_),
    .Q(\mem.mem_internal.code_mem[203][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[204][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2280),
    .D(_01042_),
    .Q_N(_14730_),
    .Q(\mem.mem_internal.code_mem[204][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[204][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2281),
    .D(_01043_),
    .Q_N(_14729_),
    .Q(\mem.mem_internal.code_mem[204][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[204][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2282),
    .D(_01044_),
    .Q_N(_14728_),
    .Q(\mem.mem_internal.code_mem[204][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[204][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2283),
    .D(_01045_),
    .Q_N(_14727_),
    .Q(\mem.mem_internal.code_mem[204][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[204][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2284),
    .D(_01046_),
    .Q_N(_14726_),
    .Q(\mem.mem_internal.code_mem[204][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[204][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2285),
    .D(_01047_),
    .Q_N(_14725_),
    .Q(\mem.mem_internal.code_mem[204][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[204][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2286),
    .D(_01048_),
    .Q_N(_14724_),
    .Q(\mem.mem_internal.code_mem[204][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[204][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2287),
    .D(_01049_),
    .Q_N(_14723_),
    .Q(\mem.mem_internal.code_mem[204][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[205][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2288),
    .D(_01050_),
    .Q_N(_14722_),
    .Q(\mem.mem_internal.code_mem[205][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[205][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2289),
    .D(_01051_),
    .Q_N(_14721_),
    .Q(\mem.mem_internal.code_mem[205][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[205][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2290),
    .D(_01052_),
    .Q_N(_14720_),
    .Q(\mem.mem_internal.code_mem[205][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[205][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2291),
    .D(_01053_),
    .Q_N(_14719_),
    .Q(\mem.mem_internal.code_mem[205][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[205][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2292),
    .D(_01054_),
    .Q_N(_14718_),
    .Q(\mem.mem_internal.code_mem[205][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[205][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2293),
    .D(_01055_),
    .Q_N(_14717_),
    .Q(\mem.mem_internal.code_mem[205][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[205][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2294),
    .D(_01056_),
    .Q_N(_14716_),
    .Q(\mem.mem_internal.code_mem[205][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[205][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2295),
    .D(_01057_),
    .Q_N(_14715_),
    .Q(\mem.mem_internal.code_mem[205][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[206][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2296),
    .D(_01058_),
    .Q_N(_14714_),
    .Q(\mem.mem_internal.code_mem[206][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[206][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2297),
    .D(_01059_),
    .Q_N(_14713_),
    .Q(\mem.mem_internal.code_mem[206][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[206][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2298),
    .D(_01060_),
    .Q_N(_14712_),
    .Q(\mem.mem_internal.code_mem[206][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[206][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2299),
    .D(_01061_),
    .Q_N(_14711_),
    .Q(\mem.mem_internal.code_mem[206][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[206][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2300),
    .D(_01062_),
    .Q_N(_14710_),
    .Q(\mem.mem_internal.code_mem[206][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[206][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2301),
    .D(_01063_),
    .Q_N(_14709_),
    .Q(\mem.mem_internal.code_mem[206][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[206][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2302),
    .D(_01064_),
    .Q_N(_14708_),
    .Q(\mem.mem_internal.code_mem[206][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[206][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2303),
    .D(_01065_),
    .Q_N(_14707_),
    .Q(\mem.mem_internal.code_mem[206][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[207][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2304),
    .D(_01066_),
    .Q_N(_14706_),
    .Q(\mem.mem_internal.code_mem[207][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[207][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2305),
    .D(_01067_),
    .Q_N(_14705_),
    .Q(\mem.mem_internal.code_mem[207][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[207][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2306),
    .D(_01068_),
    .Q_N(_14704_),
    .Q(\mem.mem_internal.code_mem[207][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[207][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2307),
    .D(_01069_),
    .Q_N(_14703_),
    .Q(\mem.mem_internal.code_mem[207][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[207][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2308),
    .D(_01070_),
    .Q_N(_14702_),
    .Q(\mem.mem_internal.code_mem[207][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[207][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2309),
    .D(_01071_),
    .Q_N(_14701_),
    .Q(\mem.mem_internal.code_mem[207][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[207][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2310),
    .D(_01072_),
    .Q_N(_14700_),
    .Q(\mem.mem_internal.code_mem[207][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[207][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2311),
    .D(_01073_),
    .Q_N(_14699_),
    .Q(\mem.mem_internal.code_mem[207][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[208][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2312),
    .D(_01074_),
    .Q_N(_14698_),
    .Q(\mem.mem_internal.code_mem[208][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[208][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2313),
    .D(_01075_),
    .Q_N(_14697_),
    .Q(\mem.mem_internal.code_mem[208][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[208][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2314),
    .D(_01076_),
    .Q_N(_14696_),
    .Q(\mem.mem_internal.code_mem[208][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[208][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2315),
    .D(_01077_),
    .Q_N(_14695_),
    .Q(\mem.mem_internal.code_mem[208][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[208][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2316),
    .D(_01078_),
    .Q_N(_14694_),
    .Q(\mem.mem_internal.code_mem[208][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[208][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2317),
    .D(_01079_),
    .Q_N(_14693_),
    .Q(\mem.mem_internal.code_mem[208][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[208][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2318),
    .D(_01080_),
    .Q_N(_14692_),
    .Q(\mem.mem_internal.code_mem[208][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[208][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2319),
    .D(_01081_),
    .Q_N(_14691_),
    .Q(\mem.mem_internal.code_mem[208][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[209][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2320),
    .D(_01082_),
    .Q_N(_14690_),
    .Q(\mem.mem_internal.code_mem[209][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[209][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2321),
    .D(_01083_),
    .Q_N(_14689_),
    .Q(\mem.mem_internal.code_mem[209][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[209][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2322),
    .D(_01084_),
    .Q_N(_14688_),
    .Q(\mem.mem_internal.code_mem[209][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[209][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2323),
    .D(_01085_),
    .Q_N(_14687_),
    .Q(\mem.mem_internal.code_mem[209][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[209][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2324),
    .D(_01086_),
    .Q_N(_14686_),
    .Q(\mem.mem_internal.code_mem[209][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[209][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2325),
    .D(_01087_),
    .Q_N(_14685_),
    .Q(\mem.mem_internal.code_mem[209][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[209][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2326),
    .D(_01088_),
    .Q_N(_14684_),
    .Q(\mem.mem_internal.code_mem[209][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[209][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2327),
    .D(_01089_),
    .Q_N(_14683_),
    .Q(\mem.mem_internal.code_mem[209][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[20][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2328),
    .D(_01090_),
    .Q_N(_14682_),
    .Q(\mem.mem_internal.code_mem[20][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[20][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2329),
    .D(_01091_),
    .Q_N(_14681_),
    .Q(\mem.mem_internal.code_mem[20][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[20][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2330),
    .D(_01092_),
    .Q_N(_14680_),
    .Q(\mem.mem_internal.code_mem[20][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[20][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2331),
    .D(_01093_),
    .Q_N(_14679_),
    .Q(\mem.mem_internal.code_mem[20][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[20][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2332),
    .D(_01094_),
    .Q_N(_14678_),
    .Q(\mem.mem_internal.code_mem[20][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[20][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2333),
    .D(_01095_),
    .Q_N(_14677_),
    .Q(\mem.mem_internal.code_mem[20][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[20][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2334),
    .D(_01096_),
    .Q_N(_14676_),
    .Q(\mem.mem_internal.code_mem[20][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[20][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2335),
    .D(_01097_),
    .Q_N(_14675_),
    .Q(\mem.mem_internal.code_mem[20][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[210][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2336),
    .D(_01098_),
    .Q_N(_14674_),
    .Q(\mem.mem_internal.code_mem[210][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[210][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2337),
    .D(_01099_),
    .Q_N(_14673_),
    .Q(\mem.mem_internal.code_mem[210][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[210][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2338),
    .D(_01100_),
    .Q_N(_14672_),
    .Q(\mem.mem_internal.code_mem[210][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[210][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2339),
    .D(_01101_),
    .Q_N(_14671_),
    .Q(\mem.mem_internal.code_mem[210][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[210][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2340),
    .D(_01102_),
    .Q_N(_14670_),
    .Q(\mem.mem_internal.code_mem[210][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[210][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2341),
    .D(_01103_),
    .Q_N(_14669_),
    .Q(\mem.mem_internal.code_mem[210][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[210][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2342),
    .D(_01104_),
    .Q_N(_14668_),
    .Q(\mem.mem_internal.code_mem[210][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[210][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2343),
    .D(_01105_),
    .Q_N(_14667_),
    .Q(\mem.mem_internal.code_mem[210][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[211][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2344),
    .D(_01106_),
    .Q_N(_14666_),
    .Q(\mem.mem_internal.code_mem[211][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[211][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2345),
    .D(_01107_),
    .Q_N(_14665_),
    .Q(\mem.mem_internal.code_mem[211][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[211][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2346),
    .D(_01108_),
    .Q_N(_14664_),
    .Q(\mem.mem_internal.code_mem[211][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[211][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2347),
    .D(_01109_),
    .Q_N(_14663_),
    .Q(\mem.mem_internal.code_mem[211][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[211][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2348),
    .D(_01110_),
    .Q_N(_14662_),
    .Q(\mem.mem_internal.code_mem[211][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[211][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2349),
    .D(_01111_),
    .Q_N(_14661_),
    .Q(\mem.mem_internal.code_mem[211][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[211][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2350),
    .D(_01112_),
    .Q_N(_14660_),
    .Q(\mem.mem_internal.code_mem[211][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[211][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2351),
    .D(_01113_),
    .Q_N(_14659_),
    .Q(\mem.mem_internal.code_mem[211][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[212][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2352),
    .D(_01114_),
    .Q_N(_14658_),
    .Q(\mem.mem_internal.code_mem[212][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[212][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2353),
    .D(_01115_),
    .Q_N(_14657_),
    .Q(\mem.mem_internal.code_mem[212][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[212][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2354),
    .D(_01116_),
    .Q_N(_14656_),
    .Q(\mem.mem_internal.code_mem[212][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[212][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2355),
    .D(_01117_),
    .Q_N(_14655_),
    .Q(\mem.mem_internal.code_mem[212][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[212][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2356),
    .D(_01118_),
    .Q_N(_14654_),
    .Q(\mem.mem_internal.code_mem[212][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[212][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2357),
    .D(_01119_),
    .Q_N(_14653_),
    .Q(\mem.mem_internal.code_mem[212][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[212][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2358),
    .D(_01120_),
    .Q_N(_14652_),
    .Q(\mem.mem_internal.code_mem[212][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[212][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2359),
    .D(_01121_),
    .Q_N(_14651_),
    .Q(\mem.mem_internal.code_mem[212][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[213][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2360),
    .D(_01122_),
    .Q_N(_14650_),
    .Q(\mem.mem_internal.code_mem[213][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[213][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2361),
    .D(_01123_),
    .Q_N(_14649_),
    .Q(\mem.mem_internal.code_mem[213][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[213][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2362),
    .D(_01124_),
    .Q_N(_14648_),
    .Q(\mem.mem_internal.code_mem[213][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[213][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2363),
    .D(_01125_),
    .Q_N(_14647_),
    .Q(\mem.mem_internal.code_mem[213][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[213][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2364),
    .D(_01126_),
    .Q_N(_14646_),
    .Q(\mem.mem_internal.code_mem[213][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[213][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2365),
    .D(_01127_),
    .Q_N(_14645_),
    .Q(\mem.mem_internal.code_mem[213][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[213][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2366),
    .D(_01128_),
    .Q_N(_14644_),
    .Q(\mem.mem_internal.code_mem[213][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[213][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2367),
    .D(_01129_),
    .Q_N(_14643_),
    .Q(\mem.mem_internal.code_mem[213][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[214][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2368),
    .D(_01130_),
    .Q_N(_14642_),
    .Q(\mem.mem_internal.code_mem[214][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[214][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2369),
    .D(_01131_),
    .Q_N(_14641_),
    .Q(\mem.mem_internal.code_mem[214][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[214][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2370),
    .D(_01132_),
    .Q_N(_14640_),
    .Q(\mem.mem_internal.code_mem[214][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[214][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2371),
    .D(_01133_),
    .Q_N(_14639_),
    .Q(\mem.mem_internal.code_mem[214][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[214][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2372),
    .D(_01134_),
    .Q_N(_14638_),
    .Q(\mem.mem_internal.code_mem[214][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[214][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2373),
    .D(_01135_),
    .Q_N(_14637_),
    .Q(\mem.mem_internal.code_mem[214][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[214][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2374),
    .D(_01136_),
    .Q_N(_14636_),
    .Q(\mem.mem_internal.code_mem[214][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[214][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2375),
    .D(_01137_),
    .Q_N(_14635_),
    .Q(\mem.mem_internal.code_mem[214][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[215][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2376),
    .D(_01138_),
    .Q_N(_14634_),
    .Q(\mem.mem_internal.code_mem[215][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[215][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2377),
    .D(_01139_),
    .Q_N(_14633_),
    .Q(\mem.mem_internal.code_mem[215][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[215][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2378),
    .D(_01140_),
    .Q_N(_14632_),
    .Q(\mem.mem_internal.code_mem[215][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[215][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2379),
    .D(_01141_),
    .Q_N(_14631_),
    .Q(\mem.mem_internal.code_mem[215][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[215][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2380),
    .D(_01142_),
    .Q_N(_14630_),
    .Q(\mem.mem_internal.code_mem[215][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[215][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2381),
    .D(_01143_),
    .Q_N(_14629_),
    .Q(\mem.mem_internal.code_mem[215][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[215][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2382),
    .D(_01144_),
    .Q_N(_14628_),
    .Q(\mem.mem_internal.code_mem[215][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[215][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2383),
    .D(_01145_),
    .Q_N(_14627_),
    .Q(\mem.mem_internal.code_mem[215][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[216][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2384),
    .D(_01146_),
    .Q_N(_14626_),
    .Q(\mem.mem_internal.code_mem[216][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[216][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2385),
    .D(_01147_),
    .Q_N(_14625_),
    .Q(\mem.mem_internal.code_mem[216][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[216][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2386),
    .D(_01148_),
    .Q_N(_14624_),
    .Q(\mem.mem_internal.code_mem[216][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[216][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2387),
    .D(_01149_),
    .Q_N(_14623_),
    .Q(\mem.mem_internal.code_mem[216][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[216][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2388),
    .D(_01150_),
    .Q_N(_14622_),
    .Q(\mem.mem_internal.code_mem[216][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[216][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2389),
    .D(_01151_),
    .Q_N(_14621_),
    .Q(\mem.mem_internal.code_mem[216][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[216][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2390),
    .D(_01152_),
    .Q_N(_14620_),
    .Q(\mem.mem_internal.code_mem[216][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[216][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2391),
    .D(_01153_),
    .Q_N(_14619_),
    .Q(\mem.mem_internal.code_mem[216][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[217][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2392),
    .D(_01154_),
    .Q_N(_14618_),
    .Q(\mem.mem_internal.code_mem[217][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[217][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2393),
    .D(_01155_),
    .Q_N(_14617_),
    .Q(\mem.mem_internal.code_mem[217][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[217][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2394),
    .D(_01156_),
    .Q_N(_14616_),
    .Q(\mem.mem_internal.code_mem[217][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[217][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2395),
    .D(_01157_),
    .Q_N(_14615_),
    .Q(\mem.mem_internal.code_mem[217][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[217][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2396),
    .D(_01158_),
    .Q_N(_14614_),
    .Q(\mem.mem_internal.code_mem[217][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[217][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2397),
    .D(_01159_),
    .Q_N(_14613_),
    .Q(\mem.mem_internal.code_mem[217][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[217][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2398),
    .D(_01160_),
    .Q_N(_14612_),
    .Q(\mem.mem_internal.code_mem[217][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[217][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2399),
    .D(_01161_),
    .Q_N(_14611_),
    .Q(\mem.mem_internal.code_mem[217][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[218][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2400),
    .D(_01162_),
    .Q_N(_14610_),
    .Q(\mem.mem_internal.code_mem[218][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[218][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2401),
    .D(_01163_),
    .Q_N(_14609_),
    .Q(\mem.mem_internal.code_mem[218][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[218][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2402),
    .D(_01164_),
    .Q_N(_14608_),
    .Q(\mem.mem_internal.code_mem[218][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[218][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2403),
    .D(_01165_),
    .Q_N(_14607_),
    .Q(\mem.mem_internal.code_mem[218][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[218][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2404),
    .D(_01166_),
    .Q_N(_14606_),
    .Q(\mem.mem_internal.code_mem[218][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[218][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2405),
    .D(_01167_),
    .Q_N(_14605_),
    .Q(\mem.mem_internal.code_mem[218][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[218][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2406),
    .D(_01168_),
    .Q_N(_14604_),
    .Q(\mem.mem_internal.code_mem[218][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[218][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2407),
    .D(_01169_),
    .Q_N(_14603_),
    .Q(\mem.mem_internal.code_mem[218][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[219][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2408),
    .D(_01170_),
    .Q_N(_14602_),
    .Q(\mem.mem_internal.code_mem[219][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[219][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2409),
    .D(_01171_),
    .Q_N(_14601_),
    .Q(\mem.mem_internal.code_mem[219][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[219][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2410),
    .D(_01172_),
    .Q_N(_14600_),
    .Q(\mem.mem_internal.code_mem[219][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[219][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2411),
    .D(_01173_),
    .Q_N(_14599_),
    .Q(\mem.mem_internal.code_mem[219][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[219][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2412),
    .D(_01174_),
    .Q_N(_14598_),
    .Q(\mem.mem_internal.code_mem[219][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[219][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2413),
    .D(_01175_),
    .Q_N(_14597_),
    .Q(\mem.mem_internal.code_mem[219][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[219][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2414),
    .D(_01176_),
    .Q_N(_14596_),
    .Q(\mem.mem_internal.code_mem[219][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[219][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2415),
    .D(_01177_),
    .Q_N(_14595_),
    .Q(\mem.mem_internal.code_mem[219][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[21][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2416),
    .D(_01178_),
    .Q_N(_14594_),
    .Q(\mem.mem_internal.code_mem[21][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[21][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2417),
    .D(_01179_),
    .Q_N(_14593_),
    .Q(\mem.mem_internal.code_mem[21][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[21][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2418),
    .D(_01180_),
    .Q_N(_14592_),
    .Q(\mem.mem_internal.code_mem[21][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[21][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2419),
    .D(_01181_),
    .Q_N(_14591_),
    .Q(\mem.mem_internal.code_mem[21][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[21][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2420),
    .D(_01182_),
    .Q_N(_14590_),
    .Q(\mem.mem_internal.code_mem[21][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[21][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2421),
    .D(_01183_),
    .Q_N(_14589_),
    .Q(\mem.mem_internal.code_mem[21][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[21][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2422),
    .D(_01184_),
    .Q_N(_14588_),
    .Q(\mem.mem_internal.code_mem[21][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[21][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2423),
    .D(_01185_),
    .Q_N(_14587_),
    .Q(\mem.mem_internal.code_mem[21][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[220][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2424),
    .D(_01186_),
    .Q_N(_14586_),
    .Q(\mem.mem_internal.code_mem[220][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[220][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2425),
    .D(_01187_),
    .Q_N(_14585_),
    .Q(\mem.mem_internal.code_mem[220][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[220][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2426),
    .D(_01188_),
    .Q_N(_14584_),
    .Q(\mem.mem_internal.code_mem[220][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[220][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2427),
    .D(_01189_),
    .Q_N(_14583_),
    .Q(\mem.mem_internal.code_mem[220][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[220][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2428),
    .D(_01190_),
    .Q_N(_14582_),
    .Q(\mem.mem_internal.code_mem[220][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[220][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2429),
    .D(_01191_),
    .Q_N(_14581_),
    .Q(\mem.mem_internal.code_mem[220][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[220][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2430),
    .D(_01192_),
    .Q_N(_14580_),
    .Q(\mem.mem_internal.code_mem[220][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[220][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2431),
    .D(_01193_),
    .Q_N(_14579_),
    .Q(\mem.mem_internal.code_mem[220][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[221][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2432),
    .D(_01194_),
    .Q_N(_14578_),
    .Q(\mem.mem_internal.code_mem[221][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[221][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2433),
    .D(_01195_),
    .Q_N(_14577_),
    .Q(\mem.mem_internal.code_mem[221][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[221][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2434),
    .D(_01196_),
    .Q_N(_14576_),
    .Q(\mem.mem_internal.code_mem[221][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[221][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2435),
    .D(_01197_),
    .Q_N(_14575_),
    .Q(\mem.mem_internal.code_mem[221][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[221][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2436),
    .D(_01198_),
    .Q_N(_14574_),
    .Q(\mem.mem_internal.code_mem[221][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[221][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2437),
    .D(_01199_),
    .Q_N(_14573_),
    .Q(\mem.mem_internal.code_mem[221][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[221][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2438),
    .D(_01200_),
    .Q_N(_14572_),
    .Q(\mem.mem_internal.code_mem[221][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[221][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2439),
    .D(_01201_),
    .Q_N(_14571_),
    .Q(\mem.mem_internal.code_mem[221][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[222][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2440),
    .D(_01202_),
    .Q_N(_14570_),
    .Q(\mem.mem_internal.code_mem[222][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[222][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2441),
    .D(_01203_),
    .Q_N(_14569_),
    .Q(\mem.mem_internal.code_mem[222][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[222][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2442),
    .D(_01204_),
    .Q_N(_14568_),
    .Q(\mem.mem_internal.code_mem[222][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[222][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2443),
    .D(_01205_),
    .Q_N(_14567_),
    .Q(\mem.mem_internal.code_mem[222][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[222][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2444),
    .D(_01206_),
    .Q_N(_14566_),
    .Q(\mem.mem_internal.code_mem[222][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[222][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2445),
    .D(_01207_),
    .Q_N(_14565_),
    .Q(\mem.mem_internal.code_mem[222][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[222][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2446),
    .D(_01208_),
    .Q_N(_14564_),
    .Q(\mem.mem_internal.code_mem[222][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[222][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2447),
    .D(_01209_),
    .Q_N(_14563_),
    .Q(\mem.mem_internal.code_mem[222][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[223][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2448),
    .D(_01210_),
    .Q_N(_14562_),
    .Q(\mem.mem_internal.code_mem[223][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[223][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2449),
    .D(_01211_),
    .Q_N(_14561_),
    .Q(\mem.mem_internal.code_mem[223][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[223][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2450),
    .D(_01212_),
    .Q_N(_14560_),
    .Q(\mem.mem_internal.code_mem[223][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[223][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2451),
    .D(_01213_),
    .Q_N(_14559_),
    .Q(\mem.mem_internal.code_mem[223][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[223][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2452),
    .D(_01214_),
    .Q_N(_14558_),
    .Q(\mem.mem_internal.code_mem[223][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[223][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2453),
    .D(_01215_),
    .Q_N(_14557_),
    .Q(\mem.mem_internal.code_mem[223][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[223][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2454),
    .D(_01216_),
    .Q_N(_14556_),
    .Q(\mem.mem_internal.code_mem[223][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[223][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2455),
    .D(_01217_),
    .Q_N(_14555_),
    .Q(\mem.mem_internal.code_mem[223][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[224][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2456),
    .D(_01218_),
    .Q_N(_14554_),
    .Q(\mem.mem_internal.code_mem[224][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[224][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2457),
    .D(_01219_),
    .Q_N(_14553_),
    .Q(\mem.mem_internal.code_mem[224][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[224][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2458),
    .D(_01220_),
    .Q_N(_14552_),
    .Q(\mem.mem_internal.code_mem[224][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[224][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2459),
    .D(_01221_),
    .Q_N(_14551_),
    .Q(\mem.mem_internal.code_mem[224][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[224][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2460),
    .D(_01222_),
    .Q_N(_14550_),
    .Q(\mem.mem_internal.code_mem[224][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[224][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2461),
    .D(_01223_),
    .Q_N(_14549_),
    .Q(\mem.mem_internal.code_mem[224][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[224][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2462),
    .D(_01224_),
    .Q_N(_14548_),
    .Q(\mem.mem_internal.code_mem[224][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[224][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2463),
    .D(_01225_),
    .Q_N(_14547_),
    .Q(\mem.mem_internal.code_mem[224][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[225][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2464),
    .D(_01226_),
    .Q_N(_14546_),
    .Q(\mem.mem_internal.code_mem[225][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[225][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2465),
    .D(_01227_),
    .Q_N(_14545_),
    .Q(\mem.mem_internal.code_mem[225][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[225][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2466),
    .D(_01228_),
    .Q_N(_14544_),
    .Q(\mem.mem_internal.code_mem[225][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[225][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2467),
    .D(_01229_),
    .Q_N(_14543_),
    .Q(\mem.mem_internal.code_mem[225][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[225][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2468),
    .D(_01230_),
    .Q_N(_14542_),
    .Q(\mem.mem_internal.code_mem[225][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[225][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2469),
    .D(_01231_),
    .Q_N(_14541_),
    .Q(\mem.mem_internal.code_mem[225][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[225][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2470),
    .D(_01232_),
    .Q_N(_14540_),
    .Q(\mem.mem_internal.code_mem[225][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[225][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2471),
    .D(_01233_),
    .Q_N(_14539_),
    .Q(\mem.mem_internal.code_mem[225][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[226][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2472),
    .D(_01234_),
    .Q_N(_14538_),
    .Q(\mem.mem_internal.code_mem[226][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[226][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2473),
    .D(_01235_),
    .Q_N(_14537_),
    .Q(\mem.mem_internal.code_mem[226][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[226][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2474),
    .D(_01236_),
    .Q_N(_14536_),
    .Q(\mem.mem_internal.code_mem[226][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[226][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2475),
    .D(_01237_),
    .Q_N(_14535_),
    .Q(\mem.mem_internal.code_mem[226][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[226][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2476),
    .D(_01238_),
    .Q_N(_14534_),
    .Q(\mem.mem_internal.code_mem[226][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[226][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2477),
    .D(_01239_),
    .Q_N(_14533_),
    .Q(\mem.mem_internal.code_mem[226][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[226][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2478),
    .D(_01240_),
    .Q_N(_14532_),
    .Q(\mem.mem_internal.code_mem[226][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[226][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2479),
    .D(_01241_),
    .Q_N(_14531_),
    .Q(\mem.mem_internal.code_mem[226][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[227][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2480),
    .D(_01242_),
    .Q_N(_14530_),
    .Q(\mem.mem_internal.code_mem[227][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[227][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2481),
    .D(_01243_),
    .Q_N(_14529_),
    .Q(\mem.mem_internal.code_mem[227][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[227][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2482),
    .D(_01244_),
    .Q_N(_14528_),
    .Q(\mem.mem_internal.code_mem[227][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[227][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2483),
    .D(_01245_),
    .Q_N(_14527_),
    .Q(\mem.mem_internal.code_mem[227][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[227][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2484),
    .D(_01246_),
    .Q_N(_14526_),
    .Q(\mem.mem_internal.code_mem[227][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[227][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2485),
    .D(_01247_),
    .Q_N(_14525_),
    .Q(\mem.mem_internal.code_mem[227][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[227][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2486),
    .D(_01248_),
    .Q_N(_14524_),
    .Q(\mem.mem_internal.code_mem[227][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[227][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2487),
    .D(_01249_),
    .Q_N(_14523_),
    .Q(\mem.mem_internal.code_mem[227][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[228][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2488),
    .D(_01250_),
    .Q_N(_14522_),
    .Q(\mem.mem_internal.code_mem[228][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[228][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2489),
    .D(_01251_),
    .Q_N(_14521_),
    .Q(\mem.mem_internal.code_mem[228][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[228][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2490),
    .D(_01252_),
    .Q_N(_14520_),
    .Q(\mem.mem_internal.code_mem[228][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[228][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2491),
    .D(_01253_),
    .Q_N(_14519_),
    .Q(\mem.mem_internal.code_mem[228][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[228][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2492),
    .D(_01254_),
    .Q_N(_14518_),
    .Q(\mem.mem_internal.code_mem[228][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[228][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2493),
    .D(_01255_),
    .Q_N(_14517_),
    .Q(\mem.mem_internal.code_mem[228][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[228][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2494),
    .D(_01256_),
    .Q_N(_14516_),
    .Q(\mem.mem_internal.code_mem[228][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[228][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2495),
    .D(_01257_),
    .Q_N(_14515_),
    .Q(\mem.mem_internal.code_mem[228][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[229][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2496),
    .D(_01258_),
    .Q_N(_14514_),
    .Q(\mem.mem_internal.code_mem[229][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[229][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2497),
    .D(_01259_),
    .Q_N(_14513_),
    .Q(\mem.mem_internal.code_mem[229][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[229][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2498),
    .D(_01260_),
    .Q_N(_14512_),
    .Q(\mem.mem_internal.code_mem[229][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[229][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2499),
    .D(_01261_),
    .Q_N(_14511_),
    .Q(\mem.mem_internal.code_mem[229][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[229][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2500),
    .D(_01262_),
    .Q_N(_14510_),
    .Q(\mem.mem_internal.code_mem[229][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[229][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2501),
    .D(_01263_),
    .Q_N(_14509_),
    .Q(\mem.mem_internal.code_mem[229][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[229][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2502),
    .D(_01264_),
    .Q_N(_14508_),
    .Q(\mem.mem_internal.code_mem[229][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[229][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2503),
    .D(_01265_),
    .Q_N(_14507_),
    .Q(\mem.mem_internal.code_mem[229][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[22][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2504),
    .D(_01266_),
    .Q_N(_14506_),
    .Q(\mem.mem_internal.code_mem[22][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[22][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2505),
    .D(_01267_),
    .Q_N(_14505_),
    .Q(\mem.mem_internal.code_mem[22][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[22][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2506),
    .D(_01268_),
    .Q_N(_14504_),
    .Q(\mem.mem_internal.code_mem[22][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[22][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2507),
    .D(_01269_),
    .Q_N(_14503_),
    .Q(\mem.mem_internal.code_mem[22][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[22][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2508),
    .D(_01270_),
    .Q_N(_14502_),
    .Q(\mem.mem_internal.code_mem[22][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[22][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2509),
    .D(_01271_),
    .Q_N(_14501_),
    .Q(\mem.mem_internal.code_mem[22][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[22][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2510),
    .D(_01272_),
    .Q_N(_14500_),
    .Q(\mem.mem_internal.code_mem[22][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[22][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2511),
    .D(_01273_),
    .Q_N(_14499_),
    .Q(\mem.mem_internal.code_mem[22][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[230][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2512),
    .D(_01274_),
    .Q_N(_14498_),
    .Q(\mem.mem_internal.code_mem[230][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[230][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2513),
    .D(_01275_),
    .Q_N(_14497_),
    .Q(\mem.mem_internal.code_mem[230][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[230][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2514),
    .D(_01276_),
    .Q_N(_14496_),
    .Q(\mem.mem_internal.code_mem[230][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[230][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2515),
    .D(_01277_),
    .Q_N(_14495_),
    .Q(\mem.mem_internal.code_mem[230][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[230][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2516),
    .D(_01278_),
    .Q_N(_14494_),
    .Q(\mem.mem_internal.code_mem[230][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[230][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2517),
    .D(_01279_),
    .Q_N(_14493_),
    .Q(\mem.mem_internal.code_mem[230][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[230][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2518),
    .D(_01280_),
    .Q_N(_14492_),
    .Q(\mem.mem_internal.code_mem[230][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[230][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2519),
    .D(_01281_),
    .Q_N(_14491_),
    .Q(\mem.mem_internal.code_mem[230][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[231][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2520),
    .D(_01282_),
    .Q_N(_14490_),
    .Q(\mem.mem_internal.code_mem[231][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[231][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2521),
    .D(_01283_),
    .Q_N(_14489_),
    .Q(\mem.mem_internal.code_mem[231][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[231][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2522),
    .D(_01284_),
    .Q_N(_14488_),
    .Q(\mem.mem_internal.code_mem[231][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[231][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2523),
    .D(_01285_),
    .Q_N(_14487_),
    .Q(\mem.mem_internal.code_mem[231][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[231][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2524),
    .D(_01286_),
    .Q_N(_14486_),
    .Q(\mem.mem_internal.code_mem[231][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[231][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2525),
    .D(_01287_),
    .Q_N(_14485_),
    .Q(\mem.mem_internal.code_mem[231][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[231][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2526),
    .D(_01288_),
    .Q_N(_14484_),
    .Q(\mem.mem_internal.code_mem[231][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[231][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2527),
    .D(_01289_),
    .Q_N(_14483_),
    .Q(\mem.mem_internal.code_mem[231][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[232][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2528),
    .D(_01290_),
    .Q_N(_14482_),
    .Q(\mem.mem_internal.code_mem[232][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[232][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2529),
    .D(_01291_),
    .Q_N(_14481_),
    .Q(\mem.mem_internal.code_mem[232][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[232][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2530),
    .D(_01292_),
    .Q_N(_14480_),
    .Q(\mem.mem_internal.code_mem[232][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[232][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2531),
    .D(_01293_),
    .Q_N(_14479_),
    .Q(\mem.mem_internal.code_mem[232][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[232][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2532),
    .D(_01294_),
    .Q_N(_14478_),
    .Q(\mem.mem_internal.code_mem[232][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[232][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2533),
    .D(_01295_),
    .Q_N(_14477_),
    .Q(\mem.mem_internal.code_mem[232][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[232][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2534),
    .D(_01296_),
    .Q_N(_14476_),
    .Q(\mem.mem_internal.code_mem[232][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[232][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2535),
    .D(_01297_),
    .Q_N(_14475_),
    .Q(\mem.mem_internal.code_mem[232][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[233][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2536),
    .D(_01298_),
    .Q_N(_14474_),
    .Q(\mem.mem_internal.code_mem[233][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[233][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2537),
    .D(_01299_),
    .Q_N(_14473_),
    .Q(\mem.mem_internal.code_mem[233][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[233][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2538),
    .D(_01300_),
    .Q_N(_14472_),
    .Q(\mem.mem_internal.code_mem[233][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[233][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2539),
    .D(_01301_),
    .Q_N(_14471_),
    .Q(\mem.mem_internal.code_mem[233][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[233][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2540),
    .D(_01302_),
    .Q_N(_14470_),
    .Q(\mem.mem_internal.code_mem[233][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[233][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2541),
    .D(_01303_),
    .Q_N(_14469_),
    .Q(\mem.mem_internal.code_mem[233][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[233][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2542),
    .D(_01304_),
    .Q_N(_14468_),
    .Q(\mem.mem_internal.code_mem[233][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[233][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2543),
    .D(_01305_),
    .Q_N(_14467_),
    .Q(\mem.mem_internal.code_mem[233][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[234][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2544),
    .D(_01306_),
    .Q_N(_14466_),
    .Q(\mem.mem_internal.code_mem[234][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[234][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2545),
    .D(_01307_),
    .Q_N(_14465_),
    .Q(\mem.mem_internal.code_mem[234][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[234][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2546),
    .D(_01308_),
    .Q_N(_14464_),
    .Q(\mem.mem_internal.code_mem[234][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[234][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2547),
    .D(_01309_),
    .Q_N(_14463_),
    .Q(\mem.mem_internal.code_mem[234][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[234][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2548),
    .D(_01310_),
    .Q_N(_14462_),
    .Q(\mem.mem_internal.code_mem[234][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[234][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2549),
    .D(_01311_),
    .Q_N(_14461_),
    .Q(\mem.mem_internal.code_mem[234][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[234][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2550),
    .D(_01312_),
    .Q_N(_14460_),
    .Q(\mem.mem_internal.code_mem[234][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[234][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2551),
    .D(_01313_),
    .Q_N(_14459_),
    .Q(\mem.mem_internal.code_mem[234][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[235][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2552),
    .D(_01314_),
    .Q_N(_14458_),
    .Q(\mem.mem_internal.code_mem[235][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[235][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2553),
    .D(_01315_),
    .Q_N(_14457_),
    .Q(\mem.mem_internal.code_mem[235][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[235][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2554),
    .D(_01316_),
    .Q_N(_14456_),
    .Q(\mem.mem_internal.code_mem[235][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[235][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2555),
    .D(_01317_),
    .Q_N(_14455_),
    .Q(\mem.mem_internal.code_mem[235][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[235][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2556),
    .D(_01318_),
    .Q_N(_14454_),
    .Q(\mem.mem_internal.code_mem[235][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[235][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2557),
    .D(_01319_),
    .Q_N(_14453_),
    .Q(\mem.mem_internal.code_mem[235][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[235][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2558),
    .D(_01320_),
    .Q_N(_14452_),
    .Q(\mem.mem_internal.code_mem[235][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[235][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2559),
    .D(_01321_),
    .Q_N(_14451_),
    .Q(\mem.mem_internal.code_mem[235][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[236][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2560),
    .D(_01322_),
    .Q_N(_14450_),
    .Q(\mem.mem_internal.code_mem[236][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[236][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2561),
    .D(_01323_),
    .Q_N(_14449_),
    .Q(\mem.mem_internal.code_mem[236][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[236][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2562),
    .D(_01324_),
    .Q_N(_14448_),
    .Q(\mem.mem_internal.code_mem[236][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[236][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2563),
    .D(_01325_),
    .Q_N(_14447_),
    .Q(\mem.mem_internal.code_mem[236][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[236][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2564),
    .D(_01326_),
    .Q_N(_14446_),
    .Q(\mem.mem_internal.code_mem[236][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[236][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2565),
    .D(_01327_),
    .Q_N(_14445_),
    .Q(\mem.mem_internal.code_mem[236][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[236][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2566),
    .D(_01328_),
    .Q_N(_14444_),
    .Q(\mem.mem_internal.code_mem[236][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[236][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2567),
    .D(_01329_),
    .Q_N(_14443_),
    .Q(\mem.mem_internal.code_mem[236][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[237][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2568),
    .D(_01330_),
    .Q_N(_14442_),
    .Q(\mem.mem_internal.code_mem[237][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[237][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2569),
    .D(_01331_),
    .Q_N(_14441_),
    .Q(\mem.mem_internal.code_mem[237][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[237][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2570),
    .D(_01332_),
    .Q_N(_14440_),
    .Q(\mem.mem_internal.code_mem[237][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[237][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2571),
    .D(_01333_),
    .Q_N(_14439_),
    .Q(\mem.mem_internal.code_mem[237][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[237][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2572),
    .D(_01334_),
    .Q_N(_14438_),
    .Q(\mem.mem_internal.code_mem[237][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[237][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2573),
    .D(_01335_),
    .Q_N(_14437_),
    .Q(\mem.mem_internal.code_mem[237][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[237][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2574),
    .D(_01336_),
    .Q_N(_14436_),
    .Q(\mem.mem_internal.code_mem[237][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[237][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2575),
    .D(_01337_),
    .Q_N(_14435_),
    .Q(\mem.mem_internal.code_mem[237][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[238][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2576),
    .D(_01338_),
    .Q_N(_14434_),
    .Q(\mem.mem_internal.code_mem[238][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[238][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2577),
    .D(_01339_),
    .Q_N(_14433_),
    .Q(\mem.mem_internal.code_mem[238][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[238][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2578),
    .D(_01340_),
    .Q_N(_14432_),
    .Q(\mem.mem_internal.code_mem[238][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[238][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2579),
    .D(_01341_),
    .Q_N(_14431_),
    .Q(\mem.mem_internal.code_mem[238][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[238][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2580),
    .D(_01342_),
    .Q_N(_14430_),
    .Q(\mem.mem_internal.code_mem[238][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[238][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2581),
    .D(_01343_),
    .Q_N(_14429_),
    .Q(\mem.mem_internal.code_mem[238][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[238][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2582),
    .D(_01344_),
    .Q_N(_14428_),
    .Q(\mem.mem_internal.code_mem[238][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[238][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2583),
    .D(_01345_),
    .Q_N(_14427_),
    .Q(\mem.mem_internal.code_mem[238][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[239][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2584),
    .D(_01346_),
    .Q_N(_14426_),
    .Q(\mem.mem_internal.code_mem[239][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[239][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2585),
    .D(_01347_),
    .Q_N(_14425_),
    .Q(\mem.mem_internal.code_mem[239][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[239][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2586),
    .D(_01348_),
    .Q_N(_14424_),
    .Q(\mem.mem_internal.code_mem[239][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[239][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2587),
    .D(_01349_),
    .Q_N(_14423_),
    .Q(\mem.mem_internal.code_mem[239][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[239][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2588),
    .D(_01350_),
    .Q_N(_14422_),
    .Q(\mem.mem_internal.code_mem[239][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[239][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2589),
    .D(_01351_),
    .Q_N(_14421_),
    .Q(\mem.mem_internal.code_mem[239][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[239][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2590),
    .D(_01352_),
    .Q_N(_14420_),
    .Q(\mem.mem_internal.code_mem[239][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[239][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2591),
    .D(_01353_),
    .Q_N(_14419_),
    .Q(\mem.mem_internal.code_mem[239][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[23][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2592),
    .D(_01354_),
    .Q_N(_14418_),
    .Q(\mem.mem_internal.code_mem[23][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[23][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2593),
    .D(_01355_),
    .Q_N(_14417_),
    .Q(\mem.mem_internal.code_mem[23][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[23][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2594),
    .D(_01356_),
    .Q_N(_14416_),
    .Q(\mem.mem_internal.code_mem[23][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[23][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2595),
    .D(_01357_),
    .Q_N(_14415_),
    .Q(\mem.mem_internal.code_mem[23][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[23][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2596),
    .D(_01358_),
    .Q_N(_14414_),
    .Q(\mem.mem_internal.code_mem[23][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[23][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2597),
    .D(_01359_),
    .Q_N(_14413_),
    .Q(\mem.mem_internal.code_mem[23][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[23][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2598),
    .D(_01360_),
    .Q_N(_14412_),
    .Q(\mem.mem_internal.code_mem[23][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[23][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2599),
    .D(_01361_),
    .Q_N(_14411_),
    .Q(\mem.mem_internal.code_mem[23][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[240][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2600),
    .D(_01362_),
    .Q_N(_14410_),
    .Q(\mem.mem_internal.code_mem[240][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[240][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2601),
    .D(_01363_),
    .Q_N(_14409_),
    .Q(\mem.mem_internal.code_mem[240][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[240][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2602),
    .D(_01364_),
    .Q_N(_14408_),
    .Q(\mem.mem_internal.code_mem[240][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[240][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2603),
    .D(_01365_),
    .Q_N(_14407_),
    .Q(\mem.mem_internal.code_mem[240][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[240][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2604),
    .D(_01366_),
    .Q_N(_14406_),
    .Q(\mem.mem_internal.code_mem[240][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[240][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2605),
    .D(_01367_),
    .Q_N(_14405_),
    .Q(\mem.mem_internal.code_mem[240][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[240][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2606),
    .D(_01368_),
    .Q_N(_14404_),
    .Q(\mem.mem_internal.code_mem[240][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[240][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2607),
    .D(_01369_),
    .Q_N(_14403_),
    .Q(\mem.mem_internal.code_mem[240][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[241][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2608),
    .D(_01370_),
    .Q_N(_14402_),
    .Q(\mem.mem_internal.code_mem[241][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[241][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2609),
    .D(_01371_),
    .Q_N(_14401_),
    .Q(\mem.mem_internal.code_mem[241][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[241][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2610),
    .D(_01372_),
    .Q_N(_14400_),
    .Q(\mem.mem_internal.code_mem[241][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[241][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2611),
    .D(_01373_),
    .Q_N(_14399_),
    .Q(\mem.mem_internal.code_mem[241][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[241][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2612),
    .D(_01374_),
    .Q_N(_14398_),
    .Q(\mem.mem_internal.code_mem[241][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[241][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2613),
    .D(_01375_),
    .Q_N(_14397_),
    .Q(\mem.mem_internal.code_mem[241][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[241][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2614),
    .D(_01376_),
    .Q_N(_14396_),
    .Q(\mem.mem_internal.code_mem[241][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[241][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2615),
    .D(_01377_),
    .Q_N(_14395_),
    .Q(\mem.mem_internal.code_mem[241][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[242][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2616),
    .D(_01378_),
    .Q_N(_14394_),
    .Q(\mem.mem_internal.code_mem[242][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[242][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2617),
    .D(_01379_),
    .Q_N(_14393_),
    .Q(\mem.mem_internal.code_mem[242][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[242][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2618),
    .D(_01380_),
    .Q_N(_14392_),
    .Q(\mem.mem_internal.code_mem[242][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[242][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2619),
    .D(_01381_),
    .Q_N(_14391_),
    .Q(\mem.mem_internal.code_mem[242][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[242][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2620),
    .D(_01382_),
    .Q_N(_14390_),
    .Q(\mem.mem_internal.code_mem[242][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[242][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2621),
    .D(_01383_),
    .Q_N(_14389_),
    .Q(\mem.mem_internal.code_mem[242][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[242][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2622),
    .D(_01384_),
    .Q_N(_14388_),
    .Q(\mem.mem_internal.code_mem[242][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[242][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2623),
    .D(_01385_),
    .Q_N(_14387_),
    .Q(\mem.mem_internal.code_mem[242][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[243][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2624),
    .D(_01386_),
    .Q_N(_14386_),
    .Q(\mem.mem_internal.code_mem[243][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[243][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2625),
    .D(_01387_),
    .Q_N(_14385_),
    .Q(\mem.mem_internal.code_mem[243][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[243][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2626),
    .D(_01388_),
    .Q_N(_14384_),
    .Q(\mem.mem_internal.code_mem[243][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[243][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2627),
    .D(_01389_),
    .Q_N(_14383_),
    .Q(\mem.mem_internal.code_mem[243][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[243][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2628),
    .D(_01390_),
    .Q_N(_14382_),
    .Q(\mem.mem_internal.code_mem[243][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[243][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2629),
    .D(_01391_),
    .Q_N(_14381_),
    .Q(\mem.mem_internal.code_mem[243][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[243][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2630),
    .D(_01392_),
    .Q_N(_14380_),
    .Q(\mem.mem_internal.code_mem[243][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[243][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2631),
    .D(_01393_),
    .Q_N(_14379_),
    .Q(\mem.mem_internal.code_mem[243][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[244][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2632),
    .D(_01394_),
    .Q_N(_14378_),
    .Q(\mem.mem_internal.code_mem[244][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[244][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2633),
    .D(_01395_),
    .Q_N(_14377_),
    .Q(\mem.mem_internal.code_mem[244][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[244][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2634),
    .D(_01396_),
    .Q_N(_14376_),
    .Q(\mem.mem_internal.code_mem[244][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[244][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2635),
    .D(_01397_),
    .Q_N(_14375_),
    .Q(\mem.mem_internal.code_mem[244][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[244][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2636),
    .D(_01398_),
    .Q_N(_14374_),
    .Q(\mem.mem_internal.code_mem[244][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[244][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2637),
    .D(_01399_),
    .Q_N(_14373_),
    .Q(\mem.mem_internal.code_mem[244][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[244][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2638),
    .D(_01400_),
    .Q_N(_14372_),
    .Q(\mem.mem_internal.code_mem[244][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[244][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2639),
    .D(_01401_),
    .Q_N(_14371_),
    .Q(\mem.mem_internal.code_mem[244][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[245][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2640),
    .D(_01402_),
    .Q_N(_14370_),
    .Q(\mem.mem_internal.code_mem[245][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[245][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2641),
    .D(_01403_),
    .Q_N(_14369_),
    .Q(\mem.mem_internal.code_mem[245][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[245][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2642),
    .D(_01404_),
    .Q_N(_14368_),
    .Q(\mem.mem_internal.code_mem[245][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[245][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2643),
    .D(_01405_),
    .Q_N(_14367_),
    .Q(\mem.mem_internal.code_mem[245][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[245][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2644),
    .D(_01406_),
    .Q_N(_14366_),
    .Q(\mem.mem_internal.code_mem[245][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[245][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2645),
    .D(_01407_),
    .Q_N(_14365_),
    .Q(\mem.mem_internal.code_mem[245][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[245][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2646),
    .D(_01408_),
    .Q_N(_14364_),
    .Q(\mem.mem_internal.code_mem[245][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[245][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2647),
    .D(_01409_),
    .Q_N(_14363_),
    .Q(\mem.mem_internal.code_mem[245][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[246][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2648),
    .D(_01410_),
    .Q_N(_14362_),
    .Q(\mem.mem_internal.code_mem[246][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[246][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2649),
    .D(_01411_),
    .Q_N(_14361_),
    .Q(\mem.mem_internal.code_mem[246][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[246][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2650),
    .D(_01412_),
    .Q_N(_14360_),
    .Q(\mem.mem_internal.code_mem[246][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[246][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2651),
    .D(_01413_),
    .Q_N(_14359_),
    .Q(\mem.mem_internal.code_mem[246][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[246][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2652),
    .D(_01414_),
    .Q_N(_14358_),
    .Q(\mem.mem_internal.code_mem[246][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[246][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2653),
    .D(_01415_),
    .Q_N(_14357_),
    .Q(\mem.mem_internal.code_mem[246][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[246][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2654),
    .D(_01416_),
    .Q_N(_14356_),
    .Q(\mem.mem_internal.code_mem[246][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[246][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2655),
    .D(_01417_),
    .Q_N(_14355_),
    .Q(\mem.mem_internal.code_mem[246][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[247][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2656),
    .D(_01418_),
    .Q_N(_14354_),
    .Q(\mem.mem_internal.code_mem[247][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[247][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2657),
    .D(_01419_),
    .Q_N(_14353_),
    .Q(\mem.mem_internal.code_mem[247][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[247][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2658),
    .D(_01420_),
    .Q_N(_14352_),
    .Q(\mem.mem_internal.code_mem[247][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[247][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2659),
    .D(_01421_),
    .Q_N(_14351_),
    .Q(\mem.mem_internal.code_mem[247][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[247][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2660),
    .D(_01422_),
    .Q_N(_14350_),
    .Q(\mem.mem_internal.code_mem[247][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[247][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2661),
    .D(_01423_),
    .Q_N(_14349_),
    .Q(\mem.mem_internal.code_mem[247][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[247][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2662),
    .D(_01424_),
    .Q_N(_14348_),
    .Q(\mem.mem_internal.code_mem[247][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[247][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2663),
    .D(_01425_),
    .Q_N(_14347_),
    .Q(\mem.mem_internal.code_mem[247][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[248][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2664),
    .D(_01426_),
    .Q_N(_14346_),
    .Q(\mem.mem_internal.code_mem[248][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[248][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2665),
    .D(_01427_),
    .Q_N(_14345_),
    .Q(\mem.mem_internal.code_mem[248][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[248][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2666),
    .D(_01428_),
    .Q_N(_14344_),
    .Q(\mem.mem_internal.code_mem[248][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[248][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2667),
    .D(_01429_),
    .Q_N(_14343_),
    .Q(\mem.mem_internal.code_mem[248][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[248][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2668),
    .D(_01430_),
    .Q_N(_14342_),
    .Q(\mem.mem_internal.code_mem[248][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[248][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2669),
    .D(_01431_),
    .Q_N(_14341_),
    .Q(\mem.mem_internal.code_mem[248][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[248][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2670),
    .D(_01432_),
    .Q_N(_14340_),
    .Q(\mem.mem_internal.code_mem[248][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[248][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2671),
    .D(_01433_),
    .Q_N(_14339_),
    .Q(\mem.mem_internal.code_mem[248][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[249][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2672),
    .D(_01434_),
    .Q_N(_14338_),
    .Q(\mem.mem_internal.code_mem[249][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[249][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2673),
    .D(_01435_),
    .Q_N(_14337_),
    .Q(\mem.mem_internal.code_mem[249][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[249][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2674),
    .D(_01436_),
    .Q_N(_14336_),
    .Q(\mem.mem_internal.code_mem[249][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[249][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2675),
    .D(_01437_),
    .Q_N(_14335_),
    .Q(\mem.mem_internal.code_mem[249][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[249][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2676),
    .D(_01438_),
    .Q_N(_14334_),
    .Q(\mem.mem_internal.code_mem[249][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[249][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2677),
    .D(_01439_),
    .Q_N(_14333_),
    .Q(\mem.mem_internal.code_mem[249][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[249][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2678),
    .D(_01440_),
    .Q_N(_14332_),
    .Q(\mem.mem_internal.code_mem[249][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[249][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2679),
    .D(_01441_),
    .Q_N(_14331_),
    .Q(\mem.mem_internal.code_mem[249][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[24][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2680),
    .D(_01442_),
    .Q_N(_14330_),
    .Q(\mem.mem_internal.code_mem[24][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[24][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2681),
    .D(_01443_),
    .Q_N(_14329_),
    .Q(\mem.mem_internal.code_mem[24][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[24][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2682),
    .D(_01444_),
    .Q_N(_14328_),
    .Q(\mem.mem_internal.code_mem[24][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[24][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2683),
    .D(_01445_),
    .Q_N(_14327_),
    .Q(\mem.mem_internal.code_mem[24][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[24][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2684),
    .D(_01446_),
    .Q_N(_14326_),
    .Q(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[24][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2685),
    .D(_01447_),
    .Q_N(_14325_),
    .Q(\mem.mem_internal.code_mem[24][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[24][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2686),
    .D(_01448_),
    .Q_N(_14324_),
    .Q(\mem.mem_internal.code_mem[24][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[24][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2687),
    .D(_01449_),
    .Q_N(_14323_),
    .Q(\mem.mem_internal.code_mem[24][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[250][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2688),
    .D(_01450_),
    .Q_N(_14322_),
    .Q(\mem.mem_internal.code_mem[250][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[250][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2689),
    .D(_01451_),
    .Q_N(_14321_),
    .Q(\mem.mem_internal.code_mem[250][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[250][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2690),
    .D(_01452_),
    .Q_N(_14320_),
    .Q(\mem.mem_internal.code_mem[250][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[250][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2691),
    .D(_01453_),
    .Q_N(_14319_),
    .Q(\mem.mem_internal.code_mem[250][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[250][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2692),
    .D(_01454_),
    .Q_N(_14318_),
    .Q(\mem.mem_internal.code_mem[250][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[250][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2693),
    .D(_01455_),
    .Q_N(_14317_),
    .Q(\mem.mem_internal.code_mem[250][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[250][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2694),
    .D(_01456_),
    .Q_N(_14316_),
    .Q(\mem.mem_internal.code_mem[250][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[250][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2695),
    .D(_01457_),
    .Q_N(_14315_),
    .Q(\mem.mem_internal.code_mem[250][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[251][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2696),
    .D(_01458_),
    .Q_N(_14314_),
    .Q(\mem.mem_internal.code_mem[251][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[251][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2697),
    .D(_01459_),
    .Q_N(_14313_),
    .Q(\mem.mem_internal.code_mem[251][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[251][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2698),
    .D(_01460_),
    .Q_N(_14312_),
    .Q(\mem.mem_internal.code_mem[251][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[251][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2699),
    .D(_01461_),
    .Q_N(_14311_),
    .Q(\mem.mem_internal.code_mem[251][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[251][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2700),
    .D(_01462_),
    .Q_N(_14310_),
    .Q(\mem.mem_internal.code_mem[251][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[251][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2701),
    .D(_01463_),
    .Q_N(_14309_),
    .Q(\mem.mem_internal.code_mem[251][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[251][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2702),
    .D(_01464_),
    .Q_N(_14308_),
    .Q(\mem.mem_internal.code_mem[251][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[251][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2703),
    .D(_01465_),
    .Q_N(_14307_),
    .Q(\mem.mem_internal.code_mem[251][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[252][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2704),
    .D(_01466_),
    .Q_N(_14306_),
    .Q(\mem.mem_internal.code_mem[252][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[252][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2705),
    .D(_01467_),
    .Q_N(_14305_),
    .Q(\mem.mem_internal.code_mem[252][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[252][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2706),
    .D(_01468_),
    .Q_N(_14304_),
    .Q(\mem.mem_internal.code_mem[252][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[252][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2707),
    .D(_01469_),
    .Q_N(_14303_),
    .Q(\mem.mem_internal.code_mem[252][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[252][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2708),
    .D(_01470_),
    .Q_N(_14302_),
    .Q(\mem.mem_internal.code_mem[252][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[252][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2709),
    .D(_01471_),
    .Q_N(_14301_),
    .Q(\mem.mem_internal.code_mem[252][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[252][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2710),
    .D(_01472_),
    .Q_N(_14300_),
    .Q(\mem.mem_internal.code_mem[252][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[252][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2711),
    .D(_01473_),
    .Q_N(_14299_),
    .Q(\mem.mem_internal.code_mem[252][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[253][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2712),
    .D(_01474_),
    .Q_N(_14298_),
    .Q(\mem.mem_internal.code_mem[253][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[253][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2713),
    .D(_01475_),
    .Q_N(_14297_),
    .Q(\mem.mem_internal.code_mem[253][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[253][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2714),
    .D(_01476_),
    .Q_N(_14296_),
    .Q(\mem.mem_internal.code_mem[253][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[253][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2715),
    .D(_01477_),
    .Q_N(_14295_),
    .Q(\mem.mem_internal.code_mem[253][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[253][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2716),
    .D(_01478_),
    .Q_N(_14294_),
    .Q(\mem.mem_internal.code_mem[253][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[253][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2717),
    .D(_01479_),
    .Q_N(_14293_),
    .Q(\mem.mem_internal.code_mem[253][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[253][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2718),
    .D(_01480_),
    .Q_N(_14292_),
    .Q(\mem.mem_internal.code_mem[253][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[253][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2719),
    .D(_01481_),
    .Q_N(_14291_),
    .Q(\mem.mem_internal.code_mem[253][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[254][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2720),
    .D(_01482_),
    .Q_N(_14290_),
    .Q(\mem.mem_internal.code_mem[254][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[254][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2721),
    .D(_01483_),
    .Q_N(_14289_),
    .Q(\mem.mem_internal.code_mem[254][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[254][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2722),
    .D(_01484_),
    .Q_N(_14288_),
    .Q(\mem.mem_internal.code_mem[254][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[254][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2723),
    .D(_01485_),
    .Q_N(_14287_),
    .Q(\mem.mem_internal.code_mem[254][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[254][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2724),
    .D(_01486_),
    .Q_N(_14286_),
    .Q(\mem.mem_internal.code_mem[254][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[254][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2725),
    .D(_01487_),
    .Q_N(_14285_),
    .Q(\mem.mem_internal.code_mem[254][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[254][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2726),
    .D(_01488_),
    .Q_N(_14284_),
    .Q(\mem.mem_internal.code_mem[254][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[254][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2727),
    .D(_01489_),
    .Q_N(_14283_),
    .Q(\mem.mem_internal.code_mem[254][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[255][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2728),
    .D(_01490_),
    .Q_N(_14282_),
    .Q(\mem.mem_internal.code_mem[255][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[255][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2729),
    .D(_01491_),
    .Q_N(_14281_),
    .Q(\mem.mem_internal.code_mem[255][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[255][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2730),
    .D(_01492_),
    .Q_N(_14280_),
    .Q(\mem.mem_internal.code_mem[255][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[255][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2731),
    .D(_01493_),
    .Q_N(_14279_),
    .Q(\mem.mem_internal.code_mem[255][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[255][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2732),
    .D(_01494_),
    .Q_N(_14278_),
    .Q(\mem.mem_internal.code_mem[255][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[255][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2733),
    .D(_01495_),
    .Q_N(_14277_),
    .Q(\mem.mem_internal.code_mem[255][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[255][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2734),
    .D(_01496_),
    .Q_N(_14276_),
    .Q(\mem.mem_internal.code_mem[255][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[255][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2735),
    .D(_01497_),
    .Q_N(_14275_),
    .Q(\mem.mem_internal.code_mem[255][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[25][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2736),
    .D(_01498_),
    .Q_N(_14274_),
    .Q(\mem.mem_internal.code_mem[25][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[25][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2737),
    .D(_01499_),
    .Q_N(_14273_),
    .Q(\mem.mem_internal.code_mem[25][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[25][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2738),
    .D(_01500_),
    .Q_N(_14272_),
    .Q(\mem.mem_internal.code_mem[25][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[25][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2739),
    .D(_01501_),
    .Q_N(_14271_),
    .Q(\mem.mem_internal.code_mem[25][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[25][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2740),
    .D(_01502_),
    .Q_N(_14270_),
    .Q(\mem.mem_internal.code_mem[25][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[25][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2741),
    .D(_01503_),
    .Q_N(_14269_),
    .Q(\mem.mem_internal.code_mem[25][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[25][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2742),
    .D(_01504_),
    .Q_N(_14268_),
    .Q(\mem.mem_internal.code_mem[25][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[25][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2743),
    .D(_01505_),
    .Q_N(_14267_),
    .Q(\mem.mem_internal.code_mem[25][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[26][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2744),
    .D(_01506_),
    .Q_N(_14266_),
    .Q(\mem.mem_internal.code_mem[26][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[26][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2745),
    .D(_01507_),
    .Q_N(_14265_),
    .Q(\mem.mem_internal.code_mem[26][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[26][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2746),
    .D(_01508_),
    .Q_N(_14264_),
    .Q(\mem.mem_internal.code_mem[26][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[26][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2747),
    .D(_01509_),
    .Q_N(_14263_),
    .Q(\mem.mem_internal.code_mem[26][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[26][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2748),
    .D(_01510_),
    .Q_N(_14262_),
    .Q(\mem.mem_internal.code_mem[26][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[26][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2749),
    .D(_01511_),
    .Q_N(_14261_),
    .Q(\mem.mem_internal.code_mem[26][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[26][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2750),
    .D(_01512_),
    .Q_N(_14260_),
    .Q(\mem.mem_internal.code_mem[26][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[26][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2751),
    .D(_01513_),
    .Q_N(_14259_),
    .Q(\mem.mem_internal.code_mem[26][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[27][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2752),
    .D(_01514_),
    .Q_N(_14258_),
    .Q(\mem.mem_internal.code_mem[27][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[27][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2753),
    .D(_01515_),
    .Q_N(_14257_),
    .Q(\mem.mem_internal.code_mem[27][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[27][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2754),
    .D(_01516_),
    .Q_N(_14256_),
    .Q(\mem.mem_internal.code_mem[27][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[27][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2755),
    .D(_01517_),
    .Q_N(_14255_),
    .Q(\mem.mem_internal.code_mem[27][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[27][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2756),
    .D(_01518_),
    .Q_N(_14254_),
    .Q(\mem.mem_internal.code_mem[27][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[27][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2757),
    .D(_01519_),
    .Q_N(_14253_),
    .Q(\mem.mem_internal.code_mem[27][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[27][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2758),
    .D(_01520_),
    .Q_N(_14252_),
    .Q(\mem.mem_internal.code_mem[27][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[27][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2759),
    .D(_01521_),
    .Q_N(_14251_),
    .Q(\mem.mem_internal.code_mem[27][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[28][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2760),
    .D(_01522_),
    .Q_N(_14250_),
    .Q(\mem.mem_internal.code_mem[28][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[28][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2761),
    .D(_01523_),
    .Q_N(_14249_),
    .Q(\mem.mem_internal.code_mem[28][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[28][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2762),
    .D(_01524_),
    .Q_N(_14248_),
    .Q(\mem.mem_internal.code_mem[28][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[28][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2763),
    .D(_01525_),
    .Q_N(_14247_),
    .Q(\mem.mem_internal.code_mem[28][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[28][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2764),
    .D(_01526_),
    .Q_N(_14246_),
    .Q(\mem.mem_internal.code_mem[28][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[28][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2765),
    .D(_01527_),
    .Q_N(_14245_),
    .Q(\mem.mem_internal.code_mem[28][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[28][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2766),
    .D(_01528_),
    .Q_N(_14244_),
    .Q(\mem.mem_internal.code_mem[28][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[28][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2767),
    .D(_01529_),
    .Q_N(_14243_),
    .Q(\mem.mem_internal.code_mem[28][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[29][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2768),
    .D(_01530_),
    .Q_N(_14242_),
    .Q(\mem.mem_internal.code_mem[29][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[29][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2769),
    .D(_01531_),
    .Q_N(_14241_),
    .Q(\mem.mem_internal.code_mem[29][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[29][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2770),
    .D(_01532_),
    .Q_N(_14240_),
    .Q(\mem.mem_internal.code_mem[29][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[29][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2771),
    .D(_01533_),
    .Q_N(_14239_),
    .Q(\mem.mem_internal.code_mem[29][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[29][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2772),
    .D(_01534_),
    .Q_N(_14238_),
    .Q(\mem.mem_internal.code_mem[29][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[29][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2773),
    .D(_01535_),
    .Q_N(_14237_),
    .Q(\mem.mem_internal.code_mem[29][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[29][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2774),
    .D(_01536_),
    .Q_N(_14236_),
    .Q(\mem.mem_internal.code_mem[29][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[29][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2775),
    .D(_01537_),
    .Q_N(_14235_),
    .Q(\mem.mem_internal.code_mem[29][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2776),
    .D(_01538_),
    .Q_N(_14234_),
    .Q(\mem.mem_internal.code_mem[2][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2777),
    .D(_01539_),
    .Q_N(_14233_),
    .Q(\mem.mem_internal.code_mem[2][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[2][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2778),
    .D(_01540_),
    .Q_N(_14232_),
    .Q(\mem.mem_internal.code_mem[2][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2779),
    .D(_01541_),
    .Q_N(_14231_),
    .Q(\mem.mem_internal.code_mem[2][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[2][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2780),
    .D(_01542_),
    .Q_N(_14230_),
    .Q(\mem.mem_internal.code_mem[2][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[2][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2781),
    .D(_01543_),
    .Q_N(_14229_),
    .Q(\mem.mem_internal.code_mem[2][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[2][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2782),
    .D(_01544_),
    .Q_N(_14228_),
    .Q(\mem.mem_internal.code_mem[2][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[2][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2783),
    .D(_01545_),
    .Q_N(_14227_),
    .Q(\mem.mem_internal.code_mem[2][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[30][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2784),
    .D(_01546_),
    .Q_N(_14226_),
    .Q(\mem.mem_internal.code_mem[30][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[30][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2785),
    .D(_01547_),
    .Q_N(_14225_),
    .Q(\mem.mem_internal.code_mem[30][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[30][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2786),
    .D(_01548_),
    .Q_N(_14224_),
    .Q(\mem.mem_internal.code_mem[30][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[30][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2787),
    .D(_01549_),
    .Q_N(_14223_),
    .Q(\mem.mem_internal.code_mem[30][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[30][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2788),
    .D(_01550_),
    .Q_N(_14222_),
    .Q(\mem.mem_internal.code_mem[30][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[30][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2789),
    .D(_01551_),
    .Q_N(_14221_),
    .Q(\mem.mem_internal.code_mem[30][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[30][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2790),
    .D(_01552_),
    .Q_N(_14220_),
    .Q(\mem.mem_internal.code_mem[30][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[30][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2791),
    .D(_01553_),
    .Q_N(_14219_),
    .Q(\mem.mem_internal.code_mem[30][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[31][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2792),
    .D(_01554_),
    .Q_N(_14218_),
    .Q(\mem.mem_internal.code_mem[31][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[31][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2793),
    .D(_01555_),
    .Q_N(_14217_),
    .Q(\mem.mem_internal.code_mem[31][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[31][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2794),
    .D(_01556_),
    .Q_N(_14216_),
    .Q(\mem.mem_internal.code_mem[31][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[31][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2795),
    .D(_01557_),
    .Q_N(_14215_),
    .Q(\mem.mem_internal.code_mem[31][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[31][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2796),
    .D(_01558_),
    .Q_N(_14214_),
    .Q(\mem.mem_internal.code_mem[31][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[31][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2797),
    .D(_01559_),
    .Q_N(_14213_),
    .Q(\mem.mem_internal.code_mem[31][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[31][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2798),
    .D(_01560_),
    .Q_N(_14212_),
    .Q(\mem.mem_internal.code_mem[31][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[31][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2799),
    .D(_01561_),
    .Q_N(_14211_),
    .Q(\mem.mem_internal.code_mem[31][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[32][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2800),
    .D(_01562_),
    .Q_N(_14210_),
    .Q(\mem.mem_internal.code_mem[32][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[32][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2801),
    .D(_01563_),
    .Q_N(_14209_),
    .Q(\mem.mem_internal.code_mem[32][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[32][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2802),
    .D(_01564_),
    .Q_N(_14208_),
    .Q(\mem.mem_internal.code_mem[32][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[32][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2803),
    .D(_01565_),
    .Q_N(_14207_),
    .Q(\mem.mem_internal.code_mem[32][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[32][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2804),
    .D(_01566_),
    .Q_N(_14206_),
    .Q(\mem.mem_internal.code_mem[32][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[32][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2805),
    .D(_01567_),
    .Q_N(_14205_),
    .Q(\mem.mem_internal.code_mem[32][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[32][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2806),
    .D(_01568_),
    .Q_N(_14204_),
    .Q(\mem.mem_internal.code_mem[32][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[32][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2807),
    .D(_01569_),
    .Q_N(_14203_),
    .Q(\mem.mem_internal.code_mem[32][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[33][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2808),
    .D(_01570_),
    .Q_N(_14202_),
    .Q(\mem.mem_internal.code_mem[33][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[33][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2809),
    .D(_01571_),
    .Q_N(_14201_),
    .Q(\mem.mem_internal.code_mem[33][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[33][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2810),
    .D(_01572_),
    .Q_N(_14200_),
    .Q(\mem.mem_internal.code_mem[33][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[33][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2811),
    .D(_01573_),
    .Q_N(_14199_),
    .Q(\mem.mem_internal.code_mem[33][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[33][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2812),
    .D(_01574_),
    .Q_N(_14198_),
    .Q(\mem.mem_internal.code_mem[33][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[33][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2813),
    .D(_01575_),
    .Q_N(_14197_),
    .Q(\mem.mem_internal.code_mem[33][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[33][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2814),
    .D(_01576_),
    .Q_N(_14196_),
    .Q(\mem.mem_internal.code_mem[33][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[33][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2815),
    .D(_01577_),
    .Q_N(_14195_),
    .Q(\mem.mem_internal.code_mem[33][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[34][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2816),
    .D(_01578_),
    .Q_N(_14194_),
    .Q(\mem.mem_internal.code_mem[34][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[34][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2817),
    .D(_01579_),
    .Q_N(_14193_),
    .Q(\mem.mem_internal.code_mem[34][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[34][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2818),
    .D(_01580_),
    .Q_N(_14192_),
    .Q(\mem.mem_internal.code_mem[34][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[34][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2819),
    .D(_01581_),
    .Q_N(_14191_),
    .Q(\mem.mem_internal.code_mem[34][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[34][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2820),
    .D(_01582_),
    .Q_N(_14190_),
    .Q(\mem.mem_internal.code_mem[34][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[34][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2821),
    .D(_01583_),
    .Q_N(_14189_),
    .Q(\mem.mem_internal.code_mem[34][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[34][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2822),
    .D(_01584_),
    .Q_N(_14188_),
    .Q(\mem.mem_internal.code_mem[34][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[34][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2823),
    .D(_01585_),
    .Q_N(_14187_),
    .Q(\mem.mem_internal.code_mem[34][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[35][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2824),
    .D(_01586_),
    .Q_N(_14186_),
    .Q(\mem.mem_internal.code_mem[35][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[35][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2825),
    .D(_01587_),
    .Q_N(_14185_),
    .Q(\mem.mem_internal.code_mem[35][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[35][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2826),
    .D(_01588_),
    .Q_N(_14184_),
    .Q(\mem.mem_internal.code_mem[35][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[35][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2827),
    .D(_01589_),
    .Q_N(_14183_),
    .Q(\mem.mem_internal.code_mem[35][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[35][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2828),
    .D(_01590_),
    .Q_N(_14182_),
    .Q(\mem.mem_internal.code_mem[35][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[35][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2829),
    .D(_01591_),
    .Q_N(_14181_),
    .Q(\mem.mem_internal.code_mem[35][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[35][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2830),
    .D(_01592_),
    .Q_N(_14180_),
    .Q(\mem.mem_internal.code_mem[35][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[35][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2831),
    .D(_01593_),
    .Q_N(_14179_),
    .Q(\mem.mem_internal.code_mem[35][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[36][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2832),
    .D(_01594_),
    .Q_N(_14178_),
    .Q(\mem.mem_internal.code_mem[36][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[36][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2833),
    .D(_01595_),
    .Q_N(_14177_),
    .Q(\mem.mem_internal.code_mem[36][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[36][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2834),
    .D(_01596_),
    .Q_N(_14176_),
    .Q(\mem.mem_internal.code_mem[36][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[36][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2835),
    .D(_01597_),
    .Q_N(_14175_),
    .Q(\mem.mem_internal.code_mem[36][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[36][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2836),
    .D(_01598_),
    .Q_N(_14174_),
    .Q(\mem.mem_internal.code_mem[36][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[36][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2837),
    .D(_01599_),
    .Q_N(_14173_),
    .Q(\mem.mem_internal.code_mem[36][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[36][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2838),
    .D(_01600_),
    .Q_N(_14172_),
    .Q(\mem.mem_internal.code_mem[36][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[36][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2839),
    .D(_01601_),
    .Q_N(_14171_),
    .Q(\mem.mem_internal.code_mem[36][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[37][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2840),
    .D(_01602_),
    .Q_N(_14170_),
    .Q(\mem.mem_internal.code_mem[37][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[37][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2841),
    .D(_01603_),
    .Q_N(_14169_),
    .Q(\mem.mem_internal.code_mem[37][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[37][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2842),
    .D(_01604_),
    .Q_N(_14168_),
    .Q(\mem.mem_internal.code_mem[37][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[37][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2843),
    .D(_01605_),
    .Q_N(_14167_),
    .Q(\mem.mem_internal.code_mem[37][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[37][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2844),
    .D(_01606_),
    .Q_N(_14166_),
    .Q(\mem.mem_internal.code_mem[37][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[37][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2845),
    .D(_01607_),
    .Q_N(_14165_),
    .Q(\mem.mem_internal.code_mem[37][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[37][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2846),
    .D(_01608_),
    .Q_N(_14164_),
    .Q(\mem.mem_internal.code_mem[37][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[37][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2847),
    .D(_01609_),
    .Q_N(_14163_),
    .Q(\mem.mem_internal.code_mem[37][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[38][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2848),
    .D(_01610_),
    .Q_N(_14162_),
    .Q(\mem.mem_internal.code_mem[38][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[38][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2849),
    .D(_01611_),
    .Q_N(_14161_),
    .Q(\mem.mem_internal.code_mem[38][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[38][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2850),
    .D(_01612_),
    .Q_N(_14160_),
    .Q(\mem.mem_internal.code_mem[38][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[38][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2851),
    .D(_01613_),
    .Q_N(_14159_),
    .Q(\mem.mem_internal.code_mem[38][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[38][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2852),
    .D(_01614_),
    .Q_N(_14158_),
    .Q(\mem.mem_internal.code_mem[38][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[38][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2853),
    .D(_01615_),
    .Q_N(_14157_),
    .Q(\mem.mem_internal.code_mem[38][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[38][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2854),
    .D(_01616_),
    .Q_N(_14156_),
    .Q(\mem.mem_internal.code_mem[38][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[38][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2855),
    .D(_01617_),
    .Q_N(_14155_),
    .Q(\mem.mem_internal.code_mem[38][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[39][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2856),
    .D(_01618_),
    .Q_N(_14154_),
    .Q(\mem.mem_internal.code_mem[39][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[39][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2857),
    .D(_01619_),
    .Q_N(_14153_),
    .Q(\mem.mem_internal.code_mem[39][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[39][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2858),
    .D(_01620_),
    .Q_N(_14152_),
    .Q(\mem.mem_internal.code_mem[39][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[39][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2859),
    .D(_01621_),
    .Q_N(_14151_),
    .Q(\mem.mem_internal.code_mem[39][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[39][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2860),
    .D(_01622_),
    .Q_N(_14150_),
    .Q(\mem.mem_internal.code_mem[39][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[39][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2861),
    .D(_01623_),
    .Q_N(_14149_),
    .Q(\mem.mem_internal.code_mem[39][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[39][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2862),
    .D(_01624_),
    .Q_N(_14148_),
    .Q(\mem.mem_internal.code_mem[39][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[39][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2863),
    .D(_01625_),
    .Q_N(_14147_),
    .Q(\mem.mem_internal.code_mem[39][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[3][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2864),
    .D(_01626_),
    .Q_N(_14146_),
    .Q(\mem.mem_internal.code_mem[3][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[3][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2865),
    .D(_01627_),
    .Q_N(_14145_),
    .Q(\mem.mem_internal.code_mem[3][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[3][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2866),
    .D(_01628_),
    .Q_N(_14144_),
    .Q(\mem.mem_internal.code_mem[3][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[3][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2867),
    .D(_01629_),
    .Q_N(_14143_),
    .Q(\mem.mem_internal.code_mem[3][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[3][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2868),
    .D(_01630_),
    .Q_N(_14142_),
    .Q(\mem.mem_internal.code_mem[3][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[3][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2869),
    .D(_01631_),
    .Q_N(_14141_),
    .Q(\mem.mem_internal.code_mem[3][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[3][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2870),
    .D(_01632_),
    .Q_N(_14140_),
    .Q(\mem.mem_internal.code_mem[3][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[3][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2871),
    .D(_01633_),
    .Q_N(_14139_),
    .Q(\mem.mem_internal.code_mem[3][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[40][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2872),
    .D(_01634_),
    .Q_N(_14138_),
    .Q(\mem.mem_internal.code_mem[40][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[40][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2873),
    .D(_01635_),
    .Q_N(_14137_),
    .Q(\mem.mem_internal.code_mem[40][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[40][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2874),
    .D(_01636_),
    .Q_N(_14136_),
    .Q(\mem.mem_internal.code_mem[40][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[40][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2875),
    .D(_01637_),
    .Q_N(_14135_),
    .Q(\mem.mem_internal.code_mem[40][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[40][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2876),
    .D(_01638_),
    .Q_N(_14134_),
    .Q(\mem.mem_internal.code_mem[40][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[40][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2877),
    .D(_01639_),
    .Q_N(_14133_),
    .Q(\mem.mem_internal.code_mem[40][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[40][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2878),
    .D(_01640_),
    .Q_N(_14132_),
    .Q(\mem.mem_internal.code_mem[40][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[40][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2879),
    .D(_01641_),
    .Q_N(_14131_),
    .Q(\mem.mem_internal.code_mem[40][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[41][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2880),
    .D(_01642_),
    .Q_N(_14130_),
    .Q(\mem.mem_internal.code_mem[41][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[41][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2881),
    .D(_01643_),
    .Q_N(_14129_),
    .Q(\mem.mem_internal.code_mem[41][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[41][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2882),
    .D(_01644_),
    .Q_N(_14128_),
    .Q(\mem.mem_internal.code_mem[41][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[41][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2883),
    .D(_01645_),
    .Q_N(_14127_),
    .Q(\mem.mem_internal.code_mem[41][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[41][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2884),
    .D(_01646_),
    .Q_N(_14126_),
    .Q(\mem.mem_internal.code_mem[41][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[41][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2885),
    .D(_01647_),
    .Q_N(_14125_),
    .Q(\mem.mem_internal.code_mem[41][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[41][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2886),
    .D(_01648_),
    .Q_N(_14124_),
    .Q(\mem.mem_internal.code_mem[41][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[41][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2887),
    .D(_01649_),
    .Q_N(_14123_),
    .Q(\mem.mem_internal.code_mem[41][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[42][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2888),
    .D(_01650_),
    .Q_N(_14122_),
    .Q(\mem.mem_internal.code_mem[42][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[42][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2889),
    .D(_01651_),
    .Q_N(_14121_),
    .Q(\mem.mem_internal.code_mem[42][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[42][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2890),
    .D(_01652_),
    .Q_N(_14120_),
    .Q(\mem.mem_internal.code_mem[42][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[42][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2891),
    .D(_01653_),
    .Q_N(_14119_),
    .Q(\mem.mem_internal.code_mem[42][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[42][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2892),
    .D(_01654_),
    .Q_N(_14118_),
    .Q(\mem.mem_internal.code_mem[42][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[42][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2893),
    .D(_01655_),
    .Q_N(_14117_),
    .Q(\mem.mem_internal.code_mem[42][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[42][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2894),
    .D(_01656_),
    .Q_N(_14116_),
    .Q(\mem.mem_internal.code_mem[42][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[42][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2895),
    .D(_01657_),
    .Q_N(_14115_),
    .Q(\mem.mem_internal.code_mem[42][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[43][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2896),
    .D(_01658_),
    .Q_N(_14114_),
    .Q(\mem.mem_internal.code_mem[43][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[43][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2897),
    .D(_01659_),
    .Q_N(_14113_),
    .Q(\mem.mem_internal.code_mem[43][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[43][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2898),
    .D(_01660_),
    .Q_N(_14112_),
    .Q(\mem.mem_internal.code_mem[43][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[43][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2899),
    .D(_01661_),
    .Q_N(_14111_),
    .Q(\mem.mem_internal.code_mem[43][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[43][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2900),
    .D(_01662_),
    .Q_N(_14110_),
    .Q(\mem.mem_internal.code_mem[43][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[43][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2901),
    .D(_01663_),
    .Q_N(_14109_),
    .Q(\mem.mem_internal.code_mem[43][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[43][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2902),
    .D(_01664_),
    .Q_N(_14108_),
    .Q(\mem.mem_internal.code_mem[43][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[43][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2903),
    .D(_01665_),
    .Q_N(_14107_),
    .Q(\mem.mem_internal.code_mem[43][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[44][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2904),
    .D(_01666_),
    .Q_N(_14106_),
    .Q(\mem.mem_internal.code_mem[44][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[44][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2905),
    .D(_01667_),
    .Q_N(_14105_),
    .Q(\mem.mem_internal.code_mem[44][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[44][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2906),
    .D(_01668_),
    .Q_N(_14104_),
    .Q(\mem.mem_internal.code_mem[44][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[44][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2907),
    .D(_01669_),
    .Q_N(_14103_),
    .Q(\mem.mem_internal.code_mem[44][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[44][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2908),
    .D(_01670_),
    .Q_N(_14102_),
    .Q(\mem.mem_internal.code_mem[44][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[44][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2909),
    .D(_01671_),
    .Q_N(_14101_),
    .Q(\mem.mem_internal.code_mem[44][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[44][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2910),
    .D(_01672_),
    .Q_N(_14100_),
    .Q(\mem.mem_internal.code_mem[44][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[44][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2911),
    .D(_01673_),
    .Q_N(_14099_),
    .Q(\mem.mem_internal.code_mem[44][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[45][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2912),
    .D(_01674_),
    .Q_N(_14098_),
    .Q(\mem.mem_internal.code_mem[45][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[45][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2913),
    .D(_01675_),
    .Q_N(_14097_),
    .Q(\mem.mem_internal.code_mem[45][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[45][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2914),
    .D(_01676_),
    .Q_N(_14096_),
    .Q(\mem.mem_internal.code_mem[45][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[45][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2915),
    .D(_01677_),
    .Q_N(_14095_),
    .Q(\mem.mem_internal.code_mem[45][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[45][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2916),
    .D(_01678_),
    .Q_N(_14094_),
    .Q(\mem.mem_internal.code_mem[45][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[45][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2917),
    .D(_01679_),
    .Q_N(_14093_),
    .Q(\mem.mem_internal.code_mem[45][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[45][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2918),
    .D(_01680_),
    .Q_N(_14092_),
    .Q(\mem.mem_internal.code_mem[45][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[45][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2919),
    .D(_01681_),
    .Q_N(_14091_),
    .Q(\mem.mem_internal.code_mem[45][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[46][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2920),
    .D(_01682_),
    .Q_N(_14090_),
    .Q(\mem.mem_internal.code_mem[46][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[46][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2921),
    .D(_01683_),
    .Q_N(_14089_),
    .Q(\mem.mem_internal.code_mem[46][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[46][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net2922),
    .D(_01684_),
    .Q_N(_14088_),
    .Q(\mem.mem_internal.code_mem[46][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[46][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2923),
    .D(_01685_),
    .Q_N(_14087_),
    .Q(\mem.mem_internal.code_mem[46][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[46][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2924),
    .D(_01686_),
    .Q_N(_14086_),
    .Q(\mem.mem_internal.code_mem[46][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[46][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2925),
    .D(_01687_),
    .Q_N(_14085_),
    .Q(\mem.mem_internal.code_mem[46][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[46][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2926),
    .D(_01688_),
    .Q_N(_14084_),
    .Q(\mem.mem_internal.code_mem[46][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[46][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2927),
    .D(_01689_),
    .Q_N(_14083_),
    .Q(\mem.mem_internal.code_mem[46][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[47][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2928),
    .D(_01690_),
    .Q_N(_14082_),
    .Q(\mem.mem_internal.code_mem[47][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[47][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2929),
    .D(_01691_),
    .Q_N(_14081_),
    .Q(\mem.mem_internal.code_mem[47][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[47][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2930),
    .D(_01692_),
    .Q_N(_14080_),
    .Q(\mem.mem_internal.code_mem[47][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[47][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2931),
    .D(_01693_),
    .Q_N(_14079_),
    .Q(\mem.mem_internal.code_mem[47][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[47][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2932),
    .D(_01694_),
    .Q_N(_14078_),
    .Q(\mem.mem_internal.code_mem[47][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[47][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2933),
    .D(_01695_),
    .Q_N(_14077_),
    .Q(\mem.mem_internal.code_mem[47][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[47][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2934),
    .D(_01696_),
    .Q_N(_14076_),
    .Q(\mem.mem_internal.code_mem[47][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[47][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2935),
    .D(_01697_),
    .Q_N(_14075_),
    .Q(\mem.mem_internal.code_mem[47][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[48][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2936),
    .D(_01698_),
    .Q_N(_14074_),
    .Q(\mem.mem_internal.code_mem[48][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[48][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2937),
    .D(_01699_),
    .Q_N(_14073_),
    .Q(\mem.mem_internal.code_mem[48][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[48][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2938),
    .D(_01700_),
    .Q_N(_14072_),
    .Q(\mem.mem_internal.code_mem[48][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[48][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2939),
    .D(_01701_),
    .Q_N(_14071_),
    .Q(\mem.mem_internal.code_mem[48][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[48][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2940),
    .D(_01702_),
    .Q_N(_14070_),
    .Q(\mem.mem_internal.code_mem[48][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[48][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2941),
    .D(_01703_),
    .Q_N(_14069_),
    .Q(\mem.mem_internal.code_mem[48][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[48][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2942),
    .D(_01704_),
    .Q_N(_14068_),
    .Q(\mem.mem_internal.code_mem[48][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[48][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2943),
    .D(_01705_),
    .Q_N(_14067_),
    .Q(\mem.mem_internal.code_mem[48][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[49][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2944),
    .D(_01706_),
    .Q_N(_14066_),
    .Q(\mem.mem_internal.code_mem[49][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[49][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2945),
    .D(_01707_),
    .Q_N(_14065_),
    .Q(\mem.mem_internal.code_mem[49][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[49][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2946),
    .D(_01708_),
    .Q_N(_14064_),
    .Q(\mem.mem_internal.code_mem[49][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[49][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2947),
    .D(_01709_),
    .Q_N(_14063_),
    .Q(\mem.mem_internal.code_mem[49][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[49][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2948),
    .D(_01710_),
    .Q_N(_14062_),
    .Q(\mem.mem_internal.code_mem[49][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[49][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2949),
    .D(_01711_),
    .Q_N(_14061_),
    .Q(\mem.mem_internal.code_mem[49][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[49][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2950),
    .D(_01712_),
    .Q_N(_14060_),
    .Q(\mem.mem_internal.code_mem[49][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[49][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2951),
    .D(_01713_),
    .Q_N(_14059_),
    .Q(\mem.mem_internal.code_mem[49][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[4][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2952),
    .D(_01714_),
    .Q_N(_14058_),
    .Q(\mem.mem_internal.code_mem[4][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[4][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2953),
    .D(_01715_),
    .Q_N(_14057_),
    .Q(\mem.mem_internal.code_mem[4][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[4][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2954),
    .D(_01716_),
    .Q_N(_14056_),
    .Q(\mem.mem_internal.code_mem[4][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[4][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2955),
    .D(_01717_),
    .Q_N(_14055_),
    .Q(\mem.mem_internal.code_mem[4][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[4][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2956),
    .D(_01718_),
    .Q_N(_14054_),
    .Q(\mem.mem_internal.code_mem[4][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[4][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2957),
    .D(_01719_),
    .Q_N(_14053_),
    .Q(\mem.mem_internal.code_mem[4][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[4][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2958),
    .D(_01720_),
    .Q_N(_14052_),
    .Q(\mem.mem_internal.code_mem[4][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[4][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2959),
    .D(_01721_),
    .Q_N(_14051_),
    .Q(\mem.mem_internal.code_mem[4][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[50][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2960),
    .D(_01722_),
    .Q_N(_14050_),
    .Q(\mem.mem_internal.code_mem[50][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[50][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2961),
    .D(_01723_),
    .Q_N(_14049_),
    .Q(\mem.mem_internal.code_mem[50][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[50][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2962),
    .D(_01724_),
    .Q_N(_14048_),
    .Q(\mem.mem_internal.code_mem[50][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[50][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2963),
    .D(_01725_),
    .Q_N(_14047_),
    .Q(\mem.mem_internal.code_mem[50][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[50][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2964),
    .D(_01726_),
    .Q_N(_14046_),
    .Q(\mem.mem_internal.code_mem[50][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[50][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2965),
    .D(_01727_),
    .Q_N(_14045_),
    .Q(\mem.mem_internal.code_mem[50][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[50][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2966),
    .D(_01728_),
    .Q_N(_14044_),
    .Q(\mem.mem_internal.code_mem[50][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[50][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2967),
    .D(_01729_),
    .Q_N(_14043_),
    .Q(\mem.mem_internal.code_mem[50][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[51][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2968),
    .D(_01730_),
    .Q_N(_14042_),
    .Q(\mem.mem_internal.code_mem[51][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[51][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2969),
    .D(_01731_),
    .Q_N(_14041_),
    .Q(\mem.mem_internal.code_mem[51][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[51][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2970),
    .D(_01732_),
    .Q_N(_14040_),
    .Q(\mem.mem_internal.code_mem[51][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[51][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2971),
    .D(_01733_),
    .Q_N(_14039_),
    .Q(\mem.mem_internal.code_mem[51][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[51][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2972),
    .D(_01734_),
    .Q_N(_14038_),
    .Q(\mem.mem_internal.code_mem[51][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[51][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2973),
    .D(_01735_),
    .Q_N(_14037_),
    .Q(\mem.mem_internal.code_mem[51][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[51][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2974),
    .D(_01736_),
    .Q_N(_14036_),
    .Q(\mem.mem_internal.code_mem[51][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[51][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2975),
    .D(_01737_),
    .Q_N(_14035_),
    .Q(\mem.mem_internal.code_mem[51][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[52][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2976),
    .D(_01738_),
    .Q_N(_14034_),
    .Q(\mem.mem_internal.code_mem[52][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[52][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2977),
    .D(_01739_),
    .Q_N(_14033_),
    .Q(\mem.mem_internal.code_mem[52][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[52][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2978),
    .D(_01740_),
    .Q_N(_14032_),
    .Q(\mem.mem_internal.code_mem[52][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[52][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2979),
    .D(_01741_),
    .Q_N(_14031_),
    .Q(\mem.mem_internal.code_mem[52][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[52][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2980),
    .D(_01742_),
    .Q_N(_14030_),
    .Q(\mem.mem_internal.code_mem[52][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[52][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2981),
    .D(_01743_),
    .Q_N(_14029_),
    .Q(\mem.mem_internal.code_mem[52][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[52][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2982),
    .D(_01744_),
    .Q_N(_14028_),
    .Q(\mem.mem_internal.code_mem[52][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[52][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2983),
    .D(_01745_),
    .Q_N(_14027_),
    .Q(\mem.mem_internal.code_mem[52][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[53][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2984),
    .D(_01746_),
    .Q_N(_14026_),
    .Q(\mem.mem_internal.code_mem[53][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[53][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2985),
    .D(_01747_),
    .Q_N(_14025_),
    .Q(\mem.mem_internal.code_mem[53][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[53][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2986),
    .D(_01748_),
    .Q_N(_14024_),
    .Q(\mem.mem_internal.code_mem[53][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[53][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2987),
    .D(_01749_),
    .Q_N(_14023_),
    .Q(\mem.mem_internal.code_mem[53][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[53][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2988),
    .D(_01750_),
    .Q_N(_14022_),
    .Q(\mem.mem_internal.code_mem[53][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[53][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2989),
    .D(_01751_),
    .Q_N(_14021_),
    .Q(\mem.mem_internal.code_mem[53][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[53][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2990),
    .D(_01752_),
    .Q_N(_14020_),
    .Q(\mem.mem_internal.code_mem[53][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[53][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2991),
    .D(_01753_),
    .Q_N(_14019_),
    .Q(\mem.mem_internal.code_mem[53][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[54][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2992),
    .D(_01754_),
    .Q_N(_14018_),
    .Q(\mem.mem_internal.code_mem[54][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[54][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2993),
    .D(_01755_),
    .Q_N(_14017_),
    .Q(\mem.mem_internal.code_mem[54][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[54][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2994),
    .D(_01756_),
    .Q_N(_14016_),
    .Q(\mem.mem_internal.code_mem[54][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[54][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2995),
    .D(_01757_),
    .Q_N(_14015_),
    .Q(\mem.mem_internal.code_mem[54][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[54][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2996),
    .D(_01758_),
    .Q_N(_14014_),
    .Q(\mem.mem_internal.code_mem[54][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[54][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2997),
    .D(_01759_),
    .Q_N(_14013_),
    .Q(\mem.mem_internal.code_mem[54][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[54][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2998),
    .D(_01760_),
    .Q_N(_14012_),
    .Q(\mem.mem_internal.code_mem[54][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[54][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2999),
    .D(_01761_),
    .Q_N(_14011_),
    .Q(\mem.mem_internal.code_mem[54][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[55][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3000),
    .D(_01762_),
    .Q_N(_14010_),
    .Q(\mem.mem_internal.code_mem[55][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[55][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3001),
    .D(_01763_),
    .Q_N(_14009_),
    .Q(\mem.mem_internal.code_mem[55][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[55][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3002),
    .D(_01764_),
    .Q_N(_14008_),
    .Q(\mem.mem_internal.code_mem[55][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[55][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3003),
    .D(_01765_),
    .Q_N(_14007_),
    .Q(\mem.mem_internal.code_mem[55][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[55][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3004),
    .D(_01766_),
    .Q_N(_14006_),
    .Q(\mem.mem_internal.code_mem[55][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[55][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3005),
    .D(_01767_),
    .Q_N(_14005_),
    .Q(\mem.mem_internal.code_mem[55][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[55][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3006),
    .D(_01768_),
    .Q_N(_14004_),
    .Q(\mem.mem_internal.code_mem[55][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[55][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3007),
    .D(_01769_),
    .Q_N(_14003_),
    .Q(\mem.mem_internal.code_mem[55][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[56][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3008),
    .D(_01770_),
    .Q_N(_14002_),
    .Q(\mem.mem_internal.code_mem[56][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[56][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3009),
    .D(_01771_),
    .Q_N(_14001_),
    .Q(\mem.mem_internal.code_mem[56][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[56][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3010),
    .D(_01772_),
    .Q_N(_14000_),
    .Q(\mem.mem_internal.code_mem[56][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[56][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3011),
    .D(_01773_),
    .Q_N(_13999_),
    .Q(\mem.mem_internal.code_mem[56][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[56][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3012),
    .D(_01774_),
    .Q_N(_13998_),
    .Q(\mem.mem_internal.code_mem[56][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[56][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3013),
    .D(_01775_),
    .Q_N(_13997_),
    .Q(\mem.mem_internal.code_mem[56][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[56][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3014),
    .D(_01776_),
    .Q_N(_13996_),
    .Q(\mem.mem_internal.code_mem[56][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[56][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3015),
    .D(_01777_),
    .Q_N(_13995_),
    .Q(\mem.mem_internal.code_mem[56][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[57][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3016),
    .D(_01778_),
    .Q_N(_13994_),
    .Q(\mem.mem_internal.code_mem[57][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[57][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3017),
    .D(_01779_),
    .Q_N(_13993_),
    .Q(\mem.mem_internal.code_mem[57][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[57][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3018),
    .D(_01780_),
    .Q_N(_13992_),
    .Q(\mem.mem_internal.code_mem[57][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[57][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3019),
    .D(_01781_),
    .Q_N(_13991_),
    .Q(\mem.mem_internal.code_mem[57][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[57][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3020),
    .D(_01782_),
    .Q_N(_13990_),
    .Q(\mem.mem_internal.code_mem[57][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[57][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3021),
    .D(_01783_),
    .Q_N(_13989_),
    .Q(\mem.mem_internal.code_mem[57][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[57][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3022),
    .D(_01784_),
    .Q_N(_13988_),
    .Q(\mem.mem_internal.code_mem[57][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[57][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3023),
    .D(_01785_),
    .Q_N(_13987_),
    .Q(\mem.mem_internal.code_mem[57][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[58][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3024),
    .D(_01786_),
    .Q_N(_13986_),
    .Q(\mem.mem_internal.code_mem[58][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[58][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net3025),
    .D(_01787_),
    .Q_N(_13985_),
    .Q(\mem.mem_internal.code_mem[58][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[58][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3026),
    .D(_01788_),
    .Q_N(_13984_),
    .Q(\mem.mem_internal.code_mem[58][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[58][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3027),
    .D(_01789_),
    .Q_N(_13983_),
    .Q(\mem.mem_internal.code_mem[58][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[58][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3028),
    .D(_01790_),
    .Q_N(_13982_),
    .Q(\mem.mem_internal.code_mem[58][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[58][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3029),
    .D(_01791_),
    .Q_N(_13981_),
    .Q(\mem.mem_internal.code_mem[58][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[58][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3030),
    .D(_01792_),
    .Q_N(_13980_),
    .Q(\mem.mem_internal.code_mem[58][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[58][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3031),
    .D(_01793_),
    .Q_N(_13979_),
    .Q(\mem.mem_internal.code_mem[58][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[59][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3032),
    .D(_01794_),
    .Q_N(_13978_),
    .Q(\mem.mem_internal.code_mem[59][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[59][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net3033),
    .D(_01795_),
    .Q_N(_13977_),
    .Q(\mem.mem_internal.code_mem[59][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[59][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3034),
    .D(_01796_),
    .Q_N(_13976_),
    .Q(\mem.mem_internal.code_mem[59][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[59][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3035),
    .D(_01797_),
    .Q_N(_13975_),
    .Q(\mem.mem_internal.code_mem[59][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[59][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3036),
    .D(_01798_),
    .Q_N(_13974_),
    .Q(\mem.mem_internal.code_mem[59][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[59][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3037),
    .D(_01799_),
    .Q_N(_13973_),
    .Q(\mem.mem_internal.code_mem[59][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[59][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3038),
    .D(_01800_),
    .Q_N(_13972_),
    .Q(\mem.mem_internal.code_mem[59][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[59][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3039),
    .D(_01801_),
    .Q_N(_13971_),
    .Q(\mem.mem_internal.code_mem[59][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[5][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3040),
    .D(_01802_),
    .Q_N(_13970_),
    .Q(\mem.mem_internal.code_mem[5][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[5][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3041),
    .D(_01803_),
    .Q_N(_13969_),
    .Q(\mem.mem_internal.code_mem[5][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[5][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3042),
    .D(_01804_),
    .Q_N(_13968_),
    .Q(\mem.mem_internal.code_mem[5][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[5][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3043),
    .D(_01805_),
    .Q_N(_13967_),
    .Q(\mem.mem_internal.code_mem[5][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[5][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3044),
    .D(_01806_),
    .Q_N(_13966_),
    .Q(\mem.mem_internal.code_mem[5][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[5][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3045),
    .D(_01807_),
    .Q_N(_13965_),
    .Q(\mem.mem_internal.code_mem[5][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[5][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3046),
    .D(_01808_),
    .Q_N(_13964_),
    .Q(\mem.mem_internal.code_mem[5][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[5][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3047),
    .D(_01809_),
    .Q_N(_13963_),
    .Q(\mem.mem_internal.code_mem[5][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[60][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net3048),
    .D(_01810_),
    .Q_N(_13962_),
    .Q(\mem.mem_internal.code_mem[60][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[60][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3049),
    .D(_01811_),
    .Q_N(_13961_),
    .Q(\mem.mem_internal.code_mem[60][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[60][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3050),
    .D(_01812_),
    .Q_N(_13960_),
    .Q(\mem.mem_internal.code_mem[60][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[60][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net3051),
    .D(_01813_),
    .Q_N(_13959_),
    .Q(\mem.mem_internal.code_mem[60][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[60][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3052),
    .D(_01814_),
    .Q_N(_13958_),
    .Q(\mem.mem_internal.code_mem[60][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[60][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3053),
    .D(_01815_),
    .Q_N(_13957_),
    .Q(\mem.mem_internal.code_mem[60][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[60][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3054),
    .D(_01816_),
    .Q_N(_13956_),
    .Q(\mem.mem_internal.code_mem[60][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[60][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net3055),
    .D(_01817_),
    .Q_N(_13955_),
    .Q(\mem.mem_internal.code_mem[60][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[61][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3056),
    .D(_01818_),
    .Q_N(_13954_),
    .Q(\mem.mem_internal.code_mem[61][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[61][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3057),
    .D(_01819_),
    .Q_N(_13953_),
    .Q(\mem.mem_internal.code_mem[61][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[61][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3058),
    .D(_01820_),
    .Q_N(_13952_),
    .Q(\mem.mem_internal.code_mem[61][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[61][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3059),
    .D(_01821_),
    .Q_N(_13951_),
    .Q(\mem.mem_internal.code_mem[61][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[61][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3060),
    .D(_01822_),
    .Q_N(_13950_),
    .Q(\mem.mem_internal.code_mem[61][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[61][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3061),
    .D(_01823_),
    .Q_N(_13949_),
    .Q(\mem.mem_internal.code_mem[61][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[61][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3062),
    .D(_01824_),
    .Q_N(_13948_),
    .Q(\mem.mem_internal.code_mem[61][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[61][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3063),
    .D(_01825_),
    .Q_N(_13947_),
    .Q(\mem.mem_internal.code_mem[61][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[62][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3064),
    .D(_01826_),
    .Q_N(_13946_),
    .Q(\mem.mem_internal.code_mem[62][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[62][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3065),
    .D(_01827_),
    .Q_N(_13945_),
    .Q(\mem.mem_internal.code_mem[62][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[62][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3066),
    .D(_01828_),
    .Q_N(_13944_),
    .Q(\mem.mem_internal.code_mem[62][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[62][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net3067),
    .D(_01829_),
    .Q_N(_13943_),
    .Q(\mem.mem_internal.code_mem[62][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[62][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3068),
    .D(_01830_),
    .Q_N(_13942_),
    .Q(\mem.mem_internal.code_mem[62][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[62][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3069),
    .D(_01831_),
    .Q_N(_13941_),
    .Q(\mem.mem_internal.code_mem[62][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[62][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3070),
    .D(_01832_),
    .Q_N(_13940_),
    .Q(\mem.mem_internal.code_mem[62][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[62][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net3071),
    .D(_01833_),
    .Q_N(_13939_),
    .Q(\mem.mem_internal.code_mem[62][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[63][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net3072),
    .D(_01834_),
    .Q_N(_13938_),
    .Q(\mem.mem_internal.code_mem[63][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[63][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3073),
    .D(_01835_),
    .Q_N(_13937_),
    .Q(\mem.mem_internal.code_mem[63][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[63][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3074),
    .D(_01836_),
    .Q_N(_13936_),
    .Q(\mem.mem_internal.code_mem[63][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[63][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3075),
    .D(_01837_),
    .Q_N(_13935_),
    .Q(\mem.mem_internal.code_mem[63][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[63][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3076),
    .D(_01838_),
    .Q_N(_13934_),
    .Q(\mem.mem_internal.code_mem[63][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[63][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3077),
    .D(_01839_),
    .Q_N(_13933_),
    .Q(\mem.mem_internal.code_mem[63][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[63][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3078),
    .D(_01840_),
    .Q_N(_13932_),
    .Q(\mem.mem_internal.code_mem[63][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[63][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3079),
    .D(_01841_),
    .Q_N(_13931_),
    .Q(\mem.mem_internal.code_mem[63][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[64][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3080),
    .D(_01842_),
    .Q_N(_13930_),
    .Q(\mem.mem_internal.code_mem[64][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[64][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3081),
    .D(_01843_),
    .Q_N(_13929_),
    .Q(\mem.mem_internal.code_mem[64][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[64][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3082),
    .D(_01844_),
    .Q_N(_13928_),
    .Q(\mem.mem_internal.code_mem[64][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[64][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3083),
    .D(_01845_),
    .Q_N(_13927_),
    .Q(\mem.mem_internal.code_mem[64][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[64][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3084),
    .D(_01846_),
    .Q_N(_13926_),
    .Q(\mem.mem_internal.code_mem[64][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[64][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3085),
    .D(_01847_),
    .Q_N(_13925_),
    .Q(\mem.mem_internal.code_mem[64][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[64][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3086),
    .D(_01848_),
    .Q_N(_13924_),
    .Q(\mem.mem_internal.code_mem[64][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[64][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3087),
    .D(_01849_),
    .Q_N(_13923_),
    .Q(\mem.mem_internal.code_mem[64][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[65][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3088),
    .D(_01850_),
    .Q_N(_13922_),
    .Q(\mem.mem_internal.code_mem[65][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[65][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3089),
    .D(_01851_),
    .Q_N(_13921_),
    .Q(\mem.mem_internal.code_mem[65][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[65][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3090),
    .D(_01852_),
    .Q_N(_13920_),
    .Q(\mem.mem_internal.code_mem[65][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[65][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3091),
    .D(_01853_),
    .Q_N(_13919_),
    .Q(\mem.mem_internal.code_mem[65][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[65][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3092),
    .D(_01854_),
    .Q_N(_13918_),
    .Q(\mem.mem_internal.code_mem[65][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[65][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3093),
    .D(_01855_),
    .Q_N(_13917_),
    .Q(\mem.mem_internal.code_mem[65][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[65][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3094),
    .D(_01856_),
    .Q_N(_13916_),
    .Q(\mem.mem_internal.code_mem[65][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[65][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3095),
    .D(_01857_),
    .Q_N(_13915_),
    .Q(\mem.mem_internal.code_mem[65][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[66][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3096),
    .D(_01858_),
    .Q_N(_13914_),
    .Q(\mem.mem_internal.code_mem[66][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[66][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3097),
    .D(_01859_),
    .Q_N(_13913_),
    .Q(\mem.mem_internal.code_mem[66][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[66][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3098),
    .D(_01860_),
    .Q_N(_13912_),
    .Q(\mem.mem_internal.code_mem[66][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[66][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3099),
    .D(_01861_),
    .Q_N(_13911_),
    .Q(\mem.mem_internal.code_mem[66][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[66][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3100),
    .D(_01862_),
    .Q_N(_13910_),
    .Q(\mem.mem_internal.code_mem[66][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[66][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3101),
    .D(_01863_),
    .Q_N(_13909_),
    .Q(\mem.mem_internal.code_mem[66][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[66][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3102),
    .D(_01864_),
    .Q_N(_13908_),
    .Q(\mem.mem_internal.code_mem[66][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[66][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3103),
    .D(_01865_),
    .Q_N(_13907_),
    .Q(\mem.mem_internal.code_mem[66][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[67][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3104),
    .D(_01866_),
    .Q_N(_13906_),
    .Q(\mem.mem_internal.code_mem[67][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[67][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3105),
    .D(_01867_),
    .Q_N(_13905_),
    .Q(\mem.mem_internal.code_mem[67][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[67][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3106),
    .D(_01868_),
    .Q_N(_13904_),
    .Q(\mem.mem_internal.code_mem[67][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[67][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3107),
    .D(_01869_),
    .Q_N(_13903_),
    .Q(\mem.mem_internal.code_mem[67][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[67][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3108),
    .D(_01870_),
    .Q_N(_13902_),
    .Q(\mem.mem_internal.code_mem[67][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[67][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3109),
    .D(_01871_),
    .Q_N(_13901_),
    .Q(\mem.mem_internal.code_mem[67][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[67][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3110),
    .D(_01872_),
    .Q_N(_13900_),
    .Q(\mem.mem_internal.code_mem[67][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[67][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3111),
    .D(_01873_),
    .Q_N(_13899_),
    .Q(\mem.mem_internal.code_mem[67][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[68][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3112),
    .D(_01874_),
    .Q_N(_13898_),
    .Q(\mem.mem_internal.code_mem[68][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[68][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3113),
    .D(_01875_),
    .Q_N(_13897_),
    .Q(\mem.mem_internal.code_mem[68][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[68][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3114),
    .D(_01876_),
    .Q_N(_13896_),
    .Q(\mem.mem_internal.code_mem[68][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[68][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3115),
    .D(_01877_),
    .Q_N(_13895_),
    .Q(\mem.mem_internal.code_mem[68][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[68][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3116),
    .D(_01878_),
    .Q_N(_13894_),
    .Q(\mem.mem_internal.code_mem[68][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[68][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3117),
    .D(_01879_),
    .Q_N(_13893_),
    .Q(\mem.mem_internal.code_mem[68][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[68][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3118),
    .D(_01880_),
    .Q_N(_13892_),
    .Q(\mem.mem_internal.code_mem[68][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[68][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3119),
    .D(_01881_),
    .Q_N(_13891_),
    .Q(\mem.mem_internal.code_mem[68][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[69][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3120),
    .D(_01882_),
    .Q_N(_13890_),
    .Q(\mem.mem_internal.code_mem[69][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[69][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3121),
    .D(_01883_),
    .Q_N(_13889_),
    .Q(\mem.mem_internal.code_mem[69][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[69][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3122),
    .D(_01884_),
    .Q_N(_13888_),
    .Q(\mem.mem_internal.code_mem[69][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[69][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3123),
    .D(_01885_),
    .Q_N(_13887_),
    .Q(\mem.mem_internal.code_mem[69][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[69][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3124),
    .D(_01886_),
    .Q_N(_13886_),
    .Q(\mem.mem_internal.code_mem[69][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[69][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3125),
    .D(_01887_),
    .Q_N(_13885_),
    .Q(\mem.mem_internal.code_mem[69][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[69][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3126),
    .D(_01888_),
    .Q_N(_13884_),
    .Q(\mem.mem_internal.code_mem[69][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[69][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3127),
    .D(_01889_),
    .Q_N(_13883_),
    .Q(\mem.mem_internal.code_mem[69][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[6][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3128),
    .D(_01890_),
    .Q_N(_13882_),
    .Q(\mem.mem_internal.code_mem[6][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[6][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3129),
    .D(_01891_),
    .Q_N(_13881_),
    .Q(\mem.mem_internal.code_mem[6][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[6][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3130),
    .D(_01892_),
    .Q_N(_13880_),
    .Q(\mem.mem_internal.code_mem[6][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[6][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3131),
    .D(_01893_),
    .Q_N(_13879_),
    .Q(\mem.mem_internal.code_mem[6][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[6][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3132),
    .D(_01894_),
    .Q_N(_13878_),
    .Q(\mem.mem_internal.code_mem[6][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[6][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3133),
    .D(_01895_),
    .Q_N(_13877_),
    .Q(\mem.mem_internal.code_mem[6][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[6][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3134),
    .D(_01896_),
    .Q_N(_13876_),
    .Q(\mem.mem_internal.code_mem[6][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[6][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3135),
    .D(_01897_),
    .Q_N(_13875_),
    .Q(\mem.mem_internal.code_mem[6][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[70][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3136),
    .D(_01898_),
    .Q_N(_13874_),
    .Q(\mem.mem_internal.code_mem[70][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[70][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3137),
    .D(_01899_),
    .Q_N(_13873_),
    .Q(\mem.mem_internal.code_mem[70][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[70][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3138),
    .D(_01900_),
    .Q_N(_13872_),
    .Q(\mem.mem_internal.code_mem[70][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[70][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3139),
    .D(_01901_),
    .Q_N(_13871_),
    .Q(\mem.mem_internal.code_mem[70][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[70][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3140),
    .D(_01902_),
    .Q_N(_13870_),
    .Q(\mem.mem_internal.code_mem[70][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[70][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3141),
    .D(_01903_),
    .Q_N(_13869_),
    .Q(\mem.mem_internal.code_mem[70][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[70][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3142),
    .D(_01904_),
    .Q_N(_13868_),
    .Q(\mem.mem_internal.code_mem[70][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[70][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3143),
    .D(_01905_),
    .Q_N(_13867_),
    .Q(\mem.mem_internal.code_mem[70][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[71][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3144),
    .D(_01906_),
    .Q_N(_13866_),
    .Q(\mem.mem_internal.code_mem[71][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[71][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3145),
    .D(_01907_),
    .Q_N(_13865_),
    .Q(\mem.mem_internal.code_mem[71][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[71][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3146),
    .D(_01908_),
    .Q_N(_13864_),
    .Q(\mem.mem_internal.code_mem[71][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[71][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3147),
    .D(_01909_),
    .Q_N(_13863_),
    .Q(\mem.mem_internal.code_mem[71][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[71][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3148),
    .D(_01910_),
    .Q_N(_13862_),
    .Q(\mem.mem_internal.code_mem[71][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[71][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3149),
    .D(_01911_),
    .Q_N(_13861_),
    .Q(\mem.mem_internal.code_mem[71][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[71][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3150),
    .D(_01912_),
    .Q_N(_13860_),
    .Q(\mem.mem_internal.code_mem[71][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[71][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3151),
    .D(_01913_),
    .Q_N(_13859_),
    .Q(\mem.mem_internal.code_mem[71][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[72][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3152),
    .D(_01914_),
    .Q_N(_13858_),
    .Q(\mem.mem_internal.code_mem[72][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[72][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3153),
    .D(_01915_),
    .Q_N(_13857_),
    .Q(\mem.mem_internal.code_mem[72][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[72][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3154),
    .D(_01916_),
    .Q_N(_13856_),
    .Q(\mem.mem_internal.code_mem[72][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[72][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3155),
    .D(_01917_),
    .Q_N(_13855_),
    .Q(\mem.mem_internal.code_mem[72][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[72][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3156),
    .D(_01918_),
    .Q_N(_13854_),
    .Q(\mem.mem_internal.code_mem[72][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[72][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3157),
    .D(_01919_),
    .Q_N(_13853_),
    .Q(\mem.mem_internal.code_mem[72][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[72][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3158),
    .D(_01920_),
    .Q_N(_13852_),
    .Q(\mem.mem_internal.code_mem[72][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[72][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3159),
    .D(_01921_),
    .Q_N(_13851_),
    .Q(\mem.mem_internal.code_mem[72][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[73][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3160),
    .D(_01922_),
    .Q_N(_13850_),
    .Q(\mem.mem_internal.code_mem[73][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[73][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3161),
    .D(_01923_),
    .Q_N(_13849_),
    .Q(\mem.mem_internal.code_mem[73][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[73][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3162),
    .D(_01924_),
    .Q_N(_13848_),
    .Q(\mem.mem_internal.code_mem[73][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[73][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3163),
    .D(_01925_),
    .Q_N(_13847_),
    .Q(\mem.mem_internal.code_mem[73][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[73][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3164),
    .D(_01926_),
    .Q_N(_13846_),
    .Q(\mem.mem_internal.code_mem[73][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[73][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3165),
    .D(_01927_),
    .Q_N(_13845_),
    .Q(\mem.mem_internal.code_mem[73][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[73][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3166),
    .D(_01928_),
    .Q_N(_13844_),
    .Q(\mem.mem_internal.code_mem[73][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[73][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3167),
    .D(_01929_),
    .Q_N(_13843_),
    .Q(\mem.mem_internal.code_mem[73][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[74][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3168),
    .D(_01930_),
    .Q_N(_13842_),
    .Q(\mem.mem_internal.code_mem[74][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[74][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3169),
    .D(_01931_),
    .Q_N(_13841_),
    .Q(\mem.mem_internal.code_mem[74][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[74][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3170),
    .D(_01932_),
    .Q_N(_13840_),
    .Q(\mem.mem_internal.code_mem[74][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[74][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3171),
    .D(_01933_),
    .Q_N(_13839_),
    .Q(\mem.mem_internal.code_mem[74][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[74][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3172),
    .D(_01934_),
    .Q_N(_13838_),
    .Q(\mem.mem_internal.code_mem[74][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[74][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3173),
    .D(_01935_),
    .Q_N(_13837_),
    .Q(\mem.mem_internal.code_mem[74][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[74][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3174),
    .D(_01936_),
    .Q_N(_13836_),
    .Q(\mem.mem_internal.code_mem[74][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[74][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3175),
    .D(_01937_),
    .Q_N(_13835_),
    .Q(\mem.mem_internal.code_mem[74][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[75][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3176),
    .D(_01938_),
    .Q_N(_13834_),
    .Q(\mem.mem_internal.code_mem[75][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[75][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3177),
    .D(_01939_),
    .Q_N(_13833_),
    .Q(\mem.mem_internal.code_mem[75][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[75][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3178),
    .D(_01940_),
    .Q_N(_13832_),
    .Q(\mem.mem_internal.code_mem[75][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[75][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3179),
    .D(_01941_),
    .Q_N(_13831_),
    .Q(\mem.mem_internal.code_mem[75][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[75][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3180),
    .D(_01942_),
    .Q_N(_13830_),
    .Q(\mem.mem_internal.code_mem[75][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[75][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3181),
    .D(_01943_),
    .Q_N(_13829_),
    .Q(\mem.mem_internal.code_mem[75][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[75][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3182),
    .D(_01944_),
    .Q_N(_13828_),
    .Q(\mem.mem_internal.code_mem[75][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[75][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3183),
    .D(_01945_),
    .Q_N(_13827_),
    .Q(\mem.mem_internal.code_mem[75][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[76][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3184),
    .D(_01946_),
    .Q_N(_13826_),
    .Q(\mem.mem_internal.code_mem[76][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[76][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3185),
    .D(_01947_),
    .Q_N(_13825_),
    .Q(\mem.mem_internal.code_mem[76][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[76][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3186),
    .D(_01948_),
    .Q_N(_13824_),
    .Q(\mem.mem_internal.code_mem[76][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[76][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3187),
    .D(_01949_),
    .Q_N(_13823_),
    .Q(\mem.mem_internal.code_mem[76][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[76][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3188),
    .D(_01950_),
    .Q_N(_13822_),
    .Q(\mem.mem_internal.code_mem[76][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[76][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3189),
    .D(_01951_),
    .Q_N(_13821_),
    .Q(\mem.mem_internal.code_mem[76][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[76][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3190),
    .D(_01952_),
    .Q_N(_13820_),
    .Q(\mem.mem_internal.code_mem[76][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[76][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3191),
    .D(_01953_),
    .Q_N(_13819_),
    .Q(\mem.mem_internal.code_mem[76][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[77][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3192),
    .D(_01954_),
    .Q_N(_13818_),
    .Q(\mem.mem_internal.code_mem[77][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[77][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3193),
    .D(_01955_),
    .Q_N(_13817_),
    .Q(\mem.mem_internal.code_mem[77][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[77][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3194),
    .D(_01956_),
    .Q_N(_13816_),
    .Q(\mem.mem_internal.code_mem[77][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[77][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net3195),
    .D(_01957_),
    .Q_N(_13815_),
    .Q(\mem.mem_internal.code_mem[77][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[77][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3196),
    .D(_01958_),
    .Q_N(_13814_),
    .Q(\mem.mem_internal.code_mem[77][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[77][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3197),
    .D(_01959_),
    .Q_N(_13813_),
    .Q(\mem.mem_internal.code_mem[77][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[77][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3198),
    .D(_01960_),
    .Q_N(_13812_),
    .Q(\mem.mem_internal.code_mem[77][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[77][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3199),
    .D(_01961_),
    .Q_N(_13811_),
    .Q(\mem.mem_internal.code_mem[77][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[78][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3200),
    .D(_01962_),
    .Q_N(_13810_),
    .Q(\mem.mem_internal.code_mem[78][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[78][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3201),
    .D(_01963_),
    .Q_N(_13809_),
    .Q(\mem.mem_internal.code_mem[78][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[78][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3202),
    .D(_01964_),
    .Q_N(_13808_),
    .Q(\mem.mem_internal.code_mem[78][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[78][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net3203),
    .D(_01965_),
    .Q_N(_13807_),
    .Q(\mem.mem_internal.code_mem[78][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[78][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3204),
    .D(_01966_),
    .Q_N(_13806_),
    .Q(\mem.mem_internal.code_mem[78][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[78][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net3205),
    .D(_01967_),
    .Q_N(_13805_),
    .Q(\mem.mem_internal.code_mem[78][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[78][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net3206),
    .D(_01968_),
    .Q_N(_13804_),
    .Q(\mem.mem_internal.code_mem[78][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[78][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3207),
    .D(_01969_),
    .Q_N(_13803_),
    .Q(\mem.mem_internal.code_mem[78][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[79][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3208),
    .D(_01970_),
    .Q_N(_13802_),
    .Q(\mem.mem_internal.code_mem[79][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[79][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3209),
    .D(_01971_),
    .Q_N(_13801_),
    .Q(\mem.mem_internal.code_mem[79][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[79][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3210),
    .D(_01972_),
    .Q_N(_13800_),
    .Q(\mem.mem_internal.code_mem[79][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[79][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net3211),
    .D(_01973_),
    .Q_N(_13799_),
    .Q(\mem.mem_internal.code_mem[79][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[79][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net3212),
    .D(_01974_),
    .Q_N(_13798_),
    .Q(\mem.mem_internal.code_mem[79][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[79][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net3213),
    .D(_01975_),
    .Q_N(_13797_),
    .Q(\mem.mem_internal.code_mem[79][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[79][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3214),
    .D(_01976_),
    .Q_N(_13796_),
    .Q(\mem.mem_internal.code_mem[79][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[79][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3215),
    .D(_01977_),
    .Q_N(_13795_),
    .Q(\mem.mem_internal.code_mem[79][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[7][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3216),
    .D(_01978_),
    .Q_N(_13794_),
    .Q(\mem.mem_internal.code_mem[7][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[7][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3217),
    .D(_01979_),
    .Q_N(_13793_),
    .Q(\mem.mem_internal.code_mem[7][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[7][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3218),
    .D(_01980_),
    .Q_N(_13792_),
    .Q(\mem.mem_internal.code_mem[7][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[7][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3219),
    .D(_01981_),
    .Q_N(_13791_),
    .Q(\mem.mem_internal.code_mem[7][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[7][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3220),
    .D(_01982_),
    .Q_N(_13790_),
    .Q(\mem.mem_internal.code_mem[7][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[7][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3221),
    .D(_01983_),
    .Q_N(_13789_),
    .Q(\mem.mem_internal.code_mem[7][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[7][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3222),
    .D(_01984_),
    .Q_N(_13788_),
    .Q(\mem.mem_internal.code_mem[7][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[7][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3223),
    .D(_01985_),
    .Q_N(_13787_),
    .Q(\mem.mem_internal.code_mem[7][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[80][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3224),
    .D(_01986_),
    .Q_N(_13786_),
    .Q(\mem.mem_internal.code_mem[80][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[80][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3225),
    .D(_01987_),
    .Q_N(_13785_),
    .Q(\mem.mem_internal.code_mem[80][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[80][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3226),
    .D(_01988_),
    .Q_N(_13784_),
    .Q(\mem.mem_internal.code_mem[80][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[80][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3227),
    .D(_01989_),
    .Q_N(_13783_),
    .Q(\mem.mem_internal.code_mem[80][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[80][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3228),
    .D(_01990_),
    .Q_N(_13782_),
    .Q(\mem.mem_internal.code_mem[80][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[80][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3229),
    .D(_01991_),
    .Q_N(_13781_),
    .Q(\mem.mem_internal.code_mem[80][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[80][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3230),
    .D(_01992_),
    .Q_N(_13780_),
    .Q(\mem.mem_internal.code_mem[80][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[80][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3231),
    .D(_01993_),
    .Q_N(_13779_),
    .Q(\mem.mem_internal.code_mem[80][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[81][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3232),
    .D(_01994_),
    .Q_N(_13778_),
    .Q(\mem.mem_internal.code_mem[81][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[81][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3233),
    .D(_01995_),
    .Q_N(_13777_),
    .Q(\mem.mem_internal.code_mem[81][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[81][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3234),
    .D(_01996_),
    .Q_N(_13776_),
    .Q(\mem.mem_internal.code_mem[81][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[81][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3235),
    .D(_01997_),
    .Q_N(_13775_),
    .Q(\mem.mem_internal.code_mem[81][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[81][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3236),
    .D(_01998_),
    .Q_N(_13774_),
    .Q(\mem.mem_internal.code_mem[81][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[81][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3237),
    .D(_01999_),
    .Q_N(_13773_),
    .Q(\mem.mem_internal.code_mem[81][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[81][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3238),
    .D(_02000_),
    .Q_N(_13772_),
    .Q(\mem.mem_internal.code_mem[81][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[81][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3239),
    .D(_02001_),
    .Q_N(_13771_),
    .Q(\mem.mem_internal.code_mem[81][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[82][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3240),
    .D(_02002_),
    .Q_N(_13770_),
    .Q(\mem.mem_internal.code_mem[82][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[82][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3241),
    .D(_02003_),
    .Q_N(_13769_),
    .Q(\mem.mem_internal.code_mem[82][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[82][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3242),
    .D(_02004_),
    .Q_N(_13768_),
    .Q(\mem.mem_internal.code_mem[82][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[82][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3243),
    .D(_02005_),
    .Q_N(_13767_),
    .Q(\mem.mem_internal.code_mem[82][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[82][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3244),
    .D(_02006_),
    .Q_N(_13766_),
    .Q(\mem.mem_internal.code_mem[82][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[82][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3245),
    .D(_02007_),
    .Q_N(_13765_),
    .Q(\mem.mem_internal.code_mem[82][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[82][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3246),
    .D(_02008_),
    .Q_N(_13764_),
    .Q(\mem.mem_internal.code_mem[82][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[82][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3247),
    .D(_02009_),
    .Q_N(_13763_),
    .Q(\mem.mem_internal.code_mem[82][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[83][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3248),
    .D(_02010_),
    .Q_N(_13762_),
    .Q(\mem.mem_internal.code_mem[83][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[83][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3249),
    .D(_02011_),
    .Q_N(_13761_),
    .Q(\mem.mem_internal.code_mem[83][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[83][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3250),
    .D(_02012_),
    .Q_N(_13760_),
    .Q(\mem.mem_internal.code_mem[83][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[83][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3251),
    .D(_02013_),
    .Q_N(_13759_),
    .Q(\mem.mem_internal.code_mem[83][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[83][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3252),
    .D(_02014_),
    .Q_N(_13758_),
    .Q(\mem.mem_internal.code_mem[83][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[83][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3253),
    .D(_02015_),
    .Q_N(_13757_),
    .Q(\mem.mem_internal.code_mem[83][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[83][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3254),
    .D(_02016_),
    .Q_N(_13756_),
    .Q(\mem.mem_internal.code_mem[83][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[83][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3255),
    .D(_02017_),
    .Q_N(_13755_),
    .Q(\mem.mem_internal.code_mem[83][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[84][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3256),
    .D(_02018_),
    .Q_N(_13754_),
    .Q(\mem.mem_internal.code_mem[84][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[84][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3257),
    .D(_02019_),
    .Q_N(_13753_),
    .Q(\mem.mem_internal.code_mem[84][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[84][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3258),
    .D(_02020_),
    .Q_N(_13752_),
    .Q(\mem.mem_internal.code_mem[84][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[84][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net3259),
    .D(_02021_),
    .Q_N(_13751_),
    .Q(\mem.mem_internal.code_mem[84][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[84][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net3260),
    .D(_02022_),
    .Q_N(_13750_),
    .Q(\mem.mem_internal.code_mem[84][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[84][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net3261),
    .D(_02023_),
    .Q_N(_13749_),
    .Q(\mem.mem_internal.code_mem[84][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[84][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3262),
    .D(_02024_),
    .Q_N(_13748_),
    .Q(\mem.mem_internal.code_mem[84][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[84][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3263),
    .D(_02025_),
    .Q_N(_13747_),
    .Q(\mem.mem_internal.code_mem[84][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[85][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3264),
    .D(_02026_),
    .Q_N(_13746_),
    .Q(\mem.mem_internal.code_mem[85][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[85][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3265),
    .D(_02027_),
    .Q_N(_13745_),
    .Q(\mem.mem_internal.code_mem[85][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[85][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3266),
    .D(_02028_),
    .Q_N(_13744_),
    .Q(\mem.mem_internal.code_mem[85][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[85][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net3267),
    .D(_02029_),
    .Q_N(_13743_),
    .Q(\mem.mem_internal.code_mem[85][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[85][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net3268),
    .D(_02030_),
    .Q_N(_13742_),
    .Q(\mem.mem_internal.code_mem[85][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[85][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net3269),
    .D(_02031_),
    .Q_N(_13741_),
    .Q(\mem.mem_internal.code_mem[85][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[85][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3270),
    .D(_02032_),
    .Q_N(_13740_),
    .Q(\mem.mem_internal.code_mem[85][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[85][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3271),
    .D(_02033_),
    .Q_N(_13739_),
    .Q(\mem.mem_internal.code_mem[85][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[86][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3272),
    .D(_02034_),
    .Q_N(_13738_),
    .Q(\mem.mem_internal.code_mem[86][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[86][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3273),
    .D(_02035_),
    .Q_N(_13737_),
    .Q(\mem.mem_internal.code_mem[86][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[86][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3274),
    .D(_02036_),
    .Q_N(_13736_),
    .Q(\mem.mem_internal.code_mem[86][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[86][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3275),
    .D(_02037_),
    .Q_N(_13735_),
    .Q(\mem.mem_internal.code_mem[86][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[86][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3276),
    .D(_02038_),
    .Q_N(_13734_),
    .Q(\mem.mem_internal.code_mem[86][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[86][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net3277),
    .D(_02039_),
    .Q_N(_13733_),
    .Q(\mem.mem_internal.code_mem[86][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[86][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3278),
    .D(_02040_),
    .Q_N(_13732_),
    .Q(\mem.mem_internal.code_mem[86][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[86][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3279),
    .D(_02041_),
    .Q_N(_13731_),
    .Q(\mem.mem_internal.code_mem[86][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[87][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3280),
    .D(_02042_),
    .Q_N(_13730_),
    .Q(\mem.mem_internal.code_mem[87][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[87][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3281),
    .D(_02043_),
    .Q_N(_13729_),
    .Q(\mem.mem_internal.code_mem[87][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[87][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3282),
    .D(_02044_),
    .Q_N(_13728_),
    .Q(\mem.mem_internal.code_mem[87][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[87][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net3283),
    .D(_02045_),
    .Q_N(_13727_),
    .Q(\mem.mem_internal.code_mem[87][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[87][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3284),
    .D(_02046_),
    .Q_N(_13726_),
    .Q(\mem.mem_internal.code_mem[87][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[87][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3285),
    .D(_02047_),
    .Q_N(_13725_),
    .Q(\mem.mem_internal.code_mem[87][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[87][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3286),
    .D(_02048_),
    .Q_N(_13724_),
    .Q(\mem.mem_internal.code_mem[87][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[87][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3287),
    .D(_02049_),
    .Q_N(_13723_),
    .Q(\mem.mem_internal.code_mem[87][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[88][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3288),
    .D(_02050_),
    .Q_N(_13722_),
    .Q(\mem.mem_internal.code_mem[88][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[88][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3289),
    .D(_02051_),
    .Q_N(_13721_),
    .Q(\mem.mem_internal.code_mem[88][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[88][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3290),
    .D(_02052_),
    .Q_N(_13720_),
    .Q(\mem.mem_internal.code_mem[88][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[88][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3291),
    .D(_02053_),
    .Q_N(_13719_),
    .Q(\mem.mem_internal.code_mem[88][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[88][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3292),
    .D(_02054_),
    .Q_N(_13718_),
    .Q(\mem.mem_internal.code_mem[88][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[88][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3293),
    .D(_02055_),
    .Q_N(_13717_),
    .Q(\mem.mem_internal.code_mem[88][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[88][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3294),
    .D(_02056_),
    .Q_N(_13716_),
    .Q(\mem.mem_internal.code_mem[88][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[88][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3295),
    .D(_02057_),
    .Q_N(_13715_),
    .Q(\mem.mem_internal.code_mem[88][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[89][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3296),
    .D(_02058_),
    .Q_N(_13714_),
    .Q(\mem.mem_internal.code_mem[89][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[89][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3297),
    .D(_02059_),
    .Q_N(_13713_),
    .Q(\mem.mem_internal.code_mem[89][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[89][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3298),
    .D(_02060_),
    .Q_N(_13712_),
    .Q(\mem.mem_internal.code_mem[89][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[89][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3299),
    .D(_02061_),
    .Q_N(_13711_),
    .Q(\mem.mem_internal.code_mem[89][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[89][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3300),
    .D(_02062_),
    .Q_N(_13710_),
    .Q(\mem.mem_internal.code_mem[89][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[89][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3301),
    .D(_02063_),
    .Q_N(_13709_),
    .Q(\mem.mem_internal.code_mem[89][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[89][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3302),
    .D(_02064_),
    .Q_N(_13708_),
    .Q(\mem.mem_internal.code_mem[89][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[89][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3303),
    .D(_02065_),
    .Q_N(_13707_),
    .Q(\mem.mem_internal.code_mem[89][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[8][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3304),
    .D(_02066_),
    .Q_N(_13706_),
    .Q(\mem.mem_internal.code_mem[8][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[8][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3305),
    .D(_02067_),
    .Q_N(_13705_),
    .Q(\mem.mem_internal.code_mem[8][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[8][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3306),
    .D(_02068_),
    .Q_N(_13704_),
    .Q(\mem.mem_internal.code_mem[8][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[8][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3307),
    .D(_02069_),
    .Q_N(_13703_),
    .Q(\mem.mem_internal.code_mem[8][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[8][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3308),
    .D(_02070_),
    .Q_N(_13702_),
    .Q(\mem.mem_internal.code_mem[8][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[8][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3309),
    .D(_02071_),
    .Q_N(_13701_),
    .Q(\mem.mem_internal.code_mem[8][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[8][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3310),
    .D(_02072_),
    .Q_N(_13700_),
    .Q(\mem.mem_internal.code_mem[8][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[8][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3311),
    .D(_02073_),
    .Q_N(_13699_),
    .Q(\mem.mem_internal.code_mem[8][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[90][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3312),
    .D(_02074_),
    .Q_N(_13698_),
    .Q(\mem.mem_internal.code_mem[90][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[90][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3313),
    .D(_02075_),
    .Q_N(_13697_),
    .Q(\mem.mem_internal.code_mem[90][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[90][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3314),
    .D(_02076_),
    .Q_N(_13696_),
    .Q(\mem.mem_internal.code_mem[90][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[90][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3315),
    .D(_02077_),
    .Q_N(_13695_),
    .Q(\mem.mem_internal.code_mem[90][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[90][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3316),
    .D(_02078_),
    .Q_N(_13694_),
    .Q(\mem.mem_internal.code_mem[90][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[90][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3317),
    .D(_02079_),
    .Q_N(_13693_),
    .Q(\mem.mem_internal.code_mem[90][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[90][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3318),
    .D(_02080_),
    .Q_N(_13692_),
    .Q(\mem.mem_internal.code_mem[90][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[90][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3319),
    .D(_02081_),
    .Q_N(_13691_),
    .Q(\mem.mem_internal.code_mem[90][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[91][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3320),
    .D(_02082_),
    .Q_N(_13690_),
    .Q(\mem.mem_internal.code_mem[91][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[91][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3321),
    .D(_02083_),
    .Q_N(_13689_),
    .Q(\mem.mem_internal.code_mem[91][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[91][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3322),
    .D(_02084_),
    .Q_N(_13688_),
    .Q(\mem.mem_internal.code_mem[91][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[91][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3323),
    .D(_02085_),
    .Q_N(_13687_),
    .Q(\mem.mem_internal.code_mem[91][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[91][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3324),
    .D(_02086_),
    .Q_N(_13686_),
    .Q(\mem.mem_internal.code_mem[91][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[91][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3325),
    .D(_02087_),
    .Q_N(_13685_),
    .Q(\mem.mem_internal.code_mem[91][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[91][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3326),
    .D(_02088_),
    .Q_N(_13684_),
    .Q(\mem.mem_internal.code_mem[91][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[91][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3327),
    .D(_02089_),
    .Q_N(_13683_),
    .Q(\mem.mem_internal.code_mem[91][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[92][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3328),
    .D(_02090_),
    .Q_N(_13682_),
    .Q(\mem.mem_internal.code_mem[92][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[92][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3329),
    .D(_02091_),
    .Q_N(_13681_),
    .Q(\mem.mem_internal.code_mem[92][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[92][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3330),
    .D(_02092_),
    .Q_N(_13680_),
    .Q(\mem.mem_internal.code_mem[92][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[92][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3331),
    .D(_02093_),
    .Q_N(_13679_),
    .Q(\mem.mem_internal.code_mem[92][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[92][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3332),
    .D(_02094_),
    .Q_N(_13678_),
    .Q(\mem.mem_internal.code_mem[92][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[92][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3333),
    .D(_02095_),
    .Q_N(_13677_),
    .Q(\mem.mem_internal.code_mem[92][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[92][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3334),
    .D(_02096_),
    .Q_N(_13676_),
    .Q(\mem.mem_internal.code_mem[92][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[92][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3335),
    .D(_02097_),
    .Q_N(_13675_),
    .Q(\mem.mem_internal.code_mem[92][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[93][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3336),
    .D(_02098_),
    .Q_N(_13674_),
    .Q(\mem.mem_internal.code_mem[93][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[93][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3337),
    .D(_02099_),
    .Q_N(_13673_),
    .Q(\mem.mem_internal.code_mem[93][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[93][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3338),
    .D(_02100_),
    .Q_N(_13672_),
    .Q(\mem.mem_internal.code_mem[93][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[93][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3339),
    .D(_02101_),
    .Q_N(_13671_),
    .Q(\mem.mem_internal.code_mem[93][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[93][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3340),
    .D(_02102_),
    .Q_N(_13670_),
    .Q(\mem.mem_internal.code_mem[93][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[93][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3341),
    .D(_02103_),
    .Q_N(_13669_),
    .Q(\mem.mem_internal.code_mem[93][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[93][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3342),
    .D(_02104_),
    .Q_N(_13668_),
    .Q(\mem.mem_internal.code_mem[93][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[93][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3343),
    .D(_02105_),
    .Q_N(_13667_),
    .Q(\mem.mem_internal.code_mem[93][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[94][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3344),
    .D(_02106_),
    .Q_N(_13666_),
    .Q(\mem.mem_internal.code_mem[94][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[94][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3345),
    .D(_02107_),
    .Q_N(_13665_),
    .Q(\mem.mem_internal.code_mem[94][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[94][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3346),
    .D(_02108_),
    .Q_N(_13664_),
    .Q(\mem.mem_internal.code_mem[94][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[94][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3347),
    .D(_02109_),
    .Q_N(_13663_),
    .Q(\mem.mem_internal.code_mem[94][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[94][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3348),
    .D(_02110_),
    .Q_N(_13662_),
    .Q(\mem.mem_internal.code_mem[94][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[94][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3349),
    .D(_02111_),
    .Q_N(_13661_),
    .Q(\mem.mem_internal.code_mem[94][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[94][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3350),
    .D(_02112_),
    .Q_N(_13660_),
    .Q(\mem.mem_internal.code_mem[94][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[94][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3351),
    .D(_02113_),
    .Q_N(_13659_),
    .Q(\mem.mem_internal.code_mem[94][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[95][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3352),
    .D(_02114_),
    .Q_N(_13658_),
    .Q(\mem.mem_internal.code_mem[95][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[95][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3353),
    .D(_02115_),
    .Q_N(_13657_),
    .Q(\mem.mem_internal.code_mem[95][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[95][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3354),
    .D(_02116_),
    .Q_N(_13656_),
    .Q(\mem.mem_internal.code_mem[95][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[95][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3355),
    .D(_02117_),
    .Q_N(_13655_),
    .Q(\mem.mem_internal.code_mem[95][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[95][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3356),
    .D(_02118_),
    .Q_N(_13654_),
    .Q(\mem.mem_internal.code_mem[95][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[95][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3357),
    .D(_02119_),
    .Q_N(_13653_),
    .Q(\mem.mem_internal.code_mem[95][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[95][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3358),
    .D(_02120_),
    .Q_N(_13652_),
    .Q(\mem.mem_internal.code_mem[95][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[95][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3359),
    .D(_02121_),
    .Q_N(_13651_),
    .Q(\mem.mem_internal.code_mem[95][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[96][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3360),
    .D(_02122_),
    .Q_N(_13650_),
    .Q(\mem.mem_internal.code_mem[96][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[96][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3361),
    .D(_02123_),
    .Q_N(_13649_),
    .Q(\mem.mem_internal.code_mem[96][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[96][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3362),
    .D(_02124_),
    .Q_N(_13648_),
    .Q(\mem.mem_internal.code_mem[96][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[96][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3363),
    .D(_02125_),
    .Q_N(_13647_),
    .Q(\mem.mem_internal.code_mem[96][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[96][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3364),
    .D(_02126_),
    .Q_N(_13646_),
    .Q(\mem.mem_internal.code_mem[96][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[96][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3365),
    .D(_02127_),
    .Q_N(_13645_),
    .Q(\mem.mem_internal.code_mem[96][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[96][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3366),
    .D(_02128_),
    .Q_N(_13644_),
    .Q(\mem.mem_internal.code_mem[96][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[96][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3367),
    .D(_02129_),
    .Q_N(_13643_),
    .Q(\mem.mem_internal.code_mem[96][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[97][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3368),
    .D(_02130_),
    .Q_N(_13642_),
    .Q(\mem.mem_internal.code_mem[97][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[97][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3369),
    .D(_02131_),
    .Q_N(_13641_),
    .Q(\mem.mem_internal.code_mem[97][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[97][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3370),
    .D(_02132_),
    .Q_N(_13640_),
    .Q(\mem.mem_internal.code_mem[97][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[97][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3371),
    .D(_02133_),
    .Q_N(_13639_),
    .Q(\mem.mem_internal.code_mem[97][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[97][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3372),
    .D(_02134_),
    .Q_N(_13638_),
    .Q(\mem.mem_internal.code_mem[97][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[97][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3373),
    .D(_02135_),
    .Q_N(_13637_),
    .Q(\mem.mem_internal.code_mem[97][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[97][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3374),
    .D(_02136_),
    .Q_N(_13636_),
    .Q(\mem.mem_internal.code_mem[97][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[97][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3375),
    .D(_02137_),
    .Q_N(_13635_),
    .Q(\mem.mem_internal.code_mem[97][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[98][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3376),
    .D(_02138_),
    .Q_N(_13634_),
    .Q(\mem.mem_internal.code_mem[98][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[98][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3377),
    .D(_02139_),
    .Q_N(_13633_),
    .Q(\mem.mem_internal.code_mem[98][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[98][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3378),
    .D(_02140_),
    .Q_N(_13632_),
    .Q(\mem.mem_internal.code_mem[98][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[98][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3379),
    .D(_02141_),
    .Q_N(_13631_),
    .Q(\mem.mem_internal.code_mem[98][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[98][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3380),
    .D(_02142_),
    .Q_N(_13630_),
    .Q(\mem.mem_internal.code_mem[98][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[98][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3381),
    .D(_02143_),
    .Q_N(_13629_),
    .Q(\mem.mem_internal.code_mem[98][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[98][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3382),
    .D(_02144_),
    .Q_N(_13628_),
    .Q(\mem.mem_internal.code_mem[98][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[98][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3383),
    .D(_02145_),
    .Q_N(_13627_),
    .Q(\mem.mem_internal.code_mem[98][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[99][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3384),
    .D(_02146_),
    .Q_N(_13626_),
    .Q(\mem.mem_internal.code_mem[99][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[99][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3385),
    .D(_02147_),
    .Q_N(_13625_),
    .Q(\mem.mem_internal.code_mem[99][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[99][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3386),
    .D(_02148_),
    .Q_N(_13624_),
    .Q(\mem.mem_internal.code_mem[99][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[99][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3387),
    .D(_02149_),
    .Q_N(_13623_),
    .Q(\mem.mem_internal.code_mem[99][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[99][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3388),
    .D(_02150_),
    .Q_N(_13622_),
    .Q(\mem.mem_internal.code_mem[99][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[99][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3389),
    .D(_02151_),
    .Q_N(_13621_),
    .Q(\mem.mem_internal.code_mem[99][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[99][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3390),
    .D(_02152_),
    .Q_N(_13620_),
    .Q(\mem.mem_internal.code_mem[99][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[99][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3391),
    .D(_02153_),
    .Q_N(_13619_),
    .Q(\mem.mem_internal.code_mem[99][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[9][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3392),
    .D(_02154_),
    .Q_N(_13618_),
    .Q(\mem.mem_internal.code_mem[9][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[9][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3393),
    .D(_02155_),
    .Q_N(_13617_),
    .Q(\mem.mem_internal.code_mem[9][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[9][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3394),
    .D(_02156_),
    .Q_N(_13616_),
    .Q(\mem.mem_internal.code_mem[9][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[9][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net3395),
    .D(_02157_),
    .Q_N(_13615_),
    .Q(\mem.mem_internal.code_mem[9][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[9][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net3396),
    .D(_02158_),
    .Q_N(_13614_),
    .Q(\mem.mem_internal.code_mem[9][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[9][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net3397),
    .D(_02159_),
    .Q_N(_13613_),
    .Q(\mem.mem_internal.code_mem[9][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[9][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net3398),
    .D(_02160_),
    .Q_N(_13612_),
    .Q(\mem.mem_internal.code_mem[9][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.code_mem[9][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3399),
    .D(_02161_),
    .Q_N(_13611_),
    .Q(\mem.mem_internal.code_mem[9][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.cycles[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3400),
    .D(_02162_),
    .Q_N(_00081_),
    .Q(\mem.mem_internal.cycles[0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.cycles[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3401),
    .D(_02163_),
    .Q_N(_13610_),
    .Q(\mem.mem_internal.cycles[1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3402),
    .D(_02164_),
    .Q_N(_13609_),
    .Q(\mem.mem_internal.data_mem[0][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3403),
    .D(_02165_),
    .Q_N(_13608_),
    .Q(\mem.mem_internal.data_mem[0][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[0][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3404),
    .D(_02166_),
    .Q_N(_13607_),
    .Q(\mem.mem_internal.data_mem[0][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3405),
    .D(_02167_),
    .Q_N(_13606_),
    .Q(\mem.mem_internal.data_mem[0][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[0][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3406),
    .D(_02168_),
    .Q_N(_13605_),
    .Q(\mem.mem_internal.data_mem[0][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[0][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3407),
    .D(_02169_),
    .Q_N(_13604_),
    .Q(\mem.mem_internal.data_mem[0][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[0][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3408),
    .D(_02170_),
    .Q_N(_13603_),
    .Q(\mem.mem_internal.data_mem[0][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[0][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3409),
    .D(_02171_),
    .Q_N(_13602_),
    .Q(\mem.mem_internal.data_mem[0][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[10][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net3410),
    .D(_02172_),
    .Q_N(_13601_),
    .Q(\mem.mem_internal.data_mem[10][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[10][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net3411),
    .D(_02173_),
    .Q_N(_13600_),
    .Q(\mem.mem_internal.data_mem[10][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[10][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3412),
    .D(_02174_),
    .Q_N(_13599_),
    .Q(\mem.mem_internal.data_mem[10][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[10][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3413),
    .D(_02175_),
    .Q_N(_13598_),
    .Q(\mem.mem_internal.data_mem[10][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[10][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3414),
    .D(_02176_),
    .Q_N(_13597_),
    .Q(\mem.mem_internal.data_mem[10][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[10][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3415),
    .D(_02177_),
    .Q_N(_13596_),
    .Q(\mem.mem_internal.data_mem[10][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[10][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3416),
    .D(_02178_),
    .Q_N(_13595_),
    .Q(\mem.mem_internal.data_mem[10][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[10][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3417),
    .D(_02179_),
    .Q_N(_13594_),
    .Q(\mem.mem_internal.data_mem[10][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[11][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3418),
    .D(_02180_),
    .Q_N(_13593_),
    .Q(\mem.mem_internal.data_mem[11][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[11][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net3419),
    .D(_02181_),
    .Q_N(_13592_),
    .Q(\mem.mem_internal.data_mem[11][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[11][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3420),
    .D(_02182_),
    .Q_N(_13591_),
    .Q(\mem.mem_internal.data_mem[11][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[11][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3421),
    .D(_02183_),
    .Q_N(_13590_),
    .Q(\mem.mem_internal.data_mem[11][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[11][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3422),
    .D(_02184_),
    .Q_N(_13589_),
    .Q(\mem.mem_internal.data_mem[11][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[11][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3423),
    .D(_02185_),
    .Q_N(_13588_),
    .Q(\mem.mem_internal.data_mem[11][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[11][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3424),
    .D(_02186_),
    .Q_N(_13587_),
    .Q(\mem.mem_internal.data_mem[11][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[11][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3425),
    .D(_02187_),
    .Q_N(_13586_),
    .Q(\mem.mem_internal.data_mem[11][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[12][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3426),
    .D(_02188_),
    .Q_N(_13585_),
    .Q(\mem.mem_internal.data_mem[12][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[12][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net3427),
    .D(_02189_),
    .Q_N(_13584_),
    .Q(\mem.mem_internal.data_mem[12][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[12][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3428),
    .D(_02190_),
    .Q_N(_13583_),
    .Q(\mem.mem_internal.data_mem[12][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[12][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net3429),
    .D(_02191_),
    .Q_N(_13582_),
    .Q(\mem.mem_internal.data_mem[12][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[12][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3430),
    .D(_02192_),
    .Q_N(_13581_),
    .Q(\mem.mem_internal.data_mem[12][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[12][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net3431),
    .D(_02193_),
    .Q_N(_13580_),
    .Q(\mem.mem_internal.data_mem[12][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[12][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3432),
    .D(_02194_),
    .Q_N(_13579_),
    .Q(\mem.mem_internal.data_mem[12][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[12][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3433),
    .D(_02195_),
    .Q_N(_13578_),
    .Q(\mem.mem_internal.data_mem[12][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[13][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3434),
    .D(_02196_),
    .Q_N(_13577_),
    .Q(\mem.mem_internal.data_mem[13][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[13][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net3435),
    .D(_02197_),
    .Q_N(_13576_),
    .Q(\mem.mem_internal.data_mem[13][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[13][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3436),
    .D(_02198_),
    .Q_N(_13575_),
    .Q(\mem.mem_internal.data_mem[13][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[13][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net3437),
    .D(_02199_),
    .Q_N(_13574_),
    .Q(\mem.mem_internal.data_mem[13][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[13][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3438),
    .D(_02200_),
    .Q_N(_13573_),
    .Q(\mem.mem_internal.data_mem[13][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[13][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3439),
    .D(_02201_),
    .Q_N(_13572_),
    .Q(\mem.mem_internal.data_mem[13][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[13][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3440),
    .D(_02202_),
    .Q_N(_13571_),
    .Q(\mem.mem_internal.data_mem[13][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[13][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3441),
    .D(_02203_),
    .Q_N(_13570_),
    .Q(\mem.mem_internal.data_mem[13][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[14][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3442),
    .D(_02204_),
    .Q_N(_13569_),
    .Q(\mem.mem_internal.data_mem[14][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[14][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net3443),
    .D(_02205_),
    .Q_N(_13568_),
    .Q(\mem.mem_internal.data_mem[14][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[14][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3444),
    .D(_02206_),
    .Q_N(_13567_),
    .Q(\mem.mem_internal.data_mem[14][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[14][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3445),
    .D(_02207_),
    .Q_N(_13566_),
    .Q(\mem.mem_internal.data_mem[14][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[14][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3446),
    .D(_02208_),
    .Q_N(_13565_),
    .Q(\mem.mem_internal.data_mem[14][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[14][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3447),
    .D(_02209_),
    .Q_N(_13564_),
    .Q(\mem.mem_internal.data_mem[14][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[14][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3448),
    .D(_02210_),
    .Q_N(_13563_),
    .Q(\mem.mem_internal.data_mem[14][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[14][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3449),
    .D(_02211_),
    .Q_N(_13562_),
    .Q(\mem.mem_internal.data_mem[14][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[15][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3450),
    .D(_02212_),
    .Q_N(_13561_),
    .Q(\mem.mem_internal.data_mem[15][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[15][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3451),
    .D(_02213_),
    .Q_N(_13560_),
    .Q(\mem.mem_internal.data_mem[15][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[15][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net3452),
    .D(_02214_),
    .Q_N(_13559_),
    .Q(\mem.mem_internal.data_mem[15][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[15][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3453),
    .D(_02215_),
    .Q_N(_13558_),
    .Q(\mem.mem_internal.data_mem[15][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[15][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3454),
    .D(_02216_),
    .Q_N(_13557_),
    .Q(\mem.mem_internal.data_mem[15][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[15][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3455),
    .D(_02217_),
    .Q_N(_13556_),
    .Q(\mem.mem_internal.data_mem[15][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[15][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3456),
    .D(_02218_),
    .Q_N(_13555_),
    .Q(\mem.mem_internal.data_mem[15][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[15][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3457),
    .D(_02219_),
    .Q_N(_13554_),
    .Q(\mem.mem_internal.data_mem[15][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[16][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3458),
    .D(_02220_),
    .Q_N(_13553_),
    .Q(\mem.mem_internal.data_mem[16][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[16][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3459),
    .D(_02221_),
    .Q_N(_13552_),
    .Q(\mem.mem_internal.data_mem[16][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[16][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3460),
    .D(_02222_),
    .Q_N(_13551_),
    .Q(\mem.mem_internal.data_mem[16][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[16][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3461),
    .D(_02223_),
    .Q_N(_13550_),
    .Q(\mem.mem_internal.data_mem[16][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[16][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3462),
    .D(_02224_),
    .Q_N(_13549_),
    .Q(\mem.mem_internal.data_mem[16][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[16][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3463),
    .D(_02225_),
    .Q_N(_13548_),
    .Q(\mem.mem_internal.data_mem[16][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[16][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3464),
    .D(_02226_),
    .Q_N(_13547_),
    .Q(\mem.mem_internal.data_mem[16][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[16][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3465),
    .D(_02227_),
    .Q_N(_13546_),
    .Q(\mem.mem_internal.data_mem[16][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[17][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3466),
    .D(_02228_),
    .Q_N(_13545_),
    .Q(\mem.mem_internal.data_mem[17][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[17][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3467),
    .D(_02229_),
    .Q_N(_13544_),
    .Q(\mem.mem_internal.data_mem[17][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[17][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3468),
    .D(_02230_),
    .Q_N(_13543_),
    .Q(\mem.mem_internal.data_mem[17][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[17][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3469),
    .D(_02231_),
    .Q_N(_13542_),
    .Q(\mem.mem_internal.data_mem[17][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[17][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3470),
    .D(_02232_),
    .Q_N(_13541_),
    .Q(\mem.mem_internal.data_mem[17][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[17][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3471),
    .D(_02233_),
    .Q_N(_13540_),
    .Q(\mem.mem_internal.data_mem[17][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[17][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3472),
    .D(_02234_),
    .Q_N(_13539_),
    .Q(\mem.mem_internal.data_mem[17][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[17][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3473),
    .D(_02235_),
    .Q_N(_13538_),
    .Q(\mem.mem_internal.data_mem[17][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[18][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3474),
    .D(_02236_),
    .Q_N(_13537_),
    .Q(\mem.mem_internal.data_mem[18][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[18][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3475),
    .D(_02237_),
    .Q_N(_13536_),
    .Q(\mem.mem_internal.data_mem[18][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[18][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3476),
    .D(_02238_),
    .Q_N(_13535_),
    .Q(\mem.mem_internal.data_mem[18][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[18][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3477),
    .D(_02239_),
    .Q_N(_13534_),
    .Q(\mem.mem_internal.data_mem[18][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[18][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3478),
    .D(_02240_),
    .Q_N(_13533_),
    .Q(\mem.mem_internal.data_mem[18][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[18][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3479),
    .D(_02241_),
    .Q_N(_13532_),
    .Q(\mem.mem_internal.data_mem[18][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[18][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3480),
    .D(_02242_),
    .Q_N(_13531_),
    .Q(\mem.mem_internal.data_mem[18][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[18][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3481),
    .D(_02243_),
    .Q_N(_13530_),
    .Q(\mem.mem_internal.data_mem[18][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[19][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3482),
    .D(_02244_),
    .Q_N(_13529_),
    .Q(\mem.mem_internal.data_mem[19][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[19][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3483),
    .D(_02245_),
    .Q_N(_13528_),
    .Q(\mem.mem_internal.data_mem[19][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[19][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3484),
    .D(_02246_),
    .Q_N(_13527_),
    .Q(\mem.mem_internal.data_mem[19][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[19][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3485),
    .D(_02247_),
    .Q_N(_13526_),
    .Q(\mem.mem_internal.data_mem[19][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[19][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3486),
    .D(_02248_),
    .Q_N(_13525_),
    .Q(\mem.mem_internal.data_mem[19][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[19][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3487),
    .D(_02249_),
    .Q_N(_13524_),
    .Q(\mem.mem_internal.data_mem[19][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[19][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3488),
    .D(_02250_),
    .Q_N(_13523_),
    .Q(\mem.mem_internal.data_mem[19][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[19][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3489),
    .D(_02251_),
    .Q_N(_13522_),
    .Q(\mem.mem_internal.data_mem[19][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3490),
    .D(_02252_),
    .Q_N(_13521_),
    .Q(\mem.mem_internal.data_mem[1][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3491),
    .D(_02253_),
    .Q_N(_13520_),
    .Q(\mem.mem_internal.data_mem[1][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[1][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3492),
    .D(_02254_),
    .Q_N(_13519_),
    .Q(\mem.mem_internal.data_mem[1][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3493),
    .D(_02255_),
    .Q_N(_13518_),
    .Q(\mem.mem_internal.data_mem[1][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[1][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3494),
    .D(_02256_),
    .Q_N(_13517_),
    .Q(\mem.mem_internal.data_mem[1][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[1][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3495),
    .D(_02257_),
    .Q_N(_13516_),
    .Q(\mem.mem_internal.data_mem[1][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[1][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3496),
    .D(_02258_),
    .Q_N(_13515_),
    .Q(\mem.mem_internal.data_mem[1][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[1][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3497),
    .D(_02259_),
    .Q_N(_13514_),
    .Q(\mem.mem_internal.data_mem[1][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[20][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3498),
    .D(_02260_),
    .Q_N(_13513_),
    .Q(\mem.mem_internal.data_mem[20][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[20][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3499),
    .D(_02261_),
    .Q_N(_13512_),
    .Q(\mem.mem_internal.data_mem[20][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[20][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3500),
    .D(_02262_),
    .Q_N(_13511_),
    .Q(\mem.mem_internal.data_mem[20][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[20][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3501),
    .D(_02263_),
    .Q_N(_13510_),
    .Q(\mem.mem_internal.data_mem[20][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[20][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3502),
    .D(_02264_),
    .Q_N(_13509_),
    .Q(\mem.mem_internal.data_mem[20][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[20][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3503),
    .D(_02265_),
    .Q_N(_13508_),
    .Q(\mem.mem_internal.data_mem[20][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[20][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3504),
    .D(_02266_),
    .Q_N(_13507_),
    .Q(\mem.mem_internal.data_mem[20][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[20][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3505),
    .D(_02267_),
    .Q_N(_13506_),
    .Q(\mem.mem_internal.data_mem[20][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[21][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3506),
    .D(_02268_),
    .Q_N(_13505_),
    .Q(\mem.mem_internal.data_mem[21][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[21][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3507),
    .D(_02269_),
    .Q_N(_13504_),
    .Q(\mem.mem_internal.data_mem[21][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[21][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3508),
    .D(_02270_),
    .Q_N(_13503_),
    .Q(\mem.mem_internal.data_mem[21][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[21][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3509),
    .D(_02271_),
    .Q_N(_13502_),
    .Q(\mem.mem_internal.data_mem[21][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[21][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3510),
    .D(_02272_),
    .Q_N(_13501_),
    .Q(\mem.mem_internal.data_mem[21][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[21][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3511),
    .D(_02273_),
    .Q_N(_13500_),
    .Q(\mem.mem_internal.data_mem[21][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[21][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3512),
    .D(_02274_),
    .Q_N(_13499_),
    .Q(\mem.mem_internal.data_mem[21][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[21][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3513),
    .D(_02275_),
    .Q_N(_13498_),
    .Q(\mem.mem_internal.data_mem[21][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[22][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3514),
    .D(_02276_),
    .Q_N(_13497_),
    .Q(\mem.mem_internal.data_mem[22][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[22][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3515),
    .D(_02277_),
    .Q_N(_13496_),
    .Q(\mem.mem_internal.data_mem[22][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[22][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3516),
    .D(_02278_),
    .Q_N(_13495_),
    .Q(\mem.mem_internal.data_mem[22][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[22][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3517),
    .D(_02279_),
    .Q_N(_13494_),
    .Q(\mem.mem_internal.data_mem[22][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[22][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3518),
    .D(_02280_),
    .Q_N(_13493_),
    .Q(\mem.mem_internal.data_mem[22][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[22][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3519),
    .D(_02281_),
    .Q_N(_13492_),
    .Q(\mem.mem_internal.data_mem[22][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[22][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3520),
    .D(_02282_),
    .Q_N(_13491_),
    .Q(\mem.mem_internal.data_mem[22][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[22][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3521),
    .D(_02283_),
    .Q_N(_13490_),
    .Q(\mem.mem_internal.data_mem[22][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[23][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3522),
    .D(_02284_),
    .Q_N(_13489_),
    .Q(\mem.mem_internal.data_mem[23][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[23][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3523),
    .D(_02285_),
    .Q_N(_13488_),
    .Q(\mem.mem_internal.data_mem[23][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[23][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3524),
    .D(_02286_),
    .Q_N(_13487_),
    .Q(\mem.mem_internal.data_mem[23][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[23][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3525),
    .D(_02287_),
    .Q_N(_13486_),
    .Q(\mem.mem_internal.data_mem[23][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[23][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3526),
    .D(_02288_),
    .Q_N(_13485_),
    .Q(\mem.mem_internal.data_mem[23][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[23][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3527),
    .D(_02289_),
    .Q_N(_13484_),
    .Q(\mem.mem_internal.data_mem[23][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[23][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3528),
    .D(_02290_),
    .Q_N(_13483_),
    .Q(\mem.mem_internal.data_mem[23][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[23][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3529),
    .D(_02291_),
    .Q_N(_13482_),
    .Q(\mem.mem_internal.data_mem[23][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[24][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_339_clk),
    .RESET_B(net3530),
    .D(_02292_),
    .Q_N(_13481_),
    .Q(\mem.mem_internal.data_mem[24][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[24][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_339_clk),
    .RESET_B(net3531),
    .D(_02293_),
    .Q_N(_13480_),
    .Q(\mem.mem_internal.data_mem[24][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[24][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3532),
    .D(_02294_),
    .Q_N(_13479_),
    .Q(\mem.mem_internal.data_mem[24][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[24][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3533),
    .D(_02295_),
    .Q_N(_13478_),
    .Q(\mem.mem_internal.data_mem[24][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[24][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3534),
    .D(_02296_),
    .Q_N(_13477_),
    .Q(\mem.mem_internal.data_mem[24][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[24][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3535),
    .D(_02297_),
    .Q_N(_13476_),
    .Q(\mem.mem_internal.data_mem[24][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[24][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3536),
    .D(_02298_),
    .Q_N(_13475_),
    .Q(\mem.mem_internal.data_mem[24][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[24][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3537),
    .D(_02299_),
    .Q_N(_13474_),
    .Q(\mem.mem_internal.data_mem[24][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[25][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_339_clk),
    .RESET_B(net3538),
    .D(_02300_),
    .Q_N(_13473_),
    .Q(\mem.mem_internal.data_mem[25][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[25][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_339_clk),
    .RESET_B(net3539),
    .D(_02301_),
    .Q_N(_13472_),
    .Q(\mem.mem_internal.data_mem[25][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[25][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3540),
    .D(_02302_),
    .Q_N(_13471_),
    .Q(\mem.mem_internal.data_mem[25][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[25][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3541),
    .D(_02303_),
    .Q_N(_13470_),
    .Q(\mem.mem_internal.data_mem[25][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[25][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3542),
    .D(_02304_),
    .Q_N(_13469_),
    .Q(\mem.mem_internal.data_mem[25][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[25][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3543),
    .D(_02305_),
    .Q_N(_13468_),
    .Q(\mem.mem_internal.data_mem[25][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[25][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3544),
    .D(_02306_),
    .Q_N(_13467_),
    .Q(\mem.mem_internal.data_mem[25][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[25][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3545),
    .D(_02307_),
    .Q_N(_13466_),
    .Q(\mem.mem_internal.data_mem[25][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[26][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_339_clk),
    .RESET_B(net3546),
    .D(_02308_),
    .Q_N(_13465_),
    .Q(\mem.mem_internal.data_mem[26][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[26][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_339_clk),
    .RESET_B(net3547),
    .D(_02309_),
    .Q_N(_13464_),
    .Q(\mem.mem_internal.data_mem[26][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[26][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3548),
    .D(_02310_),
    .Q_N(_13463_),
    .Q(\mem.mem_internal.data_mem[26][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[26][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3549),
    .D(_02311_),
    .Q_N(_13462_),
    .Q(\mem.mem_internal.data_mem[26][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[26][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3550),
    .D(_02312_),
    .Q_N(_13461_),
    .Q(\mem.mem_internal.data_mem[26][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[26][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3551),
    .D(_02313_),
    .Q_N(_13460_),
    .Q(\mem.mem_internal.data_mem[26][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[26][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3552),
    .D(_02314_),
    .Q_N(_13459_),
    .Q(\mem.mem_internal.data_mem[26][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[26][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3553),
    .D(_02315_),
    .Q_N(_13458_),
    .Q(\mem.mem_internal.data_mem[26][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[27][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_339_clk),
    .RESET_B(net3554),
    .D(_02316_),
    .Q_N(_13457_),
    .Q(\mem.mem_internal.data_mem[27][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[27][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net3555),
    .D(_02317_),
    .Q_N(_13456_),
    .Q(\mem.mem_internal.data_mem[27][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[27][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3556),
    .D(_02318_),
    .Q_N(_13455_),
    .Q(\mem.mem_internal.data_mem[27][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[27][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3557),
    .D(_02319_),
    .Q_N(_13454_),
    .Q(\mem.mem_internal.data_mem[27][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[27][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3558),
    .D(_02320_),
    .Q_N(_13453_),
    .Q(\mem.mem_internal.data_mem[27][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[27][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3559),
    .D(_02321_),
    .Q_N(_13452_),
    .Q(\mem.mem_internal.data_mem[27][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[27][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3560),
    .D(_02322_),
    .Q_N(_13451_),
    .Q(\mem.mem_internal.data_mem[27][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[27][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3561),
    .D(_02323_),
    .Q_N(_13450_),
    .Q(\mem.mem_internal.data_mem[27][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[28][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3562),
    .D(_02324_),
    .Q_N(_13449_),
    .Q(\mem.mem_internal.data_mem[28][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[28][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3563),
    .D(_02325_),
    .Q_N(_13448_),
    .Q(\mem.mem_internal.data_mem[28][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[28][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_339_clk),
    .RESET_B(net3564),
    .D(_02326_),
    .Q_N(_13447_),
    .Q(\mem.mem_internal.data_mem[28][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[28][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3565),
    .D(_02327_),
    .Q_N(_13446_),
    .Q(\mem.mem_internal.data_mem[28][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[28][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net3566),
    .D(_02328_),
    .Q_N(_13445_),
    .Q(\mem.mem_internal.data_mem[28][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[28][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net3567),
    .D(_02329_),
    .Q_N(_13444_),
    .Q(\mem.mem_internal.data_mem[28][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[28][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3568),
    .D(_02330_),
    .Q_N(_13443_),
    .Q(\mem.mem_internal.data_mem[28][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[28][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3569),
    .D(_02331_),
    .Q_N(_13442_),
    .Q(\mem.mem_internal.data_mem[28][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[29][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3570),
    .D(_02332_),
    .Q_N(_13441_),
    .Q(\mem.mem_internal.data_mem[29][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[29][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3571),
    .D(_02333_),
    .Q_N(_13440_),
    .Q(\mem.mem_internal.data_mem[29][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[29][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net3572),
    .D(_02334_),
    .Q_N(_13439_),
    .Q(\mem.mem_internal.data_mem[29][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[29][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3573),
    .D(_02335_),
    .Q_N(_13438_),
    .Q(\mem.mem_internal.data_mem[29][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[29][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net3574),
    .D(_02336_),
    .Q_N(_13437_),
    .Q(\mem.mem_internal.data_mem[29][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[29][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net3575),
    .D(_02337_),
    .Q_N(_13436_),
    .Q(\mem.mem_internal.data_mem[29][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[29][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3576),
    .D(_02338_),
    .Q_N(_13435_),
    .Q(\mem.mem_internal.data_mem[29][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[29][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3577),
    .D(_02339_),
    .Q_N(_13434_),
    .Q(\mem.mem_internal.data_mem[29][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3578),
    .D(_02340_),
    .Q_N(_13433_),
    .Q(\mem.mem_internal.data_mem[2][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3579),
    .D(_02341_),
    .Q_N(_13432_),
    .Q(\mem.mem_internal.data_mem[2][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[2][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3580),
    .D(_02342_),
    .Q_N(_13431_),
    .Q(\mem.mem_internal.data_mem[2][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3581),
    .D(_02343_),
    .Q_N(_13430_),
    .Q(\mem.mem_internal.data_mem[2][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[2][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3582),
    .D(_02344_),
    .Q_N(_13429_),
    .Q(\mem.mem_internal.data_mem[2][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[2][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3583),
    .D(_02345_),
    .Q_N(_13428_),
    .Q(\mem.mem_internal.data_mem[2][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[2][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3584),
    .D(_02346_),
    .Q_N(_13427_),
    .Q(\mem.mem_internal.data_mem[2][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[2][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3585),
    .D(_02347_),
    .Q_N(_13426_),
    .Q(\mem.mem_internal.data_mem[2][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[30][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3586),
    .D(_02348_),
    .Q_N(_13425_),
    .Q(\mem.mem_internal.data_mem[30][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[30][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3587),
    .D(_02349_),
    .Q_N(_13424_),
    .Q(\mem.mem_internal.data_mem[30][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[30][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net3588),
    .D(_02350_),
    .Q_N(_13423_),
    .Q(\mem.mem_internal.data_mem[30][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[30][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net3589),
    .D(_02351_),
    .Q_N(_13422_),
    .Q(\mem.mem_internal.data_mem[30][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[30][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net3590),
    .D(_02352_),
    .Q_N(_13421_),
    .Q(\mem.mem_internal.data_mem[30][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[30][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net3591),
    .D(_02353_),
    .Q_N(_13420_),
    .Q(\mem.mem_internal.data_mem[30][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[30][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3592),
    .D(_02354_),
    .Q_N(_13419_),
    .Q(\mem.mem_internal.data_mem[30][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[30][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3593),
    .D(_02355_),
    .Q_N(_13418_),
    .Q(\mem.mem_internal.data_mem[30][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[31][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3594),
    .D(_02356_),
    .Q_N(_13417_),
    .Q(\mem.mem_internal.data_mem[31][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[31][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3595),
    .D(_02357_),
    .Q_N(_13416_),
    .Q(\mem.mem_internal.data_mem[31][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[31][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net3596),
    .D(_02358_),
    .Q_N(_13415_),
    .Q(\mem.mem_internal.data_mem[31][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[31][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net3597),
    .D(_02359_),
    .Q_N(_13414_),
    .Q(\mem.mem_internal.data_mem[31][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[31][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net3598),
    .D(_02360_),
    .Q_N(_13413_),
    .Q(\mem.mem_internal.data_mem[31][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[31][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net3599),
    .D(_02361_),
    .Q_N(_13412_),
    .Q(\mem.mem_internal.data_mem[31][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[31][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3600),
    .D(_02362_),
    .Q_N(_13411_),
    .Q(\mem.mem_internal.data_mem[31][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[31][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3601),
    .D(_02363_),
    .Q_N(_13410_),
    .Q(\mem.mem_internal.data_mem[31][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[3][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3602),
    .D(_02364_),
    .Q_N(_13409_),
    .Q(\mem.mem_internal.data_mem[3][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[3][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3603),
    .D(_02365_),
    .Q_N(_13408_),
    .Q(\mem.mem_internal.data_mem[3][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[3][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3604),
    .D(_02366_),
    .Q_N(_13407_),
    .Q(\mem.mem_internal.data_mem[3][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[3][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3605),
    .D(_02367_),
    .Q_N(_13406_),
    .Q(\mem.mem_internal.data_mem[3][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[3][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3606),
    .D(_02368_),
    .Q_N(_13405_),
    .Q(\mem.mem_internal.data_mem[3][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[3][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3607),
    .D(_02369_),
    .Q_N(_13404_),
    .Q(\mem.mem_internal.data_mem[3][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[3][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3608),
    .D(_02370_),
    .Q_N(_13403_),
    .Q(\mem.mem_internal.data_mem[3][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[3][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3609),
    .D(_02371_),
    .Q_N(_13402_),
    .Q(\mem.mem_internal.data_mem[3][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[4][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3610),
    .D(_02372_),
    .Q_N(_13401_),
    .Q(\mem.mem_internal.data_mem[4][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[4][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3611),
    .D(_02373_),
    .Q_N(_13400_),
    .Q(\mem.mem_internal.data_mem[4][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[4][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3612),
    .D(_02374_),
    .Q_N(_13399_),
    .Q(\mem.mem_internal.data_mem[4][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[4][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3613),
    .D(_02375_),
    .Q_N(_13398_),
    .Q(\mem.mem_internal.data_mem[4][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[4][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3614),
    .D(_02376_),
    .Q_N(_13397_),
    .Q(\mem.mem_internal.data_mem[4][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[4][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3615),
    .D(_02377_),
    .Q_N(_13396_),
    .Q(\mem.mem_internal.data_mem[4][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[4][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3616),
    .D(_02378_),
    .Q_N(_13395_),
    .Q(\mem.mem_internal.data_mem[4][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[4][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3617),
    .D(_02379_),
    .Q_N(_13394_),
    .Q(\mem.mem_internal.data_mem[4][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[5][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3618),
    .D(_02380_),
    .Q_N(_13393_),
    .Q(\mem.mem_internal.data_mem[5][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[5][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3619),
    .D(_02381_),
    .Q_N(_13392_),
    .Q(\mem.mem_internal.data_mem[5][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[5][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3620),
    .D(_02382_),
    .Q_N(_13391_),
    .Q(\mem.mem_internal.data_mem[5][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[5][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3621),
    .D(_02383_),
    .Q_N(_13390_),
    .Q(\mem.mem_internal.data_mem[5][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[5][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3622),
    .D(_02384_),
    .Q_N(_13389_),
    .Q(\mem.mem_internal.data_mem[5][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[5][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3623),
    .D(_02385_),
    .Q_N(_13388_),
    .Q(\mem.mem_internal.data_mem[5][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[5][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3624),
    .D(_02386_),
    .Q_N(_13387_),
    .Q(\mem.mem_internal.data_mem[5][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[5][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3625),
    .D(_02387_),
    .Q_N(_13386_),
    .Q(\mem.mem_internal.data_mem[5][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[6][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3626),
    .D(_02388_),
    .Q_N(_13385_),
    .Q(\mem.mem_internal.data_mem[6][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[6][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3627),
    .D(_02389_),
    .Q_N(_13384_),
    .Q(\mem.mem_internal.data_mem[6][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[6][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3628),
    .D(_02390_),
    .Q_N(_13383_),
    .Q(\mem.mem_internal.data_mem[6][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[6][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3629),
    .D(_02391_),
    .Q_N(_13382_),
    .Q(\mem.mem_internal.data_mem[6][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[6][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3630),
    .D(_02392_),
    .Q_N(_13381_),
    .Q(\mem.mem_internal.data_mem[6][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[6][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3631),
    .D(_02393_),
    .Q_N(_13380_),
    .Q(\mem.mem_internal.data_mem[6][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[6][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3632),
    .D(_02394_),
    .Q_N(_13379_),
    .Q(\mem.mem_internal.data_mem[6][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[6][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3633),
    .D(_02395_),
    .Q_N(_13378_),
    .Q(\mem.mem_internal.data_mem[6][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[7][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3634),
    .D(_02396_),
    .Q_N(_13377_),
    .Q(\mem.mem_internal.data_mem[7][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[7][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3635),
    .D(_02397_),
    .Q_N(_13376_),
    .Q(\mem.mem_internal.data_mem[7][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[7][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3636),
    .D(_02398_),
    .Q_N(_13375_),
    .Q(\mem.mem_internal.data_mem[7][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[7][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3637),
    .D(_02399_),
    .Q_N(_13374_),
    .Q(\mem.mem_internal.data_mem[7][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[7][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3638),
    .D(_02400_),
    .Q_N(_13373_),
    .Q(\mem.mem_internal.data_mem[7][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[7][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3639),
    .D(_02401_),
    .Q_N(_13372_),
    .Q(\mem.mem_internal.data_mem[7][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[7][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3640),
    .D(_02402_),
    .Q_N(_13371_),
    .Q(\mem.mem_internal.data_mem[7][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[7][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3641),
    .D(_02403_),
    .Q_N(_13370_),
    .Q(\mem.mem_internal.data_mem[7][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[8][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net3642),
    .D(_02404_),
    .Q_N(_13369_),
    .Q(\mem.mem_internal.data_mem[8][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[8][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net3643),
    .D(_02405_),
    .Q_N(_13368_),
    .Q(\mem.mem_internal.data_mem[8][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[8][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3644),
    .D(_02406_),
    .Q_N(_13367_),
    .Q(\mem.mem_internal.data_mem[8][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[8][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3645),
    .D(_02407_),
    .Q_N(_13366_),
    .Q(\mem.mem_internal.data_mem[8][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[8][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3646),
    .D(_02408_),
    .Q_N(_13365_),
    .Q(\mem.mem_internal.data_mem[8][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[8][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3647),
    .D(_02409_),
    .Q_N(_13364_),
    .Q(\mem.mem_internal.data_mem[8][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[8][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3648),
    .D(_02410_),
    .Q_N(_13363_),
    .Q(\mem.mem_internal.data_mem[8][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[8][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3649),
    .D(_02411_),
    .Q_N(_13362_),
    .Q(\mem.mem_internal.data_mem[8][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[9][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net3650),
    .D(_02412_),
    .Q_N(_13361_),
    .Q(\mem.mem_internal.data_mem[9][0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[9][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net3651),
    .D(_02413_),
    .Q_N(_13360_),
    .Q(\mem.mem_internal.data_mem[9][1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[9][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3652),
    .D(_02414_),
    .Q_N(_13359_),
    .Q(\mem.mem_internal.data_mem[9][2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[9][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3653),
    .D(_02415_),
    .Q_N(_13358_),
    .Q(\mem.mem_internal.data_mem[9][3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[9][4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3654),
    .D(_02416_),
    .Q_N(_13357_),
    .Q(\mem.mem_internal.data_mem[9][4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[9][5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3655),
    .D(_02417_),
    .Q_N(_13356_),
    .Q(\mem.mem_internal.data_mem[9][5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[9][6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net3656),
    .D(_02418_),
    .Q_N(_13355_),
    .Q(\mem.mem_internal.data_mem[9][6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_mem[9][7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3657),
    .D(_02419_),
    .Q_N(_13354_),
    .Q(\mem.mem_internal.data_mem[9][7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3658),
    .D(_02420_),
    .Q_N(_13353_),
    .Q(\mem.internal_data_out[0] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3659),
    .D(_02421_),
    .Q_N(_13352_),
    .Q(\mem.internal_data_out[1] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3660),
    .D(_02422_),
    .Q_N(_13351_),
    .Q(\mem.internal_data_out[2] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3661),
    .D(_02423_),
    .Q_N(_13350_),
    .Q(\mem.internal_data_out[3] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3662),
    .D(_02424_),
    .Q_N(_13349_),
    .Q(\mem.internal_data_out[4] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3663),
    .D(_02425_),
    .Q_N(_13348_),
    .Q(\mem.internal_data_out[5] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3664),
    .D(_02426_),
    .Q_N(_13347_),
    .Q(\mem.internal_data_out[6] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3665),
    .D(_02427_),
    .Q_N(_13346_),
    .Q(\mem.internal_data_out[7] ));
 sg13g2_dfrbp_1 \mem.mem_internal.data_ready$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3666),
    .D(_02428_),
    .Q_N(_13345_),
    .Q(\mem.internal_data_ready ));
 sg13g2_dfrbp_1 \mem.mem_io.data_out[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3667),
    .D(_02429_),
    .Q_N(_13344_),
    .Q(\mem.io_data_out[0] ));
 sg13g2_dfrbp_1 \mem.mem_io.data_out[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3668),
    .D(_02430_),
    .Q_N(_13343_),
    .Q(\mem.io_data_out[1] ));
 sg13g2_dfrbp_1 \mem.mem_io.data_out[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3669),
    .D(_02431_),
    .Q_N(_13342_),
    .Q(\mem.io_data_out[2] ));
 sg13g2_dfrbp_1 \mem.mem_io.data_out[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3670),
    .D(_02432_),
    .Q_N(_13341_),
    .Q(\mem.io_data_out[3] ));
 sg13g2_dfrbp_1 \mem.mem_io.data_out[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3671),
    .D(_02433_),
    .Q_N(_13340_),
    .Q(\mem.io_data_out[4] ));
 sg13g2_dfrbp_1 \mem.mem_io.data_out[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3672),
    .D(_02434_),
    .Q_N(_13339_),
    .Q(\mem.io_data_out[5] ));
 sg13g2_dfrbp_1 \mem.mem_io.data_out[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3673),
    .D(_02435_),
    .Q_N(_13338_),
    .Q(\mem.io_data_out[6] ));
 sg13g2_dfrbp_1 \mem.mem_io.data_out[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3674),
    .D(_02436_),
    .Q_N(_13337_),
    .Q(\mem.io_data_out[7] ));
 sg13g2_dfrbp_1 \mem.mem_io.data_ready$_SDFF_PN0_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3675),
    .D(_02437_),
    .Q_N(_13336_),
    .Q(\mem.io_data_ready ));
 sg13g2_dfrbp_1 \mem.mem_io.past_write$_SDFF_PN0_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3676),
    .D(_02438_),
    .Q_N(_13335_),
    .Q(\mem.mem_io.past_write ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3677),
    .D(_02439_),
    .Q_N(_13334_),
    .Q(\mem.mem_io.porta_oe[0] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net3678),
    .D(_02440_),
    .Q_N(_13333_),
    .Q(\mem.mem_io.porta_oe[1] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_oe[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3679),
    .D(_02441_),
    .Q_N(_13332_),
    .Q(\mem.mem_io.porta_oe[2] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_oe[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3680),
    .D(_02442_),
    .Q_N(_13331_),
    .Q(\mem.mem_io.porta_oe[3] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_oe[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3681),
    .D(_02443_),
    .Q_N(_13330_),
    .Q(\mem.mem_io.porta_oe[4] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_oe[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3682),
    .D(_02444_),
    .Q_N(_13329_),
    .Q(\mem.mem_io.porta_oe[5] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_oe[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3683),
    .D(_02445_),
    .Q_N(_13328_),
    .Q(\mem.mem_io.porta_oe[6] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_oe[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net3684),
    .D(_02446_),
    .Q_N(_13327_),
    .Q(\mem.mem_io.porta_oe[7] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_out[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3685),
    .D(_02447_),
    .Q_N(_13326_),
    .Q(\mem.mem_io.porta_out[0] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_out[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3686),
    .D(_02448_),
    .Q_N(_13325_),
    .Q(\mem.mem_io.porta_out[1] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_out[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3687),
    .D(_02449_),
    .Q_N(_13324_),
    .Q(\mem.mem_io.porta_out[2] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_out[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3688),
    .D(_02450_),
    .Q_N(_13323_),
    .Q(\mem.mem_io.porta_out[3] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_out[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3689),
    .D(_02451_),
    .Q_N(_13322_),
    .Q(\mem.mem_io.porta_out[4] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_out[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3690),
    .D(_02452_),
    .Q_N(_13321_),
    .Q(\mem.mem_io.porta_out[5] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_out[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3691),
    .D(_02453_),
    .Q_N(_13320_),
    .Q(\mem.mem_io.porta_out[6] ));
 sg13g2_dfrbp_1 \mem.mem_io.porta_out[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3692),
    .D(_02454_),
    .Q_N(_13319_),
    .Q(\mem.mem_io.porta_out[7] ));
 sg13g2_dfrbp_1 \mem.mem_io.portb_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3693),
    .D(_02455_),
    .Q_N(_13318_),
    .Q(net13));
 sg13g2_dfrbp_1 \mem.mem_io.portb_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3694),
    .D(_02456_),
    .Q_N(_13317_),
    .Q(net14));
 sg13g2_dfrbp_1 \mem.mem_io.portb_oe[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3695),
    .D(_02457_),
    .Q_N(_13316_),
    .Q(net15));
 sg13g2_dfrbp_1 \mem.mem_io.portb_oe[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3696),
    .D(_02458_),
    .Q_N(_13315_),
    .Q(net16));
 sg13g2_dfrbp_1 \mem.mem_io.portb_oe[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3697),
    .D(_02459_),
    .Q_N(_13314_),
    .Q(net17));
 sg13g2_dfrbp_1 \mem.mem_io.portb_oe[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net3698),
    .D(_02460_),
    .Q_N(_13313_),
    .Q(net18));
 sg13g2_dfrbp_1 \mem.mem_io.portb_oe[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net3699),
    .D(_02461_),
    .Q_N(_13312_),
    .Q(net19));
 sg13g2_dfrbp_1 \mem.mem_io.portb_oe[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net3700),
    .D(_02462_),
    .Q_N(_13311_),
    .Q(net20));
 sg13g2_dfrbp_1 \mem.mem_io.portb_out[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3701),
    .D(_02463_),
    .Q_N(_13310_),
    .Q(net21));
 sg13g2_dfrbp_1 \mem.mem_io.portb_out[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3702),
    .D(_02464_),
    .Q_N(_13309_),
    .Q(net22));
 sg13g2_dfrbp_1 \mem.mem_io.portb_out[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3703),
    .D(_02465_),
    .Q_N(_13308_),
    .Q(net23));
 sg13g2_dfrbp_1 \mem.mem_io.portb_out[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3704),
    .D(_02466_),
    .Q_N(_13307_),
    .Q(net24));
 sg13g2_dfrbp_1 \mem.mem_io.portb_out[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3705),
    .D(_02467_),
    .Q_N(_13306_),
    .Q(net25));
 sg13g2_dfrbp_1 \mem.mem_io.portb_out[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3706),
    .D(_02468_),
    .Q_N(_13305_),
    .Q(net26));
 sg13g2_dfrbp_1 \mem.mem_io.portb_out[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3707),
    .D(_02469_),
    .Q_N(_13304_),
    .Q(net27));
 sg13g2_dfrbp_1 \mem.mem_io.portb_out[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3708),
    .D(_02470_),
    .Q_N(_13303_),
    .Q(net28));
 sg13g2_dfrbp_1 \mem_addr[0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3709),
    .D(_00015_),
    .Q_N(_13302_),
    .Q(\mem.addr[0] ));
 sg13g2_dfrbp_1 \mem_addr[1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3710),
    .D(_00016_),
    .Q_N(_13301_),
    .Q(\mem.addr[1] ));
 sg13g2_dfrbp_1 \mem_addr[2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3711),
    .D(_00017_),
    .Q_N(_00071_),
    .Q(\mem.addr[2] ));
 sg13g2_dfrbp_1 \mem_addr[3]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3712),
    .D(_00018_),
    .Q_N(_13300_),
    .Q(\mem.addr[3] ));
 sg13g2_dfrbp_1 \mem_addr[4]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3713),
    .D(_00019_),
    .Q_N(_13299_),
    .Q(\mem.addr[4] ));
 sg13g2_dfrbp_1 \mem_addr[5]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3714),
    .D(_00020_),
    .Q_N(_13298_),
    .Q(\mem.addr[5] ));
 sg13g2_dfrbp_1 \mem_addr[6]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3715),
    .D(_00021_),
    .Q_N(_13297_),
    .Q(\mem.addr[6] ));
 sg13g2_dfrbp_1 \mem_addr[7]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3716),
    .D(_00022_),
    .Q_N(_13296_),
    .Q(\mem.addr[7] ));
 sg13g2_dfrbp_1 \mem_select$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3717),
    .D(_02471_),
    .Q_N(_13295_),
    .Q(\mem.select ));
 sg13g2_dfrbp_1 \mem_type_data$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3718),
    .D(_02472_),
    .Q_N(_00080_),
    .Q(\mem.mem_internal.memory_type_data ));
 sg13g2_dfrbp_1 \mem_write_en$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3719),
    .D(_02473_),
    .Q_N(_00070_),
    .Q(\mem.mem_internal.write ));
 sg13g2_dfrbp_1 \mem_write_value[0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net3720),
    .D(_02474_),
    .Q_N(_00023_),
    .Q(\mem.data_in[0] ));
 sg13g2_dfrbp_1 \mem_write_value[1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3721),
    .D(_02475_),
    .Q_N(_00024_),
    .Q(\mem.data_in[1] ));
 sg13g2_dfrbp_1 \mem_write_value[2]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3722),
    .D(_02476_),
    .Q_N(_00025_),
    .Q(\mem.data_in[2] ));
 sg13g2_dfrbp_1 \mem_write_value[3]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3723),
    .D(_02477_),
    .Q_N(_00026_),
    .Q(\mem.data_in[3] ));
 sg13g2_dfrbp_1 \mem_write_value[4]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3724),
    .D(_02478_),
    .Q_N(_00027_),
    .Q(\mem.data_in[4] ));
 sg13g2_dfrbp_1 \mem_write_value[5]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3725),
    .D(_02479_),
    .Q_N(_00028_),
    .Q(\mem.data_in[5] ));
 sg13g2_dfrbp_1 \mem_write_value[6]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3726),
    .D(_02480_),
    .Q_N(_00029_),
    .Q(\mem.data_in[6] ));
 sg13g2_dfrbp_1 \mem_write_value[7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3727),
    .D(_02481_),
    .Q_N(_00030_),
    .Q(\mem.data_in[7] ));
 sg13g2_dfrbp_1 \memory_input[0]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3728),
    .D(_02482_),
    .Q_N(_13294_),
    .Q(\exec.memory_input[0] ));
 sg13g2_dfrbp_1 \memory_input[1]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3729),
    .D(_02483_),
    .Q_N(_13293_),
    .Q(\exec.memory_input[1] ));
 sg13g2_dfrbp_1 \memory_input[2]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net3730),
    .D(_02484_),
    .Q_N(_13292_),
    .Q(\exec.memory_input[2] ));
 sg13g2_dfrbp_1 \memory_input[3]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3731),
    .D(_02485_),
    .Q_N(_13291_),
    .Q(\exec.memory_input[3] ));
 sg13g2_dfrbp_1 \memory_input[4]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net3732),
    .D(_02486_),
    .Q_N(_13290_),
    .Q(\exec.memory_input[4] ));
 sg13g2_dfrbp_1 \memory_input[5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3733),
    .D(_02487_),
    .Q_N(_13289_),
    .Q(\exec.memory_input[5] ));
 sg13g2_dfrbp_1 \memory_input[6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net3734),
    .D(_02488_),
    .Q_N(_13288_),
    .Q(\exec.memory_input[6] ));
 sg13g2_dfrbp_1 \memory_input[7]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net3735),
    .D(_02489_),
    .Q_N(_13287_),
    .Q(\exec.memory_input[7] ));
 sg13g2_dfrbp_1 \o_shift_out$_SDFF_PN0_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3736),
    .D(_02490_),
    .Q_N(_13286_),
    .Q(o_shift_out));
 sg13g2_dfrbp_1 \opcode[0]$_SDFF_PN0_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3737),
    .D(_02491_),
    .Q_N(_13285_),
    .Q(\exec.opcode[0] ));
 sg13g2_dfrbp_1 \opcode[1]$_SDFF_PN0_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3738),
    .D(_02492_),
    .Q_N(_13284_),
    .Q(\exec.opcode[1] ));
 sg13g2_dfrbp_1 \opcode[2]$_SDFF_PN0_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3739),
    .D(_02493_),
    .Q_N(_13283_),
    .Q(\exec.opcode[2] ));
 sg13g2_dfrbp_1 \opcode[3]$_SDFF_PN0_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3740),
    .D(_02494_),
    .Q_N(_13282_),
    .Q(\exec.opcode[3] ));
 sg13g2_dfrbp_1 \opcode[4]$_SDFF_PN0_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3741),
    .D(_02495_),
    .Q_N(_13281_),
    .Q(\exec.opcode[4] ));
 sg13g2_dfrbp_1 \opcode[5]$_SDFF_PN0_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3742),
    .D(_02496_),
    .Q_N(_13280_),
    .Q(\exec.opcode[5] ));
 sg13g2_dfrbp_1 \opcode[6]$_SDFF_PN0_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3743),
    .D(_02497_),
    .Q_N(_13279_),
    .Q(\exec.opcode[6] ));
 sg13g2_dfrbp_1 \opcode[7]$_SDFF_PN0_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3744),
    .D(_02498_),
    .Q_N(_13278_),
    .Q(\exec.opcode[7] ));
 sg13g2_dfrbp_1 \out_of_order_exec$_SDFFE_PP0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3745),
    .D(_02499_),
    .Q_N(_13277_),
    .Q(\exec.out_of_order_exec ));
 sg13g2_dfrbp_1 \past_i_run$_SDFF_PN0_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net3746),
    .D(_02500_),
    .Q_N(_13276_),
    .Q(past_i_run));
 sg13g2_dfrbp_1 \pc[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3747),
    .D(_02501_),
    .Q_N(_13275_),
    .Q(\exec.pc[0] ));
 sg13g2_dfrbp_1 \pc[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3748),
    .D(_02502_),
    .Q_N(_00073_),
    .Q(\exec.pc[1] ));
 sg13g2_dfrbp_1 \pc[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3749),
    .D(_02503_),
    .Q_N(_00074_),
    .Q(\exec.pc[2] ));
 sg13g2_dfrbp_1 \pc[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3750),
    .D(_02504_),
    .Q_N(_00075_),
    .Q(\exec.pc[3] ));
 sg13g2_dfrbp_1 \pc[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3751),
    .D(_02505_),
    .Q_N(_00076_),
    .Q(\exec.pc[4] ));
 sg13g2_dfrbp_1 \pc[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3752),
    .D(_02506_),
    .Q_N(_00077_),
    .Q(\exec.pc[5] ));
 sg13g2_dfrbp_1 \pc[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3753),
    .D(_02507_),
    .Q_N(_00078_),
    .Q(\exec.pc[6] ));
 sg13g2_dfrbp_1 \pc[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3754),
    .D(_02508_),
    .Q_N(_00079_),
    .Q(\exec.pc[7] ));
 sg13g2_dfrbp_1 \shift_reg[0]$_SDFF_PN0_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3755),
    .D(_02509_),
    .Q_N(_13274_),
    .Q(\shift_reg[0] ));
 sg13g2_dfrbp_1 \shift_reg[1]$_SDFF_PN0_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3756),
    .D(_02510_),
    .Q_N(_13273_),
    .Q(\shift_reg[1] ));
 sg13g2_dfrbp_1 \shift_reg[2]$_SDFF_PN0_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3757),
    .D(_02511_),
    .Q_N(_13272_),
    .Q(\shift_reg[2] ));
 sg13g2_dfrbp_1 \shift_reg[3]$_SDFF_PN0_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3758),
    .D(_02512_),
    .Q_N(_13271_),
    .Q(\shift_reg[3] ));
 sg13g2_dfrbp_1 \shift_reg[4]$_SDFF_PN0_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3759),
    .D(_02513_),
    .Q_N(_13270_),
    .Q(\shift_reg[4] ));
 sg13g2_dfrbp_1 \shift_reg[5]$_SDFF_PN0_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3760),
    .D(_02514_),
    .Q_N(_13269_),
    .Q(\shift_reg[5] ));
 sg13g2_dfrbp_1 \shift_reg[6]$_SDFF_PN0_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3761),
    .D(_02515_),
    .Q_N(_13268_),
    .Q(\shift_reg[6] ));
 sg13g2_dfrbp_1 \shift_reg[7]$_SDFF_PN0_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3762),
    .D(_02516_),
    .Q_N(_13267_),
    .Q(\shift_reg[7] ));
 sg13g2_dfrbp_1 \single_step$_SDFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net3763),
    .D(_02517_),
    .Q_N(_00069_),
    .Q(single_step));
 sg13g2_dfrbp_1 \sp[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3764),
    .D(_02518_),
    .Q_N(_00065_),
    .Q(\exec.sp[0] ));
 sg13g2_dfrbp_1 \sp[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3765),
    .D(_02519_),
    .Q_N(_00066_),
    .Q(\exec.sp[1] ));
 sg13g2_dfrbp_1 \sp[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3766),
    .D(_02520_),
    .Q_N(_00067_),
    .Q(\exec.sp[2] ));
 sg13g2_dfrbp_1 \sp[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3767),
    .D(_02521_),
    .Q_N(_00039_),
    .Q(\exec.sp[3] ));
 sg13g2_dfrbp_1 \sp[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3768),
    .D(_02522_),
    .Q_N(_00048_),
    .Q(\exec.sp[4] ));
 sg13g2_dfrbp_1 \stack[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net3769),
    .D(_02523_),
    .Q_N(_00031_),
    .Q(\stack[0][0] ));
 sg13g2_dfrbp_1 \stack[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3770),
    .D(_02524_),
    .Q_N(_13266_),
    .Q(\stack[0][1] ));
 sg13g2_dfrbp_1 \stack[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3771),
    .D(_02525_),
    .Q_N(_13265_),
    .Q(\stack[0][2] ));
 sg13g2_dfrbp_1 \stack[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3772),
    .D(_02526_),
    .Q_N(_13264_),
    .Q(\stack[0][3] ));
 sg13g2_dfrbp_1 \stack[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net3773),
    .D(_02527_),
    .Q_N(_13263_),
    .Q(\stack[0][4] ));
 sg13g2_dfrbp_1 \stack[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3774),
    .D(_02528_),
    .Q_N(_13262_),
    .Q(\stack[0][5] ));
 sg13g2_dfrbp_1 \stack[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3775),
    .D(_02529_),
    .Q_N(_13261_),
    .Q(\stack[0][6] ));
 sg13g2_dfrbp_1 \stack[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3776),
    .D(_02530_),
    .Q_N(_13260_),
    .Q(\stack[0][7] ));
 sg13g2_dfrbp_1 \stack[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net3777),
    .D(_02531_),
    .Q_N(_00042_),
    .Q(\stack[10][0] ));
 sg13g2_dfrbp_1 \stack[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net3778),
    .D(_02532_),
    .Q_N(_13259_),
    .Q(\stack[10][1] ));
 sg13g2_dfrbp_1 \stack[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net3779),
    .D(_02533_),
    .Q_N(_13258_),
    .Q(\stack[10][2] ));
 sg13g2_dfrbp_1 \stack[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net3780),
    .D(_02534_),
    .Q_N(_13257_),
    .Q(\stack[10][3] ));
 sg13g2_dfrbp_1 \stack[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net3781),
    .D(_02535_),
    .Q_N(_13256_),
    .Q(\stack[10][4] ));
 sg13g2_dfrbp_1 \stack[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net3782),
    .D(_02536_),
    .Q_N(_13255_),
    .Q(\stack[10][5] ));
 sg13g2_dfrbp_1 \stack[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net3783),
    .D(_02537_),
    .Q_N(_13254_),
    .Q(\stack[10][6] ));
 sg13g2_dfrbp_1 \stack[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net3784),
    .D(_02538_),
    .Q_N(_13253_),
    .Q(\stack[10][7] ));
 sg13g2_dfrbp_1 \stack[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net3785),
    .D(_02539_),
    .Q_N(_00043_),
    .Q(\stack[11][0] ));
 sg13g2_dfrbp_1 \stack[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net3786),
    .D(_02540_),
    .Q_N(_13252_),
    .Q(\stack[11][1] ));
 sg13g2_dfrbp_1 \stack[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net3787),
    .D(_02541_),
    .Q_N(_13251_),
    .Q(\stack[11][2] ));
 sg13g2_dfrbp_1 \stack[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net3788),
    .D(_02542_),
    .Q_N(_13250_),
    .Q(\stack[11][3] ));
 sg13g2_dfrbp_1 \stack[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net3789),
    .D(_02543_),
    .Q_N(_13249_),
    .Q(\stack[11][4] ));
 sg13g2_dfrbp_1 \stack[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net3790),
    .D(_02544_),
    .Q_N(_13248_),
    .Q(\stack[11][5] ));
 sg13g2_dfrbp_1 \stack[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net3791),
    .D(_02545_),
    .Q_N(_13247_),
    .Q(\stack[11][6] ));
 sg13g2_dfrbp_1 \stack[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net3792),
    .D(_02546_),
    .Q_N(_13246_),
    .Q(\stack[11][7] ));
 sg13g2_dfrbp_1 \stack[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net3793),
    .D(_02547_),
    .Q_N(_00044_),
    .Q(\stack[12][0] ));
 sg13g2_dfrbp_1 \stack[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net3794),
    .D(_02548_),
    .Q_N(_13245_),
    .Q(\stack[12][1] ));
 sg13g2_dfrbp_1 \stack[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net3795),
    .D(_02549_),
    .Q_N(_13244_),
    .Q(\stack[12][2] ));
 sg13g2_dfrbp_1 \stack[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net3796),
    .D(_02550_),
    .Q_N(_13243_),
    .Q(\stack[12][3] ));
 sg13g2_dfrbp_1 \stack[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net3797),
    .D(_02551_),
    .Q_N(_13242_),
    .Q(\stack[12][4] ));
 sg13g2_dfrbp_1 \stack[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net3798),
    .D(_02552_),
    .Q_N(_13241_),
    .Q(\stack[12][5] ));
 sg13g2_dfrbp_1 \stack[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net3799),
    .D(_02553_),
    .Q_N(_13240_),
    .Q(\stack[12][6] ));
 sg13g2_dfrbp_1 \stack[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net3800),
    .D(_02554_),
    .Q_N(_13239_),
    .Q(\stack[12][7] ));
 sg13g2_dfrbp_1 \stack[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net3801),
    .D(_02555_),
    .Q_N(_00045_),
    .Q(\stack[13][0] ));
 sg13g2_dfrbp_1 \stack[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net3802),
    .D(_02556_),
    .Q_N(_13238_),
    .Q(\stack[13][1] ));
 sg13g2_dfrbp_1 \stack[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net3803),
    .D(_02557_),
    .Q_N(_13237_),
    .Q(\stack[13][2] ));
 sg13g2_dfrbp_1 \stack[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net3804),
    .D(_02558_),
    .Q_N(_13236_),
    .Q(\stack[13][3] ));
 sg13g2_dfrbp_1 \stack[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net3805),
    .D(_02559_),
    .Q_N(_13235_),
    .Q(\stack[13][4] ));
 sg13g2_dfrbp_1 \stack[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net3806),
    .D(_02560_),
    .Q_N(_13234_),
    .Q(\stack[13][5] ));
 sg13g2_dfrbp_1 \stack[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net3807),
    .D(_02561_),
    .Q_N(_13233_),
    .Q(\stack[13][6] ));
 sg13g2_dfrbp_1 \stack[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net3808),
    .D(_02562_),
    .Q_N(_13232_),
    .Q(\stack[13][7] ));
 sg13g2_dfrbp_1 \stack[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net3809),
    .D(_02563_),
    .Q_N(_00046_),
    .Q(\stack[14][0] ));
 sg13g2_dfrbp_1 \stack[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net3810),
    .D(_02564_),
    .Q_N(_13231_),
    .Q(\stack[14][1] ));
 sg13g2_dfrbp_1 \stack[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net3811),
    .D(_02565_),
    .Q_N(_13230_),
    .Q(\stack[14][2] ));
 sg13g2_dfrbp_1 \stack[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net3812),
    .D(_02566_),
    .Q_N(_13229_),
    .Q(\stack[14][3] ));
 sg13g2_dfrbp_1 \stack[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net3813),
    .D(_02567_),
    .Q_N(_13228_),
    .Q(\stack[14][4] ));
 sg13g2_dfrbp_1 \stack[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net3814),
    .D(_02568_),
    .Q_N(_13227_),
    .Q(\stack[14][5] ));
 sg13g2_dfrbp_1 \stack[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net3815),
    .D(_02569_),
    .Q_N(_13226_),
    .Q(\stack[14][6] ));
 sg13g2_dfrbp_1 \stack[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net3816),
    .D(_02570_),
    .Q_N(_13225_),
    .Q(\stack[14][7] ));
 sg13g2_dfrbp_1 \stack[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net3817),
    .D(_02571_),
    .Q_N(_00047_),
    .Q(\stack[15][0] ));
 sg13g2_dfrbp_1 \stack[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net3818),
    .D(_02572_),
    .Q_N(_13224_),
    .Q(\stack[15][1] ));
 sg13g2_dfrbp_1 \stack[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net3819),
    .D(_02573_),
    .Q_N(_13223_),
    .Q(\stack[15][2] ));
 sg13g2_dfrbp_1 \stack[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net3820),
    .D(_02574_),
    .Q_N(_13222_),
    .Q(\stack[15][3] ));
 sg13g2_dfrbp_1 \stack[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net3821),
    .D(_02575_),
    .Q_N(_13221_),
    .Q(\stack[15][4] ));
 sg13g2_dfrbp_1 \stack[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net3822),
    .D(_02576_),
    .Q_N(_13220_),
    .Q(\stack[15][5] ));
 sg13g2_dfrbp_1 \stack[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net3823),
    .D(_02577_),
    .Q_N(_13219_),
    .Q(\stack[15][6] ));
 sg13g2_dfrbp_1 \stack[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net3824),
    .D(_02578_),
    .Q_N(_13218_),
    .Q(\stack[15][7] ));
 sg13g2_dfrbp_1 \stack[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3825),
    .D(_02579_),
    .Q_N(_00049_),
    .Q(\stack[16][0] ));
 sg13g2_dfrbp_1 \stack[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3826),
    .D(_02580_),
    .Q_N(_13217_),
    .Q(\stack[16][1] ));
 sg13g2_dfrbp_1 \stack[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3827),
    .D(_02581_),
    .Q_N(_13216_),
    .Q(\stack[16][2] ));
 sg13g2_dfrbp_1 \stack[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3828),
    .D(_02582_),
    .Q_N(_13215_),
    .Q(\stack[16][3] ));
 sg13g2_dfrbp_1 \stack[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3829),
    .D(_02583_),
    .Q_N(_13214_),
    .Q(\stack[16][4] ));
 sg13g2_dfrbp_1 \stack[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3830),
    .D(_02584_),
    .Q_N(_13213_),
    .Q(\stack[16][5] ));
 sg13g2_dfrbp_1 \stack[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3831),
    .D(_02585_),
    .Q_N(_13212_),
    .Q(\stack[16][6] ));
 sg13g2_dfrbp_1 \stack[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3832),
    .D(_02586_),
    .Q_N(_13211_),
    .Q(\stack[16][7] ));
 sg13g2_dfrbp_1 \stack[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3833),
    .D(_02587_),
    .Q_N(_00050_),
    .Q(\stack[17][0] ));
 sg13g2_dfrbp_1 \stack[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3834),
    .D(_02588_),
    .Q_N(_13210_),
    .Q(\stack[17][1] ));
 sg13g2_dfrbp_1 \stack[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3835),
    .D(_02589_),
    .Q_N(_13209_),
    .Q(\stack[17][2] ));
 sg13g2_dfrbp_1 \stack[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net3836),
    .D(_02590_),
    .Q_N(_13208_),
    .Q(\stack[17][3] ));
 sg13g2_dfrbp_1 \stack[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3837),
    .D(_02591_),
    .Q_N(_13207_),
    .Q(\stack[17][4] ));
 sg13g2_dfrbp_1 \stack[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3838),
    .D(_02592_),
    .Q_N(_13206_),
    .Q(\stack[17][5] ));
 sg13g2_dfrbp_1 \stack[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net3839),
    .D(_02593_),
    .Q_N(_13205_),
    .Q(\stack[17][6] ));
 sg13g2_dfrbp_1 \stack[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net3840),
    .D(_02594_),
    .Q_N(_13204_),
    .Q(\stack[17][7] ));
 sg13g2_dfrbp_1 \stack[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net3841),
    .D(_02595_),
    .Q_N(_00051_),
    .Q(\stack[18][0] ));
 sg13g2_dfrbp_1 \stack[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net3842),
    .D(_02596_),
    .Q_N(_13203_),
    .Q(\stack[18][1] ));
 sg13g2_dfrbp_1 \stack[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net3843),
    .D(_02597_),
    .Q_N(_13202_),
    .Q(\stack[18][2] ));
 sg13g2_dfrbp_1 \stack[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net3844),
    .D(_02598_),
    .Q_N(_13201_),
    .Q(\stack[18][3] ));
 sg13g2_dfrbp_1 \stack[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net3845),
    .D(_02599_),
    .Q_N(_13200_),
    .Q(\stack[18][4] ));
 sg13g2_dfrbp_1 \stack[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net3846),
    .D(_02600_),
    .Q_N(_13199_),
    .Q(\stack[18][5] ));
 sg13g2_dfrbp_1 \stack[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net3847),
    .D(_02601_),
    .Q_N(_13198_),
    .Q(\stack[18][6] ));
 sg13g2_dfrbp_1 \stack[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net3848),
    .D(_02602_),
    .Q_N(_13197_),
    .Q(\stack[18][7] ));
 sg13g2_dfrbp_1 \stack[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3849),
    .D(_02603_),
    .Q_N(_00052_),
    .Q(\stack[19][0] ));
 sg13g2_dfrbp_1 \stack[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3850),
    .D(_02604_),
    .Q_N(_13196_),
    .Q(\stack[19][1] ));
 sg13g2_dfrbp_1 \stack[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3851),
    .D(_02605_),
    .Q_N(_13195_),
    .Q(\stack[19][2] ));
 sg13g2_dfrbp_1 \stack[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3852),
    .D(_02606_),
    .Q_N(_13194_),
    .Q(\stack[19][3] ));
 sg13g2_dfrbp_1 \stack[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3853),
    .D(_02607_),
    .Q_N(_13193_),
    .Q(\stack[19][4] ));
 sg13g2_dfrbp_1 \stack[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3854),
    .D(_02608_),
    .Q_N(_13192_),
    .Q(\stack[19][5] ));
 sg13g2_dfrbp_1 \stack[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3855),
    .D(_02609_),
    .Q_N(_13191_),
    .Q(\stack[19][6] ));
 sg13g2_dfrbp_1 \stack[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3856),
    .D(_02610_),
    .Q_N(_13190_),
    .Q(\stack[19][7] ));
 sg13g2_dfrbp_1 \stack[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net3857),
    .D(_02611_),
    .Q_N(_00032_),
    .Q(\stack[1][0] ));
 sg13g2_dfrbp_1 \stack[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net3858),
    .D(_02612_),
    .Q_N(_13189_),
    .Q(\stack[1][1] ));
 sg13g2_dfrbp_1 \stack[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net3859),
    .D(_02613_),
    .Q_N(_13188_),
    .Q(\stack[1][2] ));
 sg13g2_dfrbp_1 \stack[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net3860),
    .D(_02614_),
    .Q_N(_13187_),
    .Q(\stack[1][3] ));
 sg13g2_dfrbp_1 \stack[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net3861),
    .D(_02615_),
    .Q_N(_13186_),
    .Q(\stack[1][4] ));
 sg13g2_dfrbp_1 \stack[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net3862),
    .D(_02616_),
    .Q_N(_13185_),
    .Q(\stack[1][5] ));
 sg13g2_dfrbp_1 \stack[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net3863),
    .D(_02617_),
    .Q_N(_13184_),
    .Q(\stack[1][6] ));
 sg13g2_dfrbp_1 \stack[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net3864),
    .D(_02618_),
    .Q_N(_13183_),
    .Q(\stack[1][7] ));
 sg13g2_dfrbp_1 \stack[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net3865),
    .D(_02619_),
    .Q_N(_00053_),
    .Q(\stack[20][0] ));
 sg13g2_dfrbp_1 \stack[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net3866),
    .D(_02620_),
    .Q_N(_13182_),
    .Q(\stack[20][1] ));
 sg13g2_dfrbp_1 \stack[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net3867),
    .D(_02621_),
    .Q_N(_13181_),
    .Q(\stack[20][2] ));
 sg13g2_dfrbp_1 \stack[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3868),
    .D(_02622_),
    .Q_N(_13180_),
    .Q(\stack[20][3] ));
 sg13g2_dfrbp_1 \stack[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3869),
    .D(_02623_),
    .Q_N(_13179_),
    .Q(\stack[20][4] ));
 sg13g2_dfrbp_1 \stack[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3870),
    .D(_02624_),
    .Q_N(_13178_),
    .Q(\stack[20][5] ));
 sg13g2_dfrbp_1 \stack[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3871),
    .D(_02625_),
    .Q_N(_13177_),
    .Q(\stack[20][6] ));
 sg13g2_dfrbp_1 \stack[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3872),
    .D(_02626_),
    .Q_N(_13176_),
    .Q(\stack[20][7] ));
 sg13g2_dfrbp_1 \stack[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net3873),
    .D(_02627_),
    .Q_N(_00054_),
    .Q(\stack[21][0] ));
 sg13g2_dfrbp_1 \stack[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net3874),
    .D(_02628_),
    .Q_N(_13175_),
    .Q(\stack[21][1] ));
 sg13g2_dfrbp_1 \stack[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net3875),
    .D(_02629_),
    .Q_N(_13174_),
    .Q(\stack[21][2] ));
 sg13g2_dfrbp_1 \stack[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3876),
    .D(_02630_),
    .Q_N(_13173_),
    .Q(\stack[21][3] ));
 sg13g2_dfrbp_1 \stack[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net3877),
    .D(_02631_),
    .Q_N(_13172_),
    .Q(\stack[21][4] ));
 sg13g2_dfrbp_1 \stack[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net3878),
    .D(_02632_),
    .Q_N(_13171_),
    .Q(\stack[21][5] ));
 sg13g2_dfrbp_1 \stack[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net3879),
    .D(_02633_),
    .Q_N(_13170_),
    .Q(\stack[21][6] ));
 sg13g2_dfrbp_1 \stack[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net3880),
    .D(_02634_),
    .Q_N(_13169_),
    .Q(\stack[21][7] ));
 sg13g2_dfrbp_1 \stack[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3881),
    .D(_02635_),
    .Q_N(_00055_),
    .Q(\stack[22][0] ));
 sg13g2_dfrbp_1 \stack[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3882),
    .D(_02636_),
    .Q_N(_13168_),
    .Q(\stack[22][1] ));
 sg13g2_dfrbp_1 \stack[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3883),
    .D(_02637_),
    .Q_N(_13167_),
    .Q(\stack[22][2] ));
 sg13g2_dfrbp_1 \stack[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3884),
    .D(_02638_),
    .Q_N(_13166_),
    .Q(\stack[22][3] ));
 sg13g2_dfrbp_1 \stack[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3885),
    .D(_02639_),
    .Q_N(_13165_),
    .Q(\stack[22][4] ));
 sg13g2_dfrbp_1 \stack[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3886),
    .D(_02640_),
    .Q_N(_13164_),
    .Q(\stack[22][5] ));
 sg13g2_dfrbp_1 \stack[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3887),
    .D(_02641_),
    .Q_N(_13163_),
    .Q(\stack[22][6] ));
 sg13g2_dfrbp_1 \stack[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3888),
    .D(_02642_),
    .Q_N(_13162_),
    .Q(\stack[22][7] ));
 sg13g2_dfrbp_1 \stack[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net3889),
    .D(_02643_),
    .Q_N(_00056_),
    .Q(\stack[23][0] ));
 sg13g2_dfrbp_1 \stack[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net3890),
    .D(_02644_),
    .Q_N(_13161_),
    .Q(\stack[23][1] ));
 sg13g2_dfrbp_1 \stack[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net3891),
    .D(_02645_),
    .Q_N(_13160_),
    .Q(\stack[23][2] ));
 sg13g2_dfrbp_1 \stack[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net3892),
    .D(_02646_),
    .Q_N(_13159_),
    .Q(\stack[23][3] ));
 sg13g2_dfrbp_1 \stack[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net3893),
    .D(_02647_),
    .Q_N(_13158_),
    .Q(\stack[23][4] ));
 sg13g2_dfrbp_1 \stack[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net3894),
    .D(_02648_),
    .Q_N(_13157_),
    .Q(\stack[23][5] ));
 sg13g2_dfrbp_1 \stack[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net3895),
    .D(_02649_),
    .Q_N(_13156_),
    .Q(\stack[23][6] ));
 sg13g2_dfrbp_1 \stack[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net3896),
    .D(_02650_),
    .Q_N(_13155_),
    .Q(\stack[23][7] ));
 sg13g2_dfrbp_1 \stack[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net3897),
    .D(_02651_),
    .Q_N(_00057_),
    .Q(\stack[24][0] ));
 sg13g2_dfrbp_1 \stack[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net3898),
    .D(_02652_),
    .Q_N(_13154_),
    .Q(\stack[24][1] ));
 sg13g2_dfrbp_1 \stack[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net3899),
    .D(_02653_),
    .Q_N(_13153_),
    .Q(\stack[24][2] ));
 sg13g2_dfrbp_1 \stack[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net3900),
    .D(_02654_),
    .Q_N(_13152_),
    .Q(\stack[24][3] ));
 sg13g2_dfrbp_1 \stack[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net3901),
    .D(_02655_),
    .Q_N(_13151_),
    .Q(\stack[24][4] ));
 sg13g2_dfrbp_1 \stack[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net3902),
    .D(_02656_),
    .Q_N(_13150_),
    .Q(\stack[24][5] ));
 sg13g2_dfrbp_1 \stack[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net3903),
    .D(_02657_),
    .Q_N(_13149_),
    .Q(\stack[24][6] ));
 sg13g2_dfrbp_1 \stack[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net3904),
    .D(_02658_),
    .Q_N(_13148_),
    .Q(\stack[24][7] ));
 sg13g2_dfrbp_1 \stack[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net3905),
    .D(_02659_),
    .Q_N(_00058_),
    .Q(\stack[25][0] ));
 sg13g2_dfrbp_1 \stack[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net3906),
    .D(_02660_),
    .Q_N(_13147_),
    .Q(\stack[25][1] ));
 sg13g2_dfrbp_1 \stack[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net3907),
    .D(_02661_),
    .Q_N(_13146_),
    .Q(\stack[25][2] ));
 sg13g2_dfrbp_1 \stack[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net3908),
    .D(_02662_),
    .Q_N(_13145_),
    .Q(\stack[25][3] ));
 sg13g2_dfrbp_1 \stack[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net3909),
    .D(_02663_),
    .Q_N(_13144_),
    .Q(\stack[25][4] ));
 sg13g2_dfrbp_1 \stack[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net3910),
    .D(_02664_),
    .Q_N(_13143_),
    .Q(\stack[25][5] ));
 sg13g2_dfrbp_1 \stack[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net3911),
    .D(_02665_),
    .Q_N(_13142_),
    .Q(\stack[25][6] ));
 sg13g2_dfrbp_1 \stack[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net3912),
    .D(_02666_),
    .Q_N(_13141_),
    .Q(\stack[25][7] ));
 sg13g2_dfrbp_1 \stack[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net3913),
    .D(_02667_),
    .Q_N(_00059_),
    .Q(\stack[26][0] ));
 sg13g2_dfrbp_1 \stack[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net3914),
    .D(_02668_),
    .Q_N(_13140_),
    .Q(\stack[26][1] ));
 sg13g2_dfrbp_1 \stack[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net3915),
    .D(_02669_),
    .Q_N(_13139_),
    .Q(\stack[26][2] ));
 sg13g2_dfrbp_1 \stack[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net3916),
    .D(_02670_),
    .Q_N(_13138_),
    .Q(\stack[26][3] ));
 sg13g2_dfrbp_1 \stack[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net3917),
    .D(_02671_),
    .Q_N(_13137_),
    .Q(\stack[26][4] ));
 sg13g2_dfrbp_1 \stack[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net3918),
    .D(_02672_),
    .Q_N(_13136_),
    .Q(\stack[26][5] ));
 sg13g2_dfrbp_1 \stack[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net3919),
    .D(_02673_),
    .Q_N(_13135_),
    .Q(\stack[26][6] ));
 sg13g2_dfrbp_1 \stack[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net3920),
    .D(_02674_),
    .Q_N(_13134_),
    .Q(\stack[26][7] ));
 sg13g2_dfrbp_1 \stack[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net3921),
    .D(_02675_),
    .Q_N(_00060_),
    .Q(\stack[27][0] ));
 sg13g2_dfrbp_1 \stack[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net3922),
    .D(_02676_),
    .Q_N(_13133_),
    .Q(\stack[27][1] ));
 sg13g2_dfrbp_1 \stack[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net3923),
    .D(_02677_),
    .Q_N(_13132_),
    .Q(\stack[27][2] ));
 sg13g2_dfrbp_1 \stack[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net3924),
    .D(_02678_),
    .Q_N(_13131_),
    .Q(\stack[27][3] ));
 sg13g2_dfrbp_1 \stack[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net3925),
    .D(_02679_),
    .Q_N(_13130_),
    .Q(\stack[27][4] ));
 sg13g2_dfrbp_1 \stack[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net3926),
    .D(_02680_),
    .Q_N(_13129_),
    .Q(\stack[27][5] ));
 sg13g2_dfrbp_1 \stack[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net3927),
    .D(_02681_),
    .Q_N(_13128_),
    .Q(\stack[27][6] ));
 sg13g2_dfrbp_1 \stack[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net3928),
    .D(_02682_),
    .Q_N(_13127_),
    .Q(\stack[27][7] ));
 sg13g2_dfrbp_1 \stack[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net3929),
    .D(_02683_),
    .Q_N(_00061_),
    .Q(\stack[28][0] ));
 sg13g2_dfrbp_1 \stack[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net3930),
    .D(_02684_),
    .Q_N(_13126_),
    .Q(\stack[28][1] ));
 sg13g2_dfrbp_1 \stack[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net3931),
    .D(_02685_),
    .Q_N(_13125_),
    .Q(\stack[28][2] ));
 sg13g2_dfrbp_1 \stack[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net3932),
    .D(_02686_),
    .Q_N(_13124_),
    .Q(\stack[28][3] ));
 sg13g2_dfrbp_1 \stack[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net3933),
    .D(_02687_),
    .Q_N(_13123_),
    .Q(\stack[28][4] ));
 sg13g2_dfrbp_1 \stack[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net3934),
    .D(_02688_),
    .Q_N(_13122_),
    .Q(\stack[28][5] ));
 sg13g2_dfrbp_1 \stack[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net3935),
    .D(_02689_),
    .Q_N(_13121_),
    .Q(\stack[28][6] ));
 sg13g2_dfrbp_1 \stack[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net3936),
    .D(_02690_),
    .Q_N(_13120_),
    .Q(\stack[28][7] ));
 sg13g2_dfrbp_1 \stack[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net3937),
    .D(_02691_),
    .Q_N(_00062_),
    .Q(\stack[29][0] ));
 sg13g2_dfrbp_1 \stack[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net3938),
    .D(_02692_),
    .Q_N(_13119_),
    .Q(\stack[29][1] ));
 sg13g2_dfrbp_1 \stack[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net3939),
    .D(_02693_),
    .Q_N(_13118_),
    .Q(\stack[29][2] ));
 sg13g2_dfrbp_1 \stack[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net3940),
    .D(_02694_),
    .Q_N(_13117_),
    .Q(\stack[29][3] ));
 sg13g2_dfrbp_1 \stack[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net3941),
    .D(_02695_),
    .Q_N(_13116_),
    .Q(\stack[29][4] ));
 sg13g2_dfrbp_1 \stack[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net3942),
    .D(_02696_),
    .Q_N(_13115_),
    .Q(\stack[29][5] ));
 sg13g2_dfrbp_1 \stack[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net3943),
    .D(_02697_),
    .Q_N(_13114_),
    .Q(\stack[29][6] ));
 sg13g2_dfrbp_1 \stack[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net3944),
    .D(_02698_),
    .Q_N(_13113_),
    .Q(\stack[29][7] ));
 sg13g2_dfrbp_1 \stack[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net3945),
    .D(_02699_),
    .Q_N(_00033_),
    .Q(\stack[2][0] ));
 sg13g2_dfrbp_1 \stack[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net3946),
    .D(_02700_),
    .Q_N(_13112_),
    .Q(\stack[2][1] ));
 sg13g2_dfrbp_1 \stack[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net3947),
    .D(_02701_),
    .Q_N(_13111_),
    .Q(\stack[2][2] ));
 sg13g2_dfrbp_1 \stack[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net3948),
    .D(_02702_),
    .Q_N(_13110_),
    .Q(\stack[2][3] ));
 sg13g2_dfrbp_1 \stack[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net3949),
    .D(_02703_),
    .Q_N(_13109_),
    .Q(\stack[2][4] ));
 sg13g2_dfrbp_1 \stack[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net3950),
    .D(_02704_),
    .Q_N(_13108_),
    .Q(\stack[2][5] ));
 sg13g2_dfrbp_1 \stack[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net3951),
    .D(_02705_),
    .Q_N(_13107_),
    .Q(\stack[2][6] ));
 sg13g2_dfrbp_1 \stack[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net3952),
    .D(_02706_),
    .Q_N(_13106_),
    .Q(\stack[2][7] ));
 sg13g2_dfrbp_1 \stack[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net3953),
    .D(_02707_),
    .Q_N(_00063_),
    .Q(\stack[30][0] ));
 sg13g2_dfrbp_1 \stack[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net3954),
    .D(_02708_),
    .Q_N(_13105_),
    .Q(\stack[30][1] ));
 sg13g2_dfrbp_1 \stack[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net3955),
    .D(_02709_),
    .Q_N(_13104_),
    .Q(\stack[30][2] ));
 sg13g2_dfrbp_1 \stack[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net3956),
    .D(_02710_),
    .Q_N(_13103_),
    .Q(\stack[30][3] ));
 sg13g2_dfrbp_1 \stack[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net3957),
    .D(_02711_),
    .Q_N(_13102_),
    .Q(\stack[30][4] ));
 sg13g2_dfrbp_1 \stack[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net3958),
    .D(_02712_),
    .Q_N(_13101_),
    .Q(\stack[30][5] ));
 sg13g2_dfrbp_1 \stack[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net3959),
    .D(_02713_),
    .Q_N(_13100_),
    .Q(\stack[30][6] ));
 sg13g2_dfrbp_1 \stack[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net3960),
    .D(_02714_),
    .Q_N(_13099_),
    .Q(\stack[30][7] ));
 sg13g2_dfrbp_1 \stack[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net3961),
    .D(_02715_),
    .Q_N(_00064_),
    .Q(\stack[31][0] ));
 sg13g2_dfrbp_1 \stack[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net3962),
    .D(_02716_),
    .Q_N(_13098_),
    .Q(\stack[31][1] ));
 sg13g2_dfrbp_1 \stack[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net3963),
    .D(_02717_),
    .Q_N(_13097_),
    .Q(\stack[31][2] ));
 sg13g2_dfrbp_1 \stack[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net3964),
    .D(_02718_),
    .Q_N(_13096_),
    .Q(\stack[31][3] ));
 sg13g2_dfrbp_1 \stack[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net3965),
    .D(_02719_),
    .Q_N(_13095_),
    .Q(\stack[31][4] ));
 sg13g2_dfrbp_1 \stack[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net3966),
    .D(_02720_),
    .Q_N(_13094_),
    .Q(\stack[31][5] ));
 sg13g2_dfrbp_1 \stack[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net3967),
    .D(_02721_),
    .Q_N(_13093_),
    .Q(\stack[31][6] ));
 sg13g2_dfrbp_1 \stack[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net3968),
    .D(_02722_),
    .Q_N(_13092_),
    .Q(\stack[31][7] ));
 sg13g2_dfrbp_1 \stack[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3969),
    .D(_02723_),
    .Q_N(_00034_),
    .Q(\stack[3][0] ));
 sg13g2_dfrbp_1 \stack[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3970),
    .D(_02724_),
    .Q_N(_13091_),
    .Q(\stack[3][1] ));
 sg13g2_dfrbp_1 \stack[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3971),
    .D(_02725_),
    .Q_N(_13090_),
    .Q(\stack[3][2] ));
 sg13g2_dfrbp_1 \stack[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3972),
    .D(_02726_),
    .Q_N(_13089_),
    .Q(\stack[3][3] ));
 sg13g2_dfrbp_1 \stack[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3973),
    .D(_02727_),
    .Q_N(_13088_),
    .Q(\stack[3][4] ));
 sg13g2_dfrbp_1 \stack[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3974),
    .D(_02728_),
    .Q_N(_13087_),
    .Q(\stack[3][5] ));
 sg13g2_dfrbp_1 \stack[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3975),
    .D(_02729_),
    .Q_N(_13086_),
    .Q(\stack[3][6] ));
 sg13g2_dfrbp_1 \stack[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3976),
    .D(_02730_),
    .Q_N(_13085_),
    .Q(\stack[3][7] ));
 sg13g2_dfrbp_1 \stack[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net3977),
    .D(_02731_),
    .Q_N(_00035_),
    .Q(\stack[4][0] ));
 sg13g2_dfrbp_1 \stack[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net3978),
    .D(_02732_),
    .Q_N(_13084_),
    .Q(\stack[4][1] ));
 sg13g2_dfrbp_1 \stack[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net3979),
    .D(_02733_),
    .Q_N(_13083_),
    .Q(\stack[4][2] ));
 sg13g2_dfrbp_1 \stack[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net3980),
    .D(_02734_),
    .Q_N(_13082_),
    .Q(\stack[4][3] ));
 sg13g2_dfrbp_1 \stack[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3981),
    .D(_02735_),
    .Q_N(_13081_),
    .Q(\stack[4][4] ));
 sg13g2_dfrbp_1 \stack[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net3982),
    .D(_02736_),
    .Q_N(_13080_),
    .Q(\stack[4][5] ));
 sg13g2_dfrbp_1 \stack[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net3983),
    .D(_02737_),
    .Q_N(_13079_),
    .Q(\stack[4][6] ));
 sg13g2_dfrbp_1 \stack[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net3984),
    .D(_02738_),
    .Q_N(_13078_),
    .Q(\stack[4][7] ));
 sg13g2_dfrbp_1 \stack[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3985),
    .D(_02739_),
    .Q_N(_00036_),
    .Q(\stack[5][0] ));
 sg13g2_dfrbp_1 \stack[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net3986),
    .D(_02740_),
    .Q_N(_13077_),
    .Q(\stack[5][1] ));
 sg13g2_dfrbp_1 \stack[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3987),
    .D(_02741_),
    .Q_N(_13076_),
    .Q(\stack[5][2] ));
 sg13g2_dfrbp_1 \stack[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net3988),
    .D(_02742_),
    .Q_N(_13075_),
    .Q(\stack[5][3] ));
 sg13g2_dfrbp_1 \stack[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3989),
    .D(_02743_),
    .Q_N(_13074_),
    .Q(\stack[5][4] ));
 sg13g2_dfrbp_1 \stack[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3990),
    .D(_02744_),
    .Q_N(_13073_),
    .Q(\stack[5][5] ));
 sg13g2_dfrbp_1 \stack[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net3991),
    .D(_02745_),
    .Q_N(_13072_),
    .Q(\stack[5][6] ));
 sg13g2_dfrbp_1 \stack[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3992),
    .D(_02746_),
    .Q_N(_13071_),
    .Q(\stack[5][7] ));
 sg13g2_dfrbp_1 \stack[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3993),
    .D(_02747_),
    .Q_N(_00037_),
    .Q(\stack[6][0] ));
 sg13g2_dfrbp_1 \stack[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net3994),
    .D(_02748_),
    .Q_N(_13070_),
    .Q(\stack[6][1] ));
 sg13g2_dfrbp_1 \stack[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net3995),
    .D(_02749_),
    .Q_N(_13069_),
    .Q(\stack[6][2] ));
 sg13g2_dfrbp_1 \stack[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3996),
    .D(_02750_),
    .Q_N(_13068_),
    .Q(\stack[6][3] ));
 sg13g2_dfrbp_1 \stack[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3997),
    .D(_02751_),
    .Q_N(_13067_),
    .Q(\stack[6][4] ));
 sg13g2_dfrbp_1 \stack[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3998),
    .D(_02752_),
    .Q_N(_13066_),
    .Q(\stack[6][5] ));
 sg13g2_dfrbp_1 \stack[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3999),
    .D(_02753_),
    .Q_N(_13065_),
    .Q(\stack[6][6] ));
 sg13g2_dfrbp_1 \stack[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net4000),
    .D(_02754_),
    .Q_N(_13064_),
    .Q(\stack[6][7] ));
 sg13g2_dfrbp_1 \stack[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net4001),
    .D(_02755_),
    .Q_N(_00038_),
    .Q(\stack[7][0] ));
 sg13g2_dfrbp_1 \stack[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net4002),
    .D(_02756_),
    .Q_N(_13063_),
    .Q(\stack[7][1] ));
 sg13g2_dfrbp_1 \stack[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net4003),
    .D(_02757_),
    .Q_N(_13062_),
    .Q(\stack[7][2] ));
 sg13g2_dfrbp_1 \stack[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net4004),
    .D(_02758_),
    .Q_N(_13061_),
    .Q(\stack[7][3] ));
 sg13g2_dfrbp_1 \stack[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net4005),
    .D(_02759_),
    .Q_N(_13060_),
    .Q(\stack[7][4] ));
 sg13g2_dfrbp_1 \stack[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net4006),
    .D(_02760_),
    .Q_N(_13059_),
    .Q(\stack[7][5] ));
 sg13g2_dfrbp_1 \stack[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net4007),
    .D(_02761_),
    .Q_N(_13058_),
    .Q(\stack[7][6] ));
 sg13g2_dfrbp_1 \stack[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net4008),
    .D(_02762_),
    .Q_N(_13057_),
    .Q(\stack[7][7] ));
 sg13g2_dfrbp_1 \stack[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net4009),
    .D(_02763_),
    .Q_N(_00040_),
    .Q(\stack[8][0] ));
 sg13g2_dfrbp_1 \stack[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net4010),
    .D(_02764_),
    .Q_N(_13056_),
    .Q(\stack[8][1] ));
 sg13g2_dfrbp_1 \stack[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net4011),
    .D(_02765_),
    .Q_N(_13055_),
    .Q(\stack[8][2] ));
 sg13g2_dfrbp_1 \stack[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net4012),
    .D(_02766_),
    .Q_N(_13054_),
    .Q(\stack[8][3] ));
 sg13g2_dfrbp_1 \stack[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net4013),
    .D(_02767_),
    .Q_N(_13053_),
    .Q(\stack[8][4] ));
 sg13g2_dfrbp_1 \stack[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net4014),
    .D(_02768_),
    .Q_N(_13052_),
    .Q(\stack[8][5] ));
 sg13g2_dfrbp_1 \stack[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net4015),
    .D(_02769_),
    .Q_N(_13051_),
    .Q(\stack[8][6] ));
 sg13g2_dfrbp_1 \stack[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net4016),
    .D(_02770_),
    .Q_N(_13050_),
    .Q(\stack[8][7] ));
 sg13g2_dfrbp_1 \stack[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net4017),
    .D(_02771_),
    .Q_N(_00041_),
    .Q(\stack[9][0] ));
 sg13g2_dfrbp_1 \stack[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net4018),
    .D(_02772_),
    .Q_N(_13049_),
    .Q(\stack[9][1] ));
 sg13g2_dfrbp_1 \stack[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net4019),
    .D(_02773_),
    .Q_N(_13048_),
    .Q(\stack[9][2] ));
 sg13g2_dfrbp_1 \stack[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net4020),
    .D(_02774_),
    .Q_N(_13047_),
    .Q(\stack[9][3] ));
 sg13g2_dfrbp_1 \stack[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net4021),
    .D(_02775_),
    .Q_N(_13046_),
    .Q(\stack[9][4] ));
 sg13g2_dfrbp_1 \stack[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net4022),
    .D(_02776_),
    .Q_N(_13045_),
    .Q(\stack[9][5] ));
 sg13g2_dfrbp_1 \stack[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net4023),
    .D(_02777_),
    .Q_N(_13044_),
    .Q(\stack[9][6] ));
 sg13g2_dfrbp_1 \stack[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net4024),
    .D(_02778_),
    .Q_N(_15699_),
    .Q(\stack[9][7] ));
 sg13g2_dfrbp_1 \state[0]$_DFF_P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net4025),
    .D(_00008_),
    .Q_N(_15700_),
    .Q(o_sleep));
 sg13g2_dfrbp_1 \state[1]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net4026),
    .D(_00009_),
    .Q_N(_15701_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 \state[2]$_DFF_P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net4027),
    .D(_00010_),
    .Q_N(_15702_),
    .Q(o_wait_delay));
 sg13g2_dfrbp_1 \state[3]$_DFF_P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net4028),
    .D(_00011_),
    .Q_N(_00068_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 \state[4]$_DFF_P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net4029),
    .D(_00012_),
    .Q_N(_15703_),
    .Q(\state[4] ));
 sg13g2_dfrbp_1 \state[5]$_DFF_P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net4030),
    .D(_00013_),
    .Q_N(_00072_),
    .Q(\state[5] ));
 sg13g2_dfrbp_1 \state[6]$_DFF_P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net4031),
    .D(_00014_),
    .Q_N(_13043_),
    .Q(\state[6] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[0]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[1]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[2]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[3]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[4]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[5]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[6]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[7]),
    .X(net12));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[0]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[1]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[2]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[3]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[4]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[5]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[6]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_oe[7]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[0]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[1]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[2]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[3]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_out[4]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[5]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[6]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uio_out[7]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[0]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[1]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[2]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[3]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uo_out[4]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[5]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[6]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout37 (.A(_08812_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_08719_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_08676_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_08636_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_08075_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_08068_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_08003_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_07965_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_07929_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_07900_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_09161_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_09119_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_09098_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_09056_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_08952_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_08840_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_08720_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_08637_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_08588_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_08561_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_08466_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_08458_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_08351_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_08274_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_08200_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_08093_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_08043_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_08040_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_07590_),
    .X(net65));
 sg13g2_buf_1 fanout66 (.A(_09230_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_09211_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_09162_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_09092_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_09025_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_08985_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_08919_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_08885_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_08844_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_08804_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_08767_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_08678_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_08554_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_08529_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_08498_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_08492_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_08431_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_08392_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_08386_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_08316_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_08236_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_08141_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_08061_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_07990_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_07849_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_07785_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_10159_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_09196_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_09127_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_09121_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_08871_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_08289_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_08115_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_08083_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_07985_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_07981_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_07824_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_07784_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_07740_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_07702_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_10151_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_09090_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_09029_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_08913_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_08807_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_08552_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_08537_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_08531_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_08490_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_08421_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_08192_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_07969_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_07739_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_07701_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_10157_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_08533_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_08360_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_08235_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_08182_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_08081_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_08029_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_08008_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_07934_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_07755_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_07746_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_07665_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_09487_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_08281_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_07664_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_07610_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_07607_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_07585_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_07559_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_07547_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_07530_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_07503_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_07558_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_07546_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_05333_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_05175_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_05154_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_05134_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_05107_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_05087_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_05067_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_05048_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_05027_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_05007_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_04988_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_04817_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_04797_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_04778_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_04758_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_04717_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_04690_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_04670_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_04650_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_04631_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_04610_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_04087_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_04059_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_04038_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_04019_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_03999_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_03978_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_03959_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_03939_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_03919_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_03900_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_03880_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_03801_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_03701_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_03554_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_03533_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_03513_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_03493_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_03474_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_03454_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_03425_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_03405_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_03385_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_03366_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_03346_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_03324_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_03176_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_03156_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_03137_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_03117_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_03097_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_03078_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_03058_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_03036_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_03008_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_02988_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_02968_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_02867_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_02798_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_13042_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_13022_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_13002_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_12983_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_12963_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_12943_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_12924_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_12904_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_12883_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_12854_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_12713_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_12693_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_12672_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_12636_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_12616_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_12596_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_12576_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_12557_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_12537_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_12517_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_12498_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_12478_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_12407_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_12306_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_12286_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_12265_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_12245_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_12217_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_12198_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_12179_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_12158_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_12138_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_12119_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_12099_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_11950_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_11927_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_11907_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_11887_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_11865_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_11845_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_11826_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_11798_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_11778_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_11759_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_11739_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_11716_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_11568_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_11549_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_11529_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_11509_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_11489_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_11469_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_11448_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_11428_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_11409_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_11381_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_11361_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_11258_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_11198_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_11162_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_11142_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_11123_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_11103_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_11083_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_11063_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_11042_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_11021_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_11001_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_10982_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_10889_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_10870_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_10850_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_10829_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_10809_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_10791_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_10770_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_10742_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_10722_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_10702_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_10613_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_10545_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_10495_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_10471_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_10448_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_10426_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_10401_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_10376_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_10353_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_10329_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_10304_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_10250_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_08347_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_08294_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_08089_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_08036_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_08006_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_07947_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_05412_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_05393_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_05373_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_05353_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_05314_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_05294_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_05274_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_05255_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_05234_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_05214_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_05195_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_04965_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_04944_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_04924_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_04897_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_04877_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_04857_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_04838_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_04737_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_04508_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_04440_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_04418_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_04398_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_04378_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_04358_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_04339_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_04319_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_04299_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_04272_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_04252_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_04231_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_04206_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_04185_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_04166_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_04146_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_04126_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_04107_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_03841_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_03820_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_03781_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_03760_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_03741_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_03721_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_03680_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_03661_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_03633_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_03612_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_03592_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_03572_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_03304_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_03285_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_03265_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_03244_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_03216_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_03196_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_02945_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_02926_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_02906_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_02886_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_02847_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_02826_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_12831_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_12811_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_12791_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_12772_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_12752_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_12732_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_12453_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_12425_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_12385_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_12365_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_12345_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_12325_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_12076_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_12056_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_12037_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_12009_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_11989_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_11970_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_11696_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_11676_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_11655_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_11635_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_11616_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_11588_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_11338_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_11318_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_11298_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_11278_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_11237_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_11217_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_10949_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_10929_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_10909_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_10683_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_10660_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_10636_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_10590_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_10568_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_10517_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_08297_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_08121_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_08105_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_08060_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_08012_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_07857_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_07453_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_06106_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_06086_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_06066_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_06046_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_06027_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_06007_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_05986_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_05966_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_05946_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_05927_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_05907_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_05880_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_05857_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_05836_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_05817_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_05797_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_05776_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_05756_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_05736_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_05717_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_05695_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_05668_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_05646_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_05626_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_05607_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_05586_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_05566_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_05546_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_05524_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_05502_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_05480_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_05439_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_04586_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_04566_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_04547_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_04527_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_04479_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_04459_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_10222_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_10128_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_10098_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_09200_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_08000_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_07978_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_07856_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_07707_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_07620_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_07497_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_07313_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_04985_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_04607_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_03877_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_03343_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_02965_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_12851_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_12475_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_12096_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_11947_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_11736_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_11358_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_10979_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_10610_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_10301_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_10247_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_10199_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_10127_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_10097_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_09660_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_08389_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_08336_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_08300_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_07960_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_07640_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_07619_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_07163_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_04228_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_10211_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_10191_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_10183_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_10096_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_09772_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_08954_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_08911_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_08319_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_07751_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_07745_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_10190_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_10178_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_10165_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_10118_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_09822_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_09340_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_09156_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_09088_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_09027_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_08842_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_08631_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_08550_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_08488_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_08423_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_08135_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_07945_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_07602_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_10177_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_09339_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_09290_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_09287_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_09058_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_08353_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_08017_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_07677_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_07629_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_09280_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_08873_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_08302_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_08133_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_07568_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_07542_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_07507_),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(_10680_));
 sg13g2_buf_2 fanout527 (.A(_10657_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_10633_),
    .X(net528));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(_10233_));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(_09627_));
 sg13g2_buf_2 fanout531 (.A(_09620_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_08183_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_07561_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_07498_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_07225_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_07155_),
    .X(net536));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(_06161_));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(_06160_));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(_06158_));
 sg13g2_buf_8 fanout540 (.A(_06157_),
    .X(net540));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(_06146_));
 sg13g2_buf_8 fanout542 (.A(_06145_),
    .X(net542));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(_06143_));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(_06139_));
 sg13g2_buf_4 fanout545 (.X(net545),
    .A(_06133_));
 sg13g2_buf_2 fanout546 (.A(_06127_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_10565_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_10514_),
    .X(net548));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(_10468_));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(_10445_));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(_10423_));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(_10398_));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(_10373_));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_10350_));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(_10326_));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(_10296_));
 sg13g2_buf_2 fanout557 (.A(_10072_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_10039_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_09897_),
    .X(net559));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(_09823_));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(_09812_));
 sg13g2_buf_2 fanout562 (.A(_09645_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_09638_),
    .X(net563));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(_09626_));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(_09619_));
 sg13g2_buf_2 fanout566 (.A(_09509_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_09449_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_09418_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_09260_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_09195_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_07263_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_07188_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_07176_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_07114_),
    .X(net574));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(_06164_));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(_06163_));
 sg13g2_buf_8 fanout577 (.A(_06142_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_06138_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_05812_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_05787_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_05763_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_05739_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_05710_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_05683_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_05655_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_05629_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_05601_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_05577_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_05553_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_05527_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_05495_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_05461_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_05418_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_05387_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_05361_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_05335_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_05304_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_05278_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_05247_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_05220_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_05189_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_05162_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_05136_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_05097_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_05071_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_05040_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_05013_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_04979_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_04952_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_04926_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_04887_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_04861_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_04830_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_04803_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_04772_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_04745_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_04719_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_04680_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_04654_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_04623_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_04593_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_04569_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_04542_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_04518_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_04486_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_04460_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_04433_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_04407_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_04383_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_04359_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_04332_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_04308_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_04278_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_04247_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_04216_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_04189_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_04158_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_04132_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_04101_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_04071_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_04041_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_04009_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_03982_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_03951_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_03925_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_03894_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_03857_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_03823_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_03791_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_03764_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_03733_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_03707_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_03681_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_03652_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_03622_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_03597_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_03573_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_03544_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_03520_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_03496_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_03469_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_03442_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_03412_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_03388_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_03361_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_03334_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_03308_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_03277_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_03251_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_03210_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_03184_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_03158_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_03127_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_03101_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_03070_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_03044_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_03002_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_02976_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_02947_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_02916_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_02890_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_02859_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_02833_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_02792_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_13030_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_13004_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_12973_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_12947_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_12916_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_12890_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_12845_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_12819_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_12793_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_12762_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_12736_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_12705_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_12679_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_12630_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_12604_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_12578_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_12547_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_12521_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_12490_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_12461_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_12429_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_12398_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_12374_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_12350_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_12326_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_12299_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_12275_),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_12250_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_12218_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_12191_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_12165_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_12141_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_12114_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_12087_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_12060_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_12027_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_11995_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_11964_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_11935_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_11909_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_11877_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_11849_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_11816_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_11784_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_11753_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_11724_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_11698_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_11666_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_11639_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_11606_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_11574_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_11543_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_11517_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_11491_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_11459_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_11432_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_11399_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_11367_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_11332_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_11306_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_11280_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_11248_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_11221_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_11186_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_11148_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_11117_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_11091_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_11065_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_11032_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_11005_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_10968_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_10938_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_10914_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_10890_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_10863_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_10839_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_10814_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_10785_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_10758_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_10729_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_10705_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_10675_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_10648_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_10620_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_10592_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_10587_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_10555_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_10523_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_10492_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_10483_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_10467_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_10454_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_10417_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_10397_),
    .X(net778));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(_10349_));
 sg13g2_buf_2 fanout780 (.A(_10085_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_10080_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_10061_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_10030_),
    .X(net783));
 sg13g2_buf_4 fanout784 (.X(net784),
    .A(_09735_));
 sg13g2_buf_2 fanout785 (.A(_09723_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_09714_),
    .X(net786));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(_09625_));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(_09618_));
 sg13g2_buf_2 fanout789 (.A(_09352_),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(_09345_));
 sg13g2_buf_4 fanout791 (.X(net791),
    .A(_09214_));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(_09194_));
 sg13g2_buf_2 fanout793 (.A(_07234_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_07179_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_07178_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_07130_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_06475_));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(_06466_));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(_06420_));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(_06410_));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(_06400_));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_06393_));
 sg13g2_buf_8 fanout803 (.A(_06389_),
    .X(net803));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(_06386_));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(_06383_));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(_06380_));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(_06365_));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(_06350_));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(_06340_));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(_06336_));
 sg13g2_buf_8 fanout811 (.A(_06335_),
    .X(net811));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(_06333_));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_06322_));
 sg13g2_buf_4 fanout814 (.X(net814),
    .A(_06232_));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(_06179_));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(_06175_));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(_06155_));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(_06151_));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(_06137_));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(_06131_));
 sg13g2_buf_2 fanout821 (.A(_06097_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_06073_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_06049_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_06022_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_05997_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_05973_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_05949_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_05922_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_05895_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_05865_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_05840_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_05432_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_05171_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_04961_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_04754_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_04202_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_03995_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_03777_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_03240_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_03032_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_02822_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_12879_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_12668_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_12403_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_11903_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_11692_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_11485_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_11274_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_11059_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_10488_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_10384_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_10355_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_10314_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_10260_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_10226_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_10089_),
    .X(net856));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(_10071_));
 sg13g2_buf_2 fanout858 (.A(_10064_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_09911_),
    .X(net859));
 sg13g2_buf_4 fanout860 (.X(net860),
    .A(_09853_));
 sg13g2_buf_2 fanout861 (.A(_09746_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_09745_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_09743_),
    .X(net863));
 sg13g2_buf_4 fanout864 (.X(net864),
    .A(_09734_));
 sg13g2_buf_2 fanout865 (.A(_09732_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_09727_),
    .X(net866));
 sg13g2_buf_4 fanout867 (.X(net867),
    .A(_09713_));
 sg13g2_buf_2 fanout868 (.A(_09712_),
    .X(net868));
 sg13g2_buf_4 fanout869 (.X(net869),
    .A(_09696_));
 sg13g2_buf_2 fanout870 (.A(_09683_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_09669_),
    .X(net871));
 sg13g2_buf_4 fanout872 (.X(net872),
    .A(_09657_));
 sg13g2_buf_4 fanout873 (.X(net873),
    .A(_09624_));
 sg13g2_buf_4 fanout874 (.X(net874),
    .A(_09617_));
 sg13g2_buf_2 fanout875 (.A(_09585_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_09484_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_09478_),
    .X(net877));
 sg13g2_buf_4 fanout878 (.X(net878),
    .A(_08390_));
 sg13g2_buf_2 fanout879 (.A(_07998_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_07854_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_07743_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_07705_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_07668_),
    .X(net883));
 sg13g2_buf_8 fanout884 (.A(_06525_),
    .X(net884));
 sg13g2_buf_8 fanout885 (.A(_06497_),
    .X(net885));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(_06494_));
 sg13g2_buf_4 fanout887 (.X(net887),
    .A(_06492_));
 sg13g2_buf_4 fanout888 (.X(net888),
    .A(_06489_));
 sg13g2_buf_4 fanout889 (.X(net889),
    .A(_06487_));
 sg13g2_buf_8 fanout890 (.A(_06486_),
    .X(net890));
 sg13g2_buf_8 fanout891 (.A(_06483_),
    .X(net891));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(_06481_));
 sg13g2_buf_8 fanout893 (.A(_06480_),
    .X(net893));
 sg13g2_buf_8 fanout894 (.A(_06478_),
    .X(net894));
 sg13g2_buf_4 fanout895 (.X(net895),
    .A(_06474_));
 sg13g2_buf_8 fanout896 (.A(_06472_),
    .X(net896));
 sg13g2_buf_8 fanout897 (.A(_06470_),
    .X(net897));
 sg13g2_buf_4 fanout898 (.X(net898),
    .A(_06468_));
 sg13g2_buf_4 fanout899 (.X(net899),
    .A(_06464_));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(_06459_));
 sg13g2_buf_4 fanout901 (.X(net901),
    .A(_06456_));
 sg13g2_buf_8 fanout902 (.A(_06455_),
    .X(net902));
 sg13g2_buf_8 fanout903 (.A(_06453_),
    .X(net903));
 sg13g2_buf_4 fanout904 (.X(net904),
    .A(_06451_));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(_06449_));
 sg13g2_buf_8 fanout906 (.A(_06448_),
    .X(net906));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(_06444_));
 sg13g2_buf_8 fanout908 (.A(_06443_),
    .X(net908));
 sg13g2_buf_4 fanout909 (.X(net909),
    .A(_06441_));
 sg13g2_buf_4 fanout910 (.X(net910),
    .A(_06439_));
 sg13g2_buf_4 fanout911 (.X(net911),
    .A(_06436_));
 sg13g2_buf_4 fanout912 (.X(net912),
    .A(_06434_));
 sg13g2_buf_8 fanout913 (.A(_06433_),
    .X(net913));
 sg13g2_buf_8 fanout914 (.A(_06431_),
    .X(net914));
 sg13g2_buf_4 fanout915 (.X(net915),
    .A(_06427_));
 sg13g2_buf_8 fanout916 (.A(_06425_),
    .X(net916));
 sg13g2_buf_4 fanout917 (.X(net917),
    .A(_06423_));
 sg13g2_buf_8 fanout918 (.A(_06422_),
    .X(net918));
 sg13g2_buf_4 fanout919 (.X(net919),
    .A(_06419_));
 sg13g2_buf_8 fanout920 (.A(_06417_),
    .X(net920));
 sg13g2_buf_4 fanout921 (.X(net921),
    .A(_06412_));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(_06407_));
 sg13g2_buf_8 fanout923 (.A(_06406_),
    .X(net923));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(_06403_));
 sg13g2_buf_8 fanout925 (.A(_06402_),
    .X(net925));
 sg13g2_buf_8 fanout926 (.A(_06399_),
    .X(net926));
 sg13g2_buf_8 fanout927 (.A(_06395_),
    .X(net927));
 sg13g2_buf_8 fanout928 (.A(_06392_),
    .X(net928));
 sg13g2_buf_8 fanout929 (.A(_06385_),
    .X(net929));
 sg13g2_buf_8 fanout930 (.A(_06382_),
    .X(net930));
 sg13g2_buf_8 fanout931 (.A(_06378_),
    .X(net931));
 sg13g2_buf_4 fanout932 (.X(net932),
    .A(_06374_));
 sg13g2_buf_8 fanout933 (.A(_06373_),
    .X(net933));
 sg13g2_buf_4 fanout934 (.X(net934),
    .A(_06371_));
 sg13g2_buf_8 fanout935 (.A(_06370_),
    .X(net935));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(_06368_));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(_06367_));
 sg13g2_buf_8 fanout938 (.A(_06363_),
    .X(net938));
 sg13g2_buf_4 fanout939 (.X(net939),
    .A(_06361_));
 sg13g2_buf_8 fanout940 (.A(_06360_),
    .X(net940));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(_06358_));
 sg13g2_buf_8 fanout942 (.A(_06356_),
    .X(net942));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(_06353_));
 sg13g2_buf_8 fanout944 (.A(_06352_),
    .X(net944));
 sg13g2_buf_8 fanout945 (.A(_06349_),
    .X(net945));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(_06347_));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(_06345_));
 sg13g2_buf_8 fanout948 (.A(_06344_),
    .X(net948));
 sg13g2_buf_8 fanout949 (.A(_06342_),
    .X(net949));
 sg13g2_buf_8 fanout950 (.A(_06338_),
    .X(net950));
 sg13g2_buf_4 fanout951 (.X(net951),
    .A(_06331_));
 sg13g2_buf_8 fanout952 (.A(_06330_),
    .X(net952));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(_06328_));
 sg13g2_buf_8 fanout954 (.A(_06327_),
    .X(net954));
 sg13g2_buf_4 fanout955 (.X(net955),
    .A(_06325_));
 sg13g2_buf_8 fanout956 (.A(_06324_),
    .X(net956));
 sg13g2_buf_8 fanout957 (.A(_06321_),
    .X(net957));
 sg13g2_buf_8 fanout958 (.A(_06319_),
    .X(net958));
 sg13g2_buf_8 fanout959 (.A(_06291_),
    .X(net959));
 sg13g2_buf_4 fanout960 (.X(net960),
    .A(_06275_));
 sg13g2_buf_4 fanout961 (.X(net961),
    .A(_06273_));
 sg13g2_buf_8 fanout962 (.A(_06254_),
    .X(net962));
 sg13g2_buf_8 fanout963 (.A(_06250_),
    .X(net963));
 sg13g2_buf_4 fanout964 (.X(net964),
    .A(_06244_));
 sg13g2_buf_8 fanout965 (.A(_06238_),
    .X(net965));
 sg13g2_buf_4 fanout966 (.X(net966),
    .A(_06235_));
 sg13g2_buf_8 fanout967 (.A(_06221_),
    .X(net967));
 sg13g2_buf_4 fanout968 (.X(net968),
    .A(_06219_));
 sg13g2_buf_8 fanout969 (.A(_06218_),
    .X(net969));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(_06213_));
 sg13g2_buf_8 fanout971 (.A(_06211_),
    .X(net971));
 sg13g2_buf_4 fanout972 (.X(net972),
    .A(_06208_));
 sg13g2_buf_8 fanout973 (.A(_06207_),
    .X(net973));
 sg13g2_buf_4 fanout974 (.X(net974),
    .A(_06204_));
 sg13g2_buf_8 fanout975 (.A(_06202_),
    .X(net975));
 sg13g2_buf_4 fanout976 (.X(net976),
    .A(_06196_));
 sg13g2_buf_8 fanout977 (.A(_06195_),
    .X(net977));
 sg13g2_buf_4 fanout978 (.X(net978),
    .A(_06191_));
 sg13g2_buf_8 fanout979 (.A(_06190_),
    .X(net979));
 sg13g2_buf_4 fanout980 (.X(net980),
    .A(_06188_));
 sg13g2_buf_8 fanout981 (.A(_06186_),
    .X(net981));
 sg13g2_buf_4 fanout982 (.X(net982),
    .A(_06184_));
 sg13g2_buf_8 fanout983 (.A(_06182_),
    .X(net983));
 sg13g2_buf_8 fanout984 (.A(_06178_),
    .X(net984));
 sg13g2_buf_8 fanout985 (.A(_06173_),
    .X(net985));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(_06170_));
 sg13g2_buf_4 fanout987 (.X(net987),
    .A(_06154_));
 sg13g2_buf_4 fanout988 (.X(net988),
    .A(_06150_));
 sg13g2_buf_4 fanout989 (.X(net989),
    .A(_06136_));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(_06130_));
 sg13g2_buf_2 fanout991 (.A(_05129_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_05126_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_05123_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_05120_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_05117_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_05114_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_05111_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_05108_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_04919_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_04916_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_04913_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_04910_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_04907_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_04904_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_04901_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_04898_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_04712_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_04709_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_04706_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_04703_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_04700_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_04697_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_04694_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_04691_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_04503_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_04500_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_04497_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_04494_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_04491_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_04488_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_04484_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_04481_),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_04295_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_04292_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_04289_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_04286_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_04283_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_04280_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_04276_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_04273_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_04082_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_04079_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_04076_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_04073_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_04069_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_04066_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_04063_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_04060_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_03872_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_03868_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_03864_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_03860_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_03855_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_03851_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_03847_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_03843_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_03657_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_03654_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_03650_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_03647_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_03644_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_03641_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_03638_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_03635_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_03450_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_03447_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_03444_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_03439_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_03436_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_03433_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_03430_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_03427_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_03238_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_03235_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_03232_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_03229_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_03226_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_03223_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_03220_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_03217_),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_03030_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_03027_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(_03024_),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_03021_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_03018_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_03015_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_03012_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_03009_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_02820_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_02817_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_02814_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_02811_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(_02808_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_02805_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(_02802_),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_02799_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_12876_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(_12873_),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_12870_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_12867_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_12864_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_12861_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_12858_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_12855_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_12666_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_12662_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(_12658_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_12654_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_12650_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_12646_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_12642_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_12638_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_12449_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_12446_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_12443_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_12440_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_12437_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_12434_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_12431_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_12427_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_12241_),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_12238_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_12235_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_12232_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_12229_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_12226_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_12223_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_12220_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_12032_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(_12029_),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(_12025_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_12022_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_12019_),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(_12016_),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_12013_),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(_12010_),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(_11821_),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(_11818_),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_11814_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(_11811_),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_11808_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(_11805_),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_11802_),
    .X(net1133));
 sg13g2_buf_2 fanout1134 (.A(_11799_),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(_11611_),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(_11608_),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(_11604_),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(_11601_),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(_11598_),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(_11595_),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(_11592_),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(_11589_),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(_11404_),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(_11401_),
    .X(net1144));
 sg13g2_buf_2 fanout1145 (.A(_11397_),
    .X(net1145));
 sg13g2_buf_2 fanout1146 (.A(_11394_),
    .X(net1146));
 sg13g2_buf_2 fanout1147 (.A(_11391_),
    .X(net1147));
 sg13g2_buf_2 fanout1148 (.A(_11388_),
    .X(net1148));
 sg13g2_buf_2 fanout1149 (.A(_11385_),
    .X(net1149));
 sg13g2_buf_2 fanout1150 (.A(_11382_),
    .X(net1150));
 sg13g2_buf_2 fanout1151 (.A(_11193_),
    .X(net1151));
 sg13g2_buf_2 fanout1152 (.A(_11189_),
    .X(net1152));
 sg13g2_buf_2 fanout1153 (.A(_11184_),
    .X(net1153));
 sg13g2_buf_2 fanout1154 (.A(_11180_),
    .X(net1154));
 sg13g2_buf_2 fanout1155 (.A(_11176_),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(_11172_),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(_11168_),
    .X(net1157));
 sg13g2_buf_2 fanout1158 (.A(_11164_),
    .X(net1158));
 sg13g2_buf_2 fanout1159 (.A(_10973_),
    .X(net1159));
 sg13g2_buf_2 fanout1160 (.A(_10970_),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(_10966_),
    .X(net1161));
 sg13g2_buf_2 fanout1162 (.A(_10963_),
    .X(net1162));
 sg13g2_buf_2 fanout1163 (.A(_10960_),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(_10957_),
    .X(net1164));
 sg13g2_buf_2 fanout1165 (.A(_10954_),
    .X(net1165));
 sg13g2_buf_2 fanout1166 (.A(_10951_),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(_10766_),
    .X(net1167));
 sg13g2_buf_2 fanout1168 (.A(_10763_),
    .X(net1168));
 sg13g2_buf_2 fanout1169 (.A(_10760_),
    .X(net1169));
 sg13g2_buf_2 fanout1170 (.A(_10756_),
    .X(net1170));
 sg13g2_buf_2 fanout1171 (.A(_10753_),
    .X(net1171));
 sg13g2_buf_2 fanout1172 (.A(_10750_),
    .X(net1172));
 sg13g2_buf_2 fanout1173 (.A(_10747_),
    .X(net1173));
 sg13g2_buf_2 fanout1174 (.A(_10744_),
    .X(net1174));
 sg13g2_buf_2 fanout1175 (.A(_10540_),
    .X(net1175));
 sg13g2_buf_2 fanout1176 (.A(_10537_),
    .X(net1176));
 sg13g2_buf_2 fanout1177 (.A(_10534_),
    .X(net1177));
 sg13g2_buf_2 fanout1178 (.A(_10531_),
    .X(net1178));
 sg13g2_buf_2 fanout1179 (.A(_10528_),
    .X(net1179));
 sg13g2_buf_2 fanout1180 (.A(_10525_),
    .X(net1180));
 sg13g2_buf_2 fanout1181 (.A(_10521_),
    .X(net1181));
 sg13g2_buf_2 fanout1182 (.A(_10518_),
    .X(net1182));
 sg13g2_buf_2 fanout1183 (.A(_10289_),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(_10284_),
    .X(net1184));
 sg13g2_buf_2 fanout1185 (.A(_10279_),
    .X(net1185));
 sg13g2_buf_2 fanout1186 (.A(_10274_),
    .X(net1186));
 sg13g2_buf_2 fanout1187 (.A(_10269_),
    .X(net1187));
 sg13g2_buf_2 fanout1188 (.A(_10264_),
    .X(net1188));
 sg13g2_buf_2 fanout1189 (.A(_10258_),
    .X(net1189));
 sg13g2_buf_2 fanout1190 (.A(_10253_),
    .X(net1190));
 sg13g2_buf_2 fanout1191 (.A(_10144_),
    .X(net1191));
 sg13g2_buf_2 fanout1192 (.A(_09995_),
    .X(net1192));
 sg13g2_buf_2 fanout1193 (.A(_09985_),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(_09927_),
    .X(net1194));
 sg13g2_buf_4 fanout1195 (.X(net1195),
    .A(_09783_));
 sg13g2_buf_4 fanout1196 (.X(net1196),
    .A(_09744_));
 sg13g2_buf_2 fanout1197 (.A(_09717_),
    .X(net1197));
 sg13g2_buf_2 fanout1198 (.A(_09711_),
    .X(net1198));
 sg13g2_buf_4 fanout1199 (.X(net1199),
    .A(_09702_));
 sg13g2_buf_4 fanout1200 (.X(net1200),
    .A(_09695_));
 sg13g2_buf_4 fanout1201 (.X(net1201),
    .A(_09678_));
 sg13g2_buf_2 fanout1202 (.A(_09676_),
    .X(net1202));
 sg13g2_buf_8 fanout1203 (.A(_09664_),
    .X(net1203));
 sg13g2_buf_4 fanout1204 (.X(net1204),
    .A(_09661_));
 sg13g2_buf_2 fanout1205 (.A(_09623_),
    .X(net1205));
 sg13g2_buf_4 fanout1206 (.X(net1206),
    .A(_09616_));
 sg13g2_buf_2 fanout1207 (.A(_09273_),
    .X(net1207));
 sg13g2_buf_2 fanout1208 (.A(_08238_),
    .X(net1208));
 sg13g2_buf_2 fanout1209 (.A(_08158_),
    .X(net1209));
 sg13g2_buf_2 fanout1210 (.A(_08117_),
    .X(net1210));
 sg13g2_buf_2 fanout1211 (.A(_08111_),
    .X(net1211));
 sg13g2_buf_2 fanout1212 (.A(_08100_),
    .X(net1212));
 sg13g2_buf_2 fanout1213 (.A(_08076_),
    .X(net1213));
 sg13g2_buf_2 fanout1214 (.A(_08062_),
    .X(net1214));
 sg13g2_buf_2 fanout1215 (.A(_08005_),
    .X(net1215));
 sg13g2_buf_2 fanout1216 (.A(_07991_),
    .X(net1216));
 sg13g2_buf_2 fanout1217 (.A(_07976_),
    .X(net1217));
 sg13g2_buf_2 fanout1218 (.A(_07961_),
    .X(net1218));
 sg13g2_buf_2 fanout1219 (.A(_07930_),
    .X(net1219));
 sg13g2_buf_2 fanout1220 (.A(_07853_),
    .X(net1220));
 sg13g2_buf_2 fanout1221 (.A(_07850_),
    .X(net1221));
 sg13g2_buf_2 fanout1222 (.A(_07787_),
    .X(net1222));
 sg13g2_buf_2 fanout1223 (.A(_07742_),
    .X(net1223));
 sg13g2_buf_2 fanout1224 (.A(_07704_),
    .X(net1224));
 sg13g2_buf_2 fanout1225 (.A(_07667_),
    .X(net1225));
 sg13g2_buf_2 fanout1226 (.A(_07591_),
    .X(net1226));
 sg13g2_buf_2 fanout1227 (.A(_07101_),
    .X(net1227));
 sg13g2_buf_4 fanout1228 (.X(net1228),
    .A(_06462_));
 sg13g2_buf_8 fanout1229 (.A(_06461_),
    .X(net1229));
 sg13g2_buf_8 fanout1230 (.A(_06458_),
    .X(net1230));
 sg13g2_buf_8 fanout1231 (.A(_06446_),
    .X(net1231));
 sg13g2_buf_4 fanout1232 (.X(net1232),
    .A(_06376_));
 sg13g2_buf_4 fanout1233 (.X(net1233),
    .A(_06225_));
 sg13g2_buf_8 fanout1234 (.A(_06223_),
    .X(net1234));
 sg13g2_buf_4 fanout1235 (.X(net1235),
    .A(_06169_));
 sg13g2_buf_4 fanout1236 (.X(net1236),
    .A(_06149_));
 sg13g2_buf_2 fanout1237 (.A(_05903_),
    .X(net1237));
 sg13g2_buf_2 fanout1238 (.A(_05900_),
    .X(net1238));
 sg13g2_buf_2 fanout1239 (.A(_05897_),
    .X(net1239));
 sg13g2_buf_2 fanout1240 (.A(_05893_),
    .X(net1240));
 sg13g2_buf_2 fanout1241 (.A(_05890_),
    .X(net1241));
 sg13g2_buf_2 fanout1242 (.A(_05887_),
    .X(net1242));
 sg13g2_buf_2 fanout1243 (.A(_05882_),
    .X(net1243));
 sg13g2_buf_2 fanout1244 (.A(_05861_),
    .X(net1244));
 sg13g2_buf_2 fanout1245 (.A(_05691_),
    .X(net1245));
 sg13g2_buf_2 fanout1246 (.A(_05688_),
    .X(net1246));
 sg13g2_buf_2 fanout1247 (.A(_05685_),
    .X(net1247));
 sg13g2_buf_2 fanout1248 (.A(_05681_),
    .X(net1248));
 sg13g2_buf_2 fanout1249 (.A(_05678_),
    .X(net1249));
 sg13g2_buf_2 fanout1250 (.A(_05675_),
    .X(net1250));
 sg13g2_buf_2 fanout1251 (.A(_05670_),
    .X(net1251));
 sg13g2_buf_2 fanout1252 (.A(_05650_),
    .X(net1252));
 sg13g2_buf_2 fanout1253 (.A(_05472_),
    .X(net1253));
 sg13g2_buf_2 fanout1254 (.A(_05468_),
    .X(net1254));
 sg13g2_buf_2 fanout1255 (.A(_05464_),
    .X(net1255));
 sg13g2_buf_2 fanout1256 (.A(_05458_),
    .X(net1256));
 sg13g2_buf_2 fanout1257 (.A(_05454_),
    .X(net1257));
 sg13g2_buf_2 fanout1258 (.A(_05450_),
    .X(net1258));
 sg13g2_buf_2 fanout1259 (.A(_05446_),
    .X(net1259));
 sg13g2_buf_2 fanout1260 (.A(_05442_),
    .X(net1260));
 sg13g2_buf_2 fanout1261 (.A(_10288_),
    .X(net1261));
 sg13g2_buf_2 fanout1262 (.A(_10283_),
    .X(net1262));
 sg13g2_buf_2 fanout1263 (.A(_10278_),
    .X(net1263));
 sg13g2_buf_2 fanout1264 (.A(_10273_),
    .X(net1264));
 sg13g2_buf_2 fanout1265 (.A(_10268_),
    .X(net1265));
 sg13g2_buf_2 fanout1266 (.A(_10263_),
    .X(net1266));
 sg13g2_buf_2 fanout1267 (.A(_10257_),
    .X(net1267));
 sg13g2_buf_2 fanout1268 (.A(_10252_),
    .X(net1268));
 sg13g2_buf_2 fanout1269 (.A(_10235_),
    .X(net1269));
 sg13g2_buf_2 fanout1270 (.A(_10143_),
    .X(net1270));
 sg13g2_buf_2 fanout1271 (.A(_10112_),
    .X(net1271));
 sg13g2_buf_2 fanout1272 (.A(_10075_),
    .X(net1272));
 sg13g2_buf_4 fanout1273 (.X(net1273),
    .A(_09984_));
 sg13g2_buf_2 fanout1274 (.A(_09965_),
    .X(net1274));
 sg13g2_buf_2 fanout1275 (.A(_09914_),
    .X(net1275));
 sg13g2_buf_2 fanout1276 (.A(_09908_),
    .X(net1276));
 sg13g2_buf_2 fanout1277 (.A(_09889_),
    .X(net1277));
 sg13g2_buf_2 fanout1278 (.A(_09877_),
    .X(net1278));
 sg13g2_buf_2 fanout1279 (.A(_09677_),
    .X(net1279));
 sg13g2_buf_4 fanout1280 (.X(net1280),
    .A(_09675_));
 sg13g2_buf_2 fanout1281 (.A(_09622_),
    .X(net1281));
 sg13g2_buf_2 fanout1282 (.A(_09615_),
    .X(net1282));
 sg13g2_buf_2 fanout1283 (.A(_09548_),
    .X(net1283));
 sg13g2_buf_2 fanout1284 (.A(_09547_),
    .X(net1284));
 sg13g2_buf_2 fanout1285 (.A(_05471_),
    .X(net1285));
 sg13g2_buf_2 fanout1286 (.A(_05467_),
    .X(net1286));
 sg13g2_buf_2 fanout1287 (.A(_05463_),
    .X(net1287));
 sg13g2_buf_2 fanout1288 (.A(_05457_),
    .X(net1288));
 sg13g2_buf_2 fanout1289 (.A(_05453_),
    .X(net1289));
 sg13g2_buf_2 fanout1290 (.A(_05449_),
    .X(net1290));
 sg13g2_buf_2 fanout1291 (.A(_05445_),
    .X(net1291));
 sg13g2_buf_2 fanout1292 (.A(_05441_),
    .X(net1292));
 sg13g2_buf_2 fanout1293 (.A(_10107_),
    .X(net1293));
 sg13g2_buf_2 fanout1294 (.A(_10102_),
    .X(net1294));
 sg13g2_buf_2 fanout1295 (.A(_10092_),
    .X(net1295));
 sg13g2_buf_2 fanout1296 (.A(_10033_),
    .X(net1296));
 sg13g2_buf_2 fanout1297 (.A(_10031_),
    .X(net1297));
 sg13g2_buf_2 fanout1298 (.A(_10023_),
    .X(net1298));
 sg13g2_buf_2 fanout1299 (.A(_10021_),
    .X(net1299));
 sg13g2_buf_2 fanout1300 (.A(_10016_),
    .X(net1300));
 sg13g2_buf_2 fanout1301 (.A(_10015_),
    .X(net1301));
 sg13g2_buf_2 fanout1302 (.A(_10014_),
    .X(net1302));
 sg13g2_buf_2 fanout1303 (.A(_09923_),
    .X(net1303));
 sg13g2_buf_2 fanout1304 (.A(_09907_),
    .X(net1304));
 sg13g2_buf_2 fanout1305 (.A(_09893_),
    .X(net1305));
 sg13g2_buf_2 fanout1306 (.A(_09878_),
    .X(net1306));
 sg13g2_buf_2 fanout1307 (.A(_09871_),
    .X(net1307));
 sg13g2_buf_2 fanout1308 (.A(_09869_),
    .X(net1308));
 sg13g2_buf_2 fanout1309 (.A(_09868_),
    .X(net1309));
 sg13g2_buf_2 fanout1310 (.A(_09634_),
    .X(net1310));
 sg13g2_buf_2 fanout1311 (.A(_09621_),
    .X(net1311));
 sg13g2_tiehi _28689__1312 (.L_HI(net1312));
 sg13g2_tiehi _28690__1313 (.L_HI(net1313));
 sg13g2_tiehi _28691__1314 (.L_HI(net1314));
 sg13g2_tiehi _28692__1315 (.L_HI(net1315));
 sg13g2_tiehi _28693__1316 (.L_HI(net1316));
 sg13g2_tiehi _28694__1317 (.L_HI(net1317));
 sg13g2_tiehi _28695__1318 (.L_HI(net1318));
 sg13g2_tiehi _28696__1319 (.L_HI(net1319));
 sg13g2_tiehi \delay_counter[0]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \delay_counter[1]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \delay_counter[2]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \delay_counter[3]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \delay_counter[4]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \delay_counter[5]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \delay_counter[6]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \delay_counter[7]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \delay_cycles[0]$_SDFFE_PN0P__1328  (.L_HI(net1328));
 sg13g2_tiehi \delay_cycles[10]$_SDFFE_PN0P__1329  (.L_HI(net1329));
 sg13g2_tiehi \delay_cycles[11]$_SDFFE_PN0P__1330  (.L_HI(net1330));
 sg13g2_tiehi \delay_cycles[12]$_SDFFE_PN0P__1331  (.L_HI(net1331));
 sg13g2_tiehi \delay_cycles[13]$_SDFFE_PN0P__1332  (.L_HI(net1332));
 sg13g2_tiehi \delay_cycles[14]$_SDFFE_PN0P__1333  (.L_HI(net1333));
 sg13g2_tiehi \delay_cycles[15]$_SDFFE_PN0P__1334  (.L_HI(net1334));
 sg13g2_tiehi \delay_cycles[16]$_SDFFE_PN0P__1335  (.L_HI(net1335));
 sg13g2_tiehi \delay_cycles[17]$_SDFFE_PN0P__1336  (.L_HI(net1336));
 sg13g2_tiehi \delay_cycles[18]$_SDFFE_PN0P__1337  (.L_HI(net1337));
 sg13g2_tiehi \delay_cycles[19]$_SDFFE_PN0P__1338  (.L_HI(net1338));
 sg13g2_tiehi \delay_cycles[1]$_SDFFE_PN0P__1339  (.L_HI(net1339));
 sg13g2_tiehi \delay_cycles[20]$_SDFFE_PN0P__1340  (.L_HI(net1340));
 sg13g2_tiehi \delay_cycles[21]$_SDFFE_PN0P__1341  (.L_HI(net1341));
 sg13g2_tiehi \delay_cycles[22]$_SDFFE_PN0P__1342  (.L_HI(net1342));
 sg13g2_tiehi \delay_cycles[23]$_SDFFE_PN0P__1343  (.L_HI(net1343));
 sg13g2_tiehi \delay_cycles[2]$_SDFFE_PN0P__1344  (.L_HI(net1344));
 sg13g2_tiehi \delay_cycles[3]$_SDFFE_PN0P__1345  (.L_HI(net1345));
 sg13g2_tiehi \delay_cycles[4]$_SDFFE_PN0P__1346  (.L_HI(net1346));
 sg13g2_tiehi \delay_cycles[5]$_SDFFE_PN0P__1347  (.L_HI(net1347));
 sg13g2_tiehi \delay_cycles[6]$_SDFFE_PN0P__1348  (.L_HI(net1348));
 sg13g2_tiehi \delay_cycles[7]$_SDFFE_PN0P__1349  (.L_HI(net1349));
 sg13g2_tiehi \delay_cycles[8]$_SDFFE_PN0P__1350  (.L_HI(net1350));
 sg13g2_tiehi \delay_cycles[9]$_SDFFE_PN0P__1351  (.L_HI(net1351));
 sg13g2_tiehi \mem.mem_internal.code_mem[0][0]$_SDFFCE_PN0P__1352  (.L_HI(net1352));
 sg13g2_tiehi \mem.mem_internal.code_mem[0][1]$_SDFFCE_PN0P__1353  (.L_HI(net1353));
 sg13g2_tiehi \mem.mem_internal.code_mem[0][2]$_SDFFCE_PN0P__1354  (.L_HI(net1354));
 sg13g2_tiehi \mem.mem_internal.code_mem[0][3]$_SDFFCE_PN0P__1355  (.L_HI(net1355));
 sg13g2_tiehi \mem.mem_internal.code_mem[0][4]$_SDFFCE_PN0P__1356  (.L_HI(net1356));
 sg13g2_tiehi \mem.mem_internal.code_mem[0][5]$_SDFFCE_PN0P__1357  (.L_HI(net1357));
 sg13g2_tiehi \mem.mem_internal.code_mem[0][6]$_SDFFCE_PN0P__1358  (.L_HI(net1358));
 sg13g2_tiehi \mem.mem_internal.code_mem[0][7]$_SDFFCE_PN0P__1359  (.L_HI(net1359));
 sg13g2_tiehi \mem.mem_internal.code_mem[100][0]$_SDFFCE_PN0P__1360  (.L_HI(net1360));
 sg13g2_tiehi \mem.mem_internal.code_mem[100][1]$_SDFFCE_PN0P__1361  (.L_HI(net1361));
 sg13g2_tiehi \mem.mem_internal.code_mem[100][2]$_SDFFCE_PN0P__1362  (.L_HI(net1362));
 sg13g2_tiehi \mem.mem_internal.code_mem[100][3]$_SDFFCE_PN0P__1363  (.L_HI(net1363));
 sg13g2_tiehi \mem.mem_internal.code_mem[100][4]$_SDFFCE_PN0P__1364  (.L_HI(net1364));
 sg13g2_tiehi \mem.mem_internal.code_mem[100][5]$_SDFFCE_PN0P__1365  (.L_HI(net1365));
 sg13g2_tiehi \mem.mem_internal.code_mem[100][6]$_SDFFCE_PN0P__1366  (.L_HI(net1366));
 sg13g2_tiehi \mem.mem_internal.code_mem[100][7]$_SDFFCE_PN0P__1367  (.L_HI(net1367));
 sg13g2_tiehi \mem.mem_internal.code_mem[101][0]$_SDFFCE_PN0P__1368  (.L_HI(net1368));
 sg13g2_tiehi \mem.mem_internal.code_mem[101][1]$_SDFFCE_PN0P__1369  (.L_HI(net1369));
 sg13g2_tiehi \mem.mem_internal.code_mem[101][2]$_SDFFCE_PN0P__1370  (.L_HI(net1370));
 sg13g2_tiehi \mem.mem_internal.code_mem[101][3]$_SDFFCE_PN0P__1371  (.L_HI(net1371));
 sg13g2_tiehi \mem.mem_internal.code_mem[101][4]$_SDFFCE_PN0P__1372  (.L_HI(net1372));
 sg13g2_tiehi \mem.mem_internal.code_mem[101][5]$_SDFFCE_PN0P__1373  (.L_HI(net1373));
 sg13g2_tiehi \mem.mem_internal.code_mem[101][6]$_SDFFCE_PN0P__1374  (.L_HI(net1374));
 sg13g2_tiehi \mem.mem_internal.code_mem[101][7]$_SDFFCE_PN0P__1375  (.L_HI(net1375));
 sg13g2_tiehi \mem.mem_internal.code_mem[102][0]$_SDFFCE_PN0P__1376  (.L_HI(net1376));
 sg13g2_tiehi \mem.mem_internal.code_mem[102][1]$_SDFFCE_PN0P__1377  (.L_HI(net1377));
 sg13g2_tiehi \mem.mem_internal.code_mem[102][2]$_SDFFCE_PN0P__1378  (.L_HI(net1378));
 sg13g2_tiehi \mem.mem_internal.code_mem[102][3]$_SDFFCE_PN0P__1379  (.L_HI(net1379));
 sg13g2_tiehi \mem.mem_internal.code_mem[102][4]$_SDFFCE_PN0P__1380  (.L_HI(net1380));
 sg13g2_tiehi \mem.mem_internal.code_mem[102][5]$_SDFFCE_PN0P__1381  (.L_HI(net1381));
 sg13g2_tiehi \mem.mem_internal.code_mem[102][6]$_SDFFCE_PN0P__1382  (.L_HI(net1382));
 sg13g2_tiehi \mem.mem_internal.code_mem[102][7]$_SDFFCE_PN0P__1383  (.L_HI(net1383));
 sg13g2_tiehi \mem.mem_internal.code_mem[103][0]$_SDFFCE_PN0P__1384  (.L_HI(net1384));
 sg13g2_tiehi \mem.mem_internal.code_mem[103][1]$_SDFFCE_PN0P__1385  (.L_HI(net1385));
 sg13g2_tiehi \mem.mem_internal.code_mem[103][2]$_SDFFCE_PN0P__1386  (.L_HI(net1386));
 sg13g2_tiehi \mem.mem_internal.code_mem[103][3]$_SDFFCE_PN0P__1387  (.L_HI(net1387));
 sg13g2_tiehi \mem.mem_internal.code_mem[103][4]$_SDFFCE_PN0P__1388  (.L_HI(net1388));
 sg13g2_tiehi \mem.mem_internal.code_mem[103][5]$_SDFFCE_PN0P__1389  (.L_HI(net1389));
 sg13g2_tiehi \mem.mem_internal.code_mem[103][6]$_SDFFCE_PN0P__1390  (.L_HI(net1390));
 sg13g2_tiehi \mem.mem_internal.code_mem[103][7]$_SDFFCE_PN0P__1391  (.L_HI(net1391));
 sg13g2_tiehi \mem.mem_internal.code_mem[104][0]$_SDFFCE_PN0P__1392  (.L_HI(net1392));
 sg13g2_tiehi \mem.mem_internal.code_mem[104][1]$_SDFFCE_PN0P__1393  (.L_HI(net1393));
 sg13g2_tiehi \mem.mem_internal.code_mem[104][2]$_SDFFCE_PN0P__1394  (.L_HI(net1394));
 sg13g2_tiehi \mem.mem_internal.code_mem[104][3]$_SDFFCE_PN0P__1395  (.L_HI(net1395));
 sg13g2_tiehi \mem.mem_internal.code_mem[104][4]$_SDFFCE_PN0P__1396  (.L_HI(net1396));
 sg13g2_tiehi \mem.mem_internal.code_mem[104][5]$_SDFFCE_PN0P__1397  (.L_HI(net1397));
 sg13g2_tiehi \mem.mem_internal.code_mem[104][6]$_SDFFCE_PN0P__1398  (.L_HI(net1398));
 sg13g2_tiehi \mem.mem_internal.code_mem[104][7]$_SDFFCE_PN0P__1399  (.L_HI(net1399));
 sg13g2_tiehi \mem.mem_internal.code_mem[105][0]$_SDFFCE_PN0P__1400  (.L_HI(net1400));
 sg13g2_tiehi \mem.mem_internal.code_mem[105][1]$_SDFFCE_PN0P__1401  (.L_HI(net1401));
 sg13g2_tiehi \mem.mem_internal.code_mem[105][2]$_SDFFCE_PN0P__1402  (.L_HI(net1402));
 sg13g2_tiehi \mem.mem_internal.code_mem[105][3]$_SDFFCE_PN0P__1403  (.L_HI(net1403));
 sg13g2_tiehi \mem.mem_internal.code_mem[105][4]$_SDFFCE_PN0P__1404  (.L_HI(net1404));
 sg13g2_tiehi \mem.mem_internal.code_mem[105][5]$_SDFFCE_PN0P__1405  (.L_HI(net1405));
 sg13g2_tiehi \mem.mem_internal.code_mem[105][6]$_SDFFCE_PN0P__1406  (.L_HI(net1406));
 sg13g2_tiehi \mem.mem_internal.code_mem[105][7]$_SDFFCE_PN0P__1407  (.L_HI(net1407));
 sg13g2_tiehi \mem.mem_internal.code_mem[106][0]$_SDFFCE_PN0P__1408  (.L_HI(net1408));
 sg13g2_tiehi \mem.mem_internal.code_mem[106][1]$_SDFFCE_PN0P__1409  (.L_HI(net1409));
 sg13g2_tiehi \mem.mem_internal.code_mem[106][2]$_SDFFCE_PN0P__1410  (.L_HI(net1410));
 sg13g2_tiehi \mem.mem_internal.code_mem[106][3]$_SDFFCE_PN0P__1411  (.L_HI(net1411));
 sg13g2_tiehi \mem.mem_internal.code_mem[106][4]$_SDFFCE_PN0P__1412  (.L_HI(net1412));
 sg13g2_tiehi \mem.mem_internal.code_mem[106][5]$_SDFFCE_PN0P__1413  (.L_HI(net1413));
 sg13g2_tiehi \mem.mem_internal.code_mem[106][6]$_SDFFCE_PN0P__1414  (.L_HI(net1414));
 sg13g2_tiehi \mem.mem_internal.code_mem[106][7]$_SDFFCE_PN0P__1415  (.L_HI(net1415));
 sg13g2_tiehi \mem.mem_internal.code_mem[107][0]$_SDFFCE_PN0P__1416  (.L_HI(net1416));
 sg13g2_tiehi \mem.mem_internal.code_mem[107][1]$_SDFFCE_PN0P__1417  (.L_HI(net1417));
 sg13g2_tiehi \mem.mem_internal.code_mem[107][2]$_SDFFCE_PN0P__1418  (.L_HI(net1418));
 sg13g2_tiehi \mem.mem_internal.code_mem[107][3]$_SDFFCE_PN0P__1419  (.L_HI(net1419));
 sg13g2_tiehi \mem.mem_internal.code_mem[107][4]$_SDFFCE_PN0P__1420  (.L_HI(net1420));
 sg13g2_tiehi \mem.mem_internal.code_mem[107][5]$_SDFFCE_PN0P__1421  (.L_HI(net1421));
 sg13g2_tiehi \mem.mem_internal.code_mem[107][6]$_SDFFCE_PN0P__1422  (.L_HI(net1422));
 sg13g2_tiehi \mem.mem_internal.code_mem[107][7]$_SDFFCE_PN0P__1423  (.L_HI(net1423));
 sg13g2_tiehi \mem.mem_internal.code_mem[108][0]$_SDFFCE_PN0P__1424  (.L_HI(net1424));
 sg13g2_tiehi \mem.mem_internal.code_mem[108][1]$_SDFFCE_PN0P__1425  (.L_HI(net1425));
 sg13g2_tiehi \mem.mem_internal.code_mem[108][2]$_SDFFCE_PN0P__1426  (.L_HI(net1426));
 sg13g2_tiehi \mem.mem_internal.code_mem[108][3]$_SDFFCE_PN0P__1427  (.L_HI(net1427));
 sg13g2_tiehi \mem.mem_internal.code_mem[108][4]$_SDFFCE_PN0P__1428  (.L_HI(net1428));
 sg13g2_tiehi \mem.mem_internal.code_mem[108][5]$_SDFFCE_PN0P__1429  (.L_HI(net1429));
 sg13g2_tiehi \mem.mem_internal.code_mem[108][6]$_SDFFCE_PN0P__1430  (.L_HI(net1430));
 sg13g2_tiehi \mem.mem_internal.code_mem[108][7]$_SDFFCE_PN0P__1431  (.L_HI(net1431));
 sg13g2_tiehi \mem.mem_internal.code_mem[109][0]$_SDFFCE_PN0P__1432  (.L_HI(net1432));
 sg13g2_tiehi \mem.mem_internal.code_mem[109][1]$_SDFFCE_PN0P__1433  (.L_HI(net1433));
 sg13g2_tiehi \mem.mem_internal.code_mem[109][2]$_SDFFCE_PN0P__1434  (.L_HI(net1434));
 sg13g2_tiehi \mem.mem_internal.code_mem[109][3]$_SDFFCE_PN0P__1435  (.L_HI(net1435));
 sg13g2_tiehi \mem.mem_internal.code_mem[109][4]$_SDFFCE_PN0P__1436  (.L_HI(net1436));
 sg13g2_tiehi \mem.mem_internal.code_mem[109][5]$_SDFFCE_PN0P__1437  (.L_HI(net1437));
 sg13g2_tiehi \mem.mem_internal.code_mem[109][6]$_SDFFCE_PN0P__1438  (.L_HI(net1438));
 sg13g2_tiehi \mem.mem_internal.code_mem[109][7]$_SDFFCE_PN0P__1439  (.L_HI(net1439));
 sg13g2_tiehi \mem.mem_internal.code_mem[10][0]$_SDFFCE_PN0P__1440  (.L_HI(net1440));
 sg13g2_tiehi \mem.mem_internal.code_mem[10][1]$_SDFFCE_PN0P__1441  (.L_HI(net1441));
 sg13g2_tiehi \mem.mem_internal.code_mem[10][2]$_SDFFCE_PN0P__1442  (.L_HI(net1442));
 sg13g2_tiehi \mem.mem_internal.code_mem[10][3]$_SDFFCE_PN0P__1443  (.L_HI(net1443));
 sg13g2_tiehi \mem.mem_internal.code_mem[10][4]$_SDFFCE_PN0P__1444  (.L_HI(net1444));
 sg13g2_tiehi \mem.mem_internal.code_mem[10][5]$_SDFFCE_PN0P__1445  (.L_HI(net1445));
 sg13g2_tiehi \mem.mem_internal.code_mem[10][6]$_SDFFCE_PN0P__1446  (.L_HI(net1446));
 sg13g2_tiehi \mem.mem_internal.code_mem[10][7]$_SDFFCE_PN0P__1447  (.L_HI(net1447));
 sg13g2_tiehi \mem.mem_internal.code_mem[110][0]$_SDFFCE_PN0P__1448  (.L_HI(net1448));
 sg13g2_tiehi \mem.mem_internal.code_mem[110][1]$_SDFFCE_PN0P__1449  (.L_HI(net1449));
 sg13g2_tiehi \mem.mem_internal.code_mem[110][2]$_SDFFCE_PN0P__1450  (.L_HI(net1450));
 sg13g2_tiehi \mem.mem_internal.code_mem[110][3]$_SDFFCE_PN0P__1451  (.L_HI(net1451));
 sg13g2_tiehi \mem.mem_internal.code_mem[110][4]$_SDFFCE_PN0P__1452  (.L_HI(net1452));
 sg13g2_tiehi \mem.mem_internal.code_mem[110][5]$_SDFFCE_PN0P__1453  (.L_HI(net1453));
 sg13g2_tiehi \mem.mem_internal.code_mem[110][6]$_SDFFCE_PN0P__1454  (.L_HI(net1454));
 sg13g2_tiehi \mem.mem_internal.code_mem[110][7]$_SDFFCE_PN0P__1455  (.L_HI(net1455));
 sg13g2_tiehi \mem.mem_internal.code_mem[111][0]$_SDFFCE_PN0P__1456  (.L_HI(net1456));
 sg13g2_tiehi \mem.mem_internal.code_mem[111][1]$_SDFFCE_PN0P__1457  (.L_HI(net1457));
 sg13g2_tiehi \mem.mem_internal.code_mem[111][2]$_SDFFCE_PN0P__1458  (.L_HI(net1458));
 sg13g2_tiehi \mem.mem_internal.code_mem[111][3]$_SDFFCE_PN0P__1459  (.L_HI(net1459));
 sg13g2_tiehi \mem.mem_internal.code_mem[111][4]$_SDFFCE_PN0P__1460  (.L_HI(net1460));
 sg13g2_tiehi \mem.mem_internal.code_mem[111][5]$_SDFFCE_PN0P__1461  (.L_HI(net1461));
 sg13g2_tiehi \mem.mem_internal.code_mem[111][6]$_SDFFCE_PN0P__1462  (.L_HI(net1462));
 sg13g2_tiehi \mem.mem_internal.code_mem[111][7]$_SDFFCE_PN0P__1463  (.L_HI(net1463));
 sg13g2_tiehi \mem.mem_internal.code_mem[112][0]$_SDFFCE_PN0P__1464  (.L_HI(net1464));
 sg13g2_tiehi \mem.mem_internal.code_mem[112][1]$_SDFFCE_PN0P__1465  (.L_HI(net1465));
 sg13g2_tiehi \mem.mem_internal.code_mem[112][2]$_SDFFCE_PN0P__1466  (.L_HI(net1466));
 sg13g2_tiehi \mem.mem_internal.code_mem[112][3]$_SDFFCE_PN0P__1467  (.L_HI(net1467));
 sg13g2_tiehi \mem.mem_internal.code_mem[112][4]$_SDFFCE_PN0P__1468  (.L_HI(net1468));
 sg13g2_tiehi \mem.mem_internal.code_mem[112][5]$_SDFFCE_PN0P__1469  (.L_HI(net1469));
 sg13g2_tiehi \mem.mem_internal.code_mem[112][6]$_SDFFCE_PN0P__1470  (.L_HI(net1470));
 sg13g2_tiehi \mem.mem_internal.code_mem[112][7]$_SDFFCE_PN0P__1471  (.L_HI(net1471));
 sg13g2_tiehi \mem.mem_internal.code_mem[113][0]$_SDFFCE_PN0P__1472  (.L_HI(net1472));
 sg13g2_tiehi \mem.mem_internal.code_mem[113][1]$_SDFFCE_PN0P__1473  (.L_HI(net1473));
 sg13g2_tiehi \mem.mem_internal.code_mem[113][2]$_SDFFCE_PN0P__1474  (.L_HI(net1474));
 sg13g2_tiehi \mem.mem_internal.code_mem[113][3]$_SDFFCE_PN0P__1475  (.L_HI(net1475));
 sg13g2_tiehi \mem.mem_internal.code_mem[113][4]$_SDFFCE_PN0P__1476  (.L_HI(net1476));
 sg13g2_tiehi \mem.mem_internal.code_mem[113][5]$_SDFFCE_PN0P__1477  (.L_HI(net1477));
 sg13g2_tiehi \mem.mem_internal.code_mem[113][6]$_SDFFCE_PN0P__1478  (.L_HI(net1478));
 sg13g2_tiehi \mem.mem_internal.code_mem[113][7]$_SDFFCE_PN0P__1479  (.L_HI(net1479));
 sg13g2_tiehi \mem.mem_internal.code_mem[114][0]$_SDFFCE_PN0P__1480  (.L_HI(net1480));
 sg13g2_tiehi \mem.mem_internal.code_mem[114][1]$_SDFFCE_PN0P__1481  (.L_HI(net1481));
 sg13g2_tiehi \mem.mem_internal.code_mem[114][2]$_SDFFCE_PN0P__1482  (.L_HI(net1482));
 sg13g2_tiehi \mem.mem_internal.code_mem[114][3]$_SDFFCE_PN0P__1483  (.L_HI(net1483));
 sg13g2_tiehi \mem.mem_internal.code_mem[114][4]$_SDFFCE_PN0P__1484  (.L_HI(net1484));
 sg13g2_tiehi \mem.mem_internal.code_mem[114][5]$_SDFFCE_PN0P__1485  (.L_HI(net1485));
 sg13g2_tiehi \mem.mem_internal.code_mem[114][6]$_SDFFCE_PN0P__1486  (.L_HI(net1486));
 sg13g2_tiehi \mem.mem_internal.code_mem[114][7]$_SDFFCE_PN0P__1487  (.L_HI(net1487));
 sg13g2_tiehi \mem.mem_internal.code_mem[115][0]$_SDFFCE_PN0P__1488  (.L_HI(net1488));
 sg13g2_tiehi \mem.mem_internal.code_mem[115][1]$_SDFFCE_PN0P__1489  (.L_HI(net1489));
 sg13g2_tiehi \mem.mem_internal.code_mem[115][2]$_SDFFCE_PN0P__1490  (.L_HI(net1490));
 sg13g2_tiehi \mem.mem_internal.code_mem[115][3]$_SDFFCE_PN0P__1491  (.L_HI(net1491));
 sg13g2_tiehi \mem.mem_internal.code_mem[115][4]$_SDFFCE_PN0P__1492  (.L_HI(net1492));
 sg13g2_tiehi \mem.mem_internal.code_mem[115][5]$_SDFFCE_PN0P__1493  (.L_HI(net1493));
 sg13g2_tiehi \mem.mem_internal.code_mem[115][6]$_SDFFCE_PN0P__1494  (.L_HI(net1494));
 sg13g2_tiehi \mem.mem_internal.code_mem[115][7]$_SDFFCE_PN0P__1495  (.L_HI(net1495));
 sg13g2_tiehi \mem.mem_internal.code_mem[116][0]$_SDFFCE_PN0P__1496  (.L_HI(net1496));
 sg13g2_tiehi \mem.mem_internal.code_mem[116][1]$_SDFFCE_PN0P__1497  (.L_HI(net1497));
 sg13g2_tiehi \mem.mem_internal.code_mem[116][2]$_SDFFCE_PN0P__1498  (.L_HI(net1498));
 sg13g2_tiehi \mem.mem_internal.code_mem[116][3]$_SDFFCE_PN0P__1499  (.L_HI(net1499));
 sg13g2_tiehi \mem.mem_internal.code_mem[116][4]$_SDFFCE_PN0P__1500  (.L_HI(net1500));
 sg13g2_tiehi \mem.mem_internal.code_mem[116][5]$_SDFFCE_PN0P__1501  (.L_HI(net1501));
 sg13g2_tiehi \mem.mem_internal.code_mem[116][6]$_SDFFCE_PN0P__1502  (.L_HI(net1502));
 sg13g2_tiehi \mem.mem_internal.code_mem[116][7]$_SDFFCE_PN0P__1503  (.L_HI(net1503));
 sg13g2_tiehi \mem.mem_internal.code_mem[117][0]$_SDFFCE_PN0P__1504  (.L_HI(net1504));
 sg13g2_tiehi \mem.mem_internal.code_mem[117][1]$_SDFFCE_PN0P__1505  (.L_HI(net1505));
 sg13g2_tiehi \mem.mem_internal.code_mem[117][2]$_SDFFCE_PN0P__1506  (.L_HI(net1506));
 sg13g2_tiehi \mem.mem_internal.code_mem[117][3]$_SDFFCE_PN0P__1507  (.L_HI(net1507));
 sg13g2_tiehi \mem.mem_internal.code_mem[117][4]$_SDFFCE_PN0P__1508  (.L_HI(net1508));
 sg13g2_tiehi \mem.mem_internal.code_mem[117][5]$_SDFFCE_PN0P__1509  (.L_HI(net1509));
 sg13g2_tiehi \mem.mem_internal.code_mem[117][6]$_SDFFCE_PN0P__1510  (.L_HI(net1510));
 sg13g2_tiehi \mem.mem_internal.code_mem[117][7]$_SDFFCE_PN0P__1511  (.L_HI(net1511));
 sg13g2_tiehi \mem.mem_internal.code_mem[118][0]$_SDFFCE_PN0P__1512  (.L_HI(net1512));
 sg13g2_tiehi \mem.mem_internal.code_mem[118][1]$_SDFFCE_PN0P__1513  (.L_HI(net1513));
 sg13g2_tiehi \mem.mem_internal.code_mem[118][2]$_SDFFCE_PN0P__1514  (.L_HI(net1514));
 sg13g2_tiehi \mem.mem_internal.code_mem[118][3]$_SDFFCE_PN0P__1515  (.L_HI(net1515));
 sg13g2_tiehi \mem.mem_internal.code_mem[118][4]$_SDFFCE_PN0P__1516  (.L_HI(net1516));
 sg13g2_tiehi \mem.mem_internal.code_mem[118][5]$_SDFFCE_PN0P__1517  (.L_HI(net1517));
 sg13g2_tiehi \mem.mem_internal.code_mem[118][6]$_SDFFCE_PN0P__1518  (.L_HI(net1518));
 sg13g2_tiehi \mem.mem_internal.code_mem[118][7]$_SDFFCE_PN0P__1519  (.L_HI(net1519));
 sg13g2_tiehi \mem.mem_internal.code_mem[119][0]$_SDFFCE_PN0P__1520  (.L_HI(net1520));
 sg13g2_tiehi \mem.mem_internal.code_mem[119][1]$_SDFFCE_PN0P__1521  (.L_HI(net1521));
 sg13g2_tiehi \mem.mem_internal.code_mem[119][2]$_SDFFCE_PN0P__1522  (.L_HI(net1522));
 sg13g2_tiehi \mem.mem_internal.code_mem[119][3]$_SDFFCE_PN0P__1523  (.L_HI(net1523));
 sg13g2_tiehi \mem.mem_internal.code_mem[119][4]$_SDFFCE_PN0P__1524  (.L_HI(net1524));
 sg13g2_tiehi \mem.mem_internal.code_mem[119][5]$_SDFFCE_PN0P__1525  (.L_HI(net1525));
 sg13g2_tiehi \mem.mem_internal.code_mem[119][6]$_SDFFCE_PN0P__1526  (.L_HI(net1526));
 sg13g2_tiehi \mem.mem_internal.code_mem[119][7]$_SDFFCE_PN0P__1527  (.L_HI(net1527));
 sg13g2_tiehi \mem.mem_internal.code_mem[11][0]$_SDFFCE_PN0P__1528  (.L_HI(net1528));
 sg13g2_tiehi \mem.mem_internal.code_mem[11][1]$_SDFFCE_PN0P__1529  (.L_HI(net1529));
 sg13g2_tiehi \mem.mem_internal.code_mem[11][2]$_SDFFCE_PN0P__1530  (.L_HI(net1530));
 sg13g2_tiehi \mem.mem_internal.code_mem[11][3]$_SDFFCE_PN0P__1531  (.L_HI(net1531));
 sg13g2_tiehi \mem.mem_internal.code_mem[11][4]$_SDFFCE_PN0P__1532  (.L_HI(net1532));
 sg13g2_tiehi \mem.mem_internal.code_mem[11][5]$_SDFFCE_PN0P__1533  (.L_HI(net1533));
 sg13g2_tiehi \mem.mem_internal.code_mem[11][6]$_SDFFCE_PN0P__1534  (.L_HI(net1534));
 sg13g2_tiehi \mem.mem_internal.code_mem[11][7]$_SDFFCE_PN0P__1535  (.L_HI(net1535));
 sg13g2_tiehi \mem.mem_internal.code_mem[120][0]$_SDFFCE_PN0P__1536  (.L_HI(net1536));
 sg13g2_tiehi \mem.mem_internal.code_mem[120][1]$_SDFFCE_PN0P__1537  (.L_HI(net1537));
 sg13g2_tiehi \mem.mem_internal.code_mem[120][2]$_SDFFCE_PN0P__1538  (.L_HI(net1538));
 sg13g2_tiehi \mem.mem_internal.code_mem[120][3]$_SDFFCE_PN0P__1539  (.L_HI(net1539));
 sg13g2_tiehi \mem.mem_internal.code_mem[120][4]$_SDFFCE_PN0P__1540  (.L_HI(net1540));
 sg13g2_tiehi \mem.mem_internal.code_mem[120][5]$_SDFFCE_PN0P__1541  (.L_HI(net1541));
 sg13g2_tiehi \mem.mem_internal.code_mem[120][6]$_SDFFCE_PN0P__1542  (.L_HI(net1542));
 sg13g2_tiehi \mem.mem_internal.code_mem[120][7]$_SDFFCE_PN0P__1543  (.L_HI(net1543));
 sg13g2_tiehi \mem.mem_internal.code_mem[121][0]$_SDFFCE_PN0P__1544  (.L_HI(net1544));
 sg13g2_tiehi \mem.mem_internal.code_mem[121][1]$_SDFFCE_PN0P__1545  (.L_HI(net1545));
 sg13g2_tiehi \mem.mem_internal.code_mem[121][2]$_SDFFCE_PN0P__1546  (.L_HI(net1546));
 sg13g2_tiehi \mem.mem_internal.code_mem[121][3]$_SDFFCE_PN0P__1547  (.L_HI(net1547));
 sg13g2_tiehi \mem.mem_internal.code_mem[121][4]$_SDFFCE_PN0P__1548  (.L_HI(net1548));
 sg13g2_tiehi \mem.mem_internal.code_mem[121][5]$_SDFFCE_PN0P__1549  (.L_HI(net1549));
 sg13g2_tiehi \mem.mem_internal.code_mem[121][6]$_SDFFCE_PN0P__1550  (.L_HI(net1550));
 sg13g2_tiehi \mem.mem_internal.code_mem[121][7]$_SDFFCE_PN0P__1551  (.L_HI(net1551));
 sg13g2_tiehi \mem.mem_internal.code_mem[122][0]$_SDFFCE_PN0P__1552  (.L_HI(net1552));
 sg13g2_tiehi \mem.mem_internal.code_mem[122][1]$_SDFFCE_PN0P__1553  (.L_HI(net1553));
 sg13g2_tiehi \mem.mem_internal.code_mem[122][2]$_SDFFCE_PN0P__1554  (.L_HI(net1554));
 sg13g2_tiehi \mem.mem_internal.code_mem[122][3]$_SDFFCE_PN0P__1555  (.L_HI(net1555));
 sg13g2_tiehi \mem.mem_internal.code_mem[122][4]$_SDFFCE_PN0P__1556  (.L_HI(net1556));
 sg13g2_tiehi \mem.mem_internal.code_mem[122][5]$_SDFFCE_PN0P__1557  (.L_HI(net1557));
 sg13g2_tiehi \mem.mem_internal.code_mem[122][6]$_SDFFCE_PN0P__1558  (.L_HI(net1558));
 sg13g2_tiehi \mem.mem_internal.code_mem[122][7]$_SDFFCE_PN0P__1559  (.L_HI(net1559));
 sg13g2_tiehi \mem.mem_internal.code_mem[123][0]$_SDFFCE_PN0P__1560  (.L_HI(net1560));
 sg13g2_tiehi \mem.mem_internal.code_mem[123][1]$_SDFFCE_PN0P__1561  (.L_HI(net1561));
 sg13g2_tiehi \mem.mem_internal.code_mem[123][2]$_SDFFCE_PN0P__1562  (.L_HI(net1562));
 sg13g2_tiehi \mem.mem_internal.code_mem[123][3]$_SDFFCE_PN0P__1563  (.L_HI(net1563));
 sg13g2_tiehi \mem.mem_internal.code_mem[123][4]$_SDFFCE_PN0P__1564  (.L_HI(net1564));
 sg13g2_tiehi \mem.mem_internal.code_mem[123][5]$_SDFFCE_PN0P__1565  (.L_HI(net1565));
 sg13g2_tiehi \mem.mem_internal.code_mem[123][6]$_SDFFCE_PN0P__1566  (.L_HI(net1566));
 sg13g2_tiehi \mem.mem_internal.code_mem[123][7]$_SDFFCE_PN0P__1567  (.L_HI(net1567));
 sg13g2_tiehi \mem.mem_internal.code_mem[124][0]$_SDFFCE_PN0P__1568  (.L_HI(net1568));
 sg13g2_tiehi \mem.mem_internal.code_mem[124][1]$_SDFFCE_PN0P__1569  (.L_HI(net1569));
 sg13g2_tiehi \mem.mem_internal.code_mem[124][2]$_SDFFCE_PN0P__1570  (.L_HI(net1570));
 sg13g2_tiehi \mem.mem_internal.code_mem[124][3]$_SDFFCE_PN0P__1571  (.L_HI(net1571));
 sg13g2_tiehi \mem.mem_internal.code_mem[124][4]$_SDFFCE_PN0P__1572  (.L_HI(net1572));
 sg13g2_tiehi \mem.mem_internal.code_mem[124][5]$_SDFFCE_PN0P__1573  (.L_HI(net1573));
 sg13g2_tiehi \mem.mem_internal.code_mem[124][6]$_SDFFCE_PN0P__1574  (.L_HI(net1574));
 sg13g2_tiehi \mem.mem_internal.code_mem[124][7]$_SDFFCE_PN0P__1575  (.L_HI(net1575));
 sg13g2_tiehi \mem.mem_internal.code_mem[125][0]$_SDFFCE_PN0P__1576  (.L_HI(net1576));
 sg13g2_tiehi \mem.mem_internal.code_mem[125][1]$_SDFFCE_PN0P__1577  (.L_HI(net1577));
 sg13g2_tiehi \mem.mem_internal.code_mem[125][2]$_SDFFCE_PN0P__1578  (.L_HI(net1578));
 sg13g2_tiehi \mem.mem_internal.code_mem[125][3]$_SDFFCE_PN0P__1579  (.L_HI(net1579));
 sg13g2_tiehi \mem.mem_internal.code_mem[125][4]$_SDFFCE_PN0P__1580  (.L_HI(net1580));
 sg13g2_tiehi \mem.mem_internal.code_mem[125][5]$_SDFFCE_PN0P__1581  (.L_HI(net1581));
 sg13g2_tiehi \mem.mem_internal.code_mem[125][6]$_SDFFCE_PN0P__1582  (.L_HI(net1582));
 sg13g2_tiehi \mem.mem_internal.code_mem[125][7]$_SDFFCE_PN0P__1583  (.L_HI(net1583));
 sg13g2_tiehi \mem.mem_internal.code_mem[126][0]$_SDFFCE_PN0P__1584  (.L_HI(net1584));
 sg13g2_tiehi \mem.mem_internal.code_mem[126][1]$_SDFFCE_PN0P__1585  (.L_HI(net1585));
 sg13g2_tiehi \mem.mem_internal.code_mem[126][2]$_SDFFCE_PN0P__1586  (.L_HI(net1586));
 sg13g2_tiehi \mem.mem_internal.code_mem[126][3]$_SDFFCE_PN0P__1587  (.L_HI(net1587));
 sg13g2_tiehi \mem.mem_internal.code_mem[126][4]$_SDFFCE_PN0P__1588  (.L_HI(net1588));
 sg13g2_tiehi \mem.mem_internal.code_mem[126][5]$_SDFFCE_PN0P__1589  (.L_HI(net1589));
 sg13g2_tiehi \mem.mem_internal.code_mem[126][6]$_SDFFCE_PN0P__1590  (.L_HI(net1590));
 sg13g2_tiehi \mem.mem_internal.code_mem[126][7]$_SDFFCE_PN0P__1591  (.L_HI(net1591));
 sg13g2_tiehi \mem.mem_internal.code_mem[127][0]$_SDFFCE_PN0P__1592  (.L_HI(net1592));
 sg13g2_tiehi \mem.mem_internal.code_mem[127][1]$_SDFFCE_PN0P__1593  (.L_HI(net1593));
 sg13g2_tiehi \mem.mem_internal.code_mem[127][2]$_SDFFCE_PN0P__1594  (.L_HI(net1594));
 sg13g2_tiehi \mem.mem_internal.code_mem[127][3]$_SDFFCE_PN0P__1595  (.L_HI(net1595));
 sg13g2_tiehi \mem.mem_internal.code_mem[127][4]$_SDFFCE_PN0P__1596  (.L_HI(net1596));
 sg13g2_tiehi \mem.mem_internal.code_mem[127][5]$_SDFFCE_PN0P__1597  (.L_HI(net1597));
 sg13g2_tiehi \mem.mem_internal.code_mem[127][6]$_SDFFCE_PN0P__1598  (.L_HI(net1598));
 sg13g2_tiehi \mem.mem_internal.code_mem[127][7]$_SDFFCE_PN0P__1599  (.L_HI(net1599));
 sg13g2_tiehi \mem.mem_internal.code_mem[128][0]$_SDFFCE_PN0P__1600  (.L_HI(net1600));
 sg13g2_tiehi \mem.mem_internal.code_mem[128][1]$_SDFFCE_PN0P__1601  (.L_HI(net1601));
 sg13g2_tiehi \mem.mem_internal.code_mem[128][2]$_SDFFCE_PN0P__1602  (.L_HI(net1602));
 sg13g2_tiehi \mem.mem_internal.code_mem[128][3]$_SDFFCE_PN0P__1603  (.L_HI(net1603));
 sg13g2_tiehi \mem.mem_internal.code_mem[128][4]$_SDFFCE_PN0P__1604  (.L_HI(net1604));
 sg13g2_tiehi \mem.mem_internal.code_mem[128][5]$_SDFFCE_PN0P__1605  (.L_HI(net1605));
 sg13g2_tiehi \mem.mem_internal.code_mem[128][6]$_SDFFCE_PN0P__1606  (.L_HI(net1606));
 sg13g2_tiehi \mem.mem_internal.code_mem[128][7]$_SDFFCE_PN0P__1607  (.L_HI(net1607));
 sg13g2_tiehi \mem.mem_internal.code_mem[129][0]$_SDFFCE_PN0P__1608  (.L_HI(net1608));
 sg13g2_tiehi \mem.mem_internal.code_mem[129][1]$_SDFFCE_PN0P__1609  (.L_HI(net1609));
 sg13g2_tiehi \mem.mem_internal.code_mem[129][2]$_SDFFCE_PN0P__1610  (.L_HI(net1610));
 sg13g2_tiehi \mem.mem_internal.code_mem[129][3]$_SDFFCE_PN0P__1611  (.L_HI(net1611));
 sg13g2_tiehi \mem.mem_internal.code_mem[129][4]$_SDFFCE_PN0P__1612  (.L_HI(net1612));
 sg13g2_tiehi \mem.mem_internal.code_mem[129][5]$_SDFFCE_PN0P__1613  (.L_HI(net1613));
 sg13g2_tiehi \mem.mem_internal.code_mem[129][6]$_SDFFCE_PN0P__1614  (.L_HI(net1614));
 sg13g2_tiehi \mem.mem_internal.code_mem[129][7]$_SDFFCE_PN0P__1615  (.L_HI(net1615));
 sg13g2_tiehi \mem.mem_internal.code_mem[12][0]$_SDFFCE_PN0P__1616  (.L_HI(net1616));
 sg13g2_tiehi \mem.mem_internal.code_mem[12][1]$_SDFFCE_PN0P__1617  (.L_HI(net1617));
 sg13g2_tiehi \mem.mem_internal.code_mem[12][2]$_SDFFCE_PN0P__1618  (.L_HI(net1618));
 sg13g2_tiehi \mem.mem_internal.code_mem[12][3]$_SDFFCE_PN0P__1619  (.L_HI(net1619));
 sg13g2_tiehi \mem.mem_internal.code_mem[12][4]$_SDFFCE_PN0P__1620  (.L_HI(net1620));
 sg13g2_tiehi \mem.mem_internal.code_mem[12][5]$_SDFFCE_PN0P__1621  (.L_HI(net1621));
 sg13g2_tiehi \mem.mem_internal.code_mem[12][6]$_SDFFCE_PN0P__1622  (.L_HI(net1622));
 sg13g2_tiehi \mem.mem_internal.code_mem[12][7]$_SDFFCE_PN0P__1623  (.L_HI(net1623));
 sg13g2_tiehi \mem.mem_internal.code_mem[130][0]$_SDFFCE_PN0P__1624  (.L_HI(net1624));
 sg13g2_tiehi \mem.mem_internal.code_mem[130][1]$_SDFFCE_PN0P__1625  (.L_HI(net1625));
 sg13g2_tiehi \mem.mem_internal.code_mem[130][2]$_SDFFCE_PN0P__1626  (.L_HI(net1626));
 sg13g2_tiehi \mem.mem_internal.code_mem[130][3]$_SDFFCE_PN0P__1627  (.L_HI(net1627));
 sg13g2_tiehi \mem.mem_internal.code_mem[130][4]$_SDFFCE_PN0P__1628  (.L_HI(net1628));
 sg13g2_tiehi \mem.mem_internal.code_mem[130][5]$_SDFFCE_PN0P__1629  (.L_HI(net1629));
 sg13g2_tiehi \mem.mem_internal.code_mem[130][6]$_SDFFCE_PN0P__1630  (.L_HI(net1630));
 sg13g2_tiehi \mem.mem_internal.code_mem[130][7]$_SDFFCE_PN0P__1631  (.L_HI(net1631));
 sg13g2_tiehi \mem.mem_internal.code_mem[131][0]$_SDFFCE_PN0P__1632  (.L_HI(net1632));
 sg13g2_tiehi \mem.mem_internal.code_mem[131][1]$_SDFFCE_PN0P__1633  (.L_HI(net1633));
 sg13g2_tiehi \mem.mem_internal.code_mem[131][2]$_SDFFCE_PN0P__1634  (.L_HI(net1634));
 sg13g2_tiehi \mem.mem_internal.code_mem[131][3]$_SDFFCE_PN0P__1635  (.L_HI(net1635));
 sg13g2_tiehi \mem.mem_internal.code_mem[131][4]$_SDFFCE_PN0P__1636  (.L_HI(net1636));
 sg13g2_tiehi \mem.mem_internal.code_mem[131][5]$_SDFFCE_PN0P__1637  (.L_HI(net1637));
 sg13g2_tiehi \mem.mem_internal.code_mem[131][6]$_SDFFCE_PN0P__1638  (.L_HI(net1638));
 sg13g2_tiehi \mem.mem_internal.code_mem[131][7]$_SDFFCE_PN0P__1639  (.L_HI(net1639));
 sg13g2_tiehi \mem.mem_internal.code_mem[132][0]$_SDFFCE_PN0P__1640  (.L_HI(net1640));
 sg13g2_tiehi \mem.mem_internal.code_mem[132][1]$_SDFFCE_PN0P__1641  (.L_HI(net1641));
 sg13g2_tiehi \mem.mem_internal.code_mem[132][2]$_SDFFCE_PN0P__1642  (.L_HI(net1642));
 sg13g2_tiehi \mem.mem_internal.code_mem[132][3]$_SDFFCE_PN0P__1643  (.L_HI(net1643));
 sg13g2_tiehi \mem.mem_internal.code_mem[132][4]$_SDFFCE_PN0P__1644  (.L_HI(net1644));
 sg13g2_tiehi \mem.mem_internal.code_mem[132][5]$_SDFFCE_PN0P__1645  (.L_HI(net1645));
 sg13g2_tiehi \mem.mem_internal.code_mem[132][6]$_SDFFCE_PN0P__1646  (.L_HI(net1646));
 sg13g2_tiehi \mem.mem_internal.code_mem[132][7]$_SDFFCE_PN0P__1647  (.L_HI(net1647));
 sg13g2_tiehi \mem.mem_internal.code_mem[133][0]$_SDFFCE_PN0P__1648  (.L_HI(net1648));
 sg13g2_tiehi \mem.mem_internal.code_mem[133][1]$_SDFFCE_PN0P__1649  (.L_HI(net1649));
 sg13g2_tiehi \mem.mem_internal.code_mem[133][2]$_SDFFCE_PN0P__1650  (.L_HI(net1650));
 sg13g2_tiehi \mem.mem_internal.code_mem[133][3]$_SDFFCE_PN0P__1651  (.L_HI(net1651));
 sg13g2_tiehi \mem.mem_internal.code_mem[133][4]$_SDFFCE_PN0P__1652  (.L_HI(net1652));
 sg13g2_tiehi \mem.mem_internal.code_mem[133][5]$_SDFFCE_PN0P__1653  (.L_HI(net1653));
 sg13g2_tiehi \mem.mem_internal.code_mem[133][6]$_SDFFCE_PN0P__1654  (.L_HI(net1654));
 sg13g2_tiehi \mem.mem_internal.code_mem[133][7]$_SDFFCE_PN0P__1655  (.L_HI(net1655));
 sg13g2_tiehi \mem.mem_internal.code_mem[134][0]$_SDFFCE_PN0P__1656  (.L_HI(net1656));
 sg13g2_tiehi \mem.mem_internal.code_mem[134][1]$_SDFFCE_PN0P__1657  (.L_HI(net1657));
 sg13g2_tiehi \mem.mem_internal.code_mem[134][2]$_SDFFCE_PN0P__1658  (.L_HI(net1658));
 sg13g2_tiehi \mem.mem_internal.code_mem[134][3]$_SDFFCE_PN0P__1659  (.L_HI(net1659));
 sg13g2_tiehi \mem.mem_internal.code_mem[134][4]$_SDFFCE_PN0P__1660  (.L_HI(net1660));
 sg13g2_tiehi \mem.mem_internal.code_mem[134][5]$_SDFFCE_PN0P__1661  (.L_HI(net1661));
 sg13g2_tiehi \mem.mem_internal.code_mem[134][6]$_SDFFCE_PN0P__1662  (.L_HI(net1662));
 sg13g2_tiehi \mem.mem_internal.code_mem[134][7]$_SDFFCE_PN0P__1663  (.L_HI(net1663));
 sg13g2_tiehi \mem.mem_internal.code_mem[135][0]$_SDFFCE_PN0P__1664  (.L_HI(net1664));
 sg13g2_tiehi \mem.mem_internal.code_mem[135][1]$_SDFFCE_PN0P__1665  (.L_HI(net1665));
 sg13g2_tiehi \mem.mem_internal.code_mem[135][2]$_SDFFCE_PN0P__1666  (.L_HI(net1666));
 sg13g2_tiehi \mem.mem_internal.code_mem[135][3]$_SDFFCE_PN0P__1667  (.L_HI(net1667));
 sg13g2_tiehi \mem.mem_internal.code_mem[135][4]$_SDFFCE_PN0P__1668  (.L_HI(net1668));
 sg13g2_tiehi \mem.mem_internal.code_mem[135][5]$_SDFFCE_PN0P__1669  (.L_HI(net1669));
 sg13g2_tiehi \mem.mem_internal.code_mem[135][6]$_SDFFCE_PN0P__1670  (.L_HI(net1670));
 sg13g2_tiehi \mem.mem_internal.code_mem[135][7]$_SDFFCE_PN0P__1671  (.L_HI(net1671));
 sg13g2_tiehi \mem.mem_internal.code_mem[136][0]$_SDFFCE_PN0P__1672  (.L_HI(net1672));
 sg13g2_tiehi \mem.mem_internal.code_mem[136][1]$_SDFFCE_PN0P__1673  (.L_HI(net1673));
 sg13g2_tiehi \mem.mem_internal.code_mem[136][2]$_SDFFCE_PN0P__1674  (.L_HI(net1674));
 sg13g2_tiehi \mem.mem_internal.code_mem[136][3]$_SDFFCE_PN0P__1675  (.L_HI(net1675));
 sg13g2_tiehi \mem.mem_internal.code_mem[136][4]$_SDFFCE_PN0P__1676  (.L_HI(net1676));
 sg13g2_tiehi \mem.mem_internal.code_mem[136][5]$_SDFFCE_PN0P__1677  (.L_HI(net1677));
 sg13g2_tiehi \mem.mem_internal.code_mem[136][6]$_SDFFCE_PN0P__1678  (.L_HI(net1678));
 sg13g2_tiehi \mem.mem_internal.code_mem[136][7]$_SDFFCE_PN0P__1679  (.L_HI(net1679));
 sg13g2_tiehi \mem.mem_internal.code_mem[137][0]$_SDFFCE_PN0P__1680  (.L_HI(net1680));
 sg13g2_tiehi \mem.mem_internal.code_mem[137][1]$_SDFFCE_PN0P__1681  (.L_HI(net1681));
 sg13g2_tiehi \mem.mem_internal.code_mem[137][2]$_SDFFCE_PN0P__1682  (.L_HI(net1682));
 sg13g2_tiehi \mem.mem_internal.code_mem[137][3]$_SDFFCE_PN0P__1683  (.L_HI(net1683));
 sg13g2_tiehi \mem.mem_internal.code_mem[137][4]$_SDFFCE_PN0P__1684  (.L_HI(net1684));
 sg13g2_tiehi \mem.mem_internal.code_mem[137][5]$_SDFFCE_PN0P__1685  (.L_HI(net1685));
 sg13g2_tiehi \mem.mem_internal.code_mem[137][6]$_SDFFCE_PN0P__1686  (.L_HI(net1686));
 sg13g2_tiehi \mem.mem_internal.code_mem[137][7]$_SDFFCE_PN0P__1687  (.L_HI(net1687));
 sg13g2_tiehi \mem.mem_internal.code_mem[138][0]$_SDFFCE_PN0P__1688  (.L_HI(net1688));
 sg13g2_tiehi \mem.mem_internal.code_mem[138][1]$_SDFFCE_PN0P__1689  (.L_HI(net1689));
 sg13g2_tiehi \mem.mem_internal.code_mem[138][2]$_SDFFCE_PN0P__1690  (.L_HI(net1690));
 sg13g2_tiehi \mem.mem_internal.code_mem[138][3]$_SDFFCE_PN0P__1691  (.L_HI(net1691));
 sg13g2_tiehi \mem.mem_internal.code_mem[138][4]$_SDFFCE_PN0P__1692  (.L_HI(net1692));
 sg13g2_tiehi \mem.mem_internal.code_mem[138][5]$_SDFFCE_PN0P__1693  (.L_HI(net1693));
 sg13g2_tiehi \mem.mem_internal.code_mem[138][6]$_SDFFCE_PN0P__1694  (.L_HI(net1694));
 sg13g2_tiehi \mem.mem_internal.code_mem[138][7]$_SDFFCE_PN0P__1695  (.L_HI(net1695));
 sg13g2_tiehi \mem.mem_internal.code_mem[139][0]$_SDFFCE_PN0P__1696  (.L_HI(net1696));
 sg13g2_tiehi \mem.mem_internal.code_mem[139][1]$_SDFFCE_PN0P__1697  (.L_HI(net1697));
 sg13g2_tiehi \mem.mem_internal.code_mem[139][2]$_SDFFCE_PN0P__1698  (.L_HI(net1698));
 sg13g2_tiehi \mem.mem_internal.code_mem[139][3]$_SDFFCE_PN0P__1699  (.L_HI(net1699));
 sg13g2_tiehi \mem.mem_internal.code_mem[139][4]$_SDFFCE_PN0P__1700  (.L_HI(net1700));
 sg13g2_tiehi \mem.mem_internal.code_mem[139][5]$_SDFFCE_PN0P__1701  (.L_HI(net1701));
 sg13g2_tiehi \mem.mem_internal.code_mem[139][6]$_SDFFCE_PN0P__1702  (.L_HI(net1702));
 sg13g2_tiehi \mem.mem_internal.code_mem[139][7]$_SDFFCE_PN0P__1703  (.L_HI(net1703));
 sg13g2_tiehi \mem.mem_internal.code_mem[13][0]$_SDFFCE_PN0P__1704  (.L_HI(net1704));
 sg13g2_tiehi \mem.mem_internal.code_mem[13][1]$_SDFFCE_PN0P__1705  (.L_HI(net1705));
 sg13g2_tiehi \mem.mem_internal.code_mem[13][2]$_SDFFCE_PN0P__1706  (.L_HI(net1706));
 sg13g2_tiehi \mem.mem_internal.code_mem[13][3]$_SDFFCE_PN0P__1707  (.L_HI(net1707));
 sg13g2_tiehi \mem.mem_internal.code_mem[13][4]$_SDFFCE_PN0P__1708  (.L_HI(net1708));
 sg13g2_tiehi \mem.mem_internal.code_mem[13][5]$_SDFFCE_PN0P__1709  (.L_HI(net1709));
 sg13g2_tiehi \mem.mem_internal.code_mem[13][6]$_SDFFCE_PN0P__1710  (.L_HI(net1710));
 sg13g2_tiehi \mem.mem_internal.code_mem[13][7]$_SDFFCE_PN0P__1711  (.L_HI(net1711));
 sg13g2_tiehi \mem.mem_internal.code_mem[140][0]$_SDFFCE_PN0P__1712  (.L_HI(net1712));
 sg13g2_tiehi \mem.mem_internal.code_mem[140][1]$_SDFFCE_PN0P__1713  (.L_HI(net1713));
 sg13g2_tiehi \mem.mem_internal.code_mem[140][2]$_SDFFCE_PN0P__1714  (.L_HI(net1714));
 sg13g2_tiehi \mem.mem_internal.code_mem[140][3]$_SDFFCE_PN0P__1715  (.L_HI(net1715));
 sg13g2_tiehi \mem.mem_internal.code_mem[140][4]$_SDFFCE_PN0P__1716  (.L_HI(net1716));
 sg13g2_tiehi \mem.mem_internal.code_mem[140][5]$_SDFFCE_PN0P__1717  (.L_HI(net1717));
 sg13g2_tiehi \mem.mem_internal.code_mem[140][6]$_SDFFCE_PN0P__1718  (.L_HI(net1718));
 sg13g2_tiehi \mem.mem_internal.code_mem[140][7]$_SDFFCE_PN0P__1719  (.L_HI(net1719));
 sg13g2_tiehi \mem.mem_internal.code_mem[141][0]$_SDFFCE_PN0P__1720  (.L_HI(net1720));
 sg13g2_tiehi \mem.mem_internal.code_mem[141][1]$_SDFFCE_PN0P__1721  (.L_HI(net1721));
 sg13g2_tiehi \mem.mem_internal.code_mem[141][2]$_SDFFCE_PN0P__1722  (.L_HI(net1722));
 sg13g2_tiehi \mem.mem_internal.code_mem[141][3]$_SDFFCE_PN0P__1723  (.L_HI(net1723));
 sg13g2_tiehi \mem.mem_internal.code_mem[141][4]$_SDFFCE_PN0P__1724  (.L_HI(net1724));
 sg13g2_tiehi \mem.mem_internal.code_mem[141][5]$_SDFFCE_PN0P__1725  (.L_HI(net1725));
 sg13g2_tiehi \mem.mem_internal.code_mem[141][6]$_SDFFCE_PN0P__1726  (.L_HI(net1726));
 sg13g2_tiehi \mem.mem_internal.code_mem[141][7]$_SDFFCE_PN0P__1727  (.L_HI(net1727));
 sg13g2_tiehi \mem.mem_internal.code_mem[142][0]$_SDFFCE_PN0P__1728  (.L_HI(net1728));
 sg13g2_tiehi \mem.mem_internal.code_mem[142][1]$_SDFFCE_PN0P__1729  (.L_HI(net1729));
 sg13g2_tiehi \mem.mem_internal.code_mem[142][2]$_SDFFCE_PN0P__1730  (.L_HI(net1730));
 sg13g2_tiehi \mem.mem_internal.code_mem[142][3]$_SDFFCE_PN0P__1731  (.L_HI(net1731));
 sg13g2_tiehi \mem.mem_internal.code_mem[142][4]$_SDFFCE_PN0P__1732  (.L_HI(net1732));
 sg13g2_tiehi \mem.mem_internal.code_mem[142][5]$_SDFFCE_PN0P__1733  (.L_HI(net1733));
 sg13g2_tiehi \mem.mem_internal.code_mem[142][6]$_SDFFCE_PN0P__1734  (.L_HI(net1734));
 sg13g2_tiehi \mem.mem_internal.code_mem[142][7]$_SDFFCE_PN0P__1735  (.L_HI(net1735));
 sg13g2_tiehi \mem.mem_internal.code_mem[143][0]$_SDFFCE_PN0P__1736  (.L_HI(net1736));
 sg13g2_tiehi \mem.mem_internal.code_mem[143][1]$_SDFFCE_PN0P__1737  (.L_HI(net1737));
 sg13g2_tiehi \mem.mem_internal.code_mem[143][2]$_SDFFCE_PN0P__1738  (.L_HI(net1738));
 sg13g2_tiehi \mem.mem_internal.code_mem[143][3]$_SDFFCE_PN0P__1739  (.L_HI(net1739));
 sg13g2_tiehi \mem.mem_internal.code_mem[143][4]$_SDFFCE_PN0P__1740  (.L_HI(net1740));
 sg13g2_tiehi \mem.mem_internal.code_mem[143][5]$_SDFFCE_PN0P__1741  (.L_HI(net1741));
 sg13g2_tiehi \mem.mem_internal.code_mem[143][6]$_SDFFCE_PN0P__1742  (.L_HI(net1742));
 sg13g2_tiehi \mem.mem_internal.code_mem[143][7]$_SDFFCE_PN0P__1743  (.L_HI(net1743));
 sg13g2_tiehi \mem.mem_internal.code_mem[144][0]$_SDFFCE_PN0P__1744  (.L_HI(net1744));
 sg13g2_tiehi \mem.mem_internal.code_mem[144][1]$_SDFFCE_PN0P__1745  (.L_HI(net1745));
 sg13g2_tiehi \mem.mem_internal.code_mem[144][2]$_SDFFCE_PN0P__1746  (.L_HI(net1746));
 sg13g2_tiehi \mem.mem_internal.code_mem[144][3]$_SDFFCE_PN0P__1747  (.L_HI(net1747));
 sg13g2_tiehi \mem.mem_internal.code_mem[144][4]$_SDFFCE_PN0P__1748  (.L_HI(net1748));
 sg13g2_tiehi \mem.mem_internal.code_mem[144][5]$_SDFFCE_PN0P__1749  (.L_HI(net1749));
 sg13g2_tiehi \mem.mem_internal.code_mem[144][6]$_SDFFCE_PN0P__1750  (.L_HI(net1750));
 sg13g2_tiehi \mem.mem_internal.code_mem[144][7]$_SDFFCE_PN0P__1751  (.L_HI(net1751));
 sg13g2_tiehi \mem.mem_internal.code_mem[145][0]$_SDFFCE_PN0P__1752  (.L_HI(net1752));
 sg13g2_tiehi \mem.mem_internal.code_mem[145][1]$_SDFFCE_PN0P__1753  (.L_HI(net1753));
 sg13g2_tiehi \mem.mem_internal.code_mem[145][2]$_SDFFCE_PN0P__1754  (.L_HI(net1754));
 sg13g2_tiehi \mem.mem_internal.code_mem[145][3]$_SDFFCE_PN0P__1755  (.L_HI(net1755));
 sg13g2_tiehi \mem.mem_internal.code_mem[145][4]$_SDFFCE_PN0P__1756  (.L_HI(net1756));
 sg13g2_tiehi \mem.mem_internal.code_mem[145][5]$_SDFFCE_PN0P__1757  (.L_HI(net1757));
 sg13g2_tiehi \mem.mem_internal.code_mem[145][6]$_SDFFCE_PN0P__1758  (.L_HI(net1758));
 sg13g2_tiehi \mem.mem_internal.code_mem[145][7]$_SDFFCE_PN0P__1759  (.L_HI(net1759));
 sg13g2_tiehi \mem.mem_internal.code_mem[146][0]$_SDFFCE_PN0P__1760  (.L_HI(net1760));
 sg13g2_tiehi \mem.mem_internal.code_mem[146][1]$_SDFFCE_PN0P__1761  (.L_HI(net1761));
 sg13g2_tiehi \mem.mem_internal.code_mem[146][2]$_SDFFCE_PN0P__1762  (.L_HI(net1762));
 sg13g2_tiehi \mem.mem_internal.code_mem[146][3]$_SDFFCE_PN0P__1763  (.L_HI(net1763));
 sg13g2_tiehi \mem.mem_internal.code_mem[146][4]$_SDFFCE_PN0P__1764  (.L_HI(net1764));
 sg13g2_tiehi \mem.mem_internal.code_mem[146][5]$_SDFFCE_PN0P__1765  (.L_HI(net1765));
 sg13g2_tiehi \mem.mem_internal.code_mem[146][6]$_SDFFCE_PN0P__1766  (.L_HI(net1766));
 sg13g2_tiehi \mem.mem_internal.code_mem[146][7]$_SDFFCE_PN0P__1767  (.L_HI(net1767));
 sg13g2_tiehi \mem.mem_internal.code_mem[147][0]$_SDFFCE_PN0P__1768  (.L_HI(net1768));
 sg13g2_tiehi \mem.mem_internal.code_mem[147][1]$_SDFFCE_PN0P__1769  (.L_HI(net1769));
 sg13g2_tiehi \mem.mem_internal.code_mem[147][2]$_SDFFCE_PN0P__1770  (.L_HI(net1770));
 sg13g2_tiehi \mem.mem_internal.code_mem[147][3]$_SDFFCE_PN0P__1771  (.L_HI(net1771));
 sg13g2_tiehi \mem.mem_internal.code_mem[147][4]$_SDFFCE_PN0P__1772  (.L_HI(net1772));
 sg13g2_tiehi \mem.mem_internal.code_mem[147][5]$_SDFFCE_PN0P__1773  (.L_HI(net1773));
 sg13g2_tiehi \mem.mem_internal.code_mem[147][6]$_SDFFCE_PN0P__1774  (.L_HI(net1774));
 sg13g2_tiehi \mem.mem_internal.code_mem[147][7]$_SDFFCE_PN0P__1775  (.L_HI(net1775));
 sg13g2_tiehi \mem.mem_internal.code_mem[148][0]$_SDFFCE_PN0P__1776  (.L_HI(net1776));
 sg13g2_tiehi \mem.mem_internal.code_mem[148][1]$_SDFFCE_PN0P__1777  (.L_HI(net1777));
 sg13g2_tiehi \mem.mem_internal.code_mem[148][2]$_SDFFCE_PN0P__1778  (.L_HI(net1778));
 sg13g2_tiehi \mem.mem_internal.code_mem[148][3]$_SDFFCE_PN0P__1779  (.L_HI(net1779));
 sg13g2_tiehi \mem.mem_internal.code_mem[148][4]$_SDFFCE_PN0P__1780  (.L_HI(net1780));
 sg13g2_tiehi \mem.mem_internal.code_mem[148][5]$_SDFFCE_PN0P__1781  (.L_HI(net1781));
 sg13g2_tiehi \mem.mem_internal.code_mem[148][6]$_SDFFCE_PN0P__1782  (.L_HI(net1782));
 sg13g2_tiehi \mem.mem_internal.code_mem[148][7]$_SDFFCE_PN0P__1783  (.L_HI(net1783));
 sg13g2_tiehi \mem.mem_internal.code_mem[149][0]$_SDFFCE_PN0P__1784  (.L_HI(net1784));
 sg13g2_tiehi \mem.mem_internal.code_mem[149][1]$_SDFFCE_PN0P__1785  (.L_HI(net1785));
 sg13g2_tiehi \mem.mem_internal.code_mem[149][2]$_SDFFCE_PN0P__1786  (.L_HI(net1786));
 sg13g2_tiehi \mem.mem_internal.code_mem[149][3]$_SDFFCE_PN0P__1787  (.L_HI(net1787));
 sg13g2_tiehi \mem.mem_internal.code_mem[149][4]$_SDFFCE_PN0P__1788  (.L_HI(net1788));
 sg13g2_tiehi \mem.mem_internal.code_mem[149][5]$_SDFFCE_PN0P__1789  (.L_HI(net1789));
 sg13g2_tiehi \mem.mem_internal.code_mem[149][6]$_SDFFCE_PN0P__1790  (.L_HI(net1790));
 sg13g2_tiehi \mem.mem_internal.code_mem[149][7]$_SDFFCE_PN0P__1791  (.L_HI(net1791));
 sg13g2_tiehi \mem.mem_internal.code_mem[14][0]$_SDFFCE_PN0P__1792  (.L_HI(net1792));
 sg13g2_tiehi \mem.mem_internal.code_mem[14][1]$_SDFFCE_PN0P__1793  (.L_HI(net1793));
 sg13g2_tiehi \mem.mem_internal.code_mem[14][2]$_SDFFCE_PN0P__1794  (.L_HI(net1794));
 sg13g2_tiehi \mem.mem_internal.code_mem[14][3]$_SDFFCE_PN0P__1795  (.L_HI(net1795));
 sg13g2_tiehi \mem.mem_internal.code_mem[14][4]$_SDFFCE_PN0P__1796  (.L_HI(net1796));
 sg13g2_tiehi \mem.mem_internal.code_mem[14][5]$_SDFFCE_PN0P__1797  (.L_HI(net1797));
 sg13g2_tiehi \mem.mem_internal.code_mem[14][6]$_SDFFCE_PN0P__1798  (.L_HI(net1798));
 sg13g2_tiehi \mem.mem_internal.code_mem[14][7]$_SDFFCE_PN0P__1799  (.L_HI(net1799));
 sg13g2_tiehi \mem.mem_internal.code_mem[150][0]$_SDFFCE_PN0P__1800  (.L_HI(net1800));
 sg13g2_tiehi \mem.mem_internal.code_mem[150][1]$_SDFFCE_PN0P__1801  (.L_HI(net1801));
 sg13g2_tiehi \mem.mem_internal.code_mem[150][2]$_SDFFCE_PN0P__1802  (.L_HI(net1802));
 sg13g2_tiehi \mem.mem_internal.code_mem[150][3]$_SDFFCE_PN0P__1803  (.L_HI(net1803));
 sg13g2_tiehi \mem.mem_internal.code_mem[150][4]$_SDFFCE_PN0P__1804  (.L_HI(net1804));
 sg13g2_tiehi \mem.mem_internal.code_mem[150][5]$_SDFFCE_PN0P__1805  (.L_HI(net1805));
 sg13g2_tiehi \mem.mem_internal.code_mem[150][6]$_SDFFCE_PN0P__1806  (.L_HI(net1806));
 sg13g2_tiehi \mem.mem_internal.code_mem[150][7]$_SDFFCE_PN0P__1807  (.L_HI(net1807));
 sg13g2_tiehi \mem.mem_internal.code_mem[151][0]$_SDFFCE_PN0P__1808  (.L_HI(net1808));
 sg13g2_tiehi \mem.mem_internal.code_mem[151][1]$_SDFFCE_PN0P__1809  (.L_HI(net1809));
 sg13g2_tiehi \mem.mem_internal.code_mem[151][2]$_SDFFCE_PN0P__1810  (.L_HI(net1810));
 sg13g2_tiehi \mem.mem_internal.code_mem[151][3]$_SDFFCE_PN0P__1811  (.L_HI(net1811));
 sg13g2_tiehi \mem.mem_internal.code_mem[151][4]$_SDFFCE_PN0P__1812  (.L_HI(net1812));
 sg13g2_tiehi \mem.mem_internal.code_mem[151][5]$_SDFFCE_PN0P__1813  (.L_HI(net1813));
 sg13g2_tiehi \mem.mem_internal.code_mem[151][6]$_SDFFCE_PN0P__1814  (.L_HI(net1814));
 sg13g2_tiehi \mem.mem_internal.code_mem[151][7]$_SDFFCE_PN0P__1815  (.L_HI(net1815));
 sg13g2_tiehi \mem.mem_internal.code_mem[152][0]$_SDFFCE_PN0P__1816  (.L_HI(net1816));
 sg13g2_tiehi \mem.mem_internal.code_mem[152][1]$_SDFFCE_PN0P__1817  (.L_HI(net1817));
 sg13g2_tiehi \mem.mem_internal.code_mem[152][2]$_SDFFCE_PN0P__1818  (.L_HI(net1818));
 sg13g2_tiehi \mem.mem_internal.code_mem[152][3]$_SDFFCE_PN0P__1819  (.L_HI(net1819));
 sg13g2_tiehi \mem.mem_internal.code_mem[152][4]$_SDFFCE_PN0P__1820  (.L_HI(net1820));
 sg13g2_tiehi \mem.mem_internal.code_mem[152][5]$_SDFFCE_PN0P__1821  (.L_HI(net1821));
 sg13g2_tiehi \mem.mem_internal.code_mem[152][6]$_SDFFCE_PN0P__1822  (.L_HI(net1822));
 sg13g2_tiehi \mem.mem_internal.code_mem[152][7]$_SDFFCE_PN0P__1823  (.L_HI(net1823));
 sg13g2_tiehi \mem.mem_internal.code_mem[153][0]$_SDFFCE_PN0P__1824  (.L_HI(net1824));
 sg13g2_tiehi \mem.mem_internal.code_mem[153][1]$_SDFFCE_PN0P__1825  (.L_HI(net1825));
 sg13g2_tiehi \mem.mem_internal.code_mem[153][2]$_SDFFCE_PN0P__1826  (.L_HI(net1826));
 sg13g2_tiehi \mem.mem_internal.code_mem[153][3]$_SDFFCE_PN0P__1827  (.L_HI(net1827));
 sg13g2_tiehi \mem.mem_internal.code_mem[153][4]$_SDFFCE_PN0P__1828  (.L_HI(net1828));
 sg13g2_tiehi \mem.mem_internal.code_mem[153][5]$_SDFFCE_PN0P__1829  (.L_HI(net1829));
 sg13g2_tiehi \mem.mem_internal.code_mem[153][6]$_SDFFCE_PN0P__1830  (.L_HI(net1830));
 sg13g2_tiehi \mem.mem_internal.code_mem[153][7]$_SDFFCE_PN0P__1831  (.L_HI(net1831));
 sg13g2_tiehi \mem.mem_internal.code_mem[154][0]$_SDFFCE_PN0P__1832  (.L_HI(net1832));
 sg13g2_tiehi \mem.mem_internal.code_mem[154][1]$_SDFFCE_PN0P__1833  (.L_HI(net1833));
 sg13g2_tiehi \mem.mem_internal.code_mem[154][2]$_SDFFCE_PN0P__1834  (.L_HI(net1834));
 sg13g2_tiehi \mem.mem_internal.code_mem[154][3]$_SDFFCE_PN0P__1835  (.L_HI(net1835));
 sg13g2_tiehi \mem.mem_internal.code_mem[154][4]$_SDFFCE_PN0P__1836  (.L_HI(net1836));
 sg13g2_tiehi \mem.mem_internal.code_mem[154][5]$_SDFFCE_PN0P__1837  (.L_HI(net1837));
 sg13g2_tiehi \mem.mem_internal.code_mem[154][6]$_SDFFCE_PN0P__1838  (.L_HI(net1838));
 sg13g2_tiehi \mem.mem_internal.code_mem[154][7]$_SDFFCE_PN0P__1839  (.L_HI(net1839));
 sg13g2_tiehi \mem.mem_internal.code_mem[155][0]$_SDFFCE_PN0P__1840  (.L_HI(net1840));
 sg13g2_tiehi \mem.mem_internal.code_mem[155][1]$_SDFFCE_PN0P__1841  (.L_HI(net1841));
 sg13g2_tiehi \mem.mem_internal.code_mem[155][2]$_SDFFCE_PN0P__1842  (.L_HI(net1842));
 sg13g2_tiehi \mem.mem_internal.code_mem[155][3]$_SDFFCE_PN0P__1843  (.L_HI(net1843));
 sg13g2_tiehi \mem.mem_internal.code_mem[155][4]$_SDFFCE_PN0P__1844  (.L_HI(net1844));
 sg13g2_tiehi \mem.mem_internal.code_mem[155][5]$_SDFFCE_PN0P__1845  (.L_HI(net1845));
 sg13g2_tiehi \mem.mem_internal.code_mem[155][6]$_SDFFCE_PN0P__1846  (.L_HI(net1846));
 sg13g2_tiehi \mem.mem_internal.code_mem[155][7]$_SDFFCE_PN0P__1847  (.L_HI(net1847));
 sg13g2_tiehi \mem.mem_internal.code_mem[156][0]$_SDFFCE_PN0P__1848  (.L_HI(net1848));
 sg13g2_tiehi \mem.mem_internal.code_mem[156][1]$_SDFFCE_PN0P__1849  (.L_HI(net1849));
 sg13g2_tiehi \mem.mem_internal.code_mem[156][2]$_SDFFCE_PN0P__1850  (.L_HI(net1850));
 sg13g2_tiehi \mem.mem_internal.code_mem[156][3]$_SDFFCE_PN0P__1851  (.L_HI(net1851));
 sg13g2_tiehi \mem.mem_internal.code_mem[156][4]$_SDFFCE_PN0P__1852  (.L_HI(net1852));
 sg13g2_tiehi \mem.mem_internal.code_mem[156][5]$_SDFFCE_PN0P__1853  (.L_HI(net1853));
 sg13g2_tiehi \mem.mem_internal.code_mem[156][6]$_SDFFCE_PN0P__1854  (.L_HI(net1854));
 sg13g2_tiehi \mem.mem_internal.code_mem[156][7]$_SDFFCE_PN0P__1855  (.L_HI(net1855));
 sg13g2_tiehi \mem.mem_internal.code_mem[157][0]$_SDFFCE_PN0P__1856  (.L_HI(net1856));
 sg13g2_tiehi \mem.mem_internal.code_mem[157][1]$_SDFFCE_PN0P__1857  (.L_HI(net1857));
 sg13g2_tiehi \mem.mem_internal.code_mem[157][2]$_SDFFCE_PN0P__1858  (.L_HI(net1858));
 sg13g2_tiehi \mem.mem_internal.code_mem[157][3]$_SDFFCE_PN0P__1859  (.L_HI(net1859));
 sg13g2_tiehi \mem.mem_internal.code_mem[157][4]$_SDFFCE_PN0P__1860  (.L_HI(net1860));
 sg13g2_tiehi \mem.mem_internal.code_mem[157][5]$_SDFFCE_PN0P__1861  (.L_HI(net1861));
 sg13g2_tiehi \mem.mem_internal.code_mem[157][6]$_SDFFCE_PN0P__1862  (.L_HI(net1862));
 sg13g2_tiehi \mem.mem_internal.code_mem[157][7]$_SDFFCE_PN0P__1863  (.L_HI(net1863));
 sg13g2_tiehi \mem.mem_internal.code_mem[158][0]$_SDFFCE_PN0P__1864  (.L_HI(net1864));
 sg13g2_tiehi \mem.mem_internal.code_mem[158][1]$_SDFFCE_PN0P__1865  (.L_HI(net1865));
 sg13g2_tiehi \mem.mem_internal.code_mem[158][2]$_SDFFCE_PN0P__1866  (.L_HI(net1866));
 sg13g2_tiehi \mem.mem_internal.code_mem[158][3]$_SDFFCE_PN0P__1867  (.L_HI(net1867));
 sg13g2_tiehi \mem.mem_internal.code_mem[158][4]$_SDFFCE_PN0P__1868  (.L_HI(net1868));
 sg13g2_tiehi \mem.mem_internal.code_mem[158][5]$_SDFFCE_PN0P__1869  (.L_HI(net1869));
 sg13g2_tiehi \mem.mem_internal.code_mem[158][6]$_SDFFCE_PN0P__1870  (.L_HI(net1870));
 sg13g2_tiehi \mem.mem_internal.code_mem[158][7]$_SDFFCE_PN0P__1871  (.L_HI(net1871));
 sg13g2_tiehi \mem.mem_internal.code_mem[159][0]$_SDFFCE_PN0P__1872  (.L_HI(net1872));
 sg13g2_tiehi \mem.mem_internal.code_mem[159][1]$_SDFFCE_PN0P__1873  (.L_HI(net1873));
 sg13g2_tiehi \mem.mem_internal.code_mem[159][2]$_SDFFCE_PN0P__1874  (.L_HI(net1874));
 sg13g2_tiehi \mem.mem_internal.code_mem[159][3]$_SDFFCE_PN0P__1875  (.L_HI(net1875));
 sg13g2_tiehi \mem.mem_internal.code_mem[159][4]$_SDFFCE_PN0P__1876  (.L_HI(net1876));
 sg13g2_tiehi \mem.mem_internal.code_mem[159][5]$_SDFFCE_PN0P__1877  (.L_HI(net1877));
 sg13g2_tiehi \mem.mem_internal.code_mem[159][6]$_SDFFCE_PN0P__1878  (.L_HI(net1878));
 sg13g2_tiehi \mem.mem_internal.code_mem[159][7]$_SDFFCE_PN0P__1879  (.L_HI(net1879));
 sg13g2_tiehi \mem.mem_internal.code_mem[15][0]$_SDFFCE_PN0P__1880  (.L_HI(net1880));
 sg13g2_tiehi \mem.mem_internal.code_mem[15][1]$_SDFFCE_PN0P__1881  (.L_HI(net1881));
 sg13g2_tiehi \mem.mem_internal.code_mem[15][2]$_SDFFCE_PN0P__1882  (.L_HI(net1882));
 sg13g2_tiehi \mem.mem_internal.code_mem[15][3]$_SDFFCE_PN0P__1883  (.L_HI(net1883));
 sg13g2_tiehi \mem.mem_internal.code_mem[15][4]$_SDFFCE_PN0P__1884  (.L_HI(net1884));
 sg13g2_tiehi \mem.mem_internal.code_mem[15][5]$_SDFFCE_PN0P__1885  (.L_HI(net1885));
 sg13g2_tiehi \mem.mem_internal.code_mem[15][6]$_SDFFCE_PN0P__1886  (.L_HI(net1886));
 sg13g2_tiehi \mem.mem_internal.code_mem[15][7]$_SDFFCE_PN0P__1887  (.L_HI(net1887));
 sg13g2_tiehi \mem.mem_internal.code_mem[160][0]$_SDFFCE_PN0P__1888  (.L_HI(net1888));
 sg13g2_tiehi \mem.mem_internal.code_mem[160][1]$_SDFFCE_PN0P__1889  (.L_HI(net1889));
 sg13g2_tiehi \mem.mem_internal.code_mem[160][2]$_SDFFCE_PN0P__1890  (.L_HI(net1890));
 sg13g2_tiehi \mem.mem_internal.code_mem[160][3]$_SDFFCE_PN0P__1891  (.L_HI(net1891));
 sg13g2_tiehi \mem.mem_internal.code_mem[160][4]$_SDFFCE_PN0P__1892  (.L_HI(net1892));
 sg13g2_tiehi \mem.mem_internal.code_mem[160][5]$_SDFFCE_PN0P__1893  (.L_HI(net1893));
 sg13g2_tiehi \mem.mem_internal.code_mem[160][6]$_SDFFCE_PN0P__1894  (.L_HI(net1894));
 sg13g2_tiehi \mem.mem_internal.code_mem[160][7]$_SDFFCE_PN0P__1895  (.L_HI(net1895));
 sg13g2_tiehi \mem.mem_internal.code_mem[161][0]$_SDFFCE_PN0P__1896  (.L_HI(net1896));
 sg13g2_tiehi \mem.mem_internal.code_mem[161][1]$_SDFFCE_PN0P__1897  (.L_HI(net1897));
 sg13g2_tiehi \mem.mem_internal.code_mem[161][2]$_SDFFCE_PN0P__1898  (.L_HI(net1898));
 sg13g2_tiehi \mem.mem_internal.code_mem[161][3]$_SDFFCE_PN0P__1899  (.L_HI(net1899));
 sg13g2_tiehi \mem.mem_internal.code_mem[161][4]$_SDFFCE_PN0P__1900  (.L_HI(net1900));
 sg13g2_tiehi \mem.mem_internal.code_mem[161][5]$_SDFFCE_PN0P__1901  (.L_HI(net1901));
 sg13g2_tiehi \mem.mem_internal.code_mem[161][6]$_SDFFCE_PN0P__1902  (.L_HI(net1902));
 sg13g2_tiehi \mem.mem_internal.code_mem[161][7]$_SDFFCE_PN0P__1903  (.L_HI(net1903));
 sg13g2_tiehi \mem.mem_internal.code_mem[162][0]$_SDFFCE_PN0P__1904  (.L_HI(net1904));
 sg13g2_tiehi \mem.mem_internal.code_mem[162][1]$_SDFFCE_PN0P__1905  (.L_HI(net1905));
 sg13g2_tiehi \mem.mem_internal.code_mem[162][2]$_SDFFCE_PN0P__1906  (.L_HI(net1906));
 sg13g2_tiehi \mem.mem_internal.code_mem[162][3]$_SDFFCE_PN0P__1907  (.L_HI(net1907));
 sg13g2_tiehi \mem.mem_internal.code_mem[162][4]$_SDFFCE_PN0P__1908  (.L_HI(net1908));
 sg13g2_tiehi \mem.mem_internal.code_mem[162][5]$_SDFFCE_PN0P__1909  (.L_HI(net1909));
 sg13g2_tiehi \mem.mem_internal.code_mem[162][6]$_SDFFCE_PN0P__1910  (.L_HI(net1910));
 sg13g2_tiehi \mem.mem_internal.code_mem[162][7]$_SDFFCE_PN0P__1911  (.L_HI(net1911));
 sg13g2_tiehi \mem.mem_internal.code_mem[163][0]$_SDFFCE_PN0P__1912  (.L_HI(net1912));
 sg13g2_tiehi \mem.mem_internal.code_mem[163][1]$_SDFFCE_PN0P__1913  (.L_HI(net1913));
 sg13g2_tiehi \mem.mem_internal.code_mem[163][2]$_SDFFCE_PN0P__1914  (.L_HI(net1914));
 sg13g2_tiehi \mem.mem_internal.code_mem[163][3]$_SDFFCE_PN0P__1915  (.L_HI(net1915));
 sg13g2_tiehi \mem.mem_internal.code_mem[163][4]$_SDFFCE_PN0P__1916  (.L_HI(net1916));
 sg13g2_tiehi \mem.mem_internal.code_mem[163][5]$_SDFFCE_PN0P__1917  (.L_HI(net1917));
 sg13g2_tiehi \mem.mem_internal.code_mem[163][6]$_SDFFCE_PN0P__1918  (.L_HI(net1918));
 sg13g2_tiehi \mem.mem_internal.code_mem[163][7]$_SDFFCE_PN0P__1919  (.L_HI(net1919));
 sg13g2_tiehi \mem.mem_internal.code_mem[164][0]$_SDFFCE_PN0P__1920  (.L_HI(net1920));
 sg13g2_tiehi \mem.mem_internal.code_mem[164][1]$_SDFFCE_PN0P__1921  (.L_HI(net1921));
 sg13g2_tiehi \mem.mem_internal.code_mem[164][2]$_SDFFCE_PN0P__1922  (.L_HI(net1922));
 sg13g2_tiehi \mem.mem_internal.code_mem[164][3]$_SDFFCE_PN0P__1923  (.L_HI(net1923));
 sg13g2_tiehi \mem.mem_internal.code_mem[164][4]$_SDFFCE_PN0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \mem.mem_internal.code_mem[164][5]$_SDFFCE_PN0P__1925  (.L_HI(net1925));
 sg13g2_tiehi \mem.mem_internal.code_mem[164][6]$_SDFFCE_PN0P__1926  (.L_HI(net1926));
 sg13g2_tiehi \mem.mem_internal.code_mem[164][7]$_SDFFCE_PN0P__1927  (.L_HI(net1927));
 sg13g2_tiehi \mem.mem_internal.code_mem[165][0]$_SDFFCE_PN0P__1928  (.L_HI(net1928));
 sg13g2_tiehi \mem.mem_internal.code_mem[165][1]$_SDFFCE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \mem.mem_internal.code_mem[165][2]$_SDFFCE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \mem.mem_internal.code_mem[165][3]$_SDFFCE_PN0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \mem.mem_internal.code_mem[165][4]$_SDFFCE_PN0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \mem.mem_internal.code_mem[165][5]$_SDFFCE_PN0P__1933  (.L_HI(net1933));
 sg13g2_tiehi \mem.mem_internal.code_mem[165][6]$_SDFFCE_PN0P__1934  (.L_HI(net1934));
 sg13g2_tiehi \mem.mem_internal.code_mem[165][7]$_SDFFCE_PN0P__1935  (.L_HI(net1935));
 sg13g2_tiehi \mem.mem_internal.code_mem[166][0]$_SDFFCE_PN0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \mem.mem_internal.code_mem[166][1]$_SDFFCE_PN0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \mem.mem_internal.code_mem[166][2]$_SDFFCE_PN0P__1938  (.L_HI(net1938));
 sg13g2_tiehi \mem.mem_internal.code_mem[166][3]$_SDFFCE_PN0P__1939  (.L_HI(net1939));
 sg13g2_tiehi \mem.mem_internal.code_mem[166][4]$_SDFFCE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \mem.mem_internal.code_mem[166][5]$_SDFFCE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \mem.mem_internal.code_mem[166][6]$_SDFFCE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \mem.mem_internal.code_mem[166][7]$_SDFFCE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \mem.mem_internal.code_mem[167][0]$_SDFFCE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \mem.mem_internal.code_mem[167][1]$_SDFFCE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \mem.mem_internal.code_mem[167][2]$_SDFFCE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \mem.mem_internal.code_mem[167][3]$_SDFFCE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \mem.mem_internal.code_mem[167][4]$_SDFFCE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \mem.mem_internal.code_mem[167][5]$_SDFFCE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \mem.mem_internal.code_mem[167][6]$_SDFFCE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \mem.mem_internal.code_mem[167][7]$_SDFFCE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \mem.mem_internal.code_mem[168][0]$_SDFFCE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \mem.mem_internal.code_mem[168][1]$_SDFFCE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \mem.mem_internal.code_mem[168][2]$_SDFFCE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \mem.mem_internal.code_mem[168][3]$_SDFFCE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \mem.mem_internal.code_mem[168][4]$_SDFFCE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \mem.mem_internal.code_mem[168][5]$_SDFFCE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \mem.mem_internal.code_mem[168][6]$_SDFFCE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \mem.mem_internal.code_mem[168][7]$_SDFFCE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \mem.mem_internal.code_mem[169][0]$_SDFFCE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \mem.mem_internal.code_mem[169][1]$_SDFFCE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \mem.mem_internal.code_mem[169][2]$_SDFFCE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \mem.mem_internal.code_mem[169][3]$_SDFFCE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \mem.mem_internal.code_mem[169][4]$_SDFFCE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \mem.mem_internal.code_mem[169][5]$_SDFFCE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \mem.mem_internal.code_mem[169][6]$_SDFFCE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \mem.mem_internal.code_mem[169][7]$_SDFFCE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \mem.mem_internal.code_mem[16][0]$_SDFFCE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \mem.mem_internal.code_mem[16][1]$_SDFFCE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \mem.mem_internal.code_mem[16][2]$_SDFFCE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \mem.mem_internal.code_mem[16][3]$_SDFFCE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \mem.mem_internal.code_mem[16][4]$_SDFFCE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \mem.mem_internal.code_mem[16][5]$_SDFFCE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \mem.mem_internal.code_mem[16][6]$_SDFFCE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \mem.mem_internal.code_mem[16][7]$_SDFFCE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \mem.mem_internal.code_mem[170][0]$_SDFFCE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \mem.mem_internal.code_mem[170][1]$_SDFFCE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \mem.mem_internal.code_mem[170][2]$_SDFFCE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \mem.mem_internal.code_mem[170][3]$_SDFFCE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \mem.mem_internal.code_mem[170][4]$_SDFFCE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \mem.mem_internal.code_mem[170][5]$_SDFFCE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \mem.mem_internal.code_mem[170][6]$_SDFFCE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \mem.mem_internal.code_mem[170][7]$_SDFFCE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \mem.mem_internal.code_mem[171][0]$_SDFFCE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \mem.mem_internal.code_mem[171][1]$_SDFFCE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \mem.mem_internal.code_mem[171][2]$_SDFFCE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \mem.mem_internal.code_mem[171][3]$_SDFFCE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \mem.mem_internal.code_mem[171][4]$_SDFFCE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \mem.mem_internal.code_mem[171][5]$_SDFFCE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \mem.mem_internal.code_mem[171][6]$_SDFFCE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \mem.mem_internal.code_mem[171][7]$_SDFFCE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \mem.mem_internal.code_mem[172][0]$_SDFFCE_PN0P__1992  (.L_HI(net1992));
 sg13g2_tiehi \mem.mem_internal.code_mem[172][1]$_SDFFCE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \mem.mem_internal.code_mem[172][2]$_SDFFCE_PN0P__1994  (.L_HI(net1994));
 sg13g2_tiehi \mem.mem_internal.code_mem[172][3]$_SDFFCE_PN0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \mem.mem_internal.code_mem[172][4]$_SDFFCE_PN0P__1996  (.L_HI(net1996));
 sg13g2_tiehi \mem.mem_internal.code_mem[172][5]$_SDFFCE_PN0P__1997  (.L_HI(net1997));
 sg13g2_tiehi \mem.mem_internal.code_mem[172][6]$_SDFFCE_PN0P__1998  (.L_HI(net1998));
 sg13g2_tiehi \mem.mem_internal.code_mem[172][7]$_SDFFCE_PN0P__1999  (.L_HI(net1999));
 sg13g2_tiehi \mem.mem_internal.code_mem[173][0]$_SDFFCE_PN0P__2000  (.L_HI(net2000));
 sg13g2_tiehi \mem.mem_internal.code_mem[173][1]$_SDFFCE_PN0P__2001  (.L_HI(net2001));
 sg13g2_tiehi \mem.mem_internal.code_mem[173][2]$_SDFFCE_PN0P__2002  (.L_HI(net2002));
 sg13g2_tiehi \mem.mem_internal.code_mem[173][3]$_SDFFCE_PN0P__2003  (.L_HI(net2003));
 sg13g2_tiehi \mem.mem_internal.code_mem[173][4]$_SDFFCE_PN0P__2004  (.L_HI(net2004));
 sg13g2_tiehi \mem.mem_internal.code_mem[173][5]$_SDFFCE_PN0P__2005  (.L_HI(net2005));
 sg13g2_tiehi \mem.mem_internal.code_mem[173][6]$_SDFFCE_PN0P__2006  (.L_HI(net2006));
 sg13g2_tiehi \mem.mem_internal.code_mem[173][7]$_SDFFCE_PN0P__2007  (.L_HI(net2007));
 sg13g2_tiehi \mem.mem_internal.code_mem[174][0]$_SDFFCE_PN0P__2008  (.L_HI(net2008));
 sg13g2_tiehi \mem.mem_internal.code_mem[174][1]$_SDFFCE_PN0P__2009  (.L_HI(net2009));
 sg13g2_tiehi \mem.mem_internal.code_mem[174][2]$_SDFFCE_PN0P__2010  (.L_HI(net2010));
 sg13g2_tiehi \mem.mem_internal.code_mem[174][3]$_SDFFCE_PN0P__2011  (.L_HI(net2011));
 sg13g2_tiehi \mem.mem_internal.code_mem[174][4]$_SDFFCE_PN0P__2012  (.L_HI(net2012));
 sg13g2_tiehi \mem.mem_internal.code_mem[174][5]$_SDFFCE_PN0P__2013  (.L_HI(net2013));
 sg13g2_tiehi \mem.mem_internal.code_mem[174][6]$_SDFFCE_PN0P__2014  (.L_HI(net2014));
 sg13g2_tiehi \mem.mem_internal.code_mem[174][7]$_SDFFCE_PN0P__2015  (.L_HI(net2015));
 sg13g2_tiehi \mem.mem_internal.code_mem[175][0]$_SDFFCE_PN0P__2016  (.L_HI(net2016));
 sg13g2_tiehi \mem.mem_internal.code_mem[175][1]$_SDFFCE_PN0P__2017  (.L_HI(net2017));
 sg13g2_tiehi \mem.mem_internal.code_mem[175][2]$_SDFFCE_PN0P__2018  (.L_HI(net2018));
 sg13g2_tiehi \mem.mem_internal.code_mem[175][3]$_SDFFCE_PN0P__2019  (.L_HI(net2019));
 sg13g2_tiehi \mem.mem_internal.code_mem[175][4]$_SDFFCE_PN0P__2020  (.L_HI(net2020));
 sg13g2_tiehi \mem.mem_internal.code_mem[175][5]$_SDFFCE_PN0P__2021  (.L_HI(net2021));
 sg13g2_tiehi \mem.mem_internal.code_mem[175][6]$_SDFFCE_PN0P__2022  (.L_HI(net2022));
 sg13g2_tiehi \mem.mem_internal.code_mem[175][7]$_SDFFCE_PN0P__2023  (.L_HI(net2023));
 sg13g2_tiehi \mem.mem_internal.code_mem[176][0]$_SDFFCE_PN0P__2024  (.L_HI(net2024));
 sg13g2_tiehi \mem.mem_internal.code_mem[176][1]$_SDFFCE_PN0P__2025  (.L_HI(net2025));
 sg13g2_tiehi \mem.mem_internal.code_mem[176][2]$_SDFFCE_PN0P__2026  (.L_HI(net2026));
 sg13g2_tiehi \mem.mem_internal.code_mem[176][3]$_SDFFCE_PN0P__2027  (.L_HI(net2027));
 sg13g2_tiehi \mem.mem_internal.code_mem[176][4]$_SDFFCE_PN0P__2028  (.L_HI(net2028));
 sg13g2_tiehi \mem.mem_internal.code_mem[176][5]$_SDFFCE_PN0P__2029  (.L_HI(net2029));
 sg13g2_tiehi \mem.mem_internal.code_mem[176][6]$_SDFFCE_PN0P__2030  (.L_HI(net2030));
 sg13g2_tiehi \mem.mem_internal.code_mem[176][7]$_SDFFCE_PN0P__2031  (.L_HI(net2031));
 sg13g2_tiehi \mem.mem_internal.code_mem[177][0]$_SDFFCE_PN0P__2032  (.L_HI(net2032));
 sg13g2_tiehi \mem.mem_internal.code_mem[177][1]$_SDFFCE_PN0P__2033  (.L_HI(net2033));
 sg13g2_tiehi \mem.mem_internal.code_mem[177][2]$_SDFFCE_PN0P__2034  (.L_HI(net2034));
 sg13g2_tiehi \mem.mem_internal.code_mem[177][3]$_SDFFCE_PN0P__2035  (.L_HI(net2035));
 sg13g2_tiehi \mem.mem_internal.code_mem[177][4]$_SDFFCE_PN0P__2036  (.L_HI(net2036));
 sg13g2_tiehi \mem.mem_internal.code_mem[177][5]$_SDFFCE_PN0P__2037  (.L_HI(net2037));
 sg13g2_tiehi \mem.mem_internal.code_mem[177][6]$_SDFFCE_PN0P__2038  (.L_HI(net2038));
 sg13g2_tiehi \mem.mem_internal.code_mem[177][7]$_SDFFCE_PN0P__2039  (.L_HI(net2039));
 sg13g2_tiehi \mem.mem_internal.code_mem[178][0]$_SDFFCE_PN0P__2040  (.L_HI(net2040));
 sg13g2_tiehi \mem.mem_internal.code_mem[178][1]$_SDFFCE_PN0P__2041  (.L_HI(net2041));
 sg13g2_tiehi \mem.mem_internal.code_mem[178][2]$_SDFFCE_PN0P__2042  (.L_HI(net2042));
 sg13g2_tiehi \mem.mem_internal.code_mem[178][3]$_SDFFCE_PN0P__2043  (.L_HI(net2043));
 sg13g2_tiehi \mem.mem_internal.code_mem[178][4]$_SDFFCE_PN0P__2044  (.L_HI(net2044));
 sg13g2_tiehi \mem.mem_internal.code_mem[178][5]$_SDFFCE_PN0P__2045  (.L_HI(net2045));
 sg13g2_tiehi \mem.mem_internal.code_mem[178][6]$_SDFFCE_PN0P__2046  (.L_HI(net2046));
 sg13g2_tiehi \mem.mem_internal.code_mem[178][7]$_SDFFCE_PN0P__2047  (.L_HI(net2047));
 sg13g2_tiehi \mem.mem_internal.code_mem[179][0]$_SDFFCE_PN0P__2048  (.L_HI(net2048));
 sg13g2_tiehi \mem.mem_internal.code_mem[179][1]$_SDFFCE_PN0P__2049  (.L_HI(net2049));
 sg13g2_tiehi \mem.mem_internal.code_mem[179][2]$_SDFFCE_PN0P__2050  (.L_HI(net2050));
 sg13g2_tiehi \mem.mem_internal.code_mem[179][3]$_SDFFCE_PN0P__2051  (.L_HI(net2051));
 sg13g2_tiehi \mem.mem_internal.code_mem[179][4]$_SDFFCE_PN0P__2052  (.L_HI(net2052));
 sg13g2_tiehi \mem.mem_internal.code_mem[179][5]$_SDFFCE_PN0P__2053  (.L_HI(net2053));
 sg13g2_tiehi \mem.mem_internal.code_mem[179][6]$_SDFFCE_PN0P__2054  (.L_HI(net2054));
 sg13g2_tiehi \mem.mem_internal.code_mem[179][7]$_SDFFCE_PN0P__2055  (.L_HI(net2055));
 sg13g2_tiehi \mem.mem_internal.code_mem[17][0]$_SDFFCE_PN0P__2056  (.L_HI(net2056));
 sg13g2_tiehi \mem.mem_internal.code_mem[17][1]$_SDFFCE_PN0P__2057  (.L_HI(net2057));
 sg13g2_tiehi \mem.mem_internal.code_mem[17][2]$_SDFFCE_PN0P__2058  (.L_HI(net2058));
 sg13g2_tiehi \mem.mem_internal.code_mem[17][3]$_SDFFCE_PN0P__2059  (.L_HI(net2059));
 sg13g2_tiehi \mem.mem_internal.code_mem[17][4]$_SDFFCE_PN0P__2060  (.L_HI(net2060));
 sg13g2_tiehi \mem.mem_internal.code_mem[17][5]$_SDFFCE_PN0P__2061  (.L_HI(net2061));
 sg13g2_tiehi \mem.mem_internal.code_mem[17][6]$_SDFFCE_PN0P__2062  (.L_HI(net2062));
 sg13g2_tiehi \mem.mem_internal.code_mem[17][7]$_SDFFCE_PN0P__2063  (.L_HI(net2063));
 sg13g2_tiehi \mem.mem_internal.code_mem[180][0]$_SDFFCE_PN0P__2064  (.L_HI(net2064));
 sg13g2_tiehi \mem.mem_internal.code_mem[180][1]$_SDFFCE_PN0P__2065  (.L_HI(net2065));
 sg13g2_tiehi \mem.mem_internal.code_mem[180][2]$_SDFFCE_PN0P__2066  (.L_HI(net2066));
 sg13g2_tiehi \mem.mem_internal.code_mem[180][3]$_SDFFCE_PN0P__2067  (.L_HI(net2067));
 sg13g2_tiehi \mem.mem_internal.code_mem[180][4]$_SDFFCE_PN0P__2068  (.L_HI(net2068));
 sg13g2_tiehi \mem.mem_internal.code_mem[180][5]$_SDFFCE_PN0P__2069  (.L_HI(net2069));
 sg13g2_tiehi \mem.mem_internal.code_mem[180][6]$_SDFFCE_PN0P__2070  (.L_HI(net2070));
 sg13g2_tiehi \mem.mem_internal.code_mem[180][7]$_SDFFCE_PN0P__2071  (.L_HI(net2071));
 sg13g2_tiehi \mem.mem_internal.code_mem[181][0]$_SDFFCE_PN0P__2072  (.L_HI(net2072));
 sg13g2_tiehi \mem.mem_internal.code_mem[181][1]$_SDFFCE_PN0P__2073  (.L_HI(net2073));
 sg13g2_tiehi \mem.mem_internal.code_mem[181][2]$_SDFFCE_PN0P__2074  (.L_HI(net2074));
 sg13g2_tiehi \mem.mem_internal.code_mem[181][3]$_SDFFCE_PN0P__2075  (.L_HI(net2075));
 sg13g2_tiehi \mem.mem_internal.code_mem[181][4]$_SDFFCE_PN0P__2076  (.L_HI(net2076));
 sg13g2_tiehi \mem.mem_internal.code_mem[181][5]$_SDFFCE_PN0P__2077  (.L_HI(net2077));
 sg13g2_tiehi \mem.mem_internal.code_mem[181][6]$_SDFFCE_PN0P__2078  (.L_HI(net2078));
 sg13g2_tiehi \mem.mem_internal.code_mem[181][7]$_SDFFCE_PN0P__2079  (.L_HI(net2079));
 sg13g2_tiehi \mem.mem_internal.code_mem[182][0]$_SDFFCE_PN0P__2080  (.L_HI(net2080));
 sg13g2_tiehi \mem.mem_internal.code_mem[182][1]$_SDFFCE_PN0P__2081  (.L_HI(net2081));
 sg13g2_tiehi \mem.mem_internal.code_mem[182][2]$_SDFFCE_PN0P__2082  (.L_HI(net2082));
 sg13g2_tiehi \mem.mem_internal.code_mem[182][3]$_SDFFCE_PN0P__2083  (.L_HI(net2083));
 sg13g2_tiehi \mem.mem_internal.code_mem[182][4]$_SDFFCE_PN0P__2084  (.L_HI(net2084));
 sg13g2_tiehi \mem.mem_internal.code_mem[182][5]$_SDFFCE_PN0P__2085  (.L_HI(net2085));
 sg13g2_tiehi \mem.mem_internal.code_mem[182][6]$_SDFFCE_PN0P__2086  (.L_HI(net2086));
 sg13g2_tiehi \mem.mem_internal.code_mem[182][7]$_SDFFCE_PN0P__2087  (.L_HI(net2087));
 sg13g2_tiehi \mem.mem_internal.code_mem[183][0]$_SDFFCE_PN0P__2088  (.L_HI(net2088));
 sg13g2_tiehi \mem.mem_internal.code_mem[183][1]$_SDFFCE_PN0P__2089  (.L_HI(net2089));
 sg13g2_tiehi \mem.mem_internal.code_mem[183][2]$_SDFFCE_PN0P__2090  (.L_HI(net2090));
 sg13g2_tiehi \mem.mem_internal.code_mem[183][3]$_SDFFCE_PN0P__2091  (.L_HI(net2091));
 sg13g2_tiehi \mem.mem_internal.code_mem[183][4]$_SDFFCE_PN0P__2092  (.L_HI(net2092));
 sg13g2_tiehi \mem.mem_internal.code_mem[183][5]$_SDFFCE_PN0P__2093  (.L_HI(net2093));
 sg13g2_tiehi \mem.mem_internal.code_mem[183][6]$_SDFFCE_PN0P__2094  (.L_HI(net2094));
 sg13g2_tiehi \mem.mem_internal.code_mem[183][7]$_SDFFCE_PN0P__2095  (.L_HI(net2095));
 sg13g2_tiehi \mem.mem_internal.code_mem[184][0]$_SDFFCE_PN0P__2096  (.L_HI(net2096));
 sg13g2_tiehi \mem.mem_internal.code_mem[184][1]$_SDFFCE_PN0P__2097  (.L_HI(net2097));
 sg13g2_tiehi \mem.mem_internal.code_mem[184][2]$_SDFFCE_PN0P__2098  (.L_HI(net2098));
 sg13g2_tiehi \mem.mem_internal.code_mem[184][3]$_SDFFCE_PN0P__2099  (.L_HI(net2099));
 sg13g2_tiehi \mem.mem_internal.code_mem[184][4]$_SDFFCE_PN0P__2100  (.L_HI(net2100));
 sg13g2_tiehi \mem.mem_internal.code_mem[184][5]$_SDFFCE_PN0P__2101  (.L_HI(net2101));
 sg13g2_tiehi \mem.mem_internal.code_mem[184][6]$_SDFFCE_PN0P__2102  (.L_HI(net2102));
 sg13g2_tiehi \mem.mem_internal.code_mem[184][7]$_SDFFCE_PN0P__2103  (.L_HI(net2103));
 sg13g2_tiehi \mem.mem_internal.code_mem[185][0]$_SDFFCE_PN0P__2104  (.L_HI(net2104));
 sg13g2_tiehi \mem.mem_internal.code_mem[185][1]$_SDFFCE_PN0P__2105  (.L_HI(net2105));
 sg13g2_tiehi \mem.mem_internal.code_mem[185][2]$_SDFFCE_PN0P__2106  (.L_HI(net2106));
 sg13g2_tiehi \mem.mem_internal.code_mem[185][3]$_SDFFCE_PN0P__2107  (.L_HI(net2107));
 sg13g2_tiehi \mem.mem_internal.code_mem[185][4]$_SDFFCE_PN0P__2108  (.L_HI(net2108));
 sg13g2_tiehi \mem.mem_internal.code_mem[185][5]$_SDFFCE_PN0P__2109  (.L_HI(net2109));
 sg13g2_tiehi \mem.mem_internal.code_mem[185][6]$_SDFFCE_PN0P__2110  (.L_HI(net2110));
 sg13g2_tiehi \mem.mem_internal.code_mem[185][7]$_SDFFCE_PN0P__2111  (.L_HI(net2111));
 sg13g2_tiehi \mem.mem_internal.code_mem[186][0]$_SDFFCE_PN0P__2112  (.L_HI(net2112));
 sg13g2_tiehi \mem.mem_internal.code_mem[186][1]$_SDFFCE_PN0P__2113  (.L_HI(net2113));
 sg13g2_tiehi \mem.mem_internal.code_mem[186][2]$_SDFFCE_PN0P__2114  (.L_HI(net2114));
 sg13g2_tiehi \mem.mem_internal.code_mem[186][3]$_SDFFCE_PN0P__2115  (.L_HI(net2115));
 sg13g2_tiehi \mem.mem_internal.code_mem[186][4]$_SDFFCE_PN0P__2116  (.L_HI(net2116));
 sg13g2_tiehi \mem.mem_internal.code_mem[186][5]$_SDFFCE_PN0P__2117  (.L_HI(net2117));
 sg13g2_tiehi \mem.mem_internal.code_mem[186][6]$_SDFFCE_PN0P__2118  (.L_HI(net2118));
 sg13g2_tiehi \mem.mem_internal.code_mem[186][7]$_SDFFCE_PN0P__2119  (.L_HI(net2119));
 sg13g2_tiehi \mem.mem_internal.code_mem[187][0]$_SDFFCE_PN0P__2120  (.L_HI(net2120));
 sg13g2_tiehi \mem.mem_internal.code_mem[187][1]$_SDFFCE_PN0P__2121  (.L_HI(net2121));
 sg13g2_tiehi \mem.mem_internal.code_mem[187][2]$_SDFFCE_PN0P__2122  (.L_HI(net2122));
 sg13g2_tiehi \mem.mem_internal.code_mem[187][3]$_SDFFCE_PN0P__2123  (.L_HI(net2123));
 sg13g2_tiehi \mem.mem_internal.code_mem[187][4]$_SDFFCE_PN0P__2124  (.L_HI(net2124));
 sg13g2_tiehi \mem.mem_internal.code_mem[187][5]$_SDFFCE_PN0P__2125  (.L_HI(net2125));
 sg13g2_tiehi \mem.mem_internal.code_mem[187][6]$_SDFFCE_PN0P__2126  (.L_HI(net2126));
 sg13g2_tiehi \mem.mem_internal.code_mem[187][7]$_SDFFCE_PN0P__2127  (.L_HI(net2127));
 sg13g2_tiehi \mem.mem_internal.code_mem[188][0]$_SDFFCE_PN0P__2128  (.L_HI(net2128));
 sg13g2_tiehi \mem.mem_internal.code_mem[188][1]$_SDFFCE_PN0P__2129  (.L_HI(net2129));
 sg13g2_tiehi \mem.mem_internal.code_mem[188][2]$_SDFFCE_PN0P__2130  (.L_HI(net2130));
 sg13g2_tiehi \mem.mem_internal.code_mem[188][3]$_SDFFCE_PN0P__2131  (.L_HI(net2131));
 sg13g2_tiehi \mem.mem_internal.code_mem[188][4]$_SDFFCE_PN0P__2132  (.L_HI(net2132));
 sg13g2_tiehi \mem.mem_internal.code_mem[188][5]$_SDFFCE_PN0P__2133  (.L_HI(net2133));
 sg13g2_tiehi \mem.mem_internal.code_mem[188][6]$_SDFFCE_PN0P__2134  (.L_HI(net2134));
 sg13g2_tiehi \mem.mem_internal.code_mem[188][7]$_SDFFCE_PN0P__2135  (.L_HI(net2135));
 sg13g2_tiehi \mem.mem_internal.code_mem[189][0]$_SDFFCE_PN0P__2136  (.L_HI(net2136));
 sg13g2_tiehi \mem.mem_internal.code_mem[189][1]$_SDFFCE_PN0P__2137  (.L_HI(net2137));
 sg13g2_tiehi \mem.mem_internal.code_mem[189][2]$_SDFFCE_PN0P__2138  (.L_HI(net2138));
 sg13g2_tiehi \mem.mem_internal.code_mem[189][3]$_SDFFCE_PN0P__2139  (.L_HI(net2139));
 sg13g2_tiehi \mem.mem_internal.code_mem[189][4]$_SDFFCE_PN0P__2140  (.L_HI(net2140));
 sg13g2_tiehi \mem.mem_internal.code_mem[189][5]$_SDFFCE_PN0P__2141  (.L_HI(net2141));
 sg13g2_tiehi \mem.mem_internal.code_mem[189][6]$_SDFFCE_PN0P__2142  (.L_HI(net2142));
 sg13g2_tiehi \mem.mem_internal.code_mem[189][7]$_SDFFCE_PN0P__2143  (.L_HI(net2143));
 sg13g2_tiehi \mem.mem_internal.code_mem[18][0]$_SDFFCE_PN0P__2144  (.L_HI(net2144));
 sg13g2_tiehi \mem.mem_internal.code_mem[18][1]$_SDFFCE_PN0P__2145  (.L_HI(net2145));
 sg13g2_tiehi \mem.mem_internal.code_mem[18][2]$_SDFFCE_PN0P__2146  (.L_HI(net2146));
 sg13g2_tiehi \mem.mem_internal.code_mem[18][3]$_SDFFCE_PN0P__2147  (.L_HI(net2147));
 sg13g2_tiehi \mem.mem_internal.code_mem[18][4]$_SDFFCE_PN0P__2148  (.L_HI(net2148));
 sg13g2_tiehi \mem.mem_internal.code_mem[18][5]$_SDFFCE_PN0P__2149  (.L_HI(net2149));
 sg13g2_tiehi \mem.mem_internal.code_mem[18][6]$_SDFFCE_PN0P__2150  (.L_HI(net2150));
 sg13g2_tiehi \mem.mem_internal.code_mem[18][7]$_SDFFCE_PN0P__2151  (.L_HI(net2151));
 sg13g2_tiehi \mem.mem_internal.code_mem[190][0]$_SDFFCE_PN0P__2152  (.L_HI(net2152));
 sg13g2_tiehi \mem.mem_internal.code_mem[190][1]$_SDFFCE_PN0P__2153  (.L_HI(net2153));
 sg13g2_tiehi \mem.mem_internal.code_mem[190][2]$_SDFFCE_PN0P__2154  (.L_HI(net2154));
 sg13g2_tiehi \mem.mem_internal.code_mem[190][3]$_SDFFCE_PN0P__2155  (.L_HI(net2155));
 sg13g2_tiehi \mem.mem_internal.code_mem[190][4]$_SDFFCE_PN0P__2156  (.L_HI(net2156));
 sg13g2_tiehi \mem.mem_internal.code_mem[190][5]$_SDFFCE_PN0P__2157  (.L_HI(net2157));
 sg13g2_tiehi \mem.mem_internal.code_mem[190][6]$_SDFFCE_PN0P__2158  (.L_HI(net2158));
 sg13g2_tiehi \mem.mem_internal.code_mem[190][7]$_SDFFCE_PN0P__2159  (.L_HI(net2159));
 sg13g2_tiehi \mem.mem_internal.code_mem[191][0]$_SDFFCE_PN0P__2160  (.L_HI(net2160));
 sg13g2_tiehi \mem.mem_internal.code_mem[191][1]$_SDFFCE_PN0P__2161  (.L_HI(net2161));
 sg13g2_tiehi \mem.mem_internal.code_mem[191][2]$_SDFFCE_PN0P__2162  (.L_HI(net2162));
 sg13g2_tiehi \mem.mem_internal.code_mem[191][3]$_SDFFCE_PN0P__2163  (.L_HI(net2163));
 sg13g2_tiehi \mem.mem_internal.code_mem[191][4]$_SDFFCE_PN0P__2164  (.L_HI(net2164));
 sg13g2_tiehi \mem.mem_internal.code_mem[191][5]$_SDFFCE_PN0P__2165  (.L_HI(net2165));
 sg13g2_tiehi \mem.mem_internal.code_mem[191][6]$_SDFFCE_PN0P__2166  (.L_HI(net2166));
 sg13g2_tiehi \mem.mem_internal.code_mem[191][7]$_SDFFCE_PN0P__2167  (.L_HI(net2167));
 sg13g2_tiehi \mem.mem_internal.code_mem[192][0]$_SDFFCE_PN0P__2168  (.L_HI(net2168));
 sg13g2_tiehi \mem.mem_internal.code_mem[192][1]$_SDFFCE_PN0P__2169  (.L_HI(net2169));
 sg13g2_tiehi \mem.mem_internal.code_mem[192][2]$_SDFFCE_PN0P__2170  (.L_HI(net2170));
 sg13g2_tiehi \mem.mem_internal.code_mem[192][3]$_SDFFCE_PN0P__2171  (.L_HI(net2171));
 sg13g2_tiehi \mem.mem_internal.code_mem[192][4]$_SDFFCE_PN0P__2172  (.L_HI(net2172));
 sg13g2_tiehi \mem.mem_internal.code_mem[192][5]$_SDFFCE_PN0P__2173  (.L_HI(net2173));
 sg13g2_tiehi \mem.mem_internal.code_mem[192][6]$_SDFFCE_PN0P__2174  (.L_HI(net2174));
 sg13g2_tiehi \mem.mem_internal.code_mem[192][7]$_SDFFCE_PN0P__2175  (.L_HI(net2175));
 sg13g2_tiehi \mem.mem_internal.code_mem[193][0]$_SDFFCE_PN0P__2176  (.L_HI(net2176));
 sg13g2_tiehi \mem.mem_internal.code_mem[193][1]$_SDFFCE_PN0P__2177  (.L_HI(net2177));
 sg13g2_tiehi \mem.mem_internal.code_mem[193][2]$_SDFFCE_PN0P__2178  (.L_HI(net2178));
 sg13g2_tiehi \mem.mem_internal.code_mem[193][3]$_SDFFCE_PN0P__2179  (.L_HI(net2179));
 sg13g2_tiehi \mem.mem_internal.code_mem[193][4]$_SDFFCE_PN0P__2180  (.L_HI(net2180));
 sg13g2_tiehi \mem.mem_internal.code_mem[193][5]$_SDFFCE_PN0P__2181  (.L_HI(net2181));
 sg13g2_tiehi \mem.mem_internal.code_mem[193][6]$_SDFFCE_PN0P__2182  (.L_HI(net2182));
 sg13g2_tiehi \mem.mem_internal.code_mem[193][7]$_SDFFCE_PN0P__2183  (.L_HI(net2183));
 sg13g2_tiehi \mem.mem_internal.code_mem[194][0]$_SDFFCE_PN0P__2184  (.L_HI(net2184));
 sg13g2_tiehi \mem.mem_internal.code_mem[194][1]$_SDFFCE_PN0P__2185  (.L_HI(net2185));
 sg13g2_tiehi \mem.mem_internal.code_mem[194][2]$_SDFFCE_PN0P__2186  (.L_HI(net2186));
 sg13g2_tiehi \mem.mem_internal.code_mem[194][3]$_SDFFCE_PN0P__2187  (.L_HI(net2187));
 sg13g2_tiehi \mem.mem_internal.code_mem[194][4]$_SDFFCE_PN0P__2188  (.L_HI(net2188));
 sg13g2_tiehi \mem.mem_internal.code_mem[194][5]$_SDFFCE_PN0P__2189  (.L_HI(net2189));
 sg13g2_tiehi \mem.mem_internal.code_mem[194][6]$_SDFFCE_PN0P__2190  (.L_HI(net2190));
 sg13g2_tiehi \mem.mem_internal.code_mem[194][7]$_SDFFCE_PN0P__2191  (.L_HI(net2191));
 sg13g2_tiehi \mem.mem_internal.code_mem[195][0]$_SDFFCE_PN0P__2192  (.L_HI(net2192));
 sg13g2_tiehi \mem.mem_internal.code_mem[195][1]$_SDFFCE_PN0P__2193  (.L_HI(net2193));
 sg13g2_tiehi \mem.mem_internal.code_mem[195][2]$_SDFFCE_PN0P__2194  (.L_HI(net2194));
 sg13g2_tiehi \mem.mem_internal.code_mem[195][3]$_SDFFCE_PN0P__2195  (.L_HI(net2195));
 sg13g2_tiehi \mem.mem_internal.code_mem[195][4]$_SDFFCE_PN0P__2196  (.L_HI(net2196));
 sg13g2_tiehi \mem.mem_internal.code_mem[195][5]$_SDFFCE_PN0P__2197  (.L_HI(net2197));
 sg13g2_tiehi \mem.mem_internal.code_mem[195][6]$_SDFFCE_PN0P__2198  (.L_HI(net2198));
 sg13g2_tiehi \mem.mem_internal.code_mem[195][7]$_SDFFCE_PN0P__2199  (.L_HI(net2199));
 sg13g2_tiehi \mem.mem_internal.code_mem[196][0]$_SDFFCE_PN0P__2200  (.L_HI(net2200));
 sg13g2_tiehi \mem.mem_internal.code_mem[196][1]$_SDFFCE_PN0P__2201  (.L_HI(net2201));
 sg13g2_tiehi \mem.mem_internal.code_mem[196][2]$_SDFFCE_PN0P__2202  (.L_HI(net2202));
 sg13g2_tiehi \mem.mem_internal.code_mem[196][3]$_SDFFCE_PN0P__2203  (.L_HI(net2203));
 sg13g2_tiehi \mem.mem_internal.code_mem[196][4]$_SDFFCE_PN0P__2204  (.L_HI(net2204));
 sg13g2_tiehi \mem.mem_internal.code_mem[196][5]$_SDFFCE_PN0P__2205  (.L_HI(net2205));
 sg13g2_tiehi \mem.mem_internal.code_mem[196][6]$_SDFFCE_PN0P__2206  (.L_HI(net2206));
 sg13g2_tiehi \mem.mem_internal.code_mem[196][7]$_SDFFCE_PN0P__2207  (.L_HI(net2207));
 sg13g2_tiehi \mem.mem_internal.code_mem[197][0]$_SDFFCE_PN0P__2208  (.L_HI(net2208));
 sg13g2_tiehi \mem.mem_internal.code_mem[197][1]$_SDFFCE_PN0P__2209  (.L_HI(net2209));
 sg13g2_tiehi \mem.mem_internal.code_mem[197][2]$_SDFFCE_PN0P__2210  (.L_HI(net2210));
 sg13g2_tiehi \mem.mem_internal.code_mem[197][3]$_SDFFCE_PN0P__2211  (.L_HI(net2211));
 sg13g2_tiehi \mem.mem_internal.code_mem[197][4]$_SDFFCE_PN0P__2212  (.L_HI(net2212));
 sg13g2_tiehi \mem.mem_internal.code_mem[197][5]$_SDFFCE_PN0P__2213  (.L_HI(net2213));
 sg13g2_tiehi \mem.mem_internal.code_mem[197][6]$_SDFFCE_PN0P__2214  (.L_HI(net2214));
 sg13g2_tiehi \mem.mem_internal.code_mem[197][7]$_SDFFCE_PN0P__2215  (.L_HI(net2215));
 sg13g2_tiehi \mem.mem_internal.code_mem[198][0]$_SDFFCE_PN0P__2216  (.L_HI(net2216));
 sg13g2_tiehi \mem.mem_internal.code_mem[198][1]$_SDFFCE_PN0P__2217  (.L_HI(net2217));
 sg13g2_tiehi \mem.mem_internal.code_mem[198][2]$_SDFFCE_PN0P__2218  (.L_HI(net2218));
 sg13g2_tiehi \mem.mem_internal.code_mem[198][3]$_SDFFCE_PN0P__2219  (.L_HI(net2219));
 sg13g2_tiehi \mem.mem_internal.code_mem[198][4]$_SDFFCE_PN0P__2220  (.L_HI(net2220));
 sg13g2_tiehi \mem.mem_internal.code_mem[198][5]$_SDFFCE_PN0P__2221  (.L_HI(net2221));
 sg13g2_tiehi \mem.mem_internal.code_mem[198][6]$_SDFFCE_PN0P__2222  (.L_HI(net2222));
 sg13g2_tiehi \mem.mem_internal.code_mem[198][7]$_SDFFCE_PN0P__2223  (.L_HI(net2223));
 sg13g2_tiehi \mem.mem_internal.code_mem[199][0]$_SDFFCE_PN0P__2224  (.L_HI(net2224));
 sg13g2_tiehi \mem.mem_internal.code_mem[199][1]$_SDFFCE_PN0P__2225  (.L_HI(net2225));
 sg13g2_tiehi \mem.mem_internal.code_mem[199][2]$_SDFFCE_PN0P__2226  (.L_HI(net2226));
 sg13g2_tiehi \mem.mem_internal.code_mem[199][3]$_SDFFCE_PN0P__2227  (.L_HI(net2227));
 sg13g2_tiehi \mem.mem_internal.code_mem[199][4]$_SDFFCE_PN0P__2228  (.L_HI(net2228));
 sg13g2_tiehi \mem.mem_internal.code_mem[199][5]$_SDFFCE_PN0P__2229  (.L_HI(net2229));
 sg13g2_tiehi \mem.mem_internal.code_mem[199][6]$_SDFFCE_PN0P__2230  (.L_HI(net2230));
 sg13g2_tiehi \mem.mem_internal.code_mem[199][7]$_SDFFCE_PN0P__2231  (.L_HI(net2231));
 sg13g2_tiehi \mem.mem_internal.code_mem[19][0]$_SDFFCE_PN0P__2232  (.L_HI(net2232));
 sg13g2_tiehi \mem.mem_internal.code_mem[19][1]$_SDFFCE_PN0P__2233  (.L_HI(net2233));
 sg13g2_tiehi \mem.mem_internal.code_mem[19][2]$_SDFFCE_PN0P__2234  (.L_HI(net2234));
 sg13g2_tiehi \mem.mem_internal.code_mem[19][3]$_SDFFCE_PN0P__2235  (.L_HI(net2235));
 sg13g2_tiehi \mem.mem_internal.code_mem[19][4]$_SDFFCE_PN0P__2236  (.L_HI(net2236));
 sg13g2_tiehi \mem.mem_internal.code_mem[19][5]$_SDFFCE_PN0P__2237  (.L_HI(net2237));
 sg13g2_tiehi \mem.mem_internal.code_mem[19][6]$_SDFFCE_PN0P__2238  (.L_HI(net2238));
 sg13g2_tiehi \mem.mem_internal.code_mem[19][7]$_SDFFCE_PN0P__2239  (.L_HI(net2239));
 sg13g2_tiehi \mem.mem_internal.code_mem[1][0]$_SDFFCE_PN0P__2240  (.L_HI(net2240));
 sg13g2_tiehi \mem.mem_internal.code_mem[1][1]$_SDFFCE_PN0P__2241  (.L_HI(net2241));
 sg13g2_tiehi \mem.mem_internal.code_mem[1][2]$_SDFFCE_PN0P__2242  (.L_HI(net2242));
 sg13g2_tiehi \mem.mem_internal.code_mem[1][3]$_SDFFCE_PN0P__2243  (.L_HI(net2243));
 sg13g2_tiehi \mem.mem_internal.code_mem[1][4]$_SDFFCE_PN0P__2244  (.L_HI(net2244));
 sg13g2_tiehi \mem.mem_internal.code_mem[1][5]$_SDFFCE_PN0P__2245  (.L_HI(net2245));
 sg13g2_tiehi \mem.mem_internal.code_mem[1][6]$_SDFFCE_PN0P__2246  (.L_HI(net2246));
 sg13g2_tiehi \mem.mem_internal.code_mem[1][7]$_SDFFCE_PN0P__2247  (.L_HI(net2247));
 sg13g2_tiehi \mem.mem_internal.code_mem[200][0]$_SDFFCE_PN0P__2248  (.L_HI(net2248));
 sg13g2_tiehi \mem.mem_internal.code_mem[200][1]$_SDFFCE_PN0P__2249  (.L_HI(net2249));
 sg13g2_tiehi \mem.mem_internal.code_mem[200][2]$_SDFFCE_PN0P__2250  (.L_HI(net2250));
 sg13g2_tiehi \mem.mem_internal.code_mem[200][3]$_SDFFCE_PN0P__2251  (.L_HI(net2251));
 sg13g2_tiehi \mem.mem_internal.code_mem[200][4]$_SDFFCE_PN0P__2252  (.L_HI(net2252));
 sg13g2_tiehi \mem.mem_internal.code_mem[200][5]$_SDFFCE_PN0P__2253  (.L_HI(net2253));
 sg13g2_tiehi \mem.mem_internal.code_mem[200][6]$_SDFFCE_PN0P__2254  (.L_HI(net2254));
 sg13g2_tiehi \mem.mem_internal.code_mem[200][7]$_SDFFCE_PN0P__2255  (.L_HI(net2255));
 sg13g2_tiehi \mem.mem_internal.code_mem[201][0]$_SDFFCE_PN0P__2256  (.L_HI(net2256));
 sg13g2_tiehi \mem.mem_internal.code_mem[201][1]$_SDFFCE_PN0P__2257  (.L_HI(net2257));
 sg13g2_tiehi \mem.mem_internal.code_mem[201][2]$_SDFFCE_PN0P__2258  (.L_HI(net2258));
 sg13g2_tiehi \mem.mem_internal.code_mem[201][3]$_SDFFCE_PN0P__2259  (.L_HI(net2259));
 sg13g2_tiehi \mem.mem_internal.code_mem[201][4]$_SDFFCE_PN0P__2260  (.L_HI(net2260));
 sg13g2_tiehi \mem.mem_internal.code_mem[201][5]$_SDFFCE_PN0P__2261  (.L_HI(net2261));
 sg13g2_tiehi \mem.mem_internal.code_mem[201][6]$_SDFFCE_PN0P__2262  (.L_HI(net2262));
 sg13g2_tiehi \mem.mem_internal.code_mem[201][7]$_SDFFCE_PN0P__2263  (.L_HI(net2263));
 sg13g2_tiehi \mem.mem_internal.code_mem[202][0]$_SDFFCE_PN0P__2264  (.L_HI(net2264));
 sg13g2_tiehi \mem.mem_internal.code_mem[202][1]$_SDFFCE_PN0P__2265  (.L_HI(net2265));
 sg13g2_tiehi \mem.mem_internal.code_mem[202][2]$_SDFFCE_PN0P__2266  (.L_HI(net2266));
 sg13g2_tiehi \mem.mem_internal.code_mem[202][3]$_SDFFCE_PN0P__2267  (.L_HI(net2267));
 sg13g2_tiehi \mem.mem_internal.code_mem[202][4]$_SDFFCE_PN0P__2268  (.L_HI(net2268));
 sg13g2_tiehi \mem.mem_internal.code_mem[202][5]$_SDFFCE_PN0P__2269  (.L_HI(net2269));
 sg13g2_tiehi \mem.mem_internal.code_mem[202][6]$_SDFFCE_PN0P__2270  (.L_HI(net2270));
 sg13g2_tiehi \mem.mem_internal.code_mem[202][7]$_SDFFCE_PN0P__2271  (.L_HI(net2271));
 sg13g2_tiehi \mem.mem_internal.code_mem[203][0]$_SDFFCE_PN0P__2272  (.L_HI(net2272));
 sg13g2_tiehi \mem.mem_internal.code_mem[203][1]$_SDFFCE_PN0P__2273  (.L_HI(net2273));
 sg13g2_tiehi \mem.mem_internal.code_mem[203][2]$_SDFFCE_PN0P__2274  (.L_HI(net2274));
 sg13g2_tiehi \mem.mem_internal.code_mem[203][3]$_SDFFCE_PN0P__2275  (.L_HI(net2275));
 sg13g2_tiehi \mem.mem_internal.code_mem[203][4]$_SDFFCE_PN0P__2276  (.L_HI(net2276));
 sg13g2_tiehi \mem.mem_internal.code_mem[203][5]$_SDFFCE_PN0P__2277  (.L_HI(net2277));
 sg13g2_tiehi \mem.mem_internal.code_mem[203][6]$_SDFFCE_PN0P__2278  (.L_HI(net2278));
 sg13g2_tiehi \mem.mem_internal.code_mem[203][7]$_SDFFCE_PN0P__2279  (.L_HI(net2279));
 sg13g2_tiehi \mem.mem_internal.code_mem[204][0]$_SDFFCE_PN0P__2280  (.L_HI(net2280));
 sg13g2_tiehi \mem.mem_internal.code_mem[204][1]$_SDFFCE_PN0P__2281  (.L_HI(net2281));
 sg13g2_tiehi \mem.mem_internal.code_mem[204][2]$_SDFFCE_PN0P__2282  (.L_HI(net2282));
 sg13g2_tiehi \mem.mem_internal.code_mem[204][3]$_SDFFCE_PN0P__2283  (.L_HI(net2283));
 sg13g2_tiehi \mem.mem_internal.code_mem[204][4]$_SDFFCE_PN0P__2284  (.L_HI(net2284));
 sg13g2_tiehi \mem.mem_internal.code_mem[204][5]$_SDFFCE_PN0P__2285  (.L_HI(net2285));
 sg13g2_tiehi \mem.mem_internal.code_mem[204][6]$_SDFFCE_PN0P__2286  (.L_HI(net2286));
 sg13g2_tiehi \mem.mem_internal.code_mem[204][7]$_SDFFCE_PN0P__2287  (.L_HI(net2287));
 sg13g2_tiehi \mem.mem_internal.code_mem[205][0]$_SDFFCE_PN0P__2288  (.L_HI(net2288));
 sg13g2_tiehi \mem.mem_internal.code_mem[205][1]$_SDFFCE_PN0P__2289  (.L_HI(net2289));
 sg13g2_tiehi \mem.mem_internal.code_mem[205][2]$_SDFFCE_PN0P__2290  (.L_HI(net2290));
 sg13g2_tiehi \mem.mem_internal.code_mem[205][3]$_SDFFCE_PN0P__2291  (.L_HI(net2291));
 sg13g2_tiehi \mem.mem_internal.code_mem[205][4]$_SDFFCE_PN0P__2292  (.L_HI(net2292));
 sg13g2_tiehi \mem.mem_internal.code_mem[205][5]$_SDFFCE_PN0P__2293  (.L_HI(net2293));
 sg13g2_tiehi \mem.mem_internal.code_mem[205][6]$_SDFFCE_PN0P__2294  (.L_HI(net2294));
 sg13g2_tiehi \mem.mem_internal.code_mem[205][7]$_SDFFCE_PN0P__2295  (.L_HI(net2295));
 sg13g2_tiehi \mem.mem_internal.code_mem[206][0]$_SDFFCE_PN0P__2296  (.L_HI(net2296));
 sg13g2_tiehi \mem.mem_internal.code_mem[206][1]$_SDFFCE_PN0P__2297  (.L_HI(net2297));
 sg13g2_tiehi \mem.mem_internal.code_mem[206][2]$_SDFFCE_PN0P__2298  (.L_HI(net2298));
 sg13g2_tiehi \mem.mem_internal.code_mem[206][3]$_SDFFCE_PN0P__2299  (.L_HI(net2299));
 sg13g2_tiehi \mem.mem_internal.code_mem[206][4]$_SDFFCE_PN0P__2300  (.L_HI(net2300));
 sg13g2_tiehi \mem.mem_internal.code_mem[206][5]$_SDFFCE_PN0P__2301  (.L_HI(net2301));
 sg13g2_tiehi \mem.mem_internal.code_mem[206][6]$_SDFFCE_PN0P__2302  (.L_HI(net2302));
 sg13g2_tiehi \mem.mem_internal.code_mem[206][7]$_SDFFCE_PN0P__2303  (.L_HI(net2303));
 sg13g2_tiehi \mem.mem_internal.code_mem[207][0]$_SDFFCE_PN0P__2304  (.L_HI(net2304));
 sg13g2_tiehi \mem.mem_internal.code_mem[207][1]$_SDFFCE_PN0P__2305  (.L_HI(net2305));
 sg13g2_tiehi \mem.mem_internal.code_mem[207][2]$_SDFFCE_PN0P__2306  (.L_HI(net2306));
 sg13g2_tiehi \mem.mem_internal.code_mem[207][3]$_SDFFCE_PN0P__2307  (.L_HI(net2307));
 sg13g2_tiehi \mem.mem_internal.code_mem[207][4]$_SDFFCE_PN0P__2308  (.L_HI(net2308));
 sg13g2_tiehi \mem.mem_internal.code_mem[207][5]$_SDFFCE_PN0P__2309  (.L_HI(net2309));
 sg13g2_tiehi \mem.mem_internal.code_mem[207][6]$_SDFFCE_PN0P__2310  (.L_HI(net2310));
 sg13g2_tiehi \mem.mem_internal.code_mem[207][7]$_SDFFCE_PN0P__2311  (.L_HI(net2311));
 sg13g2_tiehi \mem.mem_internal.code_mem[208][0]$_SDFFCE_PN0P__2312  (.L_HI(net2312));
 sg13g2_tiehi \mem.mem_internal.code_mem[208][1]$_SDFFCE_PN0P__2313  (.L_HI(net2313));
 sg13g2_tiehi \mem.mem_internal.code_mem[208][2]$_SDFFCE_PN0P__2314  (.L_HI(net2314));
 sg13g2_tiehi \mem.mem_internal.code_mem[208][3]$_SDFFCE_PN0P__2315  (.L_HI(net2315));
 sg13g2_tiehi \mem.mem_internal.code_mem[208][4]$_SDFFCE_PN0P__2316  (.L_HI(net2316));
 sg13g2_tiehi \mem.mem_internal.code_mem[208][5]$_SDFFCE_PN0P__2317  (.L_HI(net2317));
 sg13g2_tiehi \mem.mem_internal.code_mem[208][6]$_SDFFCE_PN0P__2318  (.L_HI(net2318));
 sg13g2_tiehi \mem.mem_internal.code_mem[208][7]$_SDFFCE_PN0P__2319  (.L_HI(net2319));
 sg13g2_tiehi \mem.mem_internal.code_mem[209][0]$_SDFFCE_PN0P__2320  (.L_HI(net2320));
 sg13g2_tiehi \mem.mem_internal.code_mem[209][1]$_SDFFCE_PN0P__2321  (.L_HI(net2321));
 sg13g2_tiehi \mem.mem_internal.code_mem[209][2]$_SDFFCE_PN0P__2322  (.L_HI(net2322));
 sg13g2_tiehi \mem.mem_internal.code_mem[209][3]$_SDFFCE_PN0P__2323  (.L_HI(net2323));
 sg13g2_tiehi \mem.mem_internal.code_mem[209][4]$_SDFFCE_PN0P__2324  (.L_HI(net2324));
 sg13g2_tiehi \mem.mem_internal.code_mem[209][5]$_SDFFCE_PN0P__2325  (.L_HI(net2325));
 sg13g2_tiehi \mem.mem_internal.code_mem[209][6]$_SDFFCE_PN0P__2326  (.L_HI(net2326));
 sg13g2_tiehi \mem.mem_internal.code_mem[209][7]$_SDFFCE_PN0P__2327  (.L_HI(net2327));
 sg13g2_tiehi \mem.mem_internal.code_mem[20][0]$_SDFFCE_PN0P__2328  (.L_HI(net2328));
 sg13g2_tiehi \mem.mem_internal.code_mem[20][1]$_SDFFCE_PN0P__2329  (.L_HI(net2329));
 sg13g2_tiehi \mem.mem_internal.code_mem[20][2]$_SDFFCE_PN0P__2330  (.L_HI(net2330));
 sg13g2_tiehi \mem.mem_internal.code_mem[20][3]$_SDFFCE_PN0P__2331  (.L_HI(net2331));
 sg13g2_tiehi \mem.mem_internal.code_mem[20][4]$_SDFFCE_PN0P__2332  (.L_HI(net2332));
 sg13g2_tiehi \mem.mem_internal.code_mem[20][5]$_SDFFCE_PN0P__2333  (.L_HI(net2333));
 sg13g2_tiehi \mem.mem_internal.code_mem[20][6]$_SDFFCE_PN0P__2334  (.L_HI(net2334));
 sg13g2_tiehi \mem.mem_internal.code_mem[20][7]$_SDFFCE_PN0P__2335  (.L_HI(net2335));
 sg13g2_tiehi \mem.mem_internal.code_mem[210][0]$_SDFFCE_PN0P__2336  (.L_HI(net2336));
 sg13g2_tiehi \mem.mem_internal.code_mem[210][1]$_SDFFCE_PN0P__2337  (.L_HI(net2337));
 sg13g2_tiehi \mem.mem_internal.code_mem[210][2]$_SDFFCE_PN0P__2338  (.L_HI(net2338));
 sg13g2_tiehi \mem.mem_internal.code_mem[210][3]$_SDFFCE_PN0P__2339  (.L_HI(net2339));
 sg13g2_tiehi \mem.mem_internal.code_mem[210][4]$_SDFFCE_PN0P__2340  (.L_HI(net2340));
 sg13g2_tiehi \mem.mem_internal.code_mem[210][5]$_SDFFCE_PN0P__2341  (.L_HI(net2341));
 sg13g2_tiehi \mem.mem_internal.code_mem[210][6]$_SDFFCE_PN0P__2342  (.L_HI(net2342));
 sg13g2_tiehi \mem.mem_internal.code_mem[210][7]$_SDFFCE_PN0P__2343  (.L_HI(net2343));
 sg13g2_tiehi \mem.mem_internal.code_mem[211][0]$_SDFFCE_PN0P__2344  (.L_HI(net2344));
 sg13g2_tiehi \mem.mem_internal.code_mem[211][1]$_SDFFCE_PN0P__2345  (.L_HI(net2345));
 sg13g2_tiehi \mem.mem_internal.code_mem[211][2]$_SDFFCE_PN0P__2346  (.L_HI(net2346));
 sg13g2_tiehi \mem.mem_internal.code_mem[211][3]$_SDFFCE_PN0P__2347  (.L_HI(net2347));
 sg13g2_tiehi \mem.mem_internal.code_mem[211][4]$_SDFFCE_PN0P__2348  (.L_HI(net2348));
 sg13g2_tiehi \mem.mem_internal.code_mem[211][5]$_SDFFCE_PN0P__2349  (.L_HI(net2349));
 sg13g2_tiehi \mem.mem_internal.code_mem[211][6]$_SDFFCE_PN0P__2350  (.L_HI(net2350));
 sg13g2_tiehi \mem.mem_internal.code_mem[211][7]$_SDFFCE_PN0P__2351  (.L_HI(net2351));
 sg13g2_tiehi \mem.mem_internal.code_mem[212][0]$_SDFFCE_PN0P__2352  (.L_HI(net2352));
 sg13g2_tiehi \mem.mem_internal.code_mem[212][1]$_SDFFCE_PN0P__2353  (.L_HI(net2353));
 sg13g2_tiehi \mem.mem_internal.code_mem[212][2]$_SDFFCE_PN0P__2354  (.L_HI(net2354));
 sg13g2_tiehi \mem.mem_internal.code_mem[212][3]$_SDFFCE_PN0P__2355  (.L_HI(net2355));
 sg13g2_tiehi \mem.mem_internal.code_mem[212][4]$_SDFFCE_PN0P__2356  (.L_HI(net2356));
 sg13g2_tiehi \mem.mem_internal.code_mem[212][5]$_SDFFCE_PN0P__2357  (.L_HI(net2357));
 sg13g2_tiehi \mem.mem_internal.code_mem[212][6]$_SDFFCE_PN0P__2358  (.L_HI(net2358));
 sg13g2_tiehi \mem.mem_internal.code_mem[212][7]$_SDFFCE_PN0P__2359  (.L_HI(net2359));
 sg13g2_tiehi \mem.mem_internal.code_mem[213][0]$_SDFFCE_PN0P__2360  (.L_HI(net2360));
 sg13g2_tiehi \mem.mem_internal.code_mem[213][1]$_SDFFCE_PN0P__2361  (.L_HI(net2361));
 sg13g2_tiehi \mem.mem_internal.code_mem[213][2]$_SDFFCE_PN0P__2362  (.L_HI(net2362));
 sg13g2_tiehi \mem.mem_internal.code_mem[213][3]$_SDFFCE_PN0P__2363  (.L_HI(net2363));
 sg13g2_tiehi \mem.mem_internal.code_mem[213][4]$_SDFFCE_PN0P__2364  (.L_HI(net2364));
 sg13g2_tiehi \mem.mem_internal.code_mem[213][5]$_SDFFCE_PN0P__2365  (.L_HI(net2365));
 sg13g2_tiehi \mem.mem_internal.code_mem[213][6]$_SDFFCE_PN0P__2366  (.L_HI(net2366));
 sg13g2_tiehi \mem.mem_internal.code_mem[213][7]$_SDFFCE_PN0P__2367  (.L_HI(net2367));
 sg13g2_tiehi \mem.mem_internal.code_mem[214][0]$_SDFFCE_PN0P__2368  (.L_HI(net2368));
 sg13g2_tiehi \mem.mem_internal.code_mem[214][1]$_SDFFCE_PN0P__2369  (.L_HI(net2369));
 sg13g2_tiehi \mem.mem_internal.code_mem[214][2]$_SDFFCE_PN0P__2370  (.L_HI(net2370));
 sg13g2_tiehi \mem.mem_internal.code_mem[214][3]$_SDFFCE_PN0P__2371  (.L_HI(net2371));
 sg13g2_tiehi \mem.mem_internal.code_mem[214][4]$_SDFFCE_PN0P__2372  (.L_HI(net2372));
 sg13g2_tiehi \mem.mem_internal.code_mem[214][5]$_SDFFCE_PN0P__2373  (.L_HI(net2373));
 sg13g2_tiehi \mem.mem_internal.code_mem[214][6]$_SDFFCE_PN0P__2374  (.L_HI(net2374));
 sg13g2_tiehi \mem.mem_internal.code_mem[214][7]$_SDFFCE_PN0P__2375  (.L_HI(net2375));
 sg13g2_tiehi \mem.mem_internal.code_mem[215][0]$_SDFFCE_PN0P__2376  (.L_HI(net2376));
 sg13g2_tiehi \mem.mem_internal.code_mem[215][1]$_SDFFCE_PN0P__2377  (.L_HI(net2377));
 sg13g2_tiehi \mem.mem_internal.code_mem[215][2]$_SDFFCE_PN0P__2378  (.L_HI(net2378));
 sg13g2_tiehi \mem.mem_internal.code_mem[215][3]$_SDFFCE_PN0P__2379  (.L_HI(net2379));
 sg13g2_tiehi \mem.mem_internal.code_mem[215][4]$_SDFFCE_PN0P__2380  (.L_HI(net2380));
 sg13g2_tiehi \mem.mem_internal.code_mem[215][5]$_SDFFCE_PN0P__2381  (.L_HI(net2381));
 sg13g2_tiehi \mem.mem_internal.code_mem[215][6]$_SDFFCE_PN0P__2382  (.L_HI(net2382));
 sg13g2_tiehi \mem.mem_internal.code_mem[215][7]$_SDFFCE_PN0P__2383  (.L_HI(net2383));
 sg13g2_tiehi \mem.mem_internal.code_mem[216][0]$_SDFFCE_PN0P__2384  (.L_HI(net2384));
 sg13g2_tiehi \mem.mem_internal.code_mem[216][1]$_SDFFCE_PN0P__2385  (.L_HI(net2385));
 sg13g2_tiehi \mem.mem_internal.code_mem[216][2]$_SDFFCE_PN0P__2386  (.L_HI(net2386));
 sg13g2_tiehi \mem.mem_internal.code_mem[216][3]$_SDFFCE_PN0P__2387  (.L_HI(net2387));
 sg13g2_tiehi \mem.mem_internal.code_mem[216][4]$_SDFFCE_PN0P__2388  (.L_HI(net2388));
 sg13g2_tiehi \mem.mem_internal.code_mem[216][5]$_SDFFCE_PN0P__2389  (.L_HI(net2389));
 sg13g2_tiehi \mem.mem_internal.code_mem[216][6]$_SDFFCE_PN0P__2390  (.L_HI(net2390));
 sg13g2_tiehi \mem.mem_internal.code_mem[216][7]$_SDFFCE_PN0P__2391  (.L_HI(net2391));
 sg13g2_tiehi \mem.mem_internal.code_mem[217][0]$_SDFFCE_PN0P__2392  (.L_HI(net2392));
 sg13g2_tiehi \mem.mem_internal.code_mem[217][1]$_SDFFCE_PN0P__2393  (.L_HI(net2393));
 sg13g2_tiehi \mem.mem_internal.code_mem[217][2]$_SDFFCE_PN0P__2394  (.L_HI(net2394));
 sg13g2_tiehi \mem.mem_internal.code_mem[217][3]$_SDFFCE_PN0P__2395  (.L_HI(net2395));
 sg13g2_tiehi \mem.mem_internal.code_mem[217][4]$_SDFFCE_PN0P__2396  (.L_HI(net2396));
 sg13g2_tiehi \mem.mem_internal.code_mem[217][5]$_SDFFCE_PN0P__2397  (.L_HI(net2397));
 sg13g2_tiehi \mem.mem_internal.code_mem[217][6]$_SDFFCE_PN0P__2398  (.L_HI(net2398));
 sg13g2_tiehi \mem.mem_internal.code_mem[217][7]$_SDFFCE_PN0P__2399  (.L_HI(net2399));
 sg13g2_tiehi \mem.mem_internal.code_mem[218][0]$_SDFFCE_PN0P__2400  (.L_HI(net2400));
 sg13g2_tiehi \mem.mem_internal.code_mem[218][1]$_SDFFCE_PN0P__2401  (.L_HI(net2401));
 sg13g2_tiehi \mem.mem_internal.code_mem[218][2]$_SDFFCE_PN0P__2402  (.L_HI(net2402));
 sg13g2_tiehi \mem.mem_internal.code_mem[218][3]$_SDFFCE_PN0P__2403  (.L_HI(net2403));
 sg13g2_tiehi \mem.mem_internal.code_mem[218][4]$_SDFFCE_PN0P__2404  (.L_HI(net2404));
 sg13g2_tiehi \mem.mem_internal.code_mem[218][5]$_SDFFCE_PN0P__2405  (.L_HI(net2405));
 sg13g2_tiehi \mem.mem_internal.code_mem[218][6]$_SDFFCE_PN0P__2406  (.L_HI(net2406));
 sg13g2_tiehi \mem.mem_internal.code_mem[218][7]$_SDFFCE_PN0P__2407  (.L_HI(net2407));
 sg13g2_tiehi \mem.mem_internal.code_mem[219][0]$_SDFFCE_PN0P__2408  (.L_HI(net2408));
 sg13g2_tiehi \mem.mem_internal.code_mem[219][1]$_SDFFCE_PN0P__2409  (.L_HI(net2409));
 sg13g2_tiehi \mem.mem_internal.code_mem[219][2]$_SDFFCE_PN0P__2410  (.L_HI(net2410));
 sg13g2_tiehi \mem.mem_internal.code_mem[219][3]$_SDFFCE_PN0P__2411  (.L_HI(net2411));
 sg13g2_tiehi \mem.mem_internal.code_mem[219][4]$_SDFFCE_PN0P__2412  (.L_HI(net2412));
 sg13g2_tiehi \mem.mem_internal.code_mem[219][5]$_SDFFCE_PN0P__2413  (.L_HI(net2413));
 sg13g2_tiehi \mem.mem_internal.code_mem[219][6]$_SDFFCE_PN0P__2414  (.L_HI(net2414));
 sg13g2_tiehi \mem.mem_internal.code_mem[219][7]$_SDFFCE_PN0P__2415  (.L_HI(net2415));
 sg13g2_tiehi \mem.mem_internal.code_mem[21][0]$_SDFFCE_PN0P__2416  (.L_HI(net2416));
 sg13g2_tiehi \mem.mem_internal.code_mem[21][1]$_SDFFCE_PN0P__2417  (.L_HI(net2417));
 sg13g2_tiehi \mem.mem_internal.code_mem[21][2]$_SDFFCE_PN0P__2418  (.L_HI(net2418));
 sg13g2_tiehi \mem.mem_internal.code_mem[21][3]$_SDFFCE_PN0P__2419  (.L_HI(net2419));
 sg13g2_tiehi \mem.mem_internal.code_mem[21][4]$_SDFFCE_PN0P__2420  (.L_HI(net2420));
 sg13g2_tiehi \mem.mem_internal.code_mem[21][5]$_SDFFCE_PN0P__2421  (.L_HI(net2421));
 sg13g2_tiehi \mem.mem_internal.code_mem[21][6]$_SDFFCE_PN0P__2422  (.L_HI(net2422));
 sg13g2_tiehi \mem.mem_internal.code_mem[21][7]$_SDFFCE_PN0P__2423  (.L_HI(net2423));
 sg13g2_tiehi \mem.mem_internal.code_mem[220][0]$_SDFFCE_PN0P__2424  (.L_HI(net2424));
 sg13g2_tiehi \mem.mem_internal.code_mem[220][1]$_SDFFCE_PN0P__2425  (.L_HI(net2425));
 sg13g2_tiehi \mem.mem_internal.code_mem[220][2]$_SDFFCE_PN0P__2426  (.L_HI(net2426));
 sg13g2_tiehi \mem.mem_internal.code_mem[220][3]$_SDFFCE_PN0P__2427  (.L_HI(net2427));
 sg13g2_tiehi \mem.mem_internal.code_mem[220][4]$_SDFFCE_PN0P__2428  (.L_HI(net2428));
 sg13g2_tiehi \mem.mem_internal.code_mem[220][5]$_SDFFCE_PN0P__2429  (.L_HI(net2429));
 sg13g2_tiehi \mem.mem_internal.code_mem[220][6]$_SDFFCE_PN0P__2430  (.L_HI(net2430));
 sg13g2_tiehi \mem.mem_internal.code_mem[220][7]$_SDFFCE_PN0P__2431  (.L_HI(net2431));
 sg13g2_tiehi \mem.mem_internal.code_mem[221][0]$_SDFFCE_PN0P__2432  (.L_HI(net2432));
 sg13g2_tiehi \mem.mem_internal.code_mem[221][1]$_SDFFCE_PN0P__2433  (.L_HI(net2433));
 sg13g2_tiehi \mem.mem_internal.code_mem[221][2]$_SDFFCE_PN0P__2434  (.L_HI(net2434));
 sg13g2_tiehi \mem.mem_internal.code_mem[221][3]$_SDFFCE_PN0P__2435  (.L_HI(net2435));
 sg13g2_tiehi \mem.mem_internal.code_mem[221][4]$_SDFFCE_PN0P__2436  (.L_HI(net2436));
 sg13g2_tiehi \mem.mem_internal.code_mem[221][5]$_SDFFCE_PN0P__2437  (.L_HI(net2437));
 sg13g2_tiehi \mem.mem_internal.code_mem[221][6]$_SDFFCE_PN0P__2438  (.L_HI(net2438));
 sg13g2_tiehi \mem.mem_internal.code_mem[221][7]$_SDFFCE_PN0P__2439  (.L_HI(net2439));
 sg13g2_tiehi \mem.mem_internal.code_mem[222][0]$_SDFFCE_PN0P__2440  (.L_HI(net2440));
 sg13g2_tiehi \mem.mem_internal.code_mem[222][1]$_SDFFCE_PN0P__2441  (.L_HI(net2441));
 sg13g2_tiehi \mem.mem_internal.code_mem[222][2]$_SDFFCE_PN0P__2442  (.L_HI(net2442));
 sg13g2_tiehi \mem.mem_internal.code_mem[222][3]$_SDFFCE_PN0P__2443  (.L_HI(net2443));
 sg13g2_tiehi \mem.mem_internal.code_mem[222][4]$_SDFFCE_PN0P__2444  (.L_HI(net2444));
 sg13g2_tiehi \mem.mem_internal.code_mem[222][5]$_SDFFCE_PN0P__2445  (.L_HI(net2445));
 sg13g2_tiehi \mem.mem_internal.code_mem[222][6]$_SDFFCE_PN0P__2446  (.L_HI(net2446));
 sg13g2_tiehi \mem.mem_internal.code_mem[222][7]$_SDFFCE_PN0P__2447  (.L_HI(net2447));
 sg13g2_tiehi \mem.mem_internal.code_mem[223][0]$_SDFFCE_PN0P__2448  (.L_HI(net2448));
 sg13g2_tiehi \mem.mem_internal.code_mem[223][1]$_SDFFCE_PN0P__2449  (.L_HI(net2449));
 sg13g2_tiehi \mem.mem_internal.code_mem[223][2]$_SDFFCE_PN0P__2450  (.L_HI(net2450));
 sg13g2_tiehi \mem.mem_internal.code_mem[223][3]$_SDFFCE_PN0P__2451  (.L_HI(net2451));
 sg13g2_tiehi \mem.mem_internal.code_mem[223][4]$_SDFFCE_PN0P__2452  (.L_HI(net2452));
 sg13g2_tiehi \mem.mem_internal.code_mem[223][5]$_SDFFCE_PN0P__2453  (.L_HI(net2453));
 sg13g2_tiehi \mem.mem_internal.code_mem[223][6]$_SDFFCE_PN0P__2454  (.L_HI(net2454));
 sg13g2_tiehi \mem.mem_internal.code_mem[223][7]$_SDFFCE_PN0P__2455  (.L_HI(net2455));
 sg13g2_tiehi \mem.mem_internal.code_mem[224][0]$_SDFFCE_PN0P__2456  (.L_HI(net2456));
 sg13g2_tiehi \mem.mem_internal.code_mem[224][1]$_SDFFCE_PN0P__2457  (.L_HI(net2457));
 sg13g2_tiehi \mem.mem_internal.code_mem[224][2]$_SDFFCE_PN0P__2458  (.L_HI(net2458));
 sg13g2_tiehi \mem.mem_internal.code_mem[224][3]$_SDFFCE_PN0P__2459  (.L_HI(net2459));
 sg13g2_tiehi \mem.mem_internal.code_mem[224][4]$_SDFFCE_PN0P__2460  (.L_HI(net2460));
 sg13g2_tiehi \mem.mem_internal.code_mem[224][5]$_SDFFCE_PN0P__2461  (.L_HI(net2461));
 sg13g2_tiehi \mem.mem_internal.code_mem[224][6]$_SDFFCE_PN0P__2462  (.L_HI(net2462));
 sg13g2_tiehi \mem.mem_internal.code_mem[224][7]$_SDFFCE_PN0P__2463  (.L_HI(net2463));
 sg13g2_tiehi \mem.mem_internal.code_mem[225][0]$_SDFFCE_PN0P__2464  (.L_HI(net2464));
 sg13g2_tiehi \mem.mem_internal.code_mem[225][1]$_SDFFCE_PN0P__2465  (.L_HI(net2465));
 sg13g2_tiehi \mem.mem_internal.code_mem[225][2]$_SDFFCE_PN0P__2466  (.L_HI(net2466));
 sg13g2_tiehi \mem.mem_internal.code_mem[225][3]$_SDFFCE_PN0P__2467  (.L_HI(net2467));
 sg13g2_tiehi \mem.mem_internal.code_mem[225][4]$_SDFFCE_PN0P__2468  (.L_HI(net2468));
 sg13g2_tiehi \mem.mem_internal.code_mem[225][5]$_SDFFCE_PN0P__2469  (.L_HI(net2469));
 sg13g2_tiehi \mem.mem_internal.code_mem[225][6]$_SDFFCE_PN0P__2470  (.L_HI(net2470));
 sg13g2_tiehi \mem.mem_internal.code_mem[225][7]$_SDFFCE_PN0P__2471  (.L_HI(net2471));
 sg13g2_tiehi \mem.mem_internal.code_mem[226][0]$_SDFFCE_PN0P__2472  (.L_HI(net2472));
 sg13g2_tiehi \mem.mem_internal.code_mem[226][1]$_SDFFCE_PN0P__2473  (.L_HI(net2473));
 sg13g2_tiehi \mem.mem_internal.code_mem[226][2]$_SDFFCE_PN0P__2474  (.L_HI(net2474));
 sg13g2_tiehi \mem.mem_internal.code_mem[226][3]$_SDFFCE_PN0P__2475  (.L_HI(net2475));
 sg13g2_tiehi \mem.mem_internal.code_mem[226][4]$_SDFFCE_PN0P__2476  (.L_HI(net2476));
 sg13g2_tiehi \mem.mem_internal.code_mem[226][5]$_SDFFCE_PN0P__2477  (.L_HI(net2477));
 sg13g2_tiehi \mem.mem_internal.code_mem[226][6]$_SDFFCE_PN0P__2478  (.L_HI(net2478));
 sg13g2_tiehi \mem.mem_internal.code_mem[226][7]$_SDFFCE_PN0P__2479  (.L_HI(net2479));
 sg13g2_tiehi \mem.mem_internal.code_mem[227][0]$_SDFFCE_PN0P__2480  (.L_HI(net2480));
 sg13g2_tiehi \mem.mem_internal.code_mem[227][1]$_SDFFCE_PN0P__2481  (.L_HI(net2481));
 sg13g2_tiehi \mem.mem_internal.code_mem[227][2]$_SDFFCE_PN0P__2482  (.L_HI(net2482));
 sg13g2_tiehi \mem.mem_internal.code_mem[227][3]$_SDFFCE_PN0P__2483  (.L_HI(net2483));
 sg13g2_tiehi \mem.mem_internal.code_mem[227][4]$_SDFFCE_PN0P__2484  (.L_HI(net2484));
 sg13g2_tiehi \mem.mem_internal.code_mem[227][5]$_SDFFCE_PN0P__2485  (.L_HI(net2485));
 sg13g2_tiehi \mem.mem_internal.code_mem[227][6]$_SDFFCE_PN0P__2486  (.L_HI(net2486));
 sg13g2_tiehi \mem.mem_internal.code_mem[227][7]$_SDFFCE_PN0P__2487  (.L_HI(net2487));
 sg13g2_tiehi \mem.mem_internal.code_mem[228][0]$_SDFFCE_PN0P__2488  (.L_HI(net2488));
 sg13g2_tiehi \mem.mem_internal.code_mem[228][1]$_SDFFCE_PN0P__2489  (.L_HI(net2489));
 sg13g2_tiehi \mem.mem_internal.code_mem[228][2]$_SDFFCE_PN0P__2490  (.L_HI(net2490));
 sg13g2_tiehi \mem.mem_internal.code_mem[228][3]$_SDFFCE_PN0P__2491  (.L_HI(net2491));
 sg13g2_tiehi \mem.mem_internal.code_mem[228][4]$_SDFFCE_PN0P__2492  (.L_HI(net2492));
 sg13g2_tiehi \mem.mem_internal.code_mem[228][5]$_SDFFCE_PN0P__2493  (.L_HI(net2493));
 sg13g2_tiehi \mem.mem_internal.code_mem[228][6]$_SDFFCE_PN0P__2494  (.L_HI(net2494));
 sg13g2_tiehi \mem.mem_internal.code_mem[228][7]$_SDFFCE_PN0P__2495  (.L_HI(net2495));
 sg13g2_tiehi \mem.mem_internal.code_mem[229][0]$_SDFFCE_PN0P__2496  (.L_HI(net2496));
 sg13g2_tiehi \mem.mem_internal.code_mem[229][1]$_SDFFCE_PN0P__2497  (.L_HI(net2497));
 sg13g2_tiehi \mem.mem_internal.code_mem[229][2]$_SDFFCE_PN0P__2498  (.L_HI(net2498));
 sg13g2_tiehi \mem.mem_internal.code_mem[229][3]$_SDFFCE_PN0P__2499  (.L_HI(net2499));
 sg13g2_tiehi \mem.mem_internal.code_mem[229][4]$_SDFFCE_PN0P__2500  (.L_HI(net2500));
 sg13g2_tiehi \mem.mem_internal.code_mem[229][5]$_SDFFCE_PN0P__2501  (.L_HI(net2501));
 sg13g2_tiehi \mem.mem_internal.code_mem[229][6]$_SDFFCE_PN0P__2502  (.L_HI(net2502));
 sg13g2_tiehi \mem.mem_internal.code_mem[229][7]$_SDFFCE_PN0P__2503  (.L_HI(net2503));
 sg13g2_tiehi \mem.mem_internal.code_mem[22][0]$_SDFFCE_PN0P__2504  (.L_HI(net2504));
 sg13g2_tiehi \mem.mem_internal.code_mem[22][1]$_SDFFCE_PN0P__2505  (.L_HI(net2505));
 sg13g2_tiehi \mem.mem_internal.code_mem[22][2]$_SDFFCE_PN0P__2506  (.L_HI(net2506));
 sg13g2_tiehi \mem.mem_internal.code_mem[22][3]$_SDFFCE_PN0P__2507  (.L_HI(net2507));
 sg13g2_tiehi \mem.mem_internal.code_mem[22][4]$_SDFFCE_PN0P__2508  (.L_HI(net2508));
 sg13g2_tiehi \mem.mem_internal.code_mem[22][5]$_SDFFCE_PN0P__2509  (.L_HI(net2509));
 sg13g2_tiehi \mem.mem_internal.code_mem[22][6]$_SDFFCE_PN0P__2510  (.L_HI(net2510));
 sg13g2_tiehi \mem.mem_internal.code_mem[22][7]$_SDFFCE_PN0P__2511  (.L_HI(net2511));
 sg13g2_tiehi \mem.mem_internal.code_mem[230][0]$_SDFFCE_PN0P__2512  (.L_HI(net2512));
 sg13g2_tiehi \mem.mem_internal.code_mem[230][1]$_SDFFCE_PN0P__2513  (.L_HI(net2513));
 sg13g2_tiehi \mem.mem_internal.code_mem[230][2]$_SDFFCE_PN0P__2514  (.L_HI(net2514));
 sg13g2_tiehi \mem.mem_internal.code_mem[230][3]$_SDFFCE_PN0P__2515  (.L_HI(net2515));
 sg13g2_tiehi \mem.mem_internal.code_mem[230][4]$_SDFFCE_PN0P__2516  (.L_HI(net2516));
 sg13g2_tiehi \mem.mem_internal.code_mem[230][5]$_SDFFCE_PN0P__2517  (.L_HI(net2517));
 sg13g2_tiehi \mem.mem_internal.code_mem[230][6]$_SDFFCE_PN0P__2518  (.L_HI(net2518));
 sg13g2_tiehi \mem.mem_internal.code_mem[230][7]$_SDFFCE_PN0P__2519  (.L_HI(net2519));
 sg13g2_tiehi \mem.mem_internal.code_mem[231][0]$_SDFFCE_PN0P__2520  (.L_HI(net2520));
 sg13g2_tiehi \mem.mem_internal.code_mem[231][1]$_SDFFCE_PN0P__2521  (.L_HI(net2521));
 sg13g2_tiehi \mem.mem_internal.code_mem[231][2]$_SDFFCE_PN0P__2522  (.L_HI(net2522));
 sg13g2_tiehi \mem.mem_internal.code_mem[231][3]$_SDFFCE_PN0P__2523  (.L_HI(net2523));
 sg13g2_tiehi \mem.mem_internal.code_mem[231][4]$_SDFFCE_PN0P__2524  (.L_HI(net2524));
 sg13g2_tiehi \mem.mem_internal.code_mem[231][5]$_SDFFCE_PN0P__2525  (.L_HI(net2525));
 sg13g2_tiehi \mem.mem_internal.code_mem[231][6]$_SDFFCE_PN0P__2526  (.L_HI(net2526));
 sg13g2_tiehi \mem.mem_internal.code_mem[231][7]$_SDFFCE_PN0P__2527  (.L_HI(net2527));
 sg13g2_tiehi \mem.mem_internal.code_mem[232][0]$_SDFFCE_PN0P__2528  (.L_HI(net2528));
 sg13g2_tiehi \mem.mem_internal.code_mem[232][1]$_SDFFCE_PN0P__2529  (.L_HI(net2529));
 sg13g2_tiehi \mem.mem_internal.code_mem[232][2]$_SDFFCE_PN0P__2530  (.L_HI(net2530));
 sg13g2_tiehi \mem.mem_internal.code_mem[232][3]$_SDFFCE_PN0P__2531  (.L_HI(net2531));
 sg13g2_tiehi \mem.mem_internal.code_mem[232][4]$_SDFFCE_PN0P__2532  (.L_HI(net2532));
 sg13g2_tiehi \mem.mem_internal.code_mem[232][5]$_SDFFCE_PN0P__2533  (.L_HI(net2533));
 sg13g2_tiehi \mem.mem_internal.code_mem[232][6]$_SDFFCE_PN0P__2534  (.L_HI(net2534));
 sg13g2_tiehi \mem.mem_internal.code_mem[232][7]$_SDFFCE_PN0P__2535  (.L_HI(net2535));
 sg13g2_tiehi \mem.mem_internal.code_mem[233][0]$_SDFFCE_PN0P__2536  (.L_HI(net2536));
 sg13g2_tiehi \mem.mem_internal.code_mem[233][1]$_SDFFCE_PN0P__2537  (.L_HI(net2537));
 sg13g2_tiehi \mem.mem_internal.code_mem[233][2]$_SDFFCE_PN0P__2538  (.L_HI(net2538));
 sg13g2_tiehi \mem.mem_internal.code_mem[233][3]$_SDFFCE_PN0P__2539  (.L_HI(net2539));
 sg13g2_tiehi \mem.mem_internal.code_mem[233][4]$_SDFFCE_PN0P__2540  (.L_HI(net2540));
 sg13g2_tiehi \mem.mem_internal.code_mem[233][5]$_SDFFCE_PN0P__2541  (.L_HI(net2541));
 sg13g2_tiehi \mem.mem_internal.code_mem[233][6]$_SDFFCE_PN0P__2542  (.L_HI(net2542));
 sg13g2_tiehi \mem.mem_internal.code_mem[233][7]$_SDFFCE_PN0P__2543  (.L_HI(net2543));
 sg13g2_tiehi \mem.mem_internal.code_mem[234][0]$_SDFFCE_PN0P__2544  (.L_HI(net2544));
 sg13g2_tiehi \mem.mem_internal.code_mem[234][1]$_SDFFCE_PN0P__2545  (.L_HI(net2545));
 sg13g2_tiehi \mem.mem_internal.code_mem[234][2]$_SDFFCE_PN0P__2546  (.L_HI(net2546));
 sg13g2_tiehi \mem.mem_internal.code_mem[234][3]$_SDFFCE_PN0P__2547  (.L_HI(net2547));
 sg13g2_tiehi \mem.mem_internal.code_mem[234][4]$_SDFFCE_PN0P__2548  (.L_HI(net2548));
 sg13g2_tiehi \mem.mem_internal.code_mem[234][5]$_SDFFCE_PN0P__2549  (.L_HI(net2549));
 sg13g2_tiehi \mem.mem_internal.code_mem[234][6]$_SDFFCE_PN0P__2550  (.L_HI(net2550));
 sg13g2_tiehi \mem.mem_internal.code_mem[234][7]$_SDFFCE_PN0P__2551  (.L_HI(net2551));
 sg13g2_tiehi \mem.mem_internal.code_mem[235][0]$_SDFFCE_PN0P__2552  (.L_HI(net2552));
 sg13g2_tiehi \mem.mem_internal.code_mem[235][1]$_SDFFCE_PN0P__2553  (.L_HI(net2553));
 sg13g2_tiehi \mem.mem_internal.code_mem[235][2]$_SDFFCE_PN0P__2554  (.L_HI(net2554));
 sg13g2_tiehi \mem.mem_internal.code_mem[235][3]$_SDFFCE_PN0P__2555  (.L_HI(net2555));
 sg13g2_tiehi \mem.mem_internal.code_mem[235][4]$_SDFFCE_PN0P__2556  (.L_HI(net2556));
 sg13g2_tiehi \mem.mem_internal.code_mem[235][5]$_SDFFCE_PN0P__2557  (.L_HI(net2557));
 sg13g2_tiehi \mem.mem_internal.code_mem[235][6]$_SDFFCE_PN0P__2558  (.L_HI(net2558));
 sg13g2_tiehi \mem.mem_internal.code_mem[235][7]$_SDFFCE_PN0P__2559  (.L_HI(net2559));
 sg13g2_tiehi \mem.mem_internal.code_mem[236][0]$_SDFFCE_PN0P__2560  (.L_HI(net2560));
 sg13g2_tiehi \mem.mem_internal.code_mem[236][1]$_SDFFCE_PN0P__2561  (.L_HI(net2561));
 sg13g2_tiehi \mem.mem_internal.code_mem[236][2]$_SDFFCE_PN0P__2562  (.L_HI(net2562));
 sg13g2_tiehi \mem.mem_internal.code_mem[236][3]$_SDFFCE_PN0P__2563  (.L_HI(net2563));
 sg13g2_tiehi \mem.mem_internal.code_mem[236][4]$_SDFFCE_PN0P__2564  (.L_HI(net2564));
 sg13g2_tiehi \mem.mem_internal.code_mem[236][5]$_SDFFCE_PN0P__2565  (.L_HI(net2565));
 sg13g2_tiehi \mem.mem_internal.code_mem[236][6]$_SDFFCE_PN0P__2566  (.L_HI(net2566));
 sg13g2_tiehi \mem.mem_internal.code_mem[236][7]$_SDFFCE_PN0P__2567  (.L_HI(net2567));
 sg13g2_tiehi \mem.mem_internal.code_mem[237][0]$_SDFFCE_PN0P__2568  (.L_HI(net2568));
 sg13g2_tiehi \mem.mem_internal.code_mem[237][1]$_SDFFCE_PN0P__2569  (.L_HI(net2569));
 sg13g2_tiehi \mem.mem_internal.code_mem[237][2]$_SDFFCE_PN0P__2570  (.L_HI(net2570));
 sg13g2_tiehi \mem.mem_internal.code_mem[237][3]$_SDFFCE_PN0P__2571  (.L_HI(net2571));
 sg13g2_tiehi \mem.mem_internal.code_mem[237][4]$_SDFFCE_PN0P__2572  (.L_HI(net2572));
 sg13g2_tiehi \mem.mem_internal.code_mem[237][5]$_SDFFCE_PN0P__2573  (.L_HI(net2573));
 sg13g2_tiehi \mem.mem_internal.code_mem[237][6]$_SDFFCE_PN0P__2574  (.L_HI(net2574));
 sg13g2_tiehi \mem.mem_internal.code_mem[237][7]$_SDFFCE_PN0P__2575  (.L_HI(net2575));
 sg13g2_tiehi \mem.mem_internal.code_mem[238][0]$_SDFFCE_PN0P__2576  (.L_HI(net2576));
 sg13g2_tiehi \mem.mem_internal.code_mem[238][1]$_SDFFCE_PN0P__2577  (.L_HI(net2577));
 sg13g2_tiehi \mem.mem_internal.code_mem[238][2]$_SDFFCE_PN0P__2578  (.L_HI(net2578));
 sg13g2_tiehi \mem.mem_internal.code_mem[238][3]$_SDFFCE_PN0P__2579  (.L_HI(net2579));
 sg13g2_tiehi \mem.mem_internal.code_mem[238][4]$_SDFFCE_PN0P__2580  (.L_HI(net2580));
 sg13g2_tiehi \mem.mem_internal.code_mem[238][5]$_SDFFCE_PN0P__2581  (.L_HI(net2581));
 sg13g2_tiehi \mem.mem_internal.code_mem[238][6]$_SDFFCE_PN0P__2582  (.L_HI(net2582));
 sg13g2_tiehi \mem.mem_internal.code_mem[238][7]$_SDFFCE_PN0P__2583  (.L_HI(net2583));
 sg13g2_tiehi \mem.mem_internal.code_mem[239][0]$_SDFFCE_PN0P__2584  (.L_HI(net2584));
 sg13g2_tiehi \mem.mem_internal.code_mem[239][1]$_SDFFCE_PN0P__2585  (.L_HI(net2585));
 sg13g2_tiehi \mem.mem_internal.code_mem[239][2]$_SDFFCE_PN0P__2586  (.L_HI(net2586));
 sg13g2_tiehi \mem.mem_internal.code_mem[239][3]$_SDFFCE_PN0P__2587  (.L_HI(net2587));
 sg13g2_tiehi \mem.mem_internal.code_mem[239][4]$_SDFFCE_PN0P__2588  (.L_HI(net2588));
 sg13g2_tiehi \mem.mem_internal.code_mem[239][5]$_SDFFCE_PN0P__2589  (.L_HI(net2589));
 sg13g2_tiehi \mem.mem_internal.code_mem[239][6]$_SDFFCE_PN0P__2590  (.L_HI(net2590));
 sg13g2_tiehi \mem.mem_internal.code_mem[239][7]$_SDFFCE_PN0P__2591  (.L_HI(net2591));
 sg13g2_tiehi \mem.mem_internal.code_mem[23][0]$_SDFFCE_PN0P__2592  (.L_HI(net2592));
 sg13g2_tiehi \mem.mem_internal.code_mem[23][1]$_SDFFCE_PN0P__2593  (.L_HI(net2593));
 sg13g2_tiehi \mem.mem_internal.code_mem[23][2]$_SDFFCE_PN0P__2594  (.L_HI(net2594));
 sg13g2_tiehi \mem.mem_internal.code_mem[23][3]$_SDFFCE_PN0P__2595  (.L_HI(net2595));
 sg13g2_tiehi \mem.mem_internal.code_mem[23][4]$_SDFFCE_PN0P__2596  (.L_HI(net2596));
 sg13g2_tiehi \mem.mem_internal.code_mem[23][5]$_SDFFCE_PN0P__2597  (.L_HI(net2597));
 sg13g2_tiehi \mem.mem_internal.code_mem[23][6]$_SDFFCE_PN0P__2598  (.L_HI(net2598));
 sg13g2_tiehi \mem.mem_internal.code_mem[23][7]$_SDFFCE_PN0P__2599  (.L_HI(net2599));
 sg13g2_tiehi \mem.mem_internal.code_mem[240][0]$_SDFFCE_PN0P__2600  (.L_HI(net2600));
 sg13g2_tiehi \mem.mem_internal.code_mem[240][1]$_SDFFCE_PN0P__2601  (.L_HI(net2601));
 sg13g2_tiehi \mem.mem_internal.code_mem[240][2]$_SDFFCE_PN0P__2602  (.L_HI(net2602));
 sg13g2_tiehi \mem.mem_internal.code_mem[240][3]$_SDFFCE_PN0P__2603  (.L_HI(net2603));
 sg13g2_tiehi \mem.mem_internal.code_mem[240][4]$_SDFFCE_PN0P__2604  (.L_HI(net2604));
 sg13g2_tiehi \mem.mem_internal.code_mem[240][5]$_SDFFCE_PN0P__2605  (.L_HI(net2605));
 sg13g2_tiehi \mem.mem_internal.code_mem[240][6]$_SDFFCE_PN0P__2606  (.L_HI(net2606));
 sg13g2_tiehi \mem.mem_internal.code_mem[240][7]$_SDFFCE_PN0P__2607  (.L_HI(net2607));
 sg13g2_tiehi \mem.mem_internal.code_mem[241][0]$_SDFFCE_PN0P__2608  (.L_HI(net2608));
 sg13g2_tiehi \mem.mem_internal.code_mem[241][1]$_SDFFCE_PN0P__2609  (.L_HI(net2609));
 sg13g2_tiehi \mem.mem_internal.code_mem[241][2]$_SDFFCE_PN0P__2610  (.L_HI(net2610));
 sg13g2_tiehi \mem.mem_internal.code_mem[241][3]$_SDFFCE_PN0P__2611  (.L_HI(net2611));
 sg13g2_tiehi \mem.mem_internal.code_mem[241][4]$_SDFFCE_PN0P__2612  (.L_HI(net2612));
 sg13g2_tiehi \mem.mem_internal.code_mem[241][5]$_SDFFCE_PN0P__2613  (.L_HI(net2613));
 sg13g2_tiehi \mem.mem_internal.code_mem[241][6]$_SDFFCE_PN0P__2614  (.L_HI(net2614));
 sg13g2_tiehi \mem.mem_internal.code_mem[241][7]$_SDFFCE_PN0P__2615  (.L_HI(net2615));
 sg13g2_tiehi \mem.mem_internal.code_mem[242][0]$_SDFFCE_PN0P__2616  (.L_HI(net2616));
 sg13g2_tiehi \mem.mem_internal.code_mem[242][1]$_SDFFCE_PN0P__2617  (.L_HI(net2617));
 sg13g2_tiehi \mem.mem_internal.code_mem[242][2]$_SDFFCE_PN0P__2618  (.L_HI(net2618));
 sg13g2_tiehi \mem.mem_internal.code_mem[242][3]$_SDFFCE_PN0P__2619  (.L_HI(net2619));
 sg13g2_tiehi \mem.mem_internal.code_mem[242][4]$_SDFFCE_PN0P__2620  (.L_HI(net2620));
 sg13g2_tiehi \mem.mem_internal.code_mem[242][5]$_SDFFCE_PN0P__2621  (.L_HI(net2621));
 sg13g2_tiehi \mem.mem_internal.code_mem[242][6]$_SDFFCE_PN0P__2622  (.L_HI(net2622));
 sg13g2_tiehi \mem.mem_internal.code_mem[242][7]$_SDFFCE_PN0P__2623  (.L_HI(net2623));
 sg13g2_tiehi \mem.mem_internal.code_mem[243][0]$_SDFFCE_PN0P__2624  (.L_HI(net2624));
 sg13g2_tiehi \mem.mem_internal.code_mem[243][1]$_SDFFCE_PN0P__2625  (.L_HI(net2625));
 sg13g2_tiehi \mem.mem_internal.code_mem[243][2]$_SDFFCE_PN0P__2626  (.L_HI(net2626));
 sg13g2_tiehi \mem.mem_internal.code_mem[243][3]$_SDFFCE_PN0P__2627  (.L_HI(net2627));
 sg13g2_tiehi \mem.mem_internal.code_mem[243][4]$_SDFFCE_PN0P__2628  (.L_HI(net2628));
 sg13g2_tiehi \mem.mem_internal.code_mem[243][5]$_SDFFCE_PN0P__2629  (.L_HI(net2629));
 sg13g2_tiehi \mem.mem_internal.code_mem[243][6]$_SDFFCE_PN0P__2630  (.L_HI(net2630));
 sg13g2_tiehi \mem.mem_internal.code_mem[243][7]$_SDFFCE_PN0P__2631  (.L_HI(net2631));
 sg13g2_tiehi \mem.mem_internal.code_mem[244][0]$_SDFFCE_PN0P__2632  (.L_HI(net2632));
 sg13g2_tiehi \mem.mem_internal.code_mem[244][1]$_SDFFCE_PN0P__2633  (.L_HI(net2633));
 sg13g2_tiehi \mem.mem_internal.code_mem[244][2]$_SDFFCE_PN0P__2634  (.L_HI(net2634));
 sg13g2_tiehi \mem.mem_internal.code_mem[244][3]$_SDFFCE_PN0P__2635  (.L_HI(net2635));
 sg13g2_tiehi \mem.mem_internal.code_mem[244][4]$_SDFFCE_PN0P__2636  (.L_HI(net2636));
 sg13g2_tiehi \mem.mem_internal.code_mem[244][5]$_SDFFCE_PN0P__2637  (.L_HI(net2637));
 sg13g2_tiehi \mem.mem_internal.code_mem[244][6]$_SDFFCE_PN0P__2638  (.L_HI(net2638));
 sg13g2_tiehi \mem.mem_internal.code_mem[244][7]$_SDFFCE_PN0P__2639  (.L_HI(net2639));
 sg13g2_tiehi \mem.mem_internal.code_mem[245][0]$_SDFFCE_PN0P__2640  (.L_HI(net2640));
 sg13g2_tiehi \mem.mem_internal.code_mem[245][1]$_SDFFCE_PN0P__2641  (.L_HI(net2641));
 sg13g2_tiehi \mem.mem_internal.code_mem[245][2]$_SDFFCE_PN0P__2642  (.L_HI(net2642));
 sg13g2_tiehi \mem.mem_internal.code_mem[245][3]$_SDFFCE_PN0P__2643  (.L_HI(net2643));
 sg13g2_tiehi \mem.mem_internal.code_mem[245][4]$_SDFFCE_PN0P__2644  (.L_HI(net2644));
 sg13g2_tiehi \mem.mem_internal.code_mem[245][5]$_SDFFCE_PN0P__2645  (.L_HI(net2645));
 sg13g2_tiehi \mem.mem_internal.code_mem[245][6]$_SDFFCE_PN0P__2646  (.L_HI(net2646));
 sg13g2_tiehi \mem.mem_internal.code_mem[245][7]$_SDFFCE_PN0P__2647  (.L_HI(net2647));
 sg13g2_tiehi \mem.mem_internal.code_mem[246][0]$_SDFFCE_PN0P__2648  (.L_HI(net2648));
 sg13g2_tiehi \mem.mem_internal.code_mem[246][1]$_SDFFCE_PN0P__2649  (.L_HI(net2649));
 sg13g2_tiehi \mem.mem_internal.code_mem[246][2]$_SDFFCE_PN0P__2650  (.L_HI(net2650));
 sg13g2_tiehi \mem.mem_internal.code_mem[246][3]$_SDFFCE_PN0P__2651  (.L_HI(net2651));
 sg13g2_tiehi \mem.mem_internal.code_mem[246][4]$_SDFFCE_PN0P__2652  (.L_HI(net2652));
 sg13g2_tiehi \mem.mem_internal.code_mem[246][5]$_SDFFCE_PN0P__2653  (.L_HI(net2653));
 sg13g2_tiehi \mem.mem_internal.code_mem[246][6]$_SDFFCE_PN0P__2654  (.L_HI(net2654));
 sg13g2_tiehi \mem.mem_internal.code_mem[246][7]$_SDFFCE_PN0P__2655  (.L_HI(net2655));
 sg13g2_tiehi \mem.mem_internal.code_mem[247][0]$_SDFFCE_PN0P__2656  (.L_HI(net2656));
 sg13g2_tiehi \mem.mem_internal.code_mem[247][1]$_SDFFCE_PN0P__2657  (.L_HI(net2657));
 sg13g2_tiehi \mem.mem_internal.code_mem[247][2]$_SDFFCE_PN0P__2658  (.L_HI(net2658));
 sg13g2_tiehi \mem.mem_internal.code_mem[247][3]$_SDFFCE_PN0P__2659  (.L_HI(net2659));
 sg13g2_tiehi \mem.mem_internal.code_mem[247][4]$_SDFFCE_PN0P__2660  (.L_HI(net2660));
 sg13g2_tiehi \mem.mem_internal.code_mem[247][5]$_SDFFCE_PN0P__2661  (.L_HI(net2661));
 sg13g2_tiehi \mem.mem_internal.code_mem[247][6]$_SDFFCE_PN0P__2662  (.L_HI(net2662));
 sg13g2_tiehi \mem.mem_internal.code_mem[247][7]$_SDFFCE_PN0P__2663  (.L_HI(net2663));
 sg13g2_tiehi \mem.mem_internal.code_mem[248][0]$_SDFFCE_PN0P__2664  (.L_HI(net2664));
 sg13g2_tiehi \mem.mem_internal.code_mem[248][1]$_SDFFCE_PN0P__2665  (.L_HI(net2665));
 sg13g2_tiehi \mem.mem_internal.code_mem[248][2]$_SDFFCE_PN0P__2666  (.L_HI(net2666));
 sg13g2_tiehi \mem.mem_internal.code_mem[248][3]$_SDFFCE_PN0P__2667  (.L_HI(net2667));
 sg13g2_tiehi \mem.mem_internal.code_mem[248][4]$_SDFFCE_PN0P__2668  (.L_HI(net2668));
 sg13g2_tiehi \mem.mem_internal.code_mem[248][5]$_SDFFCE_PN0P__2669  (.L_HI(net2669));
 sg13g2_tiehi \mem.mem_internal.code_mem[248][6]$_SDFFCE_PN0P__2670  (.L_HI(net2670));
 sg13g2_tiehi \mem.mem_internal.code_mem[248][7]$_SDFFCE_PN0P__2671  (.L_HI(net2671));
 sg13g2_tiehi \mem.mem_internal.code_mem[249][0]$_SDFFCE_PN0P__2672  (.L_HI(net2672));
 sg13g2_tiehi \mem.mem_internal.code_mem[249][1]$_SDFFCE_PN0P__2673  (.L_HI(net2673));
 sg13g2_tiehi \mem.mem_internal.code_mem[249][2]$_SDFFCE_PN0P__2674  (.L_HI(net2674));
 sg13g2_tiehi \mem.mem_internal.code_mem[249][3]$_SDFFCE_PN0P__2675  (.L_HI(net2675));
 sg13g2_tiehi \mem.mem_internal.code_mem[249][4]$_SDFFCE_PN0P__2676  (.L_HI(net2676));
 sg13g2_tiehi \mem.mem_internal.code_mem[249][5]$_SDFFCE_PN0P__2677  (.L_HI(net2677));
 sg13g2_tiehi \mem.mem_internal.code_mem[249][6]$_SDFFCE_PN0P__2678  (.L_HI(net2678));
 sg13g2_tiehi \mem.mem_internal.code_mem[249][7]$_SDFFCE_PN0P__2679  (.L_HI(net2679));
 sg13g2_tiehi \mem.mem_internal.code_mem[24][0]$_SDFFCE_PN0P__2680  (.L_HI(net2680));
 sg13g2_tiehi \mem.mem_internal.code_mem[24][1]$_SDFFCE_PN0P__2681  (.L_HI(net2681));
 sg13g2_tiehi \mem.mem_internal.code_mem[24][2]$_SDFFCE_PN0P__2682  (.L_HI(net2682));
 sg13g2_tiehi \mem.mem_internal.code_mem[24][3]$_SDFFCE_PN0P__2683  (.L_HI(net2683));
 sg13g2_tiehi \mem.mem_internal.code_mem[24][4]$_SDFFCE_PN0P__2684  (.L_HI(net2684));
 sg13g2_tiehi \mem.mem_internal.code_mem[24][5]$_SDFFCE_PN0P__2685  (.L_HI(net2685));
 sg13g2_tiehi \mem.mem_internal.code_mem[24][6]$_SDFFCE_PN0P__2686  (.L_HI(net2686));
 sg13g2_tiehi \mem.mem_internal.code_mem[24][7]$_SDFFCE_PN0P__2687  (.L_HI(net2687));
 sg13g2_tiehi \mem.mem_internal.code_mem[250][0]$_SDFFCE_PN0P__2688  (.L_HI(net2688));
 sg13g2_tiehi \mem.mem_internal.code_mem[250][1]$_SDFFCE_PN0P__2689  (.L_HI(net2689));
 sg13g2_tiehi \mem.mem_internal.code_mem[250][2]$_SDFFCE_PN0P__2690  (.L_HI(net2690));
 sg13g2_tiehi \mem.mem_internal.code_mem[250][3]$_SDFFCE_PN0P__2691  (.L_HI(net2691));
 sg13g2_tiehi \mem.mem_internal.code_mem[250][4]$_SDFFCE_PN0P__2692  (.L_HI(net2692));
 sg13g2_tiehi \mem.mem_internal.code_mem[250][5]$_SDFFCE_PN0P__2693  (.L_HI(net2693));
 sg13g2_tiehi \mem.mem_internal.code_mem[250][6]$_SDFFCE_PN0P__2694  (.L_HI(net2694));
 sg13g2_tiehi \mem.mem_internal.code_mem[250][7]$_SDFFCE_PN0P__2695  (.L_HI(net2695));
 sg13g2_tiehi \mem.mem_internal.code_mem[251][0]$_SDFFCE_PN0P__2696  (.L_HI(net2696));
 sg13g2_tiehi \mem.mem_internal.code_mem[251][1]$_SDFFCE_PN0P__2697  (.L_HI(net2697));
 sg13g2_tiehi \mem.mem_internal.code_mem[251][2]$_SDFFCE_PN0P__2698  (.L_HI(net2698));
 sg13g2_tiehi \mem.mem_internal.code_mem[251][3]$_SDFFCE_PN0P__2699  (.L_HI(net2699));
 sg13g2_tiehi \mem.mem_internal.code_mem[251][4]$_SDFFCE_PN0P__2700  (.L_HI(net2700));
 sg13g2_tiehi \mem.mem_internal.code_mem[251][5]$_SDFFCE_PN0P__2701  (.L_HI(net2701));
 sg13g2_tiehi \mem.mem_internal.code_mem[251][6]$_SDFFCE_PN0P__2702  (.L_HI(net2702));
 sg13g2_tiehi \mem.mem_internal.code_mem[251][7]$_SDFFCE_PN0P__2703  (.L_HI(net2703));
 sg13g2_tiehi \mem.mem_internal.code_mem[252][0]$_SDFFCE_PN0P__2704  (.L_HI(net2704));
 sg13g2_tiehi \mem.mem_internal.code_mem[252][1]$_SDFFCE_PN0P__2705  (.L_HI(net2705));
 sg13g2_tiehi \mem.mem_internal.code_mem[252][2]$_SDFFCE_PN0P__2706  (.L_HI(net2706));
 sg13g2_tiehi \mem.mem_internal.code_mem[252][3]$_SDFFCE_PN0P__2707  (.L_HI(net2707));
 sg13g2_tiehi \mem.mem_internal.code_mem[252][4]$_SDFFCE_PN0P__2708  (.L_HI(net2708));
 sg13g2_tiehi \mem.mem_internal.code_mem[252][5]$_SDFFCE_PN0P__2709  (.L_HI(net2709));
 sg13g2_tiehi \mem.mem_internal.code_mem[252][6]$_SDFFCE_PN0P__2710  (.L_HI(net2710));
 sg13g2_tiehi \mem.mem_internal.code_mem[252][7]$_SDFFCE_PN0P__2711  (.L_HI(net2711));
 sg13g2_tiehi \mem.mem_internal.code_mem[253][0]$_SDFFCE_PN0P__2712  (.L_HI(net2712));
 sg13g2_tiehi \mem.mem_internal.code_mem[253][1]$_SDFFCE_PN0P__2713  (.L_HI(net2713));
 sg13g2_tiehi \mem.mem_internal.code_mem[253][2]$_SDFFCE_PN0P__2714  (.L_HI(net2714));
 sg13g2_tiehi \mem.mem_internal.code_mem[253][3]$_SDFFCE_PN0P__2715  (.L_HI(net2715));
 sg13g2_tiehi \mem.mem_internal.code_mem[253][4]$_SDFFCE_PN0P__2716  (.L_HI(net2716));
 sg13g2_tiehi \mem.mem_internal.code_mem[253][5]$_SDFFCE_PN0P__2717  (.L_HI(net2717));
 sg13g2_tiehi \mem.mem_internal.code_mem[253][6]$_SDFFCE_PN0P__2718  (.L_HI(net2718));
 sg13g2_tiehi \mem.mem_internal.code_mem[253][7]$_SDFFCE_PN0P__2719  (.L_HI(net2719));
 sg13g2_tiehi \mem.mem_internal.code_mem[254][0]$_SDFFCE_PN0P__2720  (.L_HI(net2720));
 sg13g2_tiehi \mem.mem_internal.code_mem[254][1]$_SDFFCE_PN0P__2721  (.L_HI(net2721));
 sg13g2_tiehi \mem.mem_internal.code_mem[254][2]$_SDFFCE_PN0P__2722  (.L_HI(net2722));
 sg13g2_tiehi \mem.mem_internal.code_mem[254][3]$_SDFFCE_PN0P__2723  (.L_HI(net2723));
 sg13g2_tiehi \mem.mem_internal.code_mem[254][4]$_SDFFCE_PN0P__2724  (.L_HI(net2724));
 sg13g2_tiehi \mem.mem_internal.code_mem[254][5]$_SDFFCE_PN0P__2725  (.L_HI(net2725));
 sg13g2_tiehi \mem.mem_internal.code_mem[254][6]$_SDFFCE_PN0P__2726  (.L_HI(net2726));
 sg13g2_tiehi \mem.mem_internal.code_mem[254][7]$_SDFFCE_PN0P__2727  (.L_HI(net2727));
 sg13g2_tiehi \mem.mem_internal.code_mem[255][0]$_SDFFCE_PN0P__2728  (.L_HI(net2728));
 sg13g2_tiehi \mem.mem_internal.code_mem[255][1]$_SDFFCE_PN0P__2729  (.L_HI(net2729));
 sg13g2_tiehi \mem.mem_internal.code_mem[255][2]$_SDFFCE_PN0P__2730  (.L_HI(net2730));
 sg13g2_tiehi \mem.mem_internal.code_mem[255][3]$_SDFFCE_PN0P__2731  (.L_HI(net2731));
 sg13g2_tiehi \mem.mem_internal.code_mem[255][4]$_SDFFCE_PN0P__2732  (.L_HI(net2732));
 sg13g2_tiehi \mem.mem_internal.code_mem[255][5]$_SDFFCE_PN0P__2733  (.L_HI(net2733));
 sg13g2_tiehi \mem.mem_internal.code_mem[255][6]$_SDFFCE_PN0P__2734  (.L_HI(net2734));
 sg13g2_tiehi \mem.mem_internal.code_mem[255][7]$_SDFFCE_PN0P__2735  (.L_HI(net2735));
 sg13g2_tiehi \mem.mem_internal.code_mem[25][0]$_SDFFCE_PN0P__2736  (.L_HI(net2736));
 sg13g2_tiehi \mem.mem_internal.code_mem[25][1]$_SDFFCE_PN0P__2737  (.L_HI(net2737));
 sg13g2_tiehi \mem.mem_internal.code_mem[25][2]$_SDFFCE_PN0P__2738  (.L_HI(net2738));
 sg13g2_tiehi \mem.mem_internal.code_mem[25][3]$_SDFFCE_PN0P__2739  (.L_HI(net2739));
 sg13g2_tiehi \mem.mem_internal.code_mem[25][4]$_SDFFCE_PN0P__2740  (.L_HI(net2740));
 sg13g2_tiehi \mem.mem_internal.code_mem[25][5]$_SDFFCE_PN0P__2741  (.L_HI(net2741));
 sg13g2_tiehi \mem.mem_internal.code_mem[25][6]$_SDFFCE_PN0P__2742  (.L_HI(net2742));
 sg13g2_tiehi \mem.mem_internal.code_mem[25][7]$_SDFFCE_PN0P__2743  (.L_HI(net2743));
 sg13g2_tiehi \mem.mem_internal.code_mem[26][0]$_SDFFCE_PN0P__2744  (.L_HI(net2744));
 sg13g2_tiehi \mem.mem_internal.code_mem[26][1]$_SDFFCE_PN0P__2745  (.L_HI(net2745));
 sg13g2_tiehi \mem.mem_internal.code_mem[26][2]$_SDFFCE_PN0P__2746  (.L_HI(net2746));
 sg13g2_tiehi \mem.mem_internal.code_mem[26][3]$_SDFFCE_PN0P__2747  (.L_HI(net2747));
 sg13g2_tiehi \mem.mem_internal.code_mem[26][4]$_SDFFCE_PN0P__2748  (.L_HI(net2748));
 sg13g2_tiehi \mem.mem_internal.code_mem[26][5]$_SDFFCE_PN0P__2749  (.L_HI(net2749));
 sg13g2_tiehi \mem.mem_internal.code_mem[26][6]$_SDFFCE_PN0P__2750  (.L_HI(net2750));
 sg13g2_tiehi \mem.mem_internal.code_mem[26][7]$_SDFFCE_PN0P__2751  (.L_HI(net2751));
 sg13g2_tiehi \mem.mem_internal.code_mem[27][0]$_SDFFCE_PN0P__2752  (.L_HI(net2752));
 sg13g2_tiehi \mem.mem_internal.code_mem[27][1]$_SDFFCE_PN0P__2753  (.L_HI(net2753));
 sg13g2_tiehi \mem.mem_internal.code_mem[27][2]$_SDFFCE_PN0P__2754  (.L_HI(net2754));
 sg13g2_tiehi \mem.mem_internal.code_mem[27][3]$_SDFFCE_PN0P__2755  (.L_HI(net2755));
 sg13g2_tiehi \mem.mem_internal.code_mem[27][4]$_SDFFCE_PN0P__2756  (.L_HI(net2756));
 sg13g2_tiehi \mem.mem_internal.code_mem[27][5]$_SDFFCE_PN0P__2757  (.L_HI(net2757));
 sg13g2_tiehi \mem.mem_internal.code_mem[27][6]$_SDFFCE_PN0P__2758  (.L_HI(net2758));
 sg13g2_tiehi \mem.mem_internal.code_mem[27][7]$_SDFFCE_PN0P__2759  (.L_HI(net2759));
 sg13g2_tiehi \mem.mem_internal.code_mem[28][0]$_SDFFCE_PN0P__2760  (.L_HI(net2760));
 sg13g2_tiehi \mem.mem_internal.code_mem[28][1]$_SDFFCE_PN0P__2761  (.L_HI(net2761));
 sg13g2_tiehi \mem.mem_internal.code_mem[28][2]$_SDFFCE_PN0P__2762  (.L_HI(net2762));
 sg13g2_tiehi \mem.mem_internal.code_mem[28][3]$_SDFFCE_PN0P__2763  (.L_HI(net2763));
 sg13g2_tiehi \mem.mem_internal.code_mem[28][4]$_SDFFCE_PN0P__2764  (.L_HI(net2764));
 sg13g2_tiehi \mem.mem_internal.code_mem[28][5]$_SDFFCE_PN0P__2765  (.L_HI(net2765));
 sg13g2_tiehi \mem.mem_internal.code_mem[28][6]$_SDFFCE_PN0P__2766  (.L_HI(net2766));
 sg13g2_tiehi \mem.mem_internal.code_mem[28][7]$_SDFFCE_PN0P__2767  (.L_HI(net2767));
 sg13g2_tiehi \mem.mem_internal.code_mem[29][0]$_SDFFCE_PN0P__2768  (.L_HI(net2768));
 sg13g2_tiehi \mem.mem_internal.code_mem[29][1]$_SDFFCE_PN0P__2769  (.L_HI(net2769));
 sg13g2_tiehi \mem.mem_internal.code_mem[29][2]$_SDFFCE_PN0P__2770  (.L_HI(net2770));
 sg13g2_tiehi \mem.mem_internal.code_mem[29][3]$_SDFFCE_PN0P__2771  (.L_HI(net2771));
 sg13g2_tiehi \mem.mem_internal.code_mem[29][4]$_SDFFCE_PN0P__2772  (.L_HI(net2772));
 sg13g2_tiehi \mem.mem_internal.code_mem[29][5]$_SDFFCE_PN0P__2773  (.L_HI(net2773));
 sg13g2_tiehi \mem.mem_internal.code_mem[29][6]$_SDFFCE_PN0P__2774  (.L_HI(net2774));
 sg13g2_tiehi \mem.mem_internal.code_mem[29][7]$_SDFFCE_PN0P__2775  (.L_HI(net2775));
 sg13g2_tiehi \mem.mem_internal.code_mem[2][0]$_SDFFCE_PN0P__2776  (.L_HI(net2776));
 sg13g2_tiehi \mem.mem_internal.code_mem[2][1]$_SDFFCE_PN0P__2777  (.L_HI(net2777));
 sg13g2_tiehi \mem.mem_internal.code_mem[2][2]$_SDFFCE_PN0P__2778  (.L_HI(net2778));
 sg13g2_tiehi \mem.mem_internal.code_mem[2][3]$_SDFFCE_PN0P__2779  (.L_HI(net2779));
 sg13g2_tiehi \mem.mem_internal.code_mem[2][4]$_SDFFCE_PN0P__2780  (.L_HI(net2780));
 sg13g2_tiehi \mem.mem_internal.code_mem[2][5]$_SDFFCE_PN0P__2781  (.L_HI(net2781));
 sg13g2_tiehi \mem.mem_internal.code_mem[2][6]$_SDFFCE_PN0P__2782  (.L_HI(net2782));
 sg13g2_tiehi \mem.mem_internal.code_mem[2][7]$_SDFFCE_PN0P__2783  (.L_HI(net2783));
 sg13g2_tiehi \mem.mem_internal.code_mem[30][0]$_SDFFCE_PN0P__2784  (.L_HI(net2784));
 sg13g2_tiehi \mem.mem_internal.code_mem[30][1]$_SDFFCE_PN0P__2785  (.L_HI(net2785));
 sg13g2_tiehi \mem.mem_internal.code_mem[30][2]$_SDFFCE_PN0P__2786  (.L_HI(net2786));
 sg13g2_tiehi \mem.mem_internal.code_mem[30][3]$_SDFFCE_PN0P__2787  (.L_HI(net2787));
 sg13g2_tiehi \mem.mem_internal.code_mem[30][4]$_SDFFCE_PN0P__2788  (.L_HI(net2788));
 sg13g2_tiehi \mem.mem_internal.code_mem[30][5]$_SDFFCE_PN0P__2789  (.L_HI(net2789));
 sg13g2_tiehi \mem.mem_internal.code_mem[30][6]$_SDFFCE_PN0P__2790  (.L_HI(net2790));
 sg13g2_tiehi \mem.mem_internal.code_mem[30][7]$_SDFFCE_PN0P__2791  (.L_HI(net2791));
 sg13g2_tiehi \mem.mem_internal.code_mem[31][0]$_SDFFCE_PN0P__2792  (.L_HI(net2792));
 sg13g2_tiehi \mem.mem_internal.code_mem[31][1]$_SDFFCE_PN0P__2793  (.L_HI(net2793));
 sg13g2_tiehi \mem.mem_internal.code_mem[31][2]$_SDFFCE_PN0P__2794  (.L_HI(net2794));
 sg13g2_tiehi \mem.mem_internal.code_mem[31][3]$_SDFFCE_PN0P__2795  (.L_HI(net2795));
 sg13g2_tiehi \mem.mem_internal.code_mem[31][4]$_SDFFCE_PN0P__2796  (.L_HI(net2796));
 sg13g2_tiehi \mem.mem_internal.code_mem[31][5]$_SDFFCE_PN0P__2797  (.L_HI(net2797));
 sg13g2_tiehi \mem.mem_internal.code_mem[31][6]$_SDFFCE_PN0P__2798  (.L_HI(net2798));
 sg13g2_tiehi \mem.mem_internal.code_mem[31][7]$_SDFFCE_PN0P__2799  (.L_HI(net2799));
 sg13g2_tiehi \mem.mem_internal.code_mem[32][0]$_SDFFCE_PN0P__2800  (.L_HI(net2800));
 sg13g2_tiehi \mem.mem_internal.code_mem[32][1]$_SDFFCE_PN0P__2801  (.L_HI(net2801));
 sg13g2_tiehi \mem.mem_internal.code_mem[32][2]$_SDFFCE_PN0P__2802  (.L_HI(net2802));
 sg13g2_tiehi \mem.mem_internal.code_mem[32][3]$_SDFFCE_PN0P__2803  (.L_HI(net2803));
 sg13g2_tiehi \mem.mem_internal.code_mem[32][4]$_SDFFCE_PN0P__2804  (.L_HI(net2804));
 sg13g2_tiehi \mem.mem_internal.code_mem[32][5]$_SDFFCE_PN0P__2805  (.L_HI(net2805));
 sg13g2_tiehi \mem.mem_internal.code_mem[32][6]$_SDFFCE_PN0P__2806  (.L_HI(net2806));
 sg13g2_tiehi \mem.mem_internal.code_mem[32][7]$_SDFFCE_PN0P__2807  (.L_HI(net2807));
 sg13g2_tiehi \mem.mem_internal.code_mem[33][0]$_SDFFCE_PN0P__2808  (.L_HI(net2808));
 sg13g2_tiehi \mem.mem_internal.code_mem[33][1]$_SDFFCE_PN0P__2809  (.L_HI(net2809));
 sg13g2_tiehi \mem.mem_internal.code_mem[33][2]$_SDFFCE_PN0P__2810  (.L_HI(net2810));
 sg13g2_tiehi \mem.mem_internal.code_mem[33][3]$_SDFFCE_PN0P__2811  (.L_HI(net2811));
 sg13g2_tiehi \mem.mem_internal.code_mem[33][4]$_SDFFCE_PN0P__2812  (.L_HI(net2812));
 sg13g2_tiehi \mem.mem_internal.code_mem[33][5]$_SDFFCE_PN0P__2813  (.L_HI(net2813));
 sg13g2_tiehi \mem.mem_internal.code_mem[33][6]$_SDFFCE_PN0P__2814  (.L_HI(net2814));
 sg13g2_tiehi \mem.mem_internal.code_mem[33][7]$_SDFFCE_PN0P__2815  (.L_HI(net2815));
 sg13g2_tiehi \mem.mem_internal.code_mem[34][0]$_SDFFCE_PN0P__2816  (.L_HI(net2816));
 sg13g2_tiehi \mem.mem_internal.code_mem[34][1]$_SDFFCE_PN0P__2817  (.L_HI(net2817));
 sg13g2_tiehi \mem.mem_internal.code_mem[34][2]$_SDFFCE_PN0P__2818  (.L_HI(net2818));
 sg13g2_tiehi \mem.mem_internal.code_mem[34][3]$_SDFFCE_PN0P__2819  (.L_HI(net2819));
 sg13g2_tiehi \mem.mem_internal.code_mem[34][4]$_SDFFCE_PN0P__2820  (.L_HI(net2820));
 sg13g2_tiehi \mem.mem_internal.code_mem[34][5]$_SDFFCE_PN0P__2821  (.L_HI(net2821));
 sg13g2_tiehi \mem.mem_internal.code_mem[34][6]$_SDFFCE_PN0P__2822  (.L_HI(net2822));
 sg13g2_tiehi \mem.mem_internal.code_mem[34][7]$_SDFFCE_PN0P__2823  (.L_HI(net2823));
 sg13g2_tiehi \mem.mem_internal.code_mem[35][0]$_SDFFCE_PN0P__2824  (.L_HI(net2824));
 sg13g2_tiehi \mem.mem_internal.code_mem[35][1]$_SDFFCE_PN0P__2825  (.L_HI(net2825));
 sg13g2_tiehi \mem.mem_internal.code_mem[35][2]$_SDFFCE_PN0P__2826  (.L_HI(net2826));
 sg13g2_tiehi \mem.mem_internal.code_mem[35][3]$_SDFFCE_PN0P__2827  (.L_HI(net2827));
 sg13g2_tiehi \mem.mem_internal.code_mem[35][4]$_SDFFCE_PN0P__2828  (.L_HI(net2828));
 sg13g2_tiehi \mem.mem_internal.code_mem[35][5]$_SDFFCE_PN0P__2829  (.L_HI(net2829));
 sg13g2_tiehi \mem.mem_internal.code_mem[35][6]$_SDFFCE_PN0P__2830  (.L_HI(net2830));
 sg13g2_tiehi \mem.mem_internal.code_mem[35][7]$_SDFFCE_PN0P__2831  (.L_HI(net2831));
 sg13g2_tiehi \mem.mem_internal.code_mem[36][0]$_SDFFCE_PN0P__2832  (.L_HI(net2832));
 sg13g2_tiehi \mem.mem_internal.code_mem[36][1]$_SDFFCE_PN0P__2833  (.L_HI(net2833));
 sg13g2_tiehi \mem.mem_internal.code_mem[36][2]$_SDFFCE_PN0P__2834  (.L_HI(net2834));
 sg13g2_tiehi \mem.mem_internal.code_mem[36][3]$_SDFFCE_PN0P__2835  (.L_HI(net2835));
 sg13g2_tiehi \mem.mem_internal.code_mem[36][4]$_SDFFCE_PN0P__2836  (.L_HI(net2836));
 sg13g2_tiehi \mem.mem_internal.code_mem[36][5]$_SDFFCE_PN0P__2837  (.L_HI(net2837));
 sg13g2_tiehi \mem.mem_internal.code_mem[36][6]$_SDFFCE_PN0P__2838  (.L_HI(net2838));
 sg13g2_tiehi \mem.mem_internal.code_mem[36][7]$_SDFFCE_PN0P__2839  (.L_HI(net2839));
 sg13g2_tiehi \mem.mem_internal.code_mem[37][0]$_SDFFCE_PN0P__2840  (.L_HI(net2840));
 sg13g2_tiehi \mem.mem_internal.code_mem[37][1]$_SDFFCE_PN0P__2841  (.L_HI(net2841));
 sg13g2_tiehi \mem.mem_internal.code_mem[37][2]$_SDFFCE_PN0P__2842  (.L_HI(net2842));
 sg13g2_tiehi \mem.mem_internal.code_mem[37][3]$_SDFFCE_PN0P__2843  (.L_HI(net2843));
 sg13g2_tiehi \mem.mem_internal.code_mem[37][4]$_SDFFCE_PN0P__2844  (.L_HI(net2844));
 sg13g2_tiehi \mem.mem_internal.code_mem[37][5]$_SDFFCE_PN0P__2845  (.L_HI(net2845));
 sg13g2_tiehi \mem.mem_internal.code_mem[37][6]$_SDFFCE_PN0P__2846  (.L_HI(net2846));
 sg13g2_tiehi \mem.mem_internal.code_mem[37][7]$_SDFFCE_PN0P__2847  (.L_HI(net2847));
 sg13g2_tiehi \mem.mem_internal.code_mem[38][0]$_SDFFCE_PN0P__2848  (.L_HI(net2848));
 sg13g2_tiehi \mem.mem_internal.code_mem[38][1]$_SDFFCE_PN0P__2849  (.L_HI(net2849));
 sg13g2_tiehi \mem.mem_internal.code_mem[38][2]$_SDFFCE_PN0P__2850  (.L_HI(net2850));
 sg13g2_tiehi \mem.mem_internal.code_mem[38][3]$_SDFFCE_PN0P__2851  (.L_HI(net2851));
 sg13g2_tiehi \mem.mem_internal.code_mem[38][4]$_SDFFCE_PN0P__2852  (.L_HI(net2852));
 sg13g2_tiehi \mem.mem_internal.code_mem[38][5]$_SDFFCE_PN0P__2853  (.L_HI(net2853));
 sg13g2_tiehi \mem.mem_internal.code_mem[38][6]$_SDFFCE_PN0P__2854  (.L_HI(net2854));
 sg13g2_tiehi \mem.mem_internal.code_mem[38][7]$_SDFFCE_PN0P__2855  (.L_HI(net2855));
 sg13g2_tiehi \mem.mem_internal.code_mem[39][0]$_SDFFCE_PN0P__2856  (.L_HI(net2856));
 sg13g2_tiehi \mem.mem_internal.code_mem[39][1]$_SDFFCE_PN0P__2857  (.L_HI(net2857));
 sg13g2_tiehi \mem.mem_internal.code_mem[39][2]$_SDFFCE_PN0P__2858  (.L_HI(net2858));
 sg13g2_tiehi \mem.mem_internal.code_mem[39][3]$_SDFFCE_PN0P__2859  (.L_HI(net2859));
 sg13g2_tiehi \mem.mem_internal.code_mem[39][4]$_SDFFCE_PN0P__2860  (.L_HI(net2860));
 sg13g2_tiehi \mem.mem_internal.code_mem[39][5]$_SDFFCE_PN0P__2861  (.L_HI(net2861));
 sg13g2_tiehi \mem.mem_internal.code_mem[39][6]$_SDFFCE_PN0P__2862  (.L_HI(net2862));
 sg13g2_tiehi \mem.mem_internal.code_mem[39][7]$_SDFFCE_PN0P__2863  (.L_HI(net2863));
 sg13g2_tiehi \mem.mem_internal.code_mem[3][0]$_SDFFCE_PN0P__2864  (.L_HI(net2864));
 sg13g2_tiehi \mem.mem_internal.code_mem[3][1]$_SDFFCE_PN0P__2865  (.L_HI(net2865));
 sg13g2_tiehi \mem.mem_internal.code_mem[3][2]$_SDFFCE_PN0P__2866  (.L_HI(net2866));
 sg13g2_tiehi \mem.mem_internal.code_mem[3][3]$_SDFFCE_PN0P__2867  (.L_HI(net2867));
 sg13g2_tiehi \mem.mem_internal.code_mem[3][4]$_SDFFCE_PN0P__2868  (.L_HI(net2868));
 sg13g2_tiehi \mem.mem_internal.code_mem[3][5]$_SDFFCE_PN0P__2869  (.L_HI(net2869));
 sg13g2_tiehi \mem.mem_internal.code_mem[3][6]$_SDFFCE_PN0P__2870  (.L_HI(net2870));
 sg13g2_tiehi \mem.mem_internal.code_mem[3][7]$_SDFFCE_PN0P__2871  (.L_HI(net2871));
 sg13g2_tiehi \mem.mem_internal.code_mem[40][0]$_SDFFCE_PN0P__2872  (.L_HI(net2872));
 sg13g2_tiehi \mem.mem_internal.code_mem[40][1]$_SDFFCE_PN0P__2873  (.L_HI(net2873));
 sg13g2_tiehi \mem.mem_internal.code_mem[40][2]$_SDFFCE_PN0P__2874  (.L_HI(net2874));
 sg13g2_tiehi \mem.mem_internal.code_mem[40][3]$_SDFFCE_PN0P__2875  (.L_HI(net2875));
 sg13g2_tiehi \mem.mem_internal.code_mem[40][4]$_SDFFCE_PN0P__2876  (.L_HI(net2876));
 sg13g2_tiehi \mem.mem_internal.code_mem[40][5]$_SDFFCE_PN0P__2877  (.L_HI(net2877));
 sg13g2_tiehi \mem.mem_internal.code_mem[40][6]$_SDFFCE_PN0P__2878  (.L_HI(net2878));
 sg13g2_tiehi \mem.mem_internal.code_mem[40][7]$_SDFFCE_PN0P__2879  (.L_HI(net2879));
 sg13g2_tiehi \mem.mem_internal.code_mem[41][0]$_SDFFCE_PN0P__2880  (.L_HI(net2880));
 sg13g2_tiehi \mem.mem_internal.code_mem[41][1]$_SDFFCE_PN0P__2881  (.L_HI(net2881));
 sg13g2_tiehi \mem.mem_internal.code_mem[41][2]$_SDFFCE_PN0P__2882  (.L_HI(net2882));
 sg13g2_tiehi \mem.mem_internal.code_mem[41][3]$_SDFFCE_PN0P__2883  (.L_HI(net2883));
 sg13g2_tiehi \mem.mem_internal.code_mem[41][4]$_SDFFCE_PN0P__2884  (.L_HI(net2884));
 sg13g2_tiehi \mem.mem_internal.code_mem[41][5]$_SDFFCE_PN0P__2885  (.L_HI(net2885));
 sg13g2_tiehi \mem.mem_internal.code_mem[41][6]$_SDFFCE_PN0P__2886  (.L_HI(net2886));
 sg13g2_tiehi \mem.mem_internal.code_mem[41][7]$_SDFFCE_PN0P__2887  (.L_HI(net2887));
 sg13g2_tiehi \mem.mem_internal.code_mem[42][0]$_SDFFCE_PN0P__2888  (.L_HI(net2888));
 sg13g2_tiehi \mem.mem_internal.code_mem[42][1]$_SDFFCE_PN0P__2889  (.L_HI(net2889));
 sg13g2_tiehi \mem.mem_internal.code_mem[42][2]$_SDFFCE_PN0P__2890  (.L_HI(net2890));
 sg13g2_tiehi \mem.mem_internal.code_mem[42][3]$_SDFFCE_PN0P__2891  (.L_HI(net2891));
 sg13g2_tiehi \mem.mem_internal.code_mem[42][4]$_SDFFCE_PN0P__2892  (.L_HI(net2892));
 sg13g2_tiehi \mem.mem_internal.code_mem[42][5]$_SDFFCE_PN0P__2893  (.L_HI(net2893));
 sg13g2_tiehi \mem.mem_internal.code_mem[42][6]$_SDFFCE_PN0P__2894  (.L_HI(net2894));
 sg13g2_tiehi \mem.mem_internal.code_mem[42][7]$_SDFFCE_PN0P__2895  (.L_HI(net2895));
 sg13g2_tiehi \mem.mem_internal.code_mem[43][0]$_SDFFCE_PN0P__2896  (.L_HI(net2896));
 sg13g2_tiehi \mem.mem_internal.code_mem[43][1]$_SDFFCE_PN0P__2897  (.L_HI(net2897));
 sg13g2_tiehi \mem.mem_internal.code_mem[43][2]$_SDFFCE_PN0P__2898  (.L_HI(net2898));
 sg13g2_tiehi \mem.mem_internal.code_mem[43][3]$_SDFFCE_PN0P__2899  (.L_HI(net2899));
 sg13g2_tiehi \mem.mem_internal.code_mem[43][4]$_SDFFCE_PN0P__2900  (.L_HI(net2900));
 sg13g2_tiehi \mem.mem_internal.code_mem[43][5]$_SDFFCE_PN0P__2901  (.L_HI(net2901));
 sg13g2_tiehi \mem.mem_internal.code_mem[43][6]$_SDFFCE_PN0P__2902  (.L_HI(net2902));
 sg13g2_tiehi \mem.mem_internal.code_mem[43][7]$_SDFFCE_PN0P__2903  (.L_HI(net2903));
 sg13g2_tiehi \mem.mem_internal.code_mem[44][0]$_SDFFCE_PN0P__2904  (.L_HI(net2904));
 sg13g2_tiehi \mem.mem_internal.code_mem[44][1]$_SDFFCE_PN0P__2905  (.L_HI(net2905));
 sg13g2_tiehi \mem.mem_internal.code_mem[44][2]$_SDFFCE_PN0P__2906  (.L_HI(net2906));
 sg13g2_tiehi \mem.mem_internal.code_mem[44][3]$_SDFFCE_PN0P__2907  (.L_HI(net2907));
 sg13g2_tiehi \mem.mem_internal.code_mem[44][4]$_SDFFCE_PN0P__2908  (.L_HI(net2908));
 sg13g2_tiehi \mem.mem_internal.code_mem[44][5]$_SDFFCE_PN0P__2909  (.L_HI(net2909));
 sg13g2_tiehi \mem.mem_internal.code_mem[44][6]$_SDFFCE_PN0P__2910  (.L_HI(net2910));
 sg13g2_tiehi \mem.mem_internal.code_mem[44][7]$_SDFFCE_PN0P__2911  (.L_HI(net2911));
 sg13g2_tiehi \mem.mem_internal.code_mem[45][0]$_SDFFCE_PN0P__2912  (.L_HI(net2912));
 sg13g2_tiehi \mem.mem_internal.code_mem[45][1]$_SDFFCE_PN0P__2913  (.L_HI(net2913));
 sg13g2_tiehi \mem.mem_internal.code_mem[45][2]$_SDFFCE_PN0P__2914  (.L_HI(net2914));
 sg13g2_tiehi \mem.mem_internal.code_mem[45][3]$_SDFFCE_PN0P__2915  (.L_HI(net2915));
 sg13g2_tiehi \mem.mem_internal.code_mem[45][4]$_SDFFCE_PN0P__2916  (.L_HI(net2916));
 sg13g2_tiehi \mem.mem_internal.code_mem[45][5]$_SDFFCE_PN0P__2917  (.L_HI(net2917));
 sg13g2_tiehi \mem.mem_internal.code_mem[45][6]$_SDFFCE_PN0P__2918  (.L_HI(net2918));
 sg13g2_tiehi \mem.mem_internal.code_mem[45][7]$_SDFFCE_PN0P__2919  (.L_HI(net2919));
 sg13g2_tiehi \mem.mem_internal.code_mem[46][0]$_SDFFCE_PN0P__2920  (.L_HI(net2920));
 sg13g2_tiehi \mem.mem_internal.code_mem[46][1]$_SDFFCE_PN0P__2921  (.L_HI(net2921));
 sg13g2_tiehi \mem.mem_internal.code_mem[46][2]$_SDFFCE_PN0P__2922  (.L_HI(net2922));
 sg13g2_tiehi \mem.mem_internal.code_mem[46][3]$_SDFFCE_PN0P__2923  (.L_HI(net2923));
 sg13g2_tiehi \mem.mem_internal.code_mem[46][4]$_SDFFCE_PN0P__2924  (.L_HI(net2924));
 sg13g2_tiehi \mem.mem_internal.code_mem[46][5]$_SDFFCE_PN0P__2925  (.L_HI(net2925));
 sg13g2_tiehi \mem.mem_internal.code_mem[46][6]$_SDFFCE_PN0P__2926  (.L_HI(net2926));
 sg13g2_tiehi \mem.mem_internal.code_mem[46][7]$_SDFFCE_PN0P__2927  (.L_HI(net2927));
 sg13g2_tiehi \mem.mem_internal.code_mem[47][0]$_SDFFCE_PN0P__2928  (.L_HI(net2928));
 sg13g2_tiehi \mem.mem_internal.code_mem[47][1]$_SDFFCE_PN0P__2929  (.L_HI(net2929));
 sg13g2_tiehi \mem.mem_internal.code_mem[47][2]$_SDFFCE_PN0P__2930  (.L_HI(net2930));
 sg13g2_tiehi \mem.mem_internal.code_mem[47][3]$_SDFFCE_PN0P__2931  (.L_HI(net2931));
 sg13g2_tiehi \mem.mem_internal.code_mem[47][4]$_SDFFCE_PN0P__2932  (.L_HI(net2932));
 sg13g2_tiehi \mem.mem_internal.code_mem[47][5]$_SDFFCE_PN0P__2933  (.L_HI(net2933));
 sg13g2_tiehi \mem.mem_internal.code_mem[47][6]$_SDFFCE_PN0P__2934  (.L_HI(net2934));
 sg13g2_tiehi \mem.mem_internal.code_mem[47][7]$_SDFFCE_PN0P__2935  (.L_HI(net2935));
 sg13g2_tiehi \mem.mem_internal.code_mem[48][0]$_SDFFCE_PN0P__2936  (.L_HI(net2936));
 sg13g2_tiehi \mem.mem_internal.code_mem[48][1]$_SDFFCE_PN0P__2937  (.L_HI(net2937));
 sg13g2_tiehi \mem.mem_internal.code_mem[48][2]$_SDFFCE_PN0P__2938  (.L_HI(net2938));
 sg13g2_tiehi \mem.mem_internal.code_mem[48][3]$_SDFFCE_PN0P__2939  (.L_HI(net2939));
 sg13g2_tiehi \mem.mem_internal.code_mem[48][4]$_SDFFCE_PN0P__2940  (.L_HI(net2940));
 sg13g2_tiehi \mem.mem_internal.code_mem[48][5]$_SDFFCE_PN0P__2941  (.L_HI(net2941));
 sg13g2_tiehi \mem.mem_internal.code_mem[48][6]$_SDFFCE_PN0P__2942  (.L_HI(net2942));
 sg13g2_tiehi \mem.mem_internal.code_mem[48][7]$_SDFFCE_PN0P__2943  (.L_HI(net2943));
 sg13g2_tiehi \mem.mem_internal.code_mem[49][0]$_SDFFCE_PN0P__2944  (.L_HI(net2944));
 sg13g2_tiehi \mem.mem_internal.code_mem[49][1]$_SDFFCE_PN0P__2945  (.L_HI(net2945));
 sg13g2_tiehi \mem.mem_internal.code_mem[49][2]$_SDFFCE_PN0P__2946  (.L_HI(net2946));
 sg13g2_tiehi \mem.mem_internal.code_mem[49][3]$_SDFFCE_PN0P__2947  (.L_HI(net2947));
 sg13g2_tiehi \mem.mem_internal.code_mem[49][4]$_SDFFCE_PN0P__2948  (.L_HI(net2948));
 sg13g2_tiehi \mem.mem_internal.code_mem[49][5]$_SDFFCE_PN0P__2949  (.L_HI(net2949));
 sg13g2_tiehi \mem.mem_internal.code_mem[49][6]$_SDFFCE_PN0P__2950  (.L_HI(net2950));
 sg13g2_tiehi \mem.mem_internal.code_mem[49][7]$_SDFFCE_PN0P__2951  (.L_HI(net2951));
 sg13g2_tiehi \mem.mem_internal.code_mem[4][0]$_SDFFCE_PN0P__2952  (.L_HI(net2952));
 sg13g2_tiehi \mem.mem_internal.code_mem[4][1]$_SDFFCE_PN0P__2953  (.L_HI(net2953));
 sg13g2_tiehi \mem.mem_internal.code_mem[4][2]$_SDFFCE_PN0P__2954  (.L_HI(net2954));
 sg13g2_tiehi \mem.mem_internal.code_mem[4][3]$_SDFFCE_PN0P__2955  (.L_HI(net2955));
 sg13g2_tiehi \mem.mem_internal.code_mem[4][4]$_SDFFCE_PN0P__2956  (.L_HI(net2956));
 sg13g2_tiehi \mem.mem_internal.code_mem[4][5]$_SDFFCE_PN0P__2957  (.L_HI(net2957));
 sg13g2_tiehi \mem.mem_internal.code_mem[4][6]$_SDFFCE_PN0P__2958  (.L_HI(net2958));
 sg13g2_tiehi \mem.mem_internal.code_mem[4][7]$_SDFFCE_PN0P__2959  (.L_HI(net2959));
 sg13g2_tiehi \mem.mem_internal.code_mem[50][0]$_SDFFCE_PN0P__2960  (.L_HI(net2960));
 sg13g2_tiehi \mem.mem_internal.code_mem[50][1]$_SDFFCE_PN0P__2961  (.L_HI(net2961));
 sg13g2_tiehi \mem.mem_internal.code_mem[50][2]$_SDFFCE_PN0P__2962  (.L_HI(net2962));
 sg13g2_tiehi \mem.mem_internal.code_mem[50][3]$_SDFFCE_PN0P__2963  (.L_HI(net2963));
 sg13g2_tiehi \mem.mem_internal.code_mem[50][4]$_SDFFCE_PN0P__2964  (.L_HI(net2964));
 sg13g2_tiehi \mem.mem_internal.code_mem[50][5]$_SDFFCE_PN0P__2965  (.L_HI(net2965));
 sg13g2_tiehi \mem.mem_internal.code_mem[50][6]$_SDFFCE_PN0P__2966  (.L_HI(net2966));
 sg13g2_tiehi \mem.mem_internal.code_mem[50][7]$_SDFFCE_PN0P__2967  (.L_HI(net2967));
 sg13g2_tiehi \mem.mem_internal.code_mem[51][0]$_SDFFCE_PN0P__2968  (.L_HI(net2968));
 sg13g2_tiehi \mem.mem_internal.code_mem[51][1]$_SDFFCE_PN0P__2969  (.L_HI(net2969));
 sg13g2_tiehi \mem.mem_internal.code_mem[51][2]$_SDFFCE_PN0P__2970  (.L_HI(net2970));
 sg13g2_tiehi \mem.mem_internal.code_mem[51][3]$_SDFFCE_PN0P__2971  (.L_HI(net2971));
 sg13g2_tiehi \mem.mem_internal.code_mem[51][4]$_SDFFCE_PN0P__2972  (.L_HI(net2972));
 sg13g2_tiehi \mem.mem_internal.code_mem[51][5]$_SDFFCE_PN0P__2973  (.L_HI(net2973));
 sg13g2_tiehi \mem.mem_internal.code_mem[51][6]$_SDFFCE_PN0P__2974  (.L_HI(net2974));
 sg13g2_tiehi \mem.mem_internal.code_mem[51][7]$_SDFFCE_PN0P__2975  (.L_HI(net2975));
 sg13g2_tiehi \mem.mem_internal.code_mem[52][0]$_SDFFCE_PN0P__2976  (.L_HI(net2976));
 sg13g2_tiehi \mem.mem_internal.code_mem[52][1]$_SDFFCE_PN0P__2977  (.L_HI(net2977));
 sg13g2_tiehi \mem.mem_internal.code_mem[52][2]$_SDFFCE_PN0P__2978  (.L_HI(net2978));
 sg13g2_tiehi \mem.mem_internal.code_mem[52][3]$_SDFFCE_PN0P__2979  (.L_HI(net2979));
 sg13g2_tiehi \mem.mem_internal.code_mem[52][4]$_SDFFCE_PN0P__2980  (.L_HI(net2980));
 sg13g2_tiehi \mem.mem_internal.code_mem[52][5]$_SDFFCE_PN0P__2981  (.L_HI(net2981));
 sg13g2_tiehi \mem.mem_internal.code_mem[52][6]$_SDFFCE_PN0P__2982  (.L_HI(net2982));
 sg13g2_tiehi \mem.mem_internal.code_mem[52][7]$_SDFFCE_PN0P__2983  (.L_HI(net2983));
 sg13g2_tiehi \mem.mem_internal.code_mem[53][0]$_SDFFCE_PN0P__2984  (.L_HI(net2984));
 sg13g2_tiehi \mem.mem_internal.code_mem[53][1]$_SDFFCE_PN0P__2985  (.L_HI(net2985));
 sg13g2_tiehi \mem.mem_internal.code_mem[53][2]$_SDFFCE_PN0P__2986  (.L_HI(net2986));
 sg13g2_tiehi \mem.mem_internal.code_mem[53][3]$_SDFFCE_PN0P__2987  (.L_HI(net2987));
 sg13g2_tiehi \mem.mem_internal.code_mem[53][4]$_SDFFCE_PN0P__2988  (.L_HI(net2988));
 sg13g2_tiehi \mem.mem_internal.code_mem[53][5]$_SDFFCE_PN0P__2989  (.L_HI(net2989));
 sg13g2_tiehi \mem.mem_internal.code_mem[53][6]$_SDFFCE_PN0P__2990  (.L_HI(net2990));
 sg13g2_tiehi \mem.mem_internal.code_mem[53][7]$_SDFFCE_PN0P__2991  (.L_HI(net2991));
 sg13g2_tiehi \mem.mem_internal.code_mem[54][0]$_SDFFCE_PN0P__2992  (.L_HI(net2992));
 sg13g2_tiehi \mem.mem_internal.code_mem[54][1]$_SDFFCE_PN0P__2993  (.L_HI(net2993));
 sg13g2_tiehi \mem.mem_internal.code_mem[54][2]$_SDFFCE_PN0P__2994  (.L_HI(net2994));
 sg13g2_tiehi \mem.mem_internal.code_mem[54][3]$_SDFFCE_PN0P__2995  (.L_HI(net2995));
 sg13g2_tiehi \mem.mem_internal.code_mem[54][4]$_SDFFCE_PN0P__2996  (.L_HI(net2996));
 sg13g2_tiehi \mem.mem_internal.code_mem[54][5]$_SDFFCE_PN0P__2997  (.L_HI(net2997));
 sg13g2_tiehi \mem.mem_internal.code_mem[54][6]$_SDFFCE_PN0P__2998  (.L_HI(net2998));
 sg13g2_tiehi \mem.mem_internal.code_mem[54][7]$_SDFFCE_PN0P__2999  (.L_HI(net2999));
 sg13g2_tiehi \mem.mem_internal.code_mem[55][0]$_SDFFCE_PN0P__3000  (.L_HI(net3000));
 sg13g2_tiehi \mem.mem_internal.code_mem[55][1]$_SDFFCE_PN0P__3001  (.L_HI(net3001));
 sg13g2_tiehi \mem.mem_internal.code_mem[55][2]$_SDFFCE_PN0P__3002  (.L_HI(net3002));
 sg13g2_tiehi \mem.mem_internal.code_mem[55][3]$_SDFFCE_PN0P__3003  (.L_HI(net3003));
 sg13g2_tiehi \mem.mem_internal.code_mem[55][4]$_SDFFCE_PN0P__3004  (.L_HI(net3004));
 sg13g2_tiehi \mem.mem_internal.code_mem[55][5]$_SDFFCE_PN0P__3005  (.L_HI(net3005));
 sg13g2_tiehi \mem.mem_internal.code_mem[55][6]$_SDFFCE_PN0P__3006  (.L_HI(net3006));
 sg13g2_tiehi \mem.mem_internal.code_mem[55][7]$_SDFFCE_PN0P__3007  (.L_HI(net3007));
 sg13g2_tiehi \mem.mem_internal.code_mem[56][0]$_SDFFCE_PN0P__3008  (.L_HI(net3008));
 sg13g2_tiehi \mem.mem_internal.code_mem[56][1]$_SDFFCE_PN0P__3009  (.L_HI(net3009));
 sg13g2_tiehi \mem.mem_internal.code_mem[56][2]$_SDFFCE_PN0P__3010  (.L_HI(net3010));
 sg13g2_tiehi \mem.mem_internal.code_mem[56][3]$_SDFFCE_PN0P__3011  (.L_HI(net3011));
 sg13g2_tiehi \mem.mem_internal.code_mem[56][4]$_SDFFCE_PN0P__3012  (.L_HI(net3012));
 sg13g2_tiehi \mem.mem_internal.code_mem[56][5]$_SDFFCE_PN0P__3013  (.L_HI(net3013));
 sg13g2_tiehi \mem.mem_internal.code_mem[56][6]$_SDFFCE_PN0P__3014  (.L_HI(net3014));
 sg13g2_tiehi \mem.mem_internal.code_mem[56][7]$_SDFFCE_PN0P__3015  (.L_HI(net3015));
 sg13g2_tiehi \mem.mem_internal.code_mem[57][0]$_SDFFCE_PN0P__3016  (.L_HI(net3016));
 sg13g2_tiehi \mem.mem_internal.code_mem[57][1]$_SDFFCE_PN0P__3017  (.L_HI(net3017));
 sg13g2_tiehi \mem.mem_internal.code_mem[57][2]$_SDFFCE_PN0P__3018  (.L_HI(net3018));
 sg13g2_tiehi \mem.mem_internal.code_mem[57][3]$_SDFFCE_PN0P__3019  (.L_HI(net3019));
 sg13g2_tiehi \mem.mem_internal.code_mem[57][4]$_SDFFCE_PN0P__3020  (.L_HI(net3020));
 sg13g2_tiehi \mem.mem_internal.code_mem[57][5]$_SDFFCE_PN0P__3021  (.L_HI(net3021));
 sg13g2_tiehi \mem.mem_internal.code_mem[57][6]$_SDFFCE_PN0P__3022  (.L_HI(net3022));
 sg13g2_tiehi \mem.mem_internal.code_mem[57][7]$_SDFFCE_PN0P__3023  (.L_HI(net3023));
 sg13g2_tiehi \mem.mem_internal.code_mem[58][0]$_SDFFCE_PN0P__3024  (.L_HI(net3024));
 sg13g2_tiehi \mem.mem_internal.code_mem[58][1]$_SDFFCE_PN0P__3025  (.L_HI(net3025));
 sg13g2_tiehi \mem.mem_internal.code_mem[58][2]$_SDFFCE_PN0P__3026  (.L_HI(net3026));
 sg13g2_tiehi \mem.mem_internal.code_mem[58][3]$_SDFFCE_PN0P__3027  (.L_HI(net3027));
 sg13g2_tiehi \mem.mem_internal.code_mem[58][4]$_SDFFCE_PN0P__3028  (.L_HI(net3028));
 sg13g2_tiehi \mem.mem_internal.code_mem[58][5]$_SDFFCE_PN0P__3029  (.L_HI(net3029));
 sg13g2_tiehi \mem.mem_internal.code_mem[58][6]$_SDFFCE_PN0P__3030  (.L_HI(net3030));
 sg13g2_tiehi \mem.mem_internal.code_mem[58][7]$_SDFFCE_PN0P__3031  (.L_HI(net3031));
 sg13g2_tiehi \mem.mem_internal.code_mem[59][0]$_SDFFCE_PN0P__3032  (.L_HI(net3032));
 sg13g2_tiehi \mem.mem_internal.code_mem[59][1]$_SDFFCE_PN0P__3033  (.L_HI(net3033));
 sg13g2_tiehi \mem.mem_internal.code_mem[59][2]$_SDFFCE_PN0P__3034  (.L_HI(net3034));
 sg13g2_tiehi \mem.mem_internal.code_mem[59][3]$_SDFFCE_PN0P__3035  (.L_HI(net3035));
 sg13g2_tiehi \mem.mem_internal.code_mem[59][4]$_SDFFCE_PN0P__3036  (.L_HI(net3036));
 sg13g2_tiehi \mem.mem_internal.code_mem[59][5]$_SDFFCE_PN0P__3037  (.L_HI(net3037));
 sg13g2_tiehi \mem.mem_internal.code_mem[59][6]$_SDFFCE_PN0P__3038  (.L_HI(net3038));
 sg13g2_tiehi \mem.mem_internal.code_mem[59][7]$_SDFFCE_PN0P__3039  (.L_HI(net3039));
 sg13g2_tiehi \mem.mem_internal.code_mem[5][0]$_SDFFCE_PN0P__3040  (.L_HI(net3040));
 sg13g2_tiehi \mem.mem_internal.code_mem[5][1]$_SDFFCE_PN0P__3041  (.L_HI(net3041));
 sg13g2_tiehi \mem.mem_internal.code_mem[5][2]$_SDFFCE_PN0P__3042  (.L_HI(net3042));
 sg13g2_tiehi \mem.mem_internal.code_mem[5][3]$_SDFFCE_PN0P__3043  (.L_HI(net3043));
 sg13g2_tiehi \mem.mem_internal.code_mem[5][4]$_SDFFCE_PN0P__3044  (.L_HI(net3044));
 sg13g2_tiehi \mem.mem_internal.code_mem[5][5]$_SDFFCE_PN0P__3045  (.L_HI(net3045));
 sg13g2_tiehi \mem.mem_internal.code_mem[5][6]$_SDFFCE_PN0P__3046  (.L_HI(net3046));
 sg13g2_tiehi \mem.mem_internal.code_mem[5][7]$_SDFFCE_PN0P__3047  (.L_HI(net3047));
 sg13g2_tiehi \mem.mem_internal.code_mem[60][0]$_SDFFCE_PN0P__3048  (.L_HI(net3048));
 sg13g2_tiehi \mem.mem_internal.code_mem[60][1]$_SDFFCE_PN0P__3049  (.L_HI(net3049));
 sg13g2_tiehi \mem.mem_internal.code_mem[60][2]$_SDFFCE_PN0P__3050  (.L_HI(net3050));
 sg13g2_tiehi \mem.mem_internal.code_mem[60][3]$_SDFFCE_PN0P__3051  (.L_HI(net3051));
 sg13g2_tiehi \mem.mem_internal.code_mem[60][4]$_SDFFCE_PN0P__3052  (.L_HI(net3052));
 sg13g2_tiehi \mem.mem_internal.code_mem[60][5]$_SDFFCE_PN0P__3053  (.L_HI(net3053));
 sg13g2_tiehi \mem.mem_internal.code_mem[60][6]$_SDFFCE_PN0P__3054  (.L_HI(net3054));
 sg13g2_tiehi \mem.mem_internal.code_mem[60][7]$_SDFFCE_PN0P__3055  (.L_HI(net3055));
 sg13g2_tiehi \mem.mem_internal.code_mem[61][0]$_SDFFCE_PN0P__3056  (.L_HI(net3056));
 sg13g2_tiehi \mem.mem_internal.code_mem[61][1]$_SDFFCE_PN0P__3057  (.L_HI(net3057));
 sg13g2_tiehi \mem.mem_internal.code_mem[61][2]$_SDFFCE_PN0P__3058  (.L_HI(net3058));
 sg13g2_tiehi \mem.mem_internal.code_mem[61][3]$_SDFFCE_PN0P__3059  (.L_HI(net3059));
 sg13g2_tiehi \mem.mem_internal.code_mem[61][4]$_SDFFCE_PN0P__3060  (.L_HI(net3060));
 sg13g2_tiehi \mem.mem_internal.code_mem[61][5]$_SDFFCE_PN0P__3061  (.L_HI(net3061));
 sg13g2_tiehi \mem.mem_internal.code_mem[61][6]$_SDFFCE_PN0P__3062  (.L_HI(net3062));
 sg13g2_tiehi \mem.mem_internal.code_mem[61][7]$_SDFFCE_PN0P__3063  (.L_HI(net3063));
 sg13g2_tiehi \mem.mem_internal.code_mem[62][0]$_SDFFCE_PN0P__3064  (.L_HI(net3064));
 sg13g2_tiehi \mem.mem_internal.code_mem[62][1]$_SDFFCE_PN0P__3065  (.L_HI(net3065));
 sg13g2_tiehi \mem.mem_internal.code_mem[62][2]$_SDFFCE_PN0P__3066  (.L_HI(net3066));
 sg13g2_tiehi \mem.mem_internal.code_mem[62][3]$_SDFFCE_PN0P__3067  (.L_HI(net3067));
 sg13g2_tiehi \mem.mem_internal.code_mem[62][4]$_SDFFCE_PN0P__3068  (.L_HI(net3068));
 sg13g2_tiehi \mem.mem_internal.code_mem[62][5]$_SDFFCE_PN0P__3069  (.L_HI(net3069));
 sg13g2_tiehi \mem.mem_internal.code_mem[62][6]$_SDFFCE_PN0P__3070  (.L_HI(net3070));
 sg13g2_tiehi \mem.mem_internal.code_mem[62][7]$_SDFFCE_PN0P__3071  (.L_HI(net3071));
 sg13g2_tiehi \mem.mem_internal.code_mem[63][0]$_SDFFCE_PN0P__3072  (.L_HI(net3072));
 sg13g2_tiehi \mem.mem_internal.code_mem[63][1]$_SDFFCE_PN0P__3073  (.L_HI(net3073));
 sg13g2_tiehi \mem.mem_internal.code_mem[63][2]$_SDFFCE_PN0P__3074  (.L_HI(net3074));
 sg13g2_tiehi \mem.mem_internal.code_mem[63][3]$_SDFFCE_PN0P__3075  (.L_HI(net3075));
 sg13g2_tiehi \mem.mem_internal.code_mem[63][4]$_SDFFCE_PN0P__3076  (.L_HI(net3076));
 sg13g2_tiehi \mem.mem_internal.code_mem[63][5]$_SDFFCE_PN0P__3077  (.L_HI(net3077));
 sg13g2_tiehi \mem.mem_internal.code_mem[63][6]$_SDFFCE_PN0P__3078  (.L_HI(net3078));
 sg13g2_tiehi \mem.mem_internal.code_mem[63][7]$_SDFFCE_PN0P__3079  (.L_HI(net3079));
 sg13g2_tiehi \mem.mem_internal.code_mem[64][0]$_SDFFCE_PN0P__3080  (.L_HI(net3080));
 sg13g2_tiehi \mem.mem_internal.code_mem[64][1]$_SDFFCE_PN0P__3081  (.L_HI(net3081));
 sg13g2_tiehi \mem.mem_internal.code_mem[64][2]$_SDFFCE_PN0P__3082  (.L_HI(net3082));
 sg13g2_tiehi \mem.mem_internal.code_mem[64][3]$_SDFFCE_PN0P__3083  (.L_HI(net3083));
 sg13g2_tiehi \mem.mem_internal.code_mem[64][4]$_SDFFCE_PN0P__3084  (.L_HI(net3084));
 sg13g2_tiehi \mem.mem_internal.code_mem[64][5]$_SDFFCE_PN0P__3085  (.L_HI(net3085));
 sg13g2_tiehi \mem.mem_internal.code_mem[64][6]$_SDFFCE_PN0P__3086  (.L_HI(net3086));
 sg13g2_tiehi \mem.mem_internal.code_mem[64][7]$_SDFFCE_PN0P__3087  (.L_HI(net3087));
 sg13g2_tiehi \mem.mem_internal.code_mem[65][0]$_SDFFCE_PN0P__3088  (.L_HI(net3088));
 sg13g2_tiehi \mem.mem_internal.code_mem[65][1]$_SDFFCE_PN0P__3089  (.L_HI(net3089));
 sg13g2_tiehi \mem.mem_internal.code_mem[65][2]$_SDFFCE_PN0P__3090  (.L_HI(net3090));
 sg13g2_tiehi \mem.mem_internal.code_mem[65][3]$_SDFFCE_PN0P__3091  (.L_HI(net3091));
 sg13g2_tiehi \mem.mem_internal.code_mem[65][4]$_SDFFCE_PN0P__3092  (.L_HI(net3092));
 sg13g2_tiehi \mem.mem_internal.code_mem[65][5]$_SDFFCE_PN0P__3093  (.L_HI(net3093));
 sg13g2_tiehi \mem.mem_internal.code_mem[65][6]$_SDFFCE_PN0P__3094  (.L_HI(net3094));
 sg13g2_tiehi \mem.mem_internal.code_mem[65][7]$_SDFFCE_PN0P__3095  (.L_HI(net3095));
 sg13g2_tiehi \mem.mem_internal.code_mem[66][0]$_SDFFCE_PN0P__3096  (.L_HI(net3096));
 sg13g2_tiehi \mem.mem_internal.code_mem[66][1]$_SDFFCE_PN0P__3097  (.L_HI(net3097));
 sg13g2_tiehi \mem.mem_internal.code_mem[66][2]$_SDFFCE_PN0P__3098  (.L_HI(net3098));
 sg13g2_tiehi \mem.mem_internal.code_mem[66][3]$_SDFFCE_PN0P__3099  (.L_HI(net3099));
 sg13g2_tiehi \mem.mem_internal.code_mem[66][4]$_SDFFCE_PN0P__3100  (.L_HI(net3100));
 sg13g2_tiehi \mem.mem_internal.code_mem[66][5]$_SDFFCE_PN0P__3101  (.L_HI(net3101));
 sg13g2_tiehi \mem.mem_internal.code_mem[66][6]$_SDFFCE_PN0P__3102  (.L_HI(net3102));
 sg13g2_tiehi \mem.mem_internal.code_mem[66][7]$_SDFFCE_PN0P__3103  (.L_HI(net3103));
 sg13g2_tiehi \mem.mem_internal.code_mem[67][0]$_SDFFCE_PN0P__3104  (.L_HI(net3104));
 sg13g2_tiehi \mem.mem_internal.code_mem[67][1]$_SDFFCE_PN0P__3105  (.L_HI(net3105));
 sg13g2_tiehi \mem.mem_internal.code_mem[67][2]$_SDFFCE_PN0P__3106  (.L_HI(net3106));
 sg13g2_tiehi \mem.mem_internal.code_mem[67][3]$_SDFFCE_PN0P__3107  (.L_HI(net3107));
 sg13g2_tiehi \mem.mem_internal.code_mem[67][4]$_SDFFCE_PN0P__3108  (.L_HI(net3108));
 sg13g2_tiehi \mem.mem_internal.code_mem[67][5]$_SDFFCE_PN0P__3109  (.L_HI(net3109));
 sg13g2_tiehi \mem.mem_internal.code_mem[67][6]$_SDFFCE_PN0P__3110  (.L_HI(net3110));
 sg13g2_tiehi \mem.mem_internal.code_mem[67][7]$_SDFFCE_PN0P__3111  (.L_HI(net3111));
 sg13g2_tiehi \mem.mem_internal.code_mem[68][0]$_SDFFCE_PN0P__3112  (.L_HI(net3112));
 sg13g2_tiehi \mem.mem_internal.code_mem[68][1]$_SDFFCE_PN0P__3113  (.L_HI(net3113));
 sg13g2_tiehi \mem.mem_internal.code_mem[68][2]$_SDFFCE_PN0P__3114  (.L_HI(net3114));
 sg13g2_tiehi \mem.mem_internal.code_mem[68][3]$_SDFFCE_PN0P__3115  (.L_HI(net3115));
 sg13g2_tiehi \mem.mem_internal.code_mem[68][4]$_SDFFCE_PN0P__3116  (.L_HI(net3116));
 sg13g2_tiehi \mem.mem_internal.code_mem[68][5]$_SDFFCE_PN0P__3117  (.L_HI(net3117));
 sg13g2_tiehi \mem.mem_internal.code_mem[68][6]$_SDFFCE_PN0P__3118  (.L_HI(net3118));
 sg13g2_tiehi \mem.mem_internal.code_mem[68][7]$_SDFFCE_PN0P__3119  (.L_HI(net3119));
 sg13g2_tiehi \mem.mem_internal.code_mem[69][0]$_SDFFCE_PN0P__3120  (.L_HI(net3120));
 sg13g2_tiehi \mem.mem_internal.code_mem[69][1]$_SDFFCE_PN0P__3121  (.L_HI(net3121));
 sg13g2_tiehi \mem.mem_internal.code_mem[69][2]$_SDFFCE_PN0P__3122  (.L_HI(net3122));
 sg13g2_tiehi \mem.mem_internal.code_mem[69][3]$_SDFFCE_PN0P__3123  (.L_HI(net3123));
 sg13g2_tiehi \mem.mem_internal.code_mem[69][4]$_SDFFCE_PN0P__3124  (.L_HI(net3124));
 sg13g2_tiehi \mem.mem_internal.code_mem[69][5]$_SDFFCE_PN0P__3125  (.L_HI(net3125));
 sg13g2_tiehi \mem.mem_internal.code_mem[69][6]$_SDFFCE_PN0P__3126  (.L_HI(net3126));
 sg13g2_tiehi \mem.mem_internal.code_mem[69][7]$_SDFFCE_PN0P__3127  (.L_HI(net3127));
 sg13g2_tiehi \mem.mem_internal.code_mem[6][0]$_SDFFCE_PN0P__3128  (.L_HI(net3128));
 sg13g2_tiehi \mem.mem_internal.code_mem[6][1]$_SDFFCE_PN0P__3129  (.L_HI(net3129));
 sg13g2_tiehi \mem.mem_internal.code_mem[6][2]$_SDFFCE_PN0P__3130  (.L_HI(net3130));
 sg13g2_tiehi \mem.mem_internal.code_mem[6][3]$_SDFFCE_PN0P__3131  (.L_HI(net3131));
 sg13g2_tiehi \mem.mem_internal.code_mem[6][4]$_SDFFCE_PN0P__3132  (.L_HI(net3132));
 sg13g2_tiehi \mem.mem_internal.code_mem[6][5]$_SDFFCE_PN0P__3133  (.L_HI(net3133));
 sg13g2_tiehi \mem.mem_internal.code_mem[6][6]$_SDFFCE_PN0P__3134  (.L_HI(net3134));
 sg13g2_tiehi \mem.mem_internal.code_mem[6][7]$_SDFFCE_PN0P__3135  (.L_HI(net3135));
 sg13g2_tiehi \mem.mem_internal.code_mem[70][0]$_SDFFCE_PN0P__3136  (.L_HI(net3136));
 sg13g2_tiehi \mem.mem_internal.code_mem[70][1]$_SDFFCE_PN0P__3137  (.L_HI(net3137));
 sg13g2_tiehi \mem.mem_internal.code_mem[70][2]$_SDFFCE_PN0P__3138  (.L_HI(net3138));
 sg13g2_tiehi \mem.mem_internal.code_mem[70][3]$_SDFFCE_PN0P__3139  (.L_HI(net3139));
 sg13g2_tiehi \mem.mem_internal.code_mem[70][4]$_SDFFCE_PN0P__3140  (.L_HI(net3140));
 sg13g2_tiehi \mem.mem_internal.code_mem[70][5]$_SDFFCE_PN0P__3141  (.L_HI(net3141));
 sg13g2_tiehi \mem.mem_internal.code_mem[70][6]$_SDFFCE_PN0P__3142  (.L_HI(net3142));
 sg13g2_tiehi \mem.mem_internal.code_mem[70][7]$_SDFFCE_PN0P__3143  (.L_HI(net3143));
 sg13g2_tiehi \mem.mem_internal.code_mem[71][0]$_SDFFCE_PN0P__3144  (.L_HI(net3144));
 sg13g2_tiehi \mem.mem_internal.code_mem[71][1]$_SDFFCE_PN0P__3145  (.L_HI(net3145));
 sg13g2_tiehi \mem.mem_internal.code_mem[71][2]$_SDFFCE_PN0P__3146  (.L_HI(net3146));
 sg13g2_tiehi \mem.mem_internal.code_mem[71][3]$_SDFFCE_PN0P__3147  (.L_HI(net3147));
 sg13g2_tiehi \mem.mem_internal.code_mem[71][4]$_SDFFCE_PN0P__3148  (.L_HI(net3148));
 sg13g2_tiehi \mem.mem_internal.code_mem[71][5]$_SDFFCE_PN0P__3149  (.L_HI(net3149));
 sg13g2_tiehi \mem.mem_internal.code_mem[71][6]$_SDFFCE_PN0P__3150  (.L_HI(net3150));
 sg13g2_tiehi \mem.mem_internal.code_mem[71][7]$_SDFFCE_PN0P__3151  (.L_HI(net3151));
 sg13g2_tiehi \mem.mem_internal.code_mem[72][0]$_SDFFCE_PN0P__3152  (.L_HI(net3152));
 sg13g2_tiehi \mem.mem_internal.code_mem[72][1]$_SDFFCE_PN0P__3153  (.L_HI(net3153));
 sg13g2_tiehi \mem.mem_internal.code_mem[72][2]$_SDFFCE_PN0P__3154  (.L_HI(net3154));
 sg13g2_tiehi \mem.mem_internal.code_mem[72][3]$_SDFFCE_PN0P__3155  (.L_HI(net3155));
 sg13g2_tiehi \mem.mem_internal.code_mem[72][4]$_SDFFCE_PN0P__3156  (.L_HI(net3156));
 sg13g2_tiehi \mem.mem_internal.code_mem[72][5]$_SDFFCE_PN0P__3157  (.L_HI(net3157));
 sg13g2_tiehi \mem.mem_internal.code_mem[72][6]$_SDFFCE_PN0P__3158  (.L_HI(net3158));
 sg13g2_tiehi \mem.mem_internal.code_mem[72][7]$_SDFFCE_PN0P__3159  (.L_HI(net3159));
 sg13g2_tiehi \mem.mem_internal.code_mem[73][0]$_SDFFCE_PN0P__3160  (.L_HI(net3160));
 sg13g2_tiehi \mem.mem_internal.code_mem[73][1]$_SDFFCE_PN0P__3161  (.L_HI(net3161));
 sg13g2_tiehi \mem.mem_internal.code_mem[73][2]$_SDFFCE_PN0P__3162  (.L_HI(net3162));
 sg13g2_tiehi \mem.mem_internal.code_mem[73][3]$_SDFFCE_PN0P__3163  (.L_HI(net3163));
 sg13g2_tiehi \mem.mem_internal.code_mem[73][4]$_SDFFCE_PN0P__3164  (.L_HI(net3164));
 sg13g2_tiehi \mem.mem_internal.code_mem[73][5]$_SDFFCE_PN0P__3165  (.L_HI(net3165));
 sg13g2_tiehi \mem.mem_internal.code_mem[73][6]$_SDFFCE_PN0P__3166  (.L_HI(net3166));
 sg13g2_tiehi \mem.mem_internal.code_mem[73][7]$_SDFFCE_PN0P__3167  (.L_HI(net3167));
 sg13g2_tiehi \mem.mem_internal.code_mem[74][0]$_SDFFCE_PN0P__3168  (.L_HI(net3168));
 sg13g2_tiehi \mem.mem_internal.code_mem[74][1]$_SDFFCE_PN0P__3169  (.L_HI(net3169));
 sg13g2_tiehi \mem.mem_internal.code_mem[74][2]$_SDFFCE_PN0P__3170  (.L_HI(net3170));
 sg13g2_tiehi \mem.mem_internal.code_mem[74][3]$_SDFFCE_PN0P__3171  (.L_HI(net3171));
 sg13g2_tiehi \mem.mem_internal.code_mem[74][4]$_SDFFCE_PN0P__3172  (.L_HI(net3172));
 sg13g2_tiehi \mem.mem_internal.code_mem[74][5]$_SDFFCE_PN0P__3173  (.L_HI(net3173));
 sg13g2_tiehi \mem.mem_internal.code_mem[74][6]$_SDFFCE_PN0P__3174  (.L_HI(net3174));
 sg13g2_tiehi \mem.mem_internal.code_mem[74][7]$_SDFFCE_PN0P__3175  (.L_HI(net3175));
 sg13g2_tiehi \mem.mem_internal.code_mem[75][0]$_SDFFCE_PN0P__3176  (.L_HI(net3176));
 sg13g2_tiehi \mem.mem_internal.code_mem[75][1]$_SDFFCE_PN0P__3177  (.L_HI(net3177));
 sg13g2_tiehi \mem.mem_internal.code_mem[75][2]$_SDFFCE_PN0P__3178  (.L_HI(net3178));
 sg13g2_tiehi \mem.mem_internal.code_mem[75][3]$_SDFFCE_PN0P__3179  (.L_HI(net3179));
 sg13g2_tiehi \mem.mem_internal.code_mem[75][4]$_SDFFCE_PN0P__3180  (.L_HI(net3180));
 sg13g2_tiehi \mem.mem_internal.code_mem[75][5]$_SDFFCE_PN0P__3181  (.L_HI(net3181));
 sg13g2_tiehi \mem.mem_internal.code_mem[75][6]$_SDFFCE_PN0P__3182  (.L_HI(net3182));
 sg13g2_tiehi \mem.mem_internal.code_mem[75][7]$_SDFFCE_PN0P__3183  (.L_HI(net3183));
 sg13g2_tiehi \mem.mem_internal.code_mem[76][0]$_SDFFCE_PN0P__3184  (.L_HI(net3184));
 sg13g2_tiehi \mem.mem_internal.code_mem[76][1]$_SDFFCE_PN0P__3185  (.L_HI(net3185));
 sg13g2_tiehi \mem.mem_internal.code_mem[76][2]$_SDFFCE_PN0P__3186  (.L_HI(net3186));
 sg13g2_tiehi \mem.mem_internal.code_mem[76][3]$_SDFFCE_PN0P__3187  (.L_HI(net3187));
 sg13g2_tiehi \mem.mem_internal.code_mem[76][4]$_SDFFCE_PN0P__3188  (.L_HI(net3188));
 sg13g2_tiehi \mem.mem_internal.code_mem[76][5]$_SDFFCE_PN0P__3189  (.L_HI(net3189));
 sg13g2_tiehi \mem.mem_internal.code_mem[76][6]$_SDFFCE_PN0P__3190  (.L_HI(net3190));
 sg13g2_tiehi \mem.mem_internal.code_mem[76][7]$_SDFFCE_PN0P__3191  (.L_HI(net3191));
 sg13g2_tiehi \mem.mem_internal.code_mem[77][0]$_SDFFCE_PN0P__3192  (.L_HI(net3192));
 sg13g2_tiehi \mem.mem_internal.code_mem[77][1]$_SDFFCE_PN0P__3193  (.L_HI(net3193));
 sg13g2_tiehi \mem.mem_internal.code_mem[77][2]$_SDFFCE_PN0P__3194  (.L_HI(net3194));
 sg13g2_tiehi \mem.mem_internal.code_mem[77][3]$_SDFFCE_PN0P__3195  (.L_HI(net3195));
 sg13g2_tiehi \mem.mem_internal.code_mem[77][4]$_SDFFCE_PN0P__3196  (.L_HI(net3196));
 sg13g2_tiehi \mem.mem_internal.code_mem[77][5]$_SDFFCE_PN0P__3197  (.L_HI(net3197));
 sg13g2_tiehi \mem.mem_internal.code_mem[77][6]$_SDFFCE_PN0P__3198  (.L_HI(net3198));
 sg13g2_tiehi \mem.mem_internal.code_mem[77][7]$_SDFFCE_PN0P__3199  (.L_HI(net3199));
 sg13g2_tiehi \mem.mem_internal.code_mem[78][0]$_SDFFCE_PN0P__3200  (.L_HI(net3200));
 sg13g2_tiehi \mem.mem_internal.code_mem[78][1]$_SDFFCE_PN0P__3201  (.L_HI(net3201));
 sg13g2_tiehi \mem.mem_internal.code_mem[78][2]$_SDFFCE_PN0P__3202  (.L_HI(net3202));
 sg13g2_tiehi \mem.mem_internal.code_mem[78][3]$_SDFFCE_PN0P__3203  (.L_HI(net3203));
 sg13g2_tiehi \mem.mem_internal.code_mem[78][4]$_SDFFCE_PN0P__3204  (.L_HI(net3204));
 sg13g2_tiehi \mem.mem_internal.code_mem[78][5]$_SDFFCE_PN0P__3205  (.L_HI(net3205));
 sg13g2_tiehi \mem.mem_internal.code_mem[78][6]$_SDFFCE_PN0P__3206  (.L_HI(net3206));
 sg13g2_tiehi \mem.mem_internal.code_mem[78][7]$_SDFFCE_PN0P__3207  (.L_HI(net3207));
 sg13g2_tiehi \mem.mem_internal.code_mem[79][0]$_SDFFCE_PN0P__3208  (.L_HI(net3208));
 sg13g2_tiehi \mem.mem_internal.code_mem[79][1]$_SDFFCE_PN0P__3209  (.L_HI(net3209));
 sg13g2_tiehi \mem.mem_internal.code_mem[79][2]$_SDFFCE_PN0P__3210  (.L_HI(net3210));
 sg13g2_tiehi \mem.mem_internal.code_mem[79][3]$_SDFFCE_PN0P__3211  (.L_HI(net3211));
 sg13g2_tiehi \mem.mem_internal.code_mem[79][4]$_SDFFCE_PN0P__3212  (.L_HI(net3212));
 sg13g2_tiehi \mem.mem_internal.code_mem[79][5]$_SDFFCE_PN0P__3213  (.L_HI(net3213));
 sg13g2_tiehi \mem.mem_internal.code_mem[79][6]$_SDFFCE_PN0P__3214  (.L_HI(net3214));
 sg13g2_tiehi \mem.mem_internal.code_mem[79][7]$_SDFFCE_PN0P__3215  (.L_HI(net3215));
 sg13g2_tiehi \mem.mem_internal.code_mem[7][0]$_SDFFCE_PN0P__3216  (.L_HI(net3216));
 sg13g2_tiehi \mem.mem_internal.code_mem[7][1]$_SDFFCE_PN0P__3217  (.L_HI(net3217));
 sg13g2_tiehi \mem.mem_internal.code_mem[7][2]$_SDFFCE_PN0P__3218  (.L_HI(net3218));
 sg13g2_tiehi \mem.mem_internal.code_mem[7][3]$_SDFFCE_PN0P__3219  (.L_HI(net3219));
 sg13g2_tiehi \mem.mem_internal.code_mem[7][4]$_SDFFCE_PN0P__3220  (.L_HI(net3220));
 sg13g2_tiehi \mem.mem_internal.code_mem[7][5]$_SDFFCE_PN0P__3221  (.L_HI(net3221));
 sg13g2_tiehi \mem.mem_internal.code_mem[7][6]$_SDFFCE_PN0P__3222  (.L_HI(net3222));
 sg13g2_tiehi \mem.mem_internal.code_mem[7][7]$_SDFFCE_PN0P__3223  (.L_HI(net3223));
 sg13g2_tiehi \mem.mem_internal.code_mem[80][0]$_SDFFCE_PN0P__3224  (.L_HI(net3224));
 sg13g2_tiehi \mem.mem_internal.code_mem[80][1]$_SDFFCE_PN0P__3225  (.L_HI(net3225));
 sg13g2_tiehi \mem.mem_internal.code_mem[80][2]$_SDFFCE_PN0P__3226  (.L_HI(net3226));
 sg13g2_tiehi \mem.mem_internal.code_mem[80][3]$_SDFFCE_PN0P__3227  (.L_HI(net3227));
 sg13g2_tiehi \mem.mem_internal.code_mem[80][4]$_SDFFCE_PN0P__3228  (.L_HI(net3228));
 sg13g2_tiehi \mem.mem_internal.code_mem[80][5]$_SDFFCE_PN0P__3229  (.L_HI(net3229));
 sg13g2_tiehi \mem.mem_internal.code_mem[80][6]$_SDFFCE_PN0P__3230  (.L_HI(net3230));
 sg13g2_tiehi \mem.mem_internal.code_mem[80][7]$_SDFFCE_PN0P__3231  (.L_HI(net3231));
 sg13g2_tiehi \mem.mem_internal.code_mem[81][0]$_SDFFCE_PN0P__3232  (.L_HI(net3232));
 sg13g2_tiehi \mem.mem_internal.code_mem[81][1]$_SDFFCE_PN0P__3233  (.L_HI(net3233));
 sg13g2_tiehi \mem.mem_internal.code_mem[81][2]$_SDFFCE_PN0P__3234  (.L_HI(net3234));
 sg13g2_tiehi \mem.mem_internal.code_mem[81][3]$_SDFFCE_PN0P__3235  (.L_HI(net3235));
 sg13g2_tiehi \mem.mem_internal.code_mem[81][4]$_SDFFCE_PN0P__3236  (.L_HI(net3236));
 sg13g2_tiehi \mem.mem_internal.code_mem[81][5]$_SDFFCE_PN0P__3237  (.L_HI(net3237));
 sg13g2_tiehi \mem.mem_internal.code_mem[81][6]$_SDFFCE_PN0P__3238  (.L_HI(net3238));
 sg13g2_tiehi \mem.mem_internal.code_mem[81][7]$_SDFFCE_PN0P__3239  (.L_HI(net3239));
 sg13g2_tiehi \mem.mem_internal.code_mem[82][0]$_SDFFCE_PN0P__3240  (.L_HI(net3240));
 sg13g2_tiehi \mem.mem_internal.code_mem[82][1]$_SDFFCE_PN0P__3241  (.L_HI(net3241));
 sg13g2_tiehi \mem.mem_internal.code_mem[82][2]$_SDFFCE_PN0P__3242  (.L_HI(net3242));
 sg13g2_tiehi \mem.mem_internal.code_mem[82][3]$_SDFFCE_PN0P__3243  (.L_HI(net3243));
 sg13g2_tiehi \mem.mem_internal.code_mem[82][4]$_SDFFCE_PN0P__3244  (.L_HI(net3244));
 sg13g2_tiehi \mem.mem_internal.code_mem[82][5]$_SDFFCE_PN0P__3245  (.L_HI(net3245));
 sg13g2_tiehi \mem.mem_internal.code_mem[82][6]$_SDFFCE_PN0P__3246  (.L_HI(net3246));
 sg13g2_tiehi \mem.mem_internal.code_mem[82][7]$_SDFFCE_PN0P__3247  (.L_HI(net3247));
 sg13g2_tiehi \mem.mem_internal.code_mem[83][0]$_SDFFCE_PN0P__3248  (.L_HI(net3248));
 sg13g2_tiehi \mem.mem_internal.code_mem[83][1]$_SDFFCE_PN0P__3249  (.L_HI(net3249));
 sg13g2_tiehi \mem.mem_internal.code_mem[83][2]$_SDFFCE_PN0P__3250  (.L_HI(net3250));
 sg13g2_tiehi \mem.mem_internal.code_mem[83][3]$_SDFFCE_PN0P__3251  (.L_HI(net3251));
 sg13g2_tiehi \mem.mem_internal.code_mem[83][4]$_SDFFCE_PN0P__3252  (.L_HI(net3252));
 sg13g2_tiehi \mem.mem_internal.code_mem[83][5]$_SDFFCE_PN0P__3253  (.L_HI(net3253));
 sg13g2_tiehi \mem.mem_internal.code_mem[83][6]$_SDFFCE_PN0P__3254  (.L_HI(net3254));
 sg13g2_tiehi \mem.mem_internal.code_mem[83][7]$_SDFFCE_PN0P__3255  (.L_HI(net3255));
 sg13g2_tiehi \mem.mem_internal.code_mem[84][0]$_SDFFCE_PN0P__3256  (.L_HI(net3256));
 sg13g2_tiehi \mem.mem_internal.code_mem[84][1]$_SDFFCE_PN0P__3257  (.L_HI(net3257));
 sg13g2_tiehi \mem.mem_internal.code_mem[84][2]$_SDFFCE_PN0P__3258  (.L_HI(net3258));
 sg13g2_tiehi \mem.mem_internal.code_mem[84][3]$_SDFFCE_PN0P__3259  (.L_HI(net3259));
 sg13g2_tiehi \mem.mem_internal.code_mem[84][4]$_SDFFCE_PN0P__3260  (.L_HI(net3260));
 sg13g2_tiehi \mem.mem_internal.code_mem[84][5]$_SDFFCE_PN0P__3261  (.L_HI(net3261));
 sg13g2_tiehi \mem.mem_internal.code_mem[84][6]$_SDFFCE_PN0P__3262  (.L_HI(net3262));
 sg13g2_tiehi \mem.mem_internal.code_mem[84][7]$_SDFFCE_PN0P__3263  (.L_HI(net3263));
 sg13g2_tiehi \mem.mem_internal.code_mem[85][0]$_SDFFCE_PN0P__3264  (.L_HI(net3264));
 sg13g2_tiehi \mem.mem_internal.code_mem[85][1]$_SDFFCE_PN0P__3265  (.L_HI(net3265));
 sg13g2_tiehi \mem.mem_internal.code_mem[85][2]$_SDFFCE_PN0P__3266  (.L_HI(net3266));
 sg13g2_tiehi \mem.mem_internal.code_mem[85][3]$_SDFFCE_PN0P__3267  (.L_HI(net3267));
 sg13g2_tiehi \mem.mem_internal.code_mem[85][4]$_SDFFCE_PN0P__3268  (.L_HI(net3268));
 sg13g2_tiehi \mem.mem_internal.code_mem[85][5]$_SDFFCE_PN0P__3269  (.L_HI(net3269));
 sg13g2_tiehi \mem.mem_internal.code_mem[85][6]$_SDFFCE_PN0P__3270  (.L_HI(net3270));
 sg13g2_tiehi \mem.mem_internal.code_mem[85][7]$_SDFFCE_PN0P__3271  (.L_HI(net3271));
 sg13g2_tiehi \mem.mem_internal.code_mem[86][0]$_SDFFCE_PN0P__3272  (.L_HI(net3272));
 sg13g2_tiehi \mem.mem_internal.code_mem[86][1]$_SDFFCE_PN0P__3273  (.L_HI(net3273));
 sg13g2_tiehi \mem.mem_internal.code_mem[86][2]$_SDFFCE_PN0P__3274  (.L_HI(net3274));
 sg13g2_tiehi \mem.mem_internal.code_mem[86][3]$_SDFFCE_PN0P__3275  (.L_HI(net3275));
 sg13g2_tiehi \mem.mem_internal.code_mem[86][4]$_SDFFCE_PN0P__3276  (.L_HI(net3276));
 sg13g2_tiehi \mem.mem_internal.code_mem[86][5]$_SDFFCE_PN0P__3277  (.L_HI(net3277));
 sg13g2_tiehi \mem.mem_internal.code_mem[86][6]$_SDFFCE_PN0P__3278  (.L_HI(net3278));
 sg13g2_tiehi \mem.mem_internal.code_mem[86][7]$_SDFFCE_PN0P__3279  (.L_HI(net3279));
 sg13g2_tiehi \mem.mem_internal.code_mem[87][0]$_SDFFCE_PN0P__3280  (.L_HI(net3280));
 sg13g2_tiehi \mem.mem_internal.code_mem[87][1]$_SDFFCE_PN0P__3281  (.L_HI(net3281));
 sg13g2_tiehi \mem.mem_internal.code_mem[87][2]$_SDFFCE_PN0P__3282  (.L_HI(net3282));
 sg13g2_tiehi \mem.mem_internal.code_mem[87][3]$_SDFFCE_PN0P__3283  (.L_HI(net3283));
 sg13g2_tiehi \mem.mem_internal.code_mem[87][4]$_SDFFCE_PN0P__3284  (.L_HI(net3284));
 sg13g2_tiehi \mem.mem_internal.code_mem[87][5]$_SDFFCE_PN0P__3285  (.L_HI(net3285));
 sg13g2_tiehi \mem.mem_internal.code_mem[87][6]$_SDFFCE_PN0P__3286  (.L_HI(net3286));
 sg13g2_tiehi \mem.mem_internal.code_mem[87][7]$_SDFFCE_PN0P__3287  (.L_HI(net3287));
 sg13g2_tiehi \mem.mem_internal.code_mem[88][0]$_SDFFCE_PN0P__3288  (.L_HI(net3288));
 sg13g2_tiehi \mem.mem_internal.code_mem[88][1]$_SDFFCE_PN0P__3289  (.L_HI(net3289));
 sg13g2_tiehi \mem.mem_internal.code_mem[88][2]$_SDFFCE_PN0P__3290  (.L_HI(net3290));
 sg13g2_tiehi \mem.mem_internal.code_mem[88][3]$_SDFFCE_PN0P__3291  (.L_HI(net3291));
 sg13g2_tiehi \mem.mem_internal.code_mem[88][4]$_SDFFCE_PN0P__3292  (.L_HI(net3292));
 sg13g2_tiehi \mem.mem_internal.code_mem[88][5]$_SDFFCE_PN0P__3293  (.L_HI(net3293));
 sg13g2_tiehi \mem.mem_internal.code_mem[88][6]$_SDFFCE_PN0P__3294  (.L_HI(net3294));
 sg13g2_tiehi \mem.mem_internal.code_mem[88][7]$_SDFFCE_PN0P__3295  (.L_HI(net3295));
 sg13g2_tiehi \mem.mem_internal.code_mem[89][0]$_SDFFCE_PN0P__3296  (.L_HI(net3296));
 sg13g2_tiehi \mem.mem_internal.code_mem[89][1]$_SDFFCE_PN0P__3297  (.L_HI(net3297));
 sg13g2_tiehi \mem.mem_internal.code_mem[89][2]$_SDFFCE_PN0P__3298  (.L_HI(net3298));
 sg13g2_tiehi \mem.mem_internal.code_mem[89][3]$_SDFFCE_PN0P__3299  (.L_HI(net3299));
 sg13g2_tiehi \mem.mem_internal.code_mem[89][4]$_SDFFCE_PN0P__3300  (.L_HI(net3300));
 sg13g2_tiehi \mem.mem_internal.code_mem[89][5]$_SDFFCE_PN0P__3301  (.L_HI(net3301));
 sg13g2_tiehi \mem.mem_internal.code_mem[89][6]$_SDFFCE_PN0P__3302  (.L_HI(net3302));
 sg13g2_tiehi \mem.mem_internal.code_mem[89][7]$_SDFFCE_PN0P__3303  (.L_HI(net3303));
 sg13g2_tiehi \mem.mem_internal.code_mem[8][0]$_SDFFCE_PN0P__3304  (.L_HI(net3304));
 sg13g2_tiehi \mem.mem_internal.code_mem[8][1]$_SDFFCE_PN0P__3305  (.L_HI(net3305));
 sg13g2_tiehi \mem.mem_internal.code_mem[8][2]$_SDFFCE_PN0P__3306  (.L_HI(net3306));
 sg13g2_tiehi \mem.mem_internal.code_mem[8][3]$_SDFFCE_PN0P__3307  (.L_HI(net3307));
 sg13g2_tiehi \mem.mem_internal.code_mem[8][4]$_SDFFCE_PN0P__3308  (.L_HI(net3308));
 sg13g2_tiehi \mem.mem_internal.code_mem[8][5]$_SDFFCE_PN0P__3309  (.L_HI(net3309));
 sg13g2_tiehi \mem.mem_internal.code_mem[8][6]$_SDFFCE_PN0P__3310  (.L_HI(net3310));
 sg13g2_tiehi \mem.mem_internal.code_mem[8][7]$_SDFFCE_PN0P__3311  (.L_HI(net3311));
 sg13g2_tiehi \mem.mem_internal.code_mem[90][0]$_SDFFCE_PN0P__3312  (.L_HI(net3312));
 sg13g2_tiehi \mem.mem_internal.code_mem[90][1]$_SDFFCE_PN0P__3313  (.L_HI(net3313));
 sg13g2_tiehi \mem.mem_internal.code_mem[90][2]$_SDFFCE_PN0P__3314  (.L_HI(net3314));
 sg13g2_tiehi \mem.mem_internal.code_mem[90][3]$_SDFFCE_PN0P__3315  (.L_HI(net3315));
 sg13g2_tiehi \mem.mem_internal.code_mem[90][4]$_SDFFCE_PN0P__3316  (.L_HI(net3316));
 sg13g2_tiehi \mem.mem_internal.code_mem[90][5]$_SDFFCE_PN0P__3317  (.L_HI(net3317));
 sg13g2_tiehi \mem.mem_internal.code_mem[90][6]$_SDFFCE_PN0P__3318  (.L_HI(net3318));
 sg13g2_tiehi \mem.mem_internal.code_mem[90][7]$_SDFFCE_PN0P__3319  (.L_HI(net3319));
 sg13g2_tiehi \mem.mem_internal.code_mem[91][0]$_SDFFCE_PN0P__3320  (.L_HI(net3320));
 sg13g2_tiehi \mem.mem_internal.code_mem[91][1]$_SDFFCE_PN0P__3321  (.L_HI(net3321));
 sg13g2_tiehi \mem.mem_internal.code_mem[91][2]$_SDFFCE_PN0P__3322  (.L_HI(net3322));
 sg13g2_tiehi \mem.mem_internal.code_mem[91][3]$_SDFFCE_PN0P__3323  (.L_HI(net3323));
 sg13g2_tiehi \mem.mem_internal.code_mem[91][4]$_SDFFCE_PN0P__3324  (.L_HI(net3324));
 sg13g2_tiehi \mem.mem_internal.code_mem[91][5]$_SDFFCE_PN0P__3325  (.L_HI(net3325));
 sg13g2_tiehi \mem.mem_internal.code_mem[91][6]$_SDFFCE_PN0P__3326  (.L_HI(net3326));
 sg13g2_tiehi \mem.mem_internal.code_mem[91][7]$_SDFFCE_PN0P__3327  (.L_HI(net3327));
 sg13g2_tiehi \mem.mem_internal.code_mem[92][0]$_SDFFCE_PN0P__3328  (.L_HI(net3328));
 sg13g2_tiehi \mem.mem_internal.code_mem[92][1]$_SDFFCE_PN0P__3329  (.L_HI(net3329));
 sg13g2_tiehi \mem.mem_internal.code_mem[92][2]$_SDFFCE_PN0P__3330  (.L_HI(net3330));
 sg13g2_tiehi \mem.mem_internal.code_mem[92][3]$_SDFFCE_PN0P__3331  (.L_HI(net3331));
 sg13g2_tiehi \mem.mem_internal.code_mem[92][4]$_SDFFCE_PN0P__3332  (.L_HI(net3332));
 sg13g2_tiehi \mem.mem_internal.code_mem[92][5]$_SDFFCE_PN0P__3333  (.L_HI(net3333));
 sg13g2_tiehi \mem.mem_internal.code_mem[92][6]$_SDFFCE_PN0P__3334  (.L_HI(net3334));
 sg13g2_tiehi \mem.mem_internal.code_mem[92][7]$_SDFFCE_PN0P__3335  (.L_HI(net3335));
 sg13g2_tiehi \mem.mem_internal.code_mem[93][0]$_SDFFCE_PN0P__3336  (.L_HI(net3336));
 sg13g2_tiehi \mem.mem_internal.code_mem[93][1]$_SDFFCE_PN0P__3337  (.L_HI(net3337));
 sg13g2_tiehi \mem.mem_internal.code_mem[93][2]$_SDFFCE_PN0P__3338  (.L_HI(net3338));
 sg13g2_tiehi \mem.mem_internal.code_mem[93][3]$_SDFFCE_PN0P__3339  (.L_HI(net3339));
 sg13g2_tiehi \mem.mem_internal.code_mem[93][4]$_SDFFCE_PN0P__3340  (.L_HI(net3340));
 sg13g2_tiehi \mem.mem_internal.code_mem[93][5]$_SDFFCE_PN0P__3341  (.L_HI(net3341));
 sg13g2_tiehi \mem.mem_internal.code_mem[93][6]$_SDFFCE_PN0P__3342  (.L_HI(net3342));
 sg13g2_tiehi \mem.mem_internal.code_mem[93][7]$_SDFFCE_PN0P__3343  (.L_HI(net3343));
 sg13g2_tiehi \mem.mem_internal.code_mem[94][0]$_SDFFCE_PN0P__3344  (.L_HI(net3344));
 sg13g2_tiehi \mem.mem_internal.code_mem[94][1]$_SDFFCE_PN0P__3345  (.L_HI(net3345));
 sg13g2_tiehi \mem.mem_internal.code_mem[94][2]$_SDFFCE_PN0P__3346  (.L_HI(net3346));
 sg13g2_tiehi \mem.mem_internal.code_mem[94][3]$_SDFFCE_PN0P__3347  (.L_HI(net3347));
 sg13g2_tiehi \mem.mem_internal.code_mem[94][4]$_SDFFCE_PN0P__3348  (.L_HI(net3348));
 sg13g2_tiehi \mem.mem_internal.code_mem[94][5]$_SDFFCE_PN0P__3349  (.L_HI(net3349));
 sg13g2_tiehi \mem.mem_internal.code_mem[94][6]$_SDFFCE_PN0P__3350  (.L_HI(net3350));
 sg13g2_tiehi \mem.mem_internal.code_mem[94][7]$_SDFFCE_PN0P__3351  (.L_HI(net3351));
 sg13g2_tiehi \mem.mem_internal.code_mem[95][0]$_SDFFCE_PN0P__3352  (.L_HI(net3352));
 sg13g2_tiehi \mem.mem_internal.code_mem[95][1]$_SDFFCE_PN0P__3353  (.L_HI(net3353));
 sg13g2_tiehi \mem.mem_internal.code_mem[95][2]$_SDFFCE_PN0P__3354  (.L_HI(net3354));
 sg13g2_tiehi \mem.mem_internal.code_mem[95][3]$_SDFFCE_PN0P__3355  (.L_HI(net3355));
 sg13g2_tiehi \mem.mem_internal.code_mem[95][4]$_SDFFCE_PN0P__3356  (.L_HI(net3356));
 sg13g2_tiehi \mem.mem_internal.code_mem[95][5]$_SDFFCE_PN0P__3357  (.L_HI(net3357));
 sg13g2_tiehi \mem.mem_internal.code_mem[95][6]$_SDFFCE_PN0P__3358  (.L_HI(net3358));
 sg13g2_tiehi \mem.mem_internal.code_mem[95][7]$_SDFFCE_PN0P__3359  (.L_HI(net3359));
 sg13g2_tiehi \mem.mem_internal.code_mem[96][0]$_SDFFCE_PN0P__3360  (.L_HI(net3360));
 sg13g2_tiehi \mem.mem_internal.code_mem[96][1]$_SDFFCE_PN0P__3361  (.L_HI(net3361));
 sg13g2_tiehi \mem.mem_internal.code_mem[96][2]$_SDFFCE_PN0P__3362  (.L_HI(net3362));
 sg13g2_tiehi \mem.mem_internal.code_mem[96][3]$_SDFFCE_PN0P__3363  (.L_HI(net3363));
 sg13g2_tiehi \mem.mem_internal.code_mem[96][4]$_SDFFCE_PN0P__3364  (.L_HI(net3364));
 sg13g2_tiehi \mem.mem_internal.code_mem[96][5]$_SDFFCE_PN0P__3365  (.L_HI(net3365));
 sg13g2_tiehi \mem.mem_internal.code_mem[96][6]$_SDFFCE_PN0P__3366  (.L_HI(net3366));
 sg13g2_tiehi \mem.mem_internal.code_mem[96][7]$_SDFFCE_PN0P__3367  (.L_HI(net3367));
 sg13g2_tiehi \mem.mem_internal.code_mem[97][0]$_SDFFCE_PN0P__3368  (.L_HI(net3368));
 sg13g2_tiehi \mem.mem_internal.code_mem[97][1]$_SDFFCE_PN0P__3369  (.L_HI(net3369));
 sg13g2_tiehi \mem.mem_internal.code_mem[97][2]$_SDFFCE_PN0P__3370  (.L_HI(net3370));
 sg13g2_tiehi \mem.mem_internal.code_mem[97][3]$_SDFFCE_PN0P__3371  (.L_HI(net3371));
 sg13g2_tiehi \mem.mem_internal.code_mem[97][4]$_SDFFCE_PN0P__3372  (.L_HI(net3372));
 sg13g2_tiehi \mem.mem_internal.code_mem[97][5]$_SDFFCE_PN0P__3373  (.L_HI(net3373));
 sg13g2_tiehi \mem.mem_internal.code_mem[97][6]$_SDFFCE_PN0P__3374  (.L_HI(net3374));
 sg13g2_tiehi \mem.mem_internal.code_mem[97][7]$_SDFFCE_PN0P__3375  (.L_HI(net3375));
 sg13g2_tiehi \mem.mem_internal.code_mem[98][0]$_SDFFCE_PN0P__3376  (.L_HI(net3376));
 sg13g2_tiehi \mem.mem_internal.code_mem[98][1]$_SDFFCE_PN0P__3377  (.L_HI(net3377));
 sg13g2_tiehi \mem.mem_internal.code_mem[98][2]$_SDFFCE_PN0P__3378  (.L_HI(net3378));
 sg13g2_tiehi \mem.mem_internal.code_mem[98][3]$_SDFFCE_PN0P__3379  (.L_HI(net3379));
 sg13g2_tiehi \mem.mem_internal.code_mem[98][4]$_SDFFCE_PN0P__3380  (.L_HI(net3380));
 sg13g2_tiehi \mem.mem_internal.code_mem[98][5]$_SDFFCE_PN0P__3381  (.L_HI(net3381));
 sg13g2_tiehi \mem.mem_internal.code_mem[98][6]$_SDFFCE_PN0P__3382  (.L_HI(net3382));
 sg13g2_tiehi \mem.mem_internal.code_mem[98][7]$_SDFFCE_PN0P__3383  (.L_HI(net3383));
 sg13g2_tiehi \mem.mem_internal.code_mem[99][0]$_SDFFCE_PN0P__3384  (.L_HI(net3384));
 sg13g2_tiehi \mem.mem_internal.code_mem[99][1]$_SDFFCE_PN0P__3385  (.L_HI(net3385));
 sg13g2_tiehi \mem.mem_internal.code_mem[99][2]$_SDFFCE_PN0P__3386  (.L_HI(net3386));
 sg13g2_tiehi \mem.mem_internal.code_mem[99][3]$_SDFFCE_PN0P__3387  (.L_HI(net3387));
 sg13g2_tiehi \mem.mem_internal.code_mem[99][4]$_SDFFCE_PN0P__3388  (.L_HI(net3388));
 sg13g2_tiehi \mem.mem_internal.code_mem[99][5]$_SDFFCE_PN0P__3389  (.L_HI(net3389));
 sg13g2_tiehi \mem.mem_internal.code_mem[99][6]$_SDFFCE_PN0P__3390  (.L_HI(net3390));
 sg13g2_tiehi \mem.mem_internal.code_mem[99][7]$_SDFFCE_PN0P__3391  (.L_HI(net3391));
 sg13g2_tiehi \mem.mem_internal.code_mem[9][0]$_SDFFCE_PN0P__3392  (.L_HI(net3392));
 sg13g2_tiehi \mem.mem_internal.code_mem[9][1]$_SDFFCE_PN0P__3393  (.L_HI(net3393));
 sg13g2_tiehi \mem.mem_internal.code_mem[9][2]$_SDFFCE_PN0P__3394  (.L_HI(net3394));
 sg13g2_tiehi \mem.mem_internal.code_mem[9][3]$_SDFFCE_PN0P__3395  (.L_HI(net3395));
 sg13g2_tiehi \mem.mem_internal.code_mem[9][4]$_SDFFCE_PN0P__3396  (.L_HI(net3396));
 sg13g2_tiehi \mem.mem_internal.code_mem[9][5]$_SDFFCE_PN0P__3397  (.L_HI(net3397));
 sg13g2_tiehi \mem.mem_internal.code_mem[9][6]$_SDFFCE_PN0P__3398  (.L_HI(net3398));
 sg13g2_tiehi \mem.mem_internal.code_mem[9][7]$_SDFFCE_PN0P__3399  (.L_HI(net3399));
 sg13g2_tiehi \mem.mem_internal.cycles[0]$_SDFFE_PN0P__3400  (.L_HI(net3400));
 sg13g2_tiehi \mem.mem_internal.cycles[1]$_SDFFE_PN0P__3401  (.L_HI(net3401));
 sg13g2_tiehi \mem.mem_internal.data_mem[0][0]$_SDFFCE_PN0P__3402  (.L_HI(net3402));
 sg13g2_tiehi \mem.mem_internal.data_mem[0][1]$_SDFFCE_PN0P__3403  (.L_HI(net3403));
 sg13g2_tiehi \mem.mem_internal.data_mem[0][2]$_SDFFCE_PN0P__3404  (.L_HI(net3404));
 sg13g2_tiehi \mem.mem_internal.data_mem[0][3]$_SDFFCE_PN0P__3405  (.L_HI(net3405));
 sg13g2_tiehi \mem.mem_internal.data_mem[0][4]$_SDFFCE_PN0P__3406  (.L_HI(net3406));
 sg13g2_tiehi \mem.mem_internal.data_mem[0][5]$_SDFFCE_PN0P__3407  (.L_HI(net3407));
 sg13g2_tiehi \mem.mem_internal.data_mem[0][6]$_SDFFCE_PN0P__3408  (.L_HI(net3408));
 sg13g2_tiehi \mem.mem_internal.data_mem[0][7]$_SDFFCE_PN0P__3409  (.L_HI(net3409));
 sg13g2_tiehi \mem.mem_internal.data_mem[10][0]$_SDFFCE_PN0P__3410  (.L_HI(net3410));
 sg13g2_tiehi \mem.mem_internal.data_mem[10][1]$_SDFFCE_PN0P__3411  (.L_HI(net3411));
 sg13g2_tiehi \mem.mem_internal.data_mem[10][2]$_SDFFCE_PN0P__3412  (.L_HI(net3412));
 sg13g2_tiehi \mem.mem_internal.data_mem[10][3]$_SDFFCE_PN0P__3413  (.L_HI(net3413));
 sg13g2_tiehi \mem.mem_internal.data_mem[10][4]$_SDFFCE_PN0P__3414  (.L_HI(net3414));
 sg13g2_tiehi \mem.mem_internal.data_mem[10][5]$_SDFFCE_PN0P__3415  (.L_HI(net3415));
 sg13g2_tiehi \mem.mem_internal.data_mem[10][6]$_SDFFCE_PN0P__3416  (.L_HI(net3416));
 sg13g2_tiehi \mem.mem_internal.data_mem[10][7]$_SDFFCE_PN0P__3417  (.L_HI(net3417));
 sg13g2_tiehi \mem.mem_internal.data_mem[11][0]$_SDFFCE_PN0P__3418  (.L_HI(net3418));
 sg13g2_tiehi \mem.mem_internal.data_mem[11][1]$_SDFFCE_PN0P__3419  (.L_HI(net3419));
 sg13g2_tiehi \mem.mem_internal.data_mem[11][2]$_SDFFCE_PN0P__3420  (.L_HI(net3420));
 sg13g2_tiehi \mem.mem_internal.data_mem[11][3]$_SDFFCE_PN0P__3421  (.L_HI(net3421));
 sg13g2_tiehi \mem.mem_internal.data_mem[11][4]$_SDFFCE_PN0P__3422  (.L_HI(net3422));
 sg13g2_tiehi \mem.mem_internal.data_mem[11][5]$_SDFFCE_PN0P__3423  (.L_HI(net3423));
 sg13g2_tiehi \mem.mem_internal.data_mem[11][6]$_SDFFCE_PN0P__3424  (.L_HI(net3424));
 sg13g2_tiehi \mem.mem_internal.data_mem[11][7]$_SDFFCE_PN0P__3425  (.L_HI(net3425));
 sg13g2_tiehi \mem.mem_internal.data_mem[12][0]$_SDFFCE_PN0P__3426  (.L_HI(net3426));
 sg13g2_tiehi \mem.mem_internal.data_mem[12][1]$_SDFFCE_PN0P__3427  (.L_HI(net3427));
 sg13g2_tiehi \mem.mem_internal.data_mem[12][2]$_SDFFCE_PN0P__3428  (.L_HI(net3428));
 sg13g2_tiehi \mem.mem_internal.data_mem[12][3]$_SDFFCE_PN0P__3429  (.L_HI(net3429));
 sg13g2_tiehi \mem.mem_internal.data_mem[12][4]$_SDFFCE_PN0P__3430  (.L_HI(net3430));
 sg13g2_tiehi \mem.mem_internal.data_mem[12][5]$_SDFFCE_PN0P__3431  (.L_HI(net3431));
 sg13g2_tiehi \mem.mem_internal.data_mem[12][6]$_SDFFCE_PN0P__3432  (.L_HI(net3432));
 sg13g2_tiehi \mem.mem_internal.data_mem[12][7]$_SDFFCE_PN0P__3433  (.L_HI(net3433));
 sg13g2_tiehi \mem.mem_internal.data_mem[13][0]$_SDFFCE_PN0P__3434  (.L_HI(net3434));
 sg13g2_tiehi \mem.mem_internal.data_mem[13][1]$_SDFFCE_PN0P__3435  (.L_HI(net3435));
 sg13g2_tiehi \mem.mem_internal.data_mem[13][2]$_SDFFCE_PN0P__3436  (.L_HI(net3436));
 sg13g2_tiehi \mem.mem_internal.data_mem[13][3]$_SDFFCE_PN0P__3437  (.L_HI(net3437));
 sg13g2_tiehi \mem.mem_internal.data_mem[13][4]$_SDFFCE_PN0P__3438  (.L_HI(net3438));
 sg13g2_tiehi \mem.mem_internal.data_mem[13][5]$_SDFFCE_PN0P__3439  (.L_HI(net3439));
 sg13g2_tiehi \mem.mem_internal.data_mem[13][6]$_SDFFCE_PN0P__3440  (.L_HI(net3440));
 sg13g2_tiehi \mem.mem_internal.data_mem[13][7]$_SDFFCE_PN0P__3441  (.L_HI(net3441));
 sg13g2_tiehi \mem.mem_internal.data_mem[14][0]$_SDFFCE_PN0P__3442  (.L_HI(net3442));
 sg13g2_tiehi \mem.mem_internal.data_mem[14][1]$_SDFFCE_PN0P__3443  (.L_HI(net3443));
 sg13g2_tiehi \mem.mem_internal.data_mem[14][2]$_SDFFCE_PN0P__3444  (.L_HI(net3444));
 sg13g2_tiehi \mem.mem_internal.data_mem[14][3]$_SDFFCE_PN0P__3445  (.L_HI(net3445));
 sg13g2_tiehi \mem.mem_internal.data_mem[14][4]$_SDFFCE_PN0P__3446  (.L_HI(net3446));
 sg13g2_tiehi \mem.mem_internal.data_mem[14][5]$_SDFFCE_PN0P__3447  (.L_HI(net3447));
 sg13g2_tiehi \mem.mem_internal.data_mem[14][6]$_SDFFCE_PN0P__3448  (.L_HI(net3448));
 sg13g2_tiehi \mem.mem_internal.data_mem[14][7]$_SDFFCE_PN0P__3449  (.L_HI(net3449));
 sg13g2_tiehi \mem.mem_internal.data_mem[15][0]$_SDFFCE_PN0P__3450  (.L_HI(net3450));
 sg13g2_tiehi \mem.mem_internal.data_mem[15][1]$_SDFFCE_PN0P__3451  (.L_HI(net3451));
 sg13g2_tiehi \mem.mem_internal.data_mem[15][2]$_SDFFCE_PN0P__3452  (.L_HI(net3452));
 sg13g2_tiehi \mem.mem_internal.data_mem[15][3]$_SDFFCE_PN0P__3453  (.L_HI(net3453));
 sg13g2_tiehi \mem.mem_internal.data_mem[15][4]$_SDFFCE_PN0P__3454  (.L_HI(net3454));
 sg13g2_tiehi \mem.mem_internal.data_mem[15][5]$_SDFFCE_PN0P__3455  (.L_HI(net3455));
 sg13g2_tiehi \mem.mem_internal.data_mem[15][6]$_SDFFCE_PN0P__3456  (.L_HI(net3456));
 sg13g2_tiehi \mem.mem_internal.data_mem[15][7]$_SDFFCE_PN0P__3457  (.L_HI(net3457));
 sg13g2_tiehi \mem.mem_internal.data_mem[16][0]$_SDFFCE_PN0P__3458  (.L_HI(net3458));
 sg13g2_tiehi \mem.mem_internal.data_mem[16][1]$_SDFFCE_PN0P__3459  (.L_HI(net3459));
 sg13g2_tiehi \mem.mem_internal.data_mem[16][2]$_SDFFCE_PN0P__3460  (.L_HI(net3460));
 sg13g2_tiehi \mem.mem_internal.data_mem[16][3]$_SDFFCE_PN0P__3461  (.L_HI(net3461));
 sg13g2_tiehi \mem.mem_internal.data_mem[16][4]$_SDFFCE_PN0P__3462  (.L_HI(net3462));
 sg13g2_tiehi \mem.mem_internal.data_mem[16][5]$_SDFFCE_PN0P__3463  (.L_HI(net3463));
 sg13g2_tiehi \mem.mem_internal.data_mem[16][6]$_SDFFCE_PN0P__3464  (.L_HI(net3464));
 sg13g2_tiehi \mem.mem_internal.data_mem[16][7]$_SDFFCE_PN0P__3465  (.L_HI(net3465));
 sg13g2_tiehi \mem.mem_internal.data_mem[17][0]$_SDFFCE_PN0P__3466  (.L_HI(net3466));
 sg13g2_tiehi \mem.mem_internal.data_mem[17][1]$_SDFFCE_PN0P__3467  (.L_HI(net3467));
 sg13g2_tiehi \mem.mem_internal.data_mem[17][2]$_SDFFCE_PN0P__3468  (.L_HI(net3468));
 sg13g2_tiehi \mem.mem_internal.data_mem[17][3]$_SDFFCE_PN0P__3469  (.L_HI(net3469));
 sg13g2_tiehi \mem.mem_internal.data_mem[17][4]$_SDFFCE_PN0P__3470  (.L_HI(net3470));
 sg13g2_tiehi \mem.mem_internal.data_mem[17][5]$_SDFFCE_PN0P__3471  (.L_HI(net3471));
 sg13g2_tiehi \mem.mem_internal.data_mem[17][6]$_SDFFCE_PN0P__3472  (.L_HI(net3472));
 sg13g2_tiehi \mem.mem_internal.data_mem[17][7]$_SDFFCE_PN0P__3473  (.L_HI(net3473));
 sg13g2_tiehi \mem.mem_internal.data_mem[18][0]$_SDFFCE_PN0P__3474  (.L_HI(net3474));
 sg13g2_tiehi \mem.mem_internal.data_mem[18][1]$_SDFFCE_PN0P__3475  (.L_HI(net3475));
 sg13g2_tiehi \mem.mem_internal.data_mem[18][2]$_SDFFCE_PN0P__3476  (.L_HI(net3476));
 sg13g2_tiehi \mem.mem_internal.data_mem[18][3]$_SDFFCE_PN0P__3477  (.L_HI(net3477));
 sg13g2_tiehi \mem.mem_internal.data_mem[18][4]$_SDFFCE_PN0P__3478  (.L_HI(net3478));
 sg13g2_tiehi \mem.mem_internal.data_mem[18][5]$_SDFFCE_PN0P__3479  (.L_HI(net3479));
 sg13g2_tiehi \mem.mem_internal.data_mem[18][6]$_SDFFCE_PN0P__3480  (.L_HI(net3480));
 sg13g2_tiehi \mem.mem_internal.data_mem[18][7]$_SDFFCE_PN0P__3481  (.L_HI(net3481));
 sg13g2_tiehi \mem.mem_internal.data_mem[19][0]$_SDFFCE_PN0P__3482  (.L_HI(net3482));
 sg13g2_tiehi \mem.mem_internal.data_mem[19][1]$_SDFFCE_PN0P__3483  (.L_HI(net3483));
 sg13g2_tiehi \mem.mem_internal.data_mem[19][2]$_SDFFCE_PN0P__3484  (.L_HI(net3484));
 sg13g2_tiehi \mem.mem_internal.data_mem[19][3]$_SDFFCE_PN0P__3485  (.L_HI(net3485));
 sg13g2_tiehi \mem.mem_internal.data_mem[19][4]$_SDFFCE_PN0P__3486  (.L_HI(net3486));
 sg13g2_tiehi \mem.mem_internal.data_mem[19][5]$_SDFFCE_PN0P__3487  (.L_HI(net3487));
 sg13g2_tiehi \mem.mem_internal.data_mem[19][6]$_SDFFCE_PN0P__3488  (.L_HI(net3488));
 sg13g2_tiehi \mem.mem_internal.data_mem[19][7]$_SDFFCE_PN0P__3489  (.L_HI(net3489));
 sg13g2_tiehi \mem.mem_internal.data_mem[1][0]$_SDFFCE_PN0P__3490  (.L_HI(net3490));
 sg13g2_tiehi \mem.mem_internal.data_mem[1][1]$_SDFFCE_PN0P__3491  (.L_HI(net3491));
 sg13g2_tiehi \mem.mem_internal.data_mem[1][2]$_SDFFCE_PN0P__3492  (.L_HI(net3492));
 sg13g2_tiehi \mem.mem_internal.data_mem[1][3]$_SDFFCE_PN0P__3493  (.L_HI(net3493));
 sg13g2_tiehi \mem.mem_internal.data_mem[1][4]$_SDFFCE_PN0P__3494  (.L_HI(net3494));
 sg13g2_tiehi \mem.mem_internal.data_mem[1][5]$_SDFFCE_PN0P__3495  (.L_HI(net3495));
 sg13g2_tiehi \mem.mem_internal.data_mem[1][6]$_SDFFCE_PN0P__3496  (.L_HI(net3496));
 sg13g2_tiehi \mem.mem_internal.data_mem[1][7]$_SDFFCE_PN0P__3497  (.L_HI(net3497));
 sg13g2_tiehi \mem.mem_internal.data_mem[20][0]$_SDFFCE_PN0P__3498  (.L_HI(net3498));
 sg13g2_tiehi \mem.mem_internal.data_mem[20][1]$_SDFFCE_PN0P__3499  (.L_HI(net3499));
 sg13g2_tiehi \mem.mem_internal.data_mem[20][2]$_SDFFCE_PN0P__3500  (.L_HI(net3500));
 sg13g2_tiehi \mem.mem_internal.data_mem[20][3]$_SDFFCE_PN0P__3501  (.L_HI(net3501));
 sg13g2_tiehi \mem.mem_internal.data_mem[20][4]$_SDFFCE_PN0P__3502  (.L_HI(net3502));
 sg13g2_tiehi \mem.mem_internal.data_mem[20][5]$_SDFFCE_PN0P__3503  (.L_HI(net3503));
 sg13g2_tiehi \mem.mem_internal.data_mem[20][6]$_SDFFCE_PN0P__3504  (.L_HI(net3504));
 sg13g2_tiehi \mem.mem_internal.data_mem[20][7]$_SDFFCE_PN0P__3505  (.L_HI(net3505));
 sg13g2_tiehi \mem.mem_internal.data_mem[21][0]$_SDFFCE_PN0P__3506  (.L_HI(net3506));
 sg13g2_tiehi \mem.mem_internal.data_mem[21][1]$_SDFFCE_PN0P__3507  (.L_HI(net3507));
 sg13g2_tiehi \mem.mem_internal.data_mem[21][2]$_SDFFCE_PN0P__3508  (.L_HI(net3508));
 sg13g2_tiehi \mem.mem_internal.data_mem[21][3]$_SDFFCE_PN0P__3509  (.L_HI(net3509));
 sg13g2_tiehi \mem.mem_internal.data_mem[21][4]$_SDFFCE_PN0P__3510  (.L_HI(net3510));
 sg13g2_tiehi \mem.mem_internal.data_mem[21][5]$_SDFFCE_PN0P__3511  (.L_HI(net3511));
 sg13g2_tiehi \mem.mem_internal.data_mem[21][6]$_SDFFCE_PN0P__3512  (.L_HI(net3512));
 sg13g2_tiehi \mem.mem_internal.data_mem[21][7]$_SDFFCE_PN0P__3513  (.L_HI(net3513));
 sg13g2_tiehi \mem.mem_internal.data_mem[22][0]$_SDFFCE_PN0P__3514  (.L_HI(net3514));
 sg13g2_tiehi \mem.mem_internal.data_mem[22][1]$_SDFFCE_PN0P__3515  (.L_HI(net3515));
 sg13g2_tiehi \mem.mem_internal.data_mem[22][2]$_SDFFCE_PN0P__3516  (.L_HI(net3516));
 sg13g2_tiehi \mem.mem_internal.data_mem[22][3]$_SDFFCE_PN0P__3517  (.L_HI(net3517));
 sg13g2_tiehi \mem.mem_internal.data_mem[22][4]$_SDFFCE_PN0P__3518  (.L_HI(net3518));
 sg13g2_tiehi \mem.mem_internal.data_mem[22][5]$_SDFFCE_PN0P__3519  (.L_HI(net3519));
 sg13g2_tiehi \mem.mem_internal.data_mem[22][6]$_SDFFCE_PN0P__3520  (.L_HI(net3520));
 sg13g2_tiehi \mem.mem_internal.data_mem[22][7]$_SDFFCE_PN0P__3521  (.L_HI(net3521));
 sg13g2_tiehi \mem.mem_internal.data_mem[23][0]$_SDFFCE_PN0P__3522  (.L_HI(net3522));
 sg13g2_tiehi \mem.mem_internal.data_mem[23][1]$_SDFFCE_PN0P__3523  (.L_HI(net3523));
 sg13g2_tiehi \mem.mem_internal.data_mem[23][2]$_SDFFCE_PN0P__3524  (.L_HI(net3524));
 sg13g2_tiehi \mem.mem_internal.data_mem[23][3]$_SDFFCE_PN0P__3525  (.L_HI(net3525));
 sg13g2_tiehi \mem.mem_internal.data_mem[23][4]$_SDFFCE_PN0P__3526  (.L_HI(net3526));
 sg13g2_tiehi \mem.mem_internal.data_mem[23][5]$_SDFFCE_PN0P__3527  (.L_HI(net3527));
 sg13g2_tiehi \mem.mem_internal.data_mem[23][6]$_SDFFCE_PN0P__3528  (.L_HI(net3528));
 sg13g2_tiehi \mem.mem_internal.data_mem[23][7]$_SDFFCE_PN0P__3529  (.L_HI(net3529));
 sg13g2_tiehi \mem.mem_internal.data_mem[24][0]$_SDFFCE_PN0P__3530  (.L_HI(net3530));
 sg13g2_tiehi \mem.mem_internal.data_mem[24][1]$_SDFFCE_PN0P__3531  (.L_HI(net3531));
 sg13g2_tiehi \mem.mem_internal.data_mem[24][2]$_SDFFCE_PN0P__3532  (.L_HI(net3532));
 sg13g2_tiehi \mem.mem_internal.data_mem[24][3]$_SDFFCE_PN0P__3533  (.L_HI(net3533));
 sg13g2_tiehi \mem.mem_internal.data_mem[24][4]$_SDFFCE_PN0P__3534  (.L_HI(net3534));
 sg13g2_tiehi \mem.mem_internal.data_mem[24][5]$_SDFFCE_PN0P__3535  (.L_HI(net3535));
 sg13g2_tiehi \mem.mem_internal.data_mem[24][6]$_SDFFCE_PN0P__3536  (.L_HI(net3536));
 sg13g2_tiehi \mem.mem_internal.data_mem[24][7]$_SDFFCE_PN0P__3537  (.L_HI(net3537));
 sg13g2_tiehi \mem.mem_internal.data_mem[25][0]$_SDFFCE_PN0P__3538  (.L_HI(net3538));
 sg13g2_tiehi \mem.mem_internal.data_mem[25][1]$_SDFFCE_PN0P__3539  (.L_HI(net3539));
 sg13g2_tiehi \mem.mem_internal.data_mem[25][2]$_SDFFCE_PN0P__3540  (.L_HI(net3540));
 sg13g2_tiehi \mem.mem_internal.data_mem[25][3]$_SDFFCE_PN0P__3541  (.L_HI(net3541));
 sg13g2_tiehi \mem.mem_internal.data_mem[25][4]$_SDFFCE_PN0P__3542  (.L_HI(net3542));
 sg13g2_tiehi \mem.mem_internal.data_mem[25][5]$_SDFFCE_PN0P__3543  (.L_HI(net3543));
 sg13g2_tiehi \mem.mem_internal.data_mem[25][6]$_SDFFCE_PN0P__3544  (.L_HI(net3544));
 sg13g2_tiehi \mem.mem_internal.data_mem[25][7]$_SDFFCE_PN0P__3545  (.L_HI(net3545));
 sg13g2_tiehi \mem.mem_internal.data_mem[26][0]$_SDFFCE_PN0P__3546  (.L_HI(net3546));
 sg13g2_tiehi \mem.mem_internal.data_mem[26][1]$_SDFFCE_PN0P__3547  (.L_HI(net3547));
 sg13g2_tiehi \mem.mem_internal.data_mem[26][2]$_SDFFCE_PN0P__3548  (.L_HI(net3548));
 sg13g2_tiehi \mem.mem_internal.data_mem[26][3]$_SDFFCE_PN0P__3549  (.L_HI(net3549));
 sg13g2_tiehi \mem.mem_internal.data_mem[26][4]$_SDFFCE_PN0P__3550  (.L_HI(net3550));
 sg13g2_tiehi \mem.mem_internal.data_mem[26][5]$_SDFFCE_PN0P__3551  (.L_HI(net3551));
 sg13g2_tiehi \mem.mem_internal.data_mem[26][6]$_SDFFCE_PN0P__3552  (.L_HI(net3552));
 sg13g2_tiehi \mem.mem_internal.data_mem[26][7]$_SDFFCE_PN0P__3553  (.L_HI(net3553));
 sg13g2_tiehi \mem.mem_internal.data_mem[27][0]$_SDFFCE_PN0P__3554  (.L_HI(net3554));
 sg13g2_tiehi \mem.mem_internal.data_mem[27][1]$_SDFFCE_PN0P__3555  (.L_HI(net3555));
 sg13g2_tiehi \mem.mem_internal.data_mem[27][2]$_SDFFCE_PN0P__3556  (.L_HI(net3556));
 sg13g2_tiehi \mem.mem_internal.data_mem[27][3]$_SDFFCE_PN0P__3557  (.L_HI(net3557));
 sg13g2_tiehi \mem.mem_internal.data_mem[27][4]$_SDFFCE_PN0P__3558  (.L_HI(net3558));
 sg13g2_tiehi \mem.mem_internal.data_mem[27][5]$_SDFFCE_PN0P__3559  (.L_HI(net3559));
 sg13g2_tiehi \mem.mem_internal.data_mem[27][6]$_SDFFCE_PN0P__3560  (.L_HI(net3560));
 sg13g2_tiehi \mem.mem_internal.data_mem[27][7]$_SDFFCE_PN0P__3561  (.L_HI(net3561));
 sg13g2_tiehi \mem.mem_internal.data_mem[28][0]$_SDFFCE_PN0P__3562  (.L_HI(net3562));
 sg13g2_tiehi \mem.mem_internal.data_mem[28][1]$_SDFFCE_PN0P__3563  (.L_HI(net3563));
 sg13g2_tiehi \mem.mem_internal.data_mem[28][2]$_SDFFCE_PN0P__3564  (.L_HI(net3564));
 sg13g2_tiehi \mem.mem_internal.data_mem[28][3]$_SDFFCE_PN0P__3565  (.L_HI(net3565));
 sg13g2_tiehi \mem.mem_internal.data_mem[28][4]$_SDFFCE_PN0P__3566  (.L_HI(net3566));
 sg13g2_tiehi \mem.mem_internal.data_mem[28][5]$_SDFFCE_PN0P__3567  (.L_HI(net3567));
 sg13g2_tiehi \mem.mem_internal.data_mem[28][6]$_SDFFCE_PN0P__3568  (.L_HI(net3568));
 sg13g2_tiehi \mem.mem_internal.data_mem[28][7]$_SDFFCE_PN0P__3569  (.L_HI(net3569));
 sg13g2_tiehi \mem.mem_internal.data_mem[29][0]$_SDFFCE_PN0P__3570  (.L_HI(net3570));
 sg13g2_tiehi \mem.mem_internal.data_mem[29][1]$_SDFFCE_PN0P__3571  (.L_HI(net3571));
 sg13g2_tiehi \mem.mem_internal.data_mem[29][2]$_SDFFCE_PN0P__3572  (.L_HI(net3572));
 sg13g2_tiehi \mem.mem_internal.data_mem[29][3]$_SDFFCE_PN0P__3573  (.L_HI(net3573));
 sg13g2_tiehi \mem.mem_internal.data_mem[29][4]$_SDFFCE_PN0P__3574  (.L_HI(net3574));
 sg13g2_tiehi \mem.mem_internal.data_mem[29][5]$_SDFFCE_PN0P__3575  (.L_HI(net3575));
 sg13g2_tiehi \mem.mem_internal.data_mem[29][6]$_SDFFCE_PN0P__3576  (.L_HI(net3576));
 sg13g2_tiehi \mem.mem_internal.data_mem[29][7]$_SDFFCE_PN0P__3577  (.L_HI(net3577));
 sg13g2_tiehi \mem.mem_internal.data_mem[2][0]$_SDFFCE_PN0P__3578  (.L_HI(net3578));
 sg13g2_tiehi \mem.mem_internal.data_mem[2][1]$_SDFFCE_PN0P__3579  (.L_HI(net3579));
 sg13g2_tiehi \mem.mem_internal.data_mem[2][2]$_SDFFCE_PN0P__3580  (.L_HI(net3580));
 sg13g2_tiehi \mem.mem_internal.data_mem[2][3]$_SDFFCE_PN0P__3581  (.L_HI(net3581));
 sg13g2_tiehi \mem.mem_internal.data_mem[2][4]$_SDFFCE_PN0P__3582  (.L_HI(net3582));
 sg13g2_tiehi \mem.mem_internal.data_mem[2][5]$_SDFFCE_PN0P__3583  (.L_HI(net3583));
 sg13g2_tiehi \mem.mem_internal.data_mem[2][6]$_SDFFCE_PN0P__3584  (.L_HI(net3584));
 sg13g2_tiehi \mem.mem_internal.data_mem[2][7]$_SDFFCE_PN0P__3585  (.L_HI(net3585));
 sg13g2_tiehi \mem.mem_internal.data_mem[30][0]$_SDFFCE_PN0P__3586  (.L_HI(net3586));
 sg13g2_tiehi \mem.mem_internal.data_mem[30][1]$_SDFFCE_PN0P__3587  (.L_HI(net3587));
 sg13g2_tiehi \mem.mem_internal.data_mem[30][2]$_SDFFCE_PN0P__3588  (.L_HI(net3588));
 sg13g2_tiehi \mem.mem_internal.data_mem[30][3]$_SDFFCE_PN0P__3589  (.L_HI(net3589));
 sg13g2_tiehi \mem.mem_internal.data_mem[30][4]$_SDFFCE_PN0P__3590  (.L_HI(net3590));
 sg13g2_tiehi \mem.mem_internal.data_mem[30][5]$_SDFFCE_PN0P__3591  (.L_HI(net3591));
 sg13g2_tiehi \mem.mem_internal.data_mem[30][6]$_SDFFCE_PN0P__3592  (.L_HI(net3592));
 sg13g2_tiehi \mem.mem_internal.data_mem[30][7]$_SDFFCE_PN0P__3593  (.L_HI(net3593));
 sg13g2_tiehi \mem.mem_internal.data_mem[31][0]$_SDFFCE_PN0P__3594  (.L_HI(net3594));
 sg13g2_tiehi \mem.mem_internal.data_mem[31][1]$_SDFFCE_PN0P__3595  (.L_HI(net3595));
 sg13g2_tiehi \mem.mem_internal.data_mem[31][2]$_SDFFCE_PN0P__3596  (.L_HI(net3596));
 sg13g2_tiehi \mem.mem_internal.data_mem[31][3]$_SDFFCE_PN0P__3597  (.L_HI(net3597));
 sg13g2_tiehi \mem.mem_internal.data_mem[31][4]$_SDFFCE_PN0P__3598  (.L_HI(net3598));
 sg13g2_tiehi \mem.mem_internal.data_mem[31][5]$_SDFFCE_PN0P__3599  (.L_HI(net3599));
 sg13g2_tiehi \mem.mem_internal.data_mem[31][6]$_SDFFCE_PN0P__3600  (.L_HI(net3600));
 sg13g2_tiehi \mem.mem_internal.data_mem[31][7]$_SDFFCE_PN0P__3601  (.L_HI(net3601));
 sg13g2_tiehi \mem.mem_internal.data_mem[3][0]$_SDFFCE_PN0P__3602  (.L_HI(net3602));
 sg13g2_tiehi \mem.mem_internal.data_mem[3][1]$_SDFFCE_PN0P__3603  (.L_HI(net3603));
 sg13g2_tiehi \mem.mem_internal.data_mem[3][2]$_SDFFCE_PN0P__3604  (.L_HI(net3604));
 sg13g2_tiehi \mem.mem_internal.data_mem[3][3]$_SDFFCE_PN0P__3605  (.L_HI(net3605));
 sg13g2_tiehi \mem.mem_internal.data_mem[3][4]$_SDFFCE_PN0P__3606  (.L_HI(net3606));
 sg13g2_tiehi \mem.mem_internal.data_mem[3][5]$_SDFFCE_PN0P__3607  (.L_HI(net3607));
 sg13g2_tiehi \mem.mem_internal.data_mem[3][6]$_SDFFCE_PN0P__3608  (.L_HI(net3608));
 sg13g2_tiehi \mem.mem_internal.data_mem[3][7]$_SDFFCE_PN0P__3609  (.L_HI(net3609));
 sg13g2_tiehi \mem.mem_internal.data_mem[4][0]$_SDFFCE_PN0P__3610  (.L_HI(net3610));
 sg13g2_tiehi \mem.mem_internal.data_mem[4][1]$_SDFFCE_PN0P__3611  (.L_HI(net3611));
 sg13g2_tiehi \mem.mem_internal.data_mem[4][2]$_SDFFCE_PN0P__3612  (.L_HI(net3612));
 sg13g2_tiehi \mem.mem_internal.data_mem[4][3]$_SDFFCE_PN0P__3613  (.L_HI(net3613));
 sg13g2_tiehi \mem.mem_internal.data_mem[4][4]$_SDFFCE_PN0P__3614  (.L_HI(net3614));
 sg13g2_tiehi \mem.mem_internal.data_mem[4][5]$_SDFFCE_PN0P__3615  (.L_HI(net3615));
 sg13g2_tiehi \mem.mem_internal.data_mem[4][6]$_SDFFCE_PN0P__3616  (.L_HI(net3616));
 sg13g2_tiehi \mem.mem_internal.data_mem[4][7]$_SDFFCE_PN0P__3617  (.L_HI(net3617));
 sg13g2_tiehi \mem.mem_internal.data_mem[5][0]$_SDFFCE_PN0P__3618  (.L_HI(net3618));
 sg13g2_tiehi \mem.mem_internal.data_mem[5][1]$_SDFFCE_PN0P__3619  (.L_HI(net3619));
 sg13g2_tiehi \mem.mem_internal.data_mem[5][2]$_SDFFCE_PN0P__3620  (.L_HI(net3620));
 sg13g2_tiehi \mem.mem_internal.data_mem[5][3]$_SDFFCE_PN0P__3621  (.L_HI(net3621));
 sg13g2_tiehi \mem.mem_internal.data_mem[5][4]$_SDFFCE_PN0P__3622  (.L_HI(net3622));
 sg13g2_tiehi \mem.mem_internal.data_mem[5][5]$_SDFFCE_PN0P__3623  (.L_HI(net3623));
 sg13g2_tiehi \mem.mem_internal.data_mem[5][6]$_SDFFCE_PN0P__3624  (.L_HI(net3624));
 sg13g2_tiehi \mem.mem_internal.data_mem[5][7]$_SDFFCE_PN0P__3625  (.L_HI(net3625));
 sg13g2_tiehi \mem.mem_internal.data_mem[6][0]$_SDFFCE_PN0P__3626  (.L_HI(net3626));
 sg13g2_tiehi \mem.mem_internal.data_mem[6][1]$_SDFFCE_PN0P__3627  (.L_HI(net3627));
 sg13g2_tiehi \mem.mem_internal.data_mem[6][2]$_SDFFCE_PN0P__3628  (.L_HI(net3628));
 sg13g2_tiehi \mem.mem_internal.data_mem[6][3]$_SDFFCE_PN0P__3629  (.L_HI(net3629));
 sg13g2_tiehi \mem.mem_internal.data_mem[6][4]$_SDFFCE_PN0P__3630  (.L_HI(net3630));
 sg13g2_tiehi \mem.mem_internal.data_mem[6][5]$_SDFFCE_PN0P__3631  (.L_HI(net3631));
 sg13g2_tiehi \mem.mem_internal.data_mem[6][6]$_SDFFCE_PN0P__3632  (.L_HI(net3632));
 sg13g2_tiehi \mem.mem_internal.data_mem[6][7]$_SDFFCE_PN0P__3633  (.L_HI(net3633));
 sg13g2_tiehi \mem.mem_internal.data_mem[7][0]$_SDFFCE_PN0P__3634  (.L_HI(net3634));
 sg13g2_tiehi \mem.mem_internal.data_mem[7][1]$_SDFFCE_PN0P__3635  (.L_HI(net3635));
 sg13g2_tiehi \mem.mem_internal.data_mem[7][2]$_SDFFCE_PN0P__3636  (.L_HI(net3636));
 sg13g2_tiehi \mem.mem_internal.data_mem[7][3]$_SDFFCE_PN0P__3637  (.L_HI(net3637));
 sg13g2_tiehi \mem.mem_internal.data_mem[7][4]$_SDFFCE_PN0P__3638  (.L_HI(net3638));
 sg13g2_tiehi \mem.mem_internal.data_mem[7][5]$_SDFFCE_PN0P__3639  (.L_HI(net3639));
 sg13g2_tiehi \mem.mem_internal.data_mem[7][6]$_SDFFCE_PN0P__3640  (.L_HI(net3640));
 sg13g2_tiehi \mem.mem_internal.data_mem[7][7]$_SDFFCE_PN0P__3641  (.L_HI(net3641));
 sg13g2_tiehi \mem.mem_internal.data_mem[8][0]$_SDFFCE_PN0P__3642  (.L_HI(net3642));
 sg13g2_tiehi \mem.mem_internal.data_mem[8][1]$_SDFFCE_PN0P__3643  (.L_HI(net3643));
 sg13g2_tiehi \mem.mem_internal.data_mem[8][2]$_SDFFCE_PN0P__3644  (.L_HI(net3644));
 sg13g2_tiehi \mem.mem_internal.data_mem[8][3]$_SDFFCE_PN0P__3645  (.L_HI(net3645));
 sg13g2_tiehi \mem.mem_internal.data_mem[8][4]$_SDFFCE_PN0P__3646  (.L_HI(net3646));
 sg13g2_tiehi \mem.mem_internal.data_mem[8][5]$_SDFFCE_PN0P__3647  (.L_HI(net3647));
 sg13g2_tiehi \mem.mem_internal.data_mem[8][6]$_SDFFCE_PN0P__3648  (.L_HI(net3648));
 sg13g2_tiehi \mem.mem_internal.data_mem[8][7]$_SDFFCE_PN0P__3649  (.L_HI(net3649));
 sg13g2_tiehi \mem.mem_internal.data_mem[9][0]$_SDFFCE_PN0P__3650  (.L_HI(net3650));
 sg13g2_tiehi \mem.mem_internal.data_mem[9][1]$_SDFFCE_PN0P__3651  (.L_HI(net3651));
 sg13g2_tiehi \mem.mem_internal.data_mem[9][2]$_SDFFCE_PN0P__3652  (.L_HI(net3652));
 sg13g2_tiehi \mem.mem_internal.data_mem[9][3]$_SDFFCE_PN0P__3653  (.L_HI(net3653));
 sg13g2_tiehi \mem.mem_internal.data_mem[9][4]$_SDFFCE_PN0P__3654  (.L_HI(net3654));
 sg13g2_tiehi \mem.mem_internal.data_mem[9][5]$_SDFFCE_PN0P__3655  (.L_HI(net3655));
 sg13g2_tiehi \mem.mem_internal.data_mem[9][6]$_SDFFCE_PN0P__3656  (.L_HI(net3656));
 sg13g2_tiehi \mem.mem_internal.data_mem[9][7]$_SDFFCE_PN0P__3657  (.L_HI(net3657));
 sg13g2_tiehi \mem.mem_internal.data_out[0]$_DFFE_PP__3658  (.L_HI(net3658));
 sg13g2_tiehi \mem.mem_internal.data_out[1]$_DFFE_PP__3659  (.L_HI(net3659));
 sg13g2_tiehi \mem.mem_internal.data_out[2]$_DFFE_PP__3660  (.L_HI(net3660));
 sg13g2_tiehi \mem.mem_internal.data_out[3]$_DFFE_PP__3661  (.L_HI(net3661));
 sg13g2_tiehi \mem.mem_internal.data_out[4]$_DFFE_PP__3662  (.L_HI(net3662));
 sg13g2_tiehi \mem.mem_internal.data_out[5]$_DFFE_PP__3663  (.L_HI(net3663));
 sg13g2_tiehi \mem.mem_internal.data_out[6]$_DFFE_PP__3664  (.L_HI(net3664));
 sg13g2_tiehi \mem.mem_internal.data_out[7]$_DFFE_PP__3665  (.L_HI(net3665));
 sg13g2_tiehi \mem.mem_internal.data_ready$_SDFFE_PN0P__3666  (.L_HI(net3666));
 sg13g2_tiehi \mem.mem_io.data_out[0]$_SDFFE_PN0P__3667  (.L_HI(net3667));
 sg13g2_tiehi \mem.mem_io.data_out[1]$_SDFFE_PN0P__3668  (.L_HI(net3668));
 sg13g2_tiehi \mem.mem_io.data_out[2]$_SDFFE_PN0P__3669  (.L_HI(net3669));
 sg13g2_tiehi \mem.mem_io.data_out[3]$_SDFFE_PN0P__3670  (.L_HI(net3670));
 sg13g2_tiehi \mem.mem_io.data_out[4]$_SDFFE_PN0P__3671  (.L_HI(net3671));
 sg13g2_tiehi \mem.mem_io.data_out[5]$_SDFFE_PN0P__3672  (.L_HI(net3672));
 sg13g2_tiehi \mem.mem_io.data_out[6]$_SDFFE_PN0P__3673  (.L_HI(net3673));
 sg13g2_tiehi \mem.mem_io.data_out[7]$_SDFFE_PN0P__3674  (.L_HI(net3674));
 sg13g2_tiehi \mem.mem_io.data_ready$_SDFF_PN0__3675  (.L_HI(net3675));
 sg13g2_tiehi \mem.mem_io.past_write$_SDFF_PN0__3676  (.L_HI(net3676));
 sg13g2_tiehi \mem.mem_io.porta_oe[0]$_SDFFE_PN0P__3677  (.L_HI(net3677));
 sg13g2_tiehi \mem.mem_io.porta_oe[1]$_SDFFE_PN0P__3678  (.L_HI(net3678));
 sg13g2_tiehi \mem.mem_io.porta_oe[2]$_SDFFE_PN0P__3679  (.L_HI(net3679));
 sg13g2_tiehi \mem.mem_io.porta_oe[3]$_SDFFE_PN0P__3680  (.L_HI(net3680));
 sg13g2_tiehi \mem.mem_io.porta_oe[4]$_SDFFE_PN0P__3681  (.L_HI(net3681));
 sg13g2_tiehi \mem.mem_io.porta_oe[5]$_SDFFE_PN0P__3682  (.L_HI(net3682));
 sg13g2_tiehi \mem.mem_io.porta_oe[6]$_SDFFE_PN0P__3683  (.L_HI(net3683));
 sg13g2_tiehi \mem.mem_io.porta_oe[7]$_SDFFE_PN0P__3684  (.L_HI(net3684));
 sg13g2_tiehi \mem.mem_io.porta_out[0]$_SDFFE_PN0P__3685  (.L_HI(net3685));
 sg13g2_tiehi \mem.mem_io.porta_out[1]$_SDFFE_PN0P__3686  (.L_HI(net3686));
 sg13g2_tiehi \mem.mem_io.porta_out[2]$_SDFFE_PN0P__3687  (.L_HI(net3687));
 sg13g2_tiehi \mem.mem_io.porta_out[3]$_SDFFE_PN0P__3688  (.L_HI(net3688));
 sg13g2_tiehi \mem.mem_io.porta_out[4]$_SDFFE_PN0P__3689  (.L_HI(net3689));
 sg13g2_tiehi \mem.mem_io.porta_out[5]$_SDFFE_PN0P__3690  (.L_HI(net3690));
 sg13g2_tiehi \mem.mem_io.porta_out[6]$_SDFFE_PN0P__3691  (.L_HI(net3691));
 sg13g2_tiehi \mem.mem_io.porta_out[7]$_SDFFE_PN0P__3692  (.L_HI(net3692));
 sg13g2_tiehi \mem.mem_io.portb_oe[0]$_SDFFE_PN0P__3693  (.L_HI(net3693));
 sg13g2_tiehi \mem.mem_io.portb_oe[1]$_SDFFE_PN0P__3694  (.L_HI(net3694));
 sg13g2_tiehi \mem.mem_io.portb_oe[2]$_SDFFE_PN0P__3695  (.L_HI(net3695));
 sg13g2_tiehi \mem.mem_io.portb_oe[3]$_SDFFE_PN0P__3696  (.L_HI(net3696));
 sg13g2_tiehi \mem.mem_io.portb_oe[4]$_SDFFE_PN0P__3697  (.L_HI(net3697));
 sg13g2_tiehi \mem.mem_io.portb_oe[5]$_SDFFE_PN0P__3698  (.L_HI(net3698));
 sg13g2_tiehi \mem.mem_io.portb_oe[6]$_SDFFE_PN0P__3699  (.L_HI(net3699));
 sg13g2_tiehi \mem.mem_io.portb_oe[7]$_SDFFE_PN0P__3700  (.L_HI(net3700));
 sg13g2_tiehi \mem.mem_io.portb_out[0]$_SDFFE_PN0P__3701  (.L_HI(net3701));
 sg13g2_tiehi \mem.mem_io.portb_out[1]$_SDFFE_PN0P__3702  (.L_HI(net3702));
 sg13g2_tiehi \mem.mem_io.portb_out[2]$_SDFFE_PN0P__3703  (.L_HI(net3703));
 sg13g2_tiehi \mem.mem_io.portb_out[3]$_SDFFE_PN0P__3704  (.L_HI(net3704));
 sg13g2_tiehi \mem.mem_io.portb_out[4]$_SDFFE_PN0P__3705  (.L_HI(net3705));
 sg13g2_tiehi \mem.mem_io.portb_out[5]$_SDFFE_PN0P__3706  (.L_HI(net3706));
 sg13g2_tiehi \mem.mem_io.portb_out[6]$_SDFFE_PN0P__3707  (.L_HI(net3707));
 sg13g2_tiehi \mem.mem_io.portb_out[7]$_SDFFE_PN0P__3708  (.L_HI(net3708));
 sg13g2_tiehi \mem_addr[0]$_DFFE_PP__3709  (.L_HI(net3709));
 sg13g2_tiehi \mem_addr[1]$_DFFE_PP__3710  (.L_HI(net3710));
 sg13g2_tiehi \mem_addr[2]$_DFFE_PP__3711  (.L_HI(net3711));
 sg13g2_tiehi \mem_addr[3]$_DFFE_PP__3712  (.L_HI(net3712));
 sg13g2_tiehi \mem_addr[4]$_DFFE_PP__3713  (.L_HI(net3713));
 sg13g2_tiehi \mem_addr[5]$_DFFE_PP__3714  (.L_HI(net3714));
 sg13g2_tiehi \mem_addr[6]$_DFFE_PP__3715  (.L_HI(net3715));
 sg13g2_tiehi \mem_addr[7]$_DFFE_PP__3716  (.L_HI(net3716));
 sg13g2_tiehi \mem_select$_SDFFE_PN0P__3717  (.L_HI(net3717));
 sg13g2_tiehi \mem_type_data$_DFFE_PP__3718  (.L_HI(net3718));
 sg13g2_tiehi \mem_write_en$_SDFFE_PN0P__3719  (.L_HI(net3719));
 sg13g2_tiehi \mem_write_value[0]$_DFFE_PP__3720  (.L_HI(net3720));
 sg13g2_tiehi \mem_write_value[1]$_DFFE_PP__3721  (.L_HI(net3721));
 sg13g2_tiehi \mem_write_value[2]$_DFFE_PP__3722  (.L_HI(net3722));
 sg13g2_tiehi \mem_write_value[3]$_DFFE_PP__3723  (.L_HI(net3723));
 sg13g2_tiehi \mem_write_value[4]$_DFFE_PP__3724  (.L_HI(net3724));
 sg13g2_tiehi \mem_write_value[5]$_DFFE_PP__3725  (.L_HI(net3725));
 sg13g2_tiehi \mem_write_value[6]$_DFFE_PP__3726  (.L_HI(net3726));
 sg13g2_tiehi \mem_write_value[7]$_DFFE_PP__3727  (.L_HI(net3727));
 sg13g2_tiehi \memory_input[0]$_DFFE_PP__3728  (.L_HI(net3728));
 sg13g2_tiehi \memory_input[1]$_DFFE_PP__3729  (.L_HI(net3729));
 sg13g2_tiehi \memory_input[2]$_DFFE_PP__3730  (.L_HI(net3730));
 sg13g2_tiehi \memory_input[3]$_DFFE_PP__3731  (.L_HI(net3731));
 sg13g2_tiehi \memory_input[4]$_DFFE_PP__3732  (.L_HI(net3732));
 sg13g2_tiehi \memory_input[5]$_DFFE_PP__3733  (.L_HI(net3733));
 sg13g2_tiehi \memory_input[6]$_DFFE_PP__3734  (.L_HI(net3734));
 sg13g2_tiehi \memory_input[7]$_DFFE_PP__3735  (.L_HI(net3735));
 sg13g2_tiehi \o_shift_out$_SDFF_PN0__3736  (.L_HI(net3736));
 sg13g2_tiehi \opcode[0]$_SDFF_PN0__3737  (.L_HI(net3737));
 sg13g2_tiehi \opcode[1]$_SDFF_PN0__3738  (.L_HI(net3738));
 sg13g2_tiehi \opcode[2]$_SDFF_PN0__3739  (.L_HI(net3739));
 sg13g2_tiehi \opcode[3]$_SDFF_PN0__3740  (.L_HI(net3740));
 sg13g2_tiehi \opcode[4]$_SDFF_PN0__3741  (.L_HI(net3741));
 sg13g2_tiehi \opcode[5]$_SDFF_PN0__3742  (.L_HI(net3742));
 sg13g2_tiehi \opcode[6]$_SDFF_PN0__3743  (.L_HI(net3743));
 sg13g2_tiehi \opcode[7]$_SDFF_PN0__3744  (.L_HI(net3744));
 sg13g2_tiehi \out_of_order_exec$_SDFFE_PP0P__3745  (.L_HI(net3745));
 sg13g2_tiehi \past_i_run$_SDFF_PN0__3746  (.L_HI(net3746));
 sg13g2_tiehi \pc[0]$_SDFFE_PN0P__3747  (.L_HI(net3747));
 sg13g2_tiehi \pc[1]$_SDFFE_PN0P__3748  (.L_HI(net3748));
 sg13g2_tiehi \pc[2]$_SDFFE_PN0P__3749  (.L_HI(net3749));
 sg13g2_tiehi \pc[3]$_SDFFE_PN0P__3750  (.L_HI(net3750));
 sg13g2_tiehi \pc[4]$_SDFFE_PN0P__3751  (.L_HI(net3751));
 sg13g2_tiehi \pc[5]$_SDFFE_PN0P__3752  (.L_HI(net3752));
 sg13g2_tiehi \pc[6]$_SDFFE_PN0P__3753  (.L_HI(net3753));
 sg13g2_tiehi \pc[7]$_SDFFE_PN0P__3754  (.L_HI(net3754));
 sg13g2_tiehi \shift_reg[0]$_SDFF_PN0__3755  (.L_HI(net3755));
 sg13g2_tiehi \shift_reg[1]$_SDFF_PN0__3756  (.L_HI(net3756));
 sg13g2_tiehi \shift_reg[2]$_SDFF_PN0__3757  (.L_HI(net3757));
 sg13g2_tiehi \shift_reg[3]$_SDFF_PN0__3758  (.L_HI(net3758));
 sg13g2_tiehi \shift_reg[4]$_SDFF_PN0__3759  (.L_HI(net3759));
 sg13g2_tiehi \shift_reg[5]$_SDFF_PN0__3760  (.L_HI(net3760));
 sg13g2_tiehi \shift_reg[6]$_SDFF_PN0__3761  (.L_HI(net3761));
 sg13g2_tiehi \shift_reg[7]$_SDFF_PN0__3762  (.L_HI(net3762));
 sg13g2_tiehi \single_step$_SDFFE_PN0P__3763  (.L_HI(net3763));
 sg13g2_tiehi \sp[0]$_SDFFE_PN0P__3764  (.L_HI(net3764));
 sg13g2_tiehi \sp[1]$_SDFFE_PN0P__3765  (.L_HI(net3765));
 sg13g2_tiehi \sp[2]$_SDFFE_PN0P__3766  (.L_HI(net3766));
 sg13g2_tiehi \sp[3]$_SDFFE_PN0P__3767  (.L_HI(net3767));
 sg13g2_tiehi \sp[4]$_SDFFE_PN0P__3768  (.L_HI(net3768));
 sg13g2_tiehi \stack[0][0]$_DFFE_PP__3769  (.L_HI(net3769));
 sg13g2_tiehi \stack[0][1]$_DFFE_PP__3770  (.L_HI(net3770));
 sg13g2_tiehi \stack[0][2]$_DFFE_PP__3771  (.L_HI(net3771));
 sg13g2_tiehi \stack[0][3]$_DFFE_PP__3772  (.L_HI(net3772));
 sg13g2_tiehi \stack[0][4]$_DFFE_PP__3773  (.L_HI(net3773));
 sg13g2_tiehi \stack[0][5]$_DFFE_PP__3774  (.L_HI(net3774));
 sg13g2_tiehi \stack[0][6]$_DFFE_PP__3775  (.L_HI(net3775));
 sg13g2_tiehi \stack[0][7]$_DFFE_PP__3776  (.L_HI(net3776));
 sg13g2_tiehi \stack[10][0]$_DFFE_PP__3777  (.L_HI(net3777));
 sg13g2_tiehi \stack[10][1]$_DFFE_PP__3778  (.L_HI(net3778));
 sg13g2_tiehi \stack[10][2]$_DFFE_PP__3779  (.L_HI(net3779));
 sg13g2_tiehi \stack[10][3]$_DFFE_PP__3780  (.L_HI(net3780));
 sg13g2_tiehi \stack[10][4]$_DFFE_PP__3781  (.L_HI(net3781));
 sg13g2_tiehi \stack[10][5]$_DFFE_PP__3782  (.L_HI(net3782));
 sg13g2_tiehi \stack[10][6]$_DFFE_PP__3783  (.L_HI(net3783));
 sg13g2_tiehi \stack[10][7]$_DFFE_PP__3784  (.L_HI(net3784));
 sg13g2_tiehi \stack[11][0]$_DFFE_PP__3785  (.L_HI(net3785));
 sg13g2_tiehi \stack[11][1]$_DFFE_PP__3786  (.L_HI(net3786));
 sg13g2_tiehi \stack[11][2]$_DFFE_PP__3787  (.L_HI(net3787));
 sg13g2_tiehi \stack[11][3]$_DFFE_PP__3788  (.L_HI(net3788));
 sg13g2_tiehi \stack[11][4]$_DFFE_PP__3789  (.L_HI(net3789));
 sg13g2_tiehi \stack[11][5]$_DFFE_PP__3790  (.L_HI(net3790));
 sg13g2_tiehi \stack[11][6]$_DFFE_PP__3791  (.L_HI(net3791));
 sg13g2_tiehi \stack[11][7]$_DFFE_PP__3792  (.L_HI(net3792));
 sg13g2_tiehi \stack[12][0]$_DFFE_PP__3793  (.L_HI(net3793));
 sg13g2_tiehi \stack[12][1]$_DFFE_PP__3794  (.L_HI(net3794));
 sg13g2_tiehi \stack[12][2]$_DFFE_PP__3795  (.L_HI(net3795));
 sg13g2_tiehi \stack[12][3]$_DFFE_PP__3796  (.L_HI(net3796));
 sg13g2_tiehi \stack[12][4]$_DFFE_PP__3797  (.L_HI(net3797));
 sg13g2_tiehi \stack[12][5]$_DFFE_PP__3798  (.L_HI(net3798));
 sg13g2_tiehi \stack[12][6]$_DFFE_PP__3799  (.L_HI(net3799));
 sg13g2_tiehi \stack[12][7]$_DFFE_PP__3800  (.L_HI(net3800));
 sg13g2_tiehi \stack[13][0]$_DFFE_PP__3801  (.L_HI(net3801));
 sg13g2_tiehi \stack[13][1]$_DFFE_PP__3802  (.L_HI(net3802));
 sg13g2_tiehi \stack[13][2]$_DFFE_PP__3803  (.L_HI(net3803));
 sg13g2_tiehi \stack[13][3]$_DFFE_PP__3804  (.L_HI(net3804));
 sg13g2_tiehi \stack[13][4]$_DFFE_PP__3805  (.L_HI(net3805));
 sg13g2_tiehi \stack[13][5]$_DFFE_PP__3806  (.L_HI(net3806));
 sg13g2_tiehi \stack[13][6]$_DFFE_PP__3807  (.L_HI(net3807));
 sg13g2_tiehi \stack[13][7]$_DFFE_PP__3808  (.L_HI(net3808));
 sg13g2_tiehi \stack[14][0]$_DFFE_PP__3809  (.L_HI(net3809));
 sg13g2_tiehi \stack[14][1]$_DFFE_PP__3810  (.L_HI(net3810));
 sg13g2_tiehi \stack[14][2]$_DFFE_PP__3811  (.L_HI(net3811));
 sg13g2_tiehi \stack[14][3]$_DFFE_PP__3812  (.L_HI(net3812));
 sg13g2_tiehi \stack[14][4]$_DFFE_PP__3813  (.L_HI(net3813));
 sg13g2_tiehi \stack[14][5]$_DFFE_PP__3814  (.L_HI(net3814));
 sg13g2_tiehi \stack[14][6]$_DFFE_PP__3815  (.L_HI(net3815));
 sg13g2_tiehi \stack[14][7]$_DFFE_PP__3816  (.L_HI(net3816));
 sg13g2_tiehi \stack[15][0]$_DFFE_PP__3817  (.L_HI(net3817));
 sg13g2_tiehi \stack[15][1]$_DFFE_PP__3818  (.L_HI(net3818));
 sg13g2_tiehi \stack[15][2]$_DFFE_PP__3819  (.L_HI(net3819));
 sg13g2_tiehi \stack[15][3]$_DFFE_PP__3820  (.L_HI(net3820));
 sg13g2_tiehi \stack[15][4]$_DFFE_PP__3821  (.L_HI(net3821));
 sg13g2_tiehi \stack[15][5]$_DFFE_PP__3822  (.L_HI(net3822));
 sg13g2_tiehi \stack[15][6]$_DFFE_PP__3823  (.L_HI(net3823));
 sg13g2_tiehi \stack[15][7]$_DFFE_PP__3824  (.L_HI(net3824));
 sg13g2_tiehi \stack[16][0]$_DFFE_PP__3825  (.L_HI(net3825));
 sg13g2_tiehi \stack[16][1]$_DFFE_PP__3826  (.L_HI(net3826));
 sg13g2_tiehi \stack[16][2]$_DFFE_PP__3827  (.L_HI(net3827));
 sg13g2_tiehi \stack[16][3]$_DFFE_PP__3828  (.L_HI(net3828));
 sg13g2_tiehi \stack[16][4]$_DFFE_PP__3829  (.L_HI(net3829));
 sg13g2_tiehi \stack[16][5]$_DFFE_PP__3830  (.L_HI(net3830));
 sg13g2_tiehi \stack[16][6]$_DFFE_PP__3831  (.L_HI(net3831));
 sg13g2_tiehi \stack[16][7]$_DFFE_PP__3832  (.L_HI(net3832));
 sg13g2_tiehi \stack[17][0]$_DFFE_PP__3833  (.L_HI(net3833));
 sg13g2_tiehi \stack[17][1]$_DFFE_PP__3834  (.L_HI(net3834));
 sg13g2_tiehi \stack[17][2]$_DFFE_PP__3835  (.L_HI(net3835));
 sg13g2_tiehi \stack[17][3]$_DFFE_PP__3836  (.L_HI(net3836));
 sg13g2_tiehi \stack[17][4]$_DFFE_PP__3837  (.L_HI(net3837));
 sg13g2_tiehi \stack[17][5]$_DFFE_PP__3838  (.L_HI(net3838));
 sg13g2_tiehi \stack[17][6]$_DFFE_PP__3839  (.L_HI(net3839));
 sg13g2_tiehi \stack[17][7]$_DFFE_PP__3840  (.L_HI(net3840));
 sg13g2_tiehi \stack[18][0]$_DFFE_PP__3841  (.L_HI(net3841));
 sg13g2_tiehi \stack[18][1]$_DFFE_PP__3842  (.L_HI(net3842));
 sg13g2_tiehi \stack[18][2]$_DFFE_PP__3843  (.L_HI(net3843));
 sg13g2_tiehi \stack[18][3]$_DFFE_PP__3844  (.L_HI(net3844));
 sg13g2_tiehi \stack[18][4]$_DFFE_PP__3845  (.L_HI(net3845));
 sg13g2_tiehi \stack[18][5]$_DFFE_PP__3846  (.L_HI(net3846));
 sg13g2_tiehi \stack[18][6]$_DFFE_PP__3847  (.L_HI(net3847));
 sg13g2_tiehi \stack[18][7]$_DFFE_PP__3848  (.L_HI(net3848));
 sg13g2_tiehi \stack[19][0]$_DFFE_PP__3849  (.L_HI(net3849));
 sg13g2_tiehi \stack[19][1]$_DFFE_PP__3850  (.L_HI(net3850));
 sg13g2_tiehi \stack[19][2]$_DFFE_PP__3851  (.L_HI(net3851));
 sg13g2_tiehi \stack[19][3]$_DFFE_PP__3852  (.L_HI(net3852));
 sg13g2_tiehi \stack[19][4]$_DFFE_PP__3853  (.L_HI(net3853));
 sg13g2_tiehi \stack[19][5]$_DFFE_PP__3854  (.L_HI(net3854));
 sg13g2_tiehi \stack[19][6]$_DFFE_PP__3855  (.L_HI(net3855));
 sg13g2_tiehi \stack[19][7]$_DFFE_PP__3856  (.L_HI(net3856));
 sg13g2_tiehi \stack[1][0]$_DFFE_PP__3857  (.L_HI(net3857));
 sg13g2_tiehi \stack[1][1]$_DFFE_PP__3858  (.L_HI(net3858));
 sg13g2_tiehi \stack[1][2]$_DFFE_PP__3859  (.L_HI(net3859));
 sg13g2_tiehi \stack[1][3]$_DFFE_PP__3860  (.L_HI(net3860));
 sg13g2_tiehi \stack[1][4]$_DFFE_PP__3861  (.L_HI(net3861));
 sg13g2_tiehi \stack[1][5]$_DFFE_PP__3862  (.L_HI(net3862));
 sg13g2_tiehi \stack[1][6]$_DFFE_PP__3863  (.L_HI(net3863));
 sg13g2_tiehi \stack[1][7]$_DFFE_PP__3864  (.L_HI(net3864));
 sg13g2_tiehi \stack[20][0]$_DFFE_PP__3865  (.L_HI(net3865));
 sg13g2_tiehi \stack[20][1]$_DFFE_PP__3866  (.L_HI(net3866));
 sg13g2_tiehi \stack[20][2]$_DFFE_PP__3867  (.L_HI(net3867));
 sg13g2_tiehi \stack[20][3]$_DFFE_PP__3868  (.L_HI(net3868));
 sg13g2_tiehi \stack[20][4]$_DFFE_PP__3869  (.L_HI(net3869));
 sg13g2_tiehi \stack[20][5]$_DFFE_PP__3870  (.L_HI(net3870));
 sg13g2_tiehi \stack[20][6]$_DFFE_PP__3871  (.L_HI(net3871));
 sg13g2_tiehi \stack[20][7]$_DFFE_PP__3872  (.L_HI(net3872));
 sg13g2_tiehi \stack[21][0]$_DFFE_PP__3873  (.L_HI(net3873));
 sg13g2_tiehi \stack[21][1]$_DFFE_PP__3874  (.L_HI(net3874));
 sg13g2_tiehi \stack[21][2]$_DFFE_PP__3875  (.L_HI(net3875));
 sg13g2_tiehi \stack[21][3]$_DFFE_PP__3876  (.L_HI(net3876));
 sg13g2_tiehi \stack[21][4]$_DFFE_PP__3877  (.L_HI(net3877));
 sg13g2_tiehi \stack[21][5]$_DFFE_PP__3878  (.L_HI(net3878));
 sg13g2_tiehi \stack[21][6]$_DFFE_PP__3879  (.L_HI(net3879));
 sg13g2_tiehi \stack[21][7]$_DFFE_PP__3880  (.L_HI(net3880));
 sg13g2_tiehi \stack[22][0]$_DFFE_PP__3881  (.L_HI(net3881));
 sg13g2_tiehi \stack[22][1]$_DFFE_PP__3882  (.L_HI(net3882));
 sg13g2_tiehi \stack[22][2]$_DFFE_PP__3883  (.L_HI(net3883));
 sg13g2_tiehi \stack[22][3]$_DFFE_PP__3884  (.L_HI(net3884));
 sg13g2_tiehi \stack[22][4]$_DFFE_PP__3885  (.L_HI(net3885));
 sg13g2_tiehi \stack[22][5]$_DFFE_PP__3886  (.L_HI(net3886));
 sg13g2_tiehi \stack[22][6]$_DFFE_PP__3887  (.L_HI(net3887));
 sg13g2_tiehi \stack[22][7]$_DFFE_PP__3888  (.L_HI(net3888));
 sg13g2_tiehi \stack[23][0]$_DFFE_PP__3889  (.L_HI(net3889));
 sg13g2_tiehi \stack[23][1]$_DFFE_PP__3890  (.L_HI(net3890));
 sg13g2_tiehi \stack[23][2]$_DFFE_PP__3891  (.L_HI(net3891));
 sg13g2_tiehi \stack[23][3]$_DFFE_PP__3892  (.L_HI(net3892));
 sg13g2_tiehi \stack[23][4]$_DFFE_PP__3893  (.L_HI(net3893));
 sg13g2_tiehi \stack[23][5]$_DFFE_PP__3894  (.L_HI(net3894));
 sg13g2_tiehi \stack[23][6]$_DFFE_PP__3895  (.L_HI(net3895));
 sg13g2_tiehi \stack[23][7]$_DFFE_PP__3896  (.L_HI(net3896));
 sg13g2_tiehi \stack[24][0]$_DFFE_PP__3897  (.L_HI(net3897));
 sg13g2_tiehi \stack[24][1]$_DFFE_PP__3898  (.L_HI(net3898));
 sg13g2_tiehi \stack[24][2]$_DFFE_PP__3899  (.L_HI(net3899));
 sg13g2_tiehi \stack[24][3]$_DFFE_PP__3900  (.L_HI(net3900));
 sg13g2_tiehi \stack[24][4]$_DFFE_PP__3901  (.L_HI(net3901));
 sg13g2_tiehi \stack[24][5]$_DFFE_PP__3902  (.L_HI(net3902));
 sg13g2_tiehi \stack[24][6]$_DFFE_PP__3903  (.L_HI(net3903));
 sg13g2_tiehi \stack[24][7]$_DFFE_PP__3904  (.L_HI(net3904));
 sg13g2_tiehi \stack[25][0]$_DFFE_PP__3905  (.L_HI(net3905));
 sg13g2_tiehi \stack[25][1]$_DFFE_PP__3906  (.L_HI(net3906));
 sg13g2_tiehi \stack[25][2]$_DFFE_PP__3907  (.L_HI(net3907));
 sg13g2_tiehi \stack[25][3]$_DFFE_PP__3908  (.L_HI(net3908));
 sg13g2_tiehi \stack[25][4]$_DFFE_PP__3909  (.L_HI(net3909));
 sg13g2_tiehi \stack[25][5]$_DFFE_PP__3910  (.L_HI(net3910));
 sg13g2_tiehi \stack[25][6]$_DFFE_PP__3911  (.L_HI(net3911));
 sg13g2_tiehi \stack[25][7]$_DFFE_PP__3912  (.L_HI(net3912));
 sg13g2_tiehi \stack[26][0]$_DFFE_PP__3913  (.L_HI(net3913));
 sg13g2_tiehi \stack[26][1]$_DFFE_PP__3914  (.L_HI(net3914));
 sg13g2_tiehi \stack[26][2]$_DFFE_PP__3915  (.L_HI(net3915));
 sg13g2_tiehi \stack[26][3]$_DFFE_PP__3916  (.L_HI(net3916));
 sg13g2_tiehi \stack[26][4]$_DFFE_PP__3917  (.L_HI(net3917));
 sg13g2_tiehi \stack[26][5]$_DFFE_PP__3918  (.L_HI(net3918));
 sg13g2_tiehi \stack[26][6]$_DFFE_PP__3919  (.L_HI(net3919));
 sg13g2_tiehi \stack[26][7]$_DFFE_PP__3920  (.L_HI(net3920));
 sg13g2_tiehi \stack[27][0]$_DFFE_PP__3921  (.L_HI(net3921));
 sg13g2_tiehi \stack[27][1]$_DFFE_PP__3922  (.L_HI(net3922));
 sg13g2_tiehi \stack[27][2]$_DFFE_PP__3923  (.L_HI(net3923));
 sg13g2_tiehi \stack[27][3]$_DFFE_PP__3924  (.L_HI(net3924));
 sg13g2_tiehi \stack[27][4]$_DFFE_PP__3925  (.L_HI(net3925));
 sg13g2_tiehi \stack[27][5]$_DFFE_PP__3926  (.L_HI(net3926));
 sg13g2_tiehi \stack[27][6]$_DFFE_PP__3927  (.L_HI(net3927));
 sg13g2_tiehi \stack[27][7]$_DFFE_PP__3928  (.L_HI(net3928));
 sg13g2_tiehi \stack[28][0]$_DFFE_PP__3929  (.L_HI(net3929));
 sg13g2_tiehi \stack[28][1]$_DFFE_PP__3930  (.L_HI(net3930));
 sg13g2_tiehi \stack[28][2]$_DFFE_PP__3931  (.L_HI(net3931));
 sg13g2_tiehi \stack[28][3]$_DFFE_PP__3932  (.L_HI(net3932));
 sg13g2_tiehi \stack[28][4]$_DFFE_PP__3933  (.L_HI(net3933));
 sg13g2_tiehi \stack[28][5]$_DFFE_PP__3934  (.L_HI(net3934));
 sg13g2_tiehi \stack[28][6]$_DFFE_PP__3935  (.L_HI(net3935));
 sg13g2_tiehi \stack[28][7]$_DFFE_PP__3936  (.L_HI(net3936));
 sg13g2_tiehi \stack[29][0]$_DFFE_PP__3937  (.L_HI(net3937));
 sg13g2_tiehi \stack[29][1]$_DFFE_PP__3938  (.L_HI(net3938));
 sg13g2_tiehi \stack[29][2]$_DFFE_PP__3939  (.L_HI(net3939));
 sg13g2_tiehi \stack[29][3]$_DFFE_PP__3940  (.L_HI(net3940));
 sg13g2_tiehi \stack[29][4]$_DFFE_PP__3941  (.L_HI(net3941));
 sg13g2_tiehi \stack[29][5]$_DFFE_PP__3942  (.L_HI(net3942));
 sg13g2_tiehi \stack[29][6]$_DFFE_PP__3943  (.L_HI(net3943));
 sg13g2_tiehi \stack[29][7]$_DFFE_PP__3944  (.L_HI(net3944));
 sg13g2_tiehi \stack[2][0]$_DFFE_PP__3945  (.L_HI(net3945));
 sg13g2_tiehi \stack[2][1]$_DFFE_PP__3946  (.L_HI(net3946));
 sg13g2_tiehi \stack[2][2]$_DFFE_PP__3947  (.L_HI(net3947));
 sg13g2_tiehi \stack[2][3]$_DFFE_PP__3948  (.L_HI(net3948));
 sg13g2_tiehi \stack[2][4]$_DFFE_PP__3949  (.L_HI(net3949));
 sg13g2_tiehi \stack[2][5]$_DFFE_PP__3950  (.L_HI(net3950));
 sg13g2_tiehi \stack[2][6]$_DFFE_PP__3951  (.L_HI(net3951));
 sg13g2_tiehi \stack[2][7]$_DFFE_PP__3952  (.L_HI(net3952));
 sg13g2_tiehi \stack[30][0]$_DFFE_PP__3953  (.L_HI(net3953));
 sg13g2_tiehi \stack[30][1]$_DFFE_PP__3954  (.L_HI(net3954));
 sg13g2_tiehi \stack[30][2]$_DFFE_PP__3955  (.L_HI(net3955));
 sg13g2_tiehi \stack[30][3]$_DFFE_PP__3956  (.L_HI(net3956));
 sg13g2_tiehi \stack[30][4]$_DFFE_PP__3957  (.L_HI(net3957));
 sg13g2_tiehi \stack[30][5]$_DFFE_PP__3958  (.L_HI(net3958));
 sg13g2_tiehi \stack[30][6]$_DFFE_PP__3959  (.L_HI(net3959));
 sg13g2_tiehi \stack[30][7]$_DFFE_PP__3960  (.L_HI(net3960));
 sg13g2_tiehi \stack[31][0]$_DFFE_PP__3961  (.L_HI(net3961));
 sg13g2_tiehi \stack[31][1]$_DFFE_PP__3962  (.L_HI(net3962));
 sg13g2_tiehi \stack[31][2]$_DFFE_PP__3963  (.L_HI(net3963));
 sg13g2_tiehi \stack[31][3]$_DFFE_PP__3964  (.L_HI(net3964));
 sg13g2_tiehi \stack[31][4]$_DFFE_PP__3965  (.L_HI(net3965));
 sg13g2_tiehi \stack[31][5]$_DFFE_PP__3966  (.L_HI(net3966));
 sg13g2_tiehi \stack[31][6]$_DFFE_PP__3967  (.L_HI(net3967));
 sg13g2_tiehi \stack[31][7]$_DFFE_PP__3968  (.L_HI(net3968));
 sg13g2_tiehi \stack[3][0]$_DFFE_PP__3969  (.L_HI(net3969));
 sg13g2_tiehi \stack[3][1]$_DFFE_PP__3970  (.L_HI(net3970));
 sg13g2_tiehi \stack[3][2]$_DFFE_PP__3971  (.L_HI(net3971));
 sg13g2_tiehi \stack[3][3]$_DFFE_PP__3972  (.L_HI(net3972));
 sg13g2_tiehi \stack[3][4]$_DFFE_PP__3973  (.L_HI(net3973));
 sg13g2_tiehi \stack[3][5]$_DFFE_PP__3974  (.L_HI(net3974));
 sg13g2_tiehi \stack[3][6]$_DFFE_PP__3975  (.L_HI(net3975));
 sg13g2_tiehi \stack[3][7]$_DFFE_PP__3976  (.L_HI(net3976));
 sg13g2_tiehi \stack[4][0]$_DFFE_PP__3977  (.L_HI(net3977));
 sg13g2_tiehi \stack[4][1]$_DFFE_PP__3978  (.L_HI(net3978));
 sg13g2_tiehi \stack[4][2]$_DFFE_PP__3979  (.L_HI(net3979));
 sg13g2_tiehi \stack[4][3]$_DFFE_PP__3980  (.L_HI(net3980));
 sg13g2_tiehi \stack[4][4]$_DFFE_PP__3981  (.L_HI(net3981));
 sg13g2_tiehi \stack[4][5]$_DFFE_PP__3982  (.L_HI(net3982));
 sg13g2_tiehi \stack[4][6]$_DFFE_PP__3983  (.L_HI(net3983));
 sg13g2_tiehi \stack[4][7]$_DFFE_PP__3984  (.L_HI(net3984));
 sg13g2_tiehi \stack[5][0]$_DFFE_PP__3985  (.L_HI(net3985));
 sg13g2_tiehi \stack[5][1]$_DFFE_PP__3986  (.L_HI(net3986));
 sg13g2_tiehi \stack[5][2]$_DFFE_PP__3987  (.L_HI(net3987));
 sg13g2_tiehi \stack[5][3]$_DFFE_PP__3988  (.L_HI(net3988));
 sg13g2_tiehi \stack[5][4]$_DFFE_PP__3989  (.L_HI(net3989));
 sg13g2_tiehi \stack[5][5]$_DFFE_PP__3990  (.L_HI(net3990));
 sg13g2_tiehi \stack[5][6]$_DFFE_PP__3991  (.L_HI(net3991));
 sg13g2_tiehi \stack[5][7]$_DFFE_PP__3992  (.L_HI(net3992));
 sg13g2_tiehi \stack[6][0]$_DFFE_PP__3993  (.L_HI(net3993));
 sg13g2_tiehi \stack[6][1]$_DFFE_PP__3994  (.L_HI(net3994));
 sg13g2_tiehi \stack[6][2]$_DFFE_PP__3995  (.L_HI(net3995));
 sg13g2_tiehi \stack[6][3]$_DFFE_PP__3996  (.L_HI(net3996));
 sg13g2_tiehi \stack[6][4]$_DFFE_PP__3997  (.L_HI(net3997));
 sg13g2_tiehi \stack[6][5]$_DFFE_PP__3998  (.L_HI(net3998));
 sg13g2_tiehi \stack[6][6]$_DFFE_PP__3999  (.L_HI(net3999));
 sg13g2_tiehi \stack[6][7]$_DFFE_PP__4000  (.L_HI(net4000));
 sg13g2_tiehi \stack[7][0]$_DFFE_PP__4001  (.L_HI(net4001));
 sg13g2_tiehi \stack[7][1]$_DFFE_PP__4002  (.L_HI(net4002));
 sg13g2_tiehi \stack[7][2]$_DFFE_PP__4003  (.L_HI(net4003));
 sg13g2_tiehi \stack[7][3]$_DFFE_PP__4004  (.L_HI(net4004));
 sg13g2_tiehi \stack[7][4]$_DFFE_PP__4005  (.L_HI(net4005));
 sg13g2_tiehi \stack[7][5]$_DFFE_PP__4006  (.L_HI(net4006));
 sg13g2_tiehi \stack[7][6]$_DFFE_PP__4007  (.L_HI(net4007));
 sg13g2_tiehi \stack[7][7]$_DFFE_PP__4008  (.L_HI(net4008));
 sg13g2_tiehi \stack[8][0]$_DFFE_PP__4009  (.L_HI(net4009));
 sg13g2_tiehi \stack[8][1]$_DFFE_PP__4010  (.L_HI(net4010));
 sg13g2_tiehi \stack[8][2]$_DFFE_PP__4011  (.L_HI(net4011));
 sg13g2_tiehi \stack[8][3]$_DFFE_PP__4012  (.L_HI(net4012));
 sg13g2_tiehi \stack[8][4]$_DFFE_PP__4013  (.L_HI(net4013));
 sg13g2_tiehi \stack[8][5]$_DFFE_PP__4014  (.L_HI(net4014));
 sg13g2_tiehi \stack[8][6]$_DFFE_PP__4015  (.L_HI(net4015));
 sg13g2_tiehi \stack[8][7]$_DFFE_PP__4016  (.L_HI(net4016));
 sg13g2_tiehi \stack[9][0]$_DFFE_PP__4017  (.L_HI(net4017));
 sg13g2_tiehi \stack[9][1]$_DFFE_PP__4018  (.L_HI(net4018));
 sg13g2_tiehi \stack[9][2]$_DFFE_PP__4019  (.L_HI(net4019));
 sg13g2_tiehi \stack[9][3]$_DFFE_PP__4020  (.L_HI(net4020));
 sg13g2_tiehi \stack[9][4]$_DFFE_PP__4021  (.L_HI(net4021));
 sg13g2_tiehi \stack[9][5]$_DFFE_PP__4022  (.L_HI(net4022));
 sg13g2_tiehi \stack[9][6]$_DFFE_PP__4023  (.L_HI(net4023));
 sg13g2_tiehi \stack[9][7]$_DFFE_PP__4024  (.L_HI(net4024));
 sg13g2_tiehi \state[0]$_DFF_P__4025  (.L_HI(net4025));
 sg13g2_tiehi \state[1]$_DFF_P__4026  (.L_HI(net4026));
 sg13g2_tiehi \state[2]$_DFF_P__4027  (.L_HI(net4027));
 sg13g2_tiehi \state[3]$_DFF_P__4028  (.L_HI(net4028));
 sg13g2_tiehi \state[4]$_DFF_P__4029  (.L_HI(net4029));
 sg13g2_tiehi \state[5]$_DFF_P__4030  (.L_HI(net4030));
 sg13g2_tiehi \state[6]$_DFF_P__4031  (.L_HI(net4031));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_8 clkbuf_leaf_313_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_8 clkbuf_leaf_314_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_314_clk));
 sg13g2_buf_8 clkbuf_leaf_315_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_315_clk));
 sg13g2_buf_8 clkbuf_leaf_316_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_316_clk));
 sg13g2_buf_8 clkbuf_leaf_317_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_317_clk));
 sg13g2_buf_8 clkbuf_leaf_318_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_318_clk));
 sg13g2_buf_8 clkbuf_leaf_319_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_319_clk));
 sg13g2_buf_8 clkbuf_leaf_320_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_320_clk));
 sg13g2_buf_8 clkbuf_leaf_321_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_321_clk));
 sg13g2_buf_8 clkbuf_leaf_322_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_322_clk));
 sg13g2_buf_8 clkbuf_leaf_323_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_323_clk));
 sg13g2_buf_8 clkbuf_leaf_324_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_324_clk));
 sg13g2_buf_8 clkbuf_leaf_325_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_325_clk));
 sg13g2_buf_8 clkbuf_leaf_326_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_326_clk));
 sg13g2_buf_8 clkbuf_leaf_327_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_327_clk));
 sg13g2_buf_8 clkbuf_leaf_328_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_328_clk));
 sg13g2_buf_8 clkbuf_leaf_329_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_329_clk));
 sg13g2_buf_8 clkbuf_leaf_330_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_330_clk));
 sg13g2_buf_8 clkbuf_leaf_331_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_331_clk));
 sg13g2_buf_8 clkbuf_leaf_332_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_332_clk));
 sg13g2_buf_8 clkbuf_leaf_333_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_333_clk));
 sg13g2_buf_8 clkbuf_leaf_334_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_334_clk));
 sg13g2_buf_8 clkbuf_leaf_335_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_335_clk));
 sg13g2_buf_8 clkbuf_leaf_336_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_336_clk));
 sg13g2_buf_8 clkbuf_leaf_337_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_337_clk));
 sg13g2_buf_8 clkbuf_leaf_338_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_338_clk));
 sg13g2_buf_8 clkbuf_leaf_339_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_339_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_1__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_5__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_6__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_9__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_10__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_13__leaf_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_6_14__leaf_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_6_17__leaf_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_6_22__leaf_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_6_25__leaf_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_6_26__leaf_clk));
 sg13g2_buf_8 clkload18 (.A(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_6_30__leaf_clk));
 sg13g2_buf_8 clkload21 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload22 (.A(clknet_6_33__leaf_clk));
 sg13g2_buf_8 clkload23 (.A(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkload24 (.A(clknet_6_37__leaf_clk));
 sg13g2_buf_8 clkload25 (.A(clknet_6_38__leaf_clk));
 sg13g2_buf_8 clkload26 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload27 (.A(clknet_6_41__leaf_clk));
 sg13g2_buf_8 clkload28 (.A(clknet_6_42__leaf_clk));
 sg13g2_buf_8 clkload29 (.A(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkload30 (.A(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkload31 (.A(clknet_6_46__leaf_clk));
 sg13g2_buf_8 clkload32 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload33 (.A(clknet_6_49__leaf_clk));
 sg13g2_buf_8 clkload34 (.A(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkload35 (.A(clknet_6_53__leaf_clk));
 sg13g2_buf_8 clkload36 (.A(clknet_6_54__leaf_clk));
 sg13g2_buf_8 clkload37 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload38 (.A(clknet_6_57__leaf_clk));
 sg13g2_buf_8 clkload39 (.A(clknet_6_58__leaf_clk));
 sg13g2_buf_8 clkload40 (.A(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkload41 (.A(clknet_6_61__leaf_clk));
 sg13g2_buf_8 clkload42 (.A(clknet_6_62__leaf_clk));
 sg13g2_buf_8 clkload43 (.A(clknet_6_63__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00017_));
 sg13g2_antennanp ANTENNA_2 (.A(_00017_));
 sg13g2_antennanp ANTENNA_3 (.A(_00017_));
 sg13g2_antennanp ANTENNA_4 (.A(_00017_));
 sg13g2_antennanp ANTENNA_5 (.A(_02490_));
 sg13g2_antennanp ANTENNA_6 (.A(_03341_));
 sg13g2_antennanp ANTENNA_7 (.A(_03444_));
 sg13g2_antennanp ANTENNA_8 (.A(_03444_));
 sg13g2_antennanp ANTENNA_9 (.A(_03444_));
 sg13g2_antennanp ANTENNA_10 (.A(_03621_));
 sg13g2_antennanp ANTENNA_11 (.A(_03621_));
 sg13g2_antennanp ANTENNA_12 (.A(_03621_));
 sg13g2_antennanp ANTENNA_13 (.A(_03621_));
 sg13g2_antennanp ANTENNA_14 (.A(_03621_));
 sg13g2_antennanp ANTENNA_15 (.A(_03621_));
 sg13g2_antennanp ANTENNA_16 (.A(_03621_));
 sg13g2_antennanp ANTENNA_17 (.A(_03621_));
 sg13g2_antennanp ANTENNA_18 (.A(_03843_));
 sg13g2_antennanp ANTENNA_19 (.A(_03843_));
 sg13g2_antennanp ANTENNA_20 (.A(_03843_));
 sg13g2_antennanp ANTENNA_21 (.A(_03843_));
 sg13g2_antennanp ANTENNA_22 (.A(_03850_));
 sg13g2_antennanp ANTENNA_23 (.A(_03850_));
 sg13g2_antennanp ANTENNA_24 (.A(_03850_));
 sg13g2_antennanp ANTENNA_25 (.A(_03850_));
 sg13g2_antennanp ANTENNA_26 (.A(_03850_));
 sg13g2_antennanp ANTENNA_27 (.A(_03850_));
 sg13g2_antennanp ANTENNA_28 (.A(_03850_));
 sg13g2_antennanp ANTENNA_29 (.A(_03850_));
 sg13g2_antennanp ANTENNA_30 (.A(_03855_));
 sg13g2_antennanp ANTENNA_31 (.A(_03855_));
 sg13g2_antennanp ANTENNA_32 (.A(_03855_));
 sg13g2_antennanp ANTENNA_33 (.A(_03875_));
 sg13g2_antennanp ANTENNA_34 (.A(_03995_));
 sg13g2_antennanp ANTENNA_35 (.A(_03995_));
 sg13g2_antennanp ANTENNA_36 (.A(_03995_));
 sg13g2_antennanp ANTENNA_37 (.A(_04431_));
 sg13g2_antennanp ANTENNA_38 (.A(_04431_));
 sg13g2_antennanp ANTENNA_39 (.A(_04431_));
 sg13g2_antennanp ANTENNA_40 (.A(_04431_));
 sg13g2_antennanp ANTENNA_41 (.A(_04431_));
 sg13g2_antennanp ANTENNA_42 (.A(_04431_));
 sg13g2_antennanp ANTENNA_43 (.A(_04431_));
 sg13g2_antennanp ANTENNA_44 (.A(_04431_));
 sg13g2_antennanp ANTENNA_45 (.A(_05432_));
 sg13g2_antennanp ANTENNA_46 (.A(_05432_));
 sg13g2_antennanp ANTENNA_47 (.A(_05432_));
 sg13g2_antennanp ANTENNA_48 (.A(_05441_));
 sg13g2_antennanp ANTENNA_49 (.A(_05441_));
 sg13g2_antennanp ANTENNA_50 (.A(_05441_));
 sg13g2_antennanp ANTENNA_51 (.A(_05446_));
 sg13g2_antennanp ANTENNA_52 (.A(_05446_));
 sg13g2_antennanp ANTENNA_53 (.A(_05446_));
 sg13g2_antennanp ANTENNA_54 (.A(_05446_));
 sg13g2_antennanp ANTENNA_55 (.A(_05449_));
 sg13g2_antennanp ANTENNA_56 (.A(_05449_));
 sg13g2_antennanp ANTENNA_57 (.A(_05449_));
 sg13g2_antennanp ANTENNA_58 (.A(_05453_));
 sg13g2_antennanp ANTENNA_59 (.A(_05453_));
 sg13g2_antennanp ANTENNA_60 (.A(_05453_));
 sg13g2_antennanp ANTENNA_61 (.A(_05453_));
 sg13g2_antennanp ANTENNA_62 (.A(_05453_));
 sg13g2_antennanp ANTENNA_63 (.A(_05453_));
 sg13g2_antennanp ANTENNA_64 (.A(_05453_));
 sg13g2_antennanp ANTENNA_65 (.A(_05453_));
 sg13g2_antennanp ANTENNA_66 (.A(_05453_));
 sg13g2_antennanp ANTENNA_67 (.A(_05453_));
 sg13g2_antennanp ANTENNA_68 (.A(_05457_));
 sg13g2_antennanp ANTENNA_69 (.A(_05457_));
 sg13g2_antennanp ANTENNA_70 (.A(_05457_));
 sg13g2_antennanp ANTENNA_71 (.A(_05457_));
 sg13g2_antennanp ANTENNA_72 (.A(_05457_));
 sg13g2_antennanp ANTENNA_73 (.A(_05457_));
 sg13g2_antennanp ANTENNA_74 (.A(_05463_));
 sg13g2_antennanp ANTENNA_75 (.A(_05463_));
 sg13g2_antennanp ANTENNA_76 (.A(_05463_));
 sg13g2_antennanp ANTENNA_77 (.A(_05463_));
 sg13g2_antennanp ANTENNA_78 (.A(_05463_));
 sg13g2_antennanp ANTENNA_79 (.A(_05463_));
 sg13g2_antennanp ANTENNA_80 (.A(_05467_));
 sg13g2_antennanp ANTENNA_81 (.A(_05467_));
 sg13g2_antennanp ANTENNA_82 (.A(_05467_));
 sg13g2_antennanp ANTENNA_83 (.A(_05467_));
 sg13g2_antennanp ANTENNA_84 (.A(_05467_));
 sg13g2_antennanp ANTENNA_85 (.A(_05467_));
 sg13g2_antennanp ANTENNA_86 (.A(_05471_));
 sg13g2_antennanp ANTENNA_87 (.A(_05471_));
 sg13g2_antennanp ANTENNA_88 (.A(_05471_));
 sg13g2_antennanp ANTENNA_89 (.A(_05471_));
 sg13g2_antennanp ANTENNA_90 (.A(_05471_));
 sg13g2_antennanp ANTENNA_91 (.A(_05471_));
 sg13g2_antennanp ANTENNA_92 (.A(_05471_));
 sg13g2_antennanp ANTENNA_93 (.A(_05471_));
 sg13g2_antennanp ANTENNA_94 (.A(_05471_));
 sg13g2_antennanp ANTENNA_95 (.A(_05471_));
 sg13g2_antennanp ANTENNA_96 (.A(_05476_));
 sg13g2_antennanp ANTENNA_97 (.A(_05476_));
 sg13g2_antennanp ANTENNA_98 (.A(_05498_));
 sg13g2_antennanp ANTENNA_99 (.A(_05498_));
 sg13g2_antennanp ANTENNA_100 (.A(_05542_));
 sg13g2_antennanp ANTENNA_101 (.A(_06148_));
 sg13g2_antennanp ANTENNA_102 (.A(_06148_));
 sg13g2_antennanp ANTENNA_103 (.A(_06148_));
 sg13g2_antennanp ANTENNA_104 (.A(_06148_));
 sg13g2_antennanp ANTENNA_105 (.A(_06148_));
 sg13g2_antennanp ANTENNA_106 (.A(_06153_));
 sg13g2_antennanp ANTENNA_107 (.A(_06153_));
 sg13g2_antennanp ANTENNA_108 (.A(_06153_));
 sg13g2_antennanp ANTENNA_109 (.A(_06153_));
 sg13g2_antennanp ANTENNA_110 (.A(_06153_));
 sg13g2_antennanp ANTENNA_111 (.A(_06153_));
 sg13g2_antennanp ANTENNA_112 (.A(_06153_));
 sg13g2_antennanp ANTENNA_113 (.A(_06153_));
 sg13g2_antennanp ANTENNA_114 (.A(_06171_));
 sg13g2_antennanp ANTENNA_115 (.A(_06189_));
 sg13g2_antennanp ANTENNA_116 (.A(_06253_));
 sg13g2_antennanp ANTENNA_117 (.A(_06255_));
 sg13g2_antennanp ANTENNA_118 (.A(_06268_));
 sg13g2_antennanp ANTENNA_119 (.A(_06293_));
 sg13g2_antennanp ANTENNA_120 (.A(_06298_));
 sg13g2_antennanp ANTENNA_121 (.A(_06311_));
 sg13g2_antennanp ANTENNA_122 (.A(_06329_));
 sg13g2_antennanp ANTENNA_123 (.A(_06339_));
 sg13g2_antennanp ANTENNA_124 (.A(_06339_));
 sg13g2_antennanp ANTENNA_125 (.A(_06339_));
 sg13g2_antennanp ANTENNA_126 (.A(_06339_));
 sg13g2_antennanp ANTENNA_127 (.A(_06339_));
 sg13g2_antennanp ANTENNA_128 (.A(_06339_));
 sg13g2_antennanp ANTENNA_129 (.A(_06339_));
 sg13g2_antennanp ANTENNA_130 (.A(_06339_));
 sg13g2_antennanp ANTENNA_131 (.A(_06339_));
 sg13g2_antennanp ANTENNA_132 (.A(_06339_));
 sg13g2_antennanp ANTENNA_133 (.A(_06339_));
 sg13g2_antennanp ANTENNA_134 (.A(_06339_));
 sg13g2_antennanp ANTENNA_135 (.A(_06339_));
 sg13g2_antennanp ANTENNA_136 (.A(_06393_));
 sg13g2_antennanp ANTENNA_137 (.A(_06393_));
 sg13g2_antennanp ANTENNA_138 (.A(_06393_));
 sg13g2_antennanp ANTENNA_139 (.A(_06393_));
 sg13g2_antennanp ANTENNA_140 (.A(_06393_));
 sg13g2_antennanp ANTENNA_141 (.A(_06393_));
 sg13g2_antennanp ANTENNA_142 (.A(_06393_));
 sg13g2_antennanp ANTENNA_143 (.A(_06393_));
 sg13g2_antennanp ANTENNA_144 (.A(_06410_));
 sg13g2_antennanp ANTENNA_145 (.A(_06410_));
 sg13g2_antennanp ANTENNA_146 (.A(_06410_));
 sg13g2_antennanp ANTENNA_147 (.A(_06410_));
 sg13g2_antennanp ANTENNA_148 (.A(_06410_));
 sg13g2_antennanp ANTENNA_149 (.A(_06416_));
 sg13g2_antennanp ANTENNA_150 (.A(_06460_));
 sg13g2_antennanp ANTENNA_151 (.A(_06493_));
 sg13g2_antennanp ANTENNA_152 (.A(_06493_));
 sg13g2_antennanp ANTENNA_153 (.A(_06516_));
 sg13g2_antennanp ANTENNA_154 (.A(_06516_));
 sg13g2_antennanp ANTENNA_155 (.A(_06518_));
 sg13g2_antennanp ANTENNA_156 (.A(_06520_));
 sg13g2_antennanp ANTENNA_157 (.A(_06559_));
 sg13g2_antennanp ANTENNA_158 (.A(_06559_));
 sg13g2_antennanp ANTENNA_159 (.A(_06595_));
 sg13g2_antennanp ANTENNA_160 (.A(_06601_));
 sg13g2_antennanp ANTENNA_161 (.A(_06616_));
 sg13g2_antennanp ANTENNA_162 (.A(_06616_));
 sg13g2_antennanp ANTENNA_163 (.A(_06618_));
 sg13g2_antennanp ANTENNA_164 (.A(_06619_));
 sg13g2_antennanp ANTENNA_165 (.A(_06620_));
 sg13g2_antennanp ANTENNA_166 (.A(_06658_));
 sg13g2_antennanp ANTENNA_167 (.A(_06694_));
 sg13g2_antennanp ANTENNA_168 (.A(_06700_));
 sg13g2_antennanp ANTENNA_169 (.A(_06715_));
 sg13g2_antennanp ANTENNA_170 (.A(_06715_));
 sg13g2_antennanp ANTENNA_171 (.A(_06718_));
 sg13g2_antennanp ANTENNA_172 (.A(_06719_));
 sg13g2_antennanp ANTENNA_173 (.A(_06757_));
 sg13g2_antennanp ANTENNA_174 (.A(_06772_));
 sg13g2_antennanp ANTENNA_175 (.A(_06772_));
 sg13g2_antennanp ANTENNA_176 (.A(_06793_));
 sg13g2_antennanp ANTENNA_177 (.A(_06793_));
 sg13g2_antennanp ANTENNA_178 (.A(_06799_));
 sg13g2_antennanp ANTENNA_179 (.A(_06814_));
 sg13g2_antennanp ANTENNA_180 (.A(_06814_));
 sg13g2_antennanp ANTENNA_181 (.A(_06818_));
 sg13g2_antennanp ANTENNA_182 (.A(_06856_));
 sg13g2_antennanp ANTENNA_183 (.A(_06870_));
 sg13g2_antennanp ANTENNA_184 (.A(_06870_));
 sg13g2_antennanp ANTENNA_185 (.A(_06871_));
 sg13g2_antennanp ANTENNA_186 (.A(_06871_));
 sg13g2_antennanp ANTENNA_187 (.A(_06913_));
 sg13g2_antennanp ANTENNA_188 (.A(_06913_));
 sg13g2_antennanp ANTENNA_189 (.A(_06917_));
 sg13g2_antennanp ANTENNA_190 (.A(_06955_));
 sg13g2_antennanp ANTENNA_191 (.A(_06975_));
 sg13g2_antennanp ANTENNA_192 (.A(_06991_));
 sg13g2_antennanp ANTENNA_193 (.A(_07012_));
 sg13g2_antennanp ANTENNA_194 (.A(_07012_));
 sg13g2_antennanp ANTENNA_195 (.A(_07016_));
 sg13g2_antennanp ANTENNA_196 (.A(_07054_));
 sg13g2_antennanp ANTENNA_197 (.A(_07069_));
 sg13g2_antennanp ANTENNA_198 (.A(_07069_));
 sg13g2_antennanp ANTENNA_199 (.A(_07074_));
 sg13g2_antennanp ANTENNA_200 (.A(_07090_));
 sg13g2_antennanp ANTENNA_201 (.A(_07090_));
 sg13g2_antennanp ANTENNA_202 (.A(_07096_));
 sg13g2_antennanp ANTENNA_203 (.A(_07105_));
 sg13g2_antennanp ANTENNA_204 (.A(_07335_));
 sg13g2_antennanp ANTENNA_205 (.A(_07416_));
 sg13g2_antennanp ANTENNA_206 (.A(_07416_));
 sg13g2_antennanp ANTENNA_207 (.A(_07416_));
 sg13g2_antennanp ANTENNA_208 (.A(_07416_));
 sg13g2_antennanp ANTENNA_209 (.A(_07416_));
 sg13g2_antennanp ANTENNA_210 (.A(_07416_));
 sg13g2_antennanp ANTENNA_211 (.A(_09194_));
 sg13g2_antennanp ANTENNA_212 (.A(_09194_));
 sg13g2_antennanp ANTENNA_213 (.A(_09194_));
 sg13g2_antennanp ANTENNA_214 (.A(_09194_));
 sg13g2_antennanp ANTENNA_215 (.A(_09260_));
 sg13g2_antennanp ANTENNA_216 (.A(_09260_));
 sg13g2_antennanp ANTENNA_217 (.A(_09260_));
 sg13g2_antennanp ANTENNA_218 (.A(_09260_));
 sg13g2_antennanp ANTENNA_219 (.A(_09260_));
 sg13g2_antennanp ANTENNA_220 (.A(_09260_));
 sg13g2_antennanp ANTENNA_221 (.A(_09260_));
 sg13g2_antennanp ANTENNA_222 (.A(_09260_));
 sg13g2_antennanp ANTENNA_223 (.A(_09260_));
 sg13g2_antennanp ANTENNA_224 (.A(_09260_));
 sg13g2_antennanp ANTENNA_225 (.A(_09260_));
 sg13g2_antennanp ANTENNA_226 (.A(_09260_));
 sg13g2_antennanp ANTENNA_227 (.A(_09260_));
 sg13g2_antennanp ANTENNA_228 (.A(_09260_));
 sg13g2_antennanp ANTENNA_229 (.A(_09260_));
 sg13g2_antennanp ANTENNA_230 (.A(_09260_));
 sg13g2_antennanp ANTENNA_231 (.A(_09260_));
 sg13g2_antennanp ANTENNA_232 (.A(_09260_));
 sg13g2_antennanp ANTENNA_233 (.A(_09273_));
 sg13g2_antennanp ANTENNA_234 (.A(_09273_));
 sg13g2_antennanp ANTENNA_235 (.A(_09273_));
 sg13g2_antennanp ANTENNA_236 (.A(_09273_));
 sg13g2_antennanp ANTENNA_237 (.A(_09273_));
 sg13g2_antennanp ANTENNA_238 (.A(_09273_));
 sg13g2_antennanp ANTENNA_239 (.A(_09273_));
 sg13g2_antennanp ANTENNA_240 (.A(_09273_));
 sg13g2_antennanp ANTENNA_241 (.A(_09273_));
 sg13g2_antennanp ANTENNA_242 (.A(_09345_));
 sg13g2_antennanp ANTENNA_243 (.A(_09345_));
 sg13g2_antennanp ANTENNA_244 (.A(_09345_));
 sg13g2_antennanp ANTENNA_245 (.A(_09345_));
 sg13g2_antennanp ANTENNA_246 (.A(_09345_));
 sg13g2_antennanp ANTENNA_247 (.A(_09345_));
 sg13g2_antennanp ANTENNA_248 (.A(_09345_));
 sg13g2_antennanp ANTENNA_249 (.A(_09345_));
 sg13g2_antennanp ANTENNA_250 (.A(_09345_));
 sg13g2_antennanp ANTENNA_251 (.A(_09418_));
 sg13g2_antennanp ANTENNA_252 (.A(_09418_));
 sg13g2_antennanp ANTENNA_253 (.A(_09418_));
 sg13g2_antennanp ANTENNA_254 (.A(_09418_));
 sg13g2_antennanp ANTENNA_255 (.A(_09418_));
 sg13g2_antennanp ANTENNA_256 (.A(_09418_));
 sg13g2_antennanp ANTENNA_257 (.A(_09418_));
 sg13g2_antennanp ANTENNA_258 (.A(_09418_));
 sg13g2_antennanp ANTENNA_259 (.A(_09418_));
 sg13g2_antennanp ANTENNA_260 (.A(_09906_));
 sg13g2_antennanp ANTENNA_261 (.A(_09906_));
 sg13g2_antennanp ANTENNA_262 (.A(_09906_));
 sg13g2_antennanp ANTENNA_263 (.A(_09906_));
 sg13g2_antennanp ANTENNA_264 (.A(_09906_));
 sg13g2_antennanp ANTENNA_265 (.A(_09906_));
 sg13g2_antennanp ANTENNA_266 (.A(_09906_));
 sg13g2_antennanp ANTENNA_267 (.A(_09906_));
 sg13g2_antennanp ANTENNA_268 (.A(_09906_));
 sg13g2_antennanp ANTENNA_269 (.A(_09906_));
 sg13g2_antennanp ANTENNA_270 (.A(_09906_));
 sg13g2_antennanp ANTENNA_271 (.A(_09906_));
 sg13g2_antennanp ANTENNA_272 (.A(_09906_));
 sg13g2_antennanp ANTENNA_273 (.A(_09906_));
 sg13g2_antennanp ANTENNA_274 (.A(_09928_));
 sg13g2_antennanp ANTENNA_275 (.A(_09928_));
 sg13g2_antennanp ANTENNA_276 (.A(_09928_));
 sg13g2_antennanp ANTENNA_277 (.A(_09928_));
 sg13g2_antennanp ANTENNA_278 (.A(_09928_));
 sg13g2_antennanp ANTENNA_279 (.A(_09928_));
 sg13g2_antennanp ANTENNA_280 (.A(_09928_));
 sg13g2_antennanp ANTENNA_281 (.A(_09928_));
 sg13g2_antennanp ANTENNA_282 (.A(_09928_));
 sg13g2_antennanp ANTENNA_283 (.A(_09928_));
 sg13g2_antennanp ANTENNA_284 (.A(_09928_));
 sg13g2_antennanp ANTENNA_285 (.A(_09928_));
 sg13g2_antennanp ANTENNA_286 (.A(_09928_));
 sg13g2_antennanp ANTENNA_287 (.A(_09928_));
 sg13g2_antennanp ANTENNA_288 (.A(_09928_));
 sg13g2_antennanp ANTENNA_289 (.A(_09928_));
 sg13g2_antennanp ANTENNA_290 (.A(_09929_));
 sg13g2_antennanp ANTENNA_291 (.A(_09929_));
 sg13g2_antennanp ANTENNA_292 (.A(_09929_));
 sg13g2_antennanp ANTENNA_293 (.A(_09929_));
 sg13g2_antennanp ANTENNA_294 (.A(_09930_));
 sg13g2_antennanp ANTENNA_295 (.A(_09930_));
 sg13g2_antennanp ANTENNA_296 (.A(_09935_));
 sg13g2_antennanp ANTENNA_297 (.A(_09935_));
 sg13g2_antennanp ANTENNA_298 (.A(_09935_));
 sg13g2_antennanp ANTENNA_299 (.A(_09935_));
 sg13g2_antennanp ANTENNA_300 (.A(_09935_));
 sg13g2_antennanp ANTENNA_301 (.A(_09935_));
 sg13g2_antennanp ANTENNA_302 (.A(_09935_));
 sg13g2_antennanp ANTENNA_303 (.A(_09935_));
 sg13g2_antennanp ANTENNA_304 (.A(_09935_));
 sg13g2_antennanp ANTENNA_305 (.A(_09935_));
 sg13g2_antennanp ANTENNA_306 (.A(_09935_));
 sg13g2_antennanp ANTENNA_307 (.A(_09935_));
 sg13g2_antennanp ANTENNA_308 (.A(_09935_));
 sg13g2_antennanp ANTENNA_309 (.A(_09935_));
 sg13g2_antennanp ANTENNA_310 (.A(_09935_));
 sg13g2_antennanp ANTENNA_311 (.A(_09935_));
 sg13g2_antennanp ANTENNA_312 (.A(_09935_));
 sg13g2_antennanp ANTENNA_313 (.A(_09935_));
 sg13g2_antennanp ANTENNA_314 (.A(_09935_));
 sg13g2_antennanp ANTENNA_315 (.A(_09935_));
 sg13g2_antennanp ANTENNA_316 (.A(_09986_));
 sg13g2_antennanp ANTENNA_317 (.A(_09986_));
 sg13g2_antennanp ANTENNA_318 (.A(_09986_));
 sg13g2_antennanp ANTENNA_319 (.A(_09986_));
 sg13g2_antennanp ANTENNA_320 (.A(_09986_));
 sg13g2_antennanp ANTENNA_321 (.A(_10040_));
 sg13g2_antennanp ANTENNA_322 (.A(_10040_));
 sg13g2_antennanp ANTENNA_323 (.A(_10040_));
 sg13g2_antennanp ANTENNA_324 (.A(_10042_));
 sg13g2_antennanp ANTENNA_325 (.A(_10042_));
 sg13g2_antennanp ANTENNA_326 (.A(_10042_));
 sg13g2_antennanp ANTENNA_327 (.A(_10042_));
 sg13g2_antennanp ANTENNA_328 (.A(_10046_));
 sg13g2_antennanp ANTENNA_329 (.A(_10048_));
 sg13g2_antennanp ANTENNA_330 (.A(_10051_));
 sg13g2_antennanp ANTENNA_331 (.A(_10053_));
 sg13g2_antennanp ANTENNA_332 (.A(_10071_));
 sg13g2_antennanp ANTENNA_333 (.A(_10071_));
 sg13g2_antennanp ANTENNA_334 (.A(_10071_));
 sg13g2_antennanp ANTENNA_335 (.A(_10071_));
 sg13g2_antennanp ANTENNA_336 (.A(_10071_));
 sg13g2_antennanp ANTENNA_337 (.A(_10071_));
 sg13g2_antennanp ANTENNA_338 (.A(_10080_));
 sg13g2_antennanp ANTENNA_339 (.A(_10080_));
 sg13g2_antennanp ANTENNA_340 (.A(_10080_));
 sg13g2_antennanp ANTENNA_341 (.A(_10080_));
 sg13g2_antennanp ANTENNA_342 (.A(_10083_));
 sg13g2_antennanp ANTENNA_343 (.A(_10091_));
 sg13g2_antennanp ANTENNA_344 (.A(_10101_));
 sg13g2_antennanp ANTENNA_345 (.A(_10106_));
 sg13g2_antennanp ANTENNA_346 (.A(_10110_));
 sg13g2_antennanp ANTENNA_347 (.A(_10121_));
 sg13g2_antennanp ANTENNA_348 (.A(_10131_));
 sg13g2_antennanp ANTENNA_349 (.A(_10136_));
 sg13g2_antennanp ANTENNA_350 (.A(_10140_));
 sg13g2_antennanp ANTENNA_351 (.A(_10226_));
 sg13g2_antennanp ANTENNA_352 (.A(_10226_));
 sg13g2_antennanp ANTENNA_353 (.A(_10226_));
 sg13g2_antennanp ANTENNA_354 (.A(_10232_));
 sg13g2_antennanp ANTENNA_355 (.A(_10232_));
 sg13g2_antennanp ANTENNA_356 (.A(_10232_));
 sg13g2_antennanp ANTENNA_357 (.A(_10232_));
 sg13g2_antennanp ANTENNA_358 (.A(_10232_));
 sg13g2_antennanp ANTENNA_359 (.A(_10232_));
 sg13g2_antennanp ANTENNA_360 (.A(_10232_));
 sg13g2_antennanp ANTENNA_361 (.A(_10235_));
 sg13g2_antennanp ANTENNA_362 (.A(_10235_));
 sg13g2_antennanp ANTENNA_363 (.A(_10235_));
 sg13g2_antennanp ANTENNA_364 (.A(_10235_));
 sg13g2_antennanp ANTENNA_365 (.A(_10236_));
 sg13g2_antennanp ANTENNA_366 (.A(_10236_));
 sg13g2_antennanp ANTENNA_367 (.A(_10236_));
 sg13g2_antennanp ANTENNA_368 (.A(_10236_));
 sg13g2_antennanp ANTENNA_369 (.A(_10236_));
 sg13g2_antennanp ANTENNA_370 (.A(_10236_));
 sg13g2_antennanp ANTENNA_371 (.A(_10243_));
 sg13g2_antennanp ANTENNA_372 (.A(_10243_));
 sg13g2_antennanp ANTENNA_373 (.A(_10243_));
 sg13g2_antennanp ANTENNA_374 (.A(_10243_));
 sg13g2_antennanp ANTENNA_375 (.A(_10243_));
 sg13g2_antennanp ANTENNA_376 (.A(_10243_));
 sg13g2_antennanp ANTENNA_377 (.A(_10256_));
 sg13g2_antennanp ANTENNA_378 (.A(_10256_));
 sg13g2_antennanp ANTENNA_379 (.A(_10256_));
 sg13g2_antennanp ANTENNA_380 (.A(_10256_));
 sg13g2_antennanp ANTENNA_381 (.A(_10287_));
 sg13g2_antennanp ANTENNA_382 (.A(_10287_));
 sg13g2_antennanp ANTENNA_383 (.A(_10287_));
 sg13g2_antennanp ANTENNA_384 (.A(_10287_));
 sg13g2_antennanp ANTENNA_385 (.A(_10287_));
 sg13g2_antennanp ANTENNA_386 (.A(_10295_));
 sg13g2_antennanp ANTENNA_387 (.A(_10295_));
 sg13g2_antennanp ANTENNA_388 (.A(_10295_));
 sg13g2_antennanp ANTENNA_389 (.A(_10295_));
 sg13g2_antennanp ANTENNA_390 (.A(_10295_));
 sg13g2_antennanp ANTENNA_391 (.A(_10295_));
 sg13g2_antennanp ANTENNA_392 (.A(_10295_));
 sg13g2_antennanp ANTENNA_393 (.A(_10295_));
 sg13g2_antennanp ANTENNA_394 (.A(_10325_));
 sg13g2_antennanp ANTENNA_395 (.A(_10325_));
 sg13g2_antennanp ANTENNA_396 (.A(_10325_));
 sg13g2_antennanp ANTENNA_397 (.A(_10325_));
 sg13g2_antennanp ANTENNA_398 (.A(_10325_));
 sg13g2_antennanp ANTENNA_399 (.A(_10325_));
 sg13g2_antennanp ANTENNA_400 (.A(_10325_));
 sg13g2_antennanp ANTENNA_401 (.A(_10325_));
 sg13g2_antennanp ANTENNA_402 (.A(_10325_));
 sg13g2_antennanp ANTENNA_403 (.A(_10325_));
 sg13g2_antennanp ANTENNA_404 (.A(_10325_));
 sg13g2_antennanp ANTENNA_405 (.A(_10325_));
 sg13g2_antennanp ANTENNA_406 (.A(_10326_));
 sg13g2_antennanp ANTENNA_407 (.A(_10326_));
 sg13g2_antennanp ANTENNA_408 (.A(_10326_));
 sg13g2_antennanp ANTENNA_409 (.A(_10349_));
 sg13g2_antennanp ANTENNA_410 (.A(_10349_));
 sg13g2_antennanp ANTENNA_411 (.A(_10349_));
 sg13g2_antennanp ANTENNA_412 (.A(_10349_));
 sg13g2_antennanp ANTENNA_413 (.A(_10350_));
 sg13g2_antennanp ANTENNA_414 (.A(_10350_));
 sg13g2_antennanp ANTENNA_415 (.A(_10350_));
 sg13g2_antennanp ANTENNA_416 (.A(_10373_));
 sg13g2_antennanp ANTENNA_417 (.A(_10373_));
 sg13g2_antennanp ANTENNA_418 (.A(_10373_));
 sg13g2_antennanp ANTENNA_419 (.A(_10373_));
 sg13g2_antennanp ANTENNA_420 (.A(_10373_));
 sg13g2_antennanp ANTENNA_421 (.A(_10373_));
 sg13g2_antennanp ANTENNA_422 (.A(_10373_));
 sg13g2_antennanp ANTENNA_423 (.A(_10373_));
 sg13g2_antennanp ANTENNA_424 (.A(_10373_));
 sg13g2_antennanp ANTENNA_425 (.A(_10373_));
 sg13g2_antennanp ANTENNA_426 (.A(_10397_));
 sg13g2_antennanp ANTENNA_427 (.A(_10397_));
 sg13g2_antennanp ANTENNA_428 (.A(_10397_));
 sg13g2_antennanp ANTENNA_429 (.A(_10397_));
 sg13g2_antennanp ANTENNA_430 (.A(_10397_));
 sg13g2_antennanp ANTENNA_431 (.A(_10397_));
 sg13g2_antennanp ANTENNA_432 (.A(_10397_));
 sg13g2_antennanp ANTENNA_433 (.A(_10397_));
 sg13g2_antennanp ANTENNA_434 (.A(_10415_));
 sg13g2_antennanp ANTENNA_435 (.A(_10415_));
 sg13g2_antennanp ANTENNA_436 (.A(_10415_));
 sg13g2_antennanp ANTENNA_437 (.A(_10415_));
 sg13g2_antennanp ANTENNA_438 (.A(_10415_));
 sg13g2_antennanp ANTENNA_439 (.A(_10415_));
 sg13g2_antennanp ANTENNA_440 (.A(_10415_));
 sg13g2_antennanp ANTENNA_441 (.A(_10415_));
 sg13g2_antennanp ANTENNA_442 (.A(_10415_));
 sg13g2_antennanp ANTENNA_443 (.A(_10415_));
 sg13g2_antennanp ANTENNA_444 (.A(_10415_));
 sg13g2_antennanp ANTENNA_445 (.A(_10415_));
 sg13g2_antennanp ANTENNA_446 (.A(_10415_));
 sg13g2_antennanp ANTENNA_447 (.A(_10415_));
 sg13g2_antennanp ANTENNA_448 (.A(_10415_));
 sg13g2_antennanp ANTENNA_449 (.A(_10415_));
 sg13g2_antennanp ANTENNA_450 (.A(_10415_));
 sg13g2_antennanp ANTENNA_451 (.A(_10415_));
 sg13g2_antennanp ANTENNA_452 (.A(_10415_));
 sg13g2_antennanp ANTENNA_453 (.A(_10415_));
 sg13g2_antennanp ANTENNA_454 (.A(_10415_));
 sg13g2_antennanp ANTENNA_455 (.A(_10415_));
 sg13g2_antennanp ANTENNA_456 (.A(_10415_));
 sg13g2_antennanp ANTENNA_457 (.A(_10415_));
 sg13g2_antennanp ANTENNA_458 (.A(_10415_));
 sg13g2_antennanp ANTENNA_459 (.A(_10415_));
 sg13g2_antennanp ANTENNA_460 (.A(_10422_));
 sg13g2_antennanp ANTENNA_461 (.A(_10422_));
 sg13g2_antennanp ANTENNA_462 (.A(_10422_));
 sg13g2_antennanp ANTENNA_463 (.A(_10422_));
 sg13g2_antennanp ANTENNA_464 (.A(_10422_));
 sg13g2_antennanp ANTENNA_465 (.A(_10422_));
 sg13g2_antennanp ANTENNA_466 (.A(_10422_));
 sg13g2_antennanp ANTENNA_467 (.A(_10422_));
 sg13g2_antennanp ANTENNA_468 (.A(_10422_));
 sg13g2_antennanp ANTENNA_469 (.A(_10422_));
 sg13g2_antennanp ANTENNA_470 (.A(_10422_));
 sg13g2_antennanp ANTENNA_471 (.A(_10422_));
 sg13g2_antennanp ANTENNA_472 (.A(_10422_));
 sg13g2_antennanp ANTENNA_473 (.A(_10422_));
 sg13g2_antennanp ANTENNA_474 (.A(_10422_));
 sg13g2_antennanp ANTENNA_475 (.A(_10422_));
 sg13g2_antennanp ANTENNA_476 (.A(_10422_));
 sg13g2_antennanp ANTENNA_477 (.A(_10444_));
 sg13g2_antennanp ANTENNA_478 (.A(_10444_));
 sg13g2_antennanp ANTENNA_479 (.A(_10444_));
 sg13g2_antennanp ANTENNA_480 (.A(_10444_));
 sg13g2_antennanp ANTENNA_481 (.A(_10444_));
 sg13g2_antennanp ANTENNA_482 (.A(_10444_));
 sg13g2_antennanp ANTENNA_483 (.A(_10444_));
 sg13g2_antennanp ANTENNA_484 (.A(_10444_));
 sg13g2_antennanp ANTENNA_485 (.A(_10444_));
 sg13g2_antennanp ANTENNA_486 (.A(_10444_));
 sg13g2_antennanp ANTENNA_487 (.A(_10444_));
 sg13g2_antennanp ANTENNA_488 (.A(_10444_));
 sg13g2_antennanp ANTENNA_489 (.A(_10444_));
 sg13g2_antennanp ANTENNA_490 (.A(_10444_));
 sg13g2_antennanp ANTENNA_491 (.A(_10444_));
 sg13g2_antennanp ANTENNA_492 (.A(_10444_));
 sg13g2_antennanp ANTENNA_493 (.A(_10444_));
 sg13g2_antennanp ANTENNA_494 (.A(_10445_));
 sg13g2_antennanp ANTENNA_495 (.A(_10445_));
 sg13g2_antennanp ANTENNA_496 (.A(_10445_));
 sg13g2_antennanp ANTENNA_497 (.A(_10468_));
 sg13g2_antennanp ANTENNA_498 (.A(_10468_));
 sg13g2_antennanp ANTENNA_499 (.A(_10468_));
 sg13g2_antennanp ANTENNA_500 (.A(_10468_));
 sg13g2_antennanp ANTENNA_501 (.A(_10468_));
 sg13g2_antennanp ANTENNA_502 (.A(_10468_));
 sg13g2_antennanp ANTENNA_503 (.A(_10468_));
 sg13g2_antennanp ANTENNA_504 (.A(_10468_));
 sg13g2_antennanp ANTENNA_505 (.A(_10468_));
 sg13g2_antennanp ANTENNA_506 (.A(_10468_));
 sg13g2_antennanp ANTENNA_507 (.A(_10491_));
 sg13g2_antennanp ANTENNA_508 (.A(_10491_));
 sg13g2_antennanp ANTENNA_509 (.A(_10491_));
 sg13g2_antennanp ANTENNA_510 (.A(_10491_));
 sg13g2_antennanp ANTENNA_511 (.A(_10491_));
 sg13g2_antennanp ANTENNA_512 (.A(_10491_));
 sg13g2_antennanp ANTENNA_513 (.A(_10491_));
 sg13g2_antennanp ANTENNA_514 (.A(_10491_));
 sg13g2_antennanp ANTENNA_515 (.A(_10491_));
 sg13g2_antennanp ANTENNA_516 (.A(_10491_));
 sg13g2_antennanp ANTENNA_517 (.A(_10491_));
 sg13g2_antennanp ANTENNA_518 (.A(_10513_));
 sg13g2_antennanp ANTENNA_519 (.A(_10513_));
 sg13g2_antennanp ANTENNA_520 (.A(_10513_));
 sg13g2_antennanp ANTENNA_521 (.A(_10513_));
 sg13g2_antennanp ANTENNA_522 (.A(_10513_));
 sg13g2_antennanp ANTENNA_523 (.A(_10513_));
 sg13g2_antennanp ANTENNA_524 (.A(_10513_));
 sg13g2_antennanp ANTENNA_525 (.A(_10514_));
 sg13g2_antennanp ANTENNA_526 (.A(_10514_));
 sg13g2_antennanp ANTENNA_527 (.A(_10514_));
 sg13g2_antennanp ANTENNA_528 (.A(_10514_));
 sg13g2_antennanp ANTENNA_529 (.A(_10514_));
 sg13g2_antennanp ANTENNA_530 (.A(_10514_));
 sg13g2_antennanp ANTENNA_531 (.A(_10514_));
 sg13g2_antennanp ANTENNA_532 (.A(_10514_));
 sg13g2_antennanp ANTENNA_533 (.A(_10514_));
 sg13g2_antennanp ANTENNA_534 (.A(_10514_));
 sg13g2_antennanp ANTENNA_535 (.A(_10564_));
 sg13g2_antennanp ANTENNA_536 (.A(_10564_));
 sg13g2_antennanp ANTENNA_537 (.A(_10564_));
 sg13g2_antennanp ANTENNA_538 (.A(_10564_));
 sg13g2_antennanp ANTENNA_539 (.A(_10564_));
 sg13g2_antennanp ANTENNA_540 (.A(_10564_));
 sg13g2_antennanp ANTENNA_541 (.A(_10564_));
 sg13g2_antennanp ANTENNA_542 (.A(_10564_));
 sg13g2_antennanp ANTENNA_543 (.A(_10564_));
 sg13g2_antennanp ANTENNA_544 (.A(_10564_));
 sg13g2_antennanp ANTENNA_545 (.A(_10564_));
 sg13g2_antennanp ANTENNA_546 (.A(_10564_));
 sg13g2_antennanp ANTENNA_547 (.A(_10564_));
 sg13g2_antennanp ANTENNA_548 (.A(_10564_));
 sg13g2_antennanp ANTENNA_549 (.A(_10564_));
 sg13g2_antennanp ANTENNA_550 (.A(_10565_));
 sg13g2_antennanp ANTENNA_551 (.A(_10565_));
 sg13g2_antennanp ANTENNA_552 (.A(_10565_));
 sg13g2_antennanp ANTENNA_553 (.A(_10565_));
 sg13g2_antennanp ANTENNA_554 (.A(_10565_));
 sg13g2_antennanp ANTENNA_555 (.A(_10565_));
 sg13g2_antennanp ANTENNA_556 (.A(_10565_));
 sg13g2_antennanp ANTENNA_557 (.A(_10565_));
 sg13g2_antennanp ANTENNA_558 (.A(_10586_));
 sg13g2_antennanp ANTENNA_559 (.A(_10586_));
 sg13g2_antennanp ANTENNA_560 (.A(_10586_));
 sg13g2_antennanp ANTENNA_561 (.A(_10586_));
 sg13g2_antennanp ANTENNA_562 (.A(_10586_));
 sg13g2_antennanp ANTENNA_563 (.A(_10586_));
 sg13g2_antennanp ANTENNA_564 (.A(_10586_));
 sg13g2_antennanp ANTENNA_565 (.A(_10586_));
 sg13g2_antennanp ANTENNA_566 (.A(_10586_));
 sg13g2_antennanp ANTENNA_567 (.A(_10586_));
 sg13g2_antennanp ANTENNA_568 (.A(_10586_));
 sg13g2_antennanp ANTENNA_569 (.A(_10586_));
 sg13g2_antennanp ANTENNA_570 (.A(_10586_));
 sg13g2_antennanp ANTENNA_571 (.A(_10586_));
 sg13g2_antennanp ANTENNA_572 (.A(_10587_));
 sg13g2_antennanp ANTENNA_573 (.A(_10587_));
 sg13g2_antennanp ANTENNA_574 (.A(_10587_));
 sg13g2_antennanp ANTENNA_575 (.A(_10587_));
 sg13g2_antennanp ANTENNA_576 (.A(_10632_));
 sg13g2_antennanp ANTENNA_577 (.A(_10632_));
 sg13g2_antennanp ANTENNA_578 (.A(_10632_));
 sg13g2_antennanp ANTENNA_579 (.A(_10632_));
 sg13g2_antennanp ANTENNA_580 (.A(_10632_));
 sg13g2_antennanp ANTENNA_581 (.A(_10632_));
 sg13g2_antennanp ANTENNA_582 (.A(_10632_));
 sg13g2_antennanp ANTENNA_583 (.A(_10632_));
 sg13g2_antennanp ANTENNA_584 (.A(_10632_));
 sg13g2_antennanp ANTENNA_585 (.A(_10632_));
 sg13g2_antennanp ANTENNA_586 (.A(_10632_));
 sg13g2_antennanp ANTENNA_587 (.A(_10632_));
 sg13g2_antennanp ANTENNA_588 (.A(_10632_));
 sg13g2_antennanp ANTENNA_589 (.A(_10632_));
 sg13g2_antennanp ANTENNA_590 (.A(_10632_));
 sg13g2_antennanp ANTENNA_591 (.A(_10633_));
 sg13g2_antennanp ANTENNA_592 (.A(_10633_));
 sg13g2_antennanp ANTENNA_593 (.A(_10633_));
 sg13g2_antennanp ANTENNA_594 (.A(_10633_));
 sg13g2_antennanp ANTENNA_595 (.A(_10633_));
 sg13g2_antennanp ANTENNA_596 (.A(_10656_));
 sg13g2_antennanp ANTENNA_597 (.A(_10656_));
 sg13g2_antennanp ANTENNA_598 (.A(_10656_));
 sg13g2_antennanp ANTENNA_599 (.A(_10656_));
 sg13g2_antennanp ANTENNA_600 (.A(_10656_));
 sg13g2_antennanp ANTENNA_601 (.A(_10656_));
 sg13g2_antennanp ANTENNA_602 (.A(_10656_));
 sg13g2_antennanp ANTENNA_603 (.A(_10657_));
 sg13g2_antennanp ANTENNA_604 (.A(_10657_));
 sg13g2_antennanp ANTENNA_605 (.A(_10657_));
 sg13g2_antennanp ANTENNA_606 (.A(_10679_));
 sg13g2_antennanp ANTENNA_607 (.A(_10679_));
 sg13g2_antennanp ANTENNA_608 (.A(_10679_));
 sg13g2_antennanp ANTENNA_609 (.A(_10679_));
 sg13g2_antennanp ANTENNA_610 (.A(_10679_));
 sg13g2_antennanp ANTENNA_611 (.A(_10679_));
 sg13g2_antennanp ANTENNA_612 (.A(_10679_));
 sg13g2_antennanp ANTENNA_613 (.A(_10679_));
 sg13g2_antennanp ANTENNA_614 (.A(_10679_));
 sg13g2_antennanp ANTENNA_615 (.A(_10679_));
 sg13g2_antennanp ANTENNA_616 (.A(_10679_));
 sg13g2_antennanp ANTENNA_617 (.A(_10679_));
 sg13g2_antennanp ANTENNA_618 (.A(_10680_));
 sg13g2_antennanp ANTENNA_619 (.A(_10680_));
 sg13g2_antennanp ANTENNA_620 (.A(_10680_));
 sg13g2_antennanp ANTENNA_621 (.A(_11171_));
 sg13g2_antennanp ANTENNA_622 (.A(_11171_));
 sg13g2_antennanp ANTENNA_623 (.A(_11171_));
 sg13g2_antennanp ANTENNA_624 (.A(_11171_));
 sg13g2_antennanp ANTENNA_625 (.A(_11171_));
 sg13g2_antennanp ANTENNA_626 (.A(_11171_));
 sg13g2_antennanp ANTENNA_627 (.A(_11171_));
 sg13g2_antennanp ANTENNA_628 (.A(_11734_));
 sg13g2_antennanp ANTENNA_629 (.A(_11875_));
 sg13g2_antennanp ANTENNA_630 (.A(_11875_));
 sg13g2_antennanp ANTENNA_631 (.A(_11875_));
 sg13g2_antennanp ANTENNA_632 (.A(_11875_));
 sg13g2_antennanp ANTENNA_633 (.A(_11875_));
 sg13g2_antennanp ANTENNA_634 (.A(_11875_));
 sg13g2_antennanp ANTENNA_635 (.A(_11875_));
 sg13g2_antennanp ANTENNA_636 (.A(_11875_));
 sg13g2_antennanp ANTENNA_637 (.A(_11875_));
 sg13g2_antennanp ANTENNA_638 (.A(_11875_));
 sg13g2_antennanp ANTENNA_639 (.A(_11875_));
 sg13g2_antennanp ANTENNA_640 (.A(_11875_));
 sg13g2_antennanp ANTENNA_641 (.A(_11875_));
 sg13g2_antennanp ANTENNA_642 (.A(_11875_));
 sg13g2_antennanp ANTENNA_643 (.A(_11875_));
 sg13g2_antennanp ANTENNA_644 (.A(_11875_));
 sg13g2_antennanp ANTENNA_645 (.A(_11875_));
 sg13g2_antennanp ANTENNA_646 (.A(_11875_));
 sg13g2_antennanp ANTENNA_647 (.A(_11875_));
 sg13g2_antennanp ANTENNA_648 (.A(_11875_));
 sg13g2_antennanp ANTENNA_649 (.A(_11875_));
 sg13g2_antennanp ANTENNA_650 (.A(_11875_));
 sg13g2_antennanp ANTENNA_651 (.A(_11875_));
 sg13g2_antennanp ANTENNA_652 (.A(_11875_));
 sg13g2_antennanp ANTENNA_653 (.A(_11875_));
 sg13g2_antennanp ANTENNA_654 (.A(_11875_));
 sg13g2_antennanp ANTENNA_655 (.A(_11875_));
 sg13g2_antennanp ANTENNA_656 (.A(_11875_));
 sg13g2_antennanp ANTENNA_657 (.A(_11875_));
 sg13g2_antennanp ANTENNA_658 (.A(_11875_));
 sg13g2_antennanp ANTENNA_659 (.A(_12403_));
 sg13g2_antennanp ANTENNA_660 (.A(_12403_));
 sg13g2_antennanp ANTENNA_661 (.A(_12403_));
 sg13g2_antennanp ANTENNA_662 (.A(_12403_));
 sg13g2_antennanp ANTENNA_663 (.A(_12431_));
 sg13g2_antennanp ANTENNA_664 (.A(_12431_));
 sg13g2_antennanp ANTENNA_665 (.A(_12431_));
 sg13g2_antennanp ANTENNA_666 (.A(_12431_));
 sg13g2_antennanp ANTENNA_667 (.A(_12434_));
 sg13g2_antennanp ANTENNA_668 (.A(_12434_));
 sg13g2_antennanp ANTENNA_669 (.A(_12434_));
 sg13g2_antennanp ANTENNA_670 (.A(_12443_));
 sg13g2_antennanp ANTENNA_671 (.A(_12443_));
 sg13g2_antennanp ANTENNA_672 (.A(_12443_));
 sg13g2_antennanp ANTENNA_673 (.A(_12630_));
 sg13g2_antennanp ANTENNA_674 (.A(_12630_));
 sg13g2_antennanp ANTENNA_675 (.A(_12630_));
 sg13g2_antennanp ANTENNA_676 (.A(_12649_));
 sg13g2_antennanp ANTENNA_677 (.A(_12649_));
 sg13g2_antennanp ANTENNA_678 (.A(_12649_));
 sg13g2_antennanp ANTENNA_679 (.A(_12649_));
 sg13g2_antennanp ANTENNA_680 (.A(_12649_));
 sg13g2_antennanp ANTENNA_681 (.A(_12649_));
 sg13g2_antennanp ANTENNA_682 (.A(_12649_));
 sg13g2_antennanp ANTENNA_683 (.A(_12649_));
 sg13g2_antennanp ANTENNA_684 (.A(_12649_));
 sg13g2_antennanp ANTENNA_685 (.A(_12649_));
 sg13g2_antennanp ANTENNA_686 (.A(_12649_));
 sg13g2_antennanp ANTENNA_687 (.A(_12649_));
 sg13g2_antennanp ANTENNA_688 (.A(_12649_));
 sg13g2_antennanp ANTENNA_689 (.A(_12653_));
 sg13g2_antennanp ANTENNA_690 (.A(_12653_));
 sg13g2_antennanp ANTENNA_691 (.A(_12653_));
 sg13g2_antennanp ANTENNA_692 (.A(_12653_));
 sg13g2_antennanp ANTENNA_693 (.A(_12653_));
 sg13g2_antennanp ANTENNA_694 (.A(_12653_));
 sg13g2_antennanp ANTENNA_695 (.A(_12653_));
 sg13g2_antennanp ANTENNA_696 (.A(_12653_));
 sg13g2_antennanp ANTENNA_697 (.A(_12654_));
 sg13g2_antennanp ANTENNA_698 (.A(_12654_));
 sg13g2_antennanp ANTENNA_699 (.A(_12654_));
 sg13g2_antennanp ANTENNA_700 (.A(_12658_));
 sg13g2_antennanp ANTENNA_701 (.A(_12658_));
 sg13g2_antennanp ANTENNA_702 (.A(_12658_));
 sg13g2_antennanp ANTENNA_703 (.A(_12658_));
 sg13g2_antennanp ANTENNA_704 (.A(_12662_));
 sg13g2_antennanp ANTENNA_705 (.A(_12662_));
 sg13g2_antennanp ANTENNA_706 (.A(_12662_));
 sg13g2_antennanp ANTENNA_707 (.A(_12662_));
 sg13g2_antennanp ANTENNA_708 (.A(_12849_));
 sg13g2_antennanp ANTENNA_709 (.A(clk));
 sg13g2_antennanp ANTENNA_710 (.A(clk));
 sg13g2_antennanp ANTENNA_711 (.A(\mem.data_in[1] ));
 sg13g2_antennanp ANTENNA_712 (.A(\mem.io_data_out[3] ));
 sg13g2_antennanp ANTENNA_713 (.A(\mem.io_data_out[3] ));
 sg13g2_antennanp ANTENNA_714 (.A(\mem.io_data_out[7] ));
 sg13g2_antennanp ANTENNA_715 (.A(\mem.io_data_out[7] ));
 sg13g2_antennanp ANTENNA_716 (.A(\mem.mem_internal.code_mem[24][0] ));
 sg13g2_antennanp ANTENNA_717 (.A(\mem.mem_internal.code_mem[24][0] ));
 sg13g2_antennanp ANTENNA_718 (.A(\mem.mem_internal.code_mem[24][0] ));
 sg13g2_antennanp ANTENNA_719 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_720 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_721 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_722 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_723 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_724 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_725 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_726 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_727 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_728 (.A(net1));
 sg13g2_antennanp ANTENNA_729 (.A(net1));
 sg13g2_antennanp ANTENNA_730 (.A(net1));
 sg13g2_antennanp ANTENNA_731 (.A(net2));
 sg13g2_antennanp ANTENNA_732 (.A(net2));
 sg13g2_antennanp ANTENNA_733 (.A(net4));
 sg13g2_antennanp ANTENNA_734 (.A(net527));
 sg13g2_antennanp ANTENNA_735 (.A(net527));
 sg13g2_antennanp ANTENNA_736 (.A(net527));
 sg13g2_antennanp ANTENNA_737 (.A(net527));
 sg13g2_antennanp ANTENNA_738 (.A(net527));
 sg13g2_antennanp ANTENNA_739 (.A(net527));
 sg13g2_antennanp ANTENNA_740 (.A(net527));
 sg13g2_antennanp ANTENNA_741 (.A(net527));
 sg13g2_antennanp ANTENNA_742 (.A(net527));
 sg13g2_antennanp ANTENNA_743 (.A(net527));
 sg13g2_antennanp ANTENNA_744 (.A(net527));
 sg13g2_antennanp ANTENNA_745 (.A(net527));
 sg13g2_antennanp ANTENNA_746 (.A(net527));
 sg13g2_antennanp ANTENNA_747 (.A(net527));
 sg13g2_antennanp ANTENNA_748 (.A(net529));
 sg13g2_antennanp ANTENNA_749 (.A(net529));
 sg13g2_antennanp ANTENNA_750 (.A(net529));
 sg13g2_antennanp ANTENNA_751 (.A(net529));
 sg13g2_antennanp ANTENNA_752 (.A(net529));
 sg13g2_antennanp ANTENNA_753 (.A(net529));
 sg13g2_antennanp ANTENNA_754 (.A(net529));
 sg13g2_antennanp ANTENNA_755 (.A(net529));
 sg13g2_antennanp ANTENNA_756 (.A(net529));
 sg13g2_antennanp ANTENNA_757 (.A(net529));
 sg13g2_antennanp ANTENNA_758 (.A(net529));
 sg13g2_antennanp ANTENNA_759 (.A(net529));
 sg13g2_antennanp ANTENNA_760 (.A(net549));
 sg13g2_antennanp ANTENNA_761 (.A(net549));
 sg13g2_antennanp ANTENNA_762 (.A(net549));
 sg13g2_antennanp ANTENNA_763 (.A(net549));
 sg13g2_antennanp ANTENNA_764 (.A(net549));
 sg13g2_antennanp ANTENNA_765 (.A(net549));
 sg13g2_antennanp ANTENNA_766 (.A(net549));
 sg13g2_antennanp ANTENNA_767 (.A(net549));
 sg13g2_antennanp ANTENNA_768 (.A(net549));
 sg13g2_antennanp ANTENNA_769 (.A(net549));
 sg13g2_antennanp ANTENNA_770 (.A(net549));
 sg13g2_antennanp ANTENNA_771 (.A(net549));
 sg13g2_antennanp ANTENNA_772 (.A(net549));
 sg13g2_antennanp ANTENNA_773 (.A(net549));
 sg13g2_antennanp ANTENNA_774 (.A(net549));
 sg13g2_antennanp ANTENNA_775 (.A(net549));
 sg13g2_antennanp ANTENNA_776 (.A(net549));
 sg13g2_antennanp ANTENNA_777 (.A(net549));
 sg13g2_antennanp ANTENNA_778 (.A(net549));
 sg13g2_antennanp ANTENNA_779 (.A(net549));
 sg13g2_antennanp ANTENNA_780 (.A(net549));
 sg13g2_antennanp ANTENNA_781 (.A(net551));
 sg13g2_antennanp ANTENNA_782 (.A(net551));
 sg13g2_antennanp ANTENNA_783 (.A(net551));
 sg13g2_antennanp ANTENNA_784 (.A(net551));
 sg13g2_antennanp ANTENNA_785 (.A(net551));
 sg13g2_antennanp ANTENNA_786 (.A(net551));
 sg13g2_antennanp ANTENNA_787 (.A(net551));
 sg13g2_antennanp ANTENNA_788 (.A(net551));
 sg13g2_antennanp ANTENNA_789 (.A(net551));
 sg13g2_antennanp ANTENNA_790 (.A(net551));
 sg13g2_antennanp ANTENNA_791 (.A(net551));
 sg13g2_antennanp ANTENNA_792 (.A(net551));
 sg13g2_antennanp ANTENNA_793 (.A(net551));
 sg13g2_antennanp ANTENNA_794 (.A(net551));
 sg13g2_antennanp ANTENNA_795 (.A(net551));
 sg13g2_antennanp ANTENNA_796 (.A(net551));
 sg13g2_antennanp ANTENNA_797 (.A(net551));
 sg13g2_antennanp ANTENNA_798 (.A(net551));
 sg13g2_antennanp ANTENNA_799 (.A(net551));
 sg13g2_antennanp ANTENNA_800 (.A(net552));
 sg13g2_antennanp ANTENNA_801 (.A(net552));
 sg13g2_antennanp ANTENNA_802 (.A(net552));
 sg13g2_antennanp ANTENNA_803 (.A(net552));
 sg13g2_antennanp ANTENNA_804 (.A(net552));
 sg13g2_antennanp ANTENNA_805 (.A(net552));
 sg13g2_antennanp ANTENNA_806 (.A(net552));
 sg13g2_antennanp ANTENNA_807 (.A(net552));
 sg13g2_antennanp ANTENNA_808 (.A(net552));
 sg13g2_antennanp ANTENNA_809 (.A(net552));
 sg13g2_antennanp ANTENNA_810 (.A(net552));
 sg13g2_antennanp ANTENNA_811 (.A(net552));
 sg13g2_antennanp ANTENNA_812 (.A(net552));
 sg13g2_antennanp ANTENNA_813 (.A(net553));
 sg13g2_antennanp ANTENNA_814 (.A(net553));
 sg13g2_antennanp ANTENNA_815 (.A(net553));
 sg13g2_antennanp ANTENNA_816 (.A(net553));
 sg13g2_antennanp ANTENNA_817 (.A(net553));
 sg13g2_antennanp ANTENNA_818 (.A(net553));
 sg13g2_antennanp ANTENNA_819 (.A(net553));
 sg13g2_antennanp ANTENNA_820 (.A(net553));
 sg13g2_antennanp ANTENNA_821 (.A(net553));
 sg13g2_antennanp ANTENNA_822 (.A(net553));
 sg13g2_antennanp ANTENNA_823 (.A(net553));
 sg13g2_antennanp ANTENNA_824 (.A(net553));
 sg13g2_antennanp ANTENNA_825 (.A(net553));
 sg13g2_antennanp ANTENNA_826 (.A(net553));
 sg13g2_antennanp ANTENNA_827 (.A(net553));
 sg13g2_antennanp ANTENNA_828 (.A(net553));
 sg13g2_antennanp ANTENNA_829 (.A(net553));
 sg13g2_antennanp ANTENNA_830 (.A(net553));
 sg13g2_antennanp ANTENNA_831 (.A(net553));
 sg13g2_antennanp ANTENNA_832 (.A(net553));
 sg13g2_antennanp ANTENNA_833 (.A(net554));
 sg13g2_antennanp ANTENNA_834 (.A(net554));
 sg13g2_antennanp ANTENNA_835 (.A(net554));
 sg13g2_antennanp ANTENNA_836 (.A(net554));
 sg13g2_antennanp ANTENNA_837 (.A(net554));
 sg13g2_antennanp ANTENNA_838 (.A(net554));
 sg13g2_antennanp ANTENNA_839 (.A(net554));
 sg13g2_antennanp ANTENNA_840 (.A(net554));
 sg13g2_antennanp ANTENNA_841 (.A(net554));
 sg13g2_antennanp ANTENNA_842 (.A(net554));
 sg13g2_antennanp ANTENNA_843 (.A(net554));
 sg13g2_antennanp ANTENNA_844 (.A(net554));
 sg13g2_antennanp ANTENNA_845 (.A(net554));
 sg13g2_antennanp ANTENNA_846 (.A(net554));
 sg13g2_antennanp ANTENNA_847 (.A(net554));
 sg13g2_antennanp ANTENNA_848 (.A(net554));
 sg13g2_antennanp ANTENNA_849 (.A(net554));
 sg13g2_antennanp ANTENNA_850 (.A(net554));
 sg13g2_antennanp ANTENNA_851 (.A(net554));
 sg13g2_antennanp ANTENNA_852 (.A(net554));
 sg13g2_antennanp ANTENNA_853 (.A(net554));
 sg13g2_antennanp ANTENNA_854 (.A(net554));
 sg13g2_antennanp ANTENNA_855 (.A(net554));
 sg13g2_antennanp ANTENNA_856 (.A(net554));
 sg13g2_antennanp ANTENNA_857 (.A(net554));
 sg13g2_antennanp ANTENNA_858 (.A(net554));
 sg13g2_antennanp ANTENNA_859 (.A(net554));
 sg13g2_antennanp ANTENNA_860 (.A(net554));
 sg13g2_antennanp ANTENNA_861 (.A(net554));
 sg13g2_antennanp ANTENNA_862 (.A(net554));
 sg13g2_antennanp ANTENNA_863 (.A(net554));
 sg13g2_antennanp ANTENNA_864 (.A(net554));
 sg13g2_antennanp ANTENNA_865 (.A(net554));
 sg13g2_antennanp ANTENNA_866 (.A(net554));
 sg13g2_antennanp ANTENNA_867 (.A(net554));
 sg13g2_antennanp ANTENNA_868 (.A(net554));
 sg13g2_antennanp ANTENNA_869 (.A(net556));
 sg13g2_antennanp ANTENNA_870 (.A(net556));
 sg13g2_antennanp ANTENNA_871 (.A(net556));
 sg13g2_antennanp ANTENNA_872 (.A(net556));
 sg13g2_antennanp ANTENNA_873 (.A(net556));
 sg13g2_antennanp ANTENNA_874 (.A(net556));
 sg13g2_antennanp ANTENNA_875 (.A(net556));
 sg13g2_antennanp ANTENNA_876 (.A(net556));
 sg13g2_antennanp ANTENNA_877 (.A(net556));
 sg13g2_antennanp ANTENNA_878 (.A(net556));
 sg13g2_antennanp ANTENNA_879 (.A(net556));
 sg13g2_antennanp ANTENNA_880 (.A(net556));
 sg13g2_antennanp ANTENNA_881 (.A(net556));
 sg13g2_antennanp ANTENNA_882 (.A(net556));
 sg13g2_antennanp ANTENNA_883 (.A(net556));
 sg13g2_antennanp ANTENNA_884 (.A(net568));
 sg13g2_antennanp ANTENNA_885 (.A(net568));
 sg13g2_antennanp ANTENNA_886 (.A(net568));
 sg13g2_antennanp ANTENNA_887 (.A(net568));
 sg13g2_antennanp ANTENNA_888 (.A(net568));
 sg13g2_antennanp ANTENNA_889 (.A(net568));
 sg13g2_antennanp ANTENNA_890 (.A(net568));
 sg13g2_antennanp ANTENNA_891 (.A(net568));
 sg13g2_antennanp ANTENNA_892 (.A(net568));
 sg13g2_antennanp ANTENNA_893 (.A(net641));
 sg13g2_antennanp ANTENNA_894 (.A(net641));
 sg13g2_antennanp ANTENNA_895 (.A(net641));
 sg13g2_antennanp ANTENNA_896 (.A(net641));
 sg13g2_antennanp ANTENNA_897 (.A(net641));
 sg13g2_antennanp ANTENNA_898 (.A(net641));
 sg13g2_antennanp ANTENNA_899 (.A(net641));
 sg13g2_antennanp ANTENNA_900 (.A(net641));
 sg13g2_antennanp ANTENNA_901 (.A(net641));
 sg13g2_antennanp ANTENNA_902 (.A(net697));
 sg13g2_antennanp ANTENNA_903 (.A(net697));
 sg13g2_antennanp ANTENNA_904 (.A(net697));
 sg13g2_antennanp ANTENNA_905 (.A(net697));
 sg13g2_antennanp ANTENNA_906 (.A(net697));
 sg13g2_antennanp ANTENNA_907 (.A(net697));
 sg13g2_antennanp ANTENNA_908 (.A(net697));
 sg13g2_antennanp ANTENNA_909 (.A(net697));
 sg13g2_antennanp ANTENNA_910 (.A(net697));
 sg13g2_antennanp ANTENNA_911 (.A(net770));
 sg13g2_antennanp ANTENNA_912 (.A(net770));
 sg13g2_antennanp ANTENNA_913 (.A(net770));
 sg13g2_antennanp ANTENNA_914 (.A(net770));
 sg13g2_antennanp ANTENNA_915 (.A(net770));
 sg13g2_antennanp ANTENNA_916 (.A(net770));
 sg13g2_antennanp ANTENNA_917 (.A(net770));
 sg13g2_antennanp ANTENNA_918 (.A(net770));
 sg13g2_antennanp ANTENNA_919 (.A(net773));
 sg13g2_antennanp ANTENNA_920 (.A(net773));
 sg13g2_antennanp ANTENNA_921 (.A(net773));
 sg13g2_antennanp ANTENNA_922 (.A(net773));
 sg13g2_antennanp ANTENNA_923 (.A(net773));
 sg13g2_antennanp ANTENNA_924 (.A(net773));
 sg13g2_antennanp ANTENNA_925 (.A(net773));
 sg13g2_antennanp ANTENNA_926 (.A(net773));
 sg13g2_antennanp ANTENNA_927 (.A(net773));
 sg13g2_antennanp ANTENNA_928 (.A(net773));
 sg13g2_antennanp ANTENNA_929 (.A(net773));
 sg13g2_antennanp ANTENNA_930 (.A(net773));
 sg13g2_antennanp ANTENNA_931 (.A(net773));
 sg13g2_antennanp ANTENNA_932 (.A(net778));
 sg13g2_antennanp ANTENNA_933 (.A(net778));
 sg13g2_antennanp ANTENNA_934 (.A(net778));
 sg13g2_antennanp ANTENNA_935 (.A(net778));
 sg13g2_antennanp ANTENNA_936 (.A(net778));
 sg13g2_antennanp ANTENNA_937 (.A(net778));
 sg13g2_antennanp ANTENNA_938 (.A(net778));
 sg13g2_antennanp ANTENNA_939 (.A(net778));
 sg13g2_antennanp ANTENNA_940 (.A(net791));
 sg13g2_antennanp ANTENNA_941 (.A(net791));
 sg13g2_antennanp ANTENNA_942 (.A(net791));
 sg13g2_antennanp ANTENNA_943 (.A(net791));
 sg13g2_antennanp ANTENNA_944 (.A(net791));
 sg13g2_antennanp ANTENNA_945 (.A(net791));
 sg13g2_antennanp ANTENNA_946 (.A(net791));
 sg13g2_antennanp ANTENNA_947 (.A(net791));
 sg13g2_antennanp ANTENNA_948 (.A(net791));
 sg13g2_antennanp ANTENNA_949 (.A(net791));
 sg13g2_antennanp ANTENNA_950 (.A(net791));
 sg13g2_antennanp ANTENNA_951 (.A(net791));
 sg13g2_antennanp ANTENNA_952 (.A(net791));
 sg13g2_antennanp ANTENNA_953 (.A(net791));
 sg13g2_antennanp ANTENNA_954 (.A(net791));
 sg13g2_antennanp ANTENNA_955 (.A(net791));
 sg13g2_antennanp ANTENNA_956 (.A(net791));
 sg13g2_antennanp ANTENNA_957 (.A(net791));
 sg13g2_antennanp ANTENNA_958 (.A(net791));
 sg13g2_antennanp ANTENNA_959 (.A(net791));
 sg13g2_antennanp ANTENNA_960 (.A(net791));
 sg13g2_antennanp ANTENNA_961 (.A(net791));
 sg13g2_antennanp ANTENNA_962 (.A(net791));
 sg13g2_antennanp ANTENNA_963 (.A(net791));
 sg13g2_antennanp ANTENNA_964 (.A(net791));
 sg13g2_antennanp ANTENNA_965 (.A(net791));
 sg13g2_antennanp ANTENNA_966 (.A(net791));
 sg13g2_antennanp ANTENNA_967 (.A(net791));
 sg13g2_antennanp ANTENNA_968 (.A(net791));
 sg13g2_antennanp ANTENNA_969 (.A(net792));
 sg13g2_antennanp ANTENNA_970 (.A(net792));
 sg13g2_antennanp ANTENNA_971 (.A(net792));
 sg13g2_antennanp ANTENNA_972 (.A(net792));
 sg13g2_antennanp ANTENNA_973 (.A(net792));
 sg13g2_antennanp ANTENNA_974 (.A(net792));
 sg13g2_antennanp ANTENNA_975 (.A(net792));
 sg13g2_antennanp ANTENNA_976 (.A(net792));
 sg13g2_antennanp ANTENNA_977 (.A(net792));
 sg13g2_antennanp ANTENNA_978 (.A(net792));
 sg13g2_antennanp ANTENNA_979 (.A(net792));
 sg13g2_antennanp ANTENNA_980 (.A(net792));
 sg13g2_antennanp ANTENNA_981 (.A(net792));
 sg13g2_antennanp ANTENNA_982 (.A(net792));
 sg13g2_antennanp ANTENNA_983 (.A(net792));
 sg13g2_antennanp ANTENNA_984 (.A(net792));
 sg13g2_antennanp ANTENNA_985 (.A(net792));
 sg13g2_antennanp ANTENNA_986 (.A(net792));
 sg13g2_antennanp ANTENNA_987 (.A(net792));
 sg13g2_antennanp ANTENNA_988 (.A(net792));
 sg13g2_antennanp ANTENNA_989 (.A(net802));
 sg13g2_antennanp ANTENNA_990 (.A(net802));
 sg13g2_antennanp ANTENNA_991 (.A(net802));
 sg13g2_antennanp ANTENNA_992 (.A(net802));
 sg13g2_antennanp ANTENNA_993 (.A(net802));
 sg13g2_antennanp ANTENNA_994 (.A(net802));
 sg13g2_antennanp ANTENNA_995 (.A(net802));
 sg13g2_antennanp ANTENNA_996 (.A(net802));
 sg13g2_antennanp ANTENNA_997 (.A(net802));
 sg13g2_antennanp ANTENNA_998 (.A(net838));
 sg13g2_antennanp ANTENNA_999 (.A(net838));
 sg13g2_antennanp ANTENNA_1000 (.A(net838));
 sg13g2_antennanp ANTENNA_1001 (.A(net838));
 sg13g2_antennanp ANTENNA_1002 (.A(net838));
 sg13g2_antennanp ANTENNA_1003 (.A(net838));
 sg13g2_antennanp ANTENNA_1004 (.A(net838));
 sg13g2_antennanp ANTENNA_1005 (.A(net838));
 sg13g2_antennanp ANTENNA_1006 (.A(net838));
 sg13g2_antennanp ANTENNA_1007 (.A(net839));
 sg13g2_antennanp ANTENNA_1008 (.A(net839));
 sg13g2_antennanp ANTENNA_1009 (.A(net839));
 sg13g2_antennanp ANTENNA_1010 (.A(net839));
 sg13g2_antennanp ANTENNA_1011 (.A(net839));
 sg13g2_antennanp ANTENNA_1012 (.A(net839));
 sg13g2_antennanp ANTENNA_1013 (.A(net839));
 sg13g2_antennanp ANTENNA_1014 (.A(net839));
 sg13g2_antennanp ANTENNA_1015 (.A(net839));
 sg13g2_antennanp ANTENNA_1016 (.A(net878));
 sg13g2_antennanp ANTENNA_1017 (.A(net878));
 sg13g2_antennanp ANTENNA_1018 (.A(net878));
 sg13g2_antennanp ANTENNA_1019 (.A(net878));
 sg13g2_antennanp ANTENNA_1020 (.A(net878));
 sg13g2_antennanp ANTENNA_1021 (.A(net878));
 sg13g2_antennanp ANTENNA_1022 (.A(net878));
 sg13g2_antennanp ANTENNA_1023 (.A(net878));
 sg13g2_antennanp ANTENNA_1024 (.A(net878));
 sg13g2_antennanp ANTENNA_1025 (.A(net878));
 sg13g2_antennanp ANTENNA_1026 (.A(net878));
 sg13g2_antennanp ANTENNA_1027 (.A(net878));
 sg13g2_antennanp ANTENNA_1028 (.A(net878));
 sg13g2_antennanp ANTENNA_1029 (.A(net878));
 sg13g2_antennanp ANTENNA_1030 (.A(net878));
 sg13g2_antennanp ANTENNA_1031 (.A(net878));
 sg13g2_antennanp ANTENNA_1032 (.A(net878));
 sg13g2_antennanp ANTENNA_1033 (.A(net878));
 sg13g2_antennanp ANTENNA_1034 (.A(net878));
 sg13g2_antennanp ANTENNA_1035 (.A(net878));
 sg13g2_antennanp ANTENNA_1036 (.A(net878));
 sg13g2_antennanp ANTENNA_1037 (.A(net878));
 sg13g2_antennanp ANTENNA_1038 (.A(net878));
 sg13g2_antennanp ANTENNA_1039 (.A(net878));
 sg13g2_antennanp ANTENNA_1040 (.A(net878));
 sg13g2_antennanp ANTENNA_1041 (.A(net878));
 sg13g2_antennanp ANTENNA_1042 (.A(net878));
 sg13g2_antennanp ANTENNA_1043 (.A(net878));
 sg13g2_antennanp ANTENNA_1044 (.A(net878));
 sg13g2_antennanp ANTENNA_1045 (.A(net878));
 sg13g2_antennanp ANTENNA_1046 (.A(net878));
 sg13g2_antennanp ANTENNA_1047 (.A(net878));
 sg13g2_antennanp ANTENNA_1048 (.A(net878));
 sg13g2_antennanp ANTENNA_1049 (.A(net878));
 sg13g2_antennanp ANTENNA_1050 (.A(net878));
 sg13g2_antennanp ANTENNA_1051 (.A(net878));
 sg13g2_antennanp ANTENNA_1052 (.A(net878));
 sg13g2_antennanp ANTENNA_1053 (.A(net878));
 sg13g2_antennanp ANTENNA_1054 (.A(net878));
 sg13g2_antennanp ANTENNA_1055 (.A(net878));
 sg13g2_antennanp ANTENNA_1056 (.A(net878));
 sg13g2_antennanp ANTENNA_1057 (.A(net878));
 sg13g2_antennanp ANTENNA_1058 (.A(net878));
 sg13g2_antennanp ANTENNA_1059 (.A(net878));
 sg13g2_antennanp ANTENNA_1060 (.A(net924));
 sg13g2_antennanp ANTENNA_1061 (.A(net924));
 sg13g2_antennanp ANTENNA_1062 (.A(net924));
 sg13g2_antennanp ANTENNA_1063 (.A(net924));
 sg13g2_antennanp ANTENNA_1064 (.A(net924));
 sg13g2_antennanp ANTENNA_1065 (.A(net924));
 sg13g2_antennanp ANTENNA_1066 (.A(net924));
 sg13g2_antennanp ANTENNA_1067 (.A(net924));
 sg13g2_antennanp ANTENNA_1068 (.A(net924));
 sg13g2_antennanp ANTENNA_1069 (.A(net925));
 sg13g2_antennanp ANTENNA_1070 (.A(net925));
 sg13g2_antennanp ANTENNA_1071 (.A(net925));
 sg13g2_antennanp ANTENNA_1072 (.A(net925));
 sg13g2_antennanp ANTENNA_1073 (.A(net925));
 sg13g2_antennanp ANTENNA_1074 (.A(net925));
 sg13g2_antennanp ANTENNA_1075 (.A(net925));
 sg13g2_antennanp ANTENNA_1076 (.A(net925));
 sg13g2_antennanp ANTENNA_1077 (.A(net925));
 sg13g2_antennanp ANTENNA_1078 (.A(net968));
 sg13g2_antennanp ANTENNA_1079 (.A(net968));
 sg13g2_antennanp ANTENNA_1080 (.A(net968));
 sg13g2_antennanp ANTENNA_1081 (.A(net968));
 sg13g2_antennanp ANTENNA_1082 (.A(net968));
 sg13g2_antennanp ANTENNA_1083 (.A(net968));
 sg13g2_antennanp ANTENNA_1084 (.A(net968));
 sg13g2_antennanp ANTENNA_1085 (.A(net968));
 sg13g2_antennanp ANTENNA_1086 (.A(net968));
 sg13g2_antennanp ANTENNA_1087 (.A(net968));
 sg13g2_antennanp ANTENNA_1088 (.A(net968));
 sg13g2_antennanp ANTENNA_1089 (.A(net968));
 sg13g2_antennanp ANTENNA_1090 (.A(net968));
 sg13g2_antennanp ANTENNA_1091 (.A(net968));
 sg13g2_antennanp ANTENNA_1092 (.A(net968));
 sg13g2_antennanp ANTENNA_1093 (.A(net968));
 sg13g2_antennanp ANTENNA_1094 (.A(net982));
 sg13g2_antennanp ANTENNA_1095 (.A(net982));
 sg13g2_antennanp ANTENNA_1096 (.A(net982));
 sg13g2_antennanp ANTENNA_1097 (.A(net982));
 sg13g2_antennanp ANTENNA_1098 (.A(net982));
 sg13g2_antennanp ANTENNA_1099 (.A(net982));
 sg13g2_antennanp ANTENNA_1100 (.A(net982));
 sg13g2_antennanp ANTENNA_1101 (.A(net982));
 sg13g2_antennanp ANTENNA_1102 (.A(net982));
 sg13g2_antennanp ANTENNA_1103 (.A(net989));
 sg13g2_antennanp ANTENNA_1104 (.A(net989));
 sg13g2_antennanp ANTENNA_1105 (.A(net989));
 sg13g2_antennanp ANTENNA_1106 (.A(net989));
 sg13g2_antennanp ANTENNA_1107 (.A(net989));
 sg13g2_antennanp ANTENNA_1108 (.A(net989));
 sg13g2_antennanp ANTENNA_1109 (.A(net989));
 sg13g2_antennanp ANTENNA_1110 (.A(net989));
 sg13g2_antennanp ANTENNA_1111 (.A(net989));
 sg13g2_antennanp ANTENNA_1112 (.A(net989));
 sg13g2_antennanp ANTENNA_1113 (.A(net989));
 sg13g2_antennanp ANTENNA_1114 (.A(net989));
 sg13g2_antennanp ANTENNA_1115 (.A(net989));
 sg13g2_antennanp ANTENNA_1116 (.A(net989));
 sg13g2_antennanp ANTENNA_1117 (.A(net990));
 sg13g2_antennanp ANTENNA_1118 (.A(net990));
 sg13g2_antennanp ANTENNA_1119 (.A(net990));
 sg13g2_antennanp ANTENNA_1120 (.A(net990));
 sg13g2_antennanp ANTENNA_1121 (.A(net990));
 sg13g2_antennanp ANTENNA_1122 (.A(net990));
 sg13g2_antennanp ANTENNA_1123 (.A(net990));
 sg13g2_antennanp ANTENNA_1124 (.A(net990));
 sg13g2_antennanp ANTENNA_1125 (.A(net990));
 sg13g2_antennanp ANTENNA_1126 (.A(net1051));
 sg13g2_antennanp ANTENNA_1127 (.A(net1051));
 sg13g2_antennanp ANTENNA_1128 (.A(net1051));
 sg13g2_antennanp ANTENNA_1129 (.A(net1051));
 sg13g2_antennanp ANTENNA_1130 (.A(net1051));
 sg13g2_antennanp ANTENNA_1131 (.A(net1051));
 sg13g2_antennanp ANTENNA_1132 (.A(net1051));
 sg13g2_antennanp ANTENNA_1133 (.A(net1051));
 sg13g2_antennanp ANTENNA_1134 (.A(net1051));
 sg13g2_antennanp ANTENNA_1135 (.A(net1054));
 sg13g2_antennanp ANTENNA_1136 (.A(net1054));
 sg13g2_antennanp ANTENNA_1137 (.A(net1054));
 sg13g2_antennanp ANTENNA_1138 (.A(net1054));
 sg13g2_antennanp ANTENNA_1139 (.A(net1054));
 sg13g2_antennanp ANTENNA_1140 (.A(net1054));
 sg13g2_antennanp ANTENNA_1141 (.A(net1054));
 sg13g2_antennanp ANTENNA_1142 (.A(net1054));
 sg13g2_antennanp ANTENNA_1143 (.A(net1099));
 sg13g2_antennanp ANTENNA_1144 (.A(net1099));
 sg13g2_antennanp ANTENNA_1145 (.A(net1099));
 sg13g2_antennanp ANTENNA_1146 (.A(net1099));
 sg13g2_antennanp ANTENNA_1147 (.A(net1099));
 sg13g2_antennanp ANTENNA_1148 (.A(net1099));
 sg13g2_antennanp ANTENNA_1149 (.A(net1099));
 sg13g2_antennanp ANTENNA_1150 (.A(net1099));
 sg13g2_antennanp ANTENNA_1151 (.A(net1099));
 sg13g2_antennanp ANTENNA_1152 (.A(net1099));
 sg13g2_antennanp ANTENNA_1153 (.A(net1099));
 sg13g2_antennanp ANTENNA_1154 (.A(net1099));
 sg13g2_antennanp ANTENNA_1155 (.A(net1099));
 sg13g2_antennanp ANTENNA_1156 (.A(net1099));
 sg13g2_antennanp ANTENNA_1157 (.A(net1099));
 sg13g2_antennanp ANTENNA_1158 (.A(net1100));
 sg13g2_antennanp ANTENNA_1159 (.A(net1100));
 sg13g2_antennanp ANTENNA_1160 (.A(net1100));
 sg13g2_antennanp ANTENNA_1161 (.A(net1100));
 sg13g2_antennanp ANTENNA_1162 (.A(net1100));
 sg13g2_antennanp ANTENNA_1163 (.A(net1100));
 sg13g2_antennanp ANTENNA_1164 (.A(net1100));
 sg13g2_antennanp ANTENNA_1165 (.A(net1100));
 sg13g2_antennanp ANTENNA_1166 (.A(net1100));
 sg13g2_antennanp ANTENNA_1167 (.A(net1100));
 sg13g2_antennanp ANTENNA_1168 (.A(net1100));
 sg13g2_antennanp ANTENNA_1169 (.A(net1100));
 sg13g2_antennanp ANTENNA_1170 (.A(net1100));
 sg13g2_antennanp ANTENNA_1171 (.A(net1100));
 sg13g2_antennanp ANTENNA_1172 (.A(net1100));
 sg13g2_antennanp ANTENNA_1173 (.A(net1100));
 sg13g2_antennanp ANTENNA_1174 (.A(net1104));
 sg13g2_antennanp ANTENNA_1175 (.A(net1104));
 sg13g2_antennanp ANTENNA_1176 (.A(net1104));
 sg13g2_antennanp ANTENNA_1177 (.A(net1104));
 sg13g2_antennanp ANTENNA_1178 (.A(net1104));
 sg13g2_antennanp ANTENNA_1179 (.A(net1104));
 sg13g2_antennanp ANTENNA_1180 (.A(net1104));
 sg13g2_antennanp ANTENNA_1181 (.A(net1104));
 sg13g2_antennanp ANTENNA_1182 (.A(net1104));
 sg13g2_antennanp ANTENNA_1183 (.A(net1192));
 sg13g2_antennanp ANTENNA_1184 (.A(net1192));
 sg13g2_antennanp ANTENNA_1185 (.A(net1192));
 sg13g2_antennanp ANTENNA_1186 (.A(net1192));
 sg13g2_antennanp ANTENNA_1187 (.A(net1192));
 sg13g2_antennanp ANTENNA_1188 (.A(net1192));
 sg13g2_antennanp ANTENNA_1189 (.A(net1192));
 sg13g2_antennanp ANTENNA_1190 (.A(net1192));
 sg13g2_antennanp ANTENNA_1191 (.A(net1192));
 sg13g2_antennanp ANTENNA_1192 (.A(net1192));
 sg13g2_antennanp ANTENNA_1193 (.A(net1192));
 sg13g2_antennanp ANTENNA_1194 (.A(net1192));
 sg13g2_antennanp ANTENNA_1195 (.A(net1192));
 sg13g2_antennanp ANTENNA_1196 (.A(net1192));
 sg13g2_antennanp ANTENNA_1197 (.A(net1192));
 sg13g2_antennanp ANTENNA_1198 (.A(net1192));
 sg13g2_antennanp ANTENNA_1199 (.A(net1192));
 sg13g2_antennanp ANTENNA_1200 (.A(net1192));
 sg13g2_antennanp ANTENNA_1201 (.A(net1192));
 sg13g2_antennanp ANTENNA_1202 (.A(net1192));
 sg13g2_antennanp ANTENNA_1203 (.A(net1192));
 sg13g2_antennanp ANTENNA_1204 (.A(net1192));
 sg13g2_antennanp ANTENNA_1205 (.A(net1192));
 sg13g2_antennanp ANTENNA_1206 (.A(net1192));
 sg13g2_antennanp ANTENNA_1207 (.A(net1192));
 sg13g2_antennanp ANTENNA_1208 (.A(net1192));
 sg13g2_antennanp ANTENNA_1209 (.A(net1192));
 sg13g2_antennanp ANTENNA_1210 (.A(net1192));
 sg13g2_antennanp ANTENNA_1211 (.A(net1192));
 sg13g2_antennanp ANTENNA_1212 (.A(net1192));
 sg13g2_antennanp ANTENNA_1213 (.A(net1192));
 sg13g2_antennanp ANTENNA_1214 (.A(net1192));
 sg13g2_antennanp ANTENNA_1215 (.A(net1192));
 sg13g2_antennanp ANTENNA_1216 (.A(net1192));
 sg13g2_antennanp ANTENNA_1217 (.A(net1193));
 sg13g2_antennanp ANTENNA_1218 (.A(net1193));
 sg13g2_antennanp ANTENNA_1219 (.A(net1193));
 sg13g2_antennanp ANTENNA_1220 (.A(net1193));
 sg13g2_antennanp ANTENNA_1221 (.A(net1193));
 sg13g2_antennanp ANTENNA_1222 (.A(net1193));
 sg13g2_antennanp ANTENNA_1223 (.A(net1193));
 sg13g2_antennanp ANTENNA_1224 (.A(net1193));
 sg13g2_antennanp ANTENNA_1225 (.A(net1193));
 sg13g2_antennanp ANTENNA_1226 (.A(net1273));
 sg13g2_antennanp ANTENNA_1227 (.A(net1273));
 sg13g2_antennanp ANTENNA_1228 (.A(net1273));
 sg13g2_antennanp ANTENNA_1229 (.A(net1273));
 sg13g2_antennanp ANTENNA_1230 (.A(net1273));
 sg13g2_antennanp ANTENNA_1231 (.A(net1273));
 sg13g2_antennanp ANTENNA_1232 (.A(net1273));
 sg13g2_antennanp ANTENNA_1233 (.A(net1273));
 sg13g2_antennanp ANTENNA_1234 (.A(net1273));
 sg13g2_antennanp ANTENNA_1235 (.A(net1273));
 sg13g2_antennanp ANTENNA_1236 (.A(net1273));
 sg13g2_antennanp ANTENNA_1237 (.A(net1273));
 sg13g2_antennanp ANTENNA_1238 (.A(net1273));
 sg13g2_antennanp ANTENNA_1239 (.A(net1273));
 sg13g2_antennanp ANTENNA_1240 (.A(net1273));
 sg13g2_antennanp ANTENNA_1241 (.A(net1273));
 sg13g2_antennanp ANTENNA_1242 (.A(net1273));
 sg13g2_antennanp ANTENNA_1243 (.A(net1273));
 sg13g2_antennanp ANTENNA_1244 (.A(net1273));
 sg13g2_antennanp ANTENNA_1245 (.A(net1273));
 sg13g2_antennanp ANTENNA_1246 (.A(net1273));
 sg13g2_antennanp ANTENNA_1247 (.A(net1273));
 sg13g2_antennanp ANTENNA_1248 (.A(net1273));
 sg13g2_antennanp ANTENNA_1249 (.A(net1273));
 sg13g2_antennanp ANTENNA_1250 (.A(net1273));
 sg13g2_antennanp ANTENNA_1251 (.A(net1273));
 sg13g2_antennanp ANTENNA_1252 (.A(net1273));
 sg13g2_antennanp ANTENNA_1253 (.A(net1273));
 sg13g2_antennanp ANTENNA_1254 (.A(net1273));
 sg13g2_antennanp ANTENNA_1255 (.A(net1276));
 sg13g2_antennanp ANTENNA_1256 (.A(net1276));
 sg13g2_antennanp ANTENNA_1257 (.A(net1276));
 sg13g2_antennanp ANTENNA_1258 (.A(net1276));
 sg13g2_antennanp ANTENNA_1259 (.A(net1276));
 sg13g2_antennanp ANTENNA_1260 (.A(net1276));
 sg13g2_antennanp ANTENNA_1261 (.A(net1276));
 sg13g2_antennanp ANTENNA_1262 (.A(net1276));
 sg13g2_antennanp ANTENNA_1263 (.A(net1276));
 sg13g2_antennanp ANTENNA_1264 (.A(net1276));
 sg13g2_antennanp ANTENNA_1265 (.A(net1276));
 sg13g2_antennanp ANTENNA_1266 (.A(net1276));
 sg13g2_antennanp ANTENNA_1267 (.A(net1276));
 sg13g2_antennanp ANTENNA_1268 (.A(net1276));
 sg13g2_antennanp ANTENNA_1269 (.A(net1276));
 sg13g2_antennanp ANTENNA_1270 (.A(net1276));
 sg13g2_antennanp ANTENNA_1271 (.A(_00017_));
 sg13g2_antennanp ANTENNA_1272 (.A(_00017_));
 sg13g2_antennanp ANTENNA_1273 (.A(_00017_));
 sg13g2_antennanp ANTENNA_1274 (.A(_00017_));
 sg13g2_antennanp ANTENNA_1275 (.A(_02490_));
 sg13g2_antennanp ANTENNA_1276 (.A(_03341_));
 sg13g2_antennanp ANTENNA_1277 (.A(_03444_));
 sg13g2_antennanp ANTENNA_1278 (.A(_03444_));
 sg13g2_antennanp ANTENNA_1279 (.A(_03444_));
 sg13g2_antennanp ANTENNA_1280 (.A(_03621_));
 sg13g2_antennanp ANTENNA_1281 (.A(_03621_));
 sg13g2_antennanp ANTENNA_1282 (.A(_03621_));
 sg13g2_antennanp ANTENNA_1283 (.A(_03621_));
 sg13g2_antennanp ANTENNA_1284 (.A(_03621_));
 sg13g2_antennanp ANTENNA_1285 (.A(_03621_));
 sg13g2_antennanp ANTENNA_1286 (.A(_03621_));
 sg13g2_antennanp ANTENNA_1287 (.A(_03621_));
 sg13g2_antennanp ANTENNA_1288 (.A(_03843_));
 sg13g2_antennanp ANTENNA_1289 (.A(_03843_));
 sg13g2_antennanp ANTENNA_1290 (.A(_03843_));
 sg13g2_antennanp ANTENNA_1291 (.A(_03843_));
 sg13g2_antennanp ANTENNA_1292 (.A(_03875_));
 sg13g2_antennanp ANTENNA_1293 (.A(_03995_));
 sg13g2_antennanp ANTENNA_1294 (.A(_03995_));
 sg13g2_antennanp ANTENNA_1295 (.A(_03995_));
 sg13g2_antennanp ANTENNA_1296 (.A(_03995_));
 sg13g2_antennanp ANTENNA_1297 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1298 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1299 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1300 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1301 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1302 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1303 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1304 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1305 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1306 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1307 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1308 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1309 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1310 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1311 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1312 (.A(_04431_));
 sg13g2_antennanp ANTENNA_1313 (.A(_05432_));
 sg13g2_antennanp ANTENNA_1314 (.A(_05432_));
 sg13g2_antennanp ANTENNA_1315 (.A(_05432_));
 sg13g2_antennanp ANTENNA_1316 (.A(_05441_));
 sg13g2_antennanp ANTENNA_1317 (.A(_05441_));
 sg13g2_antennanp ANTENNA_1318 (.A(_05441_));
 sg13g2_antennanp ANTENNA_1319 (.A(_05446_));
 sg13g2_antennanp ANTENNA_1320 (.A(_05446_));
 sg13g2_antennanp ANTENNA_1321 (.A(_05446_));
 sg13g2_antennanp ANTENNA_1322 (.A(_05446_));
 sg13g2_antennanp ANTENNA_1323 (.A(_05449_));
 sg13g2_antennanp ANTENNA_1324 (.A(_05449_));
 sg13g2_antennanp ANTENNA_1325 (.A(_05449_));
 sg13g2_antennanp ANTENNA_1326 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1327 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1328 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1329 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1330 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1331 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1332 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1333 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1334 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1335 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1336 (.A(_05457_));
 sg13g2_antennanp ANTENNA_1337 (.A(_05457_));
 sg13g2_antennanp ANTENNA_1338 (.A(_05457_));
 sg13g2_antennanp ANTENNA_1339 (.A(_05457_));
 sg13g2_antennanp ANTENNA_1340 (.A(_05457_));
 sg13g2_antennanp ANTENNA_1341 (.A(_05457_));
 sg13g2_antennanp ANTENNA_1342 (.A(_05463_));
 sg13g2_antennanp ANTENNA_1343 (.A(_05463_));
 sg13g2_antennanp ANTENNA_1344 (.A(_05463_));
 sg13g2_antennanp ANTENNA_1345 (.A(_05463_));
 sg13g2_antennanp ANTENNA_1346 (.A(_05463_));
 sg13g2_antennanp ANTENNA_1347 (.A(_05463_));
 sg13g2_antennanp ANTENNA_1348 (.A(_05467_));
 sg13g2_antennanp ANTENNA_1349 (.A(_05467_));
 sg13g2_antennanp ANTENNA_1350 (.A(_05467_));
 sg13g2_antennanp ANTENNA_1351 (.A(_05467_));
 sg13g2_antennanp ANTENNA_1352 (.A(_05467_));
 sg13g2_antennanp ANTENNA_1353 (.A(_05467_));
 sg13g2_antennanp ANTENNA_1354 (.A(_05471_));
 sg13g2_antennanp ANTENNA_1355 (.A(_05471_));
 sg13g2_antennanp ANTENNA_1356 (.A(_05471_));
 sg13g2_antennanp ANTENNA_1357 (.A(_05471_));
 sg13g2_antennanp ANTENNA_1358 (.A(_05471_));
 sg13g2_antennanp ANTENNA_1359 (.A(_05471_));
 sg13g2_antennanp ANTENNA_1360 (.A(_05471_));
 sg13g2_antennanp ANTENNA_1361 (.A(_05471_));
 sg13g2_antennanp ANTENNA_1362 (.A(_05471_));
 sg13g2_antennanp ANTENNA_1363 (.A(_05476_));
 sg13g2_antennanp ANTENNA_1364 (.A(_05476_));
 sg13g2_antennanp ANTENNA_1365 (.A(_05498_));
 sg13g2_antennanp ANTENNA_1366 (.A(_05498_));
 sg13g2_antennanp ANTENNA_1367 (.A(_06148_));
 sg13g2_antennanp ANTENNA_1368 (.A(_06148_));
 sg13g2_antennanp ANTENNA_1369 (.A(_06148_));
 sg13g2_antennanp ANTENNA_1370 (.A(_06148_));
 sg13g2_antennanp ANTENNA_1371 (.A(_06148_));
 sg13g2_antennanp ANTENNA_1372 (.A(_06148_));
 sg13g2_antennanp ANTENNA_1373 (.A(_06148_));
 sg13g2_antennanp ANTENNA_1374 (.A(_06148_));
 sg13g2_antennanp ANTENNA_1375 (.A(_06148_));
 sg13g2_antennanp ANTENNA_1376 (.A(_06171_));
 sg13g2_antennanp ANTENNA_1377 (.A(_06189_));
 sg13g2_antennanp ANTENNA_1378 (.A(_06253_));
 sg13g2_antennanp ANTENNA_1379 (.A(_06253_));
 sg13g2_antennanp ANTENNA_1380 (.A(_06255_));
 sg13g2_antennanp ANTENNA_1381 (.A(_06268_));
 sg13g2_antennanp ANTENNA_1382 (.A(_06293_));
 sg13g2_antennanp ANTENNA_1383 (.A(_06298_));
 sg13g2_antennanp ANTENNA_1384 (.A(_06311_));
 sg13g2_antennanp ANTENNA_1385 (.A(_06318_));
 sg13g2_antennanp ANTENNA_1386 (.A(_06329_));
 sg13g2_antennanp ANTENNA_1387 (.A(_06393_));
 sg13g2_antennanp ANTENNA_1388 (.A(_06393_));
 sg13g2_antennanp ANTENNA_1389 (.A(_06393_));
 sg13g2_antennanp ANTENNA_1390 (.A(_06393_));
 sg13g2_antennanp ANTENNA_1391 (.A(_06416_));
 sg13g2_antennanp ANTENNA_1392 (.A(_06460_));
 sg13g2_antennanp ANTENNA_1393 (.A(_06460_));
 sg13g2_antennanp ANTENNA_1394 (.A(_06493_));
 sg13g2_antennanp ANTENNA_1395 (.A(_06493_));
 sg13g2_antennanp ANTENNA_1396 (.A(_06516_));
 sg13g2_antennanp ANTENNA_1397 (.A(_06516_));
 sg13g2_antennanp ANTENNA_1398 (.A(_06520_));
 sg13g2_antennanp ANTENNA_1399 (.A(_06559_));
 sg13g2_antennanp ANTENNA_1400 (.A(_06560_));
 sg13g2_antennanp ANTENNA_1401 (.A(_06595_));
 sg13g2_antennanp ANTENNA_1402 (.A(_06601_));
 sg13g2_antennanp ANTENNA_1403 (.A(_06616_));
 sg13g2_antennanp ANTENNA_1404 (.A(_06618_));
 sg13g2_antennanp ANTENNA_1405 (.A(_06620_));
 sg13g2_antennanp ANTENNA_1406 (.A(_06658_));
 sg13g2_antennanp ANTENNA_1407 (.A(_06694_));
 sg13g2_antennanp ANTENNA_1408 (.A(_06719_));
 sg13g2_antennanp ANTENNA_1409 (.A(_06757_));
 sg13g2_antennanp ANTENNA_1410 (.A(_06772_));
 sg13g2_antennanp ANTENNA_1411 (.A(_06772_));
 sg13g2_antennanp ANTENNA_1412 (.A(_06793_));
 sg13g2_antennanp ANTENNA_1413 (.A(_06793_));
 sg13g2_antennanp ANTENNA_1414 (.A(_06799_));
 sg13g2_antennanp ANTENNA_1415 (.A(_06814_));
 sg13g2_antennanp ANTENNA_1416 (.A(_06814_));
 sg13g2_antennanp ANTENNA_1417 (.A(_06818_));
 sg13g2_antennanp ANTENNA_1418 (.A(_06856_));
 sg13g2_antennanp ANTENNA_1419 (.A(_06870_));
 sg13g2_antennanp ANTENNA_1420 (.A(_06870_));
 sg13g2_antennanp ANTENNA_1421 (.A(_06871_));
 sg13g2_antennanp ANTENNA_1422 (.A(_06871_));
 sg13g2_antennanp ANTENNA_1423 (.A(_06913_));
 sg13g2_antennanp ANTENNA_1424 (.A(_06917_));
 sg13g2_antennanp ANTENNA_1425 (.A(_06955_));
 sg13g2_antennanp ANTENNA_1426 (.A(_06975_));
 sg13g2_antennanp ANTENNA_1427 (.A(_06991_));
 sg13g2_antennanp ANTENNA_1428 (.A(_06991_));
 sg13g2_antennanp ANTENNA_1429 (.A(_07012_));
 sg13g2_antennanp ANTENNA_1430 (.A(_07012_));
 sg13g2_antennanp ANTENNA_1431 (.A(_07016_));
 sg13g2_antennanp ANTENNA_1432 (.A(_07054_));
 sg13g2_antennanp ANTENNA_1433 (.A(_07054_));
 sg13g2_antennanp ANTENNA_1434 (.A(_07074_));
 sg13g2_antennanp ANTENNA_1435 (.A(_07074_));
 sg13g2_antennanp ANTENNA_1436 (.A(_07090_));
 sg13g2_antennanp ANTENNA_1437 (.A(_07105_));
 sg13g2_antennanp ANTENNA_1438 (.A(_07335_));
 sg13g2_antennanp ANTENNA_1439 (.A(_09194_));
 sg13g2_antennanp ANTENNA_1440 (.A(_09194_));
 sg13g2_antennanp ANTENNA_1441 (.A(_09194_));
 sg13g2_antennanp ANTENNA_1442 (.A(_09194_));
 sg13g2_antennanp ANTENNA_1443 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1444 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1445 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1446 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1447 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1448 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1449 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1450 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1451 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1452 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1453 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1454 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1455 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1456 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1457 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1458 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1459 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1460 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1461 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1462 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1463 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1464 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1465 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1466 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1467 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1468 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1469 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1470 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1471 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1472 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1473 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1474 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1475 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1476 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1477 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1478 (.A(_09345_));
 sg13g2_antennanp ANTENNA_1479 (.A(_09418_));
 sg13g2_antennanp ANTENNA_1480 (.A(_09418_));
 sg13g2_antennanp ANTENNA_1481 (.A(_09418_));
 sg13g2_antennanp ANTENNA_1482 (.A(_09418_));
 sg13g2_antennanp ANTENNA_1483 (.A(_09418_));
 sg13g2_antennanp ANTENNA_1484 (.A(_09418_));
 sg13g2_antennanp ANTENNA_1485 (.A(_09418_));
 sg13g2_antennanp ANTENNA_1486 (.A(_09418_));
 sg13g2_antennanp ANTENNA_1487 (.A(_09418_));
 sg13g2_antennanp ANTENNA_1488 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1489 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1490 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1491 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1492 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1493 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1494 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1495 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1496 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1497 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1498 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1499 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1500 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1501 (.A(_09906_));
 sg13g2_antennanp ANTENNA_1502 (.A(_09928_));
 sg13g2_antennanp ANTENNA_1503 (.A(_09928_));
 sg13g2_antennanp ANTENNA_1504 (.A(_09928_));
 sg13g2_antennanp ANTENNA_1505 (.A(_09928_));
 sg13g2_antennanp ANTENNA_1506 (.A(_09928_));
 sg13g2_antennanp ANTENNA_1507 (.A(_09929_));
 sg13g2_antennanp ANTENNA_1508 (.A(_09929_));
 sg13g2_antennanp ANTENNA_1509 (.A(_09929_));
 sg13g2_antennanp ANTENNA_1510 (.A(_09929_));
 sg13g2_antennanp ANTENNA_1511 (.A(_09930_));
 sg13g2_antennanp ANTENNA_1512 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1513 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1514 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1515 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1516 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1517 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1518 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1519 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1520 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1521 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1522 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1523 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1524 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1525 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1526 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1527 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1528 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1529 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1530 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1531 (.A(_09935_));
 sg13g2_antennanp ANTENNA_1532 (.A(_09986_));
 sg13g2_antennanp ANTENNA_1533 (.A(_09986_));
 sg13g2_antennanp ANTENNA_1534 (.A(_09986_));
 sg13g2_antennanp ANTENNA_1535 (.A(_09986_));
 sg13g2_antennanp ANTENNA_1536 (.A(_09986_));
 sg13g2_antennanp ANTENNA_1537 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1538 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1539 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1540 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1541 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1542 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1543 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1544 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1545 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1546 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1547 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1548 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1549 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1550 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1551 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1552 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1553 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1554 (.A(_10046_));
 sg13g2_antennanp ANTENNA_1555 (.A(_10048_));
 sg13g2_antennanp ANTENNA_1556 (.A(_10051_));
 sg13g2_antennanp ANTENNA_1557 (.A(_10053_));
 sg13g2_antennanp ANTENNA_1558 (.A(_10071_));
 sg13g2_antennanp ANTENNA_1559 (.A(_10071_));
 sg13g2_antennanp ANTENNA_1560 (.A(_10071_));
 sg13g2_antennanp ANTENNA_1561 (.A(_10071_));
 sg13g2_antennanp ANTENNA_1562 (.A(_10071_));
 sg13g2_antennanp ANTENNA_1563 (.A(_10071_));
 sg13g2_antennanp ANTENNA_1564 (.A(_10071_));
 sg13g2_antennanp ANTENNA_1565 (.A(_10071_));
 sg13g2_antennanp ANTENNA_1566 (.A(_10071_));
 sg13g2_antennanp ANTENNA_1567 (.A(_10083_));
 sg13g2_antennanp ANTENNA_1568 (.A(_10091_));
 sg13g2_antennanp ANTENNA_1569 (.A(_10091_));
 sg13g2_antennanp ANTENNA_1570 (.A(_10092_));
 sg13g2_antennanp ANTENNA_1571 (.A(_10092_));
 sg13g2_antennanp ANTENNA_1572 (.A(_10092_));
 sg13g2_antennanp ANTENNA_1573 (.A(_10101_));
 sg13g2_antennanp ANTENNA_1574 (.A(_10101_));
 sg13g2_antennanp ANTENNA_1575 (.A(_10106_));
 sg13g2_antennanp ANTENNA_1576 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1577 (.A(_10121_));
 sg13g2_antennanp ANTENNA_1578 (.A(_10131_));
 sg13g2_antennanp ANTENNA_1579 (.A(_10136_));
 sg13g2_antennanp ANTENNA_1580 (.A(_10140_));
 sg13g2_antennanp ANTENNA_1581 (.A(_10226_));
 sg13g2_antennanp ANTENNA_1582 (.A(_10226_));
 sg13g2_antennanp ANTENNA_1583 (.A(_10226_));
 sg13g2_antennanp ANTENNA_1584 (.A(_10235_));
 sg13g2_antennanp ANTENNA_1585 (.A(_10235_));
 sg13g2_antennanp ANTENNA_1586 (.A(_10235_));
 sg13g2_antennanp ANTENNA_1587 (.A(_10235_));
 sg13g2_antennanp ANTENNA_1588 (.A(_10236_));
 sg13g2_antennanp ANTENNA_1589 (.A(_10236_));
 sg13g2_antennanp ANTENNA_1590 (.A(_10236_));
 sg13g2_antennanp ANTENNA_1591 (.A(_10236_));
 sg13g2_antennanp ANTENNA_1592 (.A(_10236_));
 sg13g2_antennanp ANTENNA_1593 (.A(_10236_));
 sg13g2_antennanp ANTENNA_1594 (.A(_10236_));
 sg13g2_antennanp ANTENNA_1595 (.A(_10243_));
 sg13g2_antennanp ANTENNA_1596 (.A(_10243_));
 sg13g2_antennanp ANTENNA_1597 (.A(_10243_));
 sg13g2_antennanp ANTENNA_1598 (.A(_10243_));
 sg13g2_antennanp ANTENNA_1599 (.A(_10243_));
 sg13g2_antennanp ANTENNA_1600 (.A(_10243_));
 sg13g2_antennanp ANTENNA_1601 (.A(_10256_));
 sg13g2_antennanp ANTENNA_1602 (.A(_10256_));
 sg13g2_antennanp ANTENNA_1603 (.A(_10256_));
 sg13g2_antennanp ANTENNA_1604 (.A(_10256_));
 sg13g2_antennanp ANTENNA_1605 (.A(_10256_));
 sg13g2_antennanp ANTENNA_1606 (.A(_10287_));
 sg13g2_antennanp ANTENNA_1607 (.A(_10287_));
 sg13g2_antennanp ANTENNA_1608 (.A(_10287_));
 sg13g2_antennanp ANTENNA_1609 (.A(_10287_));
 sg13g2_antennanp ANTENNA_1610 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1611 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1612 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1613 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1614 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1615 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1616 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1617 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1618 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1619 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1620 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1621 (.A(_10295_));
 sg13g2_antennanp ANTENNA_1622 (.A(_10296_));
 sg13g2_antennanp ANTENNA_1623 (.A(_10296_));
 sg13g2_antennanp ANTENNA_1624 (.A(_10296_));
 sg13g2_antennanp ANTENNA_1625 (.A(_10325_));
 sg13g2_antennanp ANTENNA_1626 (.A(_10325_));
 sg13g2_antennanp ANTENNA_1627 (.A(_10325_));
 sg13g2_antennanp ANTENNA_1628 (.A(_10325_));
 sg13g2_antennanp ANTENNA_1629 (.A(_10325_));
 sg13g2_antennanp ANTENNA_1630 (.A(_10325_));
 sg13g2_antennanp ANTENNA_1631 (.A(_10325_));
 sg13g2_antennanp ANTENNA_1632 (.A(_10349_));
 sg13g2_antennanp ANTENNA_1633 (.A(_10349_));
 sg13g2_antennanp ANTENNA_1634 (.A(_10349_));
 sg13g2_antennanp ANTENNA_1635 (.A(_10349_));
 sg13g2_antennanp ANTENNA_1636 (.A(_10350_));
 sg13g2_antennanp ANTENNA_1637 (.A(_10350_));
 sg13g2_antennanp ANTENNA_1638 (.A(_10350_));
 sg13g2_antennanp ANTENNA_1639 (.A(_10350_));
 sg13g2_antennanp ANTENNA_1640 (.A(_10350_));
 sg13g2_antennanp ANTENNA_1641 (.A(_10350_));
 sg13g2_antennanp ANTENNA_1642 (.A(_10350_));
 sg13g2_antennanp ANTENNA_1643 (.A(_10350_));
 sg13g2_antennanp ANTENNA_1644 (.A(_10350_));
 sg13g2_antennanp ANTENNA_1645 (.A(_10397_));
 sg13g2_antennanp ANTENNA_1646 (.A(_10397_));
 sg13g2_antennanp ANTENNA_1647 (.A(_10397_));
 sg13g2_antennanp ANTENNA_1648 (.A(_10397_));
 sg13g2_antennanp ANTENNA_1649 (.A(_10397_));
 sg13g2_antennanp ANTENNA_1650 (.A(_10397_));
 sg13g2_antennanp ANTENNA_1651 (.A(_10397_));
 sg13g2_antennanp ANTENNA_1652 (.A(_10397_));
 sg13g2_antennanp ANTENNA_1653 (.A(_10397_));
 sg13g2_antennanp ANTENNA_1654 (.A(_10415_));
 sg13g2_antennanp ANTENNA_1655 (.A(_10415_));
 sg13g2_antennanp ANTENNA_1656 (.A(_10415_));
 sg13g2_antennanp ANTENNA_1657 (.A(_10415_));
 sg13g2_antennanp ANTENNA_1658 (.A(_10415_));
 sg13g2_antennanp ANTENNA_1659 (.A(_10415_));
 sg13g2_antennanp ANTENNA_1660 (.A(_10415_));
 sg13g2_antennanp ANTENNA_1661 (.A(_10415_));
 sg13g2_antennanp ANTENNA_1662 (.A(_10415_));
 sg13g2_antennanp ANTENNA_1663 (.A(_10422_));
 sg13g2_antennanp ANTENNA_1664 (.A(_10422_));
 sg13g2_antennanp ANTENNA_1665 (.A(_10422_));
 sg13g2_antennanp ANTENNA_1666 (.A(_10422_));
 sg13g2_antennanp ANTENNA_1667 (.A(_10422_));
 sg13g2_antennanp ANTENNA_1668 (.A(_10422_));
 sg13g2_antennanp ANTENNA_1669 (.A(_10422_));
 sg13g2_antennanp ANTENNA_1670 (.A(_10422_));
 sg13g2_antennanp ANTENNA_1671 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1672 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1673 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1674 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1675 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1676 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1677 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1678 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1679 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1680 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1681 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1682 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1683 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1684 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1685 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1686 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1687 (.A(_10444_));
 sg13g2_antennanp ANTENNA_1688 (.A(_10468_));
 sg13g2_antennanp ANTENNA_1689 (.A(_10468_));
 sg13g2_antennanp ANTENNA_1690 (.A(_10468_));
 sg13g2_antennanp ANTENNA_1691 (.A(_10468_));
 sg13g2_antennanp ANTENNA_1692 (.A(_10468_));
 sg13g2_antennanp ANTENNA_1693 (.A(_10468_));
 sg13g2_antennanp ANTENNA_1694 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1695 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1696 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1697 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1698 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1699 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1700 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1701 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1702 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1703 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1704 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1705 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1706 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1707 (.A(_10513_));
 sg13g2_antennanp ANTENNA_1708 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1709 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1710 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1711 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1712 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1713 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1714 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1715 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1716 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1717 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1718 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1719 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1720 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1721 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1722 (.A(_10564_));
 sg13g2_antennanp ANTENNA_1723 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1724 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1725 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1726 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1727 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1728 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1729 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1730 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1731 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1732 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1733 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1734 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1735 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1736 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1737 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1738 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1739 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1740 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1741 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1742 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1743 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1744 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1745 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1746 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1747 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1748 (.A(_10586_));
 sg13g2_antennanp ANTENNA_1749 (.A(_10587_));
 sg13g2_antennanp ANTENNA_1750 (.A(_10587_));
 sg13g2_antennanp ANTENNA_1751 (.A(_10587_));
 sg13g2_antennanp ANTENNA_1752 (.A(_10587_));
 sg13g2_antennanp ANTENNA_1753 (.A(_10632_));
 sg13g2_antennanp ANTENNA_1754 (.A(_10632_));
 sg13g2_antennanp ANTENNA_1755 (.A(_10632_));
 sg13g2_antennanp ANTENNA_1756 (.A(_10632_));
 sg13g2_antennanp ANTENNA_1757 (.A(_10632_));
 sg13g2_antennanp ANTENNA_1758 (.A(_10632_));
 sg13g2_antennanp ANTENNA_1759 (.A(_10632_));
 sg13g2_antennanp ANTENNA_1760 (.A(_10633_));
 sg13g2_antennanp ANTENNA_1761 (.A(_10633_));
 sg13g2_antennanp ANTENNA_1762 (.A(_10633_));
 sg13g2_antennanp ANTENNA_1763 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1764 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1765 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1766 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1767 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1768 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1769 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1770 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1771 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1772 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1773 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1774 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1775 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1776 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1777 (.A(_10656_));
 sg13g2_antennanp ANTENNA_1778 (.A(_10679_));
 sg13g2_antennanp ANTENNA_1779 (.A(_10679_));
 sg13g2_antennanp ANTENNA_1780 (.A(_10679_));
 sg13g2_antennanp ANTENNA_1781 (.A(_10679_));
 sg13g2_antennanp ANTENNA_1782 (.A(_10679_));
 sg13g2_antennanp ANTENNA_1783 (.A(_10679_));
 sg13g2_antennanp ANTENNA_1784 (.A(_10679_));
 sg13g2_antennanp ANTENNA_1785 (.A(_10679_));
 sg13g2_antennanp ANTENNA_1786 (.A(_11947_));
 sg13g2_antennanp ANTENNA_1787 (.A(_11947_));
 sg13g2_antennanp ANTENNA_1788 (.A(_11947_));
 sg13g2_antennanp ANTENNA_1789 (.A(_11947_));
 sg13g2_antennanp ANTENNA_1790 (.A(_12437_));
 sg13g2_antennanp ANTENNA_1791 (.A(_12437_));
 sg13g2_antennanp ANTENNA_1792 (.A(_12437_));
 sg13g2_antennanp ANTENNA_1793 (.A(_12630_));
 sg13g2_antennanp ANTENNA_1794 (.A(_12630_));
 sg13g2_antennanp ANTENNA_1795 (.A(_12630_));
 sg13g2_antennanp ANTENNA_1796 (.A(_12653_));
 sg13g2_antennanp ANTENNA_1797 (.A(_12653_));
 sg13g2_antennanp ANTENNA_1798 (.A(_12653_));
 sg13g2_antennanp ANTENNA_1799 (.A(_12653_));
 sg13g2_antennanp ANTENNA_1800 (.A(_12653_));
 sg13g2_antennanp ANTENNA_1801 (.A(_12653_));
 sg13g2_antennanp ANTENNA_1802 (.A(_12653_));
 sg13g2_antennanp ANTENNA_1803 (.A(_12653_));
 sg13g2_antennanp ANTENNA_1804 (.A(clk));
 sg13g2_antennanp ANTENNA_1805 (.A(clk));
 sg13g2_antennanp ANTENNA_1806 (.A(\mem.data_in[1] ));
 sg13g2_antennanp ANTENNA_1807 (.A(\mem.io_data_out[0] ));
 sg13g2_antennanp ANTENNA_1808 (.A(\mem.io_data_out[0] ));
 sg13g2_antennanp ANTENNA_1809 (.A(\mem.io_data_out[3] ));
 sg13g2_antennanp ANTENNA_1810 (.A(\mem.io_data_out[3] ));
 sg13g2_antennanp ANTENNA_1811 (.A(\mem.io_data_out[4] ));
 sg13g2_antennanp ANTENNA_1812 (.A(\mem.io_data_out[4] ));
 sg13g2_antennanp ANTENNA_1813 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_1814 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_1815 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_1816 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_1817 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_1818 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_1819 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_1820 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_1821 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_1822 (.A(net1));
 sg13g2_antennanp ANTENNA_1823 (.A(net1));
 sg13g2_antennanp ANTENNA_1824 (.A(net1));
 sg13g2_antennanp ANTENNA_1825 (.A(net2));
 sg13g2_antennanp ANTENNA_1826 (.A(net4));
 sg13g2_antennanp ANTENNA_1827 (.A(net464));
 sg13g2_antennanp ANTENNA_1828 (.A(net464));
 sg13g2_antennanp ANTENNA_1829 (.A(net464));
 sg13g2_antennanp ANTENNA_1830 (.A(net464));
 sg13g2_antennanp ANTENNA_1831 (.A(net464));
 sg13g2_antennanp ANTENNA_1832 (.A(net464));
 sg13g2_antennanp ANTENNA_1833 (.A(net464));
 sg13g2_antennanp ANTENNA_1834 (.A(net464));
 sg13g2_antennanp ANTENNA_1835 (.A(net464));
 sg13g2_antennanp ANTENNA_1836 (.A(net528));
 sg13g2_antennanp ANTENNA_1837 (.A(net528));
 sg13g2_antennanp ANTENNA_1838 (.A(net528));
 sg13g2_antennanp ANTENNA_1839 (.A(net528));
 sg13g2_antennanp ANTENNA_1840 (.A(net528));
 sg13g2_antennanp ANTENNA_1841 (.A(net528));
 sg13g2_antennanp ANTENNA_1842 (.A(net528));
 sg13g2_antennanp ANTENNA_1843 (.A(net528));
 sg13g2_antennanp ANTENNA_1844 (.A(net528));
 sg13g2_antennanp ANTENNA_1845 (.A(net528));
 sg13g2_antennanp ANTENNA_1846 (.A(net528));
 sg13g2_antennanp ANTENNA_1847 (.A(net528));
 sg13g2_antennanp ANTENNA_1848 (.A(net528));
 sg13g2_antennanp ANTENNA_1849 (.A(net528));
 sg13g2_antennanp ANTENNA_1850 (.A(net528));
 sg13g2_antennanp ANTENNA_1851 (.A(net529));
 sg13g2_antennanp ANTENNA_1852 (.A(net529));
 sg13g2_antennanp ANTENNA_1853 (.A(net529));
 sg13g2_antennanp ANTENNA_1854 (.A(net529));
 sg13g2_antennanp ANTENNA_1855 (.A(net529));
 sg13g2_antennanp ANTENNA_1856 (.A(net529));
 sg13g2_antennanp ANTENNA_1857 (.A(net529));
 sg13g2_antennanp ANTENNA_1858 (.A(net529));
 sg13g2_antennanp ANTENNA_1859 (.A(net529));
 sg13g2_antennanp ANTENNA_1860 (.A(net529));
 sg13g2_antennanp ANTENNA_1861 (.A(net529));
 sg13g2_antennanp ANTENNA_1862 (.A(net529));
 sg13g2_antennanp ANTENNA_1863 (.A(net529));
 sg13g2_antennanp ANTENNA_1864 (.A(net529));
 sg13g2_antennanp ANTENNA_1865 (.A(net529));
 sg13g2_antennanp ANTENNA_1866 (.A(net549));
 sg13g2_antennanp ANTENNA_1867 (.A(net549));
 sg13g2_antennanp ANTENNA_1868 (.A(net549));
 sg13g2_antennanp ANTENNA_1869 (.A(net549));
 sg13g2_antennanp ANTENNA_1870 (.A(net549));
 sg13g2_antennanp ANTENNA_1871 (.A(net549));
 sg13g2_antennanp ANTENNA_1872 (.A(net549));
 sg13g2_antennanp ANTENNA_1873 (.A(net549));
 sg13g2_antennanp ANTENNA_1874 (.A(net549));
 sg13g2_antennanp ANTENNA_1875 (.A(net549));
 sg13g2_antennanp ANTENNA_1876 (.A(net549));
 sg13g2_antennanp ANTENNA_1877 (.A(net549));
 sg13g2_antennanp ANTENNA_1878 (.A(net549));
 sg13g2_antennanp ANTENNA_1879 (.A(net549));
 sg13g2_antennanp ANTENNA_1880 (.A(net549));
 sg13g2_antennanp ANTENNA_1881 (.A(net549));
 sg13g2_antennanp ANTENNA_1882 (.A(net549));
 sg13g2_antennanp ANTENNA_1883 (.A(net549));
 sg13g2_antennanp ANTENNA_1884 (.A(net549));
 sg13g2_antennanp ANTENNA_1885 (.A(net549));
 sg13g2_antennanp ANTENNA_1886 (.A(net549));
 sg13g2_antennanp ANTENNA_1887 (.A(net549));
 sg13g2_antennanp ANTENNA_1888 (.A(net549));
 sg13g2_antennanp ANTENNA_1889 (.A(net551));
 sg13g2_antennanp ANTENNA_1890 (.A(net551));
 sg13g2_antennanp ANTENNA_1891 (.A(net551));
 sg13g2_antennanp ANTENNA_1892 (.A(net551));
 sg13g2_antennanp ANTENNA_1893 (.A(net551));
 sg13g2_antennanp ANTENNA_1894 (.A(net551));
 sg13g2_antennanp ANTENNA_1895 (.A(net551));
 sg13g2_antennanp ANTENNA_1896 (.A(net551));
 sg13g2_antennanp ANTENNA_1897 (.A(net551));
 sg13g2_antennanp ANTENNA_1898 (.A(net553));
 sg13g2_antennanp ANTENNA_1899 (.A(net553));
 sg13g2_antennanp ANTENNA_1900 (.A(net553));
 sg13g2_antennanp ANTENNA_1901 (.A(net553));
 sg13g2_antennanp ANTENNA_1902 (.A(net553));
 sg13g2_antennanp ANTENNA_1903 (.A(net553));
 sg13g2_antennanp ANTENNA_1904 (.A(net553));
 sg13g2_antennanp ANTENNA_1905 (.A(net553));
 sg13g2_antennanp ANTENNA_1906 (.A(net554));
 sg13g2_antennanp ANTENNA_1907 (.A(net554));
 sg13g2_antennanp ANTENNA_1908 (.A(net554));
 sg13g2_antennanp ANTENNA_1909 (.A(net554));
 sg13g2_antennanp ANTENNA_1910 (.A(net554));
 sg13g2_antennanp ANTENNA_1911 (.A(net554));
 sg13g2_antennanp ANTENNA_1912 (.A(net554));
 sg13g2_antennanp ANTENNA_1913 (.A(net554));
 sg13g2_antennanp ANTENNA_1914 (.A(net554));
 sg13g2_antennanp ANTENNA_1915 (.A(net554));
 sg13g2_antennanp ANTENNA_1916 (.A(net554));
 sg13g2_antennanp ANTENNA_1917 (.A(net554));
 sg13g2_antennanp ANTENNA_1918 (.A(net554));
 sg13g2_antennanp ANTENNA_1919 (.A(net554));
 sg13g2_antennanp ANTENNA_1920 (.A(net554));
 sg13g2_antennanp ANTENNA_1921 (.A(net554));
 sg13g2_antennanp ANTENNA_1922 (.A(net554));
 sg13g2_antennanp ANTENNA_1923 (.A(net554));
 sg13g2_antennanp ANTENNA_1924 (.A(net554));
 sg13g2_antennanp ANTENNA_1925 (.A(net554));
 sg13g2_antennanp ANTENNA_1926 (.A(net554));
 sg13g2_antennanp ANTENNA_1927 (.A(net554));
 sg13g2_antennanp ANTENNA_1928 (.A(net554));
 sg13g2_antennanp ANTENNA_1929 (.A(net554));
 sg13g2_antennanp ANTENNA_1930 (.A(net554));
 sg13g2_antennanp ANTENNA_1931 (.A(net641));
 sg13g2_antennanp ANTENNA_1932 (.A(net641));
 sg13g2_antennanp ANTENNA_1933 (.A(net641));
 sg13g2_antennanp ANTENNA_1934 (.A(net641));
 sg13g2_antennanp ANTENNA_1935 (.A(net641));
 sg13g2_antennanp ANTENNA_1936 (.A(net641));
 sg13g2_antennanp ANTENNA_1937 (.A(net641));
 sg13g2_antennanp ANTENNA_1938 (.A(net641));
 sg13g2_antennanp ANTENNA_1939 (.A(net641));
 sg13g2_antennanp ANTENNA_1940 (.A(net697));
 sg13g2_antennanp ANTENNA_1941 (.A(net697));
 sg13g2_antennanp ANTENNA_1942 (.A(net697));
 sg13g2_antennanp ANTENNA_1943 (.A(net697));
 sg13g2_antennanp ANTENNA_1944 (.A(net697));
 sg13g2_antennanp ANTENNA_1945 (.A(net697));
 sg13g2_antennanp ANTENNA_1946 (.A(net697));
 sg13g2_antennanp ANTENNA_1947 (.A(net697));
 sg13g2_antennanp ANTENNA_1948 (.A(net697));
 sg13g2_antennanp ANTENNA_1949 (.A(net773));
 sg13g2_antennanp ANTENNA_1950 (.A(net773));
 sg13g2_antennanp ANTENNA_1951 (.A(net773));
 sg13g2_antennanp ANTENNA_1952 (.A(net773));
 sg13g2_antennanp ANTENNA_1953 (.A(net773));
 sg13g2_antennanp ANTENNA_1954 (.A(net773));
 sg13g2_antennanp ANTENNA_1955 (.A(net773));
 sg13g2_antennanp ANTENNA_1956 (.A(net773));
 sg13g2_antennanp ANTENNA_1957 (.A(net773));
 sg13g2_antennanp ANTENNA_1958 (.A(net775));
 sg13g2_antennanp ANTENNA_1959 (.A(net775));
 sg13g2_antennanp ANTENNA_1960 (.A(net775));
 sg13g2_antennanp ANTENNA_1961 (.A(net775));
 sg13g2_antennanp ANTENNA_1962 (.A(net775));
 sg13g2_antennanp ANTENNA_1963 (.A(net775));
 sg13g2_antennanp ANTENNA_1964 (.A(net775));
 sg13g2_antennanp ANTENNA_1965 (.A(net775));
 sg13g2_antennanp ANTENNA_1966 (.A(net775));
 sg13g2_antennanp ANTENNA_1967 (.A(net775));
 sg13g2_antennanp ANTENNA_1968 (.A(net775));
 sg13g2_antennanp ANTENNA_1969 (.A(net775));
 sg13g2_antennanp ANTENNA_1970 (.A(net775));
 sg13g2_antennanp ANTENNA_1971 (.A(net775));
 sg13g2_antennanp ANTENNA_1972 (.A(net778));
 sg13g2_antennanp ANTENNA_1973 (.A(net778));
 sg13g2_antennanp ANTENNA_1974 (.A(net778));
 sg13g2_antennanp ANTENNA_1975 (.A(net778));
 sg13g2_antennanp ANTENNA_1976 (.A(net778));
 sg13g2_antennanp ANTENNA_1977 (.A(net778));
 sg13g2_antennanp ANTENNA_1978 (.A(net778));
 sg13g2_antennanp ANTENNA_1979 (.A(net778));
 sg13g2_antennanp ANTENNA_1980 (.A(net778));
 sg13g2_antennanp ANTENNA_1981 (.A(net778));
 sg13g2_antennanp ANTENNA_1982 (.A(net778));
 sg13g2_antennanp ANTENNA_1983 (.A(net778));
 sg13g2_antennanp ANTENNA_1984 (.A(net778));
 sg13g2_antennanp ANTENNA_1985 (.A(net778));
 sg13g2_antennanp ANTENNA_1986 (.A(net778));
 sg13g2_antennanp ANTENNA_1987 (.A(net778));
 sg13g2_antennanp ANTENNA_1988 (.A(net791));
 sg13g2_antennanp ANTENNA_1989 (.A(net791));
 sg13g2_antennanp ANTENNA_1990 (.A(net791));
 sg13g2_antennanp ANTENNA_1991 (.A(net791));
 sg13g2_antennanp ANTENNA_1992 (.A(net791));
 sg13g2_antennanp ANTENNA_1993 (.A(net791));
 sg13g2_antennanp ANTENNA_1994 (.A(net791));
 sg13g2_antennanp ANTENNA_1995 (.A(net791));
 sg13g2_antennanp ANTENNA_1996 (.A(net791));
 sg13g2_antennanp ANTENNA_1997 (.A(net791));
 sg13g2_antennanp ANTENNA_1998 (.A(net791));
 sg13g2_antennanp ANTENNA_1999 (.A(net791));
 sg13g2_antennanp ANTENNA_2000 (.A(net791));
 sg13g2_antennanp ANTENNA_2001 (.A(net791));
 sg13g2_antennanp ANTENNA_2002 (.A(net791));
 sg13g2_antennanp ANTENNA_2003 (.A(net791));
 sg13g2_antennanp ANTENNA_2004 (.A(net791));
 sg13g2_antennanp ANTENNA_2005 (.A(net791));
 sg13g2_antennanp ANTENNA_2006 (.A(net791));
 sg13g2_antennanp ANTENNA_2007 (.A(net791));
 sg13g2_antennanp ANTENNA_2008 (.A(net791));
 sg13g2_antennanp ANTENNA_2009 (.A(net791));
 sg13g2_antennanp ANTENNA_2010 (.A(net791));
 sg13g2_antennanp ANTENNA_2011 (.A(net791));
 sg13g2_antennanp ANTENNA_2012 (.A(net791));
 sg13g2_antennanp ANTENNA_2013 (.A(net791));
 sg13g2_antennanp ANTENNA_2014 (.A(net791));
 sg13g2_antennanp ANTENNA_2015 (.A(net791));
 sg13g2_antennanp ANTENNA_2016 (.A(net791));
 sg13g2_antennanp ANTENNA_2017 (.A(net792));
 sg13g2_antennanp ANTENNA_2018 (.A(net792));
 sg13g2_antennanp ANTENNA_2019 (.A(net792));
 sg13g2_antennanp ANTENNA_2020 (.A(net792));
 sg13g2_antennanp ANTENNA_2021 (.A(net792));
 sg13g2_antennanp ANTENNA_2022 (.A(net792));
 sg13g2_antennanp ANTENNA_2023 (.A(net792));
 sg13g2_antennanp ANTENNA_2024 (.A(net792));
 sg13g2_antennanp ANTENNA_2025 (.A(net802));
 sg13g2_antennanp ANTENNA_2026 (.A(net802));
 sg13g2_antennanp ANTENNA_2027 (.A(net802));
 sg13g2_antennanp ANTENNA_2028 (.A(net802));
 sg13g2_antennanp ANTENNA_2029 (.A(net802));
 sg13g2_antennanp ANTENNA_2030 (.A(net802));
 sg13g2_antennanp ANTENNA_2031 (.A(net802));
 sg13g2_antennanp ANTENNA_2032 (.A(net802));
 sg13g2_antennanp ANTENNA_2033 (.A(net802));
 sg13g2_antennanp ANTENNA_2034 (.A(net838));
 sg13g2_antennanp ANTENNA_2035 (.A(net838));
 sg13g2_antennanp ANTENNA_2036 (.A(net838));
 sg13g2_antennanp ANTENNA_2037 (.A(net838));
 sg13g2_antennanp ANTENNA_2038 (.A(net838));
 sg13g2_antennanp ANTENNA_2039 (.A(net838));
 sg13g2_antennanp ANTENNA_2040 (.A(net838));
 sg13g2_antennanp ANTENNA_2041 (.A(net838));
 sg13g2_antennanp ANTENNA_2042 (.A(net838));
 sg13g2_antennanp ANTENNA_2043 (.A(net839));
 sg13g2_antennanp ANTENNA_2044 (.A(net839));
 sg13g2_antennanp ANTENNA_2045 (.A(net839));
 sg13g2_antennanp ANTENNA_2046 (.A(net839));
 sg13g2_antennanp ANTENNA_2047 (.A(net839));
 sg13g2_antennanp ANTENNA_2048 (.A(net839));
 sg13g2_antennanp ANTENNA_2049 (.A(net839));
 sg13g2_antennanp ANTENNA_2050 (.A(net839));
 sg13g2_antennanp ANTENNA_2051 (.A(net839));
 sg13g2_antennanp ANTENNA_2052 (.A(net878));
 sg13g2_antennanp ANTENNA_2053 (.A(net878));
 sg13g2_antennanp ANTENNA_2054 (.A(net878));
 sg13g2_antennanp ANTENNA_2055 (.A(net878));
 sg13g2_antennanp ANTENNA_2056 (.A(net878));
 sg13g2_antennanp ANTENNA_2057 (.A(net878));
 sg13g2_antennanp ANTENNA_2058 (.A(net878));
 sg13g2_antennanp ANTENNA_2059 (.A(net878));
 sg13g2_antennanp ANTENNA_2060 (.A(net878));
 sg13g2_antennanp ANTENNA_2061 (.A(net878));
 sg13g2_antennanp ANTENNA_2062 (.A(net878));
 sg13g2_antennanp ANTENNA_2063 (.A(net878));
 sg13g2_antennanp ANTENNA_2064 (.A(net878));
 sg13g2_antennanp ANTENNA_2065 (.A(net878));
 sg13g2_antennanp ANTENNA_2066 (.A(net878));
 sg13g2_antennanp ANTENNA_2067 (.A(net878));
 sg13g2_antennanp ANTENNA_2068 (.A(net878));
 sg13g2_antennanp ANTENNA_2069 (.A(net878));
 sg13g2_antennanp ANTENNA_2070 (.A(net878));
 sg13g2_antennanp ANTENNA_2071 (.A(net878));
 sg13g2_antennanp ANTENNA_2072 (.A(net878));
 sg13g2_antennanp ANTENNA_2073 (.A(net878));
 sg13g2_antennanp ANTENNA_2074 (.A(net878));
 sg13g2_antennanp ANTENNA_2075 (.A(net878));
 sg13g2_antennanp ANTENNA_2076 (.A(net878));
 sg13g2_antennanp ANTENNA_2077 (.A(net878));
 sg13g2_antennanp ANTENNA_2078 (.A(net878));
 sg13g2_antennanp ANTENNA_2079 (.A(net878));
 sg13g2_antennanp ANTENNA_2080 (.A(net878));
 sg13g2_antennanp ANTENNA_2081 (.A(net878));
 sg13g2_antennanp ANTENNA_2082 (.A(net878));
 sg13g2_antennanp ANTENNA_2083 (.A(net878));
 sg13g2_antennanp ANTENNA_2084 (.A(net878));
 sg13g2_antennanp ANTENNA_2085 (.A(net878));
 sg13g2_antennanp ANTENNA_2086 (.A(net878));
 sg13g2_antennanp ANTENNA_2087 (.A(net878));
 sg13g2_antennanp ANTENNA_2088 (.A(net878));
 sg13g2_antennanp ANTENNA_2089 (.A(net878));
 sg13g2_antennanp ANTENNA_2090 (.A(net878));
 sg13g2_antennanp ANTENNA_2091 (.A(net878));
 sg13g2_antennanp ANTENNA_2092 (.A(net878));
 sg13g2_antennanp ANTENNA_2093 (.A(net878));
 sg13g2_antennanp ANTENNA_2094 (.A(net878));
 sg13g2_antennanp ANTENNA_2095 (.A(net878));
 sg13g2_antennanp ANTENNA_2096 (.A(net878));
 sg13g2_antennanp ANTENNA_2097 (.A(net878));
 sg13g2_antennanp ANTENNA_2098 (.A(net878));
 sg13g2_antennanp ANTENNA_2099 (.A(net878));
 sg13g2_antennanp ANTENNA_2100 (.A(net924));
 sg13g2_antennanp ANTENNA_2101 (.A(net924));
 sg13g2_antennanp ANTENNA_2102 (.A(net924));
 sg13g2_antennanp ANTENNA_2103 (.A(net924));
 sg13g2_antennanp ANTENNA_2104 (.A(net924));
 sg13g2_antennanp ANTENNA_2105 (.A(net924));
 sg13g2_antennanp ANTENNA_2106 (.A(net924));
 sg13g2_antennanp ANTENNA_2107 (.A(net924));
 sg13g2_antennanp ANTENNA_2108 (.A(net924));
 sg13g2_antennanp ANTENNA_2109 (.A(net925));
 sg13g2_antennanp ANTENNA_2110 (.A(net925));
 sg13g2_antennanp ANTENNA_2111 (.A(net925));
 sg13g2_antennanp ANTENNA_2112 (.A(net925));
 sg13g2_antennanp ANTENNA_2113 (.A(net925));
 sg13g2_antennanp ANTENNA_2114 (.A(net925));
 sg13g2_antennanp ANTENNA_2115 (.A(net925));
 sg13g2_antennanp ANTENNA_2116 (.A(net925));
 sg13g2_antennanp ANTENNA_2117 (.A(net925));
 sg13g2_antennanp ANTENNA_2118 (.A(net982));
 sg13g2_antennanp ANTENNA_2119 (.A(net982));
 sg13g2_antennanp ANTENNA_2120 (.A(net982));
 sg13g2_antennanp ANTENNA_2121 (.A(net982));
 sg13g2_antennanp ANTENNA_2122 (.A(net982));
 sg13g2_antennanp ANTENNA_2123 (.A(net982));
 sg13g2_antennanp ANTENNA_2124 (.A(net982));
 sg13g2_antennanp ANTENNA_2125 (.A(net982));
 sg13g2_antennanp ANTENNA_2126 (.A(net982));
 sg13g2_antennanp ANTENNA_2127 (.A(net989));
 sg13g2_antennanp ANTENNA_2128 (.A(net989));
 sg13g2_antennanp ANTENNA_2129 (.A(net989));
 sg13g2_antennanp ANTENNA_2130 (.A(net989));
 sg13g2_antennanp ANTENNA_2131 (.A(net989));
 sg13g2_antennanp ANTENNA_2132 (.A(net989));
 sg13g2_antennanp ANTENNA_2133 (.A(net989));
 sg13g2_antennanp ANTENNA_2134 (.A(net989));
 sg13g2_antennanp ANTENNA_2135 (.A(net989));
 sg13g2_antennanp ANTENNA_2136 (.A(net990));
 sg13g2_antennanp ANTENNA_2137 (.A(net990));
 sg13g2_antennanp ANTENNA_2138 (.A(net990));
 sg13g2_antennanp ANTENNA_2139 (.A(net990));
 sg13g2_antennanp ANTENNA_2140 (.A(net990));
 sg13g2_antennanp ANTENNA_2141 (.A(net990));
 sg13g2_antennanp ANTENNA_2142 (.A(net990));
 sg13g2_antennanp ANTENNA_2143 (.A(net990));
 sg13g2_antennanp ANTENNA_2144 (.A(net990));
 sg13g2_antennanp ANTENNA_2145 (.A(net990));
 sg13g2_antennanp ANTENNA_2146 (.A(net990));
 sg13g2_antennanp ANTENNA_2147 (.A(net990));
 sg13g2_antennanp ANTENNA_2148 (.A(net990));
 sg13g2_antennanp ANTENNA_2149 (.A(net990));
 sg13g2_antennanp ANTENNA_2150 (.A(net990));
 sg13g2_antennanp ANTENNA_2151 (.A(net990));
 sg13g2_antennanp ANTENNA_2152 (.A(net990));
 sg13g2_antennanp ANTENNA_2153 (.A(net990));
 sg13g2_antennanp ANTENNA_2154 (.A(net990));
 sg13g2_antennanp ANTENNA_2155 (.A(net990));
 sg13g2_antennanp ANTENNA_2156 (.A(net990));
 sg13g2_antennanp ANTENNA_2157 (.A(net1051));
 sg13g2_antennanp ANTENNA_2158 (.A(net1051));
 sg13g2_antennanp ANTENNA_2159 (.A(net1051));
 sg13g2_antennanp ANTENNA_2160 (.A(net1051));
 sg13g2_antennanp ANTENNA_2161 (.A(net1051));
 sg13g2_antennanp ANTENNA_2162 (.A(net1051));
 sg13g2_antennanp ANTENNA_2163 (.A(net1051));
 sg13g2_antennanp ANTENNA_2164 (.A(net1051));
 sg13g2_antennanp ANTENNA_2165 (.A(net1051));
 sg13g2_antennanp ANTENNA_2166 (.A(net1099));
 sg13g2_antennanp ANTENNA_2167 (.A(net1099));
 sg13g2_antennanp ANTENNA_2168 (.A(net1099));
 sg13g2_antennanp ANTENNA_2169 (.A(net1099));
 sg13g2_antennanp ANTENNA_2170 (.A(net1099));
 sg13g2_antennanp ANTENNA_2171 (.A(net1099));
 sg13g2_antennanp ANTENNA_2172 (.A(net1099));
 sg13g2_antennanp ANTENNA_2173 (.A(net1099));
 sg13g2_antennanp ANTENNA_2174 (.A(net1100));
 sg13g2_antennanp ANTENNA_2175 (.A(net1100));
 sg13g2_antennanp ANTENNA_2176 (.A(net1100));
 sg13g2_antennanp ANTENNA_2177 (.A(net1100));
 sg13g2_antennanp ANTENNA_2178 (.A(net1100));
 sg13g2_antennanp ANTENNA_2179 (.A(net1100));
 sg13g2_antennanp ANTENNA_2180 (.A(net1100));
 sg13g2_antennanp ANTENNA_2181 (.A(net1100));
 sg13g2_antennanp ANTENNA_2182 (.A(net1100));
 sg13g2_antennanp ANTENNA_2183 (.A(net1192));
 sg13g2_antennanp ANTENNA_2184 (.A(net1192));
 sg13g2_antennanp ANTENNA_2185 (.A(net1192));
 sg13g2_antennanp ANTENNA_2186 (.A(net1192));
 sg13g2_antennanp ANTENNA_2187 (.A(net1192));
 sg13g2_antennanp ANTENNA_2188 (.A(net1192));
 sg13g2_antennanp ANTENNA_2189 (.A(net1192));
 sg13g2_antennanp ANTENNA_2190 (.A(net1192));
 sg13g2_antennanp ANTENNA_2191 (.A(net1192));
 sg13g2_antennanp ANTENNA_2192 (.A(net1192));
 sg13g2_antennanp ANTENNA_2193 (.A(net1192));
 sg13g2_antennanp ANTENNA_2194 (.A(net1192));
 sg13g2_antennanp ANTENNA_2195 (.A(net1192));
 sg13g2_antennanp ANTENNA_2196 (.A(net1192));
 sg13g2_antennanp ANTENNA_2197 (.A(net1192));
 sg13g2_antennanp ANTENNA_2198 (.A(net1192));
 sg13g2_antennanp ANTENNA_2199 (.A(net1192));
 sg13g2_antennanp ANTENNA_2200 (.A(net1192));
 sg13g2_antennanp ANTENNA_2201 (.A(net1192));
 sg13g2_antennanp ANTENNA_2202 (.A(net1192));
 sg13g2_antennanp ANTENNA_2203 (.A(net1193));
 sg13g2_antennanp ANTENNA_2204 (.A(net1193));
 sg13g2_antennanp ANTENNA_2205 (.A(net1193));
 sg13g2_antennanp ANTENNA_2206 (.A(net1193));
 sg13g2_antennanp ANTENNA_2207 (.A(net1193));
 sg13g2_antennanp ANTENNA_2208 (.A(net1193));
 sg13g2_antennanp ANTENNA_2209 (.A(net1193));
 sg13g2_antennanp ANTENNA_2210 (.A(net1193));
 sg13g2_antennanp ANTENNA_2211 (.A(net1193));
 sg13g2_antennanp ANTENNA_2212 (.A(net1273));
 sg13g2_antennanp ANTENNA_2213 (.A(net1273));
 sg13g2_antennanp ANTENNA_2214 (.A(net1273));
 sg13g2_antennanp ANTENNA_2215 (.A(net1273));
 sg13g2_antennanp ANTENNA_2216 (.A(net1273));
 sg13g2_antennanp ANTENNA_2217 (.A(net1273));
 sg13g2_antennanp ANTENNA_2218 (.A(net1273));
 sg13g2_antennanp ANTENNA_2219 (.A(net1273));
 sg13g2_antennanp ANTENNA_2220 (.A(net1273));
 sg13g2_antennanp ANTENNA_2221 (.A(net1273));
 sg13g2_antennanp ANTENNA_2222 (.A(net1273));
 sg13g2_antennanp ANTENNA_2223 (.A(net1273));
 sg13g2_antennanp ANTENNA_2224 (.A(net1273));
 sg13g2_antennanp ANTENNA_2225 (.A(net1273));
 sg13g2_antennanp ANTENNA_2226 (.A(net1273));
 sg13g2_antennanp ANTENNA_2227 (.A(net1273));
 sg13g2_antennanp ANTENNA_2228 (.A(net1273));
 sg13g2_antennanp ANTENNA_2229 (.A(net1273));
 sg13g2_antennanp ANTENNA_2230 (.A(net1276));
 sg13g2_antennanp ANTENNA_2231 (.A(net1276));
 sg13g2_antennanp ANTENNA_2232 (.A(net1276));
 sg13g2_antennanp ANTENNA_2233 (.A(net1276));
 sg13g2_antennanp ANTENNA_2234 (.A(net1276));
 sg13g2_antennanp ANTENNA_2235 (.A(net1276));
 sg13g2_antennanp ANTENNA_2236 (.A(net1276));
 sg13g2_antennanp ANTENNA_2237 (.A(net1276));
 sg13g2_antennanp ANTENNA_2238 (.A(net1276));
 sg13g2_antennanp ANTENNA_2239 (.A(net1276));
 sg13g2_antennanp ANTENNA_2240 (.A(net1276));
 sg13g2_antennanp ANTENNA_2241 (.A(net1276));
 sg13g2_antennanp ANTENNA_2242 (.A(_00017_));
 sg13g2_antennanp ANTENNA_2243 (.A(_00017_));
 sg13g2_antennanp ANTENNA_2244 (.A(_00017_));
 sg13g2_antennanp ANTENNA_2245 (.A(_00017_));
 sg13g2_antennanp ANTENNA_2246 (.A(_02490_));
 sg13g2_antennanp ANTENNA_2247 (.A(_02963_));
 sg13g2_antennanp ANTENNA_2248 (.A(_03341_));
 sg13g2_antennanp ANTENNA_2249 (.A(_03341_));
 sg13g2_antennanp ANTENNA_2250 (.A(_03444_));
 sg13g2_antennanp ANTENNA_2251 (.A(_03444_));
 sg13g2_antennanp ANTENNA_2252 (.A(_03444_));
 sg13g2_antennanp ANTENNA_2253 (.A(_03444_));
 sg13g2_antennanp ANTENNA_2254 (.A(_03621_));
 sg13g2_antennanp ANTENNA_2255 (.A(_03621_));
 sg13g2_antennanp ANTENNA_2256 (.A(_03621_));
 sg13g2_antennanp ANTENNA_2257 (.A(_03621_));
 sg13g2_antennanp ANTENNA_2258 (.A(_03621_));
 sg13g2_antennanp ANTENNA_2259 (.A(_03621_));
 sg13g2_antennanp ANTENNA_2260 (.A(_03621_));
 sg13g2_antennanp ANTENNA_2261 (.A(_03621_));
 sg13g2_antennanp ANTENNA_2262 (.A(_03843_));
 sg13g2_antennanp ANTENNA_2263 (.A(_03843_));
 sg13g2_antennanp ANTENNA_2264 (.A(_03843_));
 sg13g2_antennanp ANTENNA_2265 (.A(_03843_));
 sg13g2_antennanp ANTENNA_2266 (.A(_03875_));
 sg13g2_antennanp ANTENNA_2267 (.A(_03995_));
 sg13g2_antennanp ANTENNA_2268 (.A(_03995_));
 sg13g2_antennanp ANTENNA_2269 (.A(_03995_));
 sg13g2_antennanp ANTENNA_2270 (.A(_03995_));
 sg13g2_antennanp ANTENNA_2271 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2272 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2273 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2274 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2275 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2276 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2277 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2278 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2279 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2280 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2281 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2282 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2283 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2284 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2285 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2286 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2287 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2288 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2289 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2290 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2291 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2292 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2293 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2294 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2295 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2296 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2297 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2298 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2299 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2300 (.A(_04431_));
 sg13g2_antennanp ANTENNA_2301 (.A(_05432_));
 sg13g2_antennanp ANTENNA_2302 (.A(_05432_));
 sg13g2_antennanp ANTENNA_2303 (.A(_05432_));
 sg13g2_antennanp ANTENNA_2304 (.A(_05441_));
 sg13g2_antennanp ANTENNA_2305 (.A(_05441_));
 sg13g2_antennanp ANTENNA_2306 (.A(_05441_));
 sg13g2_antennanp ANTENNA_2307 (.A(_05449_));
 sg13g2_antennanp ANTENNA_2308 (.A(_05449_));
 sg13g2_antennanp ANTENNA_2309 (.A(_05449_));
 sg13g2_antennanp ANTENNA_2310 (.A(_05449_));
 sg13g2_antennanp ANTENNA_2311 (.A(_05449_));
 sg13g2_antennanp ANTENNA_2312 (.A(_05449_));
 sg13g2_antennanp ANTENNA_2313 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2314 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2315 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2316 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2317 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2318 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2319 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2320 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2321 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2322 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2323 (.A(_05457_));
 sg13g2_antennanp ANTENNA_2324 (.A(_05457_));
 sg13g2_antennanp ANTENNA_2325 (.A(_05457_));
 sg13g2_antennanp ANTENNA_2326 (.A(_05457_));
 sg13g2_antennanp ANTENNA_2327 (.A(_05457_));
 sg13g2_antennanp ANTENNA_2328 (.A(_05457_));
 sg13g2_antennanp ANTENNA_2329 (.A(_05463_));
 sg13g2_antennanp ANTENNA_2330 (.A(_05463_));
 sg13g2_antennanp ANTENNA_2331 (.A(_05463_));
 sg13g2_antennanp ANTENNA_2332 (.A(_05463_));
 sg13g2_antennanp ANTENNA_2333 (.A(_05463_));
 sg13g2_antennanp ANTENNA_2334 (.A(_05463_));
 sg13g2_antennanp ANTENNA_2335 (.A(_05467_));
 sg13g2_antennanp ANTENNA_2336 (.A(_05467_));
 sg13g2_antennanp ANTENNA_2337 (.A(_05467_));
 sg13g2_antennanp ANTENNA_2338 (.A(_05467_));
 sg13g2_antennanp ANTENNA_2339 (.A(_05467_));
 sg13g2_antennanp ANTENNA_2340 (.A(_05467_));
 sg13g2_antennanp ANTENNA_2341 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2342 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2343 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2344 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2345 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2346 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2347 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2348 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2349 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2350 (.A(_05471_));
 sg13g2_antennanp ANTENNA_2351 (.A(_05476_));
 sg13g2_antennanp ANTENNA_2352 (.A(_05476_));
 sg13g2_antennanp ANTENNA_2353 (.A(_05498_));
 sg13g2_antennanp ANTENNA_2354 (.A(_05498_));
 sg13g2_antennanp ANTENNA_2355 (.A(_05542_));
 sg13g2_antennanp ANTENNA_2356 (.A(_06148_));
 sg13g2_antennanp ANTENNA_2357 (.A(_06148_));
 sg13g2_antennanp ANTENNA_2358 (.A(_06148_));
 sg13g2_antennanp ANTENNA_2359 (.A(_06148_));
 sg13g2_antennanp ANTENNA_2360 (.A(_06148_));
 sg13g2_antennanp ANTENNA_2361 (.A(_06171_));
 sg13g2_antennanp ANTENNA_2362 (.A(_06189_));
 sg13g2_antennanp ANTENNA_2363 (.A(_06253_));
 sg13g2_antennanp ANTENNA_2364 (.A(_06253_));
 sg13g2_antennanp ANTENNA_2365 (.A(_06255_));
 sg13g2_antennanp ANTENNA_2366 (.A(_06268_));
 sg13g2_antennanp ANTENNA_2367 (.A(_06293_));
 sg13g2_antennanp ANTENNA_2368 (.A(_06298_));
 sg13g2_antennanp ANTENNA_2369 (.A(_06311_));
 sg13g2_antennanp ANTENNA_2370 (.A(_06318_));
 sg13g2_antennanp ANTENNA_2371 (.A(_06329_));
 sg13g2_antennanp ANTENNA_2372 (.A(_06393_));
 sg13g2_antennanp ANTENNA_2373 (.A(_06393_));
 sg13g2_antennanp ANTENNA_2374 (.A(_06393_));
 sg13g2_antennanp ANTENNA_2375 (.A(_06393_));
 sg13g2_antennanp ANTENNA_2376 (.A(_06416_));
 sg13g2_antennanp ANTENNA_2377 (.A(_06460_));
 sg13g2_antennanp ANTENNA_2378 (.A(_06460_));
 sg13g2_antennanp ANTENNA_2379 (.A(_06493_));
 sg13g2_antennanp ANTENNA_2380 (.A(_06493_));
 sg13g2_antennanp ANTENNA_2381 (.A(_06516_));
 sg13g2_antennanp ANTENNA_2382 (.A(_06520_));
 sg13g2_antennanp ANTENNA_2383 (.A(_06559_));
 sg13g2_antennanp ANTENNA_2384 (.A(_06560_));
 sg13g2_antennanp ANTENNA_2385 (.A(_06595_));
 sg13g2_antennanp ANTENNA_2386 (.A(_06601_));
 sg13g2_antennanp ANTENNA_2387 (.A(_06601_));
 sg13g2_antennanp ANTENNA_2388 (.A(_06616_));
 sg13g2_antennanp ANTENNA_2389 (.A(_06620_));
 sg13g2_antennanp ANTENNA_2390 (.A(_06620_));
 sg13g2_antennanp ANTENNA_2391 (.A(_06658_));
 sg13g2_antennanp ANTENNA_2392 (.A(_06694_));
 sg13g2_antennanp ANTENNA_2393 (.A(_06700_));
 sg13g2_antennanp ANTENNA_2394 (.A(_06717_));
 sg13g2_antennanp ANTENNA_2395 (.A(_06719_));
 sg13g2_antennanp ANTENNA_2396 (.A(_06719_));
 sg13g2_antennanp ANTENNA_2397 (.A(_06757_));
 sg13g2_antennanp ANTENNA_2398 (.A(_06772_));
 sg13g2_antennanp ANTENNA_2399 (.A(_06772_));
 sg13g2_antennanp ANTENNA_2400 (.A(_06793_));
 sg13g2_antennanp ANTENNA_2401 (.A(_06793_));
 sg13g2_antennanp ANTENNA_2402 (.A(_06799_));
 sg13g2_antennanp ANTENNA_2403 (.A(_06799_));
 sg13g2_antennanp ANTENNA_2404 (.A(_06814_));
 sg13g2_antennanp ANTENNA_2405 (.A(_06814_));
 sg13g2_antennanp ANTENNA_2406 (.A(_06818_));
 sg13g2_antennanp ANTENNA_2407 (.A(_06856_));
 sg13g2_antennanp ANTENNA_2408 (.A(_06871_));
 sg13g2_antennanp ANTENNA_2409 (.A(_06871_));
 sg13g2_antennanp ANTENNA_2410 (.A(_06913_));
 sg13g2_antennanp ANTENNA_2411 (.A(_06917_));
 sg13g2_antennanp ANTENNA_2412 (.A(_06955_));
 sg13g2_antennanp ANTENNA_2413 (.A(_06955_));
 sg13g2_antennanp ANTENNA_2414 (.A(_06975_));
 sg13g2_antennanp ANTENNA_2415 (.A(_06991_));
 sg13g2_antennanp ANTENNA_2416 (.A(_07012_));
 sg13g2_antennanp ANTENNA_2417 (.A(_07012_));
 sg13g2_antennanp ANTENNA_2418 (.A(_07016_));
 sg13g2_antennanp ANTENNA_2419 (.A(_07054_));
 sg13g2_antennanp ANTENNA_2420 (.A(_07054_));
 sg13g2_antennanp ANTENNA_2421 (.A(_07074_));
 sg13g2_antennanp ANTENNA_2422 (.A(_07074_));
 sg13g2_antennanp ANTENNA_2423 (.A(_07090_));
 sg13g2_antennanp ANTENNA_2424 (.A(_07105_));
 sg13g2_antennanp ANTENNA_2425 (.A(_07105_));
 sg13g2_antennanp ANTENNA_2426 (.A(_07335_));
 sg13g2_antennanp ANTENNA_2427 (.A(_09194_));
 sg13g2_antennanp ANTENNA_2428 (.A(_09194_));
 sg13g2_antennanp ANTENNA_2429 (.A(_09194_));
 sg13g2_antennanp ANTENNA_2430 (.A(_09194_));
 sg13g2_antennanp ANTENNA_2431 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2432 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2433 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2434 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2435 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2436 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2437 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2438 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2439 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2440 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2441 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2442 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2443 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2444 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2445 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2446 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2447 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2448 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2449 (.A(_09418_));
 sg13g2_antennanp ANTENNA_2450 (.A(_09418_));
 sg13g2_antennanp ANTENNA_2451 (.A(_09418_));
 sg13g2_antennanp ANTENNA_2452 (.A(_09418_));
 sg13g2_antennanp ANTENNA_2453 (.A(_09418_));
 sg13g2_antennanp ANTENNA_2454 (.A(_09418_));
 sg13g2_antennanp ANTENNA_2455 (.A(_09418_));
 sg13g2_antennanp ANTENNA_2456 (.A(_09418_));
 sg13g2_antennanp ANTENNA_2457 (.A(_09418_));
 sg13g2_antennanp ANTENNA_2458 (.A(_09906_));
 sg13g2_antennanp ANTENNA_2459 (.A(_09906_));
 sg13g2_antennanp ANTENNA_2460 (.A(_09906_));
 sg13g2_antennanp ANTENNA_2461 (.A(_09906_));
 sg13g2_antennanp ANTENNA_2462 (.A(_09906_));
 sg13g2_antennanp ANTENNA_2463 (.A(_09906_));
 sg13g2_antennanp ANTENNA_2464 (.A(_09906_));
 sg13g2_antennanp ANTENNA_2465 (.A(_09906_));
 sg13g2_antennanp ANTENNA_2466 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2467 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2468 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2469 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2470 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2471 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2472 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2473 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2474 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2475 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2476 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2477 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2478 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2479 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2480 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2481 (.A(_09928_));
 sg13g2_antennanp ANTENNA_2482 (.A(_09929_));
 sg13g2_antennanp ANTENNA_2483 (.A(_09929_));
 sg13g2_antennanp ANTENNA_2484 (.A(_09929_));
 sg13g2_antennanp ANTENNA_2485 (.A(_09929_));
 sg13g2_antennanp ANTENNA_2486 (.A(_10040_));
 sg13g2_antennanp ANTENNA_2487 (.A(_10040_));
 sg13g2_antennanp ANTENNA_2488 (.A(_10040_));
 sg13g2_antennanp ANTENNA_2489 (.A(_10042_));
 sg13g2_antennanp ANTENNA_2490 (.A(_10042_));
 sg13g2_antennanp ANTENNA_2491 (.A(_10042_));
 sg13g2_antennanp ANTENNA_2492 (.A(_10042_));
 sg13g2_antennanp ANTENNA_2493 (.A(_10046_));
 sg13g2_antennanp ANTENNA_2494 (.A(_10048_));
 sg13g2_antennanp ANTENNA_2495 (.A(_10051_));
 sg13g2_antennanp ANTENNA_2496 (.A(_10053_));
 sg13g2_antennanp ANTENNA_2497 (.A(_10083_));
 sg13g2_antennanp ANTENNA_2498 (.A(_10083_));
 sg13g2_antennanp ANTENNA_2499 (.A(_10091_));
 sg13g2_antennanp ANTENNA_2500 (.A(_10091_));
 sg13g2_antennanp ANTENNA_2501 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2502 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2503 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2504 (.A(_10101_));
 sg13g2_antennanp ANTENNA_2505 (.A(_10106_));
 sg13g2_antennanp ANTENNA_2506 (.A(_10110_));
 sg13g2_antennanp ANTENNA_2507 (.A(_10121_));
 sg13g2_antennanp ANTENNA_2508 (.A(_10131_));
 sg13g2_antennanp ANTENNA_2509 (.A(_10136_));
 sg13g2_antennanp ANTENNA_2510 (.A(_10140_));
 sg13g2_antennanp ANTENNA_2511 (.A(_10226_));
 sg13g2_antennanp ANTENNA_2512 (.A(_10226_));
 sg13g2_antennanp ANTENNA_2513 (.A(_10226_));
 sg13g2_antennanp ANTENNA_2514 (.A(_10235_));
 sg13g2_antennanp ANTENNA_2515 (.A(_10235_));
 sg13g2_antennanp ANTENNA_2516 (.A(_10235_));
 sg13g2_antennanp ANTENNA_2517 (.A(_10235_));
 sg13g2_antennanp ANTENNA_2518 (.A(_10236_));
 sg13g2_antennanp ANTENNA_2519 (.A(_10236_));
 sg13g2_antennanp ANTENNA_2520 (.A(_10236_));
 sg13g2_antennanp ANTENNA_2521 (.A(_10236_));
 sg13g2_antennanp ANTENNA_2522 (.A(_10236_));
 sg13g2_antennanp ANTENNA_2523 (.A(_10236_));
 sg13g2_antennanp ANTENNA_2524 (.A(_10236_));
 sg13g2_antennanp ANTENNA_2525 (.A(_10243_));
 sg13g2_antennanp ANTENNA_2526 (.A(_10243_));
 sg13g2_antennanp ANTENNA_2527 (.A(_10243_));
 sg13g2_antennanp ANTENNA_2528 (.A(_10243_));
 sg13g2_antennanp ANTENNA_2529 (.A(_10243_));
 sg13g2_antennanp ANTENNA_2530 (.A(_10243_));
 sg13g2_antennanp ANTENNA_2531 (.A(_10256_));
 sg13g2_antennanp ANTENNA_2532 (.A(_10256_));
 sg13g2_antennanp ANTENNA_2533 (.A(_10256_));
 sg13g2_antennanp ANTENNA_2534 (.A(_10256_));
 sg13g2_antennanp ANTENNA_2535 (.A(_10256_));
 sg13g2_antennanp ANTENNA_2536 (.A(_10287_));
 sg13g2_antennanp ANTENNA_2537 (.A(_10287_));
 sg13g2_antennanp ANTENNA_2538 (.A(_10287_));
 sg13g2_antennanp ANTENNA_2539 (.A(_10287_));
 sg13g2_antennanp ANTENNA_2540 (.A(_10295_));
 sg13g2_antennanp ANTENNA_2541 (.A(_10295_));
 sg13g2_antennanp ANTENNA_2542 (.A(_10295_));
 sg13g2_antennanp ANTENNA_2543 (.A(_10295_));
 sg13g2_antennanp ANTENNA_2544 (.A(_10295_));
 sg13g2_antennanp ANTENNA_2545 (.A(_10295_));
 sg13g2_antennanp ANTENNA_2546 (.A(_10295_));
 sg13g2_antennanp ANTENNA_2547 (.A(_10295_));
 sg13g2_antennanp ANTENNA_2548 (.A(_10296_));
 sg13g2_antennanp ANTENNA_2549 (.A(_10296_));
 sg13g2_antennanp ANTENNA_2550 (.A(_10296_));
 sg13g2_antennanp ANTENNA_2551 (.A(_10296_));
 sg13g2_antennanp ANTENNA_2552 (.A(_10296_));
 sg13g2_antennanp ANTENNA_2553 (.A(_10325_));
 sg13g2_antennanp ANTENNA_2554 (.A(_10325_));
 sg13g2_antennanp ANTENNA_2555 (.A(_10325_));
 sg13g2_antennanp ANTENNA_2556 (.A(_10325_));
 sg13g2_antennanp ANTENNA_2557 (.A(_10325_));
 sg13g2_antennanp ANTENNA_2558 (.A(_10325_));
 sg13g2_antennanp ANTENNA_2559 (.A(_10325_));
 sg13g2_antennanp ANTENNA_2560 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2561 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2562 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2563 (.A(_10349_));
 sg13g2_antennanp ANTENNA_2564 (.A(_10349_));
 sg13g2_antennanp ANTENNA_2565 (.A(_10349_));
 sg13g2_antennanp ANTENNA_2566 (.A(_10349_));
 sg13g2_antennanp ANTENNA_2567 (.A(_10397_));
 sg13g2_antennanp ANTENNA_2568 (.A(_10397_));
 sg13g2_antennanp ANTENNA_2569 (.A(_10397_));
 sg13g2_antennanp ANTENNA_2570 (.A(_10397_));
 sg13g2_antennanp ANTENNA_2571 (.A(_10397_));
 sg13g2_antennanp ANTENNA_2572 (.A(_10397_));
 sg13g2_antennanp ANTENNA_2573 (.A(_10397_));
 sg13g2_antennanp ANTENNA_2574 (.A(_10397_));
 sg13g2_antennanp ANTENNA_2575 (.A(_10415_));
 sg13g2_antennanp ANTENNA_2576 (.A(_10415_));
 sg13g2_antennanp ANTENNA_2577 (.A(_10415_));
 sg13g2_antennanp ANTENNA_2578 (.A(_10415_));
 sg13g2_antennanp ANTENNA_2579 (.A(_10415_));
 sg13g2_antennanp ANTENNA_2580 (.A(_10415_));
 sg13g2_antennanp ANTENNA_2581 (.A(_10415_));
 sg13g2_antennanp ANTENNA_2582 (.A(_10415_));
 sg13g2_antennanp ANTENNA_2583 (.A(_10415_));
 sg13g2_antennanp ANTENNA_2584 (.A(_10422_));
 sg13g2_antennanp ANTENNA_2585 (.A(_10422_));
 sg13g2_antennanp ANTENNA_2586 (.A(_10422_));
 sg13g2_antennanp ANTENNA_2587 (.A(_10422_));
 sg13g2_antennanp ANTENNA_2588 (.A(_10422_));
 sg13g2_antennanp ANTENNA_2589 (.A(_10422_));
 sg13g2_antennanp ANTENNA_2590 (.A(_10422_));
 sg13g2_antennanp ANTENNA_2591 (.A(_10422_));
 sg13g2_antennanp ANTENNA_2592 (.A(_10422_));
 sg13g2_antennanp ANTENNA_2593 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2594 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2595 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2596 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2597 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2598 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2599 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2600 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2601 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2602 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2603 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2604 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2605 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2606 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2607 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2608 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2609 (.A(_10444_));
 sg13g2_antennanp ANTENNA_2610 (.A(_10468_));
 sg13g2_antennanp ANTENNA_2611 (.A(_10468_));
 sg13g2_antennanp ANTENNA_2612 (.A(_10468_));
 sg13g2_antennanp ANTENNA_2613 (.A(_10468_));
 sg13g2_antennanp ANTENNA_2614 (.A(_10468_));
 sg13g2_antennanp ANTENNA_2615 (.A(_10468_));
 sg13g2_antennanp ANTENNA_2616 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2617 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2618 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2619 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2620 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2621 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2622 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2623 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2624 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2625 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2626 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2627 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2628 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2629 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2630 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2631 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2632 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2633 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2634 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2635 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2636 (.A(_10513_));
 sg13g2_antennanp ANTENNA_2637 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2638 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2639 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2640 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2641 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2642 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2643 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2644 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2645 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2646 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2647 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2648 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2649 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2650 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2651 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2652 (.A(_10564_));
 sg13g2_antennanp ANTENNA_2653 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2654 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2655 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2656 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2657 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2658 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2659 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2660 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2661 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2662 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2663 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2664 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2665 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2666 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2667 (.A(_10586_));
 sg13g2_antennanp ANTENNA_2668 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2669 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2670 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2671 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2672 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2673 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2674 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2675 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2676 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2677 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2678 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2679 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2680 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2681 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2682 (.A(_10632_));
 sg13g2_antennanp ANTENNA_2683 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2684 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2685 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2686 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2687 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2688 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2689 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2690 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2691 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2692 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2693 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2694 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2695 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2696 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2697 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2698 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2699 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2700 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2701 (.A(_10656_));
 sg13g2_antennanp ANTENNA_2702 (.A(_10679_));
 sg13g2_antennanp ANTENNA_2703 (.A(_10679_));
 sg13g2_antennanp ANTENNA_2704 (.A(_10679_));
 sg13g2_antennanp ANTENNA_2705 (.A(_10679_));
 sg13g2_antennanp ANTENNA_2706 (.A(_10679_));
 sg13g2_antennanp ANTENNA_2707 (.A(_10679_));
 sg13g2_antennanp ANTENNA_2708 (.A(_10679_));
 sg13g2_antennanp ANTENNA_2709 (.A(_10679_));
 sg13g2_antennanp ANTENNA_2710 (.A(_11171_));
 sg13g2_antennanp ANTENNA_2711 (.A(_11171_));
 sg13g2_antennanp ANTENNA_2712 (.A(_11171_));
 sg13g2_antennanp ANTENNA_2713 (.A(_11171_));
 sg13g2_antennanp ANTENNA_2714 (.A(_11171_));
 sg13g2_antennanp ANTENNA_2715 (.A(_11171_));
 sg13g2_antennanp ANTENNA_2716 (.A(_11171_));
 sg13g2_antennanp ANTENNA_2717 (.A(_11875_));
 sg13g2_antennanp ANTENNA_2718 (.A(_11875_));
 sg13g2_antennanp ANTENNA_2719 (.A(_11875_));
 sg13g2_antennanp ANTENNA_2720 (.A(_11875_));
 sg13g2_antennanp ANTENNA_2721 (.A(_11875_));
 sg13g2_antennanp ANTENNA_2722 (.A(_11875_));
 sg13g2_antennanp ANTENNA_2723 (.A(_11875_));
 sg13g2_antennanp ANTENNA_2724 (.A(_11947_));
 sg13g2_antennanp ANTENNA_2725 (.A(_11947_));
 sg13g2_antennanp ANTENNA_2726 (.A(_11947_));
 sg13g2_antennanp ANTENNA_2727 (.A(_11947_));
 sg13g2_antennanp ANTENNA_2728 (.A(_12437_));
 sg13g2_antennanp ANTENNA_2729 (.A(_12437_));
 sg13g2_antennanp ANTENNA_2730 (.A(_12437_));
 sg13g2_antennanp ANTENNA_2731 (.A(_12437_));
 sg13g2_antennanp ANTENNA_2732 (.A(_12437_));
 sg13g2_antennanp ANTENNA_2733 (.A(_12437_));
 sg13g2_antennanp ANTENNA_2734 (.A(_12437_));
 sg13g2_antennanp ANTENNA_2735 (.A(_12437_));
 sg13g2_antennanp ANTENNA_2736 (.A(_12443_));
 sg13g2_antennanp ANTENNA_2737 (.A(_12443_));
 sg13g2_antennanp ANTENNA_2738 (.A(_12443_));
 sg13g2_antennanp ANTENNA_2739 (.A(_12630_));
 sg13g2_antennanp ANTENNA_2740 (.A(_12630_));
 sg13g2_antennanp ANTENNA_2741 (.A(_12630_));
 sg13g2_antennanp ANTENNA_2742 (.A(_12653_));
 sg13g2_antennanp ANTENNA_2743 (.A(_12653_));
 sg13g2_antennanp ANTENNA_2744 (.A(_12653_));
 sg13g2_antennanp ANTENNA_2745 (.A(_12653_));
 sg13g2_antennanp ANTENNA_2746 (.A(_12653_));
 sg13g2_antennanp ANTENNA_2747 (.A(_12653_));
 sg13g2_antennanp ANTENNA_2748 (.A(_12653_));
 sg13g2_antennanp ANTENNA_2749 (.A(clk));
 sg13g2_antennanp ANTENNA_2750 (.A(clk));
 sg13g2_antennanp ANTENNA_2751 (.A(\mem.data_in[1] ));
 sg13g2_antennanp ANTENNA_2752 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_2753 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_2754 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_2755 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_2756 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_2757 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_2758 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_2759 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_2760 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_2761 (.A(net1));
 sg13g2_antennanp ANTENNA_2762 (.A(net1));
 sg13g2_antennanp ANTENNA_2763 (.A(net1));
 sg13g2_antennanp ANTENNA_2764 (.A(net2));
 sg13g2_antennanp ANTENNA_2765 (.A(net4));
 sg13g2_antennanp ANTENNA_2766 (.A(net464));
 sg13g2_antennanp ANTENNA_2767 (.A(net464));
 sg13g2_antennanp ANTENNA_2768 (.A(net464));
 sg13g2_antennanp ANTENNA_2769 (.A(net464));
 sg13g2_antennanp ANTENNA_2770 (.A(net464));
 sg13g2_antennanp ANTENNA_2771 (.A(net464));
 sg13g2_antennanp ANTENNA_2772 (.A(net464));
 sg13g2_antennanp ANTENNA_2773 (.A(net464));
 sg13g2_antennanp ANTENNA_2774 (.A(net464));
 sg13g2_antennanp ANTENNA_2775 (.A(net526));
 sg13g2_antennanp ANTENNA_2776 (.A(net526));
 sg13g2_antennanp ANTENNA_2777 (.A(net526));
 sg13g2_antennanp ANTENNA_2778 (.A(net526));
 sg13g2_antennanp ANTENNA_2779 (.A(net526));
 sg13g2_antennanp ANTENNA_2780 (.A(net526));
 sg13g2_antennanp ANTENNA_2781 (.A(net526));
 sg13g2_antennanp ANTENNA_2782 (.A(net526));
 sg13g2_antennanp ANTENNA_2783 (.A(net526));
 sg13g2_antennanp ANTENNA_2784 (.A(net528));
 sg13g2_antennanp ANTENNA_2785 (.A(net528));
 sg13g2_antennanp ANTENNA_2786 (.A(net528));
 sg13g2_antennanp ANTENNA_2787 (.A(net528));
 sg13g2_antennanp ANTENNA_2788 (.A(net528));
 sg13g2_antennanp ANTENNA_2789 (.A(net528));
 sg13g2_antennanp ANTENNA_2790 (.A(net528));
 sg13g2_antennanp ANTENNA_2791 (.A(net528));
 sg13g2_antennanp ANTENNA_2792 (.A(net528));
 sg13g2_antennanp ANTENNA_2793 (.A(net528));
 sg13g2_antennanp ANTENNA_2794 (.A(net528));
 sg13g2_antennanp ANTENNA_2795 (.A(net528));
 sg13g2_antennanp ANTENNA_2796 (.A(net528));
 sg13g2_antennanp ANTENNA_2797 (.A(net528));
 sg13g2_antennanp ANTENNA_2798 (.A(net528));
 sg13g2_antennanp ANTENNA_2799 (.A(net529));
 sg13g2_antennanp ANTENNA_2800 (.A(net529));
 sg13g2_antennanp ANTENNA_2801 (.A(net529));
 sg13g2_antennanp ANTENNA_2802 (.A(net529));
 sg13g2_antennanp ANTENNA_2803 (.A(net529));
 sg13g2_antennanp ANTENNA_2804 (.A(net529));
 sg13g2_antennanp ANTENNA_2805 (.A(net529));
 sg13g2_antennanp ANTENNA_2806 (.A(net529));
 sg13g2_antennanp ANTENNA_2807 (.A(net529));
 sg13g2_antennanp ANTENNA_2808 (.A(net529));
 sg13g2_antennanp ANTENNA_2809 (.A(net529));
 sg13g2_antennanp ANTENNA_2810 (.A(net529));
 sg13g2_antennanp ANTENNA_2811 (.A(net529));
 sg13g2_antennanp ANTENNA_2812 (.A(net529));
 sg13g2_antennanp ANTENNA_2813 (.A(net529));
 sg13g2_antennanp ANTENNA_2814 (.A(net529));
 sg13g2_antennanp ANTENNA_2815 (.A(net549));
 sg13g2_antennanp ANTENNA_2816 (.A(net549));
 sg13g2_antennanp ANTENNA_2817 (.A(net549));
 sg13g2_antennanp ANTENNA_2818 (.A(net549));
 sg13g2_antennanp ANTENNA_2819 (.A(net549));
 sg13g2_antennanp ANTENNA_2820 (.A(net549));
 sg13g2_antennanp ANTENNA_2821 (.A(net549));
 sg13g2_antennanp ANTENNA_2822 (.A(net549));
 sg13g2_antennanp ANTENNA_2823 (.A(net551));
 sg13g2_antennanp ANTENNA_2824 (.A(net551));
 sg13g2_antennanp ANTENNA_2825 (.A(net551));
 sg13g2_antennanp ANTENNA_2826 (.A(net551));
 sg13g2_antennanp ANTENNA_2827 (.A(net551));
 sg13g2_antennanp ANTENNA_2828 (.A(net551));
 sg13g2_antennanp ANTENNA_2829 (.A(net551));
 sg13g2_antennanp ANTENNA_2830 (.A(net551));
 sg13g2_antennanp ANTENNA_2831 (.A(net551));
 sg13g2_antennanp ANTENNA_2832 (.A(net553));
 sg13g2_antennanp ANTENNA_2833 (.A(net553));
 sg13g2_antennanp ANTENNA_2834 (.A(net553));
 sg13g2_antennanp ANTENNA_2835 (.A(net553));
 sg13g2_antennanp ANTENNA_2836 (.A(net553));
 sg13g2_antennanp ANTENNA_2837 (.A(net553));
 sg13g2_antennanp ANTENNA_2838 (.A(net553));
 sg13g2_antennanp ANTENNA_2839 (.A(net553));
 sg13g2_antennanp ANTENNA_2840 (.A(net553));
 sg13g2_antennanp ANTENNA_2841 (.A(net553));
 sg13g2_antennanp ANTENNA_2842 (.A(net553));
 sg13g2_antennanp ANTENNA_2843 (.A(net553));
 sg13g2_antennanp ANTENNA_2844 (.A(net553));
 sg13g2_antennanp ANTENNA_2845 (.A(net554));
 sg13g2_antennanp ANTENNA_2846 (.A(net554));
 sg13g2_antennanp ANTENNA_2847 (.A(net554));
 sg13g2_antennanp ANTENNA_2848 (.A(net554));
 sg13g2_antennanp ANTENNA_2849 (.A(net554));
 sg13g2_antennanp ANTENNA_2850 (.A(net554));
 sg13g2_antennanp ANTENNA_2851 (.A(net554));
 sg13g2_antennanp ANTENNA_2852 (.A(net554));
 sg13g2_antennanp ANTENNA_2853 (.A(net554));
 sg13g2_antennanp ANTENNA_2854 (.A(net554));
 sg13g2_antennanp ANTENNA_2855 (.A(net554));
 sg13g2_antennanp ANTENNA_2856 (.A(net554));
 sg13g2_antennanp ANTENNA_2857 (.A(net554));
 sg13g2_antennanp ANTENNA_2858 (.A(net554));
 sg13g2_antennanp ANTENNA_2859 (.A(net554));
 sg13g2_antennanp ANTENNA_2860 (.A(net554));
 sg13g2_antennanp ANTENNA_2861 (.A(net568));
 sg13g2_antennanp ANTENNA_2862 (.A(net568));
 sg13g2_antennanp ANTENNA_2863 (.A(net568));
 sg13g2_antennanp ANTENNA_2864 (.A(net568));
 sg13g2_antennanp ANTENNA_2865 (.A(net568));
 sg13g2_antennanp ANTENNA_2866 (.A(net568));
 sg13g2_antennanp ANTENNA_2867 (.A(net568));
 sg13g2_antennanp ANTENNA_2868 (.A(net568));
 sg13g2_antennanp ANTENNA_2869 (.A(net568));
 sg13g2_antennanp ANTENNA_2870 (.A(net641));
 sg13g2_antennanp ANTENNA_2871 (.A(net641));
 sg13g2_antennanp ANTENNA_2872 (.A(net641));
 sg13g2_antennanp ANTENNA_2873 (.A(net641));
 sg13g2_antennanp ANTENNA_2874 (.A(net641));
 sg13g2_antennanp ANTENNA_2875 (.A(net641));
 sg13g2_antennanp ANTENNA_2876 (.A(net641));
 sg13g2_antennanp ANTENNA_2877 (.A(net641));
 sg13g2_antennanp ANTENNA_2878 (.A(net641));
 sg13g2_antennanp ANTENNA_2879 (.A(net697));
 sg13g2_antennanp ANTENNA_2880 (.A(net697));
 sg13g2_antennanp ANTENNA_2881 (.A(net697));
 sg13g2_antennanp ANTENNA_2882 (.A(net697));
 sg13g2_antennanp ANTENNA_2883 (.A(net697));
 sg13g2_antennanp ANTENNA_2884 (.A(net697));
 sg13g2_antennanp ANTENNA_2885 (.A(net697));
 sg13g2_antennanp ANTENNA_2886 (.A(net697));
 sg13g2_antennanp ANTENNA_2887 (.A(net697));
 sg13g2_antennanp ANTENNA_2888 (.A(net770));
 sg13g2_antennanp ANTENNA_2889 (.A(net770));
 sg13g2_antennanp ANTENNA_2890 (.A(net770));
 sg13g2_antennanp ANTENNA_2891 (.A(net770));
 sg13g2_antennanp ANTENNA_2892 (.A(net770));
 sg13g2_antennanp ANTENNA_2893 (.A(net770));
 sg13g2_antennanp ANTENNA_2894 (.A(net770));
 sg13g2_antennanp ANTENNA_2895 (.A(net770));
 sg13g2_antennanp ANTENNA_2896 (.A(net773));
 sg13g2_antennanp ANTENNA_2897 (.A(net773));
 sg13g2_antennanp ANTENNA_2898 (.A(net773));
 sg13g2_antennanp ANTENNA_2899 (.A(net773));
 sg13g2_antennanp ANTENNA_2900 (.A(net773));
 sg13g2_antennanp ANTENNA_2901 (.A(net773));
 sg13g2_antennanp ANTENNA_2902 (.A(net773));
 sg13g2_antennanp ANTENNA_2903 (.A(net773));
 sg13g2_antennanp ANTENNA_2904 (.A(net773));
 sg13g2_antennanp ANTENNA_2905 (.A(net778));
 sg13g2_antennanp ANTENNA_2906 (.A(net778));
 sg13g2_antennanp ANTENNA_2907 (.A(net778));
 sg13g2_antennanp ANTENNA_2908 (.A(net778));
 sg13g2_antennanp ANTENNA_2909 (.A(net778));
 sg13g2_antennanp ANTENNA_2910 (.A(net778));
 sg13g2_antennanp ANTENNA_2911 (.A(net778));
 sg13g2_antennanp ANTENNA_2912 (.A(net778));
 sg13g2_antennanp ANTENNA_2913 (.A(net778));
 sg13g2_antennanp ANTENNA_2914 (.A(net779));
 sg13g2_antennanp ANTENNA_2915 (.A(net779));
 sg13g2_antennanp ANTENNA_2916 (.A(net779));
 sg13g2_antennanp ANTENNA_2917 (.A(net779));
 sg13g2_antennanp ANTENNA_2918 (.A(net779));
 sg13g2_antennanp ANTENNA_2919 (.A(net779));
 sg13g2_antennanp ANTENNA_2920 (.A(net779));
 sg13g2_antennanp ANTENNA_2921 (.A(net779));
 sg13g2_antennanp ANTENNA_2922 (.A(net791));
 sg13g2_antennanp ANTENNA_2923 (.A(net791));
 sg13g2_antennanp ANTENNA_2924 (.A(net791));
 sg13g2_antennanp ANTENNA_2925 (.A(net791));
 sg13g2_antennanp ANTENNA_2926 (.A(net791));
 sg13g2_antennanp ANTENNA_2927 (.A(net791));
 sg13g2_antennanp ANTENNA_2928 (.A(net791));
 sg13g2_antennanp ANTENNA_2929 (.A(net791));
 sg13g2_antennanp ANTENNA_2930 (.A(net791));
 sg13g2_antennanp ANTENNA_2931 (.A(net791));
 sg13g2_antennanp ANTENNA_2932 (.A(net791));
 sg13g2_antennanp ANTENNA_2933 (.A(net791));
 sg13g2_antennanp ANTENNA_2934 (.A(net791));
 sg13g2_antennanp ANTENNA_2935 (.A(net791));
 sg13g2_antennanp ANTENNA_2936 (.A(net791));
 sg13g2_antennanp ANTENNA_2937 (.A(net791));
 sg13g2_antennanp ANTENNA_2938 (.A(net791));
 sg13g2_antennanp ANTENNA_2939 (.A(net791));
 sg13g2_antennanp ANTENNA_2940 (.A(net791));
 sg13g2_antennanp ANTENNA_2941 (.A(net791));
 sg13g2_antennanp ANTENNA_2942 (.A(net802));
 sg13g2_antennanp ANTENNA_2943 (.A(net802));
 sg13g2_antennanp ANTENNA_2944 (.A(net802));
 sg13g2_antennanp ANTENNA_2945 (.A(net802));
 sg13g2_antennanp ANTENNA_2946 (.A(net802));
 sg13g2_antennanp ANTENNA_2947 (.A(net802));
 sg13g2_antennanp ANTENNA_2948 (.A(net802));
 sg13g2_antennanp ANTENNA_2949 (.A(net802));
 sg13g2_antennanp ANTENNA_2950 (.A(net802));
 sg13g2_antennanp ANTENNA_2951 (.A(net838));
 sg13g2_antennanp ANTENNA_2952 (.A(net838));
 sg13g2_antennanp ANTENNA_2953 (.A(net838));
 sg13g2_antennanp ANTENNA_2954 (.A(net838));
 sg13g2_antennanp ANTENNA_2955 (.A(net838));
 sg13g2_antennanp ANTENNA_2956 (.A(net838));
 sg13g2_antennanp ANTENNA_2957 (.A(net838));
 sg13g2_antennanp ANTENNA_2958 (.A(net838));
 sg13g2_antennanp ANTENNA_2959 (.A(net838));
 sg13g2_antennanp ANTENNA_2960 (.A(net839));
 sg13g2_antennanp ANTENNA_2961 (.A(net839));
 sg13g2_antennanp ANTENNA_2962 (.A(net839));
 sg13g2_antennanp ANTENNA_2963 (.A(net839));
 sg13g2_antennanp ANTENNA_2964 (.A(net839));
 sg13g2_antennanp ANTENNA_2965 (.A(net839));
 sg13g2_antennanp ANTENNA_2966 (.A(net839));
 sg13g2_antennanp ANTENNA_2967 (.A(net839));
 sg13g2_antennanp ANTENNA_2968 (.A(net839));
 sg13g2_antennanp ANTENNA_2969 (.A(net878));
 sg13g2_antennanp ANTENNA_2970 (.A(net878));
 sg13g2_antennanp ANTENNA_2971 (.A(net878));
 sg13g2_antennanp ANTENNA_2972 (.A(net878));
 sg13g2_antennanp ANTENNA_2973 (.A(net878));
 sg13g2_antennanp ANTENNA_2974 (.A(net878));
 sg13g2_antennanp ANTENNA_2975 (.A(net878));
 sg13g2_antennanp ANTENNA_2976 (.A(net878));
 sg13g2_antennanp ANTENNA_2977 (.A(net878));
 sg13g2_antennanp ANTENNA_2978 (.A(net878));
 sg13g2_antennanp ANTENNA_2979 (.A(net878));
 sg13g2_antennanp ANTENNA_2980 (.A(net878));
 sg13g2_antennanp ANTENNA_2981 (.A(net878));
 sg13g2_antennanp ANTENNA_2982 (.A(net878));
 sg13g2_antennanp ANTENNA_2983 (.A(net878));
 sg13g2_antennanp ANTENNA_2984 (.A(net878));
 sg13g2_antennanp ANTENNA_2985 (.A(net878));
 sg13g2_antennanp ANTENNA_2986 (.A(net878));
 sg13g2_antennanp ANTENNA_2987 (.A(net878));
 sg13g2_antennanp ANTENNA_2988 (.A(net878));
 sg13g2_antennanp ANTENNA_2989 (.A(net878));
 sg13g2_antennanp ANTENNA_2990 (.A(net878));
 sg13g2_antennanp ANTENNA_2991 (.A(net878));
 sg13g2_antennanp ANTENNA_2992 (.A(net878));
 sg13g2_antennanp ANTENNA_2993 (.A(net878));
 sg13g2_antennanp ANTENNA_2994 (.A(net878));
 sg13g2_antennanp ANTENNA_2995 (.A(net878));
 sg13g2_antennanp ANTENNA_2996 (.A(net878));
 sg13g2_antennanp ANTENNA_2997 (.A(net878));
 sg13g2_antennanp ANTENNA_2998 (.A(net878));
 sg13g2_antennanp ANTENNA_2999 (.A(net878));
 sg13g2_antennanp ANTENNA_3000 (.A(net878));
 sg13g2_antennanp ANTENNA_3001 (.A(net878));
 sg13g2_antennanp ANTENNA_3002 (.A(net878));
 sg13g2_antennanp ANTENNA_3003 (.A(net878));
 sg13g2_antennanp ANTENNA_3004 (.A(net878));
 sg13g2_antennanp ANTENNA_3005 (.A(net878));
 sg13g2_antennanp ANTENNA_3006 (.A(net878));
 sg13g2_antennanp ANTENNA_3007 (.A(net878));
 sg13g2_antennanp ANTENNA_3008 (.A(net878));
 sg13g2_antennanp ANTENNA_3009 (.A(net878));
 sg13g2_antennanp ANTENNA_3010 (.A(net878));
 sg13g2_antennanp ANTENNA_3011 (.A(net878));
 sg13g2_antennanp ANTENNA_3012 (.A(net878));
 sg13g2_antennanp ANTENNA_3013 (.A(net878));
 sg13g2_antennanp ANTENNA_3014 (.A(net878));
 sg13g2_antennanp ANTENNA_3015 (.A(net878));
 sg13g2_antennanp ANTENNA_3016 (.A(net878));
 sg13g2_antennanp ANTENNA_3017 (.A(net924));
 sg13g2_antennanp ANTENNA_3018 (.A(net924));
 sg13g2_antennanp ANTENNA_3019 (.A(net924));
 sg13g2_antennanp ANTENNA_3020 (.A(net924));
 sg13g2_antennanp ANTENNA_3021 (.A(net924));
 sg13g2_antennanp ANTENNA_3022 (.A(net924));
 sg13g2_antennanp ANTENNA_3023 (.A(net924));
 sg13g2_antennanp ANTENNA_3024 (.A(net924));
 sg13g2_antennanp ANTENNA_3025 (.A(net924));
 sg13g2_antennanp ANTENNA_3026 (.A(net982));
 sg13g2_antennanp ANTENNA_3027 (.A(net982));
 sg13g2_antennanp ANTENNA_3028 (.A(net982));
 sg13g2_antennanp ANTENNA_3029 (.A(net982));
 sg13g2_antennanp ANTENNA_3030 (.A(net982));
 sg13g2_antennanp ANTENNA_3031 (.A(net982));
 sg13g2_antennanp ANTENNA_3032 (.A(net982));
 sg13g2_antennanp ANTENNA_3033 (.A(net982));
 sg13g2_antennanp ANTENNA_3034 (.A(net982));
 sg13g2_antennanp ANTENNA_3035 (.A(net982));
 sg13g2_antennanp ANTENNA_3036 (.A(net982));
 sg13g2_antennanp ANTENNA_3037 (.A(net982));
 sg13g2_antennanp ANTENNA_3038 (.A(net982));
 sg13g2_antennanp ANTENNA_3039 (.A(net982));
 sg13g2_antennanp ANTENNA_3040 (.A(net982));
 sg13g2_antennanp ANTENNA_3041 (.A(net982));
 sg13g2_antennanp ANTENNA_3042 (.A(net982));
 sg13g2_antennanp ANTENNA_3043 (.A(net982));
 sg13g2_antennanp ANTENNA_3044 (.A(net982));
 sg13g2_antennanp ANTENNA_3045 (.A(net982));
 sg13g2_antennanp ANTENNA_3046 (.A(net982));
 sg13g2_antennanp ANTENNA_3047 (.A(net982));
 sg13g2_antennanp ANTENNA_3048 (.A(net982));
 sg13g2_antennanp ANTENNA_3049 (.A(net989));
 sg13g2_antennanp ANTENNA_3050 (.A(net989));
 sg13g2_antennanp ANTENNA_3051 (.A(net989));
 sg13g2_antennanp ANTENNA_3052 (.A(net989));
 sg13g2_antennanp ANTENNA_3053 (.A(net989));
 sg13g2_antennanp ANTENNA_3054 (.A(net989));
 sg13g2_antennanp ANTENNA_3055 (.A(net989));
 sg13g2_antennanp ANTENNA_3056 (.A(net989));
 sg13g2_antennanp ANTENNA_3057 (.A(net989));
 sg13g2_antennanp ANTENNA_3058 (.A(net990));
 sg13g2_antennanp ANTENNA_3059 (.A(net990));
 sg13g2_antennanp ANTENNA_3060 (.A(net990));
 sg13g2_antennanp ANTENNA_3061 (.A(net990));
 sg13g2_antennanp ANTENNA_3062 (.A(net990));
 sg13g2_antennanp ANTENNA_3063 (.A(net990));
 sg13g2_antennanp ANTENNA_3064 (.A(net990));
 sg13g2_antennanp ANTENNA_3065 (.A(net990));
 sg13g2_antennanp ANTENNA_3066 (.A(net990));
 sg13g2_antennanp ANTENNA_3067 (.A(net990));
 sg13g2_antennanp ANTENNA_3068 (.A(net990));
 sg13g2_antennanp ANTENNA_3069 (.A(net990));
 sg13g2_antennanp ANTENNA_3070 (.A(net990));
 sg13g2_antennanp ANTENNA_3071 (.A(net990));
 sg13g2_antennanp ANTENNA_3072 (.A(net990));
 sg13g2_antennanp ANTENNA_3073 (.A(net990));
 sg13g2_antennanp ANTENNA_3074 (.A(net990));
 sg13g2_antennanp ANTENNA_3075 (.A(net990));
 sg13g2_antennanp ANTENNA_3076 (.A(net990));
 sg13g2_antennanp ANTENNA_3077 (.A(net990));
 sg13g2_antennanp ANTENNA_3078 (.A(net990));
 sg13g2_antennanp ANTENNA_3079 (.A(net1051));
 sg13g2_antennanp ANTENNA_3080 (.A(net1051));
 sg13g2_antennanp ANTENNA_3081 (.A(net1051));
 sg13g2_antennanp ANTENNA_3082 (.A(net1051));
 sg13g2_antennanp ANTENNA_3083 (.A(net1051));
 sg13g2_antennanp ANTENNA_3084 (.A(net1051));
 sg13g2_antennanp ANTENNA_3085 (.A(net1051));
 sg13g2_antennanp ANTENNA_3086 (.A(net1051));
 sg13g2_antennanp ANTENNA_3087 (.A(net1051));
 sg13g2_antennanp ANTENNA_3088 (.A(net1099));
 sg13g2_antennanp ANTENNA_3089 (.A(net1099));
 sg13g2_antennanp ANTENNA_3090 (.A(net1099));
 sg13g2_antennanp ANTENNA_3091 (.A(net1099));
 sg13g2_antennanp ANTENNA_3092 (.A(net1099));
 sg13g2_antennanp ANTENNA_3093 (.A(net1099));
 sg13g2_antennanp ANTENNA_3094 (.A(net1099));
 sg13g2_antennanp ANTENNA_3095 (.A(net1099));
 sg13g2_antennanp ANTENNA_3096 (.A(net1099));
 sg13g2_antennanp ANTENNA_3097 (.A(net1100));
 sg13g2_antennanp ANTENNA_3098 (.A(net1100));
 sg13g2_antennanp ANTENNA_3099 (.A(net1100));
 sg13g2_antennanp ANTENNA_3100 (.A(net1100));
 sg13g2_antennanp ANTENNA_3101 (.A(net1100));
 sg13g2_antennanp ANTENNA_3102 (.A(net1100));
 sg13g2_antennanp ANTENNA_3103 (.A(net1100));
 sg13g2_antennanp ANTENNA_3104 (.A(net1100));
 sg13g2_antennanp ANTENNA_3105 (.A(net1100));
 sg13g2_antennanp ANTENNA_3106 (.A(net1192));
 sg13g2_antennanp ANTENNA_3107 (.A(net1192));
 sg13g2_antennanp ANTENNA_3108 (.A(net1192));
 sg13g2_antennanp ANTENNA_3109 (.A(net1192));
 sg13g2_antennanp ANTENNA_3110 (.A(net1192));
 sg13g2_antennanp ANTENNA_3111 (.A(net1192));
 sg13g2_antennanp ANTENNA_3112 (.A(net1192));
 sg13g2_antennanp ANTENNA_3113 (.A(net1192));
 sg13g2_antennanp ANTENNA_3114 (.A(net1192));
 sg13g2_antennanp ANTENNA_3115 (.A(net1192));
 sg13g2_antennanp ANTENNA_3116 (.A(net1192));
 sg13g2_antennanp ANTENNA_3117 (.A(net1192));
 sg13g2_antennanp ANTENNA_3118 (.A(net1192));
 sg13g2_antennanp ANTENNA_3119 (.A(net1192));
 sg13g2_antennanp ANTENNA_3120 (.A(net1192));
 sg13g2_antennanp ANTENNA_3121 (.A(net1192));
 sg13g2_antennanp ANTENNA_3122 (.A(net1192));
 sg13g2_antennanp ANTENNA_3123 (.A(net1192));
 sg13g2_antennanp ANTENNA_3124 (.A(net1192));
 sg13g2_antennanp ANTENNA_3125 (.A(net1192));
 sg13g2_antennanp ANTENNA_3126 (.A(net1193));
 sg13g2_antennanp ANTENNA_3127 (.A(net1193));
 sg13g2_antennanp ANTENNA_3128 (.A(net1193));
 sg13g2_antennanp ANTENNA_3129 (.A(net1193));
 sg13g2_antennanp ANTENNA_3130 (.A(net1193));
 sg13g2_antennanp ANTENNA_3131 (.A(net1193));
 sg13g2_antennanp ANTENNA_3132 (.A(net1193));
 sg13g2_antennanp ANTENNA_3133 (.A(net1193));
 sg13g2_antennanp ANTENNA_3134 (.A(net1193));
 sg13g2_antennanp ANTENNA_3135 (.A(net1273));
 sg13g2_antennanp ANTENNA_3136 (.A(net1273));
 sg13g2_antennanp ANTENNA_3137 (.A(net1273));
 sg13g2_antennanp ANTENNA_3138 (.A(net1273));
 sg13g2_antennanp ANTENNA_3139 (.A(net1273));
 sg13g2_antennanp ANTENNA_3140 (.A(net1273));
 sg13g2_antennanp ANTENNA_3141 (.A(net1273));
 sg13g2_antennanp ANTENNA_3142 (.A(net1273));
 sg13g2_antennanp ANTENNA_3143 (.A(net1273));
 sg13g2_antennanp ANTENNA_3144 (.A(net1273));
 sg13g2_antennanp ANTENNA_3145 (.A(net1273));
 sg13g2_antennanp ANTENNA_3146 (.A(net1273));
 sg13g2_antennanp ANTENNA_3147 (.A(net1273));
 sg13g2_antennanp ANTENNA_3148 (.A(net1273));
 sg13g2_antennanp ANTENNA_3149 (.A(net1273));
 sg13g2_antennanp ANTENNA_3150 (.A(net1273));
 sg13g2_antennanp ANTENNA_3151 (.A(net1273));
 sg13g2_antennanp ANTENNA_3152 (.A(net1273));
 sg13g2_antennanp ANTENNA_3153 (.A(net1276));
 sg13g2_antennanp ANTENNA_3154 (.A(net1276));
 sg13g2_antennanp ANTENNA_3155 (.A(net1276));
 sg13g2_antennanp ANTENNA_3156 (.A(net1276));
 sg13g2_antennanp ANTENNA_3157 (.A(net1276));
 sg13g2_antennanp ANTENNA_3158 (.A(net1276));
 sg13g2_antennanp ANTENNA_3159 (.A(net1276));
 sg13g2_antennanp ANTENNA_3160 (.A(net1276));
 sg13g2_antennanp ANTENNA_3161 (.A(net1276));
 sg13g2_antennanp ANTENNA_3162 (.A(net1276));
 sg13g2_antennanp ANTENNA_3163 (.A(net1276));
 sg13g2_antennanp ANTENNA_3164 (.A(net1276));
 sg13g2_antennanp ANTENNA_3165 (.A(net1276));
 sg13g2_antennanp ANTENNA_3166 (.A(_00017_));
 sg13g2_antennanp ANTENNA_3167 (.A(_00017_));
 sg13g2_antennanp ANTENNA_3168 (.A(_00017_));
 sg13g2_antennanp ANTENNA_3169 (.A(_00017_));
 sg13g2_antennanp ANTENNA_3170 (.A(_02490_));
 sg13g2_antennanp ANTENNA_3171 (.A(_03341_));
 sg13g2_antennanp ANTENNA_3172 (.A(_03444_));
 sg13g2_antennanp ANTENNA_3173 (.A(_03444_));
 sg13g2_antennanp ANTENNA_3174 (.A(_03444_));
 sg13g2_antennanp ANTENNA_3175 (.A(_03444_));
 sg13g2_antennanp ANTENNA_3176 (.A(_03621_));
 sg13g2_antennanp ANTENNA_3177 (.A(_03621_));
 sg13g2_antennanp ANTENNA_3178 (.A(_03621_));
 sg13g2_antennanp ANTENNA_3179 (.A(_03621_));
 sg13g2_antennanp ANTENNA_3180 (.A(_03621_));
 sg13g2_antennanp ANTENNA_3181 (.A(_03621_));
 sg13g2_antennanp ANTENNA_3182 (.A(_03621_));
 sg13g2_antennanp ANTENNA_3183 (.A(_03621_));
 sg13g2_antennanp ANTENNA_3184 (.A(_03843_));
 sg13g2_antennanp ANTENNA_3185 (.A(_03843_));
 sg13g2_antennanp ANTENNA_3186 (.A(_03843_));
 sg13g2_antennanp ANTENNA_3187 (.A(_03843_));
 sg13g2_antennanp ANTENNA_3188 (.A(_03875_));
 sg13g2_antennanp ANTENNA_3189 (.A(_03995_));
 sg13g2_antennanp ANTENNA_3190 (.A(_03995_));
 sg13g2_antennanp ANTENNA_3191 (.A(_03995_));
 sg13g2_antennanp ANTENNA_3192 (.A(_03995_));
 sg13g2_antennanp ANTENNA_3193 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3194 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3195 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3196 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3197 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3198 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3199 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3200 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3201 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3202 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3203 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3204 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3205 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3206 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3207 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3208 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3209 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3210 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3211 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3212 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3213 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3214 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3215 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3216 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3217 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3218 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3219 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3220 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3221 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3222 (.A(_04431_));
 sg13g2_antennanp ANTENNA_3223 (.A(_05432_));
 sg13g2_antennanp ANTENNA_3224 (.A(_05432_));
 sg13g2_antennanp ANTENNA_3225 (.A(_05432_));
 sg13g2_antennanp ANTENNA_3226 (.A(_05435_));
 sg13g2_antennanp ANTENNA_3227 (.A(_05441_));
 sg13g2_antennanp ANTENNA_3228 (.A(_05441_));
 sg13g2_antennanp ANTENNA_3229 (.A(_05441_));
 sg13g2_antennanp ANTENNA_3230 (.A(_05441_));
 sg13g2_antennanp ANTENNA_3231 (.A(_05441_));
 sg13g2_antennanp ANTENNA_3232 (.A(_05441_));
 sg13g2_antennanp ANTENNA_3233 (.A(_05449_));
 sg13g2_antennanp ANTENNA_3234 (.A(_05449_));
 sg13g2_antennanp ANTENNA_3235 (.A(_05449_));
 sg13g2_antennanp ANTENNA_3236 (.A(_05449_));
 sg13g2_antennanp ANTENNA_3237 (.A(_05449_));
 sg13g2_antennanp ANTENNA_3238 (.A(_05449_));
 sg13g2_antennanp ANTENNA_3239 (.A(_05457_));
 sg13g2_antennanp ANTENNA_3240 (.A(_05457_));
 sg13g2_antennanp ANTENNA_3241 (.A(_05457_));
 sg13g2_antennanp ANTENNA_3242 (.A(_05457_));
 sg13g2_antennanp ANTENNA_3243 (.A(_05457_));
 sg13g2_antennanp ANTENNA_3244 (.A(_05457_));
 sg13g2_antennanp ANTENNA_3245 (.A(_05463_));
 sg13g2_antennanp ANTENNA_3246 (.A(_05463_));
 sg13g2_antennanp ANTENNA_3247 (.A(_05463_));
 sg13g2_antennanp ANTENNA_3248 (.A(_05463_));
 sg13g2_antennanp ANTENNA_3249 (.A(_05463_));
 sg13g2_antennanp ANTENNA_3250 (.A(_05463_));
 sg13g2_antennanp ANTENNA_3251 (.A(_05463_));
 sg13g2_antennanp ANTENNA_3252 (.A(_05463_));
 sg13g2_antennanp ANTENNA_3253 (.A(_05463_));
 sg13g2_antennanp ANTENNA_3254 (.A(_05467_));
 sg13g2_antennanp ANTENNA_3255 (.A(_05467_));
 sg13g2_antennanp ANTENNA_3256 (.A(_05467_));
 sg13g2_antennanp ANTENNA_3257 (.A(_05471_));
 sg13g2_antennanp ANTENNA_3258 (.A(_05471_));
 sg13g2_antennanp ANTENNA_3259 (.A(_05471_));
 sg13g2_antennanp ANTENNA_3260 (.A(_05471_));
 sg13g2_antennanp ANTENNA_3261 (.A(_05471_));
 sg13g2_antennanp ANTENNA_3262 (.A(_05471_));
 sg13g2_antennanp ANTENNA_3263 (.A(_05471_));
 sg13g2_antennanp ANTENNA_3264 (.A(_05471_));
 sg13g2_antennanp ANTENNA_3265 (.A(_05471_));
 sg13g2_antennanp ANTENNA_3266 (.A(_05476_));
 sg13g2_antennanp ANTENNA_3267 (.A(_05476_));
 sg13g2_antennanp ANTENNA_3268 (.A(_05498_));
 sg13g2_antennanp ANTENNA_3269 (.A(_05498_));
 sg13g2_antennanp ANTENNA_3270 (.A(_06148_));
 sg13g2_antennanp ANTENNA_3271 (.A(_06148_));
 sg13g2_antennanp ANTENNA_3272 (.A(_06148_));
 sg13g2_antennanp ANTENNA_3273 (.A(_06148_));
 sg13g2_antennanp ANTENNA_3274 (.A(_06148_));
 sg13g2_antennanp ANTENNA_3275 (.A(_06171_));
 sg13g2_antennanp ANTENNA_3276 (.A(_06189_));
 sg13g2_antennanp ANTENNA_3277 (.A(_06253_));
 sg13g2_antennanp ANTENNA_3278 (.A(_06253_));
 sg13g2_antennanp ANTENNA_3279 (.A(_06255_));
 sg13g2_antennanp ANTENNA_3280 (.A(_06268_));
 sg13g2_antennanp ANTENNA_3281 (.A(_06293_));
 sg13g2_antennanp ANTENNA_3282 (.A(_06293_));
 sg13g2_antennanp ANTENNA_3283 (.A(_06298_));
 sg13g2_antennanp ANTENNA_3284 (.A(_06298_));
 sg13g2_antennanp ANTENNA_3285 (.A(_06318_));
 sg13g2_antennanp ANTENNA_3286 (.A(_06329_));
 sg13g2_antennanp ANTENNA_3287 (.A(_06416_));
 sg13g2_antennanp ANTENNA_3288 (.A(_06416_));
 sg13g2_antennanp ANTENNA_3289 (.A(_06460_));
 sg13g2_antennanp ANTENNA_3290 (.A(_06493_));
 sg13g2_antennanp ANTENNA_3291 (.A(_06493_));
 sg13g2_antennanp ANTENNA_3292 (.A(_06520_));
 sg13g2_antennanp ANTENNA_3293 (.A(_06559_));
 sg13g2_antennanp ANTENNA_3294 (.A(_06595_));
 sg13g2_antennanp ANTENNA_3295 (.A(_06616_));
 sg13g2_antennanp ANTENNA_3296 (.A(_06620_));
 sg13g2_antennanp ANTENNA_3297 (.A(_06620_));
 sg13g2_antennanp ANTENNA_3298 (.A(_06658_));
 sg13g2_antennanp ANTENNA_3299 (.A(_06694_));
 sg13g2_antennanp ANTENNA_3300 (.A(_06700_));
 sg13g2_antennanp ANTENNA_3301 (.A(_06715_));
 sg13g2_antennanp ANTENNA_3302 (.A(_06719_));
 sg13g2_antennanp ANTENNA_3303 (.A(_06757_));
 sg13g2_antennanp ANTENNA_3304 (.A(_06772_));
 sg13g2_antennanp ANTENNA_3305 (.A(_06772_));
 sg13g2_antennanp ANTENNA_3306 (.A(_06793_));
 sg13g2_antennanp ANTENNA_3307 (.A(_06793_));
 sg13g2_antennanp ANTENNA_3308 (.A(_06799_));
 sg13g2_antennanp ANTENNA_3309 (.A(_06799_));
 sg13g2_antennanp ANTENNA_3310 (.A(_06814_));
 sg13g2_antennanp ANTENNA_3311 (.A(_06818_));
 sg13g2_antennanp ANTENNA_3312 (.A(_06818_));
 sg13g2_antennanp ANTENNA_3313 (.A(_06856_));
 sg13g2_antennanp ANTENNA_3314 (.A(_06871_));
 sg13g2_antennanp ANTENNA_3315 (.A(_06871_));
 sg13g2_antennanp ANTENNA_3316 (.A(_06913_));
 sg13g2_antennanp ANTENNA_3317 (.A(_06955_));
 sg13g2_antennanp ANTENNA_3318 (.A(_06955_));
 sg13g2_antennanp ANTENNA_3319 (.A(_06975_));
 sg13g2_antennanp ANTENNA_3320 (.A(_07012_));
 sg13g2_antennanp ANTENNA_3321 (.A(_07012_));
 sg13g2_antennanp ANTENNA_3322 (.A(_07016_));
 sg13g2_antennanp ANTENNA_3323 (.A(_07054_));
 sg13g2_antennanp ANTENNA_3324 (.A(_07054_));
 sg13g2_antennanp ANTENNA_3325 (.A(_07074_));
 sg13g2_antennanp ANTENNA_3326 (.A(_07074_));
 sg13g2_antennanp ANTENNA_3327 (.A(_07090_));
 sg13g2_antennanp ANTENNA_3328 (.A(_07105_));
 sg13g2_antennanp ANTENNA_3329 (.A(_07105_));
 sg13g2_antennanp ANTENNA_3330 (.A(_07335_));
 sg13g2_antennanp ANTENNA_3331 (.A(_07416_));
 sg13g2_antennanp ANTENNA_3332 (.A(_07416_));
 sg13g2_antennanp ANTENNA_3333 (.A(_07416_));
 sg13g2_antennanp ANTENNA_3334 (.A(_07416_));
 sg13g2_antennanp ANTENNA_3335 (.A(_07416_));
 sg13g2_antennanp ANTENNA_3336 (.A(_07416_));
 sg13g2_antennanp ANTENNA_3337 (.A(_09194_));
 sg13g2_antennanp ANTENNA_3338 (.A(_09194_));
 sg13g2_antennanp ANTENNA_3339 (.A(_09194_));
 sg13g2_antennanp ANTENNA_3340 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3341 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3342 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3343 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3344 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3345 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3346 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3347 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3348 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3349 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3350 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3351 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3352 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3353 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3354 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3355 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3356 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3357 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3358 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3359 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3360 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3361 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3362 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3363 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3364 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3365 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3366 (.A(_09260_));
 sg13g2_antennanp ANTENNA_3367 (.A(_09273_));
 sg13g2_antennanp ANTENNA_3368 (.A(_09273_));
 sg13g2_antennanp ANTENNA_3369 (.A(_09273_));
 sg13g2_antennanp ANTENNA_3370 (.A(_09273_));
 sg13g2_antennanp ANTENNA_3371 (.A(_09273_));
 sg13g2_antennanp ANTENNA_3372 (.A(_09273_));
 sg13g2_antennanp ANTENNA_3373 (.A(_09273_));
 sg13g2_antennanp ANTENNA_3374 (.A(_09273_));
 sg13g2_antennanp ANTENNA_3375 (.A(_09273_));
 sg13g2_antennanp ANTENNA_3376 (.A(_09418_));
 sg13g2_antennanp ANTENNA_3377 (.A(_09418_));
 sg13g2_antennanp ANTENNA_3378 (.A(_09418_));
 sg13g2_antennanp ANTENNA_3379 (.A(_09418_));
 sg13g2_antennanp ANTENNA_3380 (.A(_09418_));
 sg13g2_antennanp ANTENNA_3381 (.A(_09418_));
 sg13g2_antennanp ANTENNA_3382 (.A(_09418_));
 sg13g2_antennanp ANTENNA_3383 (.A(_09418_));
 sg13g2_antennanp ANTENNA_3384 (.A(_09418_));
 sg13g2_antennanp ANTENNA_3385 (.A(_09906_));
 sg13g2_antennanp ANTENNA_3386 (.A(_09906_));
 sg13g2_antennanp ANTENNA_3387 (.A(_09906_));
 sg13g2_antennanp ANTENNA_3388 (.A(_09906_));
 sg13g2_antennanp ANTENNA_3389 (.A(_09906_));
 sg13g2_antennanp ANTENNA_3390 (.A(_09906_));
 sg13g2_antennanp ANTENNA_3391 (.A(_09906_));
 sg13g2_antennanp ANTENNA_3392 (.A(_09906_));
 sg13g2_antennanp ANTENNA_3393 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3394 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3395 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3396 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3397 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3398 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3399 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3400 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3401 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3402 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3403 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3404 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3405 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3406 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3407 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3408 (.A(_09928_));
 sg13g2_antennanp ANTENNA_3409 (.A(_09929_));
 sg13g2_antennanp ANTENNA_3410 (.A(_09929_));
 sg13g2_antennanp ANTENNA_3411 (.A(_09929_));
 sg13g2_antennanp ANTENNA_3412 (.A(_09929_));
 sg13g2_antennanp ANTENNA_3413 (.A(_09935_));
 sg13g2_antennanp ANTENNA_3414 (.A(_09935_));
 sg13g2_antennanp ANTENNA_3415 (.A(_09935_));
 sg13g2_antennanp ANTENNA_3416 (.A(_09935_));
 sg13g2_antennanp ANTENNA_3417 (.A(_09935_));
 sg13g2_antennanp ANTENNA_3418 (.A(_09935_));
 sg13g2_antennanp ANTENNA_3419 (.A(_09935_));
 sg13g2_antennanp ANTENNA_3420 (.A(_09935_));
 sg13g2_antennanp ANTENNA_3421 (.A(_09935_));
 sg13g2_antennanp ANTENNA_3422 (.A(_10040_));
 sg13g2_antennanp ANTENNA_3423 (.A(_10040_));
 sg13g2_antennanp ANTENNA_3424 (.A(_10040_));
 sg13g2_antennanp ANTENNA_3425 (.A(_10040_));
 sg13g2_antennanp ANTENNA_3426 (.A(_10040_));
 sg13g2_antennanp ANTENNA_3427 (.A(_10040_));
 sg13g2_antennanp ANTENNA_3428 (.A(_10042_));
 sg13g2_antennanp ANTENNA_3429 (.A(_10042_));
 sg13g2_antennanp ANTENNA_3430 (.A(_10042_));
 sg13g2_antennanp ANTENNA_3431 (.A(_10042_));
 sg13g2_antennanp ANTENNA_3432 (.A(_10046_));
 sg13g2_antennanp ANTENNA_3433 (.A(_10048_));
 sg13g2_antennanp ANTENNA_3434 (.A(_10051_));
 sg13g2_antennanp ANTENNA_3435 (.A(_10053_));
 sg13g2_antennanp ANTENNA_3436 (.A(_10071_));
 sg13g2_antennanp ANTENNA_3437 (.A(_10071_));
 sg13g2_antennanp ANTENNA_3438 (.A(_10071_));
 sg13g2_antennanp ANTENNA_3439 (.A(_10071_));
 sg13g2_antennanp ANTENNA_3440 (.A(_10083_));
 sg13g2_antennanp ANTENNA_3441 (.A(_10092_));
 sg13g2_antennanp ANTENNA_3442 (.A(_10092_));
 sg13g2_antennanp ANTENNA_3443 (.A(_10092_));
 sg13g2_antennanp ANTENNA_3444 (.A(_10101_));
 sg13g2_antennanp ANTENNA_3445 (.A(_10106_));
 sg13g2_antennanp ANTENNA_3446 (.A(_10110_));
 sg13g2_antennanp ANTENNA_3447 (.A(_10131_));
 sg13g2_antennanp ANTENNA_3448 (.A(_10131_));
 sg13g2_antennanp ANTENNA_3449 (.A(_10136_));
 sg13g2_antennanp ANTENNA_3450 (.A(_10140_));
 sg13g2_antennanp ANTENNA_3451 (.A(_10226_));
 sg13g2_antennanp ANTENNA_3452 (.A(_10226_));
 sg13g2_antennanp ANTENNA_3453 (.A(_10226_));
 sg13g2_antennanp ANTENNA_3454 (.A(_10243_));
 sg13g2_antennanp ANTENNA_3455 (.A(_10243_));
 sg13g2_antennanp ANTENNA_3456 (.A(_10243_));
 sg13g2_antennanp ANTENNA_3457 (.A(_10243_));
 sg13g2_antennanp ANTENNA_3458 (.A(_10243_));
 sg13g2_antennanp ANTENNA_3459 (.A(_10243_));
 sg13g2_antennanp ANTENNA_3460 (.A(_10256_));
 sg13g2_antennanp ANTENNA_3461 (.A(_10256_));
 sg13g2_antennanp ANTENNA_3462 (.A(_10256_));
 sg13g2_antennanp ANTENNA_3463 (.A(_10256_));
 sg13g2_antennanp ANTENNA_3464 (.A(_10256_));
 sg13g2_antennanp ANTENNA_3465 (.A(_10287_));
 sg13g2_antennanp ANTENNA_3466 (.A(_10287_));
 sg13g2_antennanp ANTENNA_3467 (.A(_10287_));
 sg13g2_antennanp ANTENNA_3468 (.A(_10287_));
 sg13g2_antennanp ANTENNA_3469 (.A(_10295_));
 sg13g2_antennanp ANTENNA_3470 (.A(_10295_));
 sg13g2_antennanp ANTENNA_3471 (.A(_10295_));
 sg13g2_antennanp ANTENNA_3472 (.A(_10295_));
 sg13g2_antennanp ANTENNA_3473 (.A(_10295_));
 sg13g2_antennanp ANTENNA_3474 (.A(_10295_));
 sg13g2_antennanp ANTENNA_3475 (.A(_10295_));
 sg13g2_antennanp ANTENNA_3476 (.A(_10295_));
 sg13g2_antennanp ANTENNA_3477 (.A(_10296_));
 sg13g2_antennanp ANTENNA_3478 (.A(_10296_));
 sg13g2_antennanp ANTENNA_3479 (.A(_10296_));
 sg13g2_antennanp ANTENNA_3480 (.A(_10296_));
 sg13g2_antennanp ANTENNA_3481 (.A(_10296_));
 sg13g2_antennanp ANTENNA_3482 (.A(_10325_));
 sg13g2_antennanp ANTENNA_3483 (.A(_10325_));
 sg13g2_antennanp ANTENNA_3484 (.A(_10325_));
 sg13g2_antennanp ANTENNA_3485 (.A(_10325_));
 sg13g2_antennanp ANTENNA_3486 (.A(_10325_));
 sg13g2_antennanp ANTENNA_3487 (.A(_10325_));
 sg13g2_antennanp ANTENNA_3488 (.A(_10325_));
 sg13g2_antennanp ANTENNA_3489 (.A(_10325_));
 sg13g2_antennanp ANTENNA_3490 (.A(_10326_));
 sg13g2_antennanp ANTENNA_3491 (.A(_10326_));
 sg13g2_antennanp ANTENNA_3492 (.A(_10326_));
 sg13g2_antennanp ANTENNA_3493 (.A(_10349_));
 sg13g2_antennanp ANTENNA_3494 (.A(_10349_));
 sg13g2_antennanp ANTENNA_3495 (.A(_10349_));
 sg13g2_antennanp ANTENNA_3496 (.A(_10349_));
 sg13g2_antennanp ANTENNA_3497 (.A(_10350_));
 sg13g2_antennanp ANTENNA_3498 (.A(_10350_));
 sg13g2_antennanp ANTENNA_3499 (.A(_10350_));
 sg13g2_antennanp ANTENNA_3500 (.A(_10350_));
 sg13g2_antennanp ANTENNA_3501 (.A(_10350_));
 sg13g2_antennanp ANTENNA_3502 (.A(_10350_));
 sg13g2_antennanp ANTENNA_3503 (.A(_10397_));
 sg13g2_antennanp ANTENNA_3504 (.A(_10397_));
 sg13g2_antennanp ANTENNA_3505 (.A(_10397_));
 sg13g2_antennanp ANTENNA_3506 (.A(_10397_));
 sg13g2_antennanp ANTENNA_3507 (.A(_10397_));
 sg13g2_antennanp ANTENNA_3508 (.A(_10397_));
 sg13g2_antennanp ANTENNA_3509 (.A(_10397_));
 sg13g2_antennanp ANTENNA_3510 (.A(_10397_));
 sg13g2_antennanp ANTENNA_3511 (.A(_10397_));
 sg13g2_antennanp ANTENNA_3512 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3513 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3514 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3515 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3516 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3517 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3518 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3519 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3520 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3521 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3522 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3523 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3524 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3525 (.A(_10422_));
 sg13g2_antennanp ANTENNA_3526 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3527 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3528 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3529 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3530 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3531 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3532 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3533 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3534 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3535 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3536 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3537 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3538 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3539 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3540 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3541 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3542 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3543 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3544 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3545 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3546 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3547 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3548 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3549 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3550 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3551 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3552 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3553 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3554 (.A(_10444_));
 sg13g2_antennanp ANTENNA_3555 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3556 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3557 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3558 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3559 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3560 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3561 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3562 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3563 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3564 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3565 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3566 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3567 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3568 (.A(_10564_));
 sg13g2_antennanp ANTENNA_3569 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3570 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3571 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3572 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3573 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3574 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3575 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3576 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3577 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3578 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3579 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3580 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3581 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3582 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3583 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3584 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3585 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3586 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3587 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3588 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3589 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3590 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3591 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3592 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3593 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3594 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3595 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3596 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3597 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3598 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3599 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3600 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3601 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3602 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3603 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3604 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3605 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3606 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3607 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3608 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3609 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3610 (.A(_10586_));
 sg13g2_antennanp ANTENNA_3611 (.A(_10632_));
 sg13g2_antennanp ANTENNA_3612 (.A(_10632_));
 sg13g2_antennanp ANTENNA_3613 (.A(_10632_));
 sg13g2_antennanp ANTENNA_3614 (.A(_10632_));
 sg13g2_antennanp ANTENNA_3615 (.A(_10632_));
 sg13g2_antennanp ANTENNA_3616 (.A(_10632_));
 sg13g2_antennanp ANTENNA_3617 (.A(_10632_));
 sg13g2_antennanp ANTENNA_3618 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3619 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3620 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3621 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3622 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3623 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3624 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3625 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3626 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3627 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3628 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3629 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3630 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3631 (.A(_10656_));
 sg13g2_antennanp ANTENNA_3632 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3633 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3634 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3635 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3636 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3637 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3638 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3639 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3640 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3641 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3642 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3643 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3644 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3645 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3646 (.A(_10679_));
 sg13g2_antennanp ANTENNA_3647 (.A(_10680_));
 sg13g2_antennanp ANTENNA_3648 (.A(_10680_));
 sg13g2_antennanp ANTENNA_3649 (.A(_10680_));
 sg13g2_antennanp ANTENNA_3650 (.A(_11875_));
 sg13g2_antennanp ANTENNA_3651 (.A(_11875_));
 sg13g2_antennanp ANTENNA_3652 (.A(_11875_));
 sg13g2_antennanp ANTENNA_3653 (.A(_11875_));
 sg13g2_antennanp ANTENNA_3654 (.A(_11875_));
 sg13g2_antennanp ANTENNA_3655 (.A(_11875_));
 sg13g2_antennanp ANTENNA_3656 (.A(_11875_));
 sg13g2_antennanp ANTENNA_3657 (.A(_11947_));
 sg13g2_antennanp ANTENNA_3658 (.A(_11947_));
 sg13g2_antennanp ANTENNA_3659 (.A(_11947_));
 sg13g2_antennanp ANTENNA_3660 (.A(_11947_));
 sg13g2_antennanp ANTENNA_3661 (.A(_12437_));
 sg13g2_antennanp ANTENNA_3662 (.A(_12437_));
 sg13g2_antennanp ANTENNA_3663 (.A(_12437_));
 sg13g2_antennanp ANTENNA_3664 (.A(_12437_));
 sg13g2_antennanp ANTENNA_3665 (.A(_12440_));
 sg13g2_antennanp ANTENNA_3666 (.A(_12440_));
 sg13g2_antennanp ANTENNA_3667 (.A(_12440_));
 sg13g2_antennanp ANTENNA_3668 (.A(_12630_));
 sg13g2_antennanp ANTENNA_3669 (.A(_12630_));
 sg13g2_antennanp ANTENNA_3670 (.A(_12630_));
 sg13g2_antennanp ANTENNA_3671 (.A(_12630_));
 sg13g2_antennanp ANTENNA_3672 (.A(_12653_));
 sg13g2_antennanp ANTENNA_3673 (.A(_12653_));
 sg13g2_antennanp ANTENNA_3674 (.A(_12653_));
 sg13g2_antennanp ANTENNA_3675 (.A(_12653_));
 sg13g2_antennanp ANTENNA_3676 (.A(_12653_));
 sg13g2_antennanp ANTENNA_3677 (.A(_12653_));
 sg13g2_antennanp ANTENNA_3678 (.A(_12653_));
 sg13g2_antennanp ANTENNA_3679 (.A(clk));
 sg13g2_antennanp ANTENNA_3680 (.A(clk));
 sg13g2_antennanp ANTENNA_3681 (.A(\mem.data_in[1] ));
 sg13g2_antennanp ANTENNA_3682 (.A(\mem.data_in[1] ));
 sg13g2_antennanp ANTENNA_3683 (.A(\mem.io_data_out[3] ));
 sg13g2_antennanp ANTENNA_3684 (.A(\mem.io_data_out[3] ));
 sg13g2_antennanp ANTENNA_3685 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_3686 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_3687 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_3688 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_3689 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_3690 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_3691 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_3692 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_3693 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_3694 (.A(net1));
 sg13g2_antennanp ANTENNA_3695 (.A(net1));
 sg13g2_antennanp ANTENNA_3696 (.A(net1));
 sg13g2_antennanp ANTENNA_3697 (.A(net464));
 sg13g2_antennanp ANTENNA_3698 (.A(net464));
 sg13g2_antennanp ANTENNA_3699 (.A(net464));
 sg13g2_antennanp ANTENNA_3700 (.A(net464));
 sg13g2_antennanp ANTENNA_3701 (.A(net464));
 sg13g2_antennanp ANTENNA_3702 (.A(net464));
 sg13g2_antennanp ANTENNA_3703 (.A(net464));
 sg13g2_antennanp ANTENNA_3704 (.A(net464));
 sg13g2_antennanp ANTENNA_3705 (.A(net464));
 sg13g2_antennanp ANTENNA_3706 (.A(net526));
 sg13g2_antennanp ANTENNA_3707 (.A(net526));
 sg13g2_antennanp ANTENNA_3708 (.A(net526));
 sg13g2_antennanp ANTENNA_3709 (.A(net526));
 sg13g2_antennanp ANTENNA_3710 (.A(net526));
 sg13g2_antennanp ANTENNA_3711 (.A(net526));
 sg13g2_antennanp ANTENNA_3712 (.A(net526));
 sg13g2_antennanp ANTENNA_3713 (.A(net526));
 sg13g2_antennanp ANTENNA_3714 (.A(net526));
 sg13g2_antennanp ANTENNA_3715 (.A(net526));
 sg13g2_antennanp ANTENNA_3716 (.A(net526));
 sg13g2_antennanp ANTENNA_3717 (.A(net526));
 sg13g2_antennanp ANTENNA_3718 (.A(net526));
 sg13g2_antennanp ANTENNA_3719 (.A(net549));
 sg13g2_antennanp ANTENNA_3720 (.A(net549));
 sg13g2_antennanp ANTENNA_3721 (.A(net549));
 sg13g2_antennanp ANTENNA_3722 (.A(net549));
 sg13g2_antennanp ANTENNA_3723 (.A(net549));
 sg13g2_antennanp ANTENNA_3724 (.A(net549));
 sg13g2_antennanp ANTENNA_3725 (.A(net549));
 sg13g2_antennanp ANTENNA_3726 (.A(net549));
 sg13g2_antennanp ANTENNA_3727 (.A(net553));
 sg13g2_antennanp ANTENNA_3728 (.A(net553));
 sg13g2_antennanp ANTENNA_3729 (.A(net553));
 sg13g2_antennanp ANTENNA_3730 (.A(net553));
 sg13g2_antennanp ANTENNA_3731 (.A(net553));
 sg13g2_antennanp ANTENNA_3732 (.A(net553));
 sg13g2_antennanp ANTENNA_3733 (.A(net553));
 sg13g2_antennanp ANTENNA_3734 (.A(net553));
 sg13g2_antennanp ANTENNA_3735 (.A(net553));
 sg13g2_antennanp ANTENNA_3736 (.A(net553));
 sg13g2_antennanp ANTENNA_3737 (.A(net553));
 sg13g2_antennanp ANTENNA_3738 (.A(net553));
 sg13g2_antennanp ANTENNA_3739 (.A(net553));
 sg13g2_antennanp ANTENNA_3740 (.A(net553));
 sg13g2_antennanp ANTENNA_3741 (.A(net554));
 sg13g2_antennanp ANTENNA_3742 (.A(net554));
 sg13g2_antennanp ANTENNA_3743 (.A(net554));
 sg13g2_antennanp ANTENNA_3744 (.A(net554));
 sg13g2_antennanp ANTENNA_3745 (.A(net554));
 sg13g2_antennanp ANTENNA_3746 (.A(net554));
 sg13g2_antennanp ANTENNA_3747 (.A(net554));
 sg13g2_antennanp ANTENNA_3748 (.A(net554));
 sg13g2_antennanp ANTENNA_3749 (.A(net554));
 sg13g2_antennanp ANTENNA_3750 (.A(net554));
 sg13g2_antennanp ANTENNA_3751 (.A(net554));
 sg13g2_antennanp ANTENNA_3752 (.A(net554));
 sg13g2_antennanp ANTENNA_3753 (.A(net554));
 sg13g2_antennanp ANTENNA_3754 (.A(net554));
 sg13g2_antennanp ANTENNA_3755 (.A(net554));
 sg13g2_antennanp ANTENNA_3756 (.A(net554));
 sg13g2_antennanp ANTENNA_3757 (.A(net554));
 sg13g2_antennanp ANTENNA_3758 (.A(net554));
 sg13g2_antennanp ANTENNA_3759 (.A(net554));
 sg13g2_antennanp ANTENNA_3760 (.A(net554));
 sg13g2_antennanp ANTENNA_3761 (.A(net554));
 sg13g2_antennanp ANTENNA_3762 (.A(net554));
 sg13g2_antennanp ANTENNA_3763 (.A(net554));
 sg13g2_antennanp ANTENNA_3764 (.A(net554));
 sg13g2_antennanp ANTENNA_3765 (.A(net554));
 sg13g2_antennanp ANTENNA_3766 (.A(net554));
 sg13g2_antennanp ANTENNA_3767 (.A(net554));
 sg13g2_antennanp ANTENNA_3768 (.A(net554));
 sg13g2_antennanp ANTENNA_3769 (.A(net556));
 sg13g2_antennanp ANTENNA_3770 (.A(net556));
 sg13g2_antennanp ANTENNA_3771 (.A(net556));
 sg13g2_antennanp ANTENNA_3772 (.A(net556));
 sg13g2_antennanp ANTENNA_3773 (.A(net556));
 sg13g2_antennanp ANTENNA_3774 (.A(net556));
 sg13g2_antennanp ANTENNA_3775 (.A(net556));
 sg13g2_antennanp ANTENNA_3776 (.A(net556));
 sg13g2_antennanp ANTENNA_3777 (.A(net556));
 sg13g2_antennanp ANTENNA_3778 (.A(net556));
 sg13g2_antennanp ANTENNA_3779 (.A(net556));
 sg13g2_antennanp ANTENNA_3780 (.A(net556));
 sg13g2_antennanp ANTENNA_3781 (.A(net556));
 sg13g2_antennanp ANTENNA_3782 (.A(net556));
 sg13g2_antennanp ANTENNA_3783 (.A(net556));
 sg13g2_antennanp ANTENNA_3784 (.A(net556));
 sg13g2_antennanp ANTENNA_3785 (.A(net641));
 sg13g2_antennanp ANTENNA_3786 (.A(net641));
 sg13g2_antennanp ANTENNA_3787 (.A(net641));
 sg13g2_antennanp ANTENNA_3788 (.A(net641));
 sg13g2_antennanp ANTENNA_3789 (.A(net641));
 sg13g2_antennanp ANTENNA_3790 (.A(net641));
 sg13g2_antennanp ANTENNA_3791 (.A(net641));
 sg13g2_antennanp ANTENNA_3792 (.A(net641));
 sg13g2_antennanp ANTENNA_3793 (.A(net641));
 sg13g2_antennanp ANTENNA_3794 (.A(net770));
 sg13g2_antennanp ANTENNA_3795 (.A(net770));
 sg13g2_antennanp ANTENNA_3796 (.A(net770));
 sg13g2_antennanp ANTENNA_3797 (.A(net770));
 sg13g2_antennanp ANTENNA_3798 (.A(net770));
 sg13g2_antennanp ANTENNA_3799 (.A(net770));
 sg13g2_antennanp ANTENNA_3800 (.A(net770));
 sg13g2_antennanp ANTENNA_3801 (.A(net770));
 sg13g2_antennanp ANTENNA_3802 (.A(net770));
 sg13g2_antennanp ANTENNA_3803 (.A(net770));
 sg13g2_antennanp ANTENNA_3804 (.A(net770));
 sg13g2_antennanp ANTENNA_3805 (.A(net770));
 sg13g2_antennanp ANTENNA_3806 (.A(net770));
 sg13g2_antennanp ANTENNA_3807 (.A(net778));
 sg13g2_antennanp ANTENNA_3808 (.A(net778));
 sg13g2_antennanp ANTENNA_3809 (.A(net778));
 sg13g2_antennanp ANTENNA_3810 (.A(net778));
 sg13g2_antennanp ANTENNA_3811 (.A(net778));
 sg13g2_antennanp ANTENNA_3812 (.A(net778));
 sg13g2_antennanp ANTENNA_3813 (.A(net778));
 sg13g2_antennanp ANTENNA_3814 (.A(net778));
 sg13g2_antennanp ANTENNA_3815 (.A(net779));
 sg13g2_antennanp ANTENNA_3816 (.A(net779));
 sg13g2_antennanp ANTENNA_3817 (.A(net779));
 sg13g2_antennanp ANTENNA_3818 (.A(net779));
 sg13g2_antennanp ANTENNA_3819 (.A(net779));
 sg13g2_antennanp ANTENNA_3820 (.A(net779));
 sg13g2_antennanp ANTENNA_3821 (.A(net779));
 sg13g2_antennanp ANTENNA_3822 (.A(net779));
 sg13g2_antennanp ANTENNA_3823 (.A(net792));
 sg13g2_antennanp ANTENNA_3824 (.A(net792));
 sg13g2_antennanp ANTENNA_3825 (.A(net792));
 sg13g2_antennanp ANTENNA_3826 (.A(net792));
 sg13g2_antennanp ANTENNA_3827 (.A(net792));
 sg13g2_antennanp ANTENNA_3828 (.A(net792));
 sg13g2_antennanp ANTENNA_3829 (.A(net792));
 sg13g2_antennanp ANTENNA_3830 (.A(net792));
 sg13g2_antennanp ANTENNA_3831 (.A(net802));
 sg13g2_antennanp ANTENNA_3832 (.A(net802));
 sg13g2_antennanp ANTENNA_3833 (.A(net802));
 sg13g2_antennanp ANTENNA_3834 (.A(net802));
 sg13g2_antennanp ANTENNA_3835 (.A(net802));
 sg13g2_antennanp ANTENNA_3836 (.A(net802));
 sg13g2_antennanp ANTENNA_3837 (.A(net802));
 sg13g2_antennanp ANTENNA_3838 (.A(net802));
 sg13g2_antennanp ANTENNA_3839 (.A(net802));
 sg13g2_antennanp ANTENNA_3840 (.A(net838));
 sg13g2_antennanp ANTENNA_3841 (.A(net838));
 sg13g2_antennanp ANTENNA_3842 (.A(net838));
 sg13g2_antennanp ANTENNA_3843 (.A(net838));
 sg13g2_antennanp ANTENNA_3844 (.A(net838));
 sg13g2_antennanp ANTENNA_3845 (.A(net838));
 sg13g2_antennanp ANTENNA_3846 (.A(net838));
 sg13g2_antennanp ANTENNA_3847 (.A(net838));
 sg13g2_antennanp ANTENNA_3848 (.A(net838));
 sg13g2_antennanp ANTENNA_3849 (.A(net878));
 sg13g2_antennanp ANTENNA_3850 (.A(net878));
 sg13g2_antennanp ANTENNA_3851 (.A(net878));
 sg13g2_antennanp ANTENNA_3852 (.A(net878));
 sg13g2_antennanp ANTENNA_3853 (.A(net878));
 sg13g2_antennanp ANTENNA_3854 (.A(net878));
 sg13g2_antennanp ANTENNA_3855 (.A(net878));
 sg13g2_antennanp ANTENNA_3856 (.A(net878));
 sg13g2_antennanp ANTENNA_3857 (.A(net878));
 sg13g2_antennanp ANTENNA_3858 (.A(net878));
 sg13g2_antennanp ANTENNA_3859 (.A(net878));
 sg13g2_antennanp ANTENNA_3860 (.A(net878));
 sg13g2_antennanp ANTENNA_3861 (.A(net878));
 sg13g2_antennanp ANTENNA_3862 (.A(net878));
 sg13g2_antennanp ANTENNA_3863 (.A(net878));
 sg13g2_antennanp ANTENNA_3864 (.A(net878));
 sg13g2_antennanp ANTENNA_3865 (.A(net878));
 sg13g2_antennanp ANTENNA_3866 (.A(net878));
 sg13g2_antennanp ANTENNA_3867 (.A(net878));
 sg13g2_antennanp ANTENNA_3868 (.A(net878));
 sg13g2_antennanp ANTENNA_3869 (.A(net878));
 sg13g2_antennanp ANTENNA_3870 (.A(net878));
 sg13g2_antennanp ANTENNA_3871 (.A(net878));
 sg13g2_antennanp ANTENNA_3872 (.A(net878));
 sg13g2_antennanp ANTENNA_3873 (.A(net878));
 sg13g2_antennanp ANTENNA_3874 (.A(net878));
 sg13g2_antennanp ANTENNA_3875 (.A(net878));
 sg13g2_antennanp ANTENNA_3876 (.A(net878));
 sg13g2_antennanp ANTENNA_3877 (.A(net878));
 sg13g2_antennanp ANTENNA_3878 (.A(net878));
 sg13g2_antennanp ANTENNA_3879 (.A(net878));
 sg13g2_antennanp ANTENNA_3880 (.A(net878));
 sg13g2_antennanp ANTENNA_3881 (.A(net878));
 sg13g2_antennanp ANTENNA_3882 (.A(net878));
 sg13g2_antennanp ANTENNA_3883 (.A(net878));
 sg13g2_antennanp ANTENNA_3884 (.A(net878));
 sg13g2_antennanp ANTENNA_3885 (.A(net878));
 sg13g2_antennanp ANTENNA_3886 (.A(net878));
 sg13g2_antennanp ANTENNA_3887 (.A(net878));
 sg13g2_antennanp ANTENNA_3888 (.A(net878));
 sg13g2_antennanp ANTENNA_3889 (.A(net878));
 sg13g2_antennanp ANTENNA_3890 (.A(net878));
 sg13g2_antennanp ANTENNA_3891 (.A(net878));
 sg13g2_antennanp ANTENNA_3892 (.A(net878));
 sg13g2_antennanp ANTENNA_3893 (.A(net878));
 sg13g2_antennanp ANTENNA_3894 (.A(net878));
 sg13g2_antennanp ANTENNA_3895 (.A(net878));
 sg13g2_antennanp ANTENNA_3896 (.A(net878));
 sg13g2_antennanp ANTENNA_3897 (.A(net924));
 sg13g2_antennanp ANTENNA_3898 (.A(net924));
 sg13g2_antennanp ANTENNA_3899 (.A(net924));
 sg13g2_antennanp ANTENNA_3900 (.A(net924));
 sg13g2_antennanp ANTENNA_3901 (.A(net924));
 sg13g2_antennanp ANTENNA_3902 (.A(net924));
 sg13g2_antennanp ANTENNA_3903 (.A(net924));
 sg13g2_antennanp ANTENNA_3904 (.A(net924));
 sg13g2_antennanp ANTENNA_3905 (.A(net924));
 sg13g2_antennanp ANTENNA_3906 (.A(net982));
 sg13g2_antennanp ANTENNA_3907 (.A(net982));
 sg13g2_antennanp ANTENNA_3908 (.A(net982));
 sg13g2_antennanp ANTENNA_3909 (.A(net982));
 sg13g2_antennanp ANTENNA_3910 (.A(net982));
 sg13g2_antennanp ANTENNA_3911 (.A(net982));
 sg13g2_antennanp ANTENNA_3912 (.A(net982));
 sg13g2_antennanp ANTENNA_3913 (.A(net982));
 sg13g2_antennanp ANTENNA_3914 (.A(net982));
 sg13g2_antennanp ANTENNA_3915 (.A(net989));
 sg13g2_antennanp ANTENNA_3916 (.A(net989));
 sg13g2_antennanp ANTENNA_3917 (.A(net989));
 sg13g2_antennanp ANTENNA_3918 (.A(net989));
 sg13g2_antennanp ANTENNA_3919 (.A(net989));
 sg13g2_antennanp ANTENNA_3920 (.A(net989));
 sg13g2_antennanp ANTENNA_3921 (.A(net989));
 sg13g2_antennanp ANTENNA_3922 (.A(net989));
 sg13g2_antennanp ANTENNA_3923 (.A(net989));
 sg13g2_antennanp ANTENNA_3924 (.A(net990));
 sg13g2_antennanp ANTENNA_3925 (.A(net990));
 sg13g2_antennanp ANTENNA_3926 (.A(net990));
 sg13g2_antennanp ANTENNA_3927 (.A(net990));
 sg13g2_antennanp ANTENNA_3928 (.A(net990));
 sg13g2_antennanp ANTENNA_3929 (.A(net990));
 sg13g2_antennanp ANTENNA_3930 (.A(net990));
 sg13g2_antennanp ANTENNA_3931 (.A(net990));
 sg13g2_antennanp ANTENNA_3932 (.A(net990));
 sg13g2_antennanp ANTENNA_3933 (.A(net1051));
 sg13g2_antennanp ANTENNA_3934 (.A(net1051));
 sg13g2_antennanp ANTENNA_3935 (.A(net1051));
 sg13g2_antennanp ANTENNA_3936 (.A(net1051));
 sg13g2_antennanp ANTENNA_3937 (.A(net1051));
 sg13g2_antennanp ANTENNA_3938 (.A(net1051));
 sg13g2_antennanp ANTENNA_3939 (.A(net1051));
 sg13g2_antennanp ANTENNA_3940 (.A(net1051));
 sg13g2_antennanp ANTENNA_3941 (.A(net1051));
 sg13g2_antennanp ANTENNA_3942 (.A(net1053));
 sg13g2_antennanp ANTENNA_3943 (.A(net1053));
 sg13g2_antennanp ANTENNA_3944 (.A(net1053));
 sg13g2_antennanp ANTENNA_3945 (.A(net1053));
 sg13g2_antennanp ANTENNA_3946 (.A(net1053));
 sg13g2_antennanp ANTENNA_3947 (.A(net1053));
 sg13g2_antennanp ANTENNA_3948 (.A(net1053));
 sg13g2_antennanp ANTENNA_3949 (.A(net1053));
 sg13g2_antennanp ANTENNA_3950 (.A(net1054));
 sg13g2_antennanp ANTENNA_3951 (.A(net1054));
 sg13g2_antennanp ANTENNA_3952 (.A(net1054));
 sg13g2_antennanp ANTENNA_3953 (.A(net1054));
 sg13g2_antennanp ANTENNA_3954 (.A(net1054));
 sg13g2_antennanp ANTENNA_3955 (.A(net1054));
 sg13g2_antennanp ANTENNA_3956 (.A(net1054));
 sg13g2_antennanp ANTENNA_3957 (.A(net1054));
 sg13g2_antennanp ANTENNA_3958 (.A(net1099));
 sg13g2_antennanp ANTENNA_3959 (.A(net1099));
 sg13g2_antennanp ANTENNA_3960 (.A(net1099));
 sg13g2_antennanp ANTENNA_3961 (.A(net1099));
 sg13g2_antennanp ANTENNA_3962 (.A(net1099));
 sg13g2_antennanp ANTENNA_3963 (.A(net1099));
 sg13g2_antennanp ANTENNA_3964 (.A(net1099));
 sg13g2_antennanp ANTENNA_3965 (.A(net1099));
 sg13g2_antennanp ANTENNA_3966 (.A(net1192));
 sg13g2_antennanp ANTENNA_3967 (.A(net1192));
 sg13g2_antennanp ANTENNA_3968 (.A(net1192));
 sg13g2_antennanp ANTENNA_3969 (.A(net1192));
 sg13g2_antennanp ANTENNA_3970 (.A(net1192));
 sg13g2_antennanp ANTENNA_3971 (.A(net1192));
 sg13g2_antennanp ANTENNA_3972 (.A(net1192));
 sg13g2_antennanp ANTENNA_3973 (.A(net1192));
 sg13g2_antennanp ANTENNA_3974 (.A(net1192));
 sg13g2_antennanp ANTENNA_3975 (.A(net1192));
 sg13g2_antennanp ANTENNA_3976 (.A(net1192));
 sg13g2_antennanp ANTENNA_3977 (.A(net1192));
 sg13g2_antennanp ANTENNA_3978 (.A(net1192));
 sg13g2_antennanp ANTENNA_3979 (.A(net1192));
 sg13g2_antennanp ANTENNA_3980 (.A(net1192));
 sg13g2_antennanp ANTENNA_3981 (.A(net1192));
 sg13g2_antennanp ANTENNA_3982 (.A(net1192));
 sg13g2_antennanp ANTENNA_3983 (.A(net1192));
 sg13g2_antennanp ANTENNA_3984 (.A(net1192));
 sg13g2_antennanp ANTENNA_3985 (.A(net1192));
 sg13g2_antennanp ANTENNA_3986 (.A(net1273));
 sg13g2_antennanp ANTENNA_3987 (.A(net1273));
 sg13g2_antennanp ANTENNA_3988 (.A(net1273));
 sg13g2_antennanp ANTENNA_3989 (.A(net1273));
 sg13g2_antennanp ANTENNA_3990 (.A(net1273));
 sg13g2_antennanp ANTENNA_3991 (.A(net1273));
 sg13g2_antennanp ANTENNA_3992 (.A(net1273));
 sg13g2_antennanp ANTENNA_3993 (.A(net1273));
 sg13g2_antennanp ANTENNA_3994 (.A(net1273));
 sg13g2_antennanp ANTENNA_3995 (.A(_02490_));
 sg13g2_antennanp ANTENNA_3996 (.A(_03341_));
 sg13g2_antennanp ANTENNA_3997 (.A(_03444_));
 sg13g2_antennanp ANTENNA_3998 (.A(_03444_));
 sg13g2_antennanp ANTENNA_3999 (.A(_03444_));
 sg13g2_antennanp ANTENNA_4000 (.A(_03444_));
 sg13g2_antennanp ANTENNA_4001 (.A(_03621_));
 sg13g2_antennanp ANTENNA_4002 (.A(_03621_));
 sg13g2_antennanp ANTENNA_4003 (.A(_03621_));
 sg13g2_antennanp ANTENNA_4004 (.A(_03621_));
 sg13g2_antennanp ANTENNA_4005 (.A(_03621_));
 sg13g2_antennanp ANTENNA_4006 (.A(_03621_));
 sg13g2_antennanp ANTENNA_4007 (.A(_03621_));
 sg13g2_antennanp ANTENNA_4008 (.A(_03621_));
 sg13g2_antennanp ANTENNA_4009 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4010 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4011 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4012 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4013 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4014 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4015 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4016 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4017 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4018 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4019 (.A(_03850_));
 sg13g2_antennanp ANTENNA_4020 (.A(_03875_));
 sg13g2_antennanp ANTENNA_4021 (.A(_03995_));
 sg13g2_antennanp ANTENNA_4022 (.A(_03995_));
 sg13g2_antennanp ANTENNA_4023 (.A(_03995_));
 sg13g2_antennanp ANTENNA_4024 (.A(_03995_));
 sg13g2_antennanp ANTENNA_4025 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4026 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4027 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4028 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4029 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4030 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4031 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4032 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4033 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4034 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4035 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4036 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4037 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4038 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4039 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4040 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4041 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4042 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4043 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4044 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4045 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4046 (.A(_04431_));
 sg13g2_antennanp ANTENNA_4047 (.A(_05435_));
 sg13g2_antennanp ANTENNA_4048 (.A(_05441_));
 sg13g2_antennanp ANTENNA_4049 (.A(_05441_));
 sg13g2_antennanp ANTENNA_4050 (.A(_05441_));
 sg13g2_antennanp ANTENNA_4051 (.A(_05449_));
 sg13g2_antennanp ANTENNA_4052 (.A(_05449_));
 sg13g2_antennanp ANTENNA_4053 (.A(_05449_));
 sg13g2_antennanp ANTENNA_4054 (.A(_05449_));
 sg13g2_antennanp ANTENNA_4055 (.A(_05449_));
 sg13g2_antennanp ANTENNA_4056 (.A(_05449_));
 sg13g2_antennanp ANTENNA_4057 (.A(_05453_));
 sg13g2_antennanp ANTENNA_4058 (.A(_05453_));
 sg13g2_antennanp ANTENNA_4059 (.A(_05453_));
 sg13g2_antennanp ANTENNA_4060 (.A(_05453_));
 sg13g2_antennanp ANTENNA_4061 (.A(_05453_));
 sg13g2_antennanp ANTENNA_4062 (.A(_05453_));
 sg13g2_antennanp ANTENNA_4063 (.A(_05453_));
 sg13g2_antennanp ANTENNA_4064 (.A(_05453_));
 sg13g2_antennanp ANTENNA_4065 (.A(_05453_));
 sg13g2_antennanp ANTENNA_4066 (.A(_05457_));
 sg13g2_antennanp ANTENNA_4067 (.A(_05457_));
 sg13g2_antennanp ANTENNA_4068 (.A(_05457_));
 sg13g2_antennanp ANTENNA_4069 (.A(_05457_));
 sg13g2_antennanp ANTENNA_4070 (.A(_05457_));
 sg13g2_antennanp ANTENNA_4071 (.A(_05457_));
 sg13g2_antennanp ANTENNA_4072 (.A(_05463_));
 sg13g2_antennanp ANTENNA_4073 (.A(_05463_));
 sg13g2_antennanp ANTENNA_4074 (.A(_05463_));
 sg13g2_antennanp ANTENNA_4075 (.A(_05463_));
 sg13g2_antennanp ANTENNA_4076 (.A(_05463_));
 sg13g2_antennanp ANTENNA_4077 (.A(_05463_));
 sg13g2_antennanp ANTENNA_4078 (.A(_05467_));
 sg13g2_antennanp ANTENNA_4079 (.A(_05467_));
 sg13g2_antennanp ANTENNA_4080 (.A(_05467_));
 sg13g2_antennanp ANTENNA_4081 (.A(_05467_));
 sg13g2_antennanp ANTENNA_4082 (.A(_05467_));
 sg13g2_antennanp ANTENNA_4083 (.A(_05467_));
 sg13g2_antennanp ANTENNA_4084 (.A(_05471_));
 sg13g2_antennanp ANTENNA_4085 (.A(_05471_));
 sg13g2_antennanp ANTENNA_4086 (.A(_05471_));
 sg13g2_antennanp ANTENNA_4087 (.A(_05471_));
 sg13g2_antennanp ANTENNA_4088 (.A(_05471_));
 sg13g2_antennanp ANTENNA_4089 (.A(_05471_));
 sg13g2_antennanp ANTENNA_4090 (.A(_05471_));
 sg13g2_antennanp ANTENNA_4091 (.A(_05471_));
 sg13g2_antennanp ANTENNA_4092 (.A(_05471_));
 sg13g2_antennanp ANTENNA_4093 (.A(_05476_));
 sg13g2_antennanp ANTENNA_4094 (.A(_05476_));
 sg13g2_antennanp ANTENNA_4095 (.A(_05498_));
 sg13g2_antennanp ANTENNA_4096 (.A(_05498_));
 sg13g2_antennanp ANTENNA_4097 (.A(_06148_));
 sg13g2_antennanp ANTENNA_4098 (.A(_06148_));
 sg13g2_antennanp ANTENNA_4099 (.A(_06148_));
 sg13g2_antennanp ANTENNA_4100 (.A(_06148_));
 sg13g2_antennanp ANTENNA_4101 (.A(_06148_));
 sg13g2_antennanp ANTENNA_4102 (.A(_06171_));
 sg13g2_antennanp ANTENNA_4103 (.A(_06189_));
 sg13g2_antennanp ANTENNA_4104 (.A(_06253_));
 sg13g2_antennanp ANTENNA_4105 (.A(_06255_));
 sg13g2_antennanp ANTENNA_4106 (.A(_06268_));
 sg13g2_antennanp ANTENNA_4107 (.A(_06293_));
 sg13g2_antennanp ANTENNA_4108 (.A(_06293_));
 sg13g2_antennanp ANTENNA_4109 (.A(_06298_));
 sg13g2_antennanp ANTENNA_4110 (.A(_06298_));
 sg13g2_antennanp ANTENNA_4111 (.A(_06311_));
 sg13g2_antennanp ANTENNA_4112 (.A(_06318_));
 sg13g2_antennanp ANTENNA_4113 (.A(_06329_));
 sg13g2_antennanp ANTENNA_4114 (.A(_06416_));
 sg13g2_antennanp ANTENNA_4115 (.A(_06416_));
 sg13g2_antennanp ANTENNA_4116 (.A(_06493_));
 sg13g2_antennanp ANTENNA_4117 (.A(_06493_));
 sg13g2_antennanp ANTENNA_4118 (.A(_06520_));
 sg13g2_antennanp ANTENNA_4119 (.A(_06559_));
 sg13g2_antennanp ANTENNA_4120 (.A(_06560_));
 sg13g2_antennanp ANTENNA_4121 (.A(_06595_));
 sg13g2_antennanp ANTENNA_4122 (.A(_06601_));
 sg13g2_antennanp ANTENNA_4123 (.A(_06616_));
 sg13g2_antennanp ANTENNA_4124 (.A(_06620_));
 sg13g2_antennanp ANTENNA_4125 (.A(_06700_));
 sg13g2_antennanp ANTENNA_4126 (.A(_06719_));
 sg13g2_antennanp ANTENNA_4127 (.A(_06757_));
 sg13g2_antennanp ANTENNA_4128 (.A(_06772_));
 sg13g2_antennanp ANTENNA_4129 (.A(_06772_));
 sg13g2_antennanp ANTENNA_4130 (.A(_06793_));
 sg13g2_antennanp ANTENNA_4131 (.A(_06799_));
 sg13g2_antennanp ANTENNA_4132 (.A(_06799_));
 sg13g2_antennanp ANTENNA_4133 (.A(_06814_));
 sg13g2_antennanp ANTENNA_4134 (.A(_06818_));
 sg13g2_antennanp ANTENNA_4135 (.A(_06856_));
 sg13g2_antennanp ANTENNA_4136 (.A(_06871_));
 sg13g2_antennanp ANTENNA_4137 (.A(_06871_));
 sg13g2_antennanp ANTENNA_4138 (.A(_06913_));
 sg13g2_antennanp ANTENNA_4139 (.A(_06917_));
 sg13g2_antennanp ANTENNA_4140 (.A(_06955_));
 sg13g2_antennanp ANTENNA_4141 (.A(_06955_));
 sg13g2_antennanp ANTENNA_4142 (.A(_06975_));
 sg13g2_antennanp ANTENNA_4143 (.A(_07012_));
 sg13g2_antennanp ANTENNA_4144 (.A(_07012_));
 sg13g2_antennanp ANTENNA_4145 (.A(_07016_));
 sg13g2_antennanp ANTENNA_4146 (.A(_07054_));
 sg13g2_antennanp ANTENNA_4147 (.A(_07074_));
 sg13g2_antennanp ANTENNA_4148 (.A(_07074_));
 sg13g2_antennanp ANTENNA_4149 (.A(_07090_));
 sg13g2_antennanp ANTENNA_4150 (.A(_07105_));
 sg13g2_antennanp ANTENNA_4151 (.A(_07105_));
 sg13g2_antennanp ANTENNA_4152 (.A(_07105_));
 sg13g2_antennanp ANTENNA_4153 (.A(_07335_));
 sg13g2_antennanp ANTENNA_4154 (.A(_07416_));
 sg13g2_antennanp ANTENNA_4155 (.A(_07416_));
 sg13g2_antennanp ANTENNA_4156 (.A(_07416_));
 sg13g2_antennanp ANTENNA_4157 (.A(_07416_));
 sg13g2_antennanp ANTENNA_4158 (.A(_07416_));
 sg13g2_antennanp ANTENNA_4159 (.A(_07416_));
 sg13g2_antennanp ANTENNA_4160 (.A(_09194_));
 sg13g2_antennanp ANTENNA_4161 (.A(_09194_));
 sg13g2_antennanp ANTENNA_4162 (.A(_09194_));
 sg13g2_antennanp ANTENNA_4163 (.A(_09194_));
 sg13g2_antennanp ANTENNA_4164 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4165 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4166 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4167 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4168 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4169 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4170 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4171 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4172 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4173 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4174 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4175 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4176 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4177 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4178 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4179 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4180 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4181 (.A(_09260_));
 sg13g2_antennanp ANTENNA_4182 (.A(_09345_));
 sg13g2_antennanp ANTENNA_4183 (.A(_09345_));
 sg13g2_antennanp ANTENNA_4184 (.A(_09345_));
 sg13g2_antennanp ANTENNA_4185 (.A(_09345_));
 sg13g2_antennanp ANTENNA_4186 (.A(_09345_));
 sg13g2_antennanp ANTENNA_4187 (.A(_09345_));
 sg13g2_antennanp ANTENNA_4188 (.A(_09345_));
 sg13g2_antennanp ANTENNA_4189 (.A(_09345_));
 sg13g2_antennanp ANTENNA_4190 (.A(_09345_));
 sg13g2_antennanp ANTENNA_4191 (.A(_09418_));
 sg13g2_antennanp ANTENNA_4192 (.A(_09418_));
 sg13g2_antennanp ANTENNA_4193 (.A(_09418_));
 sg13g2_antennanp ANTENNA_4194 (.A(_09418_));
 sg13g2_antennanp ANTENNA_4195 (.A(_09418_));
 sg13g2_antennanp ANTENNA_4196 (.A(_09418_));
 sg13g2_antennanp ANTENNA_4197 (.A(_09418_));
 sg13g2_antennanp ANTENNA_4198 (.A(_09418_));
 sg13g2_antennanp ANTENNA_4199 (.A(_09418_));
 sg13g2_antennanp ANTENNA_4200 (.A(_09906_));
 sg13g2_antennanp ANTENNA_4201 (.A(_09906_));
 sg13g2_antennanp ANTENNA_4202 (.A(_09906_));
 sg13g2_antennanp ANTENNA_4203 (.A(_09906_));
 sg13g2_antennanp ANTENNA_4204 (.A(_09906_));
 sg13g2_antennanp ANTENNA_4205 (.A(_09906_));
 sg13g2_antennanp ANTENNA_4206 (.A(_09906_));
 sg13g2_antennanp ANTENNA_4207 (.A(_09906_));
 sg13g2_antennanp ANTENNA_4208 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4209 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4210 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4211 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4212 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4213 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4214 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4215 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4216 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4217 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4218 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4219 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4220 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4221 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4222 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4223 (.A(_09928_));
 sg13g2_antennanp ANTENNA_4224 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4225 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4226 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4227 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4228 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4229 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4230 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4231 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4232 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4233 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4234 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4235 (.A(_09929_));
 sg13g2_antennanp ANTENNA_4236 (.A(_09930_));
 sg13g2_antennanp ANTENNA_4237 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4238 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4239 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4240 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4241 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4242 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4243 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4244 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4245 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4246 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4247 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4248 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4249 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4250 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4251 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4252 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4253 (.A(_09935_));
 sg13g2_antennanp ANTENNA_4254 (.A(_10040_));
 sg13g2_antennanp ANTENNA_4255 (.A(_10040_));
 sg13g2_antennanp ANTENNA_4256 (.A(_10040_));
 sg13g2_antennanp ANTENNA_4257 (.A(_10040_));
 sg13g2_antennanp ANTENNA_4258 (.A(_10040_));
 sg13g2_antennanp ANTENNA_4259 (.A(_10040_));
 sg13g2_antennanp ANTENNA_4260 (.A(_10040_));
 sg13g2_antennanp ANTENNA_4261 (.A(_10040_));
 sg13g2_antennanp ANTENNA_4262 (.A(_10040_));
 sg13g2_antennanp ANTENNA_4263 (.A(_10042_));
 sg13g2_antennanp ANTENNA_4264 (.A(_10042_));
 sg13g2_antennanp ANTENNA_4265 (.A(_10042_));
 sg13g2_antennanp ANTENNA_4266 (.A(_10042_));
 sg13g2_antennanp ANTENNA_4267 (.A(_10046_));
 sg13g2_antennanp ANTENNA_4268 (.A(_10048_));
 sg13g2_antennanp ANTENNA_4269 (.A(_10051_));
 sg13g2_antennanp ANTENNA_4270 (.A(_10053_));
 sg13g2_antennanp ANTENNA_4271 (.A(_10071_));
 sg13g2_antennanp ANTENNA_4272 (.A(_10071_));
 sg13g2_antennanp ANTENNA_4273 (.A(_10071_));
 sg13g2_antennanp ANTENNA_4274 (.A(_10071_));
 sg13g2_antennanp ANTENNA_4275 (.A(_10071_));
 sg13g2_antennanp ANTENNA_4276 (.A(_10071_));
 sg13g2_antennanp ANTENNA_4277 (.A(_10083_));
 sg13g2_antennanp ANTENNA_4278 (.A(_10091_));
 sg13g2_antennanp ANTENNA_4279 (.A(_10092_));
 sg13g2_antennanp ANTENNA_4280 (.A(_10092_));
 sg13g2_antennanp ANTENNA_4281 (.A(_10092_));
 sg13g2_antennanp ANTENNA_4282 (.A(_10101_));
 sg13g2_antennanp ANTENNA_4283 (.A(_10106_));
 sg13g2_antennanp ANTENNA_4284 (.A(_10110_));
 sg13g2_antennanp ANTENNA_4285 (.A(_10121_));
 sg13g2_antennanp ANTENNA_4286 (.A(_10121_));
 sg13g2_antennanp ANTENNA_4287 (.A(_10131_));
 sg13g2_antennanp ANTENNA_4288 (.A(_10131_));
 sg13g2_antennanp ANTENNA_4289 (.A(_10136_));
 sg13g2_antennanp ANTENNA_4290 (.A(_10140_));
 sg13g2_antennanp ANTENNA_4291 (.A(_10140_));
 sg13g2_antennanp ANTENNA_4292 (.A(_10226_));
 sg13g2_antennanp ANTENNA_4293 (.A(_10226_));
 sg13g2_antennanp ANTENNA_4294 (.A(_10226_));
 sg13g2_antennanp ANTENNA_4295 (.A(_10226_));
 sg13g2_antennanp ANTENNA_4296 (.A(_10226_));
 sg13g2_antennanp ANTENNA_4297 (.A(_10226_));
 sg13g2_antennanp ANTENNA_4298 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4299 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4300 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4301 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4302 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4303 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4304 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4305 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4306 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4307 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4308 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4309 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4310 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4311 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4312 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4313 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4314 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4315 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4316 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4317 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4318 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4319 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4320 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4321 (.A(_10232_));
 sg13g2_antennanp ANTENNA_4322 (.A(_10236_));
 sg13g2_antennanp ANTENNA_4323 (.A(_10236_));
 sg13g2_antennanp ANTENNA_4324 (.A(_10236_));
 sg13g2_antennanp ANTENNA_4325 (.A(_10236_));
 sg13g2_antennanp ANTENNA_4326 (.A(_10236_));
 sg13g2_antennanp ANTENNA_4327 (.A(_10236_));
 sg13g2_antennanp ANTENNA_4328 (.A(_10236_));
 sg13g2_antennanp ANTENNA_4329 (.A(_10243_));
 sg13g2_antennanp ANTENNA_4330 (.A(_10243_));
 sg13g2_antennanp ANTENNA_4331 (.A(_10243_));
 sg13g2_antennanp ANTENNA_4332 (.A(_10243_));
 sg13g2_antennanp ANTENNA_4333 (.A(_10243_));
 sg13g2_antennanp ANTENNA_4334 (.A(_10243_));
 sg13g2_antennanp ANTENNA_4335 (.A(_10256_));
 sg13g2_antennanp ANTENNA_4336 (.A(_10256_));
 sg13g2_antennanp ANTENNA_4337 (.A(_10256_));
 sg13g2_antennanp ANTENNA_4338 (.A(_10256_));
 sg13g2_antennanp ANTENNA_4339 (.A(_10256_));
 sg13g2_antennanp ANTENNA_4340 (.A(_10287_));
 sg13g2_antennanp ANTENNA_4341 (.A(_10287_));
 sg13g2_antennanp ANTENNA_4342 (.A(_10287_));
 sg13g2_antennanp ANTENNA_4343 (.A(_10287_));
 sg13g2_antennanp ANTENNA_4344 (.A(_10287_));
 sg13g2_antennanp ANTENNA_4345 (.A(_10295_));
 sg13g2_antennanp ANTENNA_4346 (.A(_10295_));
 sg13g2_antennanp ANTENNA_4347 (.A(_10295_));
 sg13g2_antennanp ANTENNA_4348 (.A(_10295_));
 sg13g2_antennanp ANTENNA_4349 (.A(_10295_));
 sg13g2_antennanp ANTENNA_4350 (.A(_10295_));
 sg13g2_antennanp ANTENNA_4351 (.A(_10295_));
 sg13g2_antennanp ANTENNA_4352 (.A(_10295_));
 sg13g2_antennanp ANTENNA_4353 (.A(_10349_));
 sg13g2_antennanp ANTENNA_4354 (.A(_10349_));
 sg13g2_antennanp ANTENNA_4355 (.A(_10349_));
 sg13g2_antennanp ANTENNA_4356 (.A(_10349_));
 sg13g2_antennanp ANTENNA_4357 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4358 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4359 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4360 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4361 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4362 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4363 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4364 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4365 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4366 (.A(_10350_));
 sg13g2_antennanp ANTENNA_4367 (.A(_10397_));
 sg13g2_antennanp ANTENNA_4368 (.A(_10397_));
 sg13g2_antennanp ANTENNA_4369 (.A(_10397_));
 sg13g2_antennanp ANTENNA_4370 (.A(_10397_));
 sg13g2_antennanp ANTENNA_4371 (.A(_10397_));
 sg13g2_antennanp ANTENNA_4372 (.A(_10397_));
 sg13g2_antennanp ANTENNA_4373 (.A(_10397_));
 sg13g2_antennanp ANTENNA_4374 (.A(_10397_));
 sg13g2_antennanp ANTENNA_4375 (.A(_10422_));
 sg13g2_antennanp ANTENNA_4376 (.A(_10422_));
 sg13g2_antennanp ANTENNA_4377 (.A(_10422_));
 sg13g2_antennanp ANTENNA_4378 (.A(_10422_));
 sg13g2_antennanp ANTENNA_4379 (.A(_10422_));
 sg13g2_antennanp ANTENNA_4380 (.A(_10422_));
 sg13g2_antennanp ANTENNA_4381 (.A(_10422_));
 sg13g2_antennanp ANTENNA_4382 (.A(_10422_));
 sg13g2_antennanp ANTENNA_4383 (.A(_10422_));
 sg13g2_antennanp ANTENNA_4384 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4385 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4386 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4387 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4388 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4389 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4390 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4391 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4392 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4393 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4394 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4395 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4396 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4397 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4398 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4399 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4400 (.A(_10444_));
 sg13g2_antennanp ANTENNA_4401 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4402 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4403 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4404 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4405 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4406 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4407 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4408 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4409 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4410 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4411 (.A(_10491_));
 sg13g2_antennanp ANTENNA_4412 (.A(_10492_));
 sg13g2_antennanp ANTENNA_4413 (.A(_10492_));
 sg13g2_antennanp ANTENNA_4414 (.A(_10492_));
 sg13g2_antennanp ANTENNA_4415 (.A(_10492_));
 sg13g2_antennanp ANTENNA_4416 (.A(_10492_));
 sg13g2_antennanp ANTENNA_4417 (.A(_10492_));
 sg13g2_antennanp ANTENNA_4418 (.A(_10492_));
 sg13g2_antennanp ANTENNA_4419 (.A(_10492_));
 sg13g2_antennanp ANTENNA_4420 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4421 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4422 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4423 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4424 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4425 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4426 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4427 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4428 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4429 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4430 (.A(_10513_));
 sg13g2_antennanp ANTENNA_4431 (.A(_10514_));
 sg13g2_antennanp ANTENNA_4432 (.A(_10514_));
 sg13g2_antennanp ANTENNA_4433 (.A(_10514_));
 sg13g2_antennanp ANTENNA_4434 (.A(_10514_));
 sg13g2_antennanp ANTENNA_4435 (.A(_10514_));
 sg13g2_antennanp ANTENNA_4436 (.A(_10514_));
 sg13g2_antennanp ANTENNA_4437 (.A(_10564_));
 sg13g2_antennanp ANTENNA_4438 (.A(_10564_));
 sg13g2_antennanp ANTENNA_4439 (.A(_10564_));
 sg13g2_antennanp ANTENNA_4440 (.A(_10564_));
 sg13g2_antennanp ANTENNA_4441 (.A(_10564_));
 sg13g2_antennanp ANTENNA_4442 (.A(_10564_));
 sg13g2_antennanp ANTENNA_4443 (.A(_10564_));
 sg13g2_antennanp ANTENNA_4444 (.A(_10586_));
 sg13g2_antennanp ANTENNA_4445 (.A(_10586_));
 sg13g2_antennanp ANTENNA_4446 (.A(_10586_));
 sg13g2_antennanp ANTENNA_4447 (.A(_10586_));
 sg13g2_antennanp ANTENNA_4448 (.A(_10586_));
 sg13g2_antennanp ANTENNA_4449 (.A(_10586_));
 sg13g2_antennanp ANTENNA_4450 (.A(_10586_));
 sg13g2_antennanp ANTENNA_4451 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4452 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4453 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4454 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4455 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4456 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4457 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4458 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4459 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4460 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4461 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4462 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4463 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4464 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4465 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4466 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4467 (.A(_10632_));
 sg13g2_antennanp ANTENNA_4468 (.A(_10656_));
 sg13g2_antennanp ANTENNA_4469 (.A(_10656_));
 sg13g2_antennanp ANTENNA_4470 (.A(_10656_));
 sg13g2_antennanp ANTENNA_4471 (.A(_10656_));
 sg13g2_antennanp ANTENNA_4472 (.A(_10656_));
 sg13g2_antennanp ANTENNA_4473 (.A(_10656_));
 sg13g2_antennanp ANTENNA_4474 (.A(_10656_));
 sg13g2_antennanp ANTENNA_4475 (.A(_10656_));
 sg13g2_antennanp ANTENNA_4476 (.A(_10657_));
 sg13g2_antennanp ANTENNA_4477 (.A(_10657_));
 sg13g2_antennanp ANTENNA_4478 (.A(_10657_));
 sg13g2_antennanp ANTENNA_4479 (.A(_10657_));
 sg13g2_antennanp ANTENNA_4480 (.A(_10657_));
 sg13g2_antennanp ANTENNA_4481 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4482 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4483 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4484 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4485 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4486 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4487 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4488 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4489 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4490 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4491 (.A(_10679_));
 sg13g2_antennanp ANTENNA_4492 (.A(_11171_));
 sg13g2_antennanp ANTENNA_4493 (.A(_11171_));
 sg13g2_antennanp ANTENNA_4494 (.A(_11171_));
 sg13g2_antennanp ANTENNA_4495 (.A(_11171_));
 sg13g2_antennanp ANTENNA_4496 (.A(_11171_));
 sg13g2_antennanp ANTENNA_4497 (.A(_11171_));
 sg13g2_antennanp ANTENNA_4498 (.A(_11171_));
 sg13g2_antennanp ANTENNA_4499 (.A(_11947_));
 sg13g2_antennanp ANTENNA_4500 (.A(_11947_));
 sg13g2_antennanp ANTENNA_4501 (.A(_11947_));
 sg13g2_antennanp ANTENNA_4502 (.A(_11947_));
 sg13g2_antennanp ANTENNA_4503 (.A(_12437_));
 sg13g2_antennanp ANTENNA_4504 (.A(_12437_));
 sg13g2_antennanp ANTENNA_4505 (.A(_12437_));
 sg13g2_antennanp ANTENNA_4506 (.A(_12653_));
 sg13g2_antennanp ANTENNA_4507 (.A(_12653_));
 sg13g2_antennanp ANTENNA_4508 (.A(_12653_));
 sg13g2_antennanp ANTENNA_4509 (.A(_12653_));
 sg13g2_antennanp ANTENNA_4510 (.A(_12653_));
 sg13g2_antennanp ANTENNA_4511 (.A(_12653_));
 sg13g2_antennanp ANTENNA_4512 (.A(_12653_));
 sg13g2_antennanp ANTENNA_4513 (.A(_12658_));
 sg13g2_antennanp ANTENNA_4514 (.A(_12658_));
 sg13g2_antennanp ANTENNA_4515 (.A(_12658_));
 sg13g2_antennanp ANTENNA_4516 (.A(_12658_));
 sg13g2_antennanp ANTENNA_4517 (.A(clk));
 sg13g2_antennanp ANTENNA_4518 (.A(clk));
 sg13g2_antennanp ANTENNA_4519 (.A(\mem.io_data_out[3] ));
 sg13g2_antennanp ANTENNA_4520 (.A(\mem.io_data_out[3] ));
 sg13g2_antennanp ANTENNA_4521 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_4522 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_4523 (.A(\mem.mem_internal.code_mem[24][4] ));
 sg13g2_antennanp ANTENNA_4524 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_4525 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_4526 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_4527 (.A(ui_in[5]));
 sg13g2_antennanp ANTENNA_4528 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_4529 (.A(ui_in[6]));
 sg13g2_antennanp ANTENNA_4530 (.A(net1));
 sg13g2_antennanp ANTENNA_4531 (.A(net1));
 sg13g2_antennanp ANTENNA_4532 (.A(net1));
 sg13g2_antennanp ANTENNA_4533 (.A(net464));
 sg13g2_antennanp ANTENNA_4534 (.A(net464));
 sg13g2_antennanp ANTENNA_4535 (.A(net464));
 sg13g2_antennanp ANTENNA_4536 (.A(net464));
 sg13g2_antennanp ANTENNA_4537 (.A(net464));
 sg13g2_antennanp ANTENNA_4538 (.A(net464));
 sg13g2_antennanp ANTENNA_4539 (.A(net464));
 sg13g2_antennanp ANTENNA_4540 (.A(net464));
 sg13g2_antennanp ANTENNA_4541 (.A(net464));
 sg13g2_antennanp ANTENNA_4542 (.A(net526));
 sg13g2_antennanp ANTENNA_4543 (.A(net526));
 sg13g2_antennanp ANTENNA_4544 (.A(net526));
 sg13g2_antennanp ANTENNA_4545 (.A(net526));
 sg13g2_antennanp ANTENNA_4546 (.A(net526));
 sg13g2_antennanp ANTENNA_4547 (.A(net526));
 sg13g2_antennanp ANTENNA_4548 (.A(net526));
 sg13g2_antennanp ANTENNA_4549 (.A(net526));
 sg13g2_antennanp ANTENNA_4550 (.A(net526));
 sg13g2_antennanp ANTENNA_4551 (.A(net526));
 sg13g2_antennanp ANTENNA_4552 (.A(net526));
 sg13g2_antennanp ANTENNA_4553 (.A(net526));
 sg13g2_antennanp ANTENNA_4554 (.A(net526));
 sg13g2_antennanp ANTENNA_4555 (.A(net526));
 sg13g2_antennanp ANTENNA_4556 (.A(net526));
 sg13g2_antennanp ANTENNA_4557 (.A(net526));
 sg13g2_antennanp ANTENNA_4558 (.A(net526));
 sg13g2_antennanp ANTENNA_4559 (.A(net526));
 sg13g2_antennanp ANTENNA_4560 (.A(net526));
 sg13g2_antennanp ANTENNA_4561 (.A(net526));
 sg13g2_antennanp ANTENNA_4562 (.A(net526));
 sg13g2_antennanp ANTENNA_4563 (.A(net526));
 sg13g2_antennanp ANTENNA_4564 (.A(net526));
 sg13g2_antennanp ANTENNA_4565 (.A(net527));
 sg13g2_antennanp ANTENNA_4566 (.A(net527));
 sg13g2_antennanp ANTENNA_4567 (.A(net527));
 sg13g2_antennanp ANTENNA_4568 (.A(net527));
 sg13g2_antennanp ANTENNA_4569 (.A(net527));
 sg13g2_antennanp ANTENNA_4570 (.A(net527));
 sg13g2_antennanp ANTENNA_4571 (.A(net527));
 sg13g2_antennanp ANTENNA_4572 (.A(net527));
 sg13g2_antennanp ANTENNA_4573 (.A(net527));
 sg13g2_antennanp ANTENNA_4574 (.A(net527));
 sg13g2_antennanp ANTENNA_4575 (.A(net527));
 sg13g2_antennanp ANTENNA_4576 (.A(net527));
 sg13g2_antennanp ANTENNA_4577 (.A(net527));
 sg13g2_antennanp ANTENNA_4578 (.A(net527));
 sg13g2_antennanp ANTENNA_4579 (.A(net529));
 sg13g2_antennanp ANTENNA_4580 (.A(net529));
 sg13g2_antennanp ANTENNA_4581 (.A(net529));
 sg13g2_antennanp ANTENNA_4582 (.A(net529));
 sg13g2_antennanp ANTENNA_4583 (.A(net529));
 sg13g2_antennanp ANTENNA_4584 (.A(net529));
 sg13g2_antennanp ANTENNA_4585 (.A(net529));
 sg13g2_antennanp ANTENNA_4586 (.A(net529));
 sg13g2_antennanp ANTENNA_4587 (.A(net529));
 sg13g2_antennanp ANTENNA_4588 (.A(net529));
 sg13g2_antennanp ANTENNA_4589 (.A(net529));
 sg13g2_antennanp ANTENNA_4590 (.A(net529));
 sg13g2_antennanp ANTENNA_4591 (.A(net529));
 sg13g2_antennanp ANTENNA_4592 (.A(net529));
 sg13g2_antennanp ANTENNA_4593 (.A(net529));
 sg13g2_antennanp ANTENNA_4594 (.A(net549));
 sg13g2_antennanp ANTENNA_4595 (.A(net549));
 sg13g2_antennanp ANTENNA_4596 (.A(net549));
 sg13g2_antennanp ANTENNA_4597 (.A(net549));
 sg13g2_antennanp ANTENNA_4598 (.A(net549));
 sg13g2_antennanp ANTENNA_4599 (.A(net549));
 sg13g2_antennanp ANTENNA_4600 (.A(net549));
 sg13g2_antennanp ANTENNA_4601 (.A(net549));
 sg13g2_antennanp ANTENNA_4602 (.A(net553));
 sg13g2_antennanp ANTENNA_4603 (.A(net553));
 sg13g2_antennanp ANTENNA_4604 (.A(net553));
 sg13g2_antennanp ANTENNA_4605 (.A(net553));
 sg13g2_antennanp ANTENNA_4606 (.A(net553));
 sg13g2_antennanp ANTENNA_4607 (.A(net553));
 sg13g2_antennanp ANTENNA_4608 (.A(net553));
 sg13g2_antennanp ANTENNA_4609 (.A(net553));
 sg13g2_antennanp ANTENNA_4610 (.A(net553));
 sg13g2_antennanp ANTENNA_4611 (.A(net553));
 sg13g2_antennanp ANTENNA_4612 (.A(net553));
 sg13g2_antennanp ANTENNA_4613 (.A(net553));
 sg13g2_antennanp ANTENNA_4614 (.A(net553));
 sg13g2_antennanp ANTENNA_4615 (.A(net553));
 sg13g2_antennanp ANTENNA_4616 (.A(net553));
 sg13g2_antennanp ANTENNA_4617 (.A(net553));
 sg13g2_antennanp ANTENNA_4618 (.A(net553));
 sg13g2_antennanp ANTENNA_4619 (.A(net554));
 sg13g2_antennanp ANTENNA_4620 (.A(net554));
 sg13g2_antennanp ANTENNA_4621 (.A(net554));
 sg13g2_antennanp ANTENNA_4622 (.A(net554));
 sg13g2_antennanp ANTENNA_4623 (.A(net554));
 sg13g2_antennanp ANTENNA_4624 (.A(net554));
 sg13g2_antennanp ANTENNA_4625 (.A(net554));
 sg13g2_antennanp ANTENNA_4626 (.A(net554));
 sg13g2_antennanp ANTENNA_4627 (.A(net554));
 sg13g2_antennanp ANTENNA_4628 (.A(net554));
 sg13g2_antennanp ANTENNA_4629 (.A(net554));
 sg13g2_antennanp ANTENNA_4630 (.A(net554));
 sg13g2_antennanp ANTENNA_4631 (.A(net554));
 sg13g2_antennanp ANTENNA_4632 (.A(net554));
 sg13g2_antennanp ANTENNA_4633 (.A(net554));
 sg13g2_antennanp ANTENNA_4634 (.A(net554));
 sg13g2_antennanp ANTENNA_4635 (.A(net554));
 sg13g2_antennanp ANTENNA_4636 (.A(net554));
 sg13g2_antennanp ANTENNA_4637 (.A(net554));
 sg13g2_antennanp ANTENNA_4638 (.A(net554));
 sg13g2_antennanp ANTENNA_4639 (.A(net554));
 sg13g2_antennanp ANTENNA_4640 (.A(net554));
 sg13g2_antennanp ANTENNA_4641 (.A(net554));
 sg13g2_antennanp ANTENNA_4642 (.A(net556));
 sg13g2_antennanp ANTENNA_4643 (.A(net556));
 sg13g2_antennanp ANTENNA_4644 (.A(net556));
 sg13g2_antennanp ANTENNA_4645 (.A(net556));
 sg13g2_antennanp ANTENNA_4646 (.A(net556));
 sg13g2_antennanp ANTENNA_4647 (.A(net556));
 sg13g2_antennanp ANTENNA_4648 (.A(net556));
 sg13g2_antennanp ANTENNA_4649 (.A(net556));
 sg13g2_antennanp ANTENNA_4650 (.A(net556));
 sg13g2_antennanp ANTENNA_4651 (.A(net641));
 sg13g2_antennanp ANTENNA_4652 (.A(net641));
 sg13g2_antennanp ANTENNA_4653 (.A(net641));
 sg13g2_antennanp ANTENNA_4654 (.A(net641));
 sg13g2_antennanp ANTENNA_4655 (.A(net641));
 sg13g2_antennanp ANTENNA_4656 (.A(net641));
 sg13g2_antennanp ANTENNA_4657 (.A(net641));
 sg13g2_antennanp ANTENNA_4658 (.A(net641));
 sg13g2_antennanp ANTENNA_4659 (.A(net641));
 sg13g2_antennanp ANTENNA_4660 (.A(net770));
 sg13g2_antennanp ANTENNA_4661 (.A(net770));
 sg13g2_antennanp ANTENNA_4662 (.A(net770));
 sg13g2_antennanp ANTENNA_4663 (.A(net770));
 sg13g2_antennanp ANTENNA_4664 (.A(net770));
 sg13g2_antennanp ANTENNA_4665 (.A(net770));
 sg13g2_antennanp ANTENNA_4666 (.A(net770));
 sg13g2_antennanp ANTENNA_4667 (.A(net770));
 sg13g2_antennanp ANTENNA_4668 (.A(net770));
 sg13g2_antennanp ANTENNA_4669 (.A(net770));
 sg13g2_antennanp ANTENNA_4670 (.A(net770));
 sg13g2_antennanp ANTENNA_4671 (.A(net770));
 sg13g2_antennanp ANTENNA_4672 (.A(net770));
 sg13g2_antennanp ANTENNA_4673 (.A(net770));
 sg13g2_antennanp ANTENNA_4674 (.A(net778));
 sg13g2_antennanp ANTENNA_4675 (.A(net778));
 sg13g2_antennanp ANTENNA_4676 (.A(net778));
 sg13g2_antennanp ANTENNA_4677 (.A(net778));
 sg13g2_antennanp ANTENNA_4678 (.A(net778));
 sg13g2_antennanp ANTENNA_4679 (.A(net778));
 sg13g2_antennanp ANTENNA_4680 (.A(net778));
 sg13g2_antennanp ANTENNA_4681 (.A(net778));
 sg13g2_antennanp ANTENNA_4682 (.A(net778));
 sg13g2_antennanp ANTENNA_4683 (.A(net779));
 sg13g2_antennanp ANTENNA_4684 (.A(net779));
 sg13g2_antennanp ANTENNA_4685 (.A(net779));
 sg13g2_antennanp ANTENNA_4686 (.A(net779));
 sg13g2_antennanp ANTENNA_4687 (.A(net779));
 sg13g2_antennanp ANTENNA_4688 (.A(net779));
 sg13g2_antennanp ANTENNA_4689 (.A(net779));
 sg13g2_antennanp ANTENNA_4690 (.A(net779));
 sg13g2_antennanp ANTENNA_4691 (.A(net779));
 sg13g2_antennanp ANTENNA_4692 (.A(net779));
 sg13g2_antennanp ANTENNA_4693 (.A(net779));
 sg13g2_antennanp ANTENNA_4694 (.A(net779));
 sg13g2_antennanp ANTENNA_4695 (.A(net779));
 sg13g2_antennanp ANTENNA_4696 (.A(net779));
 sg13g2_antennanp ANTENNA_4697 (.A(net792));
 sg13g2_antennanp ANTENNA_4698 (.A(net792));
 sg13g2_antennanp ANTENNA_4699 (.A(net792));
 sg13g2_antennanp ANTENNA_4700 (.A(net792));
 sg13g2_antennanp ANTENNA_4701 (.A(net792));
 sg13g2_antennanp ANTENNA_4702 (.A(net792));
 sg13g2_antennanp ANTENNA_4703 (.A(net792));
 sg13g2_antennanp ANTENNA_4704 (.A(net792));
 sg13g2_antennanp ANTENNA_4705 (.A(net802));
 sg13g2_antennanp ANTENNA_4706 (.A(net802));
 sg13g2_antennanp ANTENNA_4707 (.A(net802));
 sg13g2_antennanp ANTENNA_4708 (.A(net802));
 sg13g2_antennanp ANTENNA_4709 (.A(net802));
 sg13g2_antennanp ANTENNA_4710 (.A(net802));
 sg13g2_antennanp ANTENNA_4711 (.A(net802));
 sg13g2_antennanp ANTENNA_4712 (.A(net802));
 sg13g2_antennanp ANTENNA_4713 (.A(net802));
 sg13g2_antennanp ANTENNA_4714 (.A(net838));
 sg13g2_antennanp ANTENNA_4715 (.A(net838));
 sg13g2_antennanp ANTENNA_4716 (.A(net838));
 sg13g2_antennanp ANTENNA_4717 (.A(net838));
 sg13g2_antennanp ANTENNA_4718 (.A(net838));
 sg13g2_antennanp ANTENNA_4719 (.A(net838));
 sg13g2_antennanp ANTENNA_4720 (.A(net838));
 sg13g2_antennanp ANTENNA_4721 (.A(net838));
 sg13g2_antennanp ANTENNA_4722 (.A(net838));
 sg13g2_antennanp ANTENNA_4723 (.A(net878));
 sg13g2_antennanp ANTENNA_4724 (.A(net878));
 sg13g2_antennanp ANTENNA_4725 (.A(net878));
 sg13g2_antennanp ANTENNA_4726 (.A(net878));
 sg13g2_antennanp ANTENNA_4727 (.A(net878));
 sg13g2_antennanp ANTENNA_4728 (.A(net878));
 sg13g2_antennanp ANTENNA_4729 (.A(net878));
 sg13g2_antennanp ANTENNA_4730 (.A(net878));
 sg13g2_antennanp ANTENNA_4731 (.A(net878));
 sg13g2_antennanp ANTENNA_4732 (.A(net878));
 sg13g2_antennanp ANTENNA_4733 (.A(net878));
 sg13g2_antennanp ANTENNA_4734 (.A(net878));
 sg13g2_antennanp ANTENNA_4735 (.A(net878));
 sg13g2_antennanp ANTENNA_4736 (.A(net878));
 sg13g2_antennanp ANTENNA_4737 (.A(net878));
 sg13g2_antennanp ANTENNA_4738 (.A(net878));
 sg13g2_antennanp ANTENNA_4739 (.A(net878));
 sg13g2_antennanp ANTENNA_4740 (.A(net878));
 sg13g2_antennanp ANTENNA_4741 (.A(net878));
 sg13g2_antennanp ANTENNA_4742 (.A(net878));
 sg13g2_antennanp ANTENNA_4743 (.A(net924));
 sg13g2_antennanp ANTENNA_4744 (.A(net924));
 sg13g2_antennanp ANTENNA_4745 (.A(net924));
 sg13g2_antennanp ANTENNA_4746 (.A(net924));
 sg13g2_antennanp ANTENNA_4747 (.A(net924));
 sg13g2_antennanp ANTENNA_4748 (.A(net924));
 sg13g2_antennanp ANTENNA_4749 (.A(net924));
 sg13g2_antennanp ANTENNA_4750 (.A(net924));
 sg13g2_antennanp ANTENNA_4751 (.A(net924));
 sg13g2_antennanp ANTENNA_4752 (.A(net982));
 sg13g2_antennanp ANTENNA_4753 (.A(net982));
 sg13g2_antennanp ANTENNA_4754 (.A(net982));
 sg13g2_antennanp ANTENNA_4755 (.A(net982));
 sg13g2_antennanp ANTENNA_4756 (.A(net982));
 sg13g2_antennanp ANTENNA_4757 (.A(net982));
 sg13g2_antennanp ANTENNA_4758 (.A(net982));
 sg13g2_antennanp ANTENNA_4759 (.A(net982));
 sg13g2_antennanp ANTENNA_4760 (.A(net982));
 sg13g2_antennanp ANTENNA_4761 (.A(net982));
 sg13g2_antennanp ANTENNA_4762 (.A(net982));
 sg13g2_antennanp ANTENNA_4763 (.A(net982));
 sg13g2_antennanp ANTENNA_4764 (.A(net982));
 sg13g2_antennanp ANTENNA_4765 (.A(net982));
 sg13g2_antennanp ANTENNA_4766 (.A(net982));
 sg13g2_antennanp ANTENNA_4767 (.A(net982));
 sg13g2_antennanp ANTENNA_4768 (.A(net982));
 sg13g2_antennanp ANTENNA_4769 (.A(net982));
 sg13g2_antennanp ANTENNA_4770 (.A(net982));
 sg13g2_antennanp ANTENNA_4771 (.A(net982));
 sg13g2_antennanp ANTENNA_4772 (.A(net982));
 sg13g2_antennanp ANTENNA_4773 (.A(net982));
 sg13g2_antennanp ANTENNA_4774 (.A(net982));
 sg13g2_antennanp ANTENNA_4775 (.A(net989));
 sg13g2_antennanp ANTENNA_4776 (.A(net989));
 sg13g2_antennanp ANTENNA_4777 (.A(net989));
 sg13g2_antennanp ANTENNA_4778 (.A(net989));
 sg13g2_antennanp ANTENNA_4779 (.A(net989));
 sg13g2_antennanp ANTENNA_4780 (.A(net989));
 sg13g2_antennanp ANTENNA_4781 (.A(net989));
 sg13g2_antennanp ANTENNA_4782 (.A(net989));
 sg13g2_antennanp ANTENNA_4783 (.A(net989));
 sg13g2_antennanp ANTENNA_4784 (.A(net990));
 sg13g2_antennanp ANTENNA_4785 (.A(net990));
 sg13g2_antennanp ANTENNA_4786 (.A(net990));
 sg13g2_antennanp ANTENNA_4787 (.A(net990));
 sg13g2_antennanp ANTENNA_4788 (.A(net990));
 sg13g2_antennanp ANTENNA_4789 (.A(net990));
 sg13g2_antennanp ANTENNA_4790 (.A(net990));
 sg13g2_antennanp ANTENNA_4791 (.A(net990));
 sg13g2_antennanp ANTENNA_4792 (.A(net990));
 sg13g2_antennanp ANTENNA_4793 (.A(net1051));
 sg13g2_antennanp ANTENNA_4794 (.A(net1051));
 sg13g2_antennanp ANTENNA_4795 (.A(net1051));
 sg13g2_antennanp ANTENNA_4796 (.A(net1051));
 sg13g2_antennanp ANTENNA_4797 (.A(net1051));
 sg13g2_antennanp ANTENNA_4798 (.A(net1051));
 sg13g2_antennanp ANTENNA_4799 (.A(net1051));
 sg13g2_antennanp ANTENNA_4800 (.A(net1051));
 sg13g2_antennanp ANTENNA_4801 (.A(net1051));
 sg13g2_antennanp ANTENNA_4802 (.A(net1053));
 sg13g2_antennanp ANTENNA_4803 (.A(net1053));
 sg13g2_antennanp ANTENNA_4804 (.A(net1053));
 sg13g2_antennanp ANTENNA_4805 (.A(net1053));
 sg13g2_antennanp ANTENNA_4806 (.A(net1053));
 sg13g2_antennanp ANTENNA_4807 (.A(net1053));
 sg13g2_antennanp ANTENNA_4808 (.A(net1053));
 sg13g2_antennanp ANTENNA_4809 (.A(net1053));
 sg13g2_antennanp ANTENNA_4810 (.A(net1053));
 sg13g2_antennanp ANTENNA_4811 (.A(net1054));
 sg13g2_antennanp ANTENNA_4812 (.A(net1054));
 sg13g2_antennanp ANTENNA_4813 (.A(net1054));
 sg13g2_antennanp ANTENNA_4814 (.A(net1054));
 sg13g2_antennanp ANTENNA_4815 (.A(net1054));
 sg13g2_antennanp ANTENNA_4816 (.A(net1054));
 sg13g2_antennanp ANTENNA_4817 (.A(net1054));
 sg13g2_antennanp ANTENNA_4818 (.A(net1054));
 sg13g2_antennanp ANTENNA_4819 (.A(net1054));
 sg13g2_antennanp ANTENNA_4820 (.A(net1100));
 sg13g2_antennanp ANTENNA_4821 (.A(net1100));
 sg13g2_antennanp ANTENNA_4822 (.A(net1100));
 sg13g2_antennanp ANTENNA_4823 (.A(net1100));
 sg13g2_antennanp ANTENNA_4824 (.A(net1100));
 sg13g2_antennanp ANTENNA_4825 (.A(net1100));
 sg13g2_antennanp ANTENNA_4826 (.A(net1100));
 sg13g2_antennanp ANTENNA_4827 (.A(net1100));
 sg13g2_antennanp ANTENNA_4828 (.A(net1100));
 sg13g2_antennanp ANTENNA_4829 (.A(net1192));
 sg13g2_antennanp ANTENNA_4830 (.A(net1192));
 sg13g2_antennanp ANTENNA_4831 (.A(net1192));
 sg13g2_antennanp ANTENNA_4832 (.A(net1192));
 sg13g2_antennanp ANTENNA_4833 (.A(net1192));
 sg13g2_antennanp ANTENNA_4834 (.A(net1192));
 sg13g2_antennanp ANTENNA_4835 (.A(net1192));
 sg13g2_antennanp ANTENNA_4836 (.A(net1192));
 sg13g2_antennanp ANTENNA_4837 (.A(net1192));
 sg13g2_antennanp ANTENNA_4838 (.A(net1192));
 sg13g2_antennanp ANTENNA_4839 (.A(net1192));
 sg13g2_antennanp ANTENNA_4840 (.A(net1192));
 sg13g2_antennanp ANTENNA_4841 (.A(net1192));
 sg13g2_antennanp ANTENNA_4842 (.A(net1192));
 sg13g2_antennanp ANTENNA_4843 (.A(net1192));
 sg13g2_antennanp ANTENNA_4844 (.A(net1192));
 sg13g2_antennanp ANTENNA_4845 (.A(net1192));
 sg13g2_antennanp ANTENNA_4846 (.A(net1192));
 sg13g2_antennanp ANTENNA_4847 (.A(net1192));
 sg13g2_antennanp ANTENNA_4848 (.A(net1192));
 sg13g2_antennanp ANTENNA_4849 (.A(net1273));
 sg13g2_antennanp ANTENNA_4850 (.A(net1273));
 sg13g2_antennanp ANTENNA_4851 (.A(net1273));
 sg13g2_antennanp ANTENNA_4852 (.A(net1273));
 sg13g2_antennanp ANTENNA_4853 (.A(net1273));
 sg13g2_antennanp ANTENNA_4854 (.A(net1273));
 sg13g2_antennanp ANTENNA_4855 (.A(net1273));
 sg13g2_antennanp ANTENNA_4856 (.A(net1273));
 sg13g2_antennanp ANTENNA_4857 (.A(net1273));
 sg13g2_antennanp ANTENNA_4858 (.A(net1276));
 sg13g2_antennanp ANTENNA_4859 (.A(net1276));
 sg13g2_antennanp ANTENNA_4860 (.A(net1276));
 sg13g2_antennanp ANTENNA_4861 (.A(net1276));
 sg13g2_antennanp ANTENNA_4862 (.A(net1276));
 sg13g2_antennanp ANTENNA_4863 (.A(net1276));
 sg13g2_antennanp ANTENNA_4864 (.A(net1276));
 sg13g2_antennanp ANTENNA_4865 (.A(net1276));
 sg13g2_antennanp ANTENNA_4866 (.A(net1276));
 sg13g2_antennanp ANTENNA_4867 (.A(net1276));
 sg13g2_antennanp ANTENNA_4868 (.A(net1276));
 sg13g2_antennanp ANTENNA_4869 (.A(net1276));
 sg13g2_antennanp ANTENNA_4870 (.A(net1276));
 sg13g2_antennanp ANTENNA_4871 (.A(net1276));
 sg13g2_antennanp ANTENNA_4872 (.A(net1276));
 sg13g2_antennanp ANTENNA_4873 (.A(net1276));
 sg13g2_antennanp ANTENNA_4874 (.A(net1276));
 sg13g2_antennanp ANTENNA_4875 (.A(net1276));
 sg13g2_antennanp ANTENNA_4876 (.A(net1276));
 sg13g2_antennanp ANTENNA_4877 (.A(net1276));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_fill_2 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_55 ();
 sg13g2_decap_8 FILLER_0_62 ();
 sg13g2_decap_8 FILLER_0_69 ();
 sg13g2_decap_8 FILLER_0_76 ();
 sg13g2_fill_2 FILLER_0_83 ();
 sg13g2_decap_8 FILLER_0_89 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_117 ();
 sg13g2_decap_4 FILLER_0_124 ();
 sg13g2_fill_2 FILLER_0_128 ();
 sg13g2_decap_4 FILLER_0_156 ();
 sg13g2_fill_2 FILLER_0_160 ();
 sg13g2_decap_4 FILLER_0_166 ();
 sg13g2_decap_4 FILLER_0_178 ();
 sg13g2_fill_1 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_4 FILLER_0_198 ();
 sg13g2_fill_1 FILLER_0_202 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_fill_1 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_fill_2 FILLER_0_256 ();
 sg13g2_fill_2 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_4 FILLER_0_275 ();
 sg13g2_fill_2 FILLER_0_279 ();
 sg13g2_decap_4 FILLER_0_285 ();
 sg13g2_fill_2 FILLER_0_289 ();
 sg13g2_decap_4 FILLER_0_295 ();
 sg13g2_fill_2 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_4 FILLER_0_352 ();
 sg13g2_fill_1 FILLER_0_356 ();
 sg13g2_fill_2 FILLER_0_361 ();
 sg13g2_decap_4 FILLER_0_367 ();
 sg13g2_fill_2 FILLER_0_371 ();
 sg13g2_fill_1 FILLER_0_376 ();
 sg13g2_fill_1 FILLER_0_454 ();
 sg13g2_fill_2 FILLER_0_483 ();
 sg13g2_fill_1 FILLER_0_493 ();
 sg13g2_decap_8 FILLER_0_520 ();
 sg13g2_decap_8 FILLER_0_527 ();
 sg13g2_decap_4 FILLER_0_534 ();
 sg13g2_decap_8 FILLER_0_542 ();
 sg13g2_fill_2 FILLER_0_549 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_4 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_617 ();
 sg13g2_decap_8 FILLER_0_624 ();
 sg13g2_decap_8 FILLER_0_631 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_671 ();
 sg13g2_decap_8 FILLER_0_678 ();
 sg13g2_decap_8 FILLER_0_685 ();
 sg13g2_fill_2 FILLER_0_692 ();
 sg13g2_decap_4 FILLER_0_698 ();
 sg13g2_decap_4 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_715 ();
 sg13g2_decap_8 FILLER_0_722 ();
 sg13g2_decap_4 FILLER_0_729 ();
 sg13g2_fill_1 FILLER_0_761 ();
 sg13g2_decap_8 FILLER_0_788 ();
 sg13g2_decap_8 FILLER_0_795 ();
 sg13g2_decap_8 FILLER_0_802 ();
 sg13g2_decap_8 FILLER_0_809 ();
 sg13g2_decap_8 FILLER_0_816 ();
 sg13g2_decap_8 FILLER_0_823 ();
 sg13g2_decap_8 FILLER_0_830 ();
 sg13g2_decap_8 FILLER_0_837 ();
 sg13g2_fill_2 FILLER_0_844 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_fill_1 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_4 FILLER_0_903 ();
 sg13g2_fill_2 FILLER_0_907 ();
 sg13g2_decap_8 FILLER_0_935 ();
 sg13g2_decap_4 FILLER_0_942 ();
 sg13g2_decap_4 FILLER_0_1006 ();
 sg13g2_fill_2 FILLER_0_1010 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_0_1029 ();
 sg13g2_decap_8 FILLER_0_1036 ();
 sg13g2_decap_8 FILLER_0_1043 ();
 sg13g2_fill_2 FILLER_0_1050 ();
 sg13g2_decap_4 FILLER_0_1082 ();
 sg13g2_fill_1 FILLER_0_1086 ();
 sg13g2_decap_8 FILLER_0_1117 ();
 sg13g2_decap_4 FILLER_0_1124 ();
 sg13g2_decap_8 FILLER_0_1133 ();
 sg13g2_decap_8 FILLER_0_1140 ();
 sg13g2_decap_4 FILLER_0_1147 ();
 sg13g2_fill_1 FILLER_0_1151 ();
 sg13g2_decap_8 FILLER_0_1156 ();
 sg13g2_decap_8 FILLER_0_1163 ();
 sg13g2_decap_8 FILLER_0_1170 ();
 sg13g2_decap_8 FILLER_0_1177 ();
 sg13g2_decap_8 FILLER_0_1184 ();
 sg13g2_decap_8 FILLER_0_1191 ();
 sg13g2_decap_4 FILLER_0_1198 ();
 sg13g2_fill_1 FILLER_0_1202 ();
 sg13g2_decap_8 FILLER_0_1216 ();
 sg13g2_decap_8 FILLER_0_1223 ();
 sg13g2_fill_2 FILLER_0_1230 ();
 sg13g2_fill_1 FILLER_0_1232 ();
 sg13g2_decap_8 FILLER_0_1263 ();
 sg13g2_fill_2 FILLER_0_1270 ();
 sg13g2_fill_1 FILLER_0_1272 ();
 sg13g2_decap_8 FILLER_0_1277 ();
 sg13g2_decap_4 FILLER_0_1284 ();
 sg13g2_fill_2 FILLER_0_1288 ();
 sg13g2_decap_8 FILLER_0_1294 ();
 sg13g2_decap_8 FILLER_0_1301 ();
 sg13g2_decap_8 FILLER_0_1308 ();
 sg13g2_decap_8 FILLER_0_1315 ();
 sg13g2_decap_8 FILLER_0_1322 ();
 sg13g2_fill_1 FILLER_0_1329 ();
 sg13g2_decap_8 FILLER_0_1334 ();
 sg13g2_decap_8 FILLER_0_1341 ();
 sg13g2_decap_4 FILLER_0_1348 ();
 sg13g2_fill_1 FILLER_0_1352 ();
 sg13g2_fill_2 FILLER_0_1366 ();
 sg13g2_fill_1 FILLER_0_1368 ();
 sg13g2_decap_8 FILLER_0_1373 ();
 sg13g2_decap_8 FILLER_0_1380 ();
 sg13g2_decap_8 FILLER_0_1387 ();
 sg13g2_decap_8 FILLER_0_1394 ();
 sg13g2_decap_4 FILLER_0_1401 ();
 sg13g2_fill_1 FILLER_0_1405 ();
 sg13g2_decap_8 FILLER_0_1432 ();
 sg13g2_fill_2 FILLER_0_1443 ();
 sg13g2_decap_8 FILLER_0_1449 ();
 sg13g2_fill_1 FILLER_0_1456 ();
 sg13g2_fill_1 FILLER_0_1465 ();
 sg13g2_decap_8 FILLER_0_1474 ();
 sg13g2_decap_8 FILLER_0_1481 ();
 sg13g2_decap_8 FILLER_0_1488 ();
 sg13g2_fill_2 FILLER_0_1495 ();
 sg13g2_decap_8 FILLER_0_1501 ();
 sg13g2_fill_1 FILLER_0_1508 ();
 sg13g2_decap_8 FILLER_0_1535 ();
 sg13g2_decap_8 FILLER_0_1542 ();
 sg13g2_decap_4 FILLER_0_1549 ();
 sg13g2_fill_2 FILLER_0_1553 ();
 sg13g2_decap_8 FILLER_0_1585 ();
 sg13g2_decap_8 FILLER_0_1592 ();
 sg13g2_decap_4 FILLER_0_1599 ();
 sg13g2_fill_2 FILLER_0_1603 ();
 sg13g2_decap_8 FILLER_0_1630 ();
 sg13g2_decap_4 FILLER_0_1637 ();
 sg13g2_fill_2 FILLER_0_1641 ();
 sg13g2_decap_8 FILLER_0_1651 ();
 sg13g2_decap_4 FILLER_0_1658 ();
 sg13g2_fill_2 FILLER_0_1662 ();
 sg13g2_decap_8 FILLER_0_1672 ();
 sg13g2_fill_2 FILLER_0_1679 ();
 sg13g2_fill_1 FILLER_0_1681 ();
 sg13g2_decap_8 FILLER_0_1686 ();
 sg13g2_decap_8 FILLER_0_1693 ();
 sg13g2_decap_8 FILLER_0_1700 ();
 sg13g2_decap_8 FILLER_0_1707 ();
 sg13g2_decap_8 FILLER_0_1714 ();
 sg13g2_fill_2 FILLER_0_1721 ();
 sg13g2_fill_1 FILLER_0_1723 ();
 sg13g2_decap_4 FILLER_0_1729 ();
 sg13g2_fill_1 FILLER_0_1733 ();
 sg13g2_fill_2 FILLER_0_1758 ();
 sg13g2_fill_1 FILLER_0_1760 ();
 sg13g2_fill_2 FILLER_0_1766 ();
 sg13g2_decap_8 FILLER_0_1776 ();
 sg13g2_decap_4 FILLER_0_1783 ();
 sg13g2_fill_1 FILLER_0_1787 ();
 sg13g2_decap_4 FILLER_0_1792 ();
 sg13g2_fill_2 FILLER_0_1796 ();
 sg13g2_decap_8 FILLER_0_1802 ();
 sg13g2_decap_8 FILLER_0_1809 ();
 sg13g2_decap_8 FILLER_0_1816 ();
 sg13g2_fill_2 FILLER_0_1823 ();
 sg13g2_decap_4 FILLER_0_1829 ();
 sg13g2_fill_1 FILLER_0_1837 ();
 sg13g2_fill_2 FILLER_0_1842 ();
 sg13g2_fill_1 FILLER_0_1844 ();
 sg13g2_decap_8 FILLER_0_1875 ();
 sg13g2_decap_8 FILLER_0_1882 ();
 sg13g2_fill_2 FILLER_0_1889 ();
 sg13g2_fill_1 FILLER_0_1895 ();
 sg13g2_decap_8 FILLER_0_1900 ();
 sg13g2_decap_4 FILLER_0_1907 ();
 sg13g2_fill_1 FILLER_0_1911 ();
 sg13g2_decap_8 FILLER_0_1929 ();
 sg13g2_decap_8 FILLER_0_1936 ();
 sg13g2_decap_8 FILLER_0_1943 ();
 sg13g2_decap_8 FILLER_0_1950 ();
 sg13g2_decap_8 FILLER_0_1957 ();
 sg13g2_decap_8 FILLER_0_1964 ();
 sg13g2_decap_4 FILLER_0_1971 ();
 sg13g2_fill_2 FILLER_0_1975 ();
 sg13g2_fill_2 FILLER_0_1981 ();
 sg13g2_decap_8 FILLER_0_1987 ();
 sg13g2_fill_2 FILLER_0_1994 ();
 sg13g2_fill_1 FILLER_0_1996 ();
 sg13g2_decap_8 FILLER_0_2031 ();
 sg13g2_decap_8 FILLER_0_2038 ();
 sg13g2_decap_8 FILLER_0_2045 ();
 sg13g2_fill_1 FILLER_0_2052 ();
 sg13g2_fill_1 FILLER_0_2057 ();
 sg13g2_decap_8 FILLER_0_2084 ();
 sg13g2_decap_4 FILLER_0_2091 ();
 sg13g2_fill_2 FILLER_0_2095 ();
 sg13g2_decap_8 FILLER_0_2105 ();
 sg13g2_decap_8 FILLER_0_2112 ();
 sg13g2_decap_8 FILLER_0_2131 ();
 sg13g2_fill_1 FILLER_0_2138 ();
 sg13g2_decap_8 FILLER_0_2148 ();
 sg13g2_decap_8 FILLER_0_2155 ();
 sg13g2_decap_8 FILLER_0_2162 ();
 sg13g2_decap_8 FILLER_0_2169 ();
 sg13g2_decap_8 FILLER_0_2176 ();
 sg13g2_decap_8 FILLER_0_2183 ();
 sg13g2_decap_8 FILLER_0_2190 ();
 sg13g2_decap_8 FILLER_0_2197 ();
 sg13g2_decap_8 FILLER_0_2204 ();
 sg13g2_decap_8 FILLER_0_2211 ();
 sg13g2_decap_8 FILLER_0_2218 ();
 sg13g2_decap_8 FILLER_0_2225 ();
 sg13g2_decap_8 FILLER_0_2232 ();
 sg13g2_decap_8 FILLER_0_2239 ();
 sg13g2_decap_8 FILLER_0_2246 ();
 sg13g2_decap_8 FILLER_0_2253 ();
 sg13g2_decap_8 FILLER_0_2260 ();
 sg13g2_decap_8 FILLER_0_2267 ();
 sg13g2_decap_8 FILLER_0_2274 ();
 sg13g2_decap_8 FILLER_0_2281 ();
 sg13g2_decap_8 FILLER_0_2288 ();
 sg13g2_decap_8 FILLER_0_2295 ();
 sg13g2_decap_8 FILLER_0_2302 ();
 sg13g2_decap_8 FILLER_0_2309 ();
 sg13g2_decap_8 FILLER_0_2316 ();
 sg13g2_decap_8 FILLER_0_2323 ();
 sg13g2_fill_2 FILLER_0_2330 ();
 sg13g2_fill_1 FILLER_0_2332 ();
 sg13g2_decap_8 FILLER_0_2359 ();
 sg13g2_decap_8 FILLER_0_2366 ();
 sg13g2_decap_4 FILLER_0_2373 ();
 sg13g2_fill_1 FILLER_0_2377 ();
 sg13g2_decap_4 FILLER_0_2382 ();
 sg13g2_fill_2 FILLER_0_2386 ();
 sg13g2_decap_8 FILLER_0_2392 ();
 sg13g2_decap_8 FILLER_0_2416 ();
 sg13g2_decap_8 FILLER_0_2423 ();
 sg13g2_decap_8 FILLER_0_2430 ();
 sg13g2_decap_8 FILLER_0_2437 ();
 sg13g2_decap_8 FILLER_0_2444 ();
 sg13g2_decap_8 FILLER_0_2451 ();
 sg13g2_decap_8 FILLER_0_2458 ();
 sg13g2_decap_8 FILLER_0_2465 ();
 sg13g2_decap_8 FILLER_0_2472 ();
 sg13g2_decap_8 FILLER_0_2483 ();
 sg13g2_decap_8 FILLER_0_2490 ();
 sg13g2_decap_8 FILLER_0_2497 ();
 sg13g2_decap_8 FILLER_0_2504 ();
 sg13g2_decap_4 FILLER_0_2511 ();
 sg13g2_decap_8 FILLER_0_2519 ();
 sg13g2_decap_8 FILLER_0_2526 ();
 sg13g2_decap_8 FILLER_0_2533 ();
 sg13g2_decap_8 FILLER_0_2540 ();
 sg13g2_decap_8 FILLER_0_2547 ();
 sg13g2_decap_8 FILLER_0_2554 ();
 sg13g2_decap_8 FILLER_0_2561 ();
 sg13g2_decap_8 FILLER_0_2568 ();
 sg13g2_decap_8 FILLER_0_2575 ();
 sg13g2_decap_8 FILLER_0_2582 ();
 sg13g2_decap_8 FILLER_0_2589 ();
 sg13g2_decap_8 FILLER_0_2596 ();
 sg13g2_decap_8 FILLER_0_2603 ();
 sg13g2_decap_8 FILLER_0_2610 ();
 sg13g2_decap_8 FILLER_0_2617 ();
 sg13g2_decap_8 FILLER_0_2624 ();
 sg13g2_decap_8 FILLER_0_2631 ();
 sg13g2_decap_8 FILLER_0_2638 ();
 sg13g2_decap_8 FILLER_0_2645 ();
 sg13g2_decap_8 FILLER_0_2652 ();
 sg13g2_decap_8 FILLER_0_2659 ();
 sg13g2_decap_4 FILLER_0_2666 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_fill_2 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_44 ();
 sg13g2_fill_2 FILLER_1_71 ();
 sg13g2_fill_1 FILLER_1_73 ();
 sg13g2_fill_2 FILLER_1_78 ();
 sg13g2_decap_8 FILLER_1_110 ();
 sg13g2_decap_8 FILLER_1_117 ();
 sg13g2_fill_2 FILLER_1_124 ();
 sg13g2_fill_1 FILLER_1_126 ();
 sg13g2_decap_4 FILLER_1_131 ();
 sg13g2_fill_2 FILLER_1_135 ();
 sg13g2_decap_8 FILLER_1_141 ();
 sg13g2_fill_2 FILLER_1_153 ();
 sg13g2_fill_2 FILLER_1_163 ();
 sg13g2_decap_4 FILLER_1_248 ();
 sg13g2_fill_2 FILLER_1_252 ();
 sg13g2_fill_1 FILLER_1_267 ();
 sg13g2_decap_4 FILLER_1_302 ();
 sg13g2_fill_1 FILLER_1_306 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_4 FILLER_1_344 ();
 sg13g2_fill_2 FILLER_1_348 ();
 sg13g2_fill_1 FILLER_1_376 ();
 sg13g2_fill_1 FILLER_1_387 ();
 sg13g2_fill_2 FILLER_1_470 ();
 sg13g2_fill_1 FILLER_1_503 ();
 sg13g2_decap_8 FILLER_1_519 ();
 sg13g2_fill_2 FILLER_1_526 ();
 sg13g2_fill_2 FILLER_1_558 ();
 sg13g2_decap_4 FILLER_1_603 ();
 sg13g2_decap_8 FILLER_1_676 ();
 sg13g2_decap_4 FILLER_1_683 ();
 sg13g2_fill_2 FILLER_1_758 ();
 sg13g2_fill_1 FILLER_1_760 ();
 sg13g2_fill_2 FILLER_1_818 ();
 sg13g2_fill_1 FILLER_1_820 ();
 sg13g2_decap_8 FILLER_1_825 ();
 sg13g2_decap_8 FILLER_1_832 ();
 sg13g2_fill_1 FILLER_1_839 ();
 sg13g2_fill_2 FILLER_1_910 ();
 sg13g2_fill_1 FILLER_1_912 ();
 sg13g2_fill_2 FILLER_1_986 ();
 sg13g2_fill_2 FILLER_1_992 ();
 sg13g2_decap_8 FILLER_1_1028 ();
 sg13g2_fill_1 FILLER_1_1035 ();
 sg13g2_fill_1 FILLER_1_1056 ();
 sg13g2_fill_2 FILLER_1_1083 ();
 sg13g2_fill_2 FILLER_1_1090 ();
 sg13g2_fill_1 FILLER_1_1132 ();
 sg13g2_decap_4 FILLER_1_1171 ();
 sg13g2_decap_4 FILLER_1_1179 ();
 sg13g2_fill_1 FILLER_1_1217 ();
 sg13g2_decap_4 FILLER_1_1223 ();
 sg13g2_fill_2 FILLER_1_1227 ();
 sg13g2_fill_1 FILLER_1_1233 ();
 sg13g2_decap_4 FILLER_1_1239 ();
 sg13g2_fill_1 FILLER_1_1243 ();
 sg13g2_fill_1 FILLER_1_1313 ();
 sg13g2_decap_8 FILLER_1_1344 ();
 sg13g2_fill_1 FILLER_1_1351 ();
 sg13g2_fill_2 FILLER_1_1356 ();
 sg13g2_fill_1 FILLER_1_1389 ();
 sg13g2_decap_8 FILLER_1_1489 ();
 sg13g2_decap_4 FILLER_1_1496 ();
 sg13g2_fill_1 FILLER_1_1513 ();
 sg13g2_fill_2 FILLER_1_1518 ();
 sg13g2_decap_8 FILLER_1_1546 ();
 sg13g2_decap_8 FILLER_1_1553 ();
 sg13g2_decap_8 FILLER_1_1564 ();
 sg13g2_decap_4 FILLER_1_1571 ();
 sg13g2_fill_1 FILLER_1_1579 ();
 sg13g2_fill_1 FILLER_1_1585 ();
 sg13g2_fill_1 FILLER_1_1625 ();
 sg13g2_fill_1 FILLER_1_1676 ();
 sg13g2_decap_8 FILLER_1_1707 ();
 sg13g2_fill_1 FILLER_1_1788 ();
 sg13g2_fill_1 FILLER_1_1815 ();
 sg13g2_fill_1 FILLER_1_1842 ();
 sg13g2_fill_2 FILLER_1_1877 ();
 sg13g2_fill_1 FILLER_1_1888 ();
 sg13g2_fill_2 FILLER_1_1915 ();
 sg13g2_fill_1 FILLER_1_1917 ();
 sg13g2_fill_1 FILLER_1_2000 ();
 sg13g2_decap_8 FILLER_1_2027 ();
 sg13g2_decap_8 FILLER_1_2034 ();
 sg13g2_fill_1 FILLER_1_2041 ();
 sg13g2_fill_2 FILLER_1_2072 ();
 sg13g2_decap_8 FILLER_1_2078 ();
 sg13g2_fill_1 FILLER_1_2085 ();
 sg13g2_decap_8 FILLER_1_2159 ();
 sg13g2_decap_8 FILLER_1_2166 ();
 sg13g2_decap_8 FILLER_1_2173 ();
 sg13g2_decap_8 FILLER_1_2180 ();
 sg13g2_decap_8 FILLER_1_2187 ();
 sg13g2_decap_8 FILLER_1_2194 ();
 sg13g2_decap_8 FILLER_1_2201 ();
 sg13g2_decap_8 FILLER_1_2208 ();
 sg13g2_decap_8 FILLER_1_2215 ();
 sg13g2_decap_8 FILLER_1_2222 ();
 sg13g2_decap_8 FILLER_1_2229 ();
 sg13g2_decap_8 FILLER_1_2236 ();
 sg13g2_decap_8 FILLER_1_2243 ();
 sg13g2_decap_8 FILLER_1_2250 ();
 sg13g2_decap_8 FILLER_1_2257 ();
 sg13g2_decap_8 FILLER_1_2264 ();
 sg13g2_decap_8 FILLER_1_2271 ();
 sg13g2_decap_8 FILLER_1_2278 ();
 sg13g2_decap_8 FILLER_1_2285 ();
 sg13g2_decap_8 FILLER_1_2292 ();
 sg13g2_decap_8 FILLER_1_2299 ();
 sg13g2_fill_1 FILLER_1_2306 ();
 sg13g2_decap_8 FILLER_1_2333 ();
 sg13g2_fill_1 FILLER_1_2418 ();
 sg13g2_decap_8 FILLER_1_2445 ();
 sg13g2_decap_8 FILLER_1_2452 ();
 sg13g2_decap_8 FILLER_1_2459 ();
 sg13g2_fill_2 FILLER_1_2466 ();
 sg13g2_fill_1 FILLER_1_2468 ();
 sg13g2_fill_2 FILLER_1_2499 ();
 sg13g2_fill_1 FILLER_1_2501 ();
 sg13g2_decap_8 FILLER_1_2532 ();
 sg13g2_decap_8 FILLER_1_2539 ();
 sg13g2_decap_8 FILLER_1_2546 ();
 sg13g2_decap_8 FILLER_1_2553 ();
 sg13g2_decap_8 FILLER_1_2560 ();
 sg13g2_decap_8 FILLER_1_2567 ();
 sg13g2_decap_8 FILLER_1_2574 ();
 sg13g2_decap_8 FILLER_1_2581 ();
 sg13g2_decap_8 FILLER_1_2588 ();
 sg13g2_decap_8 FILLER_1_2595 ();
 sg13g2_decap_8 FILLER_1_2602 ();
 sg13g2_decap_8 FILLER_1_2609 ();
 sg13g2_decap_8 FILLER_1_2616 ();
 sg13g2_decap_8 FILLER_1_2623 ();
 sg13g2_decap_8 FILLER_1_2630 ();
 sg13g2_decap_8 FILLER_1_2637 ();
 sg13g2_decap_8 FILLER_1_2644 ();
 sg13g2_decap_8 FILLER_1_2651 ();
 sg13g2_decap_8 FILLER_1_2658 ();
 sg13g2_decap_4 FILLER_1_2665 ();
 sg13g2_fill_1 FILLER_1_2669 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_38 ();
 sg13g2_fill_1 FILLER_2_74 ();
 sg13g2_fill_1 FILLER_2_80 ();
 sg13g2_fill_1 FILLER_2_86 ();
 sg13g2_fill_2 FILLER_2_91 ();
 sg13g2_fill_2 FILLER_2_185 ();
 sg13g2_fill_2 FILLER_2_192 ();
 sg13g2_fill_1 FILLER_2_194 ();
 sg13g2_decap_4 FILLER_2_221 ();
 sg13g2_fill_1 FILLER_2_225 ();
 sg13g2_fill_2 FILLER_2_256 ();
 sg13g2_fill_1 FILLER_2_258 ();
 sg13g2_fill_2 FILLER_2_263 ();
 sg13g2_fill_1 FILLER_2_291 ();
 sg13g2_fill_2 FILLER_2_297 ();
 sg13g2_fill_1 FILLER_2_299 ();
 sg13g2_fill_2 FILLER_2_305 ();
 sg13g2_fill_1 FILLER_2_307 ();
 sg13g2_fill_2 FILLER_2_321 ();
 sg13g2_fill_2 FILLER_2_353 ();
 sg13g2_fill_1 FILLER_2_355 ();
 sg13g2_fill_2 FILLER_2_382 ();
 sg13g2_fill_1 FILLER_2_414 ();
 sg13g2_fill_1 FILLER_2_444 ();
 sg13g2_fill_2 FILLER_2_551 ();
 sg13g2_fill_2 FILLER_2_557 ();
 sg13g2_fill_1 FILLER_2_559 ();
 sg13g2_fill_1 FILLER_2_603 ();
 sg13g2_fill_1 FILLER_2_609 ();
 sg13g2_fill_1 FILLER_2_636 ();
 sg13g2_fill_2 FILLER_2_641 ();
 sg13g2_fill_1 FILLER_2_648 ();
 sg13g2_fill_2 FILLER_2_653 ();
 sg13g2_decap_4 FILLER_2_659 ();
 sg13g2_fill_1 FILLER_2_724 ();
 sg13g2_fill_1 FILLER_2_751 ();
 sg13g2_fill_1 FILLER_2_765 ();
 sg13g2_fill_2 FILLER_2_784 ();
 sg13g2_fill_1 FILLER_2_786 ();
 sg13g2_fill_1 FILLER_2_813 ();
 sg13g2_fill_2 FILLER_2_893 ();
 sg13g2_fill_1 FILLER_2_895 ();
 sg13g2_fill_2 FILLER_2_904 ();
 sg13g2_decap_4 FILLER_2_920 ();
 sg13g2_fill_2 FILLER_2_928 ();
 sg13g2_fill_2 FILLER_2_981 ();
 sg13g2_fill_2 FILLER_2_1015 ();
 sg13g2_fill_2 FILLER_2_1074 ();
 sg13g2_fill_2 FILLER_2_1102 ();
 sg13g2_fill_1 FILLER_2_1104 ();
 sg13g2_decap_4 FILLER_2_1182 ();
 sg13g2_fill_2 FILLER_2_1186 ();
 sg13g2_fill_2 FILLER_2_1222 ();
 sg13g2_decap_4 FILLER_2_1229 ();
 sg13g2_fill_2 FILLER_2_1233 ();
 sg13g2_fill_1 FILLER_2_1239 ();
 sg13g2_fill_2 FILLER_2_1278 ();
 sg13g2_fill_2 FILLER_2_1324 ();
 sg13g2_fill_1 FILLER_2_1326 ();
 sg13g2_fill_2 FILLER_2_1392 ();
 sg13g2_fill_2 FILLER_2_1441 ();
 sg13g2_fill_1 FILLER_2_1443 ();
 sg13g2_fill_2 FILLER_2_1449 ();
 sg13g2_fill_2 FILLER_2_1456 ();
 sg13g2_fill_1 FILLER_2_1489 ();
 sg13g2_fill_1 FILLER_2_1525 ();
 sg13g2_fill_1 FILLER_2_1569 ();
 sg13g2_fill_2 FILLER_2_1596 ();
 sg13g2_fill_2 FILLER_2_1624 ();
 sg13g2_fill_1 FILLER_2_1626 ();
 sg13g2_fill_1 FILLER_2_1662 ();
 sg13g2_fill_1 FILLER_2_1667 ();
 sg13g2_decap_8 FILLER_2_1699 ();
 sg13g2_fill_2 FILLER_2_1706 ();
 sg13g2_fill_1 FILLER_2_1708 ();
 sg13g2_fill_1 FILLER_2_1813 ();
 sg13g2_fill_2 FILLER_2_1840 ();
 sg13g2_fill_1 FILLER_2_1842 ();
 sg13g2_fill_2 FILLER_2_1869 ();
 sg13g2_fill_2 FILLER_2_1910 ();
 sg13g2_fill_1 FILLER_2_1912 ();
 sg13g2_fill_2 FILLER_2_1939 ();
 sg13g2_fill_1 FILLER_2_1941 ();
 sg13g2_fill_1 FILLER_2_1972 ();
 sg13g2_fill_1 FILLER_2_1987 ();
 sg13g2_fill_1 FILLER_2_1993 ();
 sg13g2_fill_1 FILLER_2_1999 ();
 sg13g2_fill_2 FILLER_2_2039 ();
 sg13g2_fill_1 FILLER_2_2055 ();
 sg13g2_fill_1 FILLER_2_2060 ();
 sg13g2_fill_1 FILLER_2_2087 ();
 sg13g2_fill_2 FILLER_2_2092 ();
 sg13g2_fill_1 FILLER_2_2120 ();
 sg13g2_fill_2 FILLER_2_2131 ();
 sg13g2_fill_1 FILLER_2_2142 ();
 sg13g2_decap_8 FILLER_2_2172 ();
 sg13g2_decap_8 FILLER_2_2179 ();
 sg13g2_decap_8 FILLER_2_2186 ();
 sg13g2_decap_8 FILLER_2_2193 ();
 sg13g2_decap_8 FILLER_2_2200 ();
 sg13g2_decap_8 FILLER_2_2207 ();
 sg13g2_decap_8 FILLER_2_2214 ();
 sg13g2_decap_8 FILLER_2_2221 ();
 sg13g2_decap_8 FILLER_2_2228 ();
 sg13g2_decap_8 FILLER_2_2235 ();
 sg13g2_decap_8 FILLER_2_2242 ();
 sg13g2_decap_8 FILLER_2_2249 ();
 sg13g2_decap_8 FILLER_2_2256 ();
 sg13g2_decap_8 FILLER_2_2263 ();
 sg13g2_decap_8 FILLER_2_2270 ();
 sg13g2_decap_4 FILLER_2_2277 ();
 sg13g2_fill_2 FILLER_2_2281 ();
 sg13g2_decap_8 FILLER_2_2317 ();
 sg13g2_fill_2 FILLER_2_2324 ();
 sg13g2_fill_1 FILLER_2_2326 ();
 sg13g2_fill_2 FILLER_2_2337 ();
 sg13g2_fill_1 FILLER_2_2339 ();
 sg13g2_fill_2 FILLER_2_2344 ();
 sg13g2_fill_1 FILLER_2_2346 ();
 sg13g2_decap_8 FILLER_2_2351 ();
 sg13g2_decap_4 FILLER_2_2383 ();
 sg13g2_fill_1 FILLER_2_2392 ();
 sg13g2_fill_1 FILLER_2_2423 ();
 sg13g2_fill_2 FILLER_2_2541 ();
 sg13g2_decap_8 FILLER_2_2547 ();
 sg13g2_decap_8 FILLER_2_2554 ();
 sg13g2_decap_8 FILLER_2_2561 ();
 sg13g2_decap_8 FILLER_2_2568 ();
 sg13g2_decap_8 FILLER_2_2575 ();
 sg13g2_decap_8 FILLER_2_2582 ();
 sg13g2_decap_8 FILLER_2_2589 ();
 sg13g2_decap_8 FILLER_2_2596 ();
 sg13g2_decap_8 FILLER_2_2603 ();
 sg13g2_decap_8 FILLER_2_2610 ();
 sg13g2_decap_8 FILLER_2_2617 ();
 sg13g2_decap_8 FILLER_2_2624 ();
 sg13g2_decap_8 FILLER_2_2631 ();
 sg13g2_decap_8 FILLER_2_2638 ();
 sg13g2_decap_8 FILLER_2_2645 ();
 sg13g2_decap_8 FILLER_2_2652 ();
 sg13g2_decap_8 FILLER_2_2659 ();
 sg13g2_decap_4 FILLER_2_2666 ();
 sg13g2_decap_4 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_4 ();
 sg13g2_fill_2 FILLER_3_76 ();
 sg13g2_fill_1 FILLER_3_108 ();
 sg13g2_decap_8 FILLER_3_114 ();
 sg13g2_fill_2 FILLER_3_121 ();
 sg13g2_fill_1 FILLER_3_123 ();
 sg13g2_fill_2 FILLER_3_180 ();
 sg13g2_fill_1 FILLER_3_255 ();
 sg13g2_fill_1 FILLER_3_282 ();
 sg13g2_fill_2 FILLER_3_304 ();
 sg13g2_fill_1 FILLER_3_337 ();
 sg13g2_fill_1 FILLER_3_351 ();
 sg13g2_fill_1 FILLER_3_425 ();
 sg13g2_fill_1 FILLER_3_431 ();
 sg13g2_fill_2 FILLER_3_518 ();
 sg13g2_fill_1 FILLER_3_520 ();
 sg13g2_fill_2 FILLER_3_547 ();
 sg13g2_fill_1 FILLER_3_575 ();
 sg13g2_fill_2 FILLER_3_669 ();
 sg13g2_fill_2 FILLER_3_726 ();
 sg13g2_fill_1 FILLER_3_728 ();
 sg13g2_fill_2 FILLER_3_755 ();
 sg13g2_fill_1 FILLER_3_765 ();
 sg13g2_decap_8 FILLER_3_804 ();
 sg13g2_decap_4 FILLER_3_811 ();
 sg13g2_fill_1 FILLER_3_815 ();
 sg13g2_decap_4 FILLER_3_842 ();
 sg13g2_fill_1 FILLER_3_846 ();
 sg13g2_decap_8 FILLER_3_851 ();
 sg13g2_fill_1 FILLER_3_867 ();
 sg13g2_fill_2 FILLER_3_936 ();
 sg13g2_fill_1 FILLER_3_1007 ();
 sg13g2_fill_1 FILLER_3_1016 ();
 sg13g2_fill_2 FILLER_3_1048 ();
 sg13g2_fill_1 FILLER_3_1050 ();
 sg13g2_fill_2 FILLER_3_1055 ();
 sg13g2_decap_4 FILLER_3_1087 ();
 sg13g2_fill_1 FILLER_3_1095 ();
 sg13g2_fill_2 FILLER_3_1130 ();
 sg13g2_fill_1 FILLER_3_1132 ();
 sg13g2_decap_4 FILLER_3_1159 ();
 sg13g2_decap_8 FILLER_3_1167 ();
 sg13g2_decap_4 FILLER_3_1174 ();
 sg13g2_fill_1 FILLER_3_1178 ();
 sg13g2_fill_1 FILLER_3_1218 ();
 sg13g2_fill_1 FILLER_3_1349 ();
 sg13g2_fill_1 FILLER_3_1354 ();
 sg13g2_fill_1 FILLER_3_1359 ();
 sg13g2_fill_2 FILLER_3_1386 ();
 sg13g2_fill_1 FILLER_3_1416 ();
 sg13g2_fill_2 FILLER_3_1429 ();
 sg13g2_fill_2 FILLER_3_1435 ();
 sg13g2_decap_8 FILLER_3_1471 ();
 sg13g2_fill_1 FILLER_3_1482 ();
 sg13g2_fill_2 FILLER_3_1509 ();
 sg13g2_decap_4 FILLER_3_1536 ();
 sg13g2_fill_2 FILLER_3_1540 ();
 sg13g2_fill_1 FILLER_3_1581 ();
 sg13g2_fill_1 FILLER_3_1632 ();
 sg13g2_fill_2 FILLER_3_1637 ();
 sg13g2_fill_2 FILLER_3_1669 ();
 sg13g2_fill_1 FILLER_3_1675 ();
 sg13g2_decap_8 FILLER_3_1706 ();
 sg13g2_fill_2 FILLER_3_1713 ();
 sg13g2_fill_1 FILLER_3_1715 ();
 sg13g2_fill_1 FILLER_3_1720 ();
 sg13g2_fill_2 FILLER_3_1725 ();
 sg13g2_fill_2 FILLER_3_1761 ();
 sg13g2_fill_1 FILLER_3_1763 ();
 sg13g2_fill_2 FILLER_3_1785 ();
 sg13g2_fill_2 FILLER_3_1792 ();
 sg13g2_decap_4 FILLER_3_1811 ();
 sg13g2_fill_1 FILLER_3_1815 ();
 sg13g2_fill_2 FILLER_3_1843 ();
 sg13g2_fill_1 FILLER_3_1845 ();
 sg13g2_fill_2 FILLER_3_1850 ();
 sg13g2_fill_1 FILLER_3_1857 ();
 sg13g2_fill_1 FILLER_3_1884 ();
 sg13g2_fill_1 FILLER_3_1898 ();
 sg13g2_fill_2 FILLER_3_1932 ();
 sg13g2_fill_2 FILLER_3_1959 ();
 sg13g2_fill_1 FILLER_3_2041 ();
 sg13g2_fill_2 FILLER_3_2051 ();
 sg13g2_fill_1 FILLER_3_2057 ();
 sg13g2_fill_1 FILLER_3_2088 ();
 sg13g2_fill_1 FILLER_3_2107 ();
 sg13g2_fill_1 FILLER_3_2137 ();
 sg13g2_decap_8 FILLER_3_2151 ();
 sg13g2_decap_8 FILLER_3_2158 ();
 sg13g2_decap_8 FILLER_3_2165 ();
 sg13g2_decap_8 FILLER_3_2172 ();
 sg13g2_decap_8 FILLER_3_2179 ();
 sg13g2_decap_8 FILLER_3_2186 ();
 sg13g2_decap_8 FILLER_3_2193 ();
 sg13g2_decap_8 FILLER_3_2200 ();
 sg13g2_decap_8 FILLER_3_2207 ();
 sg13g2_decap_8 FILLER_3_2214 ();
 sg13g2_decap_8 FILLER_3_2221 ();
 sg13g2_decap_8 FILLER_3_2228 ();
 sg13g2_decap_8 FILLER_3_2235 ();
 sg13g2_decap_8 FILLER_3_2242 ();
 sg13g2_decap_8 FILLER_3_2249 ();
 sg13g2_decap_4 FILLER_3_2256 ();
 sg13g2_decap_8 FILLER_3_2264 ();
 sg13g2_decap_8 FILLER_3_2271 ();
 sg13g2_fill_2 FILLER_3_2278 ();
 sg13g2_fill_2 FILLER_3_2283 ();
 sg13g2_decap_8 FILLER_3_2315 ();
 sg13g2_decap_8 FILLER_3_2322 ();
 sg13g2_fill_1 FILLER_3_2329 ();
 sg13g2_decap_4 FILLER_3_2340 ();
 sg13g2_fill_1 FILLER_3_2344 ();
 sg13g2_decap_4 FILLER_3_2376 ();
 sg13g2_fill_1 FILLER_3_2380 ();
 sg13g2_fill_1 FILLER_3_2386 ();
 sg13g2_decap_4 FILLER_3_2423 ();
 sg13g2_decap_8 FILLER_3_2435 ();
 sg13g2_decap_8 FILLER_3_2442 ();
 sg13g2_decap_8 FILLER_3_2449 ();
 sg13g2_fill_2 FILLER_3_2456 ();
 sg13g2_fill_2 FILLER_3_2471 ();
 sg13g2_fill_1 FILLER_3_2499 ();
 sg13g2_fill_1 FILLER_3_2504 ();
 sg13g2_fill_2 FILLER_3_2509 ();
 sg13g2_fill_1 FILLER_3_2524 ();
 sg13g2_decap_8 FILLER_3_2551 ();
 sg13g2_decap_8 FILLER_3_2558 ();
 sg13g2_decap_8 FILLER_3_2565 ();
 sg13g2_decap_8 FILLER_3_2572 ();
 sg13g2_decap_8 FILLER_3_2579 ();
 sg13g2_decap_8 FILLER_3_2586 ();
 sg13g2_decap_8 FILLER_3_2593 ();
 sg13g2_decap_8 FILLER_3_2600 ();
 sg13g2_decap_8 FILLER_3_2607 ();
 sg13g2_decap_8 FILLER_3_2614 ();
 sg13g2_decap_8 FILLER_3_2621 ();
 sg13g2_decap_8 FILLER_3_2628 ();
 sg13g2_decap_8 FILLER_3_2635 ();
 sg13g2_decap_8 FILLER_3_2642 ();
 sg13g2_decap_8 FILLER_3_2649 ();
 sg13g2_decap_8 FILLER_3_2656 ();
 sg13g2_decap_8 FILLER_3_2663 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_4 ();
 sg13g2_fill_2 FILLER_4_23 ();
 sg13g2_fill_1 FILLER_4_90 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_fill_2 FILLER_4_139 ();
 sg13g2_fill_1 FILLER_4_141 ();
 sg13g2_decap_4 FILLER_4_206 ();
 sg13g2_fill_1 FILLER_4_210 ();
 sg13g2_fill_1 FILLER_4_219 ();
 sg13g2_fill_1 FILLER_4_224 ();
 sg13g2_fill_2 FILLER_4_234 ();
 sg13g2_fill_1 FILLER_4_240 ();
 sg13g2_decap_4 FILLER_4_245 ();
 sg13g2_fill_1 FILLER_4_249 ();
 sg13g2_decap_4 FILLER_4_254 ();
 sg13g2_fill_2 FILLER_4_258 ();
 sg13g2_decap_4 FILLER_4_265 ();
 sg13g2_decap_4 FILLER_4_273 ();
 sg13g2_fill_2 FILLER_4_277 ();
 sg13g2_fill_2 FILLER_4_283 ();
 sg13g2_fill_1 FILLER_4_285 ();
 sg13g2_fill_1 FILLER_4_295 ();
 sg13g2_decap_4 FILLER_4_300 ();
 sg13g2_fill_2 FILLER_4_304 ();
 sg13g2_fill_1 FILLER_4_310 ();
 sg13g2_fill_1 FILLER_4_345 ();
 sg13g2_fill_1 FILLER_4_351 ();
 sg13g2_fill_2 FILLER_4_434 ();
 sg13g2_fill_1 FILLER_4_475 ();
 sg13g2_fill_2 FILLER_4_520 ();
 sg13g2_fill_1 FILLER_4_543 ();
 sg13g2_fill_1 FILLER_4_553 ();
 sg13g2_fill_1 FILLER_4_558 ();
 sg13g2_fill_2 FILLER_4_563 ();
 sg13g2_fill_1 FILLER_4_565 ();
 sg13g2_fill_1 FILLER_4_616 ();
 sg13g2_fill_1 FILLER_4_645 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_fill_2 FILLER_4_679 ();
 sg13g2_decap_4 FILLER_4_690 ();
 sg13g2_fill_1 FILLER_4_694 ();
 sg13g2_fill_1 FILLER_4_720 ();
 sg13g2_fill_2 FILLER_4_738 ();
 sg13g2_fill_1 FILLER_4_740 ();
 sg13g2_fill_1 FILLER_4_771 ();
 sg13g2_fill_1 FILLER_4_780 ();
 sg13g2_decap_8 FILLER_4_802 ();
 sg13g2_decap_8 FILLER_4_809 ();
 sg13g2_fill_2 FILLER_4_829 ();
 sg13g2_decap_4 FILLER_4_840 ();
 sg13g2_fill_1 FILLER_4_844 ();
 sg13g2_decap_8 FILLER_4_849 ();
 sg13g2_decap_8 FILLER_4_856 ();
 sg13g2_decap_4 FILLER_4_863 ();
 sg13g2_fill_1 FILLER_4_867 ();
 sg13g2_decap_8 FILLER_4_872 ();
 sg13g2_fill_2 FILLER_4_879 ();
 sg13g2_fill_1 FILLER_4_881 ();
 sg13g2_fill_1 FILLER_4_892 ();
 sg13g2_fill_2 FILLER_4_897 ();
 sg13g2_fill_1 FILLER_4_916 ();
 sg13g2_fill_1 FILLER_4_943 ();
 sg13g2_fill_1 FILLER_4_980 ();
 sg13g2_fill_1 FILLER_4_994 ();
 sg13g2_fill_2 FILLER_4_1021 ();
 sg13g2_fill_2 FILLER_4_1027 ();
 sg13g2_fill_2 FILLER_4_1072 ();
 sg13g2_fill_1 FILLER_4_1083 ();
 sg13g2_fill_1 FILLER_4_1101 ();
 sg13g2_fill_2 FILLER_4_1106 ();
 sg13g2_decap_8 FILLER_4_1112 ();
 sg13g2_fill_2 FILLER_4_1136 ();
 sg13g2_fill_1 FILLER_4_1138 ();
 sg13g2_decap_4 FILLER_4_1144 ();
 sg13g2_fill_1 FILLER_4_1148 ();
 sg13g2_fill_2 FILLER_4_1153 ();
 sg13g2_decap_8 FILLER_4_1176 ();
 sg13g2_decap_4 FILLER_4_1183 ();
 sg13g2_fill_2 FILLER_4_1187 ();
 sg13g2_fill_1 FILLER_4_1193 ();
 sg13g2_fill_2 FILLER_4_1267 ();
 sg13g2_fill_1 FILLER_4_1269 ();
 sg13g2_decap_4 FILLER_4_1304 ();
 sg13g2_fill_1 FILLER_4_1308 ();
 sg13g2_fill_1 FILLER_4_1322 ();
 sg13g2_fill_1 FILLER_4_1331 ();
 sg13g2_fill_1 FILLER_4_1341 ();
 sg13g2_decap_8 FILLER_4_1346 ();
 sg13g2_decap_4 FILLER_4_1353 ();
 sg13g2_fill_2 FILLER_4_1357 ();
 sg13g2_decap_8 FILLER_4_1372 ();
 sg13g2_decap_8 FILLER_4_1379 ();
 sg13g2_decap_4 FILLER_4_1386 ();
 sg13g2_fill_1 FILLER_4_1454 ();
 sg13g2_fill_1 FILLER_4_1460 ();
 sg13g2_fill_1 FILLER_4_1465 ();
 sg13g2_decap_8 FILLER_4_1500 ();
 sg13g2_fill_2 FILLER_4_1511 ();
 sg13g2_decap_4 FILLER_4_1534 ();
 sg13g2_fill_2 FILLER_4_1538 ();
 sg13g2_fill_1 FILLER_4_1562 ();
 sg13g2_fill_2 FILLER_4_1588 ();
 sg13g2_fill_1 FILLER_4_1616 ();
 sg13g2_fill_2 FILLER_4_1634 ();
 sg13g2_decap_4 FILLER_4_1640 ();
 sg13g2_fill_2 FILLER_4_1644 ();
 sg13g2_decap_8 FILLER_4_1650 ();
 sg13g2_decap_4 FILLER_4_1657 ();
 sg13g2_fill_1 FILLER_4_1665 ();
 sg13g2_decap_8 FILLER_4_1679 ();
 sg13g2_decap_8 FILLER_4_1712 ();
 sg13g2_decap_4 FILLER_4_1719 ();
 sg13g2_fill_1 FILLER_4_1732 ();
 sg13g2_fill_1 FILLER_4_1741 ();
 sg13g2_decap_8 FILLER_4_1777 ();
 sg13g2_decap_4 FILLER_4_1784 ();
 sg13g2_decap_8 FILLER_4_1792 ();
 sg13g2_decap_8 FILLER_4_1799 ();
 sg13g2_fill_1 FILLER_4_1806 ();
 sg13g2_fill_1 FILLER_4_1811 ();
 sg13g2_decap_8 FILLER_4_1820 ();
 sg13g2_decap_4 FILLER_4_1840 ();
 sg13g2_fill_1 FILLER_4_1844 ();
 sg13g2_decap_4 FILLER_4_1854 ();
 sg13g2_fill_1 FILLER_4_1858 ();
 sg13g2_fill_1 FILLER_4_1871 ();
 sg13g2_decap_8 FILLER_4_1876 ();
 sg13g2_decap_8 FILLER_4_1883 ();
 sg13g2_decap_8 FILLER_4_1890 ();
 sg13g2_decap_8 FILLER_4_1897 ();
 sg13g2_decap_8 FILLER_4_1904 ();
 sg13g2_fill_1 FILLER_4_1915 ();
 sg13g2_fill_2 FILLER_4_1921 ();
 sg13g2_fill_2 FILLER_4_1928 ();
 sg13g2_fill_2 FILLER_4_2007 ();
 sg13g2_fill_1 FILLER_4_2009 ();
 sg13g2_fill_2 FILLER_4_2027 ();
 sg13g2_fill_2 FILLER_4_2038 ();
 sg13g2_fill_1 FILLER_4_2083 ();
 sg13g2_fill_1 FILLER_4_2093 ();
 sg13g2_fill_1 FILLER_4_2099 ();
 sg13g2_fill_2 FILLER_4_2108 ();
 sg13g2_fill_2 FILLER_4_2132 ();
 sg13g2_decap_8 FILLER_4_2160 ();
 sg13g2_decap_8 FILLER_4_2167 ();
 sg13g2_decap_8 FILLER_4_2174 ();
 sg13g2_decap_8 FILLER_4_2181 ();
 sg13g2_decap_8 FILLER_4_2188 ();
 sg13g2_decap_8 FILLER_4_2195 ();
 sg13g2_decap_8 FILLER_4_2202 ();
 sg13g2_decap_8 FILLER_4_2209 ();
 sg13g2_fill_2 FILLER_4_2216 ();
 sg13g2_fill_2 FILLER_4_2222 ();
 sg13g2_decap_4 FILLER_4_2250 ();
 sg13g2_decap_8 FILLER_4_2313 ();
 sg13g2_fill_2 FILLER_4_2320 ();
 sg13g2_fill_1 FILLER_4_2322 ();
 sg13g2_decap_8 FILLER_4_2359 ();
 sg13g2_decap_4 FILLER_4_2366 ();
 sg13g2_fill_1 FILLER_4_2370 ();
 sg13g2_fill_1 FILLER_4_2402 ();
 sg13g2_decap_4 FILLER_4_2407 ();
 sg13g2_fill_2 FILLER_4_2411 ();
 sg13g2_decap_8 FILLER_4_2428 ();
 sg13g2_decap_8 FILLER_4_2435 ();
 sg13g2_decap_8 FILLER_4_2442 ();
 sg13g2_decap_8 FILLER_4_2449 ();
 sg13g2_decap_8 FILLER_4_2456 ();
 sg13g2_decap_4 FILLER_4_2463 ();
 sg13g2_fill_2 FILLER_4_2467 ();
 sg13g2_fill_2 FILLER_4_2479 ();
 sg13g2_fill_1 FILLER_4_2481 ();
 sg13g2_fill_2 FILLER_4_2508 ();
 sg13g2_fill_1 FILLER_4_2510 ();
 sg13g2_fill_1 FILLER_4_2516 ();
 sg13g2_fill_1 FILLER_4_2527 ();
 sg13g2_decap_4 FILLER_4_2549 ();
 sg13g2_fill_1 FILLER_4_2553 ();
 sg13g2_fill_2 FILLER_4_2563 ();
 sg13g2_decap_8 FILLER_4_2578 ();
 sg13g2_decap_4 FILLER_4_2585 ();
 sg13g2_decap_8 FILLER_4_2597 ();
 sg13g2_decap_8 FILLER_4_2604 ();
 sg13g2_decap_8 FILLER_4_2611 ();
 sg13g2_decap_8 FILLER_4_2618 ();
 sg13g2_decap_8 FILLER_4_2625 ();
 sg13g2_decap_8 FILLER_4_2632 ();
 sg13g2_decap_8 FILLER_4_2639 ();
 sg13g2_decap_8 FILLER_4_2646 ();
 sg13g2_decap_8 FILLER_4_2653 ();
 sg13g2_decap_8 FILLER_4_2660 ();
 sg13g2_fill_2 FILLER_4_2667 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_11 ();
 sg13g2_decap_4 FILLER_5_17 ();
 sg13g2_fill_2 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_31 ();
 sg13g2_fill_2 FILLER_5_38 ();
 sg13g2_fill_1 FILLER_5_40 ();
 sg13g2_decap_8 FILLER_5_75 ();
 sg13g2_fill_2 FILLER_5_82 ();
 sg13g2_decap_4 FILLER_5_89 ();
 sg13g2_fill_1 FILLER_5_93 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_4 FILLER_5_105 ();
 sg13g2_fill_2 FILLER_5_109 ();
 sg13g2_decap_4 FILLER_5_115 ();
 sg13g2_fill_2 FILLER_5_123 ();
 sg13g2_fill_2 FILLER_5_138 ();
 sg13g2_fill_1 FILLER_5_140 ();
 sg13g2_fill_2 FILLER_5_149 ();
 sg13g2_fill_1 FILLER_5_168 ();
 sg13g2_fill_2 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_188 ();
 sg13g2_fill_2 FILLER_5_198 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_205 ();
 sg13g2_fill_2 FILLER_5_212 ();
 sg13g2_fill_1 FILLER_5_214 ();
 sg13g2_fill_2 FILLER_5_241 ();
 sg13g2_fill_1 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_fill_1 FILLER_5_341 ();
 sg13g2_fill_2 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_5_456 ();
 sg13g2_fill_1 FILLER_5_462 ();
 sg13g2_fill_1 FILLER_5_472 ();
 sg13g2_fill_2 FILLER_5_503 ();
 sg13g2_fill_1 FILLER_5_505 ();
 sg13g2_decap_8 FILLER_5_510 ();
 sg13g2_decap_4 FILLER_5_517 ();
 sg13g2_fill_1 FILLER_5_521 ();
 sg13g2_decap_8 FILLER_5_543 ();
 sg13g2_decap_8 FILLER_5_550 ();
 sg13g2_fill_1 FILLER_5_557 ();
 sg13g2_fill_2 FILLER_5_571 ();
 sg13g2_fill_1 FILLER_5_573 ();
 sg13g2_fill_1 FILLER_5_637 ();
 sg13g2_fill_1 FILLER_5_647 ();
 sg13g2_fill_1 FILLER_5_652 ();
 sg13g2_decap_8 FILLER_5_660 ();
 sg13g2_decap_8 FILLER_5_667 ();
 sg13g2_decap_8 FILLER_5_674 ();
 sg13g2_decap_4 FILLER_5_689 ();
 sg13g2_fill_1 FILLER_5_693 ();
 sg13g2_decap_4 FILLER_5_698 ();
 sg13g2_fill_1 FILLER_5_702 ();
 sg13g2_fill_2 FILLER_5_716 ();
 sg13g2_fill_1 FILLER_5_718 ();
 sg13g2_fill_2 FILLER_5_732 ();
 sg13g2_fill_1 FILLER_5_734 ();
 sg13g2_fill_2 FILLER_5_739 ();
 sg13g2_fill_1 FILLER_5_741 ();
 sg13g2_decap_8 FILLER_5_750 ();
 sg13g2_fill_2 FILLER_5_769 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_835 ();
 sg13g2_decap_8 FILLER_5_842 ();
 sg13g2_fill_2 FILLER_5_849 ();
 sg13g2_fill_1 FILLER_5_851 ();
 sg13g2_decap_4 FILLER_5_877 ();
 sg13g2_fill_1 FILLER_5_881 ();
 sg13g2_decap_8 FILLER_5_895 ();
 sg13g2_decap_4 FILLER_5_902 ();
 sg13g2_fill_2 FILLER_5_906 ();
 sg13g2_decap_4 FILLER_5_930 ();
 sg13g2_fill_1 FILLER_5_934 ();
 sg13g2_decap_8 FILLER_5_939 ();
 sg13g2_decap_4 FILLER_5_946 ();
 sg13g2_fill_1 FILLER_5_950 ();
 sg13g2_decap_8 FILLER_5_1068 ();
 sg13g2_fill_1 FILLER_5_1075 ();
 sg13g2_fill_1 FILLER_5_1080 ();
 sg13g2_fill_1 FILLER_5_1089 ();
 sg13g2_fill_2 FILLER_5_1095 ();
 sg13g2_decap_4 FILLER_5_1101 ();
 sg13g2_fill_2 FILLER_5_1105 ();
 sg13g2_decap_4 FILLER_5_1111 ();
 sg13g2_fill_2 FILLER_5_1119 ();
 sg13g2_decap_8 FILLER_5_1125 ();
 sg13g2_fill_2 FILLER_5_1132 ();
 sg13g2_decap_8 FILLER_5_1172 ();
 sg13g2_fill_1 FILLER_5_1179 ();
 sg13g2_fill_1 FILLER_5_1223 ();
 sg13g2_fill_2 FILLER_5_1229 ();
 sg13g2_fill_1 FILLER_5_1231 ();
 sg13g2_fill_1 FILLER_5_1236 ();
 sg13g2_fill_2 FILLER_5_1250 ();
 sg13g2_decap_8 FILLER_5_1256 ();
 sg13g2_fill_2 FILLER_5_1263 ();
 sg13g2_fill_1 FILLER_5_1265 ();
 sg13g2_fill_2 FILLER_5_1270 ();
 sg13g2_decap_8 FILLER_5_1293 ();
 sg13g2_decap_8 FILLER_5_1300 ();
 sg13g2_decap_4 FILLER_5_1307 ();
 sg13g2_decap_4 FILLER_5_1315 ();
 sg13g2_fill_2 FILLER_5_1324 ();
 sg13g2_fill_2 FILLER_5_1356 ();
 sg13g2_fill_1 FILLER_5_1358 ();
 sg13g2_fill_2 FILLER_5_1367 ();
 sg13g2_fill_1 FILLER_5_1369 ();
 sg13g2_decap_8 FILLER_5_1374 ();
 sg13g2_decap_8 FILLER_5_1381 ();
 sg13g2_decap_8 FILLER_5_1388 ();
 sg13g2_fill_2 FILLER_5_1395 ();
 sg13g2_fill_1 FILLER_5_1397 ();
 sg13g2_fill_2 FILLER_5_1406 ();
 sg13g2_decap_8 FILLER_5_1447 ();
 sg13g2_decap_8 FILLER_5_1454 ();
 sg13g2_fill_2 FILLER_5_1491 ();
 sg13g2_fill_1 FILLER_5_1493 ();
 sg13g2_decap_4 FILLER_5_1502 ();
 sg13g2_fill_1 FILLER_5_1506 ();
 sg13g2_decap_8 FILLER_5_1533 ();
 sg13g2_fill_1 FILLER_5_1574 ();
 sg13g2_fill_2 FILLER_5_1596 ();
 sg13g2_fill_1 FILLER_5_1602 ();
 sg13g2_fill_2 FILLER_5_1615 ();
 sg13g2_decap_8 FILLER_5_1652 ();
 sg13g2_fill_2 FILLER_5_1664 ();
 sg13g2_fill_1 FILLER_5_1666 ();
 sg13g2_fill_1 FILLER_5_1675 ();
 sg13g2_fill_2 FILLER_5_1681 ();
 sg13g2_fill_1 FILLER_5_1683 ();
 sg13g2_decap_8 FILLER_5_1710 ();
 sg13g2_fill_1 FILLER_5_1717 ();
 sg13g2_fill_2 FILLER_5_1783 ();
 sg13g2_fill_2 FILLER_5_1789 ();
 sg13g2_fill_1 FILLER_5_1791 ();
 sg13g2_fill_2 FILLER_5_1797 ();
 sg13g2_fill_1 FILLER_5_1799 ();
 sg13g2_fill_2 FILLER_5_1804 ();
 sg13g2_fill_1 FILLER_5_1806 ();
 sg13g2_fill_2 FILLER_5_1817 ();
 sg13g2_decap_4 FILLER_5_1827 ();
 sg13g2_fill_1 FILLER_5_1831 ();
 sg13g2_fill_1 FILLER_5_1840 ();
 sg13g2_fill_1 FILLER_5_1850 ();
 sg13g2_fill_2 FILLER_5_1895 ();
 sg13g2_fill_1 FILLER_5_1901 ();
 sg13g2_fill_1 FILLER_5_1906 ();
 sg13g2_fill_1 FILLER_5_1911 ();
 sg13g2_fill_1 FILLER_5_1921 ();
 sg13g2_fill_2 FILLER_5_1926 ();
 sg13g2_fill_2 FILLER_5_1932 ();
 sg13g2_fill_2 FILLER_5_1944 ();
 sg13g2_fill_2 FILLER_5_1950 ();
 sg13g2_fill_1 FILLER_5_1973 ();
 sg13g2_fill_1 FILLER_5_2000 ();
 sg13g2_decap_8 FILLER_5_2012 ();
 sg13g2_decap_8 FILLER_5_2019 ();
 sg13g2_fill_2 FILLER_5_2026 ();
 sg13g2_fill_1 FILLER_5_2028 ();
 sg13g2_fill_1 FILLER_5_2055 ();
 sg13g2_fill_2 FILLER_5_2087 ();
 sg13g2_fill_1 FILLER_5_2089 ();
 sg13g2_fill_1 FILLER_5_2121 ();
 sg13g2_decap_8 FILLER_5_2168 ();
 sg13g2_decap_8 FILLER_5_2175 ();
 sg13g2_decap_8 FILLER_5_2182 ();
 sg13g2_decap_8 FILLER_5_2189 ();
 sg13g2_decap_8 FILLER_5_2196 ();
 sg13g2_decap_8 FILLER_5_2203 ();
 sg13g2_decap_4 FILLER_5_2210 ();
 sg13g2_fill_1 FILLER_5_2214 ();
 sg13g2_fill_2 FILLER_5_2254 ();
 sg13g2_fill_1 FILLER_5_2256 ();
 sg13g2_decap_8 FILLER_5_2262 ();
 sg13g2_fill_2 FILLER_5_2269 ();
 sg13g2_fill_1 FILLER_5_2271 ();
 sg13g2_decap_8 FILLER_5_2302 ();
 sg13g2_fill_1 FILLER_5_2309 ();
 sg13g2_decap_8 FILLER_5_2343 ();
 sg13g2_decap_4 FILLER_5_2350 ();
 sg13g2_fill_2 FILLER_5_2354 ();
 sg13g2_fill_1 FILLER_5_2361 ();
 sg13g2_fill_1 FILLER_5_2366 ();
 sg13g2_fill_1 FILLER_5_2377 ();
 sg13g2_fill_2 FILLER_5_2393 ();
 sg13g2_fill_1 FILLER_5_2402 ();
 sg13g2_fill_1 FILLER_5_2407 ();
 sg13g2_fill_1 FILLER_5_2411 ();
 sg13g2_fill_1 FILLER_5_2453 ();
 sg13g2_decap_8 FILLER_5_2457 ();
 sg13g2_decap_8 FILLER_5_2464 ();
 sg13g2_fill_1 FILLER_5_2471 ();
 sg13g2_decap_8 FILLER_5_2502 ();
 sg13g2_fill_1 FILLER_5_2509 ();
 sg13g2_decap_4 FILLER_5_2535 ();
 sg13g2_fill_1 FILLER_5_2539 ();
 sg13g2_fill_1 FILLER_5_2575 ();
 sg13g2_decap_8 FILLER_5_2607 ();
 sg13g2_decap_4 FILLER_5_2614 ();
 sg13g2_fill_2 FILLER_5_2618 ();
 sg13g2_decap_8 FILLER_5_2633 ();
 sg13g2_decap_8 FILLER_5_2640 ();
 sg13g2_decap_8 FILLER_5_2647 ();
 sg13g2_decap_8 FILLER_5_2654 ();
 sg13g2_decap_8 FILLER_5_2661 ();
 sg13g2_fill_2 FILLER_5_2668 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_13 ();
 sg13g2_fill_1 FILLER_6_17 ();
 sg13g2_decap_8 FILLER_6_27 ();
 sg13g2_decap_8 FILLER_6_34 ();
 sg13g2_fill_2 FILLER_6_85 ();
 sg13g2_decap_8 FILLER_6_113 ();
 sg13g2_decap_8 FILLER_6_120 ();
 sg13g2_decap_4 FILLER_6_127 ();
 sg13g2_fill_1 FILLER_6_148 ();
 sg13g2_fill_2 FILLER_6_158 ();
 sg13g2_fill_2 FILLER_6_173 ();
 sg13g2_fill_2 FILLER_6_209 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_fill_2 FILLER_6_226 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_fill_2 FILLER_6_261 ();
 sg13g2_fill_2 FILLER_6_268 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_fill_2 FILLER_6_297 ();
 sg13g2_decap_8 FILLER_6_303 ();
 sg13g2_fill_2 FILLER_6_310 ();
 sg13g2_fill_1 FILLER_6_312 ();
 sg13g2_fill_2 FILLER_6_330 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_fill_1 FILLER_6_369 ();
 sg13g2_fill_1 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_456 ();
 sg13g2_fill_1 FILLER_6_468 ();
 sg13g2_fill_2 FILLER_6_489 ();
 sg13g2_fill_1 FILLER_6_495 ();
 sg13g2_fill_1 FILLER_6_505 ();
 sg13g2_decap_8 FILLER_6_510 ();
 sg13g2_fill_2 FILLER_6_526 ();
 sg13g2_decap_8 FILLER_6_537 ();
 sg13g2_decap_4 FILLER_6_544 ();
 sg13g2_fill_2 FILLER_6_548 ();
 sg13g2_fill_2 FILLER_6_598 ();
 sg13g2_fill_2 FILLER_6_604 ();
 sg13g2_fill_2 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_fill_2 FILLER_6_669 ();
 sg13g2_fill_2 FILLER_6_728 ();
 sg13g2_decap_4 FILLER_6_748 ();
 sg13g2_fill_1 FILLER_6_752 ();
 sg13g2_fill_2 FILLER_6_766 ();
 sg13g2_fill_2 FILLER_6_798 ();
 sg13g2_fill_1 FILLER_6_809 ();
 sg13g2_fill_1 FILLER_6_814 ();
 sg13g2_fill_1 FILLER_6_819 ();
 sg13g2_fill_2 FILLER_6_846 ();
 sg13g2_fill_2 FILLER_6_874 ();
 sg13g2_fill_2 FILLER_6_902 ();
 sg13g2_decap_8 FILLER_6_908 ();
 sg13g2_fill_2 FILLER_6_915 ();
 sg13g2_fill_1 FILLER_6_917 ();
 sg13g2_decap_8 FILLER_6_922 ();
 sg13g2_decap_8 FILLER_6_929 ();
 sg13g2_decap_8 FILLER_6_936 ();
 sg13g2_fill_2 FILLER_6_943 ();
 sg13g2_fill_1 FILLER_6_945 ();
 sg13g2_fill_1 FILLER_6_962 ();
 sg13g2_fill_2 FILLER_6_972 ();
 sg13g2_fill_2 FILLER_6_982 ();
 sg13g2_fill_2 FILLER_6_988 ();
 sg13g2_fill_2 FILLER_6_1063 ();
 sg13g2_fill_2 FILLER_6_1083 ();
 sg13g2_fill_2 FILLER_6_1089 ();
 sg13g2_fill_1 FILLER_6_1122 ();
 sg13g2_decap_8 FILLER_6_1184 ();
 sg13g2_decap_8 FILLER_6_1191 ();
 sg13g2_decap_4 FILLER_6_1198 ();
 sg13g2_fill_2 FILLER_6_1249 ();
 sg13g2_fill_1 FILLER_6_1251 ();
 sg13g2_decap_8 FILLER_6_1256 ();
 sg13g2_decap_8 FILLER_6_1263 ();
 sg13g2_fill_2 FILLER_6_1270 ();
 sg13g2_decap_8 FILLER_6_1276 ();
 sg13g2_fill_2 FILLER_6_1283 ();
 sg13g2_fill_1 FILLER_6_1285 ();
 sg13g2_fill_2 FILLER_6_1320 ();
 sg13g2_fill_1 FILLER_6_1322 ();
 sg13g2_decap_8 FILLER_6_1331 ();
 sg13g2_fill_2 FILLER_6_1338 ();
 sg13g2_fill_1 FILLER_6_1340 ();
 sg13g2_fill_2 FILLER_6_1346 ();
 sg13g2_fill_1 FILLER_6_1352 ();
 sg13g2_fill_2 FILLER_6_1357 ();
 sg13g2_decap_8 FILLER_6_1385 ();
 sg13g2_decap_4 FILLER_6_1392 ();
 sg13g2_fill_2 FILLER_6_1396 ();
 sg13g2_decap_8 FILLER_6_1403 ();
 sg13g2_decap_8 FILLER_6_1414 ();
 sg13g2_fill_1 FILLER_6_1421 ();
 sg13g2_fill_2 FILLER_6_1427 ();
 sg13g2_fill_2 FILLER_6_1442 ();
 sg13g2_decap_8 FILLER_6_1448 ();
 sg13g2_fill_2 FILLER_6_1455 ();
 sg13g2_decap_4 FILLER_6_1466 ();
 sg13g2_fill_1 FILLER_6_1470 ();
 sg13g2_fill_1 FILLER_6_1480 ();
 sg13g2_fill_2 FILLER_6_1489 ();
 sg13g2_fill_1 FILLER_6_1491 ();
 sg13g2_decap_8 FILLER_6_1531 ();
 sg13g2_decap_4 FILLER_6_1552 ();
 sg13g2_decap_4 FILLER_6_1616 ();
 sg13g2_fill_1 FILLER_6_1620 ();
 sg13g2_fill_2 FILLER_6_1626 ();
 sg13g2_fill_1 FILLER_6_1658 ();
 sg13g2_fill_2 FILLER_6_1676 ();
 sg13g2_fill_1 FILLER_6_1678 ();
 sg13g2_fill_1 FILLER_6_1684 ();
 sg13g2_decap_8 FILLER_6_1706 ();
 sg13g2_decap_4 FILLER_6_1713 ();
 sg13g2_fill_1 FILLER_6_1717 ();
 sg13g2_fill_2 FILLER_6_1749 ();
 sg13g2_fill_1 FILLER_6_1751 ();
 sg13g2_fill_1 FILLER_6_1791 ();
 sg13g2_fill_2 FILLER_6_1796 ();
 sg13g2_fill_1 FILLER_6_1798 ();
 sg13g2_fill_2 FILLER_6_1916 ();
 sg13g2_fill_1 FILLER_6_1987 ();
 sg13g2_fill_1 FILLER_6_2014 ();
 sg13g2_fill_2 FILLER_6_2024 ();
 sg13g2_fill_1 FILLER_6_2037 ();
 sg13g2_decap_8 FILLER_6_2055 ();
 sg13g2_decap_4 FILLER_6_2062 ();
 sg13g2_fill_1 FILLER_6_2074 ();
 sg13g2_decap_4 FILLER_6_2084 ();
 sg13g2_fill_2 FILLER_6_2101 ();
 sg13g2_decap_4 FILLER_6_2132 ();
 sg13g2_decap_8 FILLER_6_2162 ();
 sg13g2_decap_8 FILLER_6_2169 ();
 sg13g2_decap_8 FILLER_6_2176 ();
 sg13g2_decap_8 FILLER_6_2183 ();
 sg13g2_decap_8 FILLER_6_2190 ();
 sg13g2_decap_8 FILLER_6_2197 ();
 sg13g2_decap_8 FILLER_6_2204 ();
 sg13g2_decap_8 FILLER_6_2211 ();
 sg13g2_fill_2 FILLER_6_2218 ();
 sg13g2_fill_1 FILLER_6_2220 ();
 sg13g2_decap_8 FILLER_6_2239 ();
 sg13g2_decap_4 FILLER_6_2246 ();
 sg13g2_fill_1 FILLER_6_2250 ();
 sg13g2_fill_2 FILLER_6_2281 ();
 sg13g2_fill_1 FILLER_6_2283 ();
 sg13g2_decap_4 FILLER_6_2321 ();
 sg13g2_fill_1 FILLER_6_2343 ();
 sg13g2_decap_4 FILLER_6_2352 ();
 sg13g2_fill_2 FILLER_6_2356 ();
 sg13g2_fill_1 FILLER_6_2366 ();
 sg13g2_fill_2 FILLER_6_2381 ();
 sg13g2_fill_1 FILLER_6_2383 ();
 sg13g2_fill_2 FILLER_6_2392 ();
 sg13g2_fill_2 FILLER_6_2433 ();
 sg13g2_fill_2 FILLER_6_2439 ();
 sg13g2_fill_1 FILLER_6_2441 ();
 sg13g2_fill_2 FILLER_6_2459 ();
 sg13g2_fill_1 FILLER_6_2461 ();
 sg13g2_decap_4 FILLER_6_2483 ();
 sg13g2_fill_2 FILLER_6_2487 ();
 sg13g2_decap_8 FILLER_6_2497 ();
 sg13g2_decap_4 FILLER_6_2512 ();
 sg13g2_fill_1 FILLER_6_2516 ();
 sg13g2_fill_2 FILLER_6_2609 ();
 sg13g2_decap_8 FILLER_6_2624 ();
 sg13g2_decap_8 FILLER_6_2631 ();
 sg13g2_decap_8 FILLER_6_2638 ();
 sg13g2_decap_8 FILLER_6_2645 ();
 sg13g2_decap_8 FILLER_6_2652 ();
 sg13g2_decap_8 FILLER_6_2659 ();
 sg13g2_decap_4 FILLER_6_2666 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_28 ();
 sg13g2_fill_1 FILLER_7_34 ();
 sg13g2_fill_1 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_66 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_decap_8 FILLER_7_94 ();
 sg13g2_fill_1 FILLER_7_101 ();
 sg13g2_decap_8 FILLER_7_110 ();
 sg13g2_decap_4 FILLER_7_117 ();
 sg13g2_fill_2 FILLER_7_121 ();
 sg13g2_fill_1 FILLER_7_132 ();
 sg13g2_fill_1 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_178 ();
 sg13g2_fill_2 FILLER_7_185 ();
 sg13g2_fill_1 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_227 ();
 sg13g2_fill_1 FILLER_7_233 ();
 sg13g2_fill_1 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_fill_1 FILLER_7_250 ();
 sg13g2_fill_1 FILLER_7_290 ();
 sg13g2_fill_2 FILLER_7_304 ();
 sg13g2_decap_4 FILLER_7_310 ();
 sg13g2_fill_2 FILLER_7_314 ();
 sg13g2_fill_1 FILLER_7_320 ();
 sg13g2_fill_1 FILLER_7_335 ();
 sg13g2_fill_1 FILLER_7_358 ();
 sg13g2_fill_2 FILLER_7_395 ();
 sg13g2_fill_1 FILLER_7_407 ();
 sg13g2_fill_2 FILLER_7_417 ();
 sg13g2_fill_1 FILLER_7_463 ();
 sg13g2_fill_2 FILLER_7_527 ();
 sg13g2_decap_4 FILLER_7_555 ();
 sg13g2_fill_2 FILLER_7_595 ();
 sg13g2_fill_2 FILLER_7_623 ();
 sg13g2_fill_1 FILLER_7_635 ();
 sg13g2_fill_2 FILLER_7_666 ();
 sg13g2_fill_2 FILLER_7_759 ();
 sg13g2_fill_1 FILLER_7_761 ();
 sg13g2_decap_8 FILLER_7_783 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_4 FILLER_7_831 ();
 sg13g2_fill_2 FILLER_7_835 ();
 sg13g2_fill_2 FILLER_7_887 ();
 sg13g2_fill_1 FILLER_7_900 ();
 sg13g2_fill_1 FILLER_7_905 ();
 sg13g2_decap_4 FILLER_7_941 ();
 sg13g2_fill_1 FILLER_7_945 ();
 sg13g2_fill_2 FILLER_7_956 ();
 sg13g2_fill_2 FILLER_7_991 ();
 sg13g2_fill_1 FILLER_7_997 ();
 sg13g2_fill_2 FILLER_7_1008 ();
 sg13g2_fill_2 FILLER_7_1018 ();
 sg13g2_fill_1 FILLER_7_1051 ();
 sg13g2_fill_2 FILLER_7_1069 ();
 sg13g2_fill_2 FILLER_7_1101 ();
 sg13g2_fill_2 FILLER_7_1147 ();
 sg13g2_fill_1 FILLER_7_1153 ();
 sg13g2_fill_1 FILLER_7_1159 ();
 sg13g2_fill_2 FILLER_7_1181 ();
 sg13g2_fill_1 FILLER_7_1183 ();
 sg13g2_fill_1 FILLER_7_1210 ();
 sg13g2_fill_2 FILLER_7_1264 ();
 sg13g2_fill_1 FILLER_7_1266 ();
 sg13g2_fill_1 FILLER_7_1272 ();
 sg13g2_fill_1 FILLER_7_1395 ();
 sg13g2_fill_1 FILLER_7_1400 ();
 sg13g2_decap_8 FILLER_7_1436 ();
 sg13g2_fill_2 FILLER_7_1443 ();
 sg13g2_fill_1 FILLER_7_1479 ();
 sg13g2_fill_2 FILLER_7_1498 ();
 sg13g2_fill_1 FILLER_7_1500 ();
 sg13g2_decap_8 FILLER_7_1518 ();
 sg13g2_decap_8 FILLER_7_1525 ();
 sg13g2_fill_1 FILLER_7_1532 ();
 sg13g2_fill_1 FILLER_7_1543 ();
 sg13g2_decap_4 FILLER_7_1557 ();
 sg13g2_fill_1 FILLER_7_1561 ();
 sg13g2_fill_1 FILLER_7_1575 ();
 sg13g2_fill_2 FILLER_7_1581 ();
 sg13g2_fill_1 FILLER_7_1592 ();
 sg13g2_fill_2 FILLER_7_1598 ();
 sg13g2_decap_8 FILLER_7_1609 ();
 sg13g2_fill_2 FILLER_7_1616 ();
 sg13g2_fill_1 FILLER_7_1618 ();
 sg13g2_fill_1 FILLER_7_1683 ();
 sg13g2_decap_8 FILLER_7_1710 ();
 sg13g2_fill_2 FILLER_7_1717 ();
 sg13g2_fill_1 FILLER_7_1732 ();
 sg13g2_fill_2 FILLER_7_1750 ();
 sg13g2_fill_2 FILLER_7_1778 ();
 sg13g2_fill_2 FILLER_7_1862 ();
 sg13g2_fill_2 FILLER_7_1911 ();
 sg13g2_fill_1 FILLER_7_1913 ();
 sg13g2_fill_1 FILLER_7_1940 ();
 sg13g2_fill_2 FILLER_7_1946 ();
 sg13g2_fill_1 FILLER_7_1977 ();
 sg13g2_decap_8 FILLER_7_2062 ();
 sg13g2_decap_8 FILLER_7_2069 ();
 sg13g2_fill_1 FILLER_7_2106 ();
 sg13g2_fill_2 FILLER_7_2128 ();
 sg13g2_fill_1 FILLER_7_2130 ();
 sg13g2_decap_8 FILLER_7_2157 ();
 sg13g2_decap_8 FILLER_7_2164 ();
 sg13g2_decap_8 FILLER_7_2171 ();
 sg13g2_decap_8 FILLER_7_2178 ();
 sg13g2_decap_8 FILLER_7_2185 ();
 sg13g2_decap_4 FILLER_7_2192 ();
 sg13g2_fill_1 FILLER_7_2196 ();
 sg13g2_decap_4 FILLER_7_2201 ();
 sg13g2_decap_4 FILLER_7_2209 ();
 sg13g2_fill_2 FILLER_7_2213 ();
 sg13g2_decap_8 FILLER_7_2241 ();
 sg13g2_decap_8 FILLER_7_2248 ();
 sg13g2_decap_8 FILLER_7_2255 ();
 sg13g2_decap_8 FILLER_7_2262 ();
 sg13g2_decap_4 FILLER_7_2269 ();
 sg13g2_fill_2 FILLER_7_2286 ();
 sg13g2_fill_1 FILLER_7_2288 ();
 sg13g2_decap_4 FILLER_7_2299 ();
 sg13g2_decap_8 FILLER_7_2351 ();
 sg13g2_fill_1 FILLER_7_2358 ();
 sg13g2_fill_2 FILLER_7_2369 ();
 sg13g2_decap_4 FILLER_7_2381 ();
 sg13g2_decap_4 FILLER_7_2405 ();
 sg13g2_fill_2 FILLER_7_2409 ();
 sg13g2_fill_1 FILLER_7_2441 ();
 sg13g2_fill_2 FILLER_7_2450 ();
 sg13g2_fill_1 FILLER_7_2452 ();
 sg13g2_decap_8 FILLER_7_2499 ();
 sg13g2_fill_2 FILLER_7_2536 ();
 sg13g2_decap_4 FILLER_7_2542 ();
 sg13g2_fill_1 FILLER_7_2546 ();
 sg13g2_fill_1 FILLER_7_2617 ();
 sg13g2_decap_4 FILLER_7_2622 ();
 sg13g2_fill_2 FILLER_7_2626 ();
 sg13g2_decap_8 FILLER_7_2636 ();
 sg13g2_decap_8 FILLER_7_2643 ();
 sg13g2_decap_8 FILLER_7_2650 ();
 sg13g2_decap_8 FILLER_7_2657 ();
 sg13g2_decap_4 FILLER_7_2664 ();
 sg13g2_fill_2 FILLER_7_2668 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_87 ();
 sg13g2_fill_1 FILLER_8_93 ();
 sg13g2_fill_1 FILLER_8_99 ();
 sg13g2_fill_2 FILLER_8_126 ();
 sg13g2_fill_1 FILLER_8_128 ();
 sg13g2_fill_2 FILLER_8_197 ();
 sg13g2_decap_4 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_229 ();
 sg13g2_decap_8 FILLER_8_236 ();
 sg13g2_decap_8 FILLER_8_243 ();
 sg13g2_decap_8 FILLER_8_250 ();
 sg13g2_fill_2 FILLER_8_257 ();
 sg13g2_fill_2 FILLER_8_311 ();
 sg13g2_fill_1 FILLER_8_313 ();
 sg13g2_fill_2 FILLER_8_319 ();
 sg13g2_fill_2 FILLER_8_380 ();
 sg13g2_fill_2 FILLER_8_392 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_2 FILLER_8_414 ();
 sg13g2_fill_1 FILLER_8_420 ();
 sg13g2_fill_1 FILLER_8_436 ();
 sg13g2_fill_1 FILLER_8_462 ();
 sg13g2_fill_2 FILLER_8_468 ();
 sg13g2_fill_1 FILLER_8_474 ();
 sg13g2_fill_1 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_519 ();
 sg13g2_fill_1 FILLER_8_526 ();
 sg13g2_fill_1 FILLER_8_536 ();
 sg13g2_fill_1 FILLER_8_558 ();
 sg13g2_fill_1 FILLER_8_563 ();
 sg13g2_fill_2 FILLER_8_598 ();
 sg13g2_fill_1 FILLER_8_626 ();
 sg13g2_fill_1 FILLER_8_633 ();
 sg13g2_fill_1 FILLER_8_637 ();
 sg13g2_fill_2 FILLER_8_731 ();
 sg13g2_fill_2 FILLER_8_804 ();
 sg13g2_fill_2 FILLER_8_841 ();
 sg13g2_fill_2 FILLER_8_852 ();
 sg13g2_fill_1 FILLER_8_871 ();
 sg13g2_fill_2 FILLER_8_897 ();
 sg13g2_fill_1 FILLER_8_903 ();
 sg13g2_fill_2 FILLER_8_943 ();
 sg13g2_fill_2 FILLER_8_971 ();
 sg13g2_fill_2 FILLER_8_1003 ();
 sg13g2_fill_2 FILLER_8_1012 ();
 sg13g2_fill_1 FILLER_8_1026 ();
 sg13g2_fill_2 FILLER_8_1101 ();
 sg13g2_fill_2 FILLER_8_1124 ();
 sg13g2_decap_8 FILLER_8_1138 ();
 sg13g2_decap_8 FILLER_8_1145 ();
 sg13g2_decap_8 FILLER_8_1152 ();
 sg13g2_decap_4 FILLER_8_1159 ();
 sg13g2_fill_2 FILLER_8_1163 ();
 sg13g2_decap_8 FILLER_8_1173 ();
 sg13g2_decap_4 FILLER_8_1180 ();
 sg13g2_fill_1 FILLER_8_1210 ();
 sg13g2_fill_1 FILLER_8_1215 ();
 sg13g2_fill_1 FILLER_8_1221 ();
 sg13g2_fill_1 FILLER_8_1252 ();
 sg13g2_fill_1 FILLER_8_1262 ();
 sg13g2_fill_2 FILLER_8_1328 ();
 sg13g2_decap_4 FILLER_8_1335 ();
 sg13g2_fill_2 FILLER_8_1343 ();
 sg13g2_fill_2 FILLER_8_1349 ();
 sg13g2_fill_2 FILLER_8_1399 ();
 sg13g2_fill_1 FILLER_8_1410 ();
 sg13g2_decap_8 FILLER_8_1437 ();
 sg13g2_decap_4 FILLER_8_1444 ();
 sg13g2_fill_1 FILLER_8_1448 ();
 sg13g2_decap_8 FILLER_8_1510 ();
 sg13g2_decap_8 FILLER_8_1517 ();
 sg13g2_fill_2 FILLER_8_1524 ();
 sg13g2_fill_2 FILLER_8_1536 ();
 sg13g2_fill_2 FILLER_8_1569 ();
 sg13g2_decap_4 FILLER_8_1604 ();
 sg13g2_fill_1 FILLER_8_1641 ();
 sg13g2_fill_1 FILLER_8_1667 ();
 sg13g2_decap_8 FILLER_8_1703 ();
 sg13g2_fill_2 FILLER_8_1710 ();
 sg13g2_fill_1 FILLER_8_1715 ();
 sg13g2_fill_2 FILLER_8_1719 ();
 sg13g2_decap_8 FILLER_8_1753 ();
 sg13g2_fill_2 FILLER_8_1769 ();
 sg13g2_fill_1 FILLER_8_1771 ();
 sg13g2_decap_8 FILLER_8_1776 ();
 sg13g2_decap_4 FILLER_8_1783 ();
 sg13g2_decap_8 FILLER_8_1791 ();
 sg13g2_fill_2 FILLER_8_1798 ();
 sg13g2_fill_1 FILLER_8_1855 ();
 sg13g2_fill_1 FILLER_8_1861 ();
 sg13g2_fill_1 FILLER_8_1888 ();
 sg13g2_fill_1 FILLER_8_1894 ();
 sg13g2_fill_2 FILLER_8_1899 ();
 sg13g2_fill_1 FILLER_8_1922 ();
 sg13g2_fill_2 FILLER_8_1928 ();
 sg13g2_fill_1 FILLER_8_1973 ();
 sg13g2_fill_1 FILLER_8_1977 ();
 sg13g2_fill_1 FILLER_8_1981 ();
 sg13g2_fill_2 FILLER_8_2071 ();
 sg13g2_fill_2 FILLER_8_2095 ();
 sg13g2_fill_1 FILLER_8_2127 ();
 sg13g2_decap_4 FILLER_8_2133 ();
 sg13g2_fill_2 FILLER_8_2141 ();
 sg13g2_decap_8 FILLER_8_2147 ();
 sg13g2_decap_8 FILLER_8_2154 ();
 sg13g2_decap_8 FILLER_8_2161 ();
 sg13g2_decap_8 FILLER_8_2168 ();
 sg13g2_decap_8 FILLER_8_2175 ();
 sg13g2_decap_8 FILLER_8_2182 ();
 sg13g2_fill_1 FILLER_8_2189 ();
 sg13g2_decap_4 FILLER_8_2216 ();
 sg13g2_fill_1 FILLER_8_2220 ();
 sg13g2_decap_4 FILLER_8_2225 ();
 sg13g2_fill_2 FILLER_8_2229 ();
 sg13g2_fill_2 FILLER_8_2261 ();
 sg13g2_fill_1 FILLER_8_2263 ();
 sg13g2_decap_4 FILLER_8_2269 ();
 sg13g2_fill_1 FILLER_8_2273 ();
 sg13g2_decap_8 FILLER_8_2300 ();
 sg13g2_fill_2 FILLER_8_2307 ();
 sg13g2_fill_1 FILLER_8_2332 ();
 sg13g2_fill_1 FILLER_8_2345 ();
 sg13g2_fill_1 FILLER_8_2360 ();
 sg13g2_fill_2 FILLER_8_2392 ();
 sg13g2_decap_8 FILLER_8_2399 ();
 sg13g2_decap_4 FILLER_8_2406 ();
 sg13g2_fill_2 FILLER_8_2415 ();
 sg13g2_fill_1 FILLER_8_2422 ();
 sg13g2_decap_8 FILLER_8_2432 ();
 sg13g2_fill_1 FILLER_8_2439 ();
 sg13g2_fill_2 FILLER_8_2461 ();
 sg13g2_fill_1 FILLER_8_2467 ();
 sg13g2_fill_1 FILLER_8_2494 ();
 sg13g2_fill_2 FILLER_8_2515 ();
 sg13g2_fill_2 FILLER_8_2521 ();
 sg13g2_fill_1 FILLER_8_2533 ();
 sg13g2_fill_2 FILLER_8_2626 ();
 sg13g2_decap_8 FILLER_8_2641 ();
 sg13g2_decap_8 FILLER_8_2648 ();
 sg13g2_decap_8 FILLER_8_2655 ();
 sg13g2_decap_8 FILLER_8_2662 ();
 sg13g2_fill_1 FILLER_8_2669 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_32 ();
 sg13g2_fill_2 FILLER_9_52 ();
 sg13g2_fill_1 FILLER_9_54 ();
 sg13g2_fill_2 FILLER_9_59 ();
 sg13g2_fill_2 FILLER_9_74 ();
 sg13g2_fill_1 FILLER_9_76 ();
 sg13g2_fill_1 FILLER_9_89 ();
 sg13g2_fill_2 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_169 ();
 sg13g2_fill_1 FILLER_9_212 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_250 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_fill_1 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_305 ();
 sg13g2_fill_1 FILLER_9_345 ();
 sg13g2_fill_2 FILLER_9_379 ();
 sg13g2_fill_1 FILLER_9_418 ();
 sg13g2_fill_2 FILLER_9_423 ();
 sg13g2_fill_1 FILLER_9_446 ();
 sg13g2_fill_2 FILLER_9_454 ();
 sg13g2_fill_2 FILLER_9_489 ();
 sg13g2_fill_1 FILLER_9_495 ();
 sg13g2_fill_2 FILLER_9_586 ();
 sg13g2_fill_1 FILLER_9_596 ();
 sg13g2_fill_2 FILLER_9_610 ();
 sg13g2_fill_1 FILLER_9_705 ();
 sg13g2_fill_1 FILLER_9_719 ();
 sg13g2_fill_1 FILLER_9_741 ();
 sg13g2_fill_1 FILLER_9_747 ();
 sg13g2_fill_1 FILLER_9_752 ();
 sg13g2_fill_1 FILLER_9_832 ();
 sg13g2_fill_2 FILLER_9_842 ();
 sg13g2_decap_4 FILLER_9_848 ();
 sg13g2_decap_8 FILLER_9_856 ();
 sg13g2_fill_1 FILLER_9_863 ();
 sg13g2_fill_2 FILLER_9_872 ();
 sg13g2_fill_1 FILLER_9_874 ();
 sg13g2_fill_1 FILLER_9_880 ();
 sg13g2_fill_2 FILLER_9_890 ();
 sg13g2_fill_1 FILLER_9_892 ();
 sg13g2_fill_2 FILLER_9_919 ();
 sg13g2_decap_4 FILLER_9_925 ();
 sg13g2_fill_2 FILLER_9_954 ();
 sg13g2_fill_1 FILLER_9_1019 ();
 sg13g2_fill_2 FILLER_9_1027 ();
 sg13g2_fill_1 FILLER_9_1039 ();
 sg13g2_fill_1 FILLER_9_1087 ();
 sg13g2_fill_2 FILLER_9_1118 ();
 sg13g2_fill_1 FILLER_9_1120 ();
 sg13g2_decap_4 FILLER_9_1143 ();
 sg13g2_fill_2 FILLER_9_1147 ();
 sg13g2_decap_4 FILLER_9_1184 ();
 sg13g2_fill_1 FILLER_9_1188 ();
 sg13g2_decap_4 FILLER_9_1197 ();
 sg13g2_fill_2 FILLER_9_1251 ();
 sg13g2_fill_1 FILLER_9_1253 ();
 sg13g2_decap_4 FILLER_9_1297 ();
 sg13g2_decap_4 FILLER_9_1305 ();
 sg13g2_decap_8 FILLER_9_1322 ();
 sg13g2_decap_8 FILLER_9_1344 ();
 sg13g2_decap_8 FILLER_9_1351 ();
 sg13g2_decap_4 FILLER_9_1358 ();
 sg13g2_fill_2 FILLER_9_1362 ();
 sg13g2_fill_1 FILLER_9_1372 ();
 sg13g2_fill_1 FILLER_9_1382 ();
 sg13g2_fill_1 FILLER_9_1413 ();
 sg13g2_fill_2 FILLER_9_1418 ();
 sg13g2_fill_1 FILLER_9_1420 ();
 sg13g2_fill_2 FILLER_9_1425 ();
 sg13g2_fill_1 FILLER_9_1427 ();
 sg13g2_fill_2 FILLER_9_1445 ();
 sg13g2_fill_1 FILLER_9_1455 ();
 sg13g2_fill_2 FILLER_9_1482 ();
 sg13g2_fill_2 FILLER_9_1488 ();
 sg13g2_fill_2 FILLER_9_1494 ();
 sg13g2_fill_1 FILLER_9_1496 ();
 sg13g2_fill_2 FILLER_9_1527 ();
 sg13g2_fill_1 FILLER_9_1529 ();
 sg13g2_fill_2 FILLER_9_1542 ();
 sg13g2_fill_1 FILLER_9_1579 ();
 sg13g2_fill_2 FILLER_9_1584 ();
 sg13g2_fill_2 FILLER_9_1611 ();
 sg13g2_fill_1 FILLER_9_1617 ();
 sg13g2_fill_1 FILLER_9_1623 ();
 sg13g2_fill_1 FILLER_9_1638 ();
 sg13g2_fill_2 FILLER_9_1651 ();
 sg13g2_fill_1 FILLER_9_1676 ();
 sg13g2_decap_8 FILLER_9_1698 ();
 sg13g2_fill_1 FILLER_9_1705 ();
 sg13g2_fill_2 FILLER_9_1735 ();
 sg13g2_decap_8 FILLER_9_1768 ();
 sg13g2_fill_2 FILLER_9_1775 ();
 sg13g2_decap_4 FILLER_9_1794 ();
 sg13g2_fill_2 FILLER_9_1798 ();
 sg13g2_decap_4 FILLER_9_1808 ();
 sg13g2_fill_1 FILLER_9_1816 ();
 sg13g2_decap_8 FILLER_9_1821 ();
 sg13g2_fill_2 FILLER_9_1828 ();
 sg13g2_fill_1 FILLER_9_1840 ();
 sg13g2_fill_2 FILLER_9_1845 ();
 sg13g2_decap_4 FILLER_9_1855 ();
 sg13g2_fill_2 FILLER_9_1859 ();
 sg13g2_decap_8 FILLER_9_1873 ();
 sg13g2_decap_8 FILLER_9_1880 ();
 sg13g2_decap_8 FILLER_9_1887 ();
 sg13g2_decap_8 FILLER_9_1894 ();
 sg13g2_decap_8 FILLER_9_1901 ();
 sg13g2_fill_1 FILLER_9_1956 ();
 sg13g2_fill_1 FILLER_9_1973 ();
 sg13g2_fill_2 FILLER_9_2005 ();
 sg13g2_fill_2 FILLER_9_2023 ();
 sg13g2_fill_2 FILLER_9_2033 ();
 sg13g2_decap_8 FILLER_9_2071 ();
 sg13g2_fill_2 FILLER_9_2078 ();
 sg13g2_decap_8 FILLER_9_2114 ();
 sg13g2_decap_8 FILLER_9_2121 ();
 sg13g2_decap_8 FILLER_9_2128 ();
 sg13g2_decap_8 FILLER_9_2135 ();
 sg13g2_fill_1 FILLER_9_2142 ();
 sg13g2_decap_8 FILLER_9_2177 ();
 sg13g2_decap_8 FILLER_9_2184 ();
 sg13g2_fill_1 FILLER_9_2191 ();
 sg13g2_decap_8 FILLER_9_2245 ();
 sg13g2_fill_1 FILLER_9_2252 ();
 sg13g2_fill_2 FILLER_9_2256 ();
 sg13g2_fill_1 FILLER_9_2258 ();
 sg13g2_decap_4 FILLER_9_2262 ();
 sg13g2_fill_1 FILLER_9_2292 ();
 sg13g2_decap_8 FILLER_9_2297 ();
 sg13g2_decap_4 FILLER_9_2360 ();
 sg13g2_fill_1 FILLER_9_2364 ();
 sg13g2_decap_4 FILLER_9_2368 ();
 sg13g2_fill_2 FILLER_9_2387 ();
 sg13g2_decap_4 FILLER_9_2394 ();
 sg13g2_decap_4 FILLER_9_2402 ();
 sg13g2_fill_1 FILLER_9_2406 ();
 sg13g2_fill_2 FILLER_9_2412 ();
 sg13g2_fill_1 FILLER_9_2414 ();
 sg13g2_fill_2 FILLER_9_2425 ();
 sg13g2_fill_1 FILLER_9_2427 ();
 sg13g2_decap_8 FILLER_9_2431 ();
 sg13g2_decap_8 FILLER_9_2443 ();
 sg13g2_decap_8 FILLER_9_2450 ();
 sg13g2_fill_1 FILLER_9_2457 ();
 sg13g2_decap_8 FILLER_9_2462 ();
 sg13g2_fill_2 FILLER_9_2469 ();
 sg13g2_fill_1 FILLER_9_2471 ();
 sg13g2_fill_2 FILLER_9_2482 ();
 sg13g2_decap_8 FILLER_9_2505 ();
 sg13g2_decap_8 FILLER_9_2512 ();
 sg13g2_fill_2 FILLER_9_2519 ();
 sg13g2_fill_2 FILLER_9_2535 ();
 sg13g2_decap_4 FILLER_9_2545 ();
 sg13g2_fill_2 FILLER_9_2549 ();
 sg13g2_decap_4 FILLER_9_2564 ();
 sg13g2_fill_2 FILLER_9_2568 ();
 sg13g2_decap_8 FILLER_9_2574 ();
 sg13g2_decap_4 FILLER_9_2581 ();
 sg13g2_fill_2 FILLER_9_2585 ();
 sg13g2_decap_8 FILLER_9_2617 ();
 sg13g2_decap_4 FILLER_9_2624 ();
 sg13g2_fill_2 FILLER_9_2628 ();
 sg13g2_decap_8 FILLER_9_2656 ();
 sg13g2_decap_8 FILLER_9_2663 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_fill_1 FILLER_10_30 ();
 sg13g2_fill_2 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_37 ();
 sg13g2_fill_1 FILLER_10_42 ();
 sg13g2_fill_1 FILLER_10_47 ();
 sg13g2_decap_8 FILLER_10_52 ();
 sg13g2_decap_8 FILLER_10_59 ();
 sg13g2_fill_2 FILLER_10_123 ();
 sg13g2_decap_4 FILLER_10_129 ();
 sg13g2_fill_2 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_139 ();
 sg13g2_fill_2 FILLER_10_155 ();
 sg13g2_fill_1 FILLER_10_157 ();
 sg13g2_fill_1 FILLER_10_166 ();
 sg13g2_fill_1 FILLER_10_214 ();
 sg13g2_fill_2 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_259 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_fill_1 FILLER_10_328 ();
 sg13g2_fill_1 FILLER_10_359 ();
 sg13g2_fill_2 FILLER_10_381 ();
 sg13g2_fill_1 FILLER_10_390 ();
 sg13g2_fill_1 FILLER_10_491 ();
 sg13g2_fill_1 FILLER_10_520 ();
 sg13g2_decap_4 FILLER_10_553 ();
 sg13g2_fill_2 FILLER_10_578 ();
 sg13g2_fill_1 FILLER_10_597 ();
 sg13g2_fill_1 FILLER_10_626 ();
 sg13g2_decap_4 FILLER_10_660 ();
 sg13g2_fill_1 FILLER_10_675 ();
 sg13g2_fill_1 FILLER_10_683 ();
 sg13g2_fill_2 FILLER_10_724 ();
 sg13g2_fill_2 FILLER_10_752 ();
 sg13g2_fill_2 FILLER_10_767 ();
 sg13g2_fill_1 FILLER_10_769 ();
 sg13g2_fill_2 FILLER_10_775 ();
 sg13g2_decap_4 FILLER_10_786 ();
 sg13g2_fill_2 FILLER_10_790 ();
 sg13g2_fill_2 FILLER_10_859 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_fill_1 FILLER_10_875 ();
 sg13g2_fill_1 FILLER_10_893 ();
 sg13g2_fill_1 FILLER_10_902 ();
 sg13g2_fill_1 FILLER_10_907 ();
 sg13g2_decap_8 FILLER_10_917 ();
 sg13g2_fill_2 FILLER_10_924 ();
 sg13g2_fill_1 FILLER_10_926 ();
 sg13g2_fill_1 FILLER_10_952 ();
 sg13g2_fill_2 FILLER_10_977 ();
 sg13g2_fill_1 FILLER_10_995 ();
 sg13g2_fill_1 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1038 ();
 sg13g2_decap_4 FILLER_10_1070 ();
 sg13g2_fill_2 FILLER_10_1074 ();
 sg13g2_decap_8 FILLER_10_1085 ();
 sg13g2_fill_2 FILLER_10_1110 ();
 sg13g2_fill_1 FILLER_10_1112 ();
 sg13g2_decap_8 FILLER_10_1181 ();
 sg13g2_decap_8 FILLER_10_1188 ();
 sg13g2_decap_8 FILLER_10_1195 ();
 sg13g2_decap_4 FILLER_10_1202 ();
 sg13g2_fill_2 FILLER_10_1206 ();
 sg13g2_fill_1 FILLER_10_1216 ();
 sg13g2_fill_1 FILLER_10_1222 ();
 sg13g2_fill_1 FILLER_10_1243 ();
 sg13g2_fill_2 FILLER_10_1270 ();
 sg13g2_fill_2 FILLER_10_1276 ();
 sg13g2_decap_8 FILLER_10_1299 ();
 sg13g2_fill_1 FILLER_10_1314 ();
 sg13g2_fill_2 FILLER_10_1324 ();
 sg13g2_fill_2 FILLER_10_1330 ();
 sg13g2_fill_2 FILLER_10_1366 ();
 sg13g2_fill_1 FILLER_10_1368 ();
 sg13g2_decap_8 FILLER_10_1399 ();
 sg13g2_decap_4 FILLER_10_1406 ();
 sg13g2_fill_2 FILLER_10_1410 ();
 sg13g2_fill_2 FILLER_10_1416 ();
 sg13g2_fill_1 FILLER_10_1431 ();
 sg13g2_fill_1 FILLER_10_1437 ();
 sg13g2_fill_2 FILLER_10_1446 ();
 sg13g2_fill_1 FILLER_10_1448 ();
 sg13g2_fill_2 FILLER_10_1467 ();
 sg13g2_fill_1 FILLER_10_1469 ();
 sg13g2_fill_2 FILLER_10_1474 ();
 sg13g2_fill_1 FILLER_10_1476 ();
 sg13g2_fill_1 FILLER_10_1489 ();
 sg13g2_fill_1 FILLER_10_1511 ();
 sg13g2_decap_8 FILLER_10_1536 ();
 sg13g2_decap_8 FILLER_10_1543 ();
 sg13g2_decap_8 FILLER_10_1558 ();
 sg13g2_fill_1 FILLER_10_1565 ();
 sg13g2_fill_2 FILLER_10_1604 ();
 sg13g2_fill_1 FILLER_10_1641 ();
 sg13g2_fill_2 FILLER_10_1800 ();
 sg13g2_decap_8 FILLER_10_1806 ();
 sg13g2_fill_2 FILLER_10_1813 ();
 sg13g2_fill_1 FILLER_10_1815 ();
 sg13g2_decap_4 FILLER_10_1854 ();
 sg13g2_decap_8 FILLER_10_1862 ();
 sg13g2_decap_8 FILLER_10_1869 ();
 sg13g2_decap_8 FILLER_10_1876 ();
 sg13g2_decap_8 FILLER_10_1883 ();
 sg13g2_decap_8 FILLER_10_1890 ();
 sg13g2_fill_2 FILLER_10_1897 ();
 sg13g2_fill_1 FILLER_10_1899 ();
 sg13g2_fill_1 FILLER_10_1930 ();
 sg13g2_fill_1 FILLER_10_1937 ();
 sg13g2_fill_1 FILLER_10_1948 ();
 sg13g2_fill_2 FILLER_10_1957 ();
 sg13g2_fill_1 FILLER_10_1974 ();
 sg13g2_fill_1 FILLER_10_1985 ();
 sg13g2_fill_2 FILLER_10_2058 ();
 sg13g2_decap_4 FILLER_10_2086 ();
 sg13g2_decap_8 FILLER_10_2094 ();
 sg13g2_decap_8 FILLER_10_2101 ();
 sg13g2_decap_8 FILLER_10_2108 ();
 sg13g2_decap_4 FILLER_10_2115 ();
 sg13g2_fill_2 FILLER_10_2119 ();
 sg13g2_fill_2 FILLER_10_2142 ();
 sg13g2_fill_2 FILLER_10_2153 ();
 sg13g2_decap_8 FILLER_10_2181 ();
 sg13g2_fill_2 FILLER_10_2192 ();
 sg13g2_fill_1 FILLER_10_2259 ();
 sg13g2_fill_1 FILLER_10_2264 ();
 sg13g2_decap_8 FILLER_10_2295 ();
 sg13g2_decap_8 FILLER_10_2302 ();
 sg13g2_decap_8 FILLER_10_2309 ();
 sg13g2_fill_1 FILLER_10_2316 ();
 sg13g2_fill_1 FILLER_10_2327 ();
 sg13g2_fill_2 FILLER_10_2331 ();
 sg13g2_decap_4 FILLER_10_2337 ();
 sg13g2_fill_2 FILLER_10_2341 ();
 sg13g2_fill_1 FILLER_10_2373 ();
 sg13g2_decap_8 FILLER_10_2379 ();
 sg13g2_fill_1 FILLER_10_2416 ();
 sg13g2_fill_1 FILLER_10_2443 ();
 sg13g2_fill_1 FILLER_10_2448 ();
 sg13g2_fill_2 FILLER_10_2453 ();
 sg13g2_fill_1 FILLER_10_2461 ();
 sg13g2_fill_1 FILLER_10_2488 ();
 sg13g2_fill_1 FILLER_10_2497 ();
 sg13g2_decap_4 FILLER_10_2524 ();
 sg13g2_fill_1 FILLER_10_2528 ();
 sg13g2_fill_2 FILLER_10_2552 ();
 sg13g2_fill_1 FILLER_10_2554 ();
 sg13g2_fill_2 FILLER_10_2559 ();
 sg13g2_fill_1 FILLER_10_2561 ();
 sg13g2_fill_2 FILLER_10_2567 ();
 sg13g2_fill_1 FILLER_10_2569 ();
 sg13g2_fill_2 FILLER_10_2596 ();
 sg13g2_decap_8 FILLER_10_2611 ();
 sg13g2_fill_1 FILLER_10_2618 ();
 sg13g2_decap_8 FILLER_10_2627 ();
 sg13g2_decap_8 FILLER_10_2634 ();
 sg13g2_decap_8 FILLER_10_2641 ();
 sg13g2_decap_8 FILLER_10_2648 ();
 sg13g2_decap_8 FILLER_10_2655 ();
 sg13g2_decap_8 FILLER_10_2662 ();
 sg13g2_fill_1 FILLER_10_2669 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_16 ();
 sg13g2_decap_4 FILLER_11_34 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_4 FILLER_11_49 ();
 sg13g2_fill_2 FILLER_11_69 ();
 sg13g2_fill_1 FILLER_11_71 ();
 sg13g2_fill_1 FILLER_11_103 ();
 sg13g2_fill_2 FILLER_11_133 ();
 sg13g2_decap_4 FILLER_11_139 ();
 sg13g2_fill_1 FILLER_11_187 ();
 sg13g2_fill_1 FILLER_11_197 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_fill_2 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_251 ();
 sg13g2_fill_2 FILLER_11_258 ();
 sg13g2_decap_4 FILLER_11_290 ();
 sg13g2_fill_1 FILLER_11_294 ();
 sg13g2_fill_2 FILLER_11_304 ();
 sg13g2_fill_1 FILLER_11_306 ();
 sg13g2_fill_2 FILLER_11_349 ();
 sg13g2_fill_1 FILLER_11_351 ();
 sg13g2_fill_2 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_389 ();
 sg13g2_fill_1 FILLER_11_417 ();
 sg13g2_fill_1 FILLER_11_422 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_fill_1 FILLER_11_475 ();
 sg13g2_fill_1 FILLER_11_480 ();
 sg13g2_fill_1 FILLER_11_486 ();
 sg13g2_fill_2 FILLER_11_500 ();
 sg13g2_decap_8 FILLER_11_509 ();
 sg13g2_decap_8 FILLER_11_516 ();
 sg13g2_fill_2 FILLER_11_523 ();
 sg13g2_decap_8 FILLER_11_528 ();
 sg13g2_decap_8 FILLER_11_535 ();
 sg13g2_decap_4 FILLER_11_542 ();
 sg13g2_fill_1 FILLER_11_626 ();
 sg13g2_fill_1 FILLER_11_636 ();
 sg13g2_fill_2 FILLER_11_645 ();
 sg13g2_fill_1 FILLER_11_647 ();
 sg13g2_decap_8 FILLER_11_652 ();
 sg13g2_decap_8 FILLER_11_659 ();
 sg13g2_decap_4 FILLER_11_666 ();
 sg13g2_fill_2 FILLER_11_670 ();
 sg13g2_fill_1 FILLER_11_712 ();
 sg13g2_fill_2 FILLER_11_743 ();
 sg13g2_fill_1 FILLER_11_745 ();
 sg13g2_fill_2 FILLER_11_755 ();
 sg13g2_fill_1 FILLER_11_757 ();
 sg13g2_fill_2 FILLER_11_770 ();
 sg13g2_fill_2 FILLER_11_776 ();
 sg13g2_fill_1 FILLER_11_778 ();
 sg13g2_decap_8 FILLER_11_783 ();
 sg13g2_fill_2 FILLER_11_790 ();
 sg13g2_fill_2 FILLER_11_823 ();
 sg13g2_fill_1 FILLER_11_837 ();
 sg13g2_fill_1 FILLER_11_867 ();
 sg13g2_decap_8 FILLER_11_894 ();
 sg13g2_decap_4 FILLER_11_901 ();
 sg13g2_decap_8 FILLER_11_940 ();
 sg13g2_decap_4 FILLER_11_947 ();
 sg13g2_fill_2 FILLER_11_951 ();
 sg13g2_fill_2 FILLER_11_956 ();
 sg13g2_fill_1 FILLER_11_958 ();
 sg13g2_fill_2 FILLER_11_967 ();
 sg13g2_fill_1 FILLER_11_983 ();
 sg13g2_fill_2 FILLER_11_1001 ();
 sg13g2_fill_2 FILLER_11_1044 ();
 sg13g2_fill_1 FILLER_11_1049 ();
 sg13g2_fill_2 FILLER_11_1066 ();
 sg13g2_fill_2 FILLER_11_1075 ();
 sg13g2_decap_8 FILLER_11_1082 ();
 sg13g2_decap_8 FILLER_11_1089 ();
 sg13g2_fill_1 FILLER_11_1096 ();
 sg13g2_decap_8 FILLER_11_1101 ();
 sg13g2_decap_8 FILLER_11_1160 ();
 sg13g2_decap_8 FILLER_11_1188 ();
 sg13g2_decap_8 FILLER_11_1195 ();
 sg13g2_fill_2 FILLER_11_1202 ();
 sg13g2_fill_1 FILLER_11_1239 ();
 sg13g2_fill_2 FILLER_11_1276 ();
 sg13g2_fill_2 FILLER_11_1297 ();
 sg13g2_fill_1 FILLER_11_1299 ();
 sg13g2_fill_2 FILLER_11_1315 ();
 sg13g2_fill_2 FILLER_11_1389 ();
 sg13g2_fill_2 FILLER_11_1412 ();
 sg13g2_fill_1 FILLER_11_1414 ();
 sg13g2_decap_8 FILLER_11_1459 ();
 sg13g2_fill_1 FILLER_11_1466 ();
 sg13g2_fill_2 FILLER_11_1472 ();
 sg13g2_decap_8 FILLER_11_1540 ();
 sg13g2_fill_2 FILLER_11_1547 ();
 sg13g2_decap_4 FILLER_11_1553 ();
 sg13g2_fill_1 FILLER_11_1557 ();
 sg13g2_fill_2 FILLER_11_1567 ();
 sg13g2_fill_1 FILLER_11_1569 ();
 sg13g2_decap_8 FILLER_11_1627 ();
 sg13g2_decap_4 FILLER_11_1634 ();
 sg13g2_fill_2 FILLER_11_1677 ();
 sg13g2_fill_1 FILLER_11_1710 ();
 sg13g2_fill_2 FILLER_11_1718 ();
 sg13g2_fill_1 FILLER_11_1750 ();
 sg13g2_fill_2 FILLER_11_1782 ();
 sg13g2_fill_1 FILLER_11_1810 ();
 sg13g2_decap_4 FILLER_11_1855 ();
 sg13g2_fill_2 FILLER_11_1859 ();
 sg13g2_fill_1 FILLER_11_1865 ();
 sg13g2_fill_2 FILLER_11_1892 ();
 sg13g2_fill_1 FILLER_11_1925 ();
 sg13g2_fill_1 FILLER_11_1930 ();
 sg13g2_fill_1 FILLER_11_1941 ();
 sg13g2_fill_1 FILLER_11_2007 ();
 sg13g2_fill_2 FILLER_11_2023 ();
 sg13g2_fill_2 FILLER_11_2063 ();
 sg13g2_decap_8 FILLER_11_2087 ();
 sg13g2_decap_8 FILLER_11_2094 ();
 sg13g2_fill_1 FILLER_11_2101 ();
 sg13g2_fill_2 FILLER_11_2132 ();
 sg13g2_fill_2 FILLER_11_2147 ();
 sg13g2_decap_4 FILLER_11_2175 ();
 sg13g2_decap_8 FILLER_11_2215 ();
 sg13g2_decap_4 FILLER_11_2222 ();
 sg13g2_fill_2 FILLER_11_2226 ();
 sg13g2_fill_1 FILLER_11_2237 ();
 sg13g2_fill_2 FILLER_11_2269 ();
 sg13g2_fill_2 FILLER_11_2282 ();
 sg13g2_decap_4 FILLER_11_2357 ();
 sg13g2_fill_2 FILLER_11_2372 ();
 sg13g2_fill_1 FILLER_11_2374 ();
 sg13g2_fill_1 FILLER_11_2407 ();
 sg13g2_decap_4 FILLER_11_2412 ();
 sg13g2_fill_1 FILLER_11_2416 ();
 sg13g2_fill_1 FILLER_11_2438 ();
 sg13g2_fill_1 FILLER_11_2444 ();
 sg13g2_fill_1 FILLER_11_2450 ();
 sg13g2_fill_1 FILLER_11_2535 ();
 sg13g2_fill_2 FILLER_11_2572 ();
 sg13g2_fill_1 FILLER_11_2604 ();
 sg13g2_decap_4 FILLER_11_2609 ();
 sg13g2_fill_2 FILLER_11_2613 ();
 sg13g2_decap_8 FILLER_11_2641 ();
 sg13g2_decap_8 FILLER_11_2648 ();
 sg13g2_decap_8 FILLER_11_2655 ();
 sg13g2_decap_8 FILLER_11_2662 ();
 sg13g2_fill_1 FILLER_11_2669 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_41 ();
 sg13g2_fill_1 FILLER_12_43 ();
 sg13g2_fill_1 FILLER_12_65 ();
 sg13g2_fill_2 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_86 ();
 sg13g2_decap_4 FILLER_12_93 ();
 sg13g2_fill_1 FILLER_12_97 ();
 sg13g2_decap_4 FILLER_12_102 ();
 sg13g2_fill_1 FILLER_12_106 ();
 sg13g2_decap_4 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_115 ();
 sg13g2_decap_8 FILLER_12_120 ();
 sg13g2_decap_8 FILLER_12_127 ();
 sg13g2_fill_2 FILLER_12_164 ();
 sg13g2_fill_2 FILLER_12_184 ();
 sg13g2_fill_2 FILLER_12_199 ();
 sg13g2_fill_1 FILLER_12_201 ();
 sg13g2_decap_4 FILLER_12_214 ();
 sg13g2_fill_2 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_224 ();
 sg13g2_fill_1 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_243 ();
 sg13g2_decap_8 FILLER_12_250 ();
 sg13g2_decap_4 FILLER_12_257 ();
 sg13g2_fill_1 FILLER_12_261 ();
 sg13g2_decap_8 FILLER_12_271 ();
 sg13g2_decap_8 FILLER_12_278 ();
 sg13g2_decap_8 FILLER_12_285 ();
 sg13g2_fill_2 FILLER_12_292 ();
 sg13g2_fill_1 FILLER_12_294 ();
 sg13g2_fill_1 FILLER_12_299 ();
 sg13g2_decap_4 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_334 ();
 sg13g2_fill_1 FILLER_12_345 ();
 sg13g2_decap_4 FILLER_12_351 ();
 sg13g2_fill_2 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_fill_2 FILLER_12_399 ();
 sg13g2_fill_1 FILLER_12_401 ();
 sg13g2_decap_8 FILLER_12_517 ();
 sg13g2_decap_8 FILLER_12_524 ();
 sg13g2_fill_2 FILLER_12_553 ();
 sg13g2_fill_1 FILLER_12_559 ();
 sg13g2_decap_8 FILLER_12_633 ();
 sg13g2_fill_2 FILLER_12_640 ();
 sg13g2_fill_2 FILLER_12_660 ();
 sg13g2_fill_1 FILLER_12_662 ();
 sg13g2_fill_2 FILLER_12_693 ();
 sg13g2_fill_1 FILLER_12_695 ();
 sg13g2_fill_2 FILLER_12_710 ();
 sg13g2_decap_4 FILLER_12_789 ();
 sg13g2_fill_1 FILLER_12_793 ();
 sg13g2_fill_2 FILLER_12_825 ();
 sg13g2_fill_1 FILLER_12_827 ();
 sg13g2_fill_2 FILLER_12_845 ();
 sg13g2_fill_1 FILLER_12_847 ();
 sg13g2_fill_2 FILLER_12_869 ();
 sg13g2_fill_2 FILLER_12_901 ();
 sg13g2_fill_1 FILLER_12_903 ();
 sg13g2_fill_2 FILLER_12_970 ();
 sg13g2_fill_2 FILLER_12_981 ();
 sg13g2_decap_4 FILLER_12_990 ();
 sg13g2_fill_1 FILLER_12_997 ();
 sg13g2_fill_1 FILLER_12_1001 ();
 sg13g2_decap_4 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_12_1038 ();
 sg13g2_fill_1 FILLER_12_1045 ();
 sg13g2_fill_2 FILLER_12_1059 ();
 sg13g2_fill_1 FILLER_12_1087 ();
 sg13g2_decap_4 FILLER_12_1092 ();
 sg13g2_decap_8 FILLER_12_1101 ();
 sg13g2_decap_4 FILLER_12_1108 ();
 sg13g2_fill_1 FILLER_12_1112 ();
 sg13g2_fill_2 FILLER_12_1134 ();
 sg13g2_fill_2 FILLER_12_1144 ();
 sg13g2_fill_1 FILLER_12_1146 ();
 sg13g2_decap_4 FILLER_12_1155 ();
 sg13g2_fill_1 FILLER_12_1209 ();
 sg13g2_fill_1 FILLER_12_1282 ();
 sg13g2_fill_1 FILLER_12_1288 ();
 sg13g2_fill_1 FILLER_12_1315 ();
 sg13g2_fill_2 FILLER_12_1359 ();
 sg13g2_decap_8 FILLER_12_1400 ();
 sg13g2_fill_2 FILLER_12_1407 ();
 sg13g2_fill_1 FILLER_12_1461 ();
 sg13g2_fill_1 FILLER_12_1470 ();
 sg13g2_fill_2 FILLER_12_1479 ();
 sg13g2_decap_4 FILLER_12_1507 ();
 sg13g2_decap_8 FILLER_12_1528 ();
 sg13g2_decap_4 FILLER_12_1535 ();
 sg13g2_fill_1 FILLER_12_1539 ();
 sg13g2_decap_8 FILLER_12_1588 ();
 sg13g2_decap_8 FILLER_12_1595 ();
 sg13g2_fill_2 FILLER_12_1602 ();
 sg13g2_fill_1 FILLER_12_1608 ();
 sg13g2_fill_1 FILLER_12_1614 ();
 sg13g2_fill_1 FILLER_12_1685 ();
 sg13g2_decap_8 FILLER_12_1715 ();
 sg13g2_decap_4 FILLER_12_1722 ();
 sg13g2_fill_1 FILLER_12_1726 ();
 sg13g2_fill_2 FILLER_12_1735 ();
 sg13g2_decap_8 FILLER_12_1762 ();
 sg13g2_fill_2 FILLER_12_1769 ();
 sg13g2_fill_2 FILLER_12_1784 ();
 sg13g2_fill_1 FILLER_12_1786 ();
 sg13g2_fill_2 FILLER_12_1791 ();
 sg13g2_fill_1 FILLER_12_1793 ();
 sg13g2_fill_2 FILLER_12_1820 ();
 sg13g2_fill_1 FILLER_12_1827 ();
 sg13g2_decap_4 FILLER_12_1836 ();
 sg13g2_fill_2 FILLER_12_1840 ();
 sg13g2_decap_8 FILLER_12_1846 ();
 sg13g2_fill_2 FILLER_12_1853 ();
 sg13g2_fill_1 FILLER_12_1855 ();
 sg13g2_fill_2 FILLER_12_1899 ();
 sg13g2_fill_2 FILLER_12_1932 ();
 sg13g2_fill_1 FILLER_12_1944 ();
 sg13g2_fill_2 FILLER_12_2046 ();
 sg13g2_fill_1 FILLER_12_2048 ();
 sg13g2_decap_8 FILLER_12_2087 ();
 sg13g2_decap_4 FILLER_12_2094 ();
 sg13g2_decap_4 FILLER_12_2124 ();
 sg13g2_fill_1 FILLER_12_2128 ();
 sg13g2_fill_1 FILLER_12_2138 ();
 sg13g2_fill_1 FILLER_12_2165 ();
 sg13g2_decap_8 FILLER_12_2170 ();
 sg13g2_decap_8 FILLER_12_2177 ();
 sg13g2_decap_8 FILLER_12_2184 ();
 sg13g2_decap_4 FILLER_12_2211 ();
 sg13g2_decap_8 FILLER_12_2233 ();
 sg13g2_decap_4 FILLER_12_2240 ();
 sg13g2_decap_8 FILLER_12_2253 ();
 sg13g2_fill_2 FILLER_12_2260 ();
 sg13g2_fill_1 FILLER_12_2262 ();
 sg13g2_decap_8 FILLER_12_2267 ();
 sg13g2_decap_8 FILLER_12_2282 ();
 sg13g2_fill_1 FILLER_12_2289 ();
 sg13g2_decap_8 FILLER_12_2300 ();
 sg13g2_fill_2 FILLER_12_2307 ();
 sg13g2_decap_8 FILLER_12_2318 ();
 sg13g2_fill_1 FILLER_12_2325 ();
 sg13g2_fill_1 FILLER_12_2398 ();
 sg13g2_fill_1 FILLER_12_2407 ();
 sg13g2_decap_4 FILLER_12_2418 ();
 sg13g2_fill_2 FILLER_12_2422 ();
 sg13g2_fill_2 FILLER_12_2436 ();
 sg13g2_fill_2 FILLER_12_2453 ();
 sg13g2_fill_1 FILLER_12_2455 ();
 sg13g2_decap_8 FILLER_12_2471 ();
 sg13g2_decap_4 FILLER_12_2478 ();
 sg13g2_fill_2 FILLER_12_2486 ();
 sg13g2_decap_8 FILLER_12_2497 ();
 sg13g2_fill_2 FILLER_12_2508 ();
 sg13g2_fill_2 FILLER_12_2519 ();
 sg13g2_fill_1 FILLER_12_2532 ();
 sg13g2_fill_1 FILLER_12_2559 ();
 sg13g2_decap_4 FILLER_12_2568 ();
 sg13g2_fill_1 FILLER_12_2572 ();
 sg13g2_fill_1 FILLER_12_2577 ();
 sg13g2_fill_1 FILLER_12_2586 ();
 sg13g2_fill_1 FILLER_12_2592 ();
 sg13g2_fill_1 FILLER_12_2619 ();
 sg13g2_decap_8 FILLER_12_2636 ();
 sg13g2_decap_8 FILLER_12_2643 ();
 sg13g2_decap_8 FILLER_12_2650 ();
 sg13g2_decap_8 FILLER_12_2657 ();
 sg13g2_decap_4 FILLER_12_2664 ();
 sg13g2_fill_2 FILLER_12_2668 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_4 ();
 sg13g2_fill_2 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_96 ();
 sg13g2_fill_1 FILLER_13_101 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_250 ();
 sg13g2_fill_2 FILLER_13_286 ();
 sg13g2_fill_1 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_320 ();
 sg13g2_fill_2 FILLER_13_382 ();
 sg13g2_decap_4 FILLER_13_388 ();
 sg13g2_fill_1 FILLER_13_392 ();
 sg13g2_fill_1 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_431 ();
 sg13g2_fill_2 FILLER_13_442 ();
 sg13g2_fill_1 FILLER_13_461 ();
 sg13g2_decap_4 FILLER_13_528 ();
 sg13g2_fill_1 FILLER_13_532 ();
 sg13g2_fill_2 FILLER_13_559 ();
 sg13g2_fill_2 FILLER_13_568 ();
 sg13g2_fill_2 FILLER_13_581 ();
 sg13g2_fill_2 FILLER_13_600 ();
 sg13g2_fill_2 FILLER_13_615 ();
 sg13g2_fill_2 FILLER_13_682 ();
 sg13g2_fill_1 FILLER_13_684 ();
 sg13g2_decap_8 FILLER_13_694 ();
 sg13g2_fill_1 FILLER_13_701 ();
 sg13g2_decap_8 FILLER_13_705 ();
 sg13g2_fill_1 FILLER_13_712 ();
 sg13g2_fill_1 FILLER_13_717 ();
 sg13g2_fill_2 FILLER_13_753 ();
 sg13g2_fill_2 FILLER_13_791 ();
 sg13g2_fill_1 FILLER_13_793 ();
 sg13g2_fill_1 FILLER_13_807 ();
 sg13g2_fill_1 FILLER_13_865 ();
 sg13g2_fill_2 FILLER_13_883 ();
 sg13g2_fill_1 FILLER_13_885 ();
 sg13g2_fill_2 FILLER_13_912 ();
 sg13g2_fill_1 FILLER_13_914 ();
 sg13g2_fill_1 FILLER_13_919 ();
 sg13g2_fill_2 FILLER_13_924 ();
 sg13g2_fill_1 FILLER_13_926 ();
 sg13g2_fill_1 FILLER_13_952 ();
 sg13g2_fill_1 FILLER_13_961 ();
 sg13g2_decap_4 FILLER_13_988 ();
 sg13g2_fill_2 FILLER_13_992 ();
 sg13g2_decap_4 FILLER_13_1020 ();
 sg13g2_fill_1 FILLER_13_1054 ();
 sg13g2_fill_1 FILLER_13_1117 ();
 sg13g2_fill_2 FILLER_13_1122 ();
 sg13g2_fill_2 FILLER_13_1129 ();
 sg13g2_fill_2 FILLER_13_1135 ();
 sg13g2_fill_1 FILLER_13_1141 ();
 sg13g2_fill_2 FILLER_13_1168 ();
 sg13g2_decap_4 FILLER_13_1191 ();
 sg13g2_fill_1 FILLER_13_1208 ();
 sg13g2_fill_1 FILLER_13_1214 ();
 sg13g2_fill_2 FILLER_13_1229 ();
 sg13g2_fill_1 FILLER_13_1231 ();
 sg13g2_fill_1 FILLER_13_1271 ();
 sg13g2_decap_4 FILLER_13_1347 ();
 sg13g2_fill_2 FILLER_13_1351 ();
 sg13g2_fill_2 FILLER_13_1440 ();
 sg13g2_fill_2 FILLER_13_1472 ();
 sg13g2_fill_1 FILLER_13_1474 ();
 sg13g2_decap_8 FILLER_13_1501 ();
 sg13g2_fill_2 FILLER_13_1534 ();
 sg13g2_fill_2 FILLER_13_1562 ();
 sg13g2_decap_8 FILLER_13_1576 ();
 sg13g2_decap_4 FILLER_13_1583 ();
 sg13g2_fill_1 FILLER_13_1587 ();
 sg13g2_decap_8 FILLER_13_1618 ();
 sg13g2_decap_4 FILLER_13_1625 ();
 sg13g2_fill_2 FILLER_13_1629 ();
 sg13g2_fill_1 FILLER_13_1647 ();
 sg13g2_fill_1 FILLER_13_1713 ();
 sg13g2_fill_1 FILLER_13_1744 ();
 sg13g2_fill_1 FILLER_13_1752 ();
 sg13g2_fill_1 FILLER_13_1786 ();
 sg13g2_decap_4 FILLER_13_1813 ();
 sg13g2_fill_2 FILLER_13_1817 ();
 sg13g2_decap_8 FILLER_13_1827 ();
 sg13g2_decap_8 FILLER_13_1834 ();
 sg13g2_decap_8 FILLER_13_1841 ();
 sg13g2_decap_8 FILLER_13_1848 ();
 sg13g2_fill_2 FILLER_13_1855 ();
 sg13g2_fill_1 FILLER_13_1857 ();
 sg13g2_fill_1 FILLER_13_1901 ();
 sg13g2_fill_1 FILLER_13_2015 ();
 sg13g2_fill_2 FILLER_13_2020 ();
 sg13g2_fill_1 FILLER_13_2048 ();
 sg13g2_fill_1 FILLER_13_2122 ();
 sg13g2_fill_1 FILLER_13_2127 ();
 sg13g2_fill_1 FILLER_13_2136 ();
 sg13g2_decap_4 FILLER_13_2142 ();
 sg13g2_fill_1 FILLER_13_2151 ();
 sg13g2_decap_8 FILLER_13_2178 ();
 sg13g2_fill_1 FILLER_13_2185 ();
 sg13g2_fill_1 FILLER_13_2200 ();
 sg13g2_fill_1 FILLER_13_2220 ();
 sg13g2_fill_1 FILLER_13_2229 ();
 sg13g2_decap_4 FILLER_13_2238 ();
 sg13g2_fill_1 FILLER_13_2242 ();
 sg13g2_fill_1 FILLER_13_2259 ();
 sg13g2_fill_1 FILLER_13_2268 ();
 sg13g2_fill_2 FILLER_13_2276 ();
 sg13g2_fill_1 FILLER_13_2278 ();
 sg13g2_fill_1 FILLER_13_2319 ();
 sg13g2_fill_1 FILLER_13_2324 ();
 sg13g2_fill_2 FILLER_13_2344 ();
 sg13g2_decap_8 FILLER_13_2356 ();
 sg13g2_decap_8 FILLER_13_2363 ();
 sg13g2_decap_8 FILLER_13_2370 ();
 sg13g2_decap_4 FILLER_13_2377 ();
 sg13g2_fill_1 FILLER_13_2385 ();
 sg13g2_decap_4 FILLER_13_2410 ();
 sg13g2_fill_2 FILLER_13_2423 ();
 sg13g2_decap_4 FILLER_13_2442 ();
 sg13g2_fill_2 FILLER_13_2446 ();
 sg13g2_decap_8 FILLER_13_2453 ();
 sg13g2_decap_8 FILLER_13_2460 ();
 sg13g2_decap_4 FILLER_13_2467 ();
 sg13g2_decap_4 FILLER_13_2476 ();
 sg13g2_fill_1 FILLER_13_2480 ();
 sg13g2_decap_8 FILLER_13_2494 ();
 sg13g2_decap_8 FILLER_13_2501 ();
 sg13g2_decap_8 FILLER_13_2508 ();
 sg13g2_decap_4 FILLER_13_2515 ();
 sg13g2_decap_8 FILLER_13_2523 ();
 sg13g2_fill_2 FILLER_13_2549 ();
 sg13g2_fill_1 FILLER_13_2559 ();
 sg13g2_decap_8 FILLER_13_2564 ();
 sg13g2_fill_1 FILLER_13_2571 ();
 sg13g2_fill_1 FILLER_13_2581 ();
 sg13g2_fill_1 FILLER_13_2587 ();
 sg13g2_fill_2 FILLER_13_2603 ();
 sg13g2_decap_4 FILLER_13_2665 ();
 sg13g2_fill_1 FILLER_13_2669 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_43 ();
 sg13g2_fill_2 FILLER_14_57 ();
 sg13g2_fill_2 FILLER_14_95 ();
 sg13g2_fill_1 FILLER_14_102 ();
 sg13g2_fill_2 FILLER_14_129 ();
 sg13g2_fill_2 FILLER_14_140 ();
 sg13g2_fill_1 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_188 ();
 sg13g2_fill_1 FILLER_14_225 ();
 sg13g2_fill_2 FILLER_14_256 ();
 sg13g2_fill_1 FILLER_14_258 ();
 sg13g2_decap_4 FILLER_14_263 ();
 sg13g2_fill_1 FILLER_14_272 ();
 sg13g2_fill_2 FILLER_14_303 ();
 sg13g2_fill_1 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_fill_2 FILLER_14_495 ();
 sg13g2_fill_1 FILLER_14_501 ();
 sg13g2_fill_1 FILLER_14_506 ();
 sg13g2_fill_1 FILLER_14_511 ();
 sg13g2_fill_1 FILLER_14_544 ();
 sg13g2_fill_2 FILLER_14_552 ();
 sg13g2_fill_2 FILLER_14_576 ();
 sg13g2_fill_1 FILLER_14_581 ();
 sg13g2_fill_2 FILLER_14_608 ();
 sg13g2_decap_4 FILLER_14_622 ();
 sg13g2_decap_4 FILLER_14_634 ();
 sg13g2_fill_2 FILLER_14_638 ();
 sg13g2_fill_2 FILLER_14_691 ();
 sg13g2_fill_1 FILLER_14_697 ();
 sg13g2_fill_2 FILLER_14_706 ();
 sg13g2_fill_1 FILLER_14_708 ();
 sg13g2_fill_2 FILLER_14_735 ();
 sg13g2_fill_2 FILLER_14_794 ();
 sg13g2_fill_1 FILLER_14_801 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_fill_1 FILLER_14_814 ();
 sg13g2_fill_1 FILLER_14_819 ();
 sg13g2_fill_1 FILLER_14_824 ();
 sg13g2_decap_4 FILLER_14_866 ();
 sg13g2_fill_2 FILLER_14_875 ();
 sg13g2_fill_1 FILLER_14_877 ();
 sg13g2_fill_2 FILLER_14_891 ();
 sg13g2_decap_4 FILLER_14_897 ();
 sg13g2_decap_4 FILLER_14_914 ();
 sg13g2_fill_1 FILLER_14_918 ();
 sg13g2_decap_8 FILLER_14_945 ();
 sg13g2_fill_2 FILLER_14_952 ();
 sg13g2_fill_1 FILLER_14_1050 ();
 sg13g2_fill_1 FILLER_14_1084 ();
 sg13g2_fill_2 FILLER_14_1097 ();
 sg13g2_decap_4 FILLER_14_1103 ();
 sg13g2_decap_8 FILLER_14_1177 ();
 sg13g2_decap_4 FILLER_14_1184 ();
 sg13g2_fill_2 FILLER_14_1213 ();
 sg13g2_fill_1 FILLER_14_1215 ();
 sg13g2_fill_1 FILLER_14_1246 ();
 sg13g2_fill_2 FILLER_14_1290 ();
 sg13g2_fill_1 FILLER_14_1292 ();
 sg13g2_decap_8 FILLER_14_1319 ();
 sg13g2_decap_4 FILLER_14_1326 ();
 sg13g2_fill_1 FILLER_14_1330 ();
 sg13g2_fill_1 FILLER_14_1336 ();
 sg13g2_decap_8 FILLER_14_1347 ();
 sg13g2_decap_8 FILLER_14_1354 ();
 sg13g2_decap_8 FILLER_14_1361 ();
 sg13g2_fill_2 FILLER_14_1368 ();
 sg13g2_decap_4 FILLER_14_1374 ();
 sg13g2_decap_4 FILLER_14_1386 ();
 sg13g2_fill_2 FILLER_14_1390 ();
 sg13g2_fill_2 FILLER_14_1406 ();
 sg13g2_fill_1 FILLER_14_1408 ();
 sg13g2_fill_2 FILLER_14_1430 ();
 sg13g2_fill_1 FILLER_14_1432 ();
 sg13g2_fill_2 FILLER_14_1498 ();
 sg13g2_decap_4 FILLER_14_1521 ();
 sg13g2_fill_1 FILLER_14_1525 ();
 sg13g2_fill_2 FILLER_14_1564 ();
 sg13g2_decap_8 FILLER_14_1598 ();
 sg13g2_decap_4 FILLER_14_1605 ();
 sg13g2_fill_1 FILLER_14_1630 ();
 sg13g2_fill_2 FILLER_14_1649 ();
 sg13g2_fill_2 FILLER_14_1663 ();
 sg13g2_fill_2 FILLER_14_1669 ();
 sg13g2_fill_2 FILLER_14_1685 ();
 sg13g2_decap_8 FILLER_14_1707 ();
 sg13g2_decap_4 FILLER_14_1714 ();
 sg13g2_fill_1 FILLER_14_1718 ();
 sg13g2_fill_2 FILLER_14_1753 ();
 sg13g2_decap_4 FILLER_14_1787 ();
 sg13g2_fill_2 FILLER_14_1795 ();
 sg13g2_fill_1 FILLER_14_1807 ();
 sg13g2_fill_2 FILLER_14_1864 ();
 sg13g2_fill_1 FILLER_14_1866 ();
 sg13g2_fill_2 FILLER_14_1892 ();
 sg13g2_fill_1 FILLER_14_1902 ();
 sg13g2_fill_2 FILLER_14_1924 ();
 sg13g2_fill_2 FILLER_14_1954 ();
 sg13g2_fill_1 FILLER_14_1960 ();
 sg13g2_fill_1 FILLER_14_1970 ();
 sg13g2_fill_1 FILLER_14_2005 ();
 sg13g2_fill_1 FILLER_14_2015 ();
 sg13g2_fill_1 FILLER_14_2020 ();
 sg13g2_fill_1 FILLER_14_2030 ();
 sg13g2_fill_1 FILLER_14_2035 ();
 sg13g2_fill_2 FILLER_14_2062 ();
 sg13g2_fill_1 FILLER_14_2098 ();
 sg13g2_fill_2 FILLER_14_2112 ();
 sg13g2_fill_1 FILLER_14_2118 ();
 sg13g2_fill_1 FILLER_14_2124 ();
 sg13g2_fill_2 FILLER_14_2150 ();
 sg13g2_fill_1 FILLER_14_2152 ();
 sg13g2_decap_8 FILLER_14_2179 ();
 sg13g2_decap_8 FILLER_14_2186 ();
 sg13g2_fill_1 FILLER_14_2193 ();
 sg13g2_fill_2 FILLER_14_2204 ();
 sg13g2_fill_2 FILLER_14_2210 ();
 sg13g2_fill_2 FILLER_14_2227 ();
 sg13g2_fill_1 FILLER_14_2229 ();
 sg13g2_fill_1 FILLER_14_2238 ();
 sg13g2_fill_1 FILLER_14_2252 ();
 sg13g2_fill_2 FILLER_14_2265 ();
 sg13g2_fill_2 FILLER_14_2283 ();
 sg13g2_fill_1 FILLER_14_2285 ();
 sg13g2_fill_2 FILLER_14_2296 ();
 sg13g2_fill_1 FILLER_14_2298 ();
 sg13g2_fill_2 FILLER_14_2309 ();
 sg13g2_fill_1 FILLER_14_2335 ();
 sg13g2_decap_8 FILLER_14_2352 ();
 sg13g2_fill_2 FILLER_14_2359 ();
 sg13g2_decap_8 FILLER_14_2365 ();
 sg13g2_decap_4 FILLER_14_2372 ();
 sg13g2_fill_1 FILLER_14_2408 ();
 sg13g2_fill_2 FILLER_14_2413 ();
 sg13g2_decap_8 FILLER_14_2432 ();
 sg13g2_decap_8 FILLER_14_2443 ();
 sg13g2_fill_2 FILLER_14_2450 ();
 sg13g2_fill_1 FILLER_14_2473 ();
 sg13g2_decap_4 FILLER_14_2482 ();
 sg13g2_fill_1 FILLER_14_2486 ();
 sg13g2_fill_2 FILLER_14_2492 ();
 sg13g2_decap_8 FILLER_14_2500 ();
 sg13g2_fill_1 FILLER_14_2515 ();
 sg13g2_fill_1 FILLER_14_2522 ();
 sg13g2_decap_8 FILLER_14_2550 ();
 sg13g2_decap_8 FILLER_14_2557 ();
 sg13g2_decap_8 FILLER_14_2564 ();
 sg13g2_decap_8 FILLER_14_2571 ();
 sg13g2_fill_1 FILLER_14_2578 ();
 sg13g2_fill_2 FILLER_14_2591 ();
 sg13g2_fill_1 FILLER_14_2593 ();
 sg13g2_fill_1 FILLER_14_2623 ();
 sg13g2_decap_8 FILLER_14_2627 ();
 sg13g2_decap_8 FILLER_14_2638 ();
 sg13g2_decap_8 FILLER_14_2645 ();
 sg13g2_decap_8 FILLER_14_2652 ();
 sg13g2_decap_8 FILLER_14_2659 ();
 sg13g2_decap_4 FILLER_14_2666 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_37 ();
 sg13g2_fill_1 FILLER_15_43 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_2 FILLER_15_71 ();
 sg13g2_fill_1 FILLER_15_99 ();
 sg13g2_fill_2 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_149 ();
 sg13g2_fill_1 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_189 ();
 sg13g2_fill_1 FILLER_15_191 ();
 sg13g2_fill_2 FILLER_15_197 ();
 sg13g2_fill_1 FILLER_15_199 ();
 sg13g2_fill_1 FILLER_15_204 ();
 sg13g2_decap_4 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_244 ();
 sg13g2_decap_8 FILLER_15_251 ();
 sg13g2_fill_2 FILLER_15_258 ();
 sg13g2_decap_8 FILLER_15_268 ();
 sg13g2_fill_2 FILLER_15_275 ();
 sg13g2_fill_1 FILLER_15_277 ();
 sg13g2_decap_8 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_289 ();
 sg13g2_decap_4 FILLER_15_296 ();
 sg13g2_fill_1 FILLER_15_300 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_fill_2 FILLER_15_330 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_344 ();
 sg13g2_fill_2 FILLER_15_376 ();
 sg13g2_fill_2 FILLER_15_399 ();
 sg13g2_fill_1 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_410 ();
 sg13g2_fill_1 FILLER_15_416 ();
 sg13g2_fill_2 FILLER_15_421 ();
 sg13g2_fill_1 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_461 ();
 sg13g2_decap_8 FILLER_15_468 ();
 sg13g2_decap_8 FILLER_15_475 ();
 sg13g2_decap_8 FILLER_15_482 ();
 sg13g2_decap_8 FILLER_15_489 ();
 sg13g2_fill_1 FILLER_15_496 ();
 sg13g2_decap_8 FILLER_15_501 ();
 sg13g2_decap_8 FILLER_15_508 ();
 sg13g2_decap_8 FILLER_15_515 ();
 sg13g2_fill_2 FILLER_15_522 ();
 sg13g2_fill_1 FILLER_15_524 ();
 sg13g2_fill_1 FILLER_15_544 ();
 sg13g2_fill_1 FILLER_15_569 ();
 sg13g2_fill_1 FILLER_15_574 ();
 sg13g2_fill_1 FILLER_15_606 ();
 sg13g2_fill_2 FILLER_15_611 ();
 sg13g2_fill_1 FILLER_15_613 ();
 sg13g2_fill_2 FILLER_15_618 ();
 sg13g2_fill_1 FILLER_15_620 ();
 sg13g2_fill_2 FILLER_15_638 ();
 sg13g2_decap_4 FILLER_15_644 ();
 sg13g2_fill_2 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_fill_2 FILLER_15_743 ();
 sg13g2_fill_1 FILLER_15_750 ();
 sg13g2_fill_2 FILLER_15_767 ();
 sg13g2_fill_2 FILLER_15_795 ();
 sg13g2_fill_2 FILLER_15_806 ();
 sg13g2_fill_1 FILLER_15_817 ();
 sg13g2_decap_4 FILLER_15_844 ();
 sg13g2_fill_1 FILLER_15_848 ();
 sg13g2_fill_2 FILLER_15_884 ();
 sg13g2_fill_1 FILLER_15_886 ();
 sg13g2_decap_8 FILLER_15_891 ();
 sg13g2_decap_8 FILLER_15_898 ();
 sg13g2_fill_1 FILLER_15_905 ();
 sg13g2_decap_4 FILLER_15_913 ();
 sg13g2_fill_1 FILLER_15_917 ();
 sg13g2_fill_2 FILLER_15_965 ();
 sg13g2_fill_2 FILLER_15_1057 ();
 sg13g2_decap_4 FILLER_15_1089 ();
 sg13g2_fill_1 FILLER_15_1093 ();
 sg13g2_fill_2 FILLER_15_1098 ();
 sg13g2_fill_1 FILLER_15_1100 ();
 sg13g2_decap_8 FILLER_15_1106 ();
 sg13g2_decap_4 FILLER_15_1113 ();
 sg13g2_fill_1 FILLER_15_1117 ();
 sg13g2_fill_1 FILLER_15_1122 ();
 sg13g2_decap_8 FILLER_15_1127 ();
 sg13g2_decap_8 FILLER_15_1134 ();
 sg13g2_fill_2 FILLER_15_1141 ();
 sg13g2_fill_1 FILLER_15_1143 ();
 sg13g2_fill_2 FILLER_15_1156 ();
 sg13g2_decap_8 FILLER_15_1162 ();
 sg13g2_decap_8 FILLER_15_1169 ();
 sg13g2_decap_8 FILLER_15_1176 ();
 sg13g2_decap_8 FILLER_15_1183 ();
 sg13g2_decap_8 FILLER_15_1190 ();
 sg13g2_fill_2 FILLER_15_1252 ();
 sg13g2_fill_1 FILLER_15_1254 ();
 sg13g2_decap_8 FILLER_15_1287 ();
 sg13g2_fill_1 FILLER_15_1294 ();
 sg13g2_fill_1 FILLER_15_1299 ();
 sg13g2_decap_8 FILLER_15_1304 ();
 sg13g2_decap_4 FILLER_15_1311 ();
 sg13g2_fill_1 FILLER_15_1315 ();
 sg13g2_fill_2 FILLER_15_1320 ();
 sg13g2_fill_1 FILLER_15_1330 ();
 sg13g2_fill_2 FILLER_15_1361 ();
 sg13g2_fill_2 FILLER_15_1367 ();
 sg13g2_fill_2 FILLER_15_1377 ();
 sg13g2_fill_1 FILLER_15_1379 ();
 sg13g2_decap_8 FILLER_15_1384 ();
 sg13g2_decap_4 FILLER_15_1391 ();
 sg13g2_fill_1 FILLER_15_1395 ();
 sg13g2_decap_4 FILLER_15_1400 ();
 sg13g2_fill_2 FILLER_15_1404 ();
 sg13g2_decap_4 FILLER_15_1438 ();
 sg13g2_decap_8 FILLER_15_1483 ();
 sg13g2_decap_4 FILLER_15_1490 ();
 sg13g2_fill_1 FILLER_15_1494 ();
 sg13g2_fill_1 FILLER_15_1501 ();
 sg13g2_decap_8 FILLER_15_1506 ();
 sg13g2_fill_2 FILLER_15_1513 ();
 sg13g2_decap_8 FILLER_15_1519 ();
 sg13g2_decap_8 FILLER_15_1526 ();
 sg13g2_decap_8 FILLER_15_1533 ();
 sg13g2_decap_4 FILLER_15_1540 ();
 sg13g2_decap_8 FILLER_15_1548 ();
 sg13g2_decap_4 FILLER_15_1555 ();
 sg13g2_decap_4 FILLER_15_1563 ();
 sg13g2_decap_4 FILLER_15_1575 ();
 sg13g2_fill_2 FILLER_15_1584 ();
 sg13g2_fill_1 FILLER_15_1586 ();
 sg13g2_fill_1 FILLER_15_1621 ();
 sg13g2_fill_1 FILLER_15_1631 ();
 sg13g2_decap_8 FILLER_15_1655 ();
 sg13g2_fill_2 FILLER_15_1662 ();
 sg13g2_fill_1 FILLER_15_1664 ();
 sg13g2_decap_8 FILLER_15_1700 ();
 sg13g2_decap_4 FILLER_15_1707 ();
 sg13g2_fill_2 FILLER_15_1711 ();
 sg13g2_decap_4 FILLER_15_1716 ();
 sg13g2_fill_1 FILLER_15_1725 ();
 sg13g2_fill_1 FILLER_15_1756 ();
 sg13g2_fill_2 FILLER_15_1762 ();
 sg13g2_fill_2 FILLER_15_1771 ();
 sg13g2_fill_2 FILLER_15_1808 ();
 sg13g2_fill_2 FILLER_15_1849 ();
 sg13g2_fill_1 FILLER_15_1851 ();
 sg13g2_fill_2 FILLER_15_1877 ();
 sg13g2_fill_1 FILLER_15_1879 ();
 sg13g2_fill_1 FILLER_15_1943 ();
 sg13g2_fill_2 FILLER_15_1976 ();
 sg13g2_fill_1 FILLER_15_1978 ();
 sg13g2_fill_2 FILLER_15_1984 ();
 sg13g2_fill_1 FILLER_15_1990 ();
 sg13g2_decap_8 FILLER_15_1995 ();
 sg13g2_fill_2 FILLER_15_2002 ();
 sg13g2_fill_1 FILLER_15_2004 ();
 sg13g2_fill_1 FILLER_15_2031 ();
 sg13g2_fill_1 FILLER_15_2101 ();
 sg13g2_fill_2 FILLER_15_2115 ();
 sg13g2_fill_2 FILLER_15_2121 ();
 sg13g2_fill_1 FILLER_15_2152 ();
 sg13g2_fill_1 FILLER_15_2162 ();
 sg13g2_decap_8 FILLER_15_2167 ();
 sg13g2_decap_4 FILLER_15_2174 ();
 sg13g2_fill_2 FILLER_15_2178 ();
 sg13g2_fill_2 FILLER_15_2276 ();
 sg13g2_decap_4 FILLER_15_2293 ();
 sg13g2_fill_1 FILLER_15_2297 ();
 sg13g2_decap_4 FILLER_15_2325 ();
 sg13g2_fill_1 FILLER_15_2329 ();
 sg13g2_decap_4 FILLER_15_2342 ();
 sg13g2_fill_1 FILLER_15_2346 ();
 sg13g2_fill_2 FILLER_15_2352 ();
 sg13g2_fill_1 FILLER_15_2393 ();
 sg13g2_decap_4 FILLER_15_2406 ();
 sg13g2_fill_2 FILLER_15_2410 ();
 sg13g2_decap_4 FILLER_15_2438 ();
 sg13g2_fill_1 FILLER_15_2442 ();
 sg13g2_fill_2 FILLER_15_2484 ();
 sg13g2_fill_1 FILLER_15_2486 ();
 sg13g2_fill_2 FILLER_15_2501 ();
 sg13g2_fill_1 FILLER_15_2515 ();
 sg13g2_fill_2 FILLER_15_2531 ();
 sg13g2_fill_2 FILLER_15_2541 ();
 sg13g2_fill_1 FILLER_15_2551 ();
 sg13g2_fill_1 FILLER_15_2557 ();
 sg13g2_fill_2 FILLER_15_2562 ();
 sg13g2_fill_1 FILLER_15_2564 ();
 sg13g2_fill_2 FILLER_15_2593 ();
 sg13g2_fill_2 FILLER_15_2599 ();
 sg13g2_fill_2 FILLER_15_2606 ();
 sg13g2_fill_1 FILLER_15_2634 ();
 sg13g2_decap_4 FILLER_15_2640 ();
 sg13g2_fill_2 FILLER_15_2644 ();
 sg13g2_decap_8 FILLER_15_2654 ();
 sg13g2_decap_8 FILLER_15_2661 ();
 sg13g2_fill_2 FILLER_15_2668 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_6 ();
 sg13g2_fill_1 FILLER_16_8 ();
 sg13g2_fill_2 FILLER_16_13 ();
 sg13g2_fill_1 FILLER_16_15 ();
 sg13g2_fill_2 FILLER_16_20 ();
 sg13g2_fill_1 FILLER_16_48 ();
 sg13g2_fill_1 FILLER_16_75 ();
 sg13g2_fill_1 FILLER_16_81 ();
 sg13g2_fill_2 FILLER_16_87 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_150 ();
 sg13g2_decap_8 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_171 ();
 sg13g2_fill_1 FILLER_16_173 ();
 sg13g2_fill_2 FILLER_16_179 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_218 ();
 sg13g2_decap_4 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_237 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_decap_4 FILLER_16_248 ();
 sg13g2_fill_1 FILLER_16_252 ();
 sg13g2_fill_2 FILLER_16_279 ();
 sg13g2_fill_1 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_293 ();
 sg13g2_fill_1 FILLER_16_299 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_fill_2 FILLER_16_313 ();
 sg13g2_fill_1 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_fill_2 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_351 ();
 sg13g2_fill_2 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_4 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_fill_2 FILLER_16_398 ();
 sg13g2_fill_1 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_413 ();
 sg13g2_fill_2 FILLER_16_425 ();
 sg13g2_fill_2 FILLER_16_435 ();
 sg13g2_decap_4 FILLER_16_441 ();
 sg13g2_fill_2 FILLER_16_445 ();
 sg13g2_decap_8 FILLER_16_477 ();
 sg13g2_fill_2 FILLER_16_484 ();
 sg13g2_fill_1 FILLER_16_486 ();
 sg13g2_fill_2 FILLER_16_495 ();
 sg13g2_decap_4 FILLER_16_501 ();
 sg13g2_fill_2 FILLER_16_526 ();
 sg13g2_fill_1 FILLER_16_528 ();
 sg13g2_fill_2 FILLER_16_533 ();
 sg13g2_fill_1 FILLER_16_535 ();
 sg13g2_fill_1 FILLER_16_551 ();
 sg13g2_fill_1 FILLER_16_556 ();
 sg13g2_fill_1 FILLER_16_567 ();
 sg13g2_fill_1 FILLER_16_574 ();
 sg13g2_fill_2 FILLER_16_596 ();
 sg13g2_fill_1 FILLER_16_628 ();
 sg13g2_decap_8 FILLER_16_659 ();
 sg13g2_decap_8 FILLER_16_666 ();
 sg13g2_decap_4 FILLER_16_673 ();
 sg13g2_fill_1 FILLER_16_698 ();
 sg13g2_fill_1 FILLER_16_725 ();
 sg13g2_decap_4 FILLER_16_730 ();
 sg13g2_fill_1 FILLER_16_738 ();
 sg13g2_fill_2 FILLER_16_747 ();
 sg13g2_decap_8 FILLER_16_779 ();
 sg13g2_fill_2 FILLER_16_786 ();
 sg13g2_fill_2 FILLER_16_813 ();
 sg13g2_fill_1 FILLER_16_854 ();
 sg13g2_fill_2 FILLER_16_874 ();
 sg13g2_fill_1 FILLER_16_876 ();
 sg13g2_decap_8 FILLER_16_930 ();
 sg13g2_decap_4 FILLER_16_937 ();
 sg13g2_fill_1 FILLER_16_941 ();
 sg13g2_decap_8 FILLER_16_946 ();
 sg13g2_decap_8 FILLER_16_953 ();
 sg13g2_decap_8 FILLER_16_960 ();
 sg13g2_decap_8 FILLER_16_967 ();
 sg13g2_fill_2 FILLER_16_974 ();
 sg13g2_fill_2 FILLER_16_1001 ();
 sg13g2_fill_1 FILLER_16_1003 ();
 sg13g2_fill_1 FILLER_16_1030 ();
 sg13g2_fill_2 FILLER_16_1036 ();
 sg13g2_fill_1 FILLER_16_1102 ();
 sg13g2_fill_2 FILLER_16_1107 ();
 sg13g2_fill_2 FILLER_16_1135 ();
 sg13g2_fill_2 FILLER_16_1141 ();
 sg13g2_decap_8 FILLER_16_1169 ();
 sg13g2_decap_8 FILLER_16_1176 ();
 sg13g2_fill_1 FILLER_16_1204 ();
 sg13g2_fill_1 FILLER_16_1244 ();
 sg13g2_fill_1 FILLER_16_1250 ();
 sg13g2_fill_1 FILLER_16_1255 ();
 sg13g2_fill_2 FILLER_16_1260 ();
 sg13g2_fill_1 FILLER_16_1267 ();
 sg13g2_decap_8 FILLER_16_1276 ();
 sg13g2_decap_8 FILLER_16_1283 ();
 sg13g2_decap_8 FILLER_16_1290 ();
 sg13g2_decap_4 FILLER_16_1297 ();
 sg13g2_fill_2 FILLER_16_1336 ();
 sg13g2_fill_1 FILLER_16_1442 ();
 sg13g2_decap_8 FILLER_16_1532 ();
 sg13g2_decap_8 FILLER_16_1539 ();
 sg13g2_decap_8 FILLER_16_1546 ();
 sg13g2_decap_8 FILLER_16_1553 ();
 sg13g2_decap_4 FILLER_16_1560 ();
 sg13g2_fill_1 FILLER_16_1624 ();
 sg13g2_fill_1 FILLER_16_1634 ();
 sg13g2_fill_1 FILLER_16_1655 ();
 sg13g2_decap_4 FILLER_16_1664 ();
 sg13g2_fill_1 FILLER_16_1668 ();
 sg13g2_fill_2 FILLER_16_1708 ();
 sg13g2_decap_4 FILLER_16_1725 ();
 sg13g2_fill_2 FILLER_16_1756 ();
 sg13g2_fill_1 FILLER_16_1758 ();
 sg13g2_fill_1 FILLER_16_1772 ();
 sg13g2_fill_2 FILLER_16_1786 ();
 sg13g2_fill_1 FILLER_16_1788 ();
 sg13g2_fill_2 FILLER_16_1814 ();
 sg13g2_fill_1 FILLER_16_1816 ();
 sg13g2_decap_4 FILLER_16_1843 ();
 sg13g2_fill_2 FILLER_16_1847 ();
 sg13g2_fill_1 FILLER_16_1853 ();
 sg13g2_decap_8 FILLER_16_1879 ();
 sg13g2_fill_2 FILLER_16_1886 ();
 sg13g2_fill_1 FILLER_16_1901 ();
 sg13g2_fill_1 FILLER_16_1912 ();
 sg13g2_fill_1 FILLER_16_1918 ();
 sg13g2_fill_1 FILLER_16_1923 ();
 sg13g2_fill_2 FILLER_16_1928 ();
 sg13g2_fill_1 FILLER_16_1930 ();
 sg13g2_decap_8 FILLER_16_1940 ();
 sg13g2_fill_2 FILLER_16_1947 ();
 sg13g2_decap_8 FILLER_16_2005 ();
 sg13g2_fill_1 FILLER_16_2012 ();
 sg13g2_decap_4 FILLER_16_2017 ();
 sg13g2_fill_1 FILLER_16_2021 ();
 sg13g2_fill_1 FILLER_16_2027 ();
 sg13g2_fill_1 FILLER_16_2032 ();
 sg13g2_fill_1 FILLER_16_2037 ();
 sg13g2_fill_1 FILLER_16_2047 ();
 sg13g2_fill_2 FILLER_16_2053 ();
 sg13g2_fill_2 FILLER_16_2060 ();
 sg13g2_fill_1 FILLER_16_2079 ();
 sg13g2_fill_2 FILLER_16_2084 ();
 sg13g2_fill_1 FILLER_16_2086 ();
 sg13g2_fill_2 FILLER_16_2091 ();
 sg13g2_fill_1 FILLER_16_2093 ();
 sg13g2_fill_1 FILLER_16_2112 ();
 sg13g2_decap_8 FILLER_16_2117 ();
 sg13g2_fill_2 FILLER_16_2124 ();
 sg13g2_decap_8 FILLER_16_2163 ();
 sg13g2_decap_8 FILLER_16_2170 ();
 sg13g2_decap_8 FILLER_16_2177 ();
 sg13g2_decap_8 FILLER_16_2184 ();
 sg13g2_fill_1 FILLER_16_2191 ();
 sg13g2_decap_8 FILLER_16_2197 ();
 sg13g2_fill_2 FILLER_16_2204 ();
 sg13g2_fill_2 FILLER_16_2225 ();
 sg13g2_fill_2 FILLER_16_2236 ();
 sg13g2_fill_1 FILLER_16_2248 ();
 sg13g2_fill_2 FILLER_16_2253 ();
 sg13g2_decap_4 FILLER_16_2281 ();
 sg13g2_decap_8 FILLER_16_2293 ();
 sg13g2_decap_4 FILLER_16_2300 ();
 sg13g2_fill_1 FILLER_16_2304 ();
 sg13g2_fill_2 FILLER_16_2318 ();
 sg13g2_decap_8 FILLER_16_2325 ();
 sg13g2_fill_2 FILLER_16_2332 ();
 sg13g2_decap_4 FILLER_16_2391 ();
 sg13g2_fill_2 FILLER_16_2395 ();
 sg13g2_fill_2 FILLER_16_2401 ();
 sg13g2_fill_1 FILLER_16_2403 ();
 sg13g2_decap_4 FILLER_16_2408 ();
 sg13g2_fill_1 FILLER_16_2412 ();
 sg13g2_fill_2 FILLER_16_2435 ();
 sg13g2_decap_8 FILLER_16_2440 ();
 sg13g2_decap_8 FILLER_16_2447 ();
 sg13g2_decap_4 FILLER_16_2454 ();
 sg13g2_fill_2 FILLER_16_2458 ();
 sg13g2_fill_2 FILLER_16_2464 ();
 sg13g2_fill_1 FILLER_16_2500 ();
 sg13g2_fill_1 FILLER_16_2513 ();
 sg13g2_fill_1 FILLER_16_2519 ();
 sg13g2_decap_8 FILLER_16_2525 ();
 sg13g2_fill_1 FILLER_16_2579 ();
 sg13g2_fill_1 FILLER_16_2592 ();
 sg13g2_fill_2 FILLER_16_2614 ();
 sg13g2_fill_1 FILLER_16_2616 ();
 sg13g2_decap_4 FILLER_16_2621 ();
 sg13g2_fill_2 FILLER_16_2630 ();
 sg13g2_fill_2 FILLER_16_2642 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_37 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_fill_2 FILLER_17_60 ();
 sg13g2_fill_1 FILLER_17_62 ();
 sg13g2_fill_1 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_99 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_fill_2 FILLER_17_128 ();
 sg13g2_fill_1 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_fill_2 FILLER_17_156 ();
 sg13g2_decap_8 FILLER_17_162 ();
 sg13g2_decap_4 FILLER_17_169 ();
 sg13g2_fill_1 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_4 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_201 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_fill_2 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_308 ();
 sg13g2_fill_1 FILLER_17_313 ();
 sg13g2_fill_2 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_4 FILLER_17_345 ();
 sg13g2_fill_2 FILLER_17_349 ();
 sg13g2_fill_2 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_fill_2 FILLER_17_394 ();
 sg13g2_fill_1 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_422 ();
 sg13g2_decap_8 FILLER_17_431 ();
 sg13g2_decap_8 FILLER_17_438 ();
 sg13g2_fill_1 FILLER_17_445 ();
 sg13g2_fill_2 FILLER_17_464 ();
 sg13g2_fill_1 FILLER_17_509 ();
 sg13g2_fill_2 FILLER_17_562 ();
 sg13g2_fill_1 FILLER_17_581 ();
 sg13g2_fill_1 FILLER_17_588 ();
 sg13g2_fill_1 FILLER_17_603 ();
 sg13g2_fill_1 FILLER_17_670 ();
 sg13g2_fill_2 FILLER_17_675 ();
 sg13g2_fill_1 FILLER_17_681 ();
 sg13g2_fill_2 FILLER_17_708 ();
 sg13g2_fill_1 FILLER_17_714 ();
 sg13g2_fill_1 FILLER_17_719 ();
 sg13g2_decap_8 FILLER_17_724 ();
 sg13g2_decap_8 FILLER_17_731 ();
 sg13g2_decap_8 FILLER_17_738 ();
 sg13g2_decap_4 FILLER_17_745 ();
 sg13g2_fill_2 FILLER_17_765 ();
 sg13g2_decap_4 FILLER_17_772 ();
 sg13g2_fill_2 FILLER_17_776 ();
 sg13g2_fill_2 FILLER_17_818 ();
 sg13g2_fill_1 FILLER_17_825 ();
 sg13g2_fill_2 FILLER_17_839 ();
 sg13g2_fill_1 FILLER_17_841 ();
 sg13g2_decap_8 FILLER_17_914 ();
 sg13g2_decap_4 FILLER_17_921 ();
 sg13g2_fill_2 FILLER_17_925 ();
 sg13g2_decap_8 FILLER_17_931 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_4 FILLER_17_945 ();
 sg13g2_fill_2 FILLER_17_949 ();
 sg13g2_decap_8 FILLER_17_968 ();
 sg13g2_decap_8 FILLER_17_975 ();
 sg13g2_fill_2 FILLER_17_982 ();
 sg13g2_decap_8 FILLER_17_988 ();
 sg13g2_decap_8 FILLER_17_995 ();
 sg13g2_fill_1 FILLER_17_1002 ();
 sg13g2_fill_2 FILLER_17_1029 ();
 sg13g2_fill_2 FILLER_17_1042 ();
 sg13g2_fill_2 FILLER_17_1053 ();
 sg13g2_fill_2 FILLER_17_1067 ();
 sg13g2_fill_1 FILLER_17_1090 ();
 sg13g2_fill_1 FILLER_17_1147 ();
 sg13g2_fill_1 FILLER_17_1152 ();
 sg13g2_fill_1 FILLER_17_1158 ();
 sg13g2_fill_1 FILLER_17_1163 ();
 sg13g2_fill_1 FILLER_17_1185 ();
 sg13g2_decap_8 FILLER_17_1190 ();
 sg13g2_decap_8 FILLER_17_1197 ();
 sg13g2_decap_4 FILLER_17_1204 ();
 sg13g2_fill_2 FILLER_17_1238 ();
 sg13g2_fill_2 FILLER_17_1245 ();
 sg13g2_decap_4 FILLER_17_1268 ();
 sg13g2_fill_2 FILLER_17_1288 ();
 sg13g2_fill_1 FILLER_17_1290 ();
 sg13g2_decap_8 FILLER_17_1299 ();
 sg13g2_fill_2 FILLER_17_1306 ();
 sg13g2_fill_2 FILLER_17_1338 ();
 sg13g2_fill_1 FILLER_17_1347 ();
 sg13g2_fill_2 FILLER_17_1353 ();
 sg13g2_fill_1 FILLER_17_1359 ();
 sg13g2_fill_1 FILLER_17_1409 ();
 sg13g2_decap_4 FILLER_17_1443 ();
 sg13g2_fill_2 FILLER_17_1447 ();
 sg13g2_fill_1 FILLER_17_1477 ();
 sg13g2_decap_8 FILLER_17_1568 ();
 sg13g2_decap_4 FILLER_17_1575 ();
 sg13g2_fill_1 FILLER_17_1609 ();
 sg13g2_fill_1 FILLER_17_1614 ();
 sg13g2_fill_1 FILLER_17_1620 ();
 sg13g2_fill_1 FILLER_17_1630 ();
 sg13g2_fill_1 FILLER_17_1635 ();
 sg13g2_fill_2 FILLER_17_1676 ();
 sg13g2_fill_1 FILLER_17_1678 ();
 sg13g2_fill_2 FILLER_17_1712 ();
 sg13g2_decap_4 FILLER_17_1737 ();
 sg13g2_fill_1 FILLER_17_1754 ();
 sg13g2_fill_2 FILLER_17_1760 ();
 sg13g2_fill_2 FILLER_17_1775 ();
 sg13g2_fill_1 FILLER_17_1821 ();
 sg13g2_fill_2 FILLER_17_1826 ();
 sg13g2_decap_8 FILLER_17_1832 ();
 sg13g2_decap_4 FILLER_17_1839 ();
 sg13g2_fill_1 FILLER_17_1873 ();
 sg13g2_decap_8 FILLER_17_1883 ();
 sg13g2_decap_4 FILLER_17_1890 ();
 sg13g2_fill_1 FILLER_17_1894 ();
 sg13g2_fill_1 FILLER_17_1898 ();
 sg13g2_fill_1 FILLER_17_1911 ();
 sg13g2_fill_1 FILLER_17_1963 ();
 sg13g2_decap_8 FILLER_17_1969 ();
 sg13g2_fill_2 FILLER_17_1976 ();
 sg13g2_decap_8 FILLER_17_1991 ();
 sg13g2_decap_4 FILLER_17_1998 ();
 sg13g2_decap_8 FILLER_17_2015 ();
 sg13g2_decap_4 FILLER_17_2022 ();
 sg13g2_decap_8 FILLER_17_2034 ();
 sg13g2_decap_8 FILLER_17_2041 ();
 sg13g2_fill_1 FILLER_17_2048 ();
 sg13g2_fill_1 FILLER_17_2062 ();
 sg13g2_decap_8 FILLER_17_2093 ();
 sg13g2_fill_2 FILLER_17_2144 ();
 sg13g2_fill_1 FILLER_17_2146 ();
 sg13g2_decap_8 FILLER_17_2173 ();
 sg13g2_decap_8 FILLER_17_2180 ();
 sg13g2_decap_8 FILLER_17_2187 ();
 sg13g2_fill_1 FILLER_17_2194 ();
 sg13g2_decap_8 FILLER_17_2200 ();
 sg13g2_decap_8 FILLER_17_2207 ();
 sg13g2_decap_4 FILLER_17_2214 ();
 sg13g2_fill_2 FILLER_17_2223 ();
 sg13g2_fill_1 FILLER_17_2225 ();
 sg13g2_fill_1 FILLER_17_2234 ();
 sg13g2_fill_1 FILLER_17_2253 ();
 sg13g2_fill_2 FILLER_17_2280 ();
 sg13g2_fill_1 FILLER_17_2282 ();
 sg13g2_decap_8 FILLER_17_2287 ();
 sg13g2_decap_8 FILLER_17_2294 ();
 sg13g2_decap_4 FILLER_17_2301 ();
 sg13g2_fill_2 FILLER_17_2305 ();
 sg13g2_fill_1 FILLER_17_2323 ();
 sg13g2_fill_2 FILLER_17_2329 ();
 sg13g2_fill_1 FILLER_17_2331 ();
 sg13g2_decap_4 FILLER_17_2337 ();
 sg13g2_decap_8 FILLER_17_2349 ();
 sg13g2_fill_2 FILLER_17_2356 ();
 sg13g2_fill_1 FILLER_17_2358 ();
 sg13g2_fill_2 FILLER_17_2384 ();
 sg13g2_fill_1 FILLER_17_2399 ();
 sg13g2_fill_2 FILLER_17_2418 ();
 sg13g2_decap_4 FILLER_17_2454 ();
 sg13g2_fill_1 FILLER_17_2458 ();
 sg13g2_fill_2 FILLER_17_2464 ();
 sg13g2_fill_2 FILLER_17_2503 ();
 sg13g2_fill_1 FILLER_17_2505 ();
 sg13g2_decap_8 FILLER_17_2510 ();
 sg13g2_decap_4 FILLER_17_2517 ();
 sg13g2_fill_2 FILLER_17_2521 ();
 sg13g2_fill_2 FILLER_17_2528 ();
 sg13g2_fill_2 FILLER_17_2546 ();
 sg13g2_decap_8 FILLER_17_2555 ();
 sg13g2_fill_1 FILLER_17_2562 ();
 sg13g2_fill_1 FILLER_17_2567 ();
 sg13g2_decap_8 FILLER_17_2572 ();
 sg13g2_fill_2 FILLER_17_2579 ();
 sg13g2_fill_1 FILLER_17_2593 ();
 sg13g2_decap_4 FILLER_17_2624 ();
 sg13g2_fill_1 FILLER_17_2628 ();
 sg13g2_decap_8 FILLER_17_2637 ();
 sg13g2_decap_8 FILLER_17_2644 ();
 sg13g2_decap_8 FILLER_17_2651 ();
 sg13g2_decap_8 FILLER_17_2658 ();
 sg13g2_decap_4 FILLER_17_2665 ();
 sg13g2_fill_1 FILLER_17_2669 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_11 ();
 sg13g2_fill_1 FILLER_18_17 ();
 sg13g2_decap_4 FILLER_18_22 ();
 sg13g2_fill_1 FILLER_18_26 ();
 sg13g2_fill_2 FILLER_18_32 ();
 sg13g2_fill_1 FILLER_18_34 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_4 FILLER_18_67 ();
 sg13g2_decap_4 FILLER_18_75 ();
 sg13g2_fill_1 FILLER_18_87 ();
 sg13g2_decap_8 FILLER_18_96 ();
 sg13g2_decap_8 FILLER_18_103 ();
 sg13g2_decap_4 FILLER_18_110 ();
 sg13g2_fill_2 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_164 ();
 sg13g2_fill_1 FILLER_18_191 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_fill_1 FILLER_18_259 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_decap_4 FILLER_18_407 ();
 sg13g2_fill_2 FILLER_18_411 ();
 sg13g2_fill_1 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_536 ();
 sg13g2_decap_4 FILLER_18_543 ();
 sg13g2_fill_1 FILLER_18_547 ();
 sg13g2_fill_2 FILLER_18_580 ();
 sg13g2_fill_1 FILLER_18_648 ();
 sg13g2_fill_2 FILLER_18_653 ();
 sg13g2_fill_1 FILLER_18_660 ();
 sg13g2_decap_8 FILLER_18_704 ();
 sg13g2_decap_8 FILLER_18_711 ();
 sg13g2_decap_4 FILLER_18_718 ();
 sg13g2_fill_1 FILLER_18_722 ();
 sg13g2_decap_8 FILLER_18_727 ();
 sg13g2_fill_2 FILLER_18_734 ();
 sg13g2_fill_1 FILLER_18_736 ();
 sg13g2_fill_2 FILLER_18_762 ();
 sg13g2_decap_4 FILLER_18_775 ();
 sg13g2_fill_1 FILLER_18_779 ();
 sg13g2_fill_1 FILLER_18_814 ();
 sg13g2_fill_2 FILLER_18_846 ();
 sg13g2_fill_1 FILLER_18_848 ();
 sg13g2_fill_2 FILLER_18_875 ();
 sg13g2_fill_2 FILLER_18_946 ();
 sg13g2_fill_1 FILLER_18_948 ();
 sg13g2_decap_4 FILLER_18_953 ();
 sg13g2_fill_2 FILLER_18_983 ();
 sg13g2_fill_1 FILLER_18_985 ();
 sg13g2_fill_1 FILLER_18_992 ();
 sg13g2_fill_2 FILLER_18_1045 ();
 sg13g2_fill_2 FILLER_18_1095 ();
 sg13g2_fill_1 FILLER_18_1097 ();
 sg13g2_fill_1 FILLER_18_1102 ();
 sg13g2_fill_2 FILLER_18_1133 ();
 sg13g2_fill_2 FILLER_18_1147 ();
 sg13g2_fill_1 FILLER_18_1149 ();
 sg13g2_decap_4 FILLER_18_1214 ();
 sg13g2_fill_1 FILLER_18_1235 ();
 sg13g2_fill_2 FILLER_18_1259 ();
 sg13g2_fill_2 FILLER_18_1287 ();
 sg13g2_fill_1 FILLER_18_1289 ();
 sg13g2_fill_1 FILLER_18_1343 ();
 sg13g2_fill_1 FILLER_18_1349 ();
 sg13g2_fill_2 FILLER_18_1354 ();
 sg13g2_fill_1 FILLER_18_1365 ();
 sg13g2_fill_1 FILLER_18_1371 ();
 sg13g2_fill_1 FILLER_18_1377 ();
 sg13g2_fill_1 FILLER_18_1404 ();
 sg13g2_fill_2 FILLER_18_1425 ();
 sg13g2_fill_2 FILLER_18_1431 ();
 sg13g2_fill_1 FILLER_18_1433 ();
 sg13g2_fill_2 FILLER_18_1459 ();
 sg13g2_fill_1 FILLER_18_1488 ();
 sg13g2_decap_8 FILLER_18_1577 ();
 sg13g2_fill_1 FILLER_18_1628 ();
 sg13g2_decap_8 FILLER_18_1663 ();
 sg13g2_decap_4 FILLER_18_1674 ();
 sg13g2_fill_2 FILLER_18_1678 ();
 sg13g2_decap_4 FILLER_18_1701 ();
 sg13g2_fill_1 FILLER_18_1714 ();
 sg13g2_fill_1 FILLER_18_1718 ();
 sg13g2_decap_8 FILLER_18_1732 ();
 sg13g2_fill_1 FILLER_18_1739 ();
 sg13g2_decap_4 FILLER_18_1766 ();
 sg13g2_fill_1 FILLER_18_1770 ();
 sg13g2_decap_8 FILLER_18_1830 ();
 sg13g2_decap_8 FILLER_18_1837 ();
 sg13g2_fill_1 FILLER_18_1844 ();
 sg13g2_fill_2 FILLER_18_1866 ();
 sg13g2_fill_2 FILLER_18_1916 ();
 sg13g2_fill_2 FILLER_18_1969 ();
 sg13g2_fill_1 FILLER_18_1975 ();
 sg13g2_decap_8 FILLER_18_2006 ();
 sg13g2_fill_1 FILLER_18_2013 ();
 sg13g2_fill_2 FILLER_18_2019 ();
 sg13g2_decap_8 FILLER_18_2095 ();
 sg13g2_fill_2 FILLER_18_2102 ();
 sg13g2_fill_1 FILLER_18_2104 ();
 sg13g2_decap_8 FILLER_18_2160 ();
 sg13g2_fill_2 FILLER_18_2167 ();
 sg13g2_fill_1 FILLER_18_2169 ();
 sg13g2_fill_2 FILLER_18_2174 ();
 sg13g2_decap_8 FILLER_18_2192 ();
 sg13g2_fill_1 FILLER_18_2199 ();
 sg13g2_fill_1 FILLER_18_2221 ();
 sg13g2_fill_1 FILLER_18_2251 ();
 sg13g2_fill_1 FILLER_18_2286 ();
 sg13g2_fill_2 FILLER_18_2344 ();
 sg13g2_fill_1 FILLER_18_2346 ();
 sg13g2_decap_8 FILLER_18_2368 ();
 sg13g2_fill_2 FILLER_18_2375 ();
 sg13g2_fill_2 FILLER_18_2431 ();
 sg13g2_fill_1 FILLER_18_2438 ();
 sg13g2_decap_8 FILLER_18_2443 ();
 sg13g2_decap_8 FILLER_18_2450 ();
 sg13g2_decap_8 FILLER_18_2457 ();
 sg13g2_decap_8 FILLER_18_2464 ();
 sg13g2_fill_2 FILLER_18_2471 ();
 sg13g2_fill_1 FILLER_18_2487 ();
 sg13g2_decap_8 FILLER_18_2492 ();
 sg13g2_decap_8 FILLER_18_2499 ();
 sg13g2_decap_4 FILLER_18_2506 ();
 sg13g2_fill_2 FILLER_18_2510 ();
 sg13g2_fill_2 FILLER_18_2517 ();
 sg13g2_decap_8 FILLER_18_2523 ();
 sg13g2_decap_8 FILLER_18_2530 ();
 sg13g2_decap_4 FILLER_18_2537 ();
 sg13g2_decap_4 FILLER_18_2556 ();
 sg13g2_decap_8 FILLER_18_2568 ();
 sg13g2_fill_2 FILLER_18_2575 ();
 sg13g2_decap_4 FILLER_18_2582 ();
 sg13g2_decap_4 FILLER_18_2590 ();
 sg13g2_fill_2 FILLER_18_2594 ();
 sg13g2_fill_1 FILLER_18_2600 ();
 sg13g2_decap_8 FILLER_18_2627 ();
 sg13g2_decap_8 FILLER_18_2634 ();
 sg13g2_decap_8 FILLER_18_2641 ();
 sg13g2_decap_8 FILLER_18_2648 ();
 sg13g2_decap_8 FILLER_18_2655 ();
 sg13g2_decap_8 FILLER_18_2662 ();
 sg13g2_fill_1 FILLER_18_2669 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_6 ();
 sg13g2_fill_1 FILLER_19_8 ();
 sg13g2_fill_2 FILLER_19_13 ();
 sg13g2_fill_1 FILLER_19_15 ();
 sg13g2_fill_2 FILLER_19_42 ();
 sg13g2_fill_1 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_118 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_fill_2 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_215 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_294 ();
 sg13g2_fill_2 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_350 ();
 sg13g2_fill_2 FILLER_19_390 ();
 sg13g2_fill_1 FILLER_19_418 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_fill_2 FILLER_19_503 ();
 sg13g2_fill_1 FILLER_19_567 ();
 sg13g2_fill_2 FILLER_19_572 ();
 sg13g2_fill_2 FILLER_19_588 ();
 sg13g2_decap_4 FILLER_19_630 ();
 sg13g2_decap_4 FILLER_19_647 ();
 sg13g2_fill_1 FILLER_19_664 ();
 sg13g2_fill_1 FILLER_19_706 ();
 sg13g2_decap_4 FILLER_19_783 ();
 sg13g2_fill_2 FILLER_19_787 ();
 sg13g2_fill_2 FILLER_19_806 ();
 sg13g2_fill_1 FILLER_19_812 ();
 sg13g2_fill_1 FILLER_19_822 ();
 sg13g2_fill_1 FILLER_19_827 ();
 sg13g2_fill_1 FILLER_19_841 ();
 sg13g2_fill_2 FILLER_19_863 ();
 sg13g2_fill_1 FILLER_19_869 ();
 sg13g2_fill_2 FILLER_19_874 ();
 sg13g2_decap_4 FILLER_19_885 ();
 sg13g2_fill_1 FILLER_19_889 ();
 sg13g2_fill_2 FILLER_19_894 ();
 sg13g2_fill_1 FILLER_19_896 ();
 sg13g2_decap_4 FILLER_19_901 ();
 sg13g2_fill_2 FILLER_19_905 ();
 sg13g2_fill_1 FILLER_19_915 ();
 sg13g2_fill_1 FILLER_19_925 ();
 sg13g2_fill_1 FILLER_19_930 ();
 sg13g2_fill_2 FILLER_19_948 ();
 sg13g2_fill_2 FILLER_19_981 ();
 sg13g2_fill_1 FILLER_19_995 ();
 sg13g2_fill_1 FILLER_19_1032 ();
 sg13g2_fill_1 FILLER_19_1054 ();
 sg13g2_decap_4 FILLER_19_1121 ();
 sg13g2_fill_1 FILLER_19_1125 ();
 sg13g2_fill_2 FILLER_19_1130 ();
 sg13g2_decap_4 FILLER_19_1162 ();
 sg13g2_decap_8 FILLER_19_1201 ();
 sg13g2_decap_8 FILLER_19_1208 ();
 sg13g2_decap_4 FILLER_19_1215 ();
 sg13g2_fill_1 FILLER_19_1219 ();
 sg13g2_fill_1 FILLER_19_1224 ();
 sg13g2_fill_2 FILLER_19_1325 ();
 sg13g2_decap_8 FILLER_19_1353 ();
 sg13g2_fill_1 FILLER_19_1360 ();
 sg13g2_fill_2 FILLER_19_1366 ();
 sg13g2_fill_1 FILLER_19_1372 ();
 sg13g2_fill_1 FILLER_19_1385 ();
 sg13g2_fill_1 FILLER_19_1427 ();
 sg13g2_fill_2 FILLER_19_1465 ();
 sg13g2_fill_2 FILLER_19_1494 ();
 sg13g2_fill_2 FILLER_19_1543 ();
 sg13g2_fill_1 FILLER_19_1545 ();
 sg13g2_decap_4 FILLER_19_1559 ();
 sg13g2_fill_2 FILLER_19_1563 ();
 sg13g2_fill_2 FILLER_19_1626 ();
 sg13g2_fill_1 FILLER_19_1628 ();
 sg13g2_fill_1 FILLER_19_1634 ();
 sg13g2_decap_8 FILLER_19_1639 ();
 sg13g2_decap_8 FILLER_19_1676 ();
 sg13g2_decap_4 FILLER_19_1687 ();
 sg13g2_fill_2 FILLER_19_1691 ();
 sg13g2_decap_8 FILLER_19_1697 ();
 sg13g2_fill_1 FILLER_19_1704 ();
 sg13g2_fill_1 FILLER_19_1708 ();
 sg13g2_fill_2 FILLER_19_1823 ();
 sg13g2_fill_1 FILLER_19_1825 ();
 sg13g2_fill_2 FILLER_19_1830 ();
 sg13g2_fill_2 FILLER_19_1858 ();
 sg13g2_fill_1 FILLER_19_1898 ();
 sg13g2_fill_2 FILLER_19_1902 ();
 sg13g2_fill_2 FILLER_19_1952 ();
 sg13g2_fill_2 FILLER_19_1964 ();
 sg13g2_fill_2 FILLER_19_2014 ();
 sg13g2_fill_1 FILLER_19_2016 ();
 sg13g2_fill_1 FILLER_19_2022 ();
 sg13g2_fill_2 FILLER_19_2027 ();
 sg13g2_fill_2 FILLER_19_2110 ();
 sg13g2_fill_1 FILLER_19_2112 ();
 sg13g2_fill_2 FILLER_19_2141 ();
 sg13g2_fill_1 FILLER_19_2143 ();
 sg13g2_fill_2 FILLER_19_2215 ();
 sg13g2_decap_8 FILLER_19_2227 ();
 sg13g2_decap_8 FILLER_19_2234 ();
 sg13g2_fill_2 FILLER_19_2241 ();
 sg13g2_fill_1 FILLER_19_2247 ();
 sg13g2_fill_2 FILLER_19_2254 ();
 sg13g2_fill_2 FILLER_19_2271 ();
 sg13g2_fill_1 FILLER_19_2278 ();
 sg13g2_decap_4 FILLER_19_2307 ();
 sg13g2_fill_1 FILLER_19_2319 ();
 sg13g2_decap_8 FILLER_19_2324 ();
 sg13g2_decap_4 FILLER_19_2331 ();
 sg13g2_fill_2 FILLER_19_2335 ();
 sg13g2_fill_2 FILLER_19_2342 ();
 sg13g2_fill_2 FILLER_19_2349 ();
 sg13g2_decap_8 FILLER_19_2372 ();
 sg13g2_decap_8 FILLER_19_2379 ();
 sg13g2_fill_1 FILLER_19_2386 ();
 sg13g2_fill_2 FILLER_19_2396 ();
 sg13g2_decap_4 FILLER_19_2402 ();
 sg13g2_decap_8 FILLER_19_2438 ();
 sg13g2_decap_8 FILLER_19_2445 ();
 sg13g2_decap_8 FILLER_19_2452 ();
 sg13g2_fill_2 FILLER_19_2459 ();
 sg13g2_fill_1 FILLER_19_2461 ();
 sg13g2_decap_4 FILLER_19_2494 ();
 sg13g2_fill_2 FILLER_19_2502 ();
 sg13g2_fill_1 FILLER_19_2504 ();
 sg13g2_decap_4 FILLER_19_2509 ();
 sg13g2_fill_1 FILLER_19_2513 ();
 sg13g2_decap_4 FILLER_19_2584 ();
 sg13g2_fill_1 FILLER_19_2588 ();
 sg13g2_decap_4 FILLER_19_2594 ();
 sg13g2_fill_2 FILLER_19_2610 ();
 sg13g2_fill_2 FILLER_19_2617 ();
 sg13g2_decap_8 FILLER_19_2645 ();
 sg13g2_decap_8 FILLER_19_2652 ();
 sg13g2_decap_8 FILLER_19_2659 ();
 sg13g2_decap_4 FILLER_19_2666 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_32 ();
 sg13g2_fill_1 FILLER_20_37 ();
 sg13g2_fill_1 FILLER_20_69 ();
 sg13g2_fill_2 FILLER_20_83 ();
 sg13g2_fill_1 FILLER_20_166 ();
 sg13g2_fill_2 FILLER_20_181 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_decap_4 FILLER_20_268 ();
 sg13g2_fill_2 FILLER_20_272 ();
 sg13g2_fill_2 FILLER_20_291 ();
 sg13g2_fill_1 FILLER_20_293 ();
 sg13g2_fill_2 FILLER_20_298 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_374 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_413 ();
 sg13g2_fill_2 FILLER_20_440 ();
 sg13g2_fill_1 FILLER_20_491 ();
 sg13g2_fill_2 FILLER_20_536 ();
 sg13g2_fill_1 FILLER_20_546 ();
 sg13g2_fill_1 FILLER_20_552 ();
 sg13g2_fill_2 FILLER_20_566 ();
 sg13g2_fill_1 FILLER_20_577 ();
 sg13g2_fill_1 FILLER_20_602 ();
 sg13g2_fill_2 FILLER_20_607 ();
 sg13g2_fill_1 FILLER_20_613 ();
 sg13g2_fill_1 FILLER_20_622 ();
 sg13g2_decap_8 FILLER_20_627 ();
 sg13g2_decap_4 FILLER_20_634 ();
 sg13g2_fill_2 FILLER_20_638 ();
 sg13g2_fill_2 FILLER_20_669 ();
 sg13g2_fill_2 FILLER_20_675 ();
 sg13g2_fill_2 FILLER_20_681 ();
 sg13g2_fill_1 FILLER_20_687 ();
 sg13g2_fill_1 FILLER_20_698 ();
 sg13g2_fill_2 FILLER_20_737 ();
 sg13g2_fill_1 FILLER_20_758 ();
 sg13g2_fill_1 FILLER_20_801 ();
 sg13g2_fill_1 FILLER_20_806 ();
 sg13g2_fill_1 FILLER_20_813 ();
 sg13g2_fill_2 FILLER_20_896 ();
 sg13g2_fill_1 FILLER_20_898 ();
 sg13g2_fill_1 FILLER_20_903 ();
 sg13g2_fill_1 FILLER_20_912 ();
 sg13g2_fill_1 FILLER_20_918 ();
 sg13g2_fill_2 FILLER_20_924 ();
 sg13g2_fill_2 FILLER_20_949 ();
 sg13g2_fill_2 FILLER_20_982 ();
 sg13g2_fill_1 FILLER_20_1042 ();
 sg13g2_fill_2 FILLER_20_1060 ();
 sg13g2_decap_8 FILLER_20_1075 ();
 sg13g2_fill_2 FILLER_20_1109 ();
 sg13g2_decap_4 FILLER_20_1181 ();
 sg13g2_fill_1 FILLER_20_1185 ();
 sg13g2_fill_2 FILLER_20_1196 ();
 sg13g2_fill_1 FILLER_20_1220 ();
 sg13g2_fill_1 FILLER_20_1225 ();
 sg13g2_fill_2 FILLER_20_1231 ();
 sg13g2_decap_4 FILLER_20_1271 ();
 sg13g2_fill_2 FILLER_20_1275 ();
 sg13g2_decap_4 FILLER_20_1307 ();
 sg13g2_fill_2 FILLER_20_1311 ();
 sg13g2_decap_8 FILLER_20_1348 ();
 sg13g2_decap_8 FILLER_20_1355 ();
 sg13g2_decap_8 FILLER_20_1362 ();
 sg13g2_decap_4 FILLER_20_1369 ();
 sg13g2_fill_1 FILLER_20_1373 ();
 sg13g2_decap_4 FILLER_20_1378 ();
 sg13g2_fill_1 FILLER_20_1398 ();
 sg13g2_fill_1 FILLER_20_1435 ();
 sg13g2_fill_2 FILLER_20_1441 ();
 sg13g2_fill_2 FILLER_20_1461 ();
 sg13g2_fill_1 FILLER_20_1477 ();
 sg13g2_fill_1 FILLER_20_1527 ();
 sg13g2_fill_2 FILLER_20_1536 ();
 sg13g2_decap_4 FILLER_20_1553 ();
 sg13g2_fill_2 FILLER_20_1557 ();
 sg13g2_fill_2 FILLER_20_1607 ();
 sg13g2_fill_1 FILLER_20_1609 ();
 sg13g2_fill_1 FILLER_20_1614 ();
 sg13g2_decap_8 FILLER_20_1620 ();
 sg13g2_decap_8 FILLER_20_1627 ();
 sg13g2_fill_1 FILLER_20_1634 ();
 sg13g2_fill_1 FILLER_20_1683 ();
 sg13g2_fill_2 FILLER_20_1718 ();
 sg13g2_fill_1 FILLER_20_1723 ();
 sg13g2_fill_2 FILLER_20_1728 ();
 sg13g2_fill_1 FILLER_20_1734 ();
 sg13g2_fill_1 FILLER_20_1739 ();
 sg13g2_fill_1 FILLER_20_1766 ();
 sg13g2_fill_1 FILLER_20_1779 ();
 sg13g2_fill_2 FILLER_20_1788 ();
 sg13g2_fill_2 FILLER_20_1798 ();
 sg13g2_fill_1 FILLER_20_1807 ();
 sg13g2_fill_1 FILLER_20_1859 ();
 sg13g2_fill_2 FILLER_20_1908 ();
 sg13g2_fill_1 FILLER_20_1928 ();
 sg13g2_fill_1 FILLER_20_1974 ();
 sg13g2_fill_1 FILLER_20_1984 ();
 sg13g2_fill_1 FILLER_20_1993 ();
 sg13g2_decap_8 FILLER_20_2050 ();
 sg13g2_decap_8 FILLER_20_2057 ();
 sg13g2_fill_1 FILLER_20_2064 ();
 sg13g2_fill_1 FILLER_20_2069 ();
 sg13g2_decap_8 FILLER_20_2153 ();
 sg13g2_decap_8 FILLER_20_2164 ();
 sg13g2_fill_2 FILLER_20_2171 ();
 sg13g2_fill_2 FILLER_20_2219 ();
 sg13g2_fill_1 FILLER_20_2225 ();
 sg13g2_fill_2 FILLER_20_2252 ();
 sg13g2_fill_1 FILLER_20_2263 ();
 sg13g2_decap_8 FILLER_20_2324 ();
 sg13g2_decap_4 FILLER_20_2331 ();
 sg13g2_fill_1 FILLER_20_2335 ();
 sg13g2_decap_8 FILLER_20_2341 ();
 sg13g2_fill_1 FILLER_20_2348 ();
 sg13g2_decap_8 FILLER_20_2375 ();
 sg13g2_fill_2 FILLER_20_2382 ();
 sg13g2_decap_8 FILLER_20_2392 ();
 sg13g2_decap_8 FILLER_20_2399 ();
 sg13g2_fill_1 FILLER_20_2427 ();
 sg13g2_fill_1 FILLER_20_2480 ();
 sg13g2_decap_8 FILLER_20_2538 ();
 sg13g2_decap_8 FILLER_20_2545 ();
 sg13g2_fill_1 FILLER_20_2552 ();
 sg13g2_fill_1 FILLER_20_2571 ();
 sg13g2_fill_1 FILLER_20_2575 ();
 sg13g2_fill_1 FILLER_20_2608 ();
 sg13g2_fill_2 FILLER_20_2622 ();
 sg13g2_fill_1 FILLER_20_2624 ();
 sg13g2_fill_1 FILLER_20_2655 ();
 sg13g2_decap_8 FILLER_20_2660 ();
 sg13g2_fill_2 FILLER_20_2667 ();
 sg13g2_fill_1 FILLER_20_2669 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_59 ();
 sg13g2_fill_2 FILLER_21_65 ();
 sg13g2_decap_8 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_1 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_fill_2 FILLER_21_304 ();
 sg13g2_fill_1 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_404 ();
 sg13g2_fill_2 FILLER_21_430 ();
 sg13g2_fill_2 FILLER_21_441 ();
 sg13g2_fill_1 FILLER_21_479 ();
 sg13g2_decap_4 FILLER_21_485 ();
 sg13g2_fill_1 FILLER_21_489 ();
 sg13g2_fill_2 FILLER_21_508 ();
 sg13g2_fill_2 FILLER_21_518 ();
 sg13g2_fill_1 FILLER_21_617 ();
 sg13g2_decap_8 FILLER_21_627 ();
 sg13g2_fill_2 FILLER_21_660 ();
 sg13g2_fill_1 FILLER_21_662 ();
 sg13g2_fill_1 FILLER_21_699 ();
 sg13g2_fill_2 FILLER_21_721 ();
 sg13g2_fill_2 FILLER_21_731 ();
 sg13g2_fill_1 FILLER_21_749 ();
 sg13g2_fill_1 FILLER_21_763 ();
 sg13g2_fill_1 FILLER_21_787 ();
 sg13g2_decap_4 FILLER_21_800 ();
 sg13g2_fill_1 FILLER_21_811 ();
 sg13g2_fill_1 FILLER_21_859 ();
 sg13g2_fill_2 FILLER_21_865 ();
 sg13g2_fill_2 FILLER_21_871 ();
 sg13g2_decap_4 FILLER_21_899 ();
 sg13g2_fill_2 FILLER_21_903 ();
 sg13g2_decap_4 FILLER_21_974 ();
 sg13g2_fill_2 FILLER_21_978 ();
 sg13g2_decap_4 FILLER_21_1000 ();
 sg13g2_fill_1 FILLER_21_1013 ();
 sg13g2_fill_2 FILLER_21_1017 ();
 sg13g2_fill_1 FILLER_21_1045 ();
 sg13g2_fill_1 FILLER_21_1070 ();
 sg13g2_fill_1 FILLER_21_1076 ();
 sg13g2_fill_2 FILLER_21_1089 ();
 sg13g2_fill_2 FILLER_21_1104 ();
 sg13g2_fill_2 FILLER_21_1111 ();
 sg13g2_fill_1 FILLER_21_1113 ();
 sg13g2_fill_2 FILLER_21_1118 ();
 sg13g2_decap_8 FILLER_21_1124 ();
 sg13g2_decap_8 FILLER_21_1131 ();
 sg13g2_fill_2 FILLER_21_1138 ();
 sg13g2_fill_2 FILLER_21_1191 ();
 sg13g2_fill_1 FILLER_21_1193 ();
 sg13g2_decap_4 FILLER_21_1202 ();
 sg13g2_fill_2 FILLER_21_1230 ();
 sg13g2_decap_4 FILLER_21_1236 ();
 sg13g2_fill_1 FILLER_21_1254 ();
 sg13g2_fill_1 FILLER_21_1258 ();
 sg13g2_decap_4 FILLER_21_1266 ();
 sg13g2_fill_2 FILLER_21_1270 ();
 sg13g2_fill_1 FILLER_21_1278 ();
 sg13g2_decap_4 FILLER_21_1323 ();
 sg13g2_fill_1 FILLER_21_1327 ();
 sg13g2_decap_8 FILLER_21_1332 ();
 sg13g2_decap_8 FILLER_21_1339 ();
 sg13g2_fill_2 FILLER_21_1346 ();
 sg13g2_decap_8 FILLER_21_1352 ();
 sg13g2_decap_4 FILLER_21_1359 ();
 sg13g2_fill_1 FILLER_21_1363 ();
 sg13g2_fill_1 FILLER_21_1383 ();
 sg13g2_fill_2 FILLER_21_1389 ();
 sg13g2_fill_2 FILLER_21_1406 ();
 sg13g2_fill_1 FILLER_21_1413 ();
 sg13g2_fill_2 FILLER_21_1423 ();
 sg13g2_fill_1 FILLER_21_1439 ();
 sg13g2_fill_2 FILLER_21_1471 ();
 sg13g2_fill_2 FILLER_21_1478 ();
 sg13g2_fill_1 FILLER_21_1480 ();
 sg13g2_fill_1 FILLER_21_1513 ();
 sg13g2_decap_8 FILLER_21_1550 ();
 sg13g2_decap_8 FILLER_21_1557 ();
 sg13g2_decap_8 FILLER_21_1564 ();
 sg13g2_fill_1 FILLER_21_1571 ();
 sg13g2_fill_1 FILLER_21_1576 ();
 sg13g2_fill_2 FILLER_21_1598 ();
 sg13g2_decap_4 FILLER_21_1625 ();
 sg13g2_fill_1 FILLER_21_1629 ();
 sg13g2_fill_2 FILLER_21_1633 ();
 sg13g2_fill_1 FILLER_21_1635 ();
 sg13g2_fill_1 FILLER_21_1640 ();
 sg13g2_fill_2 FILLER_21_1646 ();
 sg13g2_fill_1 FILLER_21_1669 ();
 sg13g2_fill_1 FILLER_21_1687 ();
 sg13g2_fill_2 FILLER_21_1721 ();
 sg13g2_fill_1 FILLER_21_1748 ();
 sg13g2_fill_2 FILLER_21_1754 ();
 sg13g2_decap_8 FILLER_21_1836 ();
 sg13g2_decap_8 FILLER_21_1843 ();
 sg13g2_fill_2 FILLER_21_1882 ();
 sg13g2_fill_1 FILLER_21_1910 ();
 sg13g2_fill_1 FILLER_21_1940 ();
 sg13g2_decap_8 FILLER_21_1989 ();
 sg13g2_decap_4 FILLER_21_1996 ();
 sg13g2_fill_1 FILLER_21_2007 ();
 sg13g2_fill_1 FILLER_21_2025 ();
 sg13g2_decap_8 FILLER_21_2043 ();
 sg13g2_decap_8 FILLER_21_2050 ();
 sg13g2_decap_8 FILLER_21_2057 ();
 sg13g2_decap_8 FILLER_21_2064 ();
 sg13g2_decap_4 FILLER_21_2071 ();
 sg13g2_fill_1 FILLER_21_2075 ();
 sg13g2_fill_2 FILLER_21_2080 ();
 sg13g2_decap_8 FILLER_21_2086 ();
 sg13g2_decap_4 FILLER_21_2093 ();
 sg13g2_fill_1 FILLER_21_2097 ();
 sg13g2_fill_1 FILLER_21_2107 ();
 sg13g2_fill_1 FILLER_21_2112 ();
 sg13g2_fill_1 FILLER_21_2117 ();
 sg13g2_fill_1 FILLER_21_2122 ();
 sg13g2_fill_1 FILLER_21_2148 ();
 sg13g2_decap_4 FILLER_21_2184 ();
 sg13g2_fill_2 FILLER_21_2215 ();
 sg13g2_decap_8 FILLER_21_2224 ();
 sg13g2_fill_2 FILLER_21_2231 ();
 sg13g2_fill_1 FILLER_21_2251 ();
 sg13g2_fill_2 FILLER_21_2283 ();
 sg13g2_decap_8 FILLER_21_2324 ();
 sg13g2_fill_2 FILLER_21_2331 ();
 sg13g2_fill_2 FILLER_21_2347 ();
 sg13g2_fill_1 FILLER_21_2349 ();
 sg13g2_fill_1 FILLER_21_2378 ();
 sg13g2_fill_1 FILLER_21_2481 ();
 sg13g2_decap_8 FILLER_21_2549 ();
 sg13g2_fill_1 FILLER_21_2583 ();
 sg13g2_decap_8 FILLER_21_2647 ();
 sg13g2_decap_8 FILLER_21_2654 ();
 sg13g2_decap_8 FILLER_21_2661 ();
 sg13g2_fill_2 FILLER_21_2668 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_decap_4 FILLER_22_13 ();
 sg13g2_fill_2 FILLER_22_21 ();
 sg13g2_decap_4 FILLER_22_27 ();
 sg13g2_fill_1 FILLER_22_31 ();
 sg13g2_decap_8 FILLER_22_36 ();
 sg13g2_fill_2 FILLER_22_43 ();
 sg13g2_decap_4 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_57 ();
 sg13g2_fill_2 FILLER_22_75 ();
 sg13g2_decap_8 FILLER_22_94 ();
 sg13g2_decap_8 FILLER_22_101 ();
 sg13g2_decap_8 FILLER_22_108 ();
 sg13g2_decap_4 FILLER_22_115 ();
 sg13g2_fill_2 FILLER_22_119 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_fill_1 FILLER_22_157 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_257 ();
 sg13g2_decap_4 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_fill_2 FILLER_22_329 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_22_412 ();
 sg13g2_decap_4 FILLER_22_419 ();
 sg13g2_fill_2 FILLER_22_423 ();
 sg13g2_fill_1 FILLER_22_442 ();
 sg13g2_fill_2 FILLER_22_460 ();
 sg13g2_decap_4 FILLER_22_474 ();
 sg13g2_decap_8 FILLER_22_482 ();
 sg13g2_fill_2 FILLER_22_489 ();
 sg13g2_fill_2 FILLER_22_495 ();
 sg13g2_decap_8 FILLER_22_557 ();
 sg13g2_fill_2 FILLER_22_607 ();
 sg13g2_fill_1 FILLER_22_670 ();
 sg13g2_decap_8 FILLER_22_680 ();
 sg13g2_fill_1 FILLER_22_687 ();
 sg13g2_fill_2 FILLER_22_698 ();
 sg13g2_fill_2 FILLER_22_709 ();
 sg13g2_fill_1 FILLER_22_721 ();
 sg13g2_fill_2 FILLER_22_739 ();
 sg13g2_fill_1 FILLER_22_748 ();
 sg13g2_fill_1 FILLER_22_753 ();
 sg13g2_fill_1 FILLER_22_759 ();
 sg13g2_decap_8 FILLER_22_807 ();
 sg13g2_decap_8 FILLER_22_814 ();
 sg13g2_fill_2 FILLER_22_821 ();
 sg13g2_fill_1 FILLER_22_823 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_decap_4 FILLER_22_861 ();
 sg13g2_fill_2 FILLER_22_865 ();
 sg13g2_decap_8 FILLER_22_884 ();
 sg13g2_decap_8 FILLER_22_891 ();
 sg13g2_decap_4 FILLER_22_898 ();
 sg13g2_fill_1 FILLER_22_902 ();
 sg13g2_fill_1 FILLER_22_950 ();
 sg13g2_decap_8 FILLER_22_955 ();
 sg13g2_decap_8 FILLER_22_962 ();
 sg13g2_decap_8 FILLER_22_969 ();
 sg13g2_decap_8 FILLER_22_976 ();
 sg13g2_decap_8 FILLER_22_983 ();
 sg13g2_fill_1 FILLER_22_990 ();
 sg13g2_decap_8 FILLER_22_995 ();
 sg13g2_fill_1 FILLER_22_1010 ();
 sg13g2_fill_1 FILLER_22_1030 ();
 sg13g2_fill_2 FILLER_22_1079 ();
 sg13g2_fill_1 FILLER_22_1081 ();
 sg13g2_decap_4 FILLER_22_1120 ();
 sg13g2_fill_1 FILLER_22_1124 ();
 sg13g2_decap_8 FILLER_22_1129 ();
 sg13g2_decap_8 FILLER_22_1136 ();
 sg13g2_decap_8 FILLER_22_1143 ();
 sg13g2_fill_1 FILLER_22_1150 ();
 sg13g2_decap_4 FILLER_22_1185 ();
 sg13g2_fill_1 FILLER_22_1189 ();
 sg13g2_decap_8 FILLER_22_1206 ();
 sg13g2_fill_2 FILLER_22_1273 ();
 sg13g2_fill_2 FILLER_22_1295 ();
 sg13g2_fill_1 FILLER_22_1297 ();
 sg13g2_decap_4 FILLER_22_1336 ();
 sg13g2_fill_2 FILLER_22_1340 ();
 sg13g2_fill_2 FILLER_22_1368 ();
 sg13g2_fill_1 FILLER_22_1462 ();
 sg13g2_fill_1 FILLER_22_1468 ();
 sg13g2_fill_1 FILLER_22_1473 ();
 sg13g2_fill_2 FILLER_22_1478 ();
 sg13g2_fill_1 FILLER_22_1506 ();
 sg13g2_decap_8 FILLER_22_1554 ();
 sg13g2_decap_8 FILLER_22_1561 ();
 sg13g2_decap_8 FILLER_22_1568 ();
 sg13g2_fill_1 FILLER_22_1575 ();
 sg13g2_fill_2 FILLER_22_1692 ();
 sg13g2_fill_1 FILLER_22_1729 ();
 sg13g2_fill_1 FILLER_22_1738 ();
 sg13g2_fill_1 FILLER_22_1744 ();
 sg13g2_fill_2 FILLER_22_1748 ();
 sg13g2_fill_2 FILLER_22_1764 ();
 sg13g2_fill_1 FILLER_22_1771 ();
 sg13g2_fill_1 FILLER_22_1819 ();
 sg13g2_fill_2 FILLER_22_1864 ();
 sg13g2_fill_1 FILLER_22_1866 ();
 sg13g2_decap_8 FILLER_22_1883 ();
 sg13g2_fill_1 FILLER_22_1890 ();
 sg13g2_decap_8 FILLER_22_1895 ();
 sg13g2_decap_4 FILLER_22_1902 ();
 sg13g2_fill_1 FILLER_22_1906 ();
 sg13g2_fill_1 FILLER_22_1918 ();
 sg13g2_fill_2 FILLER_22_1967 ();
 sg13g2_fill_2 FILLER_22_1999 ();
 sg13g2_decap_8 FILLER_22_2032 ();
 sg13g2_decap_8 FILLER_22_2039 ();
 sg13g2_decap_8 FILLER_22_2046 ();
 sg13g2_decap_4 FILLER_22_2053 ();
 sg13g2_fill_2 FILLER_22_2057 ();
 sg13g2_fill_2 FILLER_22_2076 ();
 sg13g2_decap_8 FILLER_22_2099 ();
 sg13g2_decap_8 FILLER_22_2106 ();
 sg13g2_decap_8 FILLER_22_2113 ();
 sg13g2_decap_8 FILLER_22_2124 ();
 sg13g2_decap_4 FILLER_22_2131 ();
 sg13g2_fill_2 FILLER_22_2135 ();
 sg13g2_decap_8 FILLER_22_2141 ();
 sg13g2_decap_4 FILLER_22_2148 ();
 sg13g2_decap_8 FILLER_22_2165 ();
 sg13g2_decap_8 FILLER_22_2172 ();
 sg13g2_decap_4 FILLER_22_2179 ();
 sg13g2_fill_2 FILLER_22_2213 ();
 sg13g2_decap_8 FILLER_22_2230 ();
 sg13g2_decap_4 FILLER_22_2237 ();
 sg13g2_fill_1 FILLER_22_2241 ();
 sg13g2_decap_4 FILLER_22_2254 ();
 sg13g2_fill_1 FILLER_22_2258 ();
 sg13g2_fill_1 FILLER_22_2277 ();
 sg13g2_decap_4 FILLER_22_2282 ();
 sg13g2_fill_1 FILLER_22_2286 ();
 sg13g2_fill_1 FILLER_22_2292 ();
 sg13g2_fill_1 FILLER_22_2408 ();
 sg13g2_fill_2 FILLER_22_2413 ();
 sg13g2_fill_1 FILLER_22_2415 ();
 sg13g2_decap_8 FILLER_22_2452 ();
 sg13g2_fill_2 FILLER_22_2459 ();
 sg13g2_fill_1 FILLER_22_2470 ();
 sg13g2_decap_8 FILLER_22_2503 ();
 sg13g2_fill_1 FILLER_22_2510 ();
 sg13g2_fill_1 FILLER_22_2517 ();
 sg13g2_fill_2 FILLER_22_2539 ();
 sg13g2_fill_1 FILLER_22_2541 ();
 sg13g2_decap_4 FILLER_22_2559 ();
 sg13g2_fill_1 FILLER_22_2563 ();
 sg13g2_fill_1 FILLER_22_2571 ();
 sg13g2_decap_8 FILLER_22_2618 ();
 sg13g2_fill_2 FILLER_22_2625 ();
 sg13g2_fill_1 FILLER_22_2627 ();
 sg13g2_decap_4 FILLER_22_2632 ();
 sg13g2_decap_8 FILLER_22_2662 ();
 sg13g2_fill_1 FILLER_22_2669 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_46 ();
 sg13g2_fill_2 FILLER_23_61 ();
 sg13g2_decap_8 FILLER_23_101 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_121 ();
 sg13g2_fill_2 FILLER_23_152 ();
 sg13g2_fill_1 FILLER_23_159 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_231 ();
 sg13g2_decap_4 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_263 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_323 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_fill_1 FILLER_23_341 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_1 FILLER_23_417 ();
 sg13g2_decap_4 FILLER_23_431 ();
 sg13g2_fill_1 FILLER_23_458 ();
 sg13g2_fill_1 FILLER_23_505 ();
 sg13g2_fill_1 FILLER_23_511 ();
 sg13g2_fill_1 FILLER_23_517 ();
 sg13g2_fill_2 FILLER_23_544 ();
 sg13g2_fill_1 FILLER_23_567 ();
 sg13g2_fill_2 FILLER_23_573 ();
 sg13g2_fill_1 FILLER_23_575 ();
 sg13g2_fill_1 FILLER_23_588 ();
 sg13g2_fill_1 FILLER_23_627 ();
 sg13g2_fill_2 FILLER_23_641 ();
 sg13g2_fill_1 FILLER_23_643 ();
 sg13g2_fill_2 FILLER_23_740 ();
 sg13g2_fill_2 FILLER_23_754 ();
 sg13g2_fill_1 FILLER_23_759 ();
 sg13g2_fill_1 FILLER_23_768 ();
 sg13g2_fill_1 FILLER_23_804 ();
 sg13g2_fill_1 FILLER_23_809 ();
 sg13g2_decap_8 FILLER_23_814 ();
 sg13g2_decap_8 FILLER_23_821 ();
 sg13g2_decap_4 FILLER_23_828 ();
 sg13g2_fill_2 FILLER_23_832 ();
 sg13g2_decap_8 FILLER_23_844 ();
 sg13g2_decap_8 FILLER_23_851 ();
 sg13g2_decap_8 FILLER_23_858 ();
 sg13g2_decap_8 FILLER_23_865 ();
 sg13g2_decap_4 FILLER_23_872 ();
 sg13g2_fill_1 FILLER_23_876 ();
 sg13g2_decap_8 FILLER_23_894 ();
 sg13g2_decap_8 FILLER_23_901 ();
 sg13g2_decap_4 FILLER_23_908 ();
 sg13g2_fill_1 FILLER_23_912 ();
 sg13g2_decap_4 FILLER_23_939 ();
 sg13g2_fill_1 FILLER_23_956 ();
 sg13g2_fill_2 FILLER_23_996 ();
 sg13g2_fill_1 FILLER_23_998 ();
 sg13g2_decap_8 FILLER_23_1032 ();
 sg13g2_decap_8 FILLER_23_1074 ();
 sg13g2_fill_1 FILLER_23_1081 ();
 sg13g2_fill_1 FILLER_23_1186 ();
 sg13g2_fill_2 FILLER_23_1295 ();
 sg13g2_fill_1 FILLER_23_1311 ();
 sg13g2_fill_1 FILLER_23_1375 ();
 sg13g2_fill_1 FILLER_23_1381 ();
 sg13g2_fill_1 FILLER_23_1386 ();
 sg13g2_fill_1 FILLER_23_1392 ();
 sg13g2_fill_2 FILLER_23_1423 ();
 sg13g2_fill_2 FILLER_23_1467 ();
 sg13g2_fill_1 FILLER_23_1478 ();
 sg13g2_decap_8 FILLER_23_1573 ();
 sg13g2_decap_4 FILLER_23_1580 ();
 sg13g2_fill_1 FILLER_23_1584 ();
 sg13g2_decap_4 FILLER_23_1589 ();
 sg13g2_fill_1 FILLER_23_1602 ();
 sg13g2_fill_2 FILLER_23_1607 ();
 sg13g2_fill_1 FILLER_23_1613 ();
 sg13g2_fill_2 FILLER_23_1627 ();
 sg13g2_fill_2 FILLER_23_1646 ();
 sg13g2_fill_1 FILLER_23_1688 ();
 sg13g2_fill_1 FILLER_23_1719 ();
 sg13g2_fill_1 FILLER_23_1724 ();
 sg13g2_fill_1 FILLER_23_1739 ();
 sg13g2_fill_1 FILLER_23_1744 ();
 sg13g2_fill_1 FILLER_23_1749 ();
 sg13g2_fill_2 FILLER_23_1754 ();
 sg13g2_fill_1 FILLER_23_1765 ();
 sg13g2_fill_1 FILLER_23_1792 ();
 sg13g2_fill_2 FILLER_23_1827 ();
 sg13g2_decap_8 FILLER_23_1833 ();
 sg13g2_fill_2 FILLER_23_1840 ();
 sg13g2_fill_1 FILLER_23_1842 ();
 sg13g2_decap_4 FILLER_23_1864 ();
 sg13g2_fill_1 FILLER_23_1868 ();
 sg13g2_fill_2 FILLER_23_1881 ();
 sg13g2_fill_1 FILLER_23_1883 ();
 sg13g2_decap_8 FILLER_23_1888 ();
 sg13g2_decap_8 FILLER_23_1895 ();
 sg13g2_decap_4 FILLER_23_1902 ();
 sg13g2_fill_1 FILLER_23_1911 ();
 sg13g2_decap_8 FILLER_23_1994 ();
 sg13g2_decap_8 FILLER_23_2018 ();
 sg13g2_decap_8 FILLER_23_2025 ();
 sg13g2_decap_4 FILLER_23_2032 ();
 sg13g2_fill_2 FILLER_23_2036 ();
 sg13g2_fill_2 FILLER_23_2046 ();
 sg13g2_fill_1 FILLER_23_2048 ();
 sg13g2_fill_1 FILLER_23_2054 ();
 sg13g2_fill_1 FILLER_23_2085 ();
 sg13g2_fill_2 FILLER_23_2137 ();
 sg13g2_decap_8 FILLER_23_2143 ();
 sg13g2_decap_8 FILLER_23_2150 ();
 sg13g2_decap_4 FILLER_23_2157 ();
 sg13g2_fill_2 FILLER_23_2161 ();
 sg13g2_fill_1 FILLER_23_2220 ();
 sg13g2_fill_1 FILLER_23_2229 ();
 sg13g2_fill_2 FILLER_23_2234 ();
 sg13g2_decap_4 FILLER_23_2266 ();
 sg13g2_fill_1 FILLER_23_2270 ();
 sg13g2_fill_2 FILLER_23_2288 ();
 sg13g2_fill_2 FILLER_23_2304 ();
 sg13g2_fill_1 FILLER_23_2336 ();
 sg13g2_decap_4 FILLER_23_2355 ();
 sg13g2_fill_1 FILLER_23_2359 ();
 sg13g2_fill_2 FILLER_23_2372 ();
 sg13g2_decap_4 FILLER_23_2383 ();
 sg13g2_fill_1 FILLER_23_2420 ();
 sg13g2_fill_1 FILLER_23_2426 ();
 sg13g2_decap_8 FILLER_23_2441 ();
 sg13g2_decap_8 FILLER_23_2448 ();
 sg13g2_decap_4 FILLER_23_2455 ();
 sg13g2_fill_2 FILLER_23_2459 ();
 sg13g2_fill_1 FILLER_23_2471 ();
 sg13g2_fill_2 FILLER_23_2477 ();
 sg13g2_decap_4 FILLER_23_2483 ();
 sg13g2_fill_1 FILLER_23_2487 ();
 sg13g2_decap_8 FILLER_23_2493 ();
 sg13g2_decap_4 FILLER_23_2500 ();
 sg13g2_fill_2 FILLER_23_2504 ();
 sg13g2_decap_4 FILLER_23_2539 ();
 sg13g2_fill_2 FILLER_23_2551 ();
 sg13g2_fill_1 FILLER_23_2553 ();
 sg13g2_fill_1 FILLER_23_2558 ();
 sg13g2_fill_2 FILLER_23_2575 ();
 sg13g2_fill_2 FILLER_23_2585 ();
 sg13g2_decap_4 FILLER_23_2624 ();
 sg13g2_fill_1 FILLER_23_2628 ();
 sg13g2_fill_2 FILLER_23_2641 ();
 sg13g2_fill_1 FILLER_23_2643 ();
 sg13g2_fill_2 FILLER_23_2648 ();
 sg13g2_fill_1 FILLER_23_2650 ();
 sg13g2_decap_4 FILLER_23_2664 ();
 sg13g2_fill_2 FILLER_23_2668 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_33 ();
 sg13g2_fill_1 FILLER_24_41 ();
 sg13g2_fill_1 FILLER_24_68 ();
 sg13g2_fill_2 FILLER_24_118 ();
 sg13g2_fill_1 FILLER_24_120 ();
 sg13g2_fill_2 FILLER_24_151 ();
 sg13g2_decap_4 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_222 ();
 sg13g2_fill_2 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_357 ();
 sg13g2_fill_1 FILLER_24_362 ();
 sg13g2_fill_1 FILLER_24_367 ();
 sg13g2_fill_2 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_24_379 ();
 sg13g2_fill_1 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_533 ();
 sg13g2_fill_2 FILLER_24_540 ();
 sg13g2_fill_1 FILLER_24_542 ();
 sg13g2_decap_8 FILLER_24_564 ();
 sg13g2_decap_8 FILLER_24_571 ();
 sg13g2_decap_8 FILLER_24_578 ();
 sg13g2_fill_2 FILLER_24_585 ();
 sg13g2_fill_1 FILLER_24_587 ();
 sg13g2_fill_1 FILLER_24_613 ();
 sg13g2_fill_2 FILLER_24_622 ();
 sg13g2_fill_1 FILLER_24_624 ();
 sg13g2_fill_2 FILLER_24_638 ();
 sg13g2_fill_1 FILLER_24_640 ();
 sg13g2_decap_8 FILLER_24_682 ();
 sg13g2_decap_4 FILLER_24_689 ();
 sg13g2_fill_2 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_fill_2 FILLER_24_707 ();
 sg13g2_fill_1 FILLER_24_709 ();
 sg13g2_fill_2 FILLER_24_745 ();
 sg13g2_fill_1 FILLER_24_763 ();
 sg13g2_fill_2 FILLER_24_782 ();
 sg13g2_fill_1 FILLER_24_788 ();
 sg13g2_fill_1 FILLER_24_793 ();
 sg13g2_fill_1 FILLER_24_803 ();
 sg13g2_fill_1 FILLER_24_830 ();
 sg13g2_decap_8 FILLER_24_852 ();
 sg13g2_decap_4 FILLER_24_859 ();
 sg13g2_fill_1 FILLER_24_863 ();
 sg13g2_fill_1 FILLER_24_873 ();
 sg13g2_fill_1 FILLER_24_878 ();
 sg13g2_decap_8 FILLER_24_909 ();
 sg13g2_fill_2 FILLER_24_916 ();
 sg13g2_fill_1 FILLER_24_918 ();
 sg13g2_decap_8 FILLER_24_927 ();
 sg13g2_fill_2 FILLER_24_934 ();
 sg13g2_fill_1 FILLER_24_936 ();
 sg13g2_decap_4 FILLER_24_963 ();
 sg13g2_fill_2 FILLER_24_967 ();
 sg13g2_fill_2 FILLER_24_973 ();
 sg13g2_decap_8 FILLER_24_1031 ();
 sg13g2_decap_4 FILLER_24_1038 ();
 sg13g2_decap_4 FILLER_24_1105 ();
 sg13g2_fill_2 FILLER_24_1109 ();
 sg13g2_decap_8 FILLER_24_1146 ();
 sg13g2_decap_8 FILLER_24_1179 ();
 sg13g2_decap_4 FILLER_24_1186 ();
 sg13g2_fill_2 FILLER_24_1190 ();
 sg13g2_fill_1 FILLER_24_1228 ();
 sg13g2_fill_2 FILLER_24_1233 ();
 sg13g2_fill_1 FILLER_24_1243 ();
 sg13g2_fill_1 FILLER_24_1310 ();
 sg13g2_fill_1 FILLER_24_1316 ();
 sg13g2_fill_2 FILLER_24_1320 ();
 sg13g2_fill_2 FILLER_24_1348 ();
 sg13g2_fill_1 FILLER_24_1380 ();
 sg13g2_fill_2 FILLER_24_1389 ();
 sg13g2_fill_1 FILLER_24_1406 ();
 sg13g2_decap_4 FILLER_24_1416 ();
 sg13g2_fill_1 FILLER_24_1436 ();
 sg13g2_fill_2 FILLER_24_1441 ();
 sg13g2_fill_1 FILLER_24_1443 ();
 sg13g2_fill_2 FILLER_24_1462 ();
 sg13g2_fill_1 FILLER_24_1464 ();
 sg13g2_fill_2 FILLER_24_1483 ();
 sg13g2_fill_1 FILLER_24_1485 ();
 sg13g2_fill_2 FILLER_24_1494 ();
 sg13g2_fill_1 FILLER_24_1500 ();
 sg13g2_fill_1 FILLER_24_1508 ();
 sg13g2_fill_2 FILLER_24_1530 ();
 sg13g2_decap_8 FILLER_24_1558 ();
 sg13g2_fill_1 FILLER_24_1565 ();
 sg13g2_decap_8 FILLER_24_1587 ();
 sg13g2_fill_2 FILLER_24_1594 ();
 sg13g2_fill_1 FILLER_24_1596 ();
 sg13g2_fill_2 FILLER_24_1666 ();
 sg13g2_fill_1 FILLER_24_1682 ();
 sg13g2_fill_1 FILLER_24_1688 ();
 sg13g2_fill_2 FILLER_24_1715 ();
 sg13g2_fill_2 FILLER_24_1747 ();
 sg13g2_decap_8 FILLER_24_1810 ();
 sg13g2_fill_2 FILLER_24_1817 ();
 sg13g2_decap_8 FILLER_24_1823 ();
 sg13g2_decap_8 FILLER_24_1830 ();
 sg13g2_fill_1 FILLER_24_1837 ();
 sg13g2_fill_2 FILLER_24_1841 ();
 sg13g2_decap_4 FILLER_24_1899 ();
 sg13g2_fill_2 FILLER_24_1903 ();
 sg13g2_fill_2 FILLER_24_1915 ();
 sg13g2_fill_2 FILLER_24_1922 ();
 sg13g2_fill_2 FILLER_24_1931 ();
 sg13g2_fill_1 FILLER_24_1937 ();
 sg13g2_fill_1 FILLER_24_1965 ();
 sg13g2_decap_4 FILLER_24_1984 ();
 sg13g2_fill_2 FILLER_24_1988 ();
 sg13g2_fill_2 FILLER_24_2060 ();
 sg13g2_decap_4 FILLER_24_2083 ();
 sg13g2_decap_4 FILLER_24_2113 ();
 sg13g2_decap_4 FILLER_24_2152 ();
 sg13g2_fill_1 FILLER_24_2156 ();
 sg13g2_fill_2 FILLER_24_2193 ();
 sg13g2_fill_1 FILLER_24_2200 ();
 sg13g2_fill_1 FILLER_24_2285 ();
 sg13g2_decap_4 FILLER_24_2343 ();
 sg13g2_fill_1 FILLER_24_2347 ();
 sg13g2_fill_1 FILLER_24_2372 ();
 sg13g2_fill_1 FILLER_24_2378 ();
 sg13g2_decap_8 FILLER_24_2427 ();
 sg13g2_fill_1 FILLER_24_2434 ();
 sg13g2_decap_4 FILLER_24_2440 ();
 sg13g2_fill_1 FILLER_24_2444 ();
 sg13g2_decap_8 FILLER_24_2485 ();
 sg13g2_decap_8 FILLER_24_2492 ();
 sg13g2_decap_4 FILLER_24_2499 ();
 sg13g2_decap_4 FILLER_24_2597 ();
 sg13g2_fill_1 FILLER_24_2601 ();
 sg13g2_fill_2 FILLER_24_2654 ();
 sg13g2_fill_1 FILLER_24_2656 ();
 sg13g2_decap_8 FILLER_24_2661 ();
 sg13g2_fill_2 FILLER_24_2668 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_69 ();
 sg13g2_fill_1 FILLER_25_71 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_4 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_256 ();
 sg13g2_decap_4 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_decap_4 FILLER_25_300 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_4 FILLER_25_372 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_2 FILLER_25_473 ();
 sg13g2_fill_1 FILLER_25_475 ();
 sg13g2_fill_2 FILLER_25_507 ();
 sg13g2_decap_8 FILLER_25_517 ();
 sg13g2_decap_8 FILLER_25_524 ();
 sg13g2_decap_8 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_559 ();
 sg13g2_decap_4 FILLER_25_566 ();
 sg13g2_fill_1 FILLER_25_570 ();
 sg13g2_decap_4 FILLER_25_575 ();
 sg13g2_fill_2 FILLER_25_579 ();
 sg13g2_fill_1 FILLER_25_615 ();
 sg13g2_fill_1 FILLER_25_637 ();
 sg13g2_fill_1 FILLER_25_659 ();
 sg13g2_fill_1 FILLER_25_665 ();
 sg13g2_fill_2 FILLER_25_670 ();
 sg13g2_fill_2 FILLER_25_803 ();
 sg13g2_fill_1 FILLER_25_831 ();
 sg13g2_fill_2 FILLER_25_890 ();
 sg13g2_fill_1 FILLER_25_892 ();
 sg13g2_decap_4 FILLER_25_902 ();
 sg13g2_fill_2 FILLER_25_911 ();
 sg13g2_fill_1 FILLER_25_913 ();
 sg13g2_fill_1 FILLER_25_922 ();
 sg13g2_fill_2 FILLER_25_941 ();
 sg13g2_decap_4 FILLER_25_1033 ();
 sg13g2_decap_4 FILLER_25_1042 ();
 sg13g2_fill_1 FILLER_25_1085 ();
 sg13g2_fill_2 FILLER_25_1090 ();
 sg13g2_fill_1 FILLER_25_1092 ();
 sg13g2_decap_8 FILLER_25_1101 ();
 sg13g2_fill_2 FILLER_25_1108 ();
 sg13g2_fill_1 FILLER_25_1110 ();
 sg13g2_fill_1 FILLER_25_1145 ();
 sg13g2_decap_8 FILLER_25_1150 ();
 sg13g2_fill_1 FILLER_25_1157 ();
 sg13g2_decap_8 FILLER_25_1162 ();
 sg13g2_fill_1 FILLER_25_1169 ();
 sg13g2_fill_1 FILLER_25_1205 ();
 sg13g2_decap_4 FILLER_25_1211 ();
 sg13g2_fill_1 FILLER_25_1215 ();
 sg13g2_fill_1 FILLER_25_1268 ();
 sg13g2_fill_2 FILLER_25_1295 ();
 sg13g2_fill_2 FILLER_25_1307 ();
 sg13g2_fill_1 FILLER_25_1313 ();
 sg13g2_fill_2 FILLER_25_1339 ();
 sg13g2_fill_1 FILLER_25_1341 ();
 sg13g2_decap_8 FILLER_25_1350 ();
 sg13g2_fill_1 FILLER_25_1357 ();
 sg13g2_decap_4 FILLER_25_1362 ();
 sg13g2_fill_1 FILLER_25_1366 ();
 sg13g2_fill_1 FILLER_25_1372 ();
 sg13g2_decap_4 FILLER_25_1377 ();
 sg13g2_decap_8 FILLER_25_1394 ();
 sg13g2_fill_1 FILLER_25_1401 ();
 sg13g2_decap_4 FILLER_25_1406 ();
 sg13g2_fill_2 FILLER_25_1419 ();
 sg13g2_fill_1 FILLER_25_1421 ();
 sg13g2_fill_2 FILLER_25_1439 ();
 sg13g2_fill_2 FILLER_25_1450 ();
 sg13g2_decap_4 FILLER_25_1457 ();
 sg13g2_fill_1 FILLER_25_1468 ();
 sg13g2_decap_8 FILLER_25_1473 ();
 sg13g2_decap_4 FILLER_25_1480 ();
 sg13g2_fill_1 FILLER_25_1484 ();
 sg13g2_decap_8 FILLER_25_1489 ();
 sg13g2_fill_1 FILLER_25_1496 ();
 sg13g2_fill_2 FILLER_25_1540 ();
 sg13g2_fill_1 FILLER_25_1542 ();
 sg13g2_decap_8 FILLER_25_1547 ();
 sg13g2_fill_2 FILLER_25_1563 ();
 sg13g2_fill_1 FILLER_25_1565 ();
 sg13g2_fill_2 FILLER_25_1591 ();
 sg13g2_fill_2 FILLER_25_1597 ();
 sg13g2_fill_1 FILLER_25_1603 ();
 sg13g2_fill_1 FILLER_25_1686 ();
 sg13g2_fill_1 FILLER_25_1715 ();
 sg13g2_decap_8 FILLER_25_1806 ();
 sg13g2_decap_8 FILLER_25_1813 ();
 sg13g2_fill_2 FILLER_25_1820 ();
 sg13g2_decap_4 FILLER_25_1826 ();
 sg13g2_fill_2 FILLER_25_1834 ();
 sg13g2_fill_1 FILLER_25_1861 ();
 sg13g2_fill_1 FILLER_25_1928 ();
 sg13g2_fill_1 FILLER_25_1944 ();
 sg13g2_decap_8 FILLER_25_1976 ();
 sg13g2_decap_4 FILLER_25_1983 ();
 sg13g2_fill_1 FILLER_25_2004 ();
 sg13g2_fill_2 FILLER_25_2010 ();
 sg13g2_fill_1 FILLER_25_2103 ();
 sg13g2_fill_2 FILLER_25_2125 ();
 sg13g2_fill_2 FILLER_25_2132 ();
 sg13g2_fill_1 FILLER_25_2160 ();
 sg13g2_fill_2 FILLER_25_2185 ();
 sg13g2_fill_1 FILLER_25_2199 ();
 sg13g2_fill_2 FILLER_25_2244 ();
 sg13g2_fill_1 FILLER_25_2246 ();
 sg13g2_fill_2 FILLER_25_2279 ();
 sg13g2_decap_8 FILLER_25_2324 ();
 sg13g2_decap_8 FILLER_25_2331 ();
 sg13g2_decap_4 FILLER_25_2338 ();
 sg13g2_decap_4 FILLER_25_2351 ();
 sg13g2_fill_2 FILLER_25_2380 ();
 sg13g2_decap_4 FILLER_25_2397 ();
 sg13g2_decap_4 FILLER_25_2410 ();
 sg13g2_fill_1 FILLER_25_2414 ();
 sg13g2_decap_8 FILLER_25_2419 ();
 sg13g2_fill_2 FILLER_25_2426 ();
 sg13g2_fill_1 FILLER_25_2428 ();
 sg13g2_fill_2 FILLER_25_2433 ();
 sg13g2_fill_1 FILLER_25_2439 ();
 sg13g2_fill_1 FILLER_25_2448 ();
 sg13g2_fill_1 FILLER_25_2478 ();
 sg13g2_decap_8 FILLER_25_2482 ();
 sg13g2_decap_4 FILLER_25_2489 ();
 sg13g2_fill_1 FILLER_25_2519 ();
 sg13g2_decap_4 FILLER_25_2524 ();
 sg13g2_fill_1 FILLER_25_2528 ();
 sg13g2_fill_1 FILLER_25_2535 ();
 sg13g2_decap_4 FILLER_25_2565 ();
 sg13g2_decap_4 FILLER_25_2581 ();
 sg13g2_fill_2 FILLER_25_2585 ();
 sg13g2_fill_2 FILLER_25_2602 ();
 sg13g2_fill_1 FILLER_25_2604 ();
 sg13g2_decap_4 FILLER_25_2634 ();
 sg13g2_decap_8 FILLER_25_2642 ();
 sg13g2_fill_1 FILLER_25_2649 ();
 sg13g2_decap_8 FILLER_25_2654 ();
 sg13g2_decap_8 FILLER_25_2661 ();
 sg13g2_fill_2 FILLER_25_2668 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_58 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_79 ();
 sg13g2_fill_2 FILLER_26_101 ();
 sg13g2_fill_1 FILLER_26_103 ();
 sg13g2_decap_8 FILLER_26_108 ();
 sg13g2_decap_8 FILLER_26_115 ();
 sg13g2_decap_8 FILLER_26_122 ();
 sg13g2_decap_4 FILLER_26_129 ();
 sg13g2_decap_4 FILLER_26_137 ();
 sg13g2_fill_1 FILLER_26_141 ();
 sg13g2_fill_2 FILLER_26_156 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_decap_4 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_225 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_fill_1 FILLER_26_240 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_4 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_293 ();
 sg13g2_decap_4 FILLER_26_303 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_fill_2 FILLER_26_313 ();
 sg13g2_fill_1 FILLER_26_315 ();
 sg13g2_fill_1 FILLER_26_321 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_fill_1 FILLER_26_379 ();
 sg13g2_decap_4 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_393 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_fill_2 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_26_410 ();
 sg13g2_decap_4 FILLER_26_514 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_fill_2 FILLER_26_590 ();
 sg13g2_fill_1 FILLER_26_597 ();
 sg13g2_fill_1 FILLER_26_602 ();
 sg13g2_fill_1 FILLER_26_608 ();
 sg13g2_fill_1 FILLER_26_613 ();
 sg13g2_fill_2 FILLER_26_667 ();
 sg13g2_fill_1 FILLER_26_669 ();
 sg13g2_decap_8 FILLER_26_696 ();
 sg13g2_decap_8 FILLER_26_703 ();
 sg13g2_fill_2 FILLER_26_710 ();
 sg13g2_decap_4 FILLER_26_721 ();
 sg13g2_decap_4 FILLER_26_729 ();
 sg13g2_fill_1 FILLER_26_733 ();
 sg13g2_fill_2 FILLER_26_738 ();
 sg13g2_fill_2 FILLER_26_783 ();
 sg13g2_fill_1 FILLER_26_785 ();
 sg13g2_fill_1 FILLER_26_794 ();
 sg13g2_fill_1 FILLER_26_799 ();
 sg13g2_fill_2 FILLER_26_805 ();
 sg13g2_fill_1 FILLER_26_807 ();
 sg13g2_fill_2 FILLER_26_812 ();
 sg13g2_fill_1 FILLER_26_862 ();
 sg13g2_fill_1 FILLER_26_868 ();
 sg13g2_fill_1 FILLER_26_899 ();
 sg13g2_decap_8 FILLER_26_934 ();
 sg13g2_fill_1 FILLER_26_949 ();
 sg13g2_fill_2 FILLER_26_959 ();
 sg13g2_fill_1 FILLER_26_961 ();
 sg13g2_decap_8 FILLER_26_972 ();
 sg13g2_decap_4 FILLER_26_979 ();
 sg13g2_fill_2 FILLER_26_987 ();
 sg13g2_fill_1 FILLER_26_1016 ();
 sg13g2_fill_2 FILLER_26_1043 ();
 sg13g2_fill_1 FILLER_26_1045 ();
 sg13g2_decap_8 FILLER_26_1072 ();
 sg13g2_decap_4 FILLER_26_1083 ();
 sg13g2_decap_8 FILLER_26_1091 ();
 sg13g2_decap_4 FILLER_26_1102 ();
 sg13g2_fill_1 FILLER_26_1132 ();
 sg13g2_fill_2 FILLER_26_1138 ();
 sg13g2_fill_1 FILLER_26_1140 ();
 sg13g2_fill_2 FILLER_26_1167 ();
 sg13g2_fill_1 FILLER_26_1169 ();
 sg13g2_fill_2 FILLER_26_1273 ();
 sg13g2_fill_1 FILLER_26_1278 ();
 sg13g2_fill_1 FILLER_26_1284 ();
 sg13g2_fill_2 FILLER_26_1334 ();
 sg13g2_fill_1 FILLER_26_1336 ();
 sg13g2_decap_8 FILLER_26_1341 ();
 sg13g2_fill_1 FILLER_26_1358 ();
 sg13g2_fill_1 FILLER_26_1363 ();
 sg13g2_fill_2 FILLER_26_1424 ();
 sg13g2_fill_1 FILLER_26_1426 ();
 sg13g2_fill_2 FILLER_26_1437 ();
 sg13g2_fill_1 FILLER_26_1465 ();
 sg13g2_fill_1 FILLER_26_1471 ();
 sg13g2_decap_8 FILLER_26_1476 ();
 sg13g2_fill_1 FILLER_26_1483 ();
 sg13g2_fill_2 FILLER_26_1493 ();
 sg13g2_fill_1 FILLER_26_1495 ();
 sg13g2_decap_4 FILLER_26_1543 ();
 sg13g2_fill_1 FILLER_26_1547 ();
 sg13g2_fill_1 FILLER_26_1613 ();
 sg13g2_fill_2 FILLER_26_1623 ();
 sg13g2_fill_2 FILLER_26_1649 ();
 sg13g2_fill_1 FILLER_26_1658 ();
 sg13g2_decap_8 FILLER_26_1685 ();
 sg13g2_decap_4 FILLER_26_1692 ();
 sg13g2_fill_1 FILLER_26_1696 ();
 sg13g2_decap_8 FILLER_26_1701 ();
 sg13g2_fill_1 FILLER_26_1708 ();
 sg13g2_decap_8 FILLER_26_1714 ();
 sg13g2_fill_2 FILLER_26_1721 ();
 sg13g2_fill_2 FILLER_26_1762 ();
 sg13g2_fill_1 FILLER_26_1773 ();
 sg13g2_fill_2 FILLER_26_1795 ();
 sg13g2_fill_1 FILLER_26_1871 ();
 sg13g2_fill_2 FILLER_26_1925 ();
 sg13g2_fill_1 FILLER_26_1927 ();
 sg13g2_decap_4 FILLER_26_1932 ();
 sg13g2_decap_8 FILLER_26_1973 ();
 sg13g2_decap_4 FILLER_26_2056 ();
 sg13g2_fill_2 FILLER_26_2091 ();
 sg13g2_fill_1 FILLER_26_2093 ();
 sg13g2_fill_1 FILLER_26_2120 ();
 sg13g2_fill_1 FILLER_26_2130 ();
 sg13g2_decap_4 FILLER_26_2157 ();
 sg13g2_decap_8 FILLER_26_2170 ();
 sg13g2_decap_8 FILLER_26_2177 ();
 sg13g2_fill_2 FILLER_26_2184 ();
 sg13g2_fill_1 FILLER_26_2204 ();
 sg13g2_fill_1 FILLER_26_2210 ();
 sg13g2_fill_1 FILLER_26_2215 ();
 sg13g2_fill_2 FILLER_26_2221 ();
 sg13g2_fill_2 FILLER_26_2231 ();
 sg13g2_fill_1 FILLER_26_2233 ();
 sg13g2_fill_1 FILLER_26_2239 ();
 sg13g2_fill_2 FILLER_26_2248 ();
 sg13g2_decap_4 FILLER_26_2276 ();
 sg13g2_decap_8 FILLER_26_2318 ();
 sg13g2_decap_8 FILLER_26_2325 ();
 sg13g2_fill_1 FILLER_26_2332 ();
 sg13g2_fill_2 FILLER_26_2345 ();
 sg13g2_fill_1 FILLER_26_2347 ();
 sg13g2_fill_2 FILLER_26_2391 ();
 sg13g2_fill_2 FILLER_26_2398 ();
 sg13g2_decap_8 FILLER_26_2410 ();
 sg13g2_decap_8 FILLER_26_2417 ();
 sg13g2_fill_2 FILLER_26_2432 ();
 sg13g2_fill_2 FILLER_26_2471 ();
 sg13g2_decap_8 FILLER_26_2478 ();
 sg13g2_fill_2 FILLER_26_2495 ();
 sg13g2_fill_1 FILLER_26_2497 ();
 sg13g2_fill_1 FILLER_26_2505 ();
 sg13g2_fill_1 FILLER_26_2511 ();
 sg13g2_fill_1 FILLER_26_2516 ();
 sg13g2_fill_2 FILLER_26_2522 ();
 sg13g2_decap_4 FILLER_26_2532 ();
 sg13g2_decap_4 FILLER_26_2545 ();
 sg13g2_decap_4 FILLER_26_2557 ();
 sg13g2_fill_2 FILLER_26_2573 ();
 sg13g2_decap_4 FILLER_26_2610 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_11 ();
 sg13g2_decap_8 FILLER_27_16 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_33 ();
 sg13g2_fill_2 FILLER_27_43 ();
 sg13g2_fill_2 FILLER_27_54 ();
 sg13g2_fill_1 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_113 ();
 sg13g2_decap_8 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_157 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_178 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_decap_4 FILLER_27_271 ();
 sg13g2_fill_2 FILLER_27_275 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_fill_2 FILLER_27_400 ();
 sg13g2_fill_1 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_27_413 ();
 sg13g2_fill_1 FILLER_27_417 ();
 sg13g2_fill_1 FILLER_27_431 ();
 sg13g2_fill_1 FILLER_27_469 ();
 sg13g2_fill_2 FILLER_27_485 ();
 sg13g2_fill_1 FILLER_27_538 ();
 sg13g2_fill_1 FILLER_27_577 ();
 sg13g2_fill_1 FILLER_27_596 ();
 sg13g2_fill_1 FILLER_27_601 ();
 sg13g2_fill_1 FILLER_27_628 ();
 sg13g2_fill_2 FILLER_27_659 ();
 sg13g2_decap_8 FILLER_27_691 ();
 sg13g2_decap_4 FILLER_27_698 ();
 sg13g2_decap_8 FILLER_27_706 ();
 sg13g2_fill_2 FILLER_27_713 ();
 sg13g2_decap_4 FILLER_27_719 ();
 sg13g2_fill_2 FILLER_27_753 ();
 sg13g2_fill_1 FILLER_27_762 ();
 sg13g2_fill_1 FILLER_27_798 ();
 sg13g2_fill_1 FILLER_27_829 ();
 sg13g2_fill_2 FILLER_27_872 ();
 sg13g2_decap_8 FILLER_27_949 ();
 sg13g2_decap_4 FILLER_27_956 ();
 sg13g2_fill_2 FILLER_27_960 ();
 sg13g2_fill_1 FILLER_27_966 ();
 sg13g2_fill_2 FILLER_27_971 ();
 sg13g2_fill_2 FILLER_27_977 ();
 sg13g2_fill_1 FILLER_27_987 ();
 sg13g2_decap_4 FILLER_27_992 ();
 sg13g2_fill_2 FILLER_27_996 ();
 sg13g2_fill_2 FILLER_27_1020 ();
 sg13g2_fill_1 FILLER_27_1030 ();
 sg13g2_fill_2 FILLER_27_1035 ();
 sg13g2_fill_2 FILLER_27_1041 ();
 sg13g2_fill_1 FILLER_27_1073 ();
 sg13g2_fill_1 FILLER_27_1105 ();
 sg13g2_decap_8 FILLER_27_1152 ();
 sg13g2_decap_8 FILLER_27_1159 ();
 sg13g2_fill_1 FILLER_27_1166 ();
 sg13g2_decap_8 FILLER_27_1170 ();
 sg13g2_fill_2 FILLER_27_1177 ();
 sg13g2_fill_1 FILLER_27_1179 ();
 sg13g2_decap_4 FILLER_27_1184 ();
 sg13g2_decap_4 FILLER_27_1191 ();
 sg13g2_fill_1 FILLER_27_1215 ();
 sg13g2_fill_2 FILLER_27_1242 ();
 sg13g2_fill_2 FILLER_27_1257 ();
 sg13g2_fill_1 FILLER_27_1283 ();
 sg13g2_fill_1 FILLER_27_1317 ();
 sg13g2_fill_2 FILLER_27_1385 ();
 sg13g2_fill_1 FILLER_27_1387 ();
 sg13g2_fill_2 FILLER_27_1432 ();
 sg13g2_fill_1 FILLER_27_1434 ();
 sg13g2_fill_1 FILLER_27_1490 ();
 sg13g2_fill_1 FILLER_27_1517 ();
 sg13g2_fill_2 FILLER_27_1568 ();
 sg13g2_fill_2 FILLER_27_1580 ();
 sg13g2_fill_1 FILLER_27_1597 ();
 sg13g2_fill_1 FILLER_27_1601 ();
 sg13g2_fill_1 FILLER_27_1607 ();
 sg13g2_fill_1 FILLER_27_1653 ();
 sg13g2_decap_4 FILLER_27_1690 ();
 sg13g2_fill_1 FILLER_27_1694 ();
 sg13g2_fill_1 FILLER_27_1700 ();
 sg13g2_decap_4 FILLER_27_1709 ();
 sg13g2_fill_1 FILLER_27_1713 ();
 sg13g2_decap_8 FILLER_27_1718 ();
 sg13g2_decap_8 FILLER_27_1742 ();
 sg13g2_decap_8 FILLER_27_1749 ();
 sg13g2_decap_8 FILLER_27_1756 ();
 sg13g2_decap_8 FILLER_27_1763 ();
 sg13g2_fill_2 FILLER_27_1770 ();
 sg13g2_fill_1 FILLER_27_1772 ();
 sg13g2_decap_8 FILLER_27_1780 ();
 sg13g2_decap_4 FILLER_27_1787 ();
 sg13g2_fill_1 FILLER_27_1791 ();
 sg13g2_fill_2 FILLER_27_1860 ();
 sg13g2_fill_1 FILLER_27_1880 ();
 sg13g2_decap_4 FILLER_27_1918 ();
 sg13g2_fill_2 FILLER_27_2013 ();
 sg13g2_fill_1 FILLER_27_2015 ();
 sg13g2_decap_4 FILLER_27_2025 ();
 sg13g2_fill_2 FILLER_27_2037 ();
 sg13g2_fill_1 FILLER_27_2039 ();
 sg13g2_fill_1 FILLER_27_2044 ();
 sg13g2_fill_2 FILLER_27_2126 ();
 sg13g2_decap_8 FILLER_27_2154 ();
 sg13g2_decap_8 FILLER_27_2161 ();
 sg13g2_decap_8 FILLER_27_2168 ();
 sg13g2_fill_2 FILLER_27_2188 ();
 sg13g2_fill_1 FILLER_27_2190 ();
 sg13g2_fill_2 FILLER_27_2208 ();
 sg13g2_decap_4 FILLER_27_2218 ();
 sg13g2_fill_1 FILLER_27_2222 ();
 sg13g2_decap_8 FILLER_27_2239 ();
 sg13g2_fill_2 FILLER_27_2251 ();
 sg13g2_decap_4 FILLER_27_2258 ();
 sg13g2_fill_1 FILLER_27_2262 ();
 sg13g2_decap_4 FILLER_27_2283 ();
 sg13g2_fill_1 FILLER_27_2300 ();
 sg13g2_decap_4 FILLER_27_2306 ();
 sg13g2_decap_4 FILLER_27_2314 ();
 sg13g2_fill_2 FILLER_27_2322 ();
 sg13g2_fill_1 FILLER_27_2324 ();
 sg13g2_fill_2 FILLER_27_2343 ();
 sg13g2_fill_2 FILLER_27_2375 ();
 sg13g2_decap_8 FILLER_27_2402 ();
 sg13g2_fill_1 FILLER_27_2409 ();
 sg13g2_decap_4 FILLER_27_2420 ();
 sg13g2_fill_1 FILLER_27_2424 ();
 sg13g2_decap_4 FILLER_27_2430 ();
 sg13g2_fill_1 FILLER_27_2486 ();
 sg13g2_fill_2 FILLER_27_2499 ();
 sg13g2_fill_1 FILLER_27_2506 ();
 sg13g2_fill_1 FILLER_27_2523 ();
 sg13g2_fill_1 FILLER_27_2529 ();
 sg13g2_fill_1 FILLER_27_2536 ();
 sg13g2_fill_1 FILLER_27_2550 ();
 sg13g2_fill_2 FILLER_27_2556 ();
 sg13g2_decap_4 FILLER_27_2588 ();
 sg13g2_fill_1 FILLER_27_2592 ();
 sg13g2_decap_8 FILLER_27_2597 ();
 sg13g2_decap_8 FILLER_27_2604 ();
 sg13g2_decap_8 FILLER_27_2618 ();
 sg13g2_fill_2 FILLER_27_2625 ();
 sg13g2_decap_4 FILLER_27_2665 ();
 sg13g2_fill_1 FILLER_27_2669 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_32 ();
 sg13g2_fill_2 FILLER_28_73 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_fill_1 FILLER_28_186 ();
 sg13g2_fill_2 FILLER_28_235 ();
 sg13g2_fill_1 FILLER_28_237 ();
 sg13g2_fill_2 FILLER_28_264 ();
 sg13g2_fill_1 FILLER_28_266 ();
 sg13g2_fill_1 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_411 ();
 sg13g2_decap_4 FILLER_28_418 ();
 sg13g2_fill_2 FILLER_28_453 ();
 sg13g2_fill_2 FILLER_28_472 ();
 sg13g2_fill_1 FILLER_28_521 ();
 sg13g2_fill_2 FILLER_28_543 ();
 sg13g2_fill_1 FILLER_28_545 ();
 sg13g2_fill_2 FILLER_28_615 ();
 sg13g2_fill_1 FILLER_28_640 ();
 sg13g2_fill_2 FILLER_28_675 ();
 sg13g2_decap_4 FILLER_28_686 ();
 sg13g2_fill_2 FILLER_28_690 ();
 sg13g2_fill_1 FILLER_28_701 ();
 sg13g2_fill_2 FILLER_28_775 ();
 sg13g2_fill_1 FILLER_28_777 ();
 sg13g2_fill_1 FILLER_28_804 ();
 sg13g2_fill_1 FILLER_28_872 ();
 sg13g2_fill_2 FILLER_28_953 ();
 sg13g2_fill_1 FILLER_28_959 ();
 sg13g2_fill_1 FILLER_28_991 ();
 sg13g2_fill_2 FILLER_28_1017 ();
 sg13g2_fill_2 FILLER_28_1037 ();
 sg13g2_fill_1 FILLER_28_1039 ();
 sg13g2_fill_1 FILLER_28_1054 ();
 sg13g2_fill_2 FILLER_28_1071 ();
 sg13g2_fill_1 FILLER_28_1073 ();
 sg13g2_decap_8 FILLER_28_1105 ();
 sg13g2_fill_1 FILLER_28_1112 ();
 sg13g2_decap_8 FILLER_28_1117 ();
 sg13g2_fill_1 FILLER_28_1145 ();
 sg13g2_fill_1 FILLER_28_1149 ();
 sg13g2_fill_1 FILLER_28_1183 ();
 sg13g2_fill_2 FILLER_28_1221 ();
 sg13g2_fill_1 FILLER_28_1265 ();
 sg13g2_fill_2 FILLER_28_1269 ();
 sg13g2_fill_1 FILLER_28_1312 ();
 sg13g2_fill_1 FILLER_28_1342 ();
 sg13g2_fill_1 FILLER_28_1352 ();
 sg13g2_fill_2 FILLER_28_1363 ();
 sg13g2_decap_8 FILLER_28_1369 ();
 sg13g2_decap_8 FILLER_28_1376 ();
 sg13g2_decap_8 FILLER_28_1383 ();
 sg13g2_fill_2 FILLER_28_1390 ();
 sg13g2_decap_4 FILLER_28_1439 ();
 sg13g2_fill_1 FILLER_28_1443 ();
 sg13g2_fill_2 FILLER_28_1452 ();
 sg13g2_decap_8 FILLER_28_1525 ();
 sg13g2_decap_4 FILLER_28_1532 ();
 sg13g2_fill_2 FILLER_28_1592 ();
 sg13g2_fill_2 FILLER_28_1601 ();
 sg13g2_fill_2 FILLER_28_1631 ();
 sg13g2_fill_1 FILLER_28_1666 ();
 sg13g2_fill_2 FILLER_28_1698 ();
 sg13g2_fill_1 FILLER_28_1700 ();
 sg13g2_decap_8 FILLER_28_1736 ();
 sg13g2_fill_2 FILLER_28_1781 ();
 sg13g2_fill_1 FILLER_28_1783 ();
 sg13g2_fill_1 FILLER_28_1814 ();
 sg13g2_fill_2 FILLER_28_1839 ();
 sg13g2_fill_1 FILLER_28_1853 ();
 sg13g2_fill_1 FILLER_28_1893 ();
 sg13g2_fill_1 FILLER_28_1960 ();
 sg13g2_decap_8 FILLER_28_1969 ();
 sg13g2_decap_4 FILLER_28_1976 ();
 sg13g2_fill_2 FILLER_28_1999 ();
 sg13g2_fill_2 FILLER_28_2030 ();
 sg13g2_fill_2 FILLER_28_2037 ();
 sg13g2_fill_1 FILLER_28_2039 ();
 sg13g2_fill_2 FILLER_28_2049 ();
 sg13g2_fill_1 FILLER_28_2051 ();
 sg13g2_fill_1 FILLER_28_2086 ();
 sg13g2_fill_2 FILLER_28_2096 ();
 sg13g2_fill_2 FILLER_28_2102 ();
 sg13g2_fill_2 FILLER_28_2108 ();
 sg13g2_fill_1 FILLER_28_2110 ();
 sg13g2_fill_2 FILLER_28_2119 ();
 sg13g2_decap_8 FILLER_28_2155 ();
 sg13g2_decap_8 FILLER_28_2162 ();
 sg13g2_fill_1 FILLER_28_2209 ();
 sg13g2_fill_2 FILLER_28_2216 ();
 sg13g2_fill_1 FILLER_28_2234 ();
 sg13g2_decap_8 FILLER_28_2240 ();
 sg13g2_decap_4 FILLER_28_2247 ();
 sg13g2_fill_2 FILLER_28_2251 ();
 sg13g2_fill_2 FILLER_28_2258 ();
 sg13g2_fill_1 FILLER_28_2260 ();
 sg13g2_decap_8 FILLER_28_2327 ();
 sg13g2_fill_1 FILLER_28_2349 ();
 sg13g2_fill_2 FILLER_28_2363 ();
 sg13g2_decap_4 FILLER_28_2393 ();
 sg13g2_fill_1 FILLER_28_2402 ();
 sg13g2_fill_1 FILLER_28_2408 ();
 sg13g2_decap_4 FILLER_28_2417 ();
 sg13g2_decap_8 FILLER_28_2434 ();
 sg13g2_decap_8 FILLER_28_2445 ();
 sg13g2_decap_4 FILLER_28_2457 ();
 sg13g2_fill_1 FILLER_28_2461 ();
 sg13g2_decap_8 FILLER_28_2474 ();
 sg13g2_decap_8 FILLER_28_2481 ();
 sg13g2_decap_4 FILLER_28_2488 ();
 sg13g2_fill_1 FILLER_28_2492 ();
 sg13g2_decap_4 FILLER_28_2498 ();
 sg13g2_decap_4 FILLER_28_2516 ();
 sg13g2_fill_2 FILLER_28_2520 ();
 sg13g2_fill_1 FILLER_28_2534 ();
 sg13g2_decap_4 FILLER_28_2544 ();
 sg13g2_fill_1 FILLER_28_2548 ();
 sg13g2_fill_2 FILLER_28_2565 ();
 sg13g2_decap_4 FILLER_28_2585 ();
 sg13g2_fill_2 FILLER_28_2610 ();
 sg13g2_fill_1 FILLER_28_2612 ();
 sg13g2_decap_4 FILLER_28_2634 ();
 sg13g2_decap_8 FILLER_28_2659 ();
 sg13g2_decap_4 FILLER_28_2666 ();
 sg13g2_fill_2 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_62 ();
 sg13g2_fill_1 FILLER_29_64 ();
 sg13g2_fill_1 FILLER_29_79 ();
 sg13g2_decap_4 FILLER_29_127 ();
 sg13g2_decap_4 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_334 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_decap_4 FILLER_29_355 ();
 sg13g2_fill_1 FILLER_29_364 ();
 sg13g2_fill_1 FILLER_29_369 ();
 sg13g2_fill_2 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_402 ();
 sg13g2_decap_4 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_29_459 ();
 sg13g2_decap_8 FILLER_29_466 ();
 sg13g2_decap_8 FILLER_29_473 ();
 sg13g2_fill_2 FILLER_29_480 ();
 sg13g2_fill_1 FILLER_29_485 ();
 sg13g2_fill_1 FILLER_29_552 ();
 sg13g2_fill_1 FILLER_29_601 ();
 sg13g2_decap_4 FILLER_29_606 ();
 sg13g2_fill_2 FILLER_29_610 ();
 sg13g2_fill_2 FILLER_29_616 ();
 sg13g2_fill_1 FILLER_29_618 ();
 sg13g2_fill_2 FILLER_29_623 ();
 sg13g2_decap_4 FILLER_29_642 ();
 sg13g2_fill_1 FILLER_29_646 ();
 sg13g2_fill_2 FILLER_29_655 ();
 sg13g2_fill_2 FILLER_29_661 ();
 sg13g2_fill_1 FILLER_29_667 ();
 sg13g2_fill_2 FILLER_29_742 ();
 sg13g2_fill_2 FILLER_29_832 ();
 sg13g2_fill_2 FILLER_29_884 ();
 sg13g2_fill_1 FILLER_29_890 ();
 sg13g2_fill_2 FILLER_29_899 ();
 sg13g2_fill_1 FILLER_29_901 ();
 sg13g2_fill_1 FILLER_29_907 ();
 sg13g2_fill_2 FILLER_29_912 ();
 sg13g2_fill_2 FILLER_29_918 ();
 sg13g2_fill_1 FILLER_29_920 ();
 sg13g2_fill_2 FILLER_29_926 ();
 sg13g2_fill_2 FILLER_29_949 ();
 sg13g2_fill_1 FILLER_29_951 ();
 sg13g2_fill_2 FILLER_29_957 ();
 sg13g2_fill_1 FILLER_29_959 ();
 sg13g2_fill_2 FILLER_29_964 ();
 sg13g2_fill_1 FILLER_29_971 ();
 sg13g2_fill_2 FILLER_29_1002 ();
 sg13g2_fill_1 FILLER_29_1030 ();
 sg13g2_fill_2 FILLER_29_1052 ();
 sg13g2_fill_1 FILLER_29_1054 ();
 sg13g2_fill_2 FILLER_29_1071 ();
 sg13g2_fill_1 FILLER_29_1073 ();
 sg13g2_decap_8 FILLER_29_1112 ();
 sg13g2_decap_4 FILLER_29_1119 ();
 sg13g2_fill_1 FILLER_29_1123 ();
 sg13g2_fill_2 FILLER_29_1218 ();
 sg13g2_fill_2 FILLER_29_1226 ();
 sg13g2_fill_2 FILLER_29_1312 ();
 sg13g2_fill_2 FILLER_29_1344 ();
 sg13g2_decap_8 FILLER_29_1367 ();
 sg13g2_decap_8 FILLER_29_1374 ();
 sg13g2_decap_8 FILLER_29_1381 ();
 sg13g2_decap_4 FILLER_29_1388 ();
 sg13g2_fill_2 FILLER_29_1392 ();
 sg13g2_decap_4 FILLER_29_1398 ();
 sg13g2_fill_2 FILLER_29_1427 ();
 sg13g2_fill_1 FILLER_29_1429 ();
 sg13g2_decap_8 FILLER_29_1434 ();
 sg13g2_fill_2 FILLER_29_1451 ();
 sg13g2_fill_1 FILLER_29_1489 ();
 sg13g2_fill_2 FILLER_29_1547 ();
 sg13g2_fill_1 FILLER_29_1566 ();
 sg13g2_fill_1 FILLER_29_1598 ();
 sg13g2_fill_2 FILLER_29_1612 ();
 sg13g2_fill_1 FILLER_29_1642 ();
 sg13g2_fill_2 FILLER_29_1699 ();
 sg13g2_fill_2 FILLER_29_1739 ();
 sg13g2_fill_1 FILLER_29_1741 ();
 sg13g2_fill_2 FILLER_29_1746 ();
 sg13g2_fill_2 FILLER_29_1753 ();
 sg13g2_fill_1 FILLER_29_1755 ();
 sg13g2_fill_1 FILLER_29_1760 ();
 sg13g2_fill_1 FILLER_29_1766 ();
 sg13g2_fill_2 FILLER_29_1806 ();
 sg13g2_fill_2 FILLER_29_1830 ();
 sg13g2_fill_1 FILLER_29_1849 ();
 sg13g2_fill_1 FILLER_29_1875 ();
 sg13g2_fill_1 FILLER_29_1918 ();
 sg13g2_fill_2 FILLER_29_1931 ();
 sg13g2_fill_2 FILLER_29_1950 ();
 sg13g2_decap_8 FILLER_29_1956 ();
 sg13g2_fill_2 FILLER_29_1963 ();
 sg13g2_fill_2 FILLER_29_1978 ();
 sg13g2_fill_1 FILLER_29_2001 ();
 sg13g2_decap_8 FILLER_29_2009 ();
 sg13g2_decap_4 FILLER_29_2016 ();
 sg13g2_fill_2 FILLER_29_2020 ();
 sg13g2_decap_4 FILLER_29_2026 ();
 sg13g2_decap_8 FILLER_29_2034 ();
 sg13g2_fill_1 FILLER_29_2045 ();
 sg13g2_decap_8 FILLER_29_2076 ();
 sg13g2_decap_8 FILLER_29_2083 ();
 sg13g2_fill_2 FILLER_29_2090 ();
 sg13g2_fill_1 FILLER_29_2092 ();
 sg13g2_decap_8 FILLER_29_2097 ();
 sg13g2_fill_2 FILLER_29_2104 ();
 sg13g2_decap_8 FILLER_29_2158 ();
 sg13g2_decap_8 FILLER_29_2165 ();
 sg13g2_decap_4 FILLER_29_2172 ();
 sg13g2_fill_2 FILLER_29_2197 ();
 sg13g2_fill_1 FILLER_29_2199 ();
 sg13g2_fill_2 FILLER_29_2239 ();
 sg13g2_fill_1 FILLER_29_2241 ();
 sg13g2_decap_8 FILLER_29_2251 ();
 sg13g2_fill_1 FILLER_29_2283 ();
 sg13g2_fill_2 FILLER_29_2332 ();
 sg13g2_fill_1 FILLER_29_2334 ();
 sg13g2_fill_1 FILLER_29_2361 ();
 sg13g2_decap_4 FILLER_29_2383 ();
 sg13g2_fill_1 FILLER_29_2387 ();
 sg13g2_fill_1 FILLER_29_2393 ();
 sg13g2_fill_1 FILLER_29_2399 ();
 sg13g2_fill_1 FILLER_29_2405 ();
 sg13g2_decap_4 FILLER_29_2411 ();
 sg13g2_fill_2 FILLER_29_2427 ();
 sg13g2_fill_1 FILLER_29_2429 ();
 sg13g2_fill_2 FILLER_29_2435 ();
 sg13g2_fill_1 FILLER_29_2441 ();
 sg13g2_fill_2 FILLER_29_2461 ();
 sg13g2_decap_8 FILLER_29_2476 ();
 sg13g2_fill_1 FILLER_29_2483 ();
 sg13g2_decap_4 FILLER_29_2489 ();
 sg13g2_fill_2 FILLER_29_2497 ();
 sg13g2_fill_1 FILLER_29_2508 ();
 sg13g2_fill_1 FILLER_29_2521 ();
 sg13g2_fill_1 FILLER_29_2531 ();
 sg13g2_decap_8 FILLER_29_2538 ();
 sg13g2_fill_1 FILLER_29_2545 ();
 sg13g2_decap_4 FILLER_29_2573 ();
 sg13g2_fill_1 FILLER_29_2577 ();
 sg13g2_fill_1 FILLER_29_2583 ();
 sg13g2_fill_1 FILLER_29_2589 ();
 sg13g2_decap_8 FILLER_29_2621 ();
 sg13g2_decap_8 FILLER_29_2628 ();
 sg13g2_decap_8 FILLER_29_2635 ();
 sg13g2_decap_8 FILLER_29_2642 ();
 sg13g2_decap_8 FILLER_29_2649 ();
 sg13g2_decap_8 FILLER_29_2656 ();
 sg13g2_decap_8 FILLER_29_2663 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_decap_4 FILLER_30_92 ();
 sg13g2_fill_1 FILLER_30_96 ();
 sg13g2_decap_8 FILLER_30_135 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_decap_4 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_185 ();
 sg13g2_decap_4 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_fill_2 FILLER_30_232 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_decap_8 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_4 FILLER_30_381 ();
 sg13g2_fill_2 FILLER_30_425 ();
 sg13g2_decap_8 FILLER_30_431 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_fill_1 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_561 ();
 sg13g2_decap_8 FILLER_30_568 ();
 sg13g2_decap_8 FILLER_30_579 ();
 sg13g2_fill_1 FILLER_30_595 ();
 sg13g2_fill_1 FILLER_30_665 ();
 sg13g2_fill_2 FILLER_30_711 ();
 sg13g2_fill_1 FILLER_30_713 ();
 sg13g2_fill_1 FILLER_30_755 ();
 sg13g2_decap_8 FILLER_30_781 ();
 sg13g2_decap_4 FILLER_30_788 ();
 sg13g2_fill_1 FILLER_30_804 ();
 sg13g2_fill_2 FILLER_30_814 ();
 sg13g2_fill_1 FILLER_30_842 ();
 sg13g2_fill_2 FILLER_30_851 ();
 sg13g2_fill_1 FILLER_30_884 ();
 sg13g2_decap_4 FILLER_30_906 ();
 sg13g2_fill_1 FILLER_30_910 ();
 sg13g2_fill_1 FILLER_30_916 ();
 sg13g2_decap_4 FILLER_30_922 ();
 sg13g2_fill_1 FILLER_30_926 ();
 sg13g2_decap_4 FILLER_30_1008 ();
 sg13g2_fill_1 FILLER_30_1012 ();
 sg13g2_decap_8 FILLER_30_1017 ();
 sg13g2_fill_2 FILLER_30_1033 ();
 sg13g2_fill_1 FILLER_30_1035 ();
 sg13g2_fill_1 FILLER_30_1057 ();
 sg13g2_fill_2 FILLER_30_1067 ();
 sg13g2_fill_1 FILLER_30_1069 ();
 sg13g2_fill_2 FILLER_30_1089 ();
 sg13g2_fill_2 FILLER_30_1121 ();
 sg13g2_fill_2 FILLER_30_1165 ();
 sg13g2_fill_2 FILLER_30_1170 ();
 sg13g2_fill_1 FILLER_30_1282 ();
 sg13g2_fill_2 FILLER_30_1305 ();
 sg13g2_fill_2 FILLER_30_1315 ();
 sg13g2_fill_1 FILLER_30_1326 ();
 sg13g2_fill_1 FILLER_30_1331 ();
 sg13g2_fill_2 FILLER_30_1336 ();
 sg13g2_fill_2 FILLER_30_1347 ();
 sg13g2_decap_4 FILLER_30_1379 ();
 sg13g2_fill_2 FILLER_30_1421 ();
 sg13g2_fill_1 FILLER_30_1432 ();
 sg13g2_fill_1 FILLER_30_1496 ();
 sg13g2_fill_2 FILLER_30_1510 ();
 sg13g2_fill_2 FILLER_30_1522 ();
 sg13g2_fill_1 FILLER_30_1524 ();
 sg13g2_fill_2 FILLER_30_1580 ();
 sg13g2_fill_2 FILLER_30_1605 ();
 sg13g2_fill_1 FILLER_30_1657 ();
 sg13g2_fill_1 FILLER_30_1694 ();
 sg13g2_fill_1 FILLER_30_1730 ();
 sg13g2_fill_1 FILLER_30_1735 ();
 sg13g2_fill_2 FILLER_30_1783 ();
 sg13g2_fill_2 FILLER_30_1822 ();
 sg13g2_fill_2 FILLER_30_1849 ();
 sg13g2_fill_2 FILLER_30_1867 ();
 sg13g2_fill_1 FILLER_30_1936 ();
 sg13g2_decap_4 FILLER_30_1945 ();
 sg13g2_fill_2 FILLER_30_1949 ();
 sg13g2_decap_4 FILLER_30_2013 ();
 sg13g2_fill_1 FILLER_30_2017 ();
 sg13g2_fill_2 FILLER_30_2022 ();
 sg13g2_fill_1 FILLER_30_2033 ();
 sg13g2_decap_4 FILLER_30_2064 ();
 sg13g2_fill_1 FILLER_30_2132 ();
 sg13g2_decap_4 FILLER_30_2137 ();
 sg13g2_decap_8 FILLER_30_2145 ();
 sg13g2_decap_8 FILLER_30_2152 ();
 sg13g2_decap_8 FILLER_30_2159 ();
 sg13g2_decap_4 FILLER_30_2166 ();
 sg13g2_fill_2 FILLER_30_2170 ();
 sg13g2_fill_2 FILLER_30_2189 ();
 sg13g2_fill_1 FILLER_30_2244 ();
 sg13g2_decap_4 FILLER_30_2293 ();
 sg13g2_fill_2 FILLER_30_2297 ();
 sg13g2_fill_1 FILLER_30_2304 ();
 sg13g2_decap_4 FILLER_30_2310 ();
 sg13g2_fill_2 FILLER_30_2318 ();
 sg13g2_fill_1 FILLER_30_2343 ();
 sg13g2_decap_8 FILLER_30_2353 ();
 sg13g2_fill_2 FILLER_30_2360 ();
 sg13g2_fill_2 FILLER_30_2378 ();
 sg13g2_fill_1 FILLER_30_2397 ();
 sg13g2_fill_1 FILLER_30_2406 ();
 sg13g2_fill_1 FILLER_30_2415 ();
 sg13g2_decap_4 FILLER_30_2424 ();
 sg13g2_decap_8 FILLER_30_2433 ();
 sg13g2_decap_4 FILLER_30_2440 ();
 sg13g2_fill_2 FILLER_30_2444 ();
 sg13g2_decap_8 FILLER_30_2488 ();
 sg13g2_decap_4 FILLER_30_2495 ();
 sg13g2_fill_2 FILLER_30_2522 ();
 sg13g2_decap_4 FILLER_30_2531 ();
 sg13g2_decap_4 FILLER_30_2559 ();
 sg13g2_decap_4 FILLER_30_2572 ();
 sg13g2_fill_1 FILLER_30_2576 ();
 sg13g2_fill_1 FILLER_30_2580 ();
 sg13g2_decap_8 FILLER_30_2584 ();
 sg13g2_fill_1 FILLER_30_2604 ();
 sg13g2_fill_2 FILLER_30_2647 ();
 sg13g2_fill_1 FILLER_30_2649 ();
 sg13g2_decap_8 FILLER_30_2655 ();
 sg13g2_decap_8 FILLER_30_2662 ();
 sg13g2_fill_1 FILLER_30_2669 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_27 ();
 sg13g2_fill_1 FILLER_31_29 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_93 ();
 sg13g2_decap_8 FILLER_31_115 ();
 sg13g2_decap_8 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_129 ();
 sg13g2_decap_8 FILLER_31_136 ();
 sg13g2_decap_8 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_173 ();
 sg13g2_decap_4 FILLER_31_182 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_fill_2 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_fill_1 FILLER_31_265 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_decap_4 FILLER_31_310 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_decap_4 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_fill_2 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_31_409 ();
 sg13g2_decap_4 FILLER_31_416 ();
 sg13g2_fill_1 FILLER_31_420 ();
 sg13g2_fill_1 FILLER_31_477 ();
 sg13g2_decap_8 FILLER_31_482 ();
 sg13g2_decap_8 FILLER_31_489 ();
 sg13g2_decap_4 FILLER_31_496 ();
 sg13g2_fill_1 FILLER_31_500 ();
 sg13g2_decap_8 FILLER_31_509 ();
 sg13g2_decap_8 FILLER_31_516 ();
 sg13g2_fill_2 FILLER_31_523 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_fill_1 FILLER_31_553 ();
 sg13g2_fill_1 FILLER_31_593 ();
 sg13g2_fill_1 FILLER_31_603 ();
 sg13g2_decap_4 FILLER_31_609 ();
 sg13g2_fill_2 FILLER_31_650 ();
 sg13g2_fill_1 FILLER_31_678 ();
 sg13g2_fill_1 FILLER_31_686 ();
 sg13g2_fill_1 FILLER_31_695 ();
 sg13g2_fill_1 FILLER_31_715 ();
 sg13g2_fill_2 FILLER_31_733 ();
 sg13g2_fill_1 FILLER_31_751 ();
 sg13g2_fill_2 FILLER_31_760 ();
 sg13g2_fill_1 FILLER_31_766 ();
 sg13g2_fill_1 FILLER_31_783 ();
 sg13g2_fill_1 FILLER_31_823 ();
 sg13g2_decap_8 FILLER_31_912 ();
 sg13g2_decap_4 FILLER_31_919 ();
 sg13g2_fill_1 FILLER_31_923 ();
 sg13g2_fill_2 FILLER_31_933 ();
 sg13g2_fill_2 FILLER_31_942 ();
 sg13g2_fill_1 FILLER_31_944 ();
 sg13g2_decap_4 FILLER_31_954 ();
 sg13g2_fill_2 FILLER_31_970 ();
 sg13g2_fill_2 FILLER_31_976 ();
 sg13g2_fill_1 FILLER_31_978 ();
 sg13g2_fill_1 FILLER_31_984 ();
 sg13g2_decap_4 FILLER_31_989 ();
 sg13g2_fill_2 FILLER_31_993 ();
 sg13g2_decap_8 FILLER_31_999 ();
 sg13g2_decap_8 FILLER_31_1006 ();
 sg13g2_decap_4 FILLER_31_1013 ();
 sg13g2_fill_2 FILLER_31_1017 ();
 sg13g2_fill_1 FILLER_31_1045 ();
 sg13g2_fill_2 FILLER_31_1111 ();
 sg13g2_fill_2 FILLER_31_1194 ();
 sg13g2_fill_1 FILLER_31_1342 ();
 sg13g2_decap_4 FILLER_31_1352 ();
 sg13g2_fill_1 FILLER_31_1356 ();
 sg13g2_decap_8 FILLER_31_1361 ();
 sg13g2_decap_4 FILLER_31_1394 ();
 sg13g2_fill_1 FILLER_31_1403 ();
 sg13g2_fill_2 FILLER_31_1408 ();
 sg13g2_fill_1 FILLER_31_1410 ();
 sg13g2_fill_1 FILLER_31_1456 ();
 sg13g2_fill_2 FILLER_31_1526 ();
 sg13g2_fill_1 FILLER_31_1528 ();
 sg13g2_decap_4 FILLER_31_1571 ();
 sg13g2_fill_1 FILLER_31_1579 ();
 sg13g2_fill_1 FILLER_31_1631 ();
 sg13g2_fill_2 FILLER_31_1637 ();
 sg13g2_fill_2 FILLER_31_1643 ();
 sg13g2_fill_1 FILLER_31_1675 ();
 sg13g2_fill_1 FILLER_31_1733 ();
 sg13g2_fill_1 FILLER_31_1790 ();
 sg13g2_fill_2 FILLER_31_1817 ();
 sg13g2_fill_1 FILLER_31_1850 ();
 sg13g2_fill_2 FILLER_31_1881 ();
 sg13g2_fill_2 FILLER_31_1990 ();
 sg13g2_fill_2 FILLER_31_2031 ();
 sg13g2_decap_8 FILLER_31_2059 ();
 sg13g2_fill_2 FILLER_31_2087 ();
 sg13g2_decap_8 FILLER_31_2093 ();
 sg13g2_decap_8 FILLER_31_2100 ();
 sg13g2_fill_2 FILLER_31_2107 ();
 sg13g2_fill_1 FILLER_31_2109 ();
 sg13g2_fill_1 FILLER_31_2131 ();
 sg13g2_decap_4 FILLER_31_2162 ();
 sg13g2_fill_1 FILLER_31_2175 ();
 sg13g2_fill_2 FILLER_31_2180 ();
 sg13g2_fill_2 FILLER_31_2187 ();
 sg13g2_fill_2 FILLER_31_2193 ();
 sg13g2_fill_2 FILLER_31_2200 ();
 sg13g2_fill_1 FILLER_31_2217 ();
 sg13g2_decap_8 FILLER_31_2222 ();
 sg13g2_fill_2 FILLER_31_2229 ();
 sg13g2_fill_1 FILLER_31_2231 ();
 sg13g2_fill_1 FILLER_31_2237 ();
 sg13g2_decap_8 FILLER_31_2242 ();
 sg13g2_fill_1 FILLER_31_2249 ();
 sg13g2_fill_2 FILLER_31_2256 ();
 sg13g2_decap_8 FILLER_31_2268 ();
 sg13g2_fill_1 FILLER_31_2275 ();
 sg13g2_decap_4 FILLER_31_2305 ();
 sg13g2_decap_8 FILLER_31_2317 ();
 sg13g2_fill_2 FILLER_31_2338 ();
 sg13g2_fill_1 FILLER_31_2340 ();
 sg13g2_decap_8 FILLER_31_2353 ();
 sg13g2_fill_1 FILLER_31_2360 ();
 sg13g2_decap_4 FILLER_31_2423 ();
 sg13g2_fill_2 FILLER_31_2427 ();
 sg13g2_decap_4 FILLER_31_2437 ();
 sg13g2_fill_2 FILLER_31_2441 ();
 sg13g2_decap_4 FILLER_31_2488 ();
 sg13g2_fill_1 FILLER_31_2492 ();
 sg13g2_decap_4 FILLER_31_2527 ();
 sg13g2_fill_1 FILLER_31_2539 ();
 sg13g2_fill_1 FILLER_31_2573 ();
 sg13g2_fill_2 FILLER_31_2605 ();
 sg13g2_decap_8 FILLER_31_2620 ();
 sg13g2_fill_1 FILLER_31_2627 ();
 sg13g2_decap_8 FILLER_31_2649 ();
 sg13g2_decap_8 FILLER_31_2656 ();
 sg13g2_decap_8 FILLER_31_2663 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_32 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_fill_2 FILLER_32_44 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_fill_2 FILLER_32_52 ();
 sg13g2_decap_4 FILLER_32_58 ();
 sg13g2_decap_8 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_92 ();
 sg13g2_fill_2 FILLER_32_135 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_290 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_321 ();
 sg13g2_decap_4 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_4 FILLER_32_434 ();
 sg13g2_fill_1 FILLER_32_438 ();
 sg13g2_decap_8 FILLER_32_443 ();
 sg13g2_fill_2 FILLER_32_450 ();
 sg13g2_fill_1 FILLER_32_452 ();
 sg13g2_decap_8 FILLER_32_470 ();
 sg13g2_decap_8 FILLER_32_477 ();
 sg13g2_decap_4 FILLER_32_484 ();
 sg13g2_decap_8 FILLER_32_518 ();
 sg13g2_decap_8 FILLER_32_525 ();
 sg13g2_decap_8 FILLER_32_532 ();
 sg13g2_fill_1 FILLER_32_539 ();
 sg13g2_decap_8 FILLER_32_582 ();
 sg13g2_fill_1 FILLER_32_619 ();
 sg13g2_fill_2 FILLER_32_648 ();
 sg13g2_fill_2 FILLER_32_660 ();
 sg13g2_fill_2 FILLER_32_678 ();
 sg13g2_fill_1 FILLER_32_680 ();
 sg13g2_fill_2 FILLER_32_686 ();
 sg13g2_fill_2 FILLER_32_709 ();
 sg13g2_fill_2 FILLER_32_715 ();
 sg13g2_fill_1 FILLER_32_717 ();
 sg13g2_fill_2 FILLER_32_723 ();
 sg13g2_fill_2 FILLER_32_729 ();
 sg13g2_fill_1 FILLER_32_735 ();
 sg13g2_fill_2 FILLER_32_745 ();
 sg13g2_fill_1 FILLER_32_819 ();
 sg13g2_fill_2 FILLER_32_851 ();
 sg13g2_fill_1 FILLER_32_857 ();
 sg13g2_fill_1 FILLER_32_862 ();
 sg13g2_fill_2 FILLER_32_876 ();
 sg13g2_fill_1 FILLER_32_878 ();
 sg13g2_fill_1 FILLER_32_905 ();
 sg13g2_fill_2 FILLER_32_915 ();
 sg13g2_fill_1 FILLER_32_917 ();
 sg13g2_fill_1 FILLER_32_962 ();
 sg13g2_fill_2 FILLER_32_971 ();
 sg13g2_fill_1 FILLER_32_992 ();
 sg13g2_fill_1 FILLER_32_1065 ();
 sg13g2_decap_4 FILLER_32_1104 ();
 sg13g2_fill_1 FILLER_32_1108 ();
 sg13g2_fill_2 FILLER_32_1141 ();
 sg13g2_fill_2 FILLER_32_1200 ();
 sg13g2_fill_2 FILLER_32_1226 ();
 sg13g2_fill_2 FILLER_32_1275 ();
 sg13g2_fill_2 FILLER_32_1307 ();
 sg13g2_fill_2 FILLER_32_1314 ();
 sg13g2_fill_2 FILLER_32_1337 ();
 sg13g2_decap_8 FILLER_32_1364 ();
 sg13g2_decap_4 FILLER_32_1371 ();
 sg13g2_fill_1 FILLER_32_1396 ();
 sg13g2_fill_1 FILLER_32_1423 ();
 sg13g2_fill_1 FILLER_32_1442 ();
 sg13g2_fill_2 FILLER_32_1448 ();
 sg13g2_fill_1 FILLER_32_1506 ();
 sg13g2_fill_1 FILLER_32_1533 ();
 sg13g2_fill_1 FILLER_32_1560 ();
 sg13g2_fill_1 FILLER_32_1612 ();
 sg13g2_fill_1 FILLER_32_1641 ();
 sg13g2_decap_8 FILLER_32_1663 ();
 sg13g2_decap_8 FILLER_32_1670 ();
 sg13g2_fill_2 FILLER_32_1677 ();
 sg13g2_decap_8 FILLER_32_1691 ();
 sg13g2_fill_2 FILLER_32_1698 ();
 sg13g2_decap_8 FILLER_32_1721 ();
 sg13g2_fill_1 FILLER_32_1741 ();
 sg13g2_fill_1 FILLER_32_1750 ();
 sg13g2_fill_2 FILLER_32_1763 ();
 sg13g2_fill_1 FILLER_32_1794 ();
 sg13g2_fill_1 FILLER_32_1799 ();
 sg13g2_fill_2 FILLER_32_1837 ();
 sg13g2_fill_1 FILLER_32_1919 ();
 sg13g2_fill_2 FILLER_32_2010 ();
 sg13g2_fill_2 FILLER_32_2046 ();
 sg13g2_fill_1 FILLER_32_2048 ();
 sg13g2_decap_8 FILLER_32_2153 ();
 sg13g2_fill_2 FILLER_32_2160 ();
 sg13g2_fill_1 FILLER_32_2162 ();
 sg13g2_fill_2 FILLER_32_2182 ();
 sg13g2_fill_1 FILLER_32_2221 ();
 sg13g2_fill_2 FILLER_32_2227 ();
 sg13g2_fill_1 FILLER_32_2229 ();
 sg13g2_fill_1 FILLER_32_2233 ();
 sg13g2_fill_2 FILLER_32_2239 ();
 sg13g2_decap_4 FILLER_32_2252 ();
 sg13g2_decap_8 FILLER_32_2306 ();
 sg13g2_decap_8 FILLER_32_2313 ();
 sg13g2_decap_4 FILLER_32_2320 ();
 sg13g2_decap_4 FILLER_32_2328 ();
 sg13g2_fill_1 FILLER_32_2332 ();
 sg13g2_fill_2 FILLER_32_2338 ();
 sg13g2_fill_1 FILLER_32_2340 ();
 sg13g2_decap_8 FILLER_32_2348 ();
 sg13g2_decap_8 FILLER_32_2355 ();
 sg13g2_decap_8 FILLER_32_2362 ();
 sg13g2_decap_4 FILLER_32_2369 ();
 sg13g2_fill_2 FILLER_32_2373 ();
 sg13g2_fill_2 FILLER_32_2434 ();
 sg13g2_decap_8 FILLER_32_2448 ();
 sg13g2_decap_4 FILLER_32_2455 ();
 sg13g2_fill_1 FILLER_32_2459 ();
 sg13g2_fill_2 FILLER_32_2479 ();
 sg13g2_fill_1 FILLER_32_2485 ();
 sg13g2_fill_2 FILLER_32_2501 ();
 sg13g2_fill_2 FILLER_32_2535 ();
 sg13g2_fill_1 FILLER_32_2537 ();
 sg13g2_fill_1 FILLER_32_2545 ();
 sg13g2_fill_2 FILLER_32_2554 ();
 sg13g2_fill_1 FILLER_32_2607 ();
 sg13g2_decap_8 FILLER_32_2658 ();
 sg13g2_decap_4 FILLER_32_2665 ();
 sg13g2_fill_1 FILLER_32_2669 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_32 ();
 sg13g2_decap_8 FILLER_33_58 ();
 sg13g2_fill_2 FILLER_33_65 ();
 sg13g2_fill_1 FILLER_33_67 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_142 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_4 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_fill_2 FILLER_33_321 ();
 sg13g2_fill_2 FILLER_33_362 ();
 sg13g2_fill_2 FILLER_33_390 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_fill_2 FILLER_33_419 ();
 sg13g2_fill_1 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_430 ();
 sg13g2_decap_8 FILLER_33_445 ();
 sg13g2_decap_4 FILLER_33_452 ();
 sg13g2_fill_1 FILLER_33_456 ();
 sg13g2_fill_2 FILLER_33_486 ();
 sg13g2_decap_8 FILLER_33_509 ();
 sg13g2_decap_4 FILLER_33_516 ();
 sg13g2_fill_2 FILLER_33_520 ();
 sg13g2_decap_4 FILLER_33_551 ();
 sg13g2_fill_1 FILLER_33_555 ();
 sg13g2_fill_1 FILLER_33_582 ();
 sg13g2_fill_2 FILLER_33_609 ();
 sg13g2_fill_1 FILLER_33_611 ();
 sg13g2_fill_1 FILLER_33_627 ();
 sg13g2_decap_8 FILLER_33_636 ();
 sg13g2_fill_1 FILLER_33_643 ();
 sg13g2_fill_2 FILLER_33_653 ();
 sg13g2_decap_4 FILLER_33_687 ();
 sg13g2_fill_2 FILLER_33_691 ();
 sg13g2_fill_2 FILLER_33_697 ();
 sg13g2_fill_1 FILLER_33_725 ();
 sg13g2_fill_1 FILLER_33_739 ();
 sg13g2_fill_1 FILLER_33_748 ();
 sg13g2_fill_1 FILLER_33_760 ();
 sg13g2_fill_1 FILLER_33_772 ();
 sg13g2_fill_1 FILLER_33_777 ();
 sg13g2_fill_1 FILLER_33_804 ();
 sg13g2_fill_2 FILLER_33_842 ();
 sg13g2_fill_1 FILLER_33_850 ();
 sg13g2_fill_1 FILLER_33_877 ();
 sg13g2_fill_1 FILLER_33_883 ();
 sg13g2_fill_1 FILLER_33_893 ();
 sg13g2_fill_2 FILLER_33_1038 ();
 sg13g2_fill_2 FILLER_33_1044 ();
 sg13g2_decap_8 FILLER_33_1072 ();
 sg13g2_fill_2 FILLER_33_1079 ();
 sg13g2_fill_1 FILLER_33_1081 ();
 sg13g2_decap_4 FILLER_33_1088 ();
 sg13g2_fill_2 FILLER_33_1092 ();
 sg13g2_decap_8 FILLER_33_1098 ();
 sg13g2_decap_8 FILLER_33_1105 ();
 sg13g2_decap_8 FILLER_33_1112 ();
 sg13g2_fill_2 FILLER_33_1119 ();
 sg13g2_fill_1 FILLER_33_1121 ();
 sg13g2_fill_1 FILLER_33_1149 ();
 sg13g2_fill_2 FILLER_33_1159 ();
 sg13g2_fill_2 FILLER_33_1194 ();
 sg13g2_fill_2 FILLER_33_1275 ();
 sg13g2_decap_8 FILLER_33_1350 ();
 sg13g2_decap_8 FILLER_33_1357 ();
 sg13g2_decap_8 FILLER_33_1364 ();
 sg13g2_decap_4 FILLER_33_1371 ();
 sg13g2_decap_8 FILLER_33_1396 ();
 sg13g2_decap_4 FILLER_33_1403 ();
 sg13g2_fill_2 FILLER_33_1424 ();
 sg13g2_fill_1 FILLER_33_1426 ();
 sg13g2_fill_2 FILLER_33_1459 ();
 sg13g2_fill_2 FILLER_33_1465 ();
 sg13g2_fill_2 FILLER_33_1472 ();
 sg13g2_fill_1 FILLER_33_1500 ();
 sg13g2_fill_1 FILLER_33_1514 ();
 sg13g2_fill_2 FILLER_33_1614 ();
 sg13g2_fill_1 FILLER_33_1640 ();
 sg13g2_fill_2 FILLER_33_1645 ();
 sg13g2_fill_2 FILLER_33_1660 ();
 sg13g2_decap_8 FILLER_33_1675 ();
 sg13g2_decap_8 FILLER_33_1682 ();
 sg13g2_decap_8 FILLER_33_1689 ();
 sg13g2_decap_8 FILLER_33_1696 ();
 sg13g2_decap_4 FILLER_33_1703 ();
 sg13g2_fill_2 FILLER_33_1740 ();
 sg13g2_fill_1 FILLER_33_1746 ();
 sg13g2_fill_1 FILLER_33_1755 ();
 sg13g2_fill_2 FILLER_33_1797 ();
 sg13g2_fill_1 FILLER_33_1861 ();
 sg13g2_fill_1 FILLER_33_1914 ();
 sg13g2_fill_1 FILLER_33_1966 ();
 sg13g2_fill_1 FILLER_33_2005 ();
 sg13g2_decap_8 FILLER_33_2055 ();
 sg13g2_fill_2 FILLER_33_2062 ();
 sg13g2_fill_1 FILLER_33_2064 ();
 sg13g2_fill_1 FILLER_33_2122 ();
 sg13g2_decap_8 FILLER_33_2149 ();
 sg13g2_decap_8 FILLER_33_2156 ();
 sg13g2_fill_2 FILLER_33_2163 ();
 sg13g2_fill_2 FILLER_33_2173 ();
 sg13g2_fill_2 FILLER_33_2192 ();
 sg13g2_fill_2 FILLER_33_2206 ();
 sg13g2_fill_1 FILLER_33_2212 ();
 sg13g2_decap_4 FILLER_33_2217 ();
 sg13g2_fill_2 FILLER_33_2221 ();
 sg13g2_fill_1 FILLER_33_2236 ();
 sg13g2_fill_2 FILLER_33_2247 ();
 sg13g2_decap_8 FILLER_33_2253 ();
 sg13g2_decap_8 FILLER_33_2260 ();
 sg13g2_fill_1 FILLER_33_2276 ();
 sg13g2_decap_4 FILLER_33_2303 ();
 sg13g2_fill_1 FILLER_33_2307 ();
 sg13g2_decap_4 FILLER_33_2318 ();
 sg13g2_decap_8 FILLER_33_2335 ();
 sg13g2_decap_8 FILLER_33_2347 ();
 sg13g2_fill_2 FILLER_33_2359 ();
 sg13g2_decap_8 FILLER_33_2366 ();
 sg13g2_fill_2 FILLER_33_2373 ();
 sg13g2_fill_1 FILLER_33_2375 ();
 sg13g2_decap_4 FILLER_33_2380 ();
 sg13g2_decap_8 FILLER_33_2394 ();
 sg13g2_fill_2 FILLER_33_2401 ();
 sg13g2_fill_1 FILLER_33_2428 ();
 sg13g2_fill_1 FILLER_33_2433 ();
 sg13g2_fill_1 FILLER_33_2438 ();
 sg13g2_decap_8 FILLER_33_2444 ();
 sg13g2_fill_1 FILLER_33_2451 ();
 sg13g2_fill_1 FILLER_33_2469 ();
 sg13g2_fill_1 FILLER_33_2489 ();
 sg13g2_fill_1 FILLER_33_2521 ();
 sg13g2_fill_2 FILLER_33_2548 ();
 sg13g2_decap_8 FILLER_33_2555 ();
 sg13g2_fill_2 FILLER_33_2562 ();
 sg13g2_fill_1 FILLER_33_2564 ();
 sg13g2_fill_1 FILLER_33_2569 ();
 sg13g2_fill_2 FILLER_33_2575 ();
 sg13g2_decap_4 FILLER_33_2589 ();
 sg13g2_decap_8 FILLER_33_2663 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_72 ();
 sg13g2_decap_8 FILLER_34_108 ();
 sg13g2_decap_8 FILLER_34_115 ();
 sg13g2_decap_8 FILLER_34_122 ();
 sg13g2_decap_8 FILLER_34_129 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_decap_4 FILLER_34_265 ();
 sg13g2_fill_2 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_fill_2 FILLER_34_387 ();
 sg13g2_fill_1 FILLER_34_389 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_fill_1 FILLER_34_416 ();
 sg13g2_fill_1 FILLER_34_447 ();
 sg13g2_fill_2 FILLER_34_503 ();
 sg13g2_fill_1 FILLER_34_505 ();
 sg13g2_decap_8 FILLER_34_540 ();
 sg13g2_fill_2 FILLER_34_547 ();
 sg13g2_fill_1 FILLER_34_549 ();
 sg13g2_decap_8 FILLER_34_571 ();
 sg13g2_fill_2 FILLER_34_578 ();
 sg13g2_fill_1 FILLER_34_580 ();
 sg13g2_fill_1 FILLER_34_591 ();
 sg13g2_fill_2 FILLER_34_601 ();
 sg13g2_fill_2 FILLER_34_620 ();
 sg13g2_fill_1 FILLER_34_622 ();
 sg13g2_decap_8 FILLER_34_629 ();
 sg13g2_decap_8 FILLER_34_636 ();
 sg13g2_fill_2 FILLER_34_643 ();
 sg13g2_fill_2 FILLER_34_660 ();
 sg13g2_fill_2 FILLER_34_692 ();
 sg13g2_fill_2 FILLER_34_702 ();
 sg13g2_fill_1 FILLER_34_704 ();
 sg13g2_fill_1 FILLER_34_718 ();
 sg13g2_fill_1 FILLER_34_724 ();
 sg13g2_fill_2 FILLER_34_730 ();
 sg13g2_fill_1 FILLER_34_732 ();
 sg13g2_fill_1 FILLER_34_771 ();
 sg13g2_fill_1 FILLER_34_788 ();
 sg13g2_fill_1 FILLER_34_838 ();
 sg13g2_fill_2 FILLER_34_850 ();
 sg13g2_fill_1 FILLER_34_878 ();
 sg13g2_fill_1 FILLER_34_884 ();
 sg13g2_fill_1 FILLER_34_919 ();
 sg13g2_fill_1 FILLER_34_1003 ();
 sg13g2_decap_8 FILLER_34_1030 ();
 sg13g2_fill_1 FILLER_34_1050 ();
 sg13g2_fill_2 FILLER_34_1068 ();
 sg13g2_fill_2 FILLER_34_1075 ();
 sg13g2_fill_1 FILLER_34_1077 ();
 sg13g2_decap_8 FILLER_34_1108 ();
 sg13g2_decap_8 FILLER_34_1115 ();
 sg13g2_fill_1 FILLER_34_1173 ();
 sg13g2_fill_1 FILLER_34_1258 ();
 sg13g2_fill_1 FILLER_34_1276 ();
 sg13g2_fill_2 FILLER_34_1290 ();
 sg13g2_decap_8 FILLER_34_1347 ();
 sg13g2_decap_8 FILLER_34_1354 ();
 sg13g2_decap_8 FILLER_34_1361 ();
 sg13g2_fill_2 FILLER_34_1368 ();
 sg13g2_decap_8 FILLER_34_1391 ();
 sg13g2_decap_4 FILLER_34_1398 ();
 sg13g2_fill_1 FILLER_34_1454 ();
 sg13g2_decap_8 FILLER_34_1462 ();
 sg13g2_decap_8 FILLER_34_1469 ();
 sg13g2_decap_4 FILLER_34_1476 ();
 sg13g2_fill_2 FILLER_34_1480 ();
 sg13g2_fill_1 FILLER_34_1492 ();
 sg13g2_fill_1 FILLER_34_1514 ();
 sg13g2_fill_1 FILLER_34_1540 ();
 sg13g2_fill_1 FILLER_34_1572 ();
 sg13g2_fill_2 FILLER_34_1584 ();
 sg13g2_fill_1 FILLER_34_1595 ();
 sg13g2_decap_8 FILLER_34_1604 ();
 sg13g2_decap_8 FILLER_34_1611 ();
 sg13g2_decap_4 FILLER_34_1618 ();
 sg13g2_fill_2 FILLER_34_1622 ();
 sg13g2_fill_1 FILLER_34_1653 ();
 sg13g2_fill_1 FILLER_34_1658 ();
 sg13g2_fill_2 FILLER_34_1663 ();
 sg13g2_fill_1 FILLER_34_1665 ();
 sg13g2_decap_8 FILLER_34_1692 ();
 sg13g2_fill_1 FILLER_34_1711 ();
 sg13g2_fill_2 FILLER_34_1733 ();
 sg13g2_fill_1 FILLER_34_1781 ();
 sg13g2_fill_2 FILLER_34_1789 ();
 sg13g2_fill_1 FILLER_34_1803 ();
 sg13g2_fill_1 FILLER_34_1813 ();
 sg13g2_fill_2 FILLER_34_1835 ();
 sg13g2_fill_2 FILLER_34_1847 ();
 sg13g2_fill_2 FILLER_34_1852 ();
 sg13g2_fill_1 FILLER_34_1857 ();
 sg13g2_fill_1 FILLER_34_1898 ();
 sg13g2_fill_2 FILLER_34_1978 ();
 sg13g2_fill_1 FILLER_34_1992 ();
 sg13g2_fill_2 FILLER_34_1998 ();
 sg13g2_fill_1 FILLER_34_2022 ();
 sg13g2_fill_2 FILLER_34_2068 ();
 sg13g2_fill_1 FILLER_34_2105 ();
 sg13g2_decap_8 FILLER_34_2139 ();
 sg13g2_decap_8 FILLER_34_2146 ();
 sg13g2_decap_8 FILLER_34_2153 ();
 sg13g2_fill_2 FILLER_34_2175 ();
 sg13g2_fill_1 FILLER_34_2193 ();
 sg13g2_fill_1 FILLER_34_2199 ();
 sg13g2_decap_4 FILLER_34_2207 ();
 sg13g2_fill_1 FILLER_34_2211 ();
 sg13g2_fill_1 FILLER_34_2222 ();
 sg13g2_decap_4 FILLER_34_2228 ();
 sg13g2_fill_1 FILLER_34_2232 ();
 sg13g2_decap_4 FILLER_34_2247 ();
 sg13g2_fill_1 FILLER_34_2251 ();
 sg13g2_fill_2 FILLER_34_2257 ();
 sg13g2_fill_1 FILLER_34_2259 ();
 sg13g2_decap_4 FILLER_34_2264 ();
 sg13g2_fill_2 FILLER_34_2281 ();
 sg13g2_fill_2 FILLER_34_2310 ();
 sg13g2_decap_4 FILLER_34_2329 ();
 sg13g2_decap_8 FILLER_34_2337 ();
 sg13g2_decap_8 FILLER_34_2344 ();
 sg13g2_decap_8 FILLER_34_2351 ();
 sg13g2_fill_1 FILLER_34_2358 ();
 sg13g2_fill_1 FILLER_34_2369 ();
 sg13g2_decap_4 FILLER_34_2391 ();
 sg13g2_fill_1 FILLER_34_2395 ();
 sg13g2_fill_2 FILLER_34_2455 ();
 sg13g2_fill_1 FILLER_34_2457 ();
 sg13g2_fill_1 FILLER_34_2463 ();
 sg13g2_fill_2 FILLER_34_2496 ();
 sg13g2_fill_1 FILLER_34_2506 ();
 sg13g2_fill_2 FILLER_34_2511 ();
 sg13g2_fill_1 FILLER_34_2513 ();
 sg13g2_decap_8 FILLER_34_2519 ();
 sg13g2_decap_4 FILLER_34_2526 ();
 sg13g2_fill_2 FILLER_34_2530 ();
 sg13g2_decap_8 FILLER_34_2541 ();
 sg13g2_decap_8 FILLER_34_2548 ();
 sg13g2_decap_8 FILLER_34_2555 ();
 sg13g2_decap_4 FILLER_34_2562 ();
 sg13g2_fill_1 FILLER_34_2566 ();
 sg13g2_decap_8 FILLER_34_2580 ();
 sg13g2_fill_2 FILLER_34_2587 ();
 sg13g2_fill_1 FILLER_34_2589 ();
 sg13g2_fill_1 FILLER_34_2621 ();
 sg13g2_fill_2 FILLER_34_2630 ();
 sg13g2_decap_8 FILLER_34_2661 ();
 sg13g2_fill_2 FILLER_34_2668 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_47 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_decap_8 FILLER_35_108 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_117 ();
 sg13g2_decap_4 FILLER_35_122 ();
 sg13g2_fill_2 FILLER_35_126 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_229 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_2 FILLER_35_262 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_277 ();
 sg13g2_fill_2 FILLER_35_282 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_289 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_361 ();
 sg13g2_decap_4 FILLER_35_370 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_fill_2 FILLER_35_387 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_395 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_2 FILLER_35_408 ();
 sg13g2_fill_2 FILLER_35_492 ();
 sg13g2_decap_8 FILLER_35_520 ();
 sg13g2_decap_8 FILLER_35_527 ();
 sg13g2_decap_8 FILLER_35_534 ();
 sg13g2_fill_2 FILLER_35_541 ();
 sg13g2_decap_8 FILLER_35_552 ();
 sg13g2_decap_8 FILLER_35_559 ();
 sg13g2_fill_2 FILLER_35_566 ();
 sg13g2_decap_8 FILLER_35_611 ();
 sg13g2_decap_4 FILLER_35_622 ();
 sg13g2_fill_1 FILLER_35_626 ();
 sg13g2_fill_1 FILLER_35_653 ();
 sg13g2_fill_2 FILLER_35_661 ();
 sg13g2_fill_2 FILLER_35_698 ();
 sg13g2_fill_1 FILLER_35_700 ();
 sg13g2_fill_2 FILLER_35_705 ();
 sg13g2_fill_1 FILLER_35_707 ();
 sg13g2_fill_2 FILLER_35_768 ();
 sg13g2_fill_2 FILLER_35_779 ();
 sg13g2_fill_1 FILLER_35_809 ();
 sg13g2_fill_1 FILLER_35_817 ();
 sg13g2_fill_2 FILLER_35_898 ();
 sg13g2_decap_8 FILLER_35_905 ();
 sg13g2_fill_1 FILLER_35_942 ();
 sg13g2_fill_1 FILLER_35_994 ();
 sg13g2_fill_1 FILLER_35_999 ();
 sg13g2_decap_8 FILLER_35_1033 ();
 sg13g2_decap_8 FILLER_35_1040 ();
 sg13g2_fill_2 FILLER_35_1072 ();
 sg13g2_fill_2 FILLER_35_1122 ();
 sg13g2_fill_1 FILLER_35_1124 ();
 sg13g2_fill_1 FILLER_35_1160 ();
 sg13g2_fill_2 FILLER_35_1184 ();
 sg13g2_fill_2 FILLER_35_1201 ();
 sg13g2_fill_1 FILLER_35_1203 ();
 sg13g2_fill_1 FILLER_35_1208 ();
 sg13g2_fill_2 FILLER_35_1215 ();
 sg13g2_fill_2 FILLER_35_1234 ();
 sg13g2_decap_4 FILLER_35_1239 ();
 sg13g2_fill_2 FILLER_35_1243 ();
 sg13g2_decap_8 FILLER_35_1249 ();
 sg13g2_fill_2 FILLER_35_1256 ();
 sg13g2_fill_1 FILLER_35_1258 ();
 sg13g2_fill_1 FILLER_35_1271 ();
 sg13g2_fill_1 FILLER_35_1281 ();
 sg13g2_fill_2 FILLER_35_1326 ();
 sg13g2_decap_8 FILLER_35_1340 ();
 sg13g2_fill_2 FILLER_35_1347 ();
 sg13g2_fill_1 FILLER_35_1349 ();
 sg13g2_decap_8 FILLER_35_1371 ();
 sg13g2_fill_1 FILLER_35_1399 ();
 sg13g2_decap_4 FILLER_35_1456 ();
 sg13g2_fill_2 FILLER_35_1499 ();
 sg13g2_fill_2 FILLER_35_1510 ();
 sg13g2_fill_1 FILLER_35_1524 ();
 sg13g2_fill_1 FILLER_35_1540 ();
 sg13g2_decap_4 FILLER_35_1599 ();
 sg13g2_fill_1 FILLER_35_1603 ();
 sg13g2_fill_2 FILLER_35_1625 ();
 sg13g2_fill_1 FILLER_35_1627 ();
 sg13g2_fill_1 FILLER_35_1654 ();
 sg13g2_fill_2 FILLER_35_1759 ();
 sg13g2_fill_1 FILLER_35_1771 ();
 sg13g2_fill_2 FILLER_35_1775 ();
 sg13g2_fill_1 FILLER_35_1794 ();
 sg13g2_fill_2 FILLER_35_1812 ();
 sg13g2_fill_1 FILLER_35_1853 ();
 sg13g2_fill_1 FILLER_35_1864 ();
 sg13g2_fill_1 FILLER_35_1891 ();
 sg13g2_fill_2 FILLER_35_1931 ();
 sg13g2_fill_1 FILLER_35_1938 ();
 sg13g2_fill_1 FILLER_35_1956 ();
 sg13g2_fill_2 FILLER_35_1961 ();
 sg13g2_fill_1 FILLER_35_1968 ();
 sg13g2_fill_1 FILLER_35_1994 ();
 sg13g2_fill_2 FILLER_35_2000 ();
 sg13g2_fill_1 FILLER_35_2032 ();
 sg13g2_fill_1 FILLER_35_2041 ();
 sg13g2_decap_8 FILLER_35_2075 ();
 sg13g2_decap_4 FILLER_35_2082 ();
 sg13g2_decap_8 FILLER_35_2090 ();
 sg13g2_decap_8 FILLER_35_2097 ();
 sg13g2_decap_8 FILLER_35_2104 ();
 sg13g2_decap_8 FILLER_35_2111 ();
 sg13g2_decap_8 FILLER_35_2118 ();
 sg13g2_decap_8 FILLER_35_2125 ();
 sg13g2_decap_8 FILLER_35_2132 ();
 sg13g2_decap_8 FILLER_35_2139 ();
 sg13g2_decap_8 FILLER_35_2146 ();
 sg13g2_decap_4 FILLER_35_2153 ();
 sg13g2_fill_2 FILLER_35_2170 ();
 sg13g2_fill_1 FILLER_35_2183 ();
 sg13g2_fill_1 FILLER_35_2212 ();
 sg13g2_fill_2 FILLER_35_2218 ();
 sg13g2_fill_1 FILLER_35_2241 ();
 sg13g2_fill_1 FILLER_35_2262 ();
 sg13g2_decap_8 FILLER_35_2268 ();
 sg13g2_decap_8 FILLER_35_2275 ();
 sg13g2_decap_8 FILLER_35_2282 ();
 sg13g2_fill_1 FILLER_35_2306 ();
 sg13g2_fill_2 FILLER_35_2311 ();
 sg13g2_decap_4 FILLER_35_2322 ();
 sg13g2_fill_2 FILLER_35_2326 ();
 sg13g2_decap_8 FILLER_35_2337 ();
 sg13g2_fill_1 FILLER_35_2344 ();
 sg13g2_fill_2 FILLER_35_2349 ();
 sg13g2_decap_8 FILLER_35_2392 ();
 sg13g2_decap_8 FILLER_35_2399 ();
 sg13g2_decap_4 FILLER_35_2406 ();
 sg13g2_fill_2 FILLER_35_2410 ();
 sg13g2_decap_8 FILLER_35_2424 ();
 sg13g2_fill_1 FILLER_35_2431 ();
 sg13g2_decap_8 FILLER_35_2450 ();
 sg13g2_fill_2 FILLER_35_2457 ();
 sg13g2_fill_1 FILLER_35_2476 ();
 sg13g2_decap_8 FILLER_35_2503 ();
 sg13g2_fill_1 FILLER_35_2510 ();
 sg13g2_fill_2 FILLER_35_2533 ();
 sg13g2_fill_1 FILLER_35_2535 ();
 sg13g2_decap_8 FILLER_35_2549 ();
 sg13g2_decap_8 FILLER_35_2556 ();
 sg13g2_fill_2 FILLER_35_2563 ();
 sg13g2_decap_8 FILLER_35_2663 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_decap_8 FILLER_36_16 ();
 sg13g2_fill_2 FILLER_36_75 ();
 sg13g2_fill_1 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_decap_4 FILLER_36_136 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_fill_1 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_243 ();
 sg13g2_fill_1 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_250 ();
 sg13g2_decap_4 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_decap_4 FILLER_36_407 ();
 sg13g2_fill_1 FILLER_36_411 ();
 sg13g2_fill_1 FILLER_36_490 ();
 sg13g2_fill_2 FILLER_36_516 ();
 sg13g2_fill_1 FILLER_36_522 ();
 sg13g2_fill_2 FILLER_36_570 ();
 sg13g2_fill_2 FILLER_36_590 ();
 sg13g2_fill_1 FILLER_36_618 ();
 sg13g2_decap_4 FILLER_36_660 ();
 sg13g2_fill_1 FILLER_36_664 ();
 sg13g2_fill_1 FILLER_36_691 ();
 sg13g2_fill_2 FILLER_36_710 ();
 sg13g2_fill_2 FILLER_36_729 ();
 sg13g2_fill_1 FILLER_36_731 ();
 sg13g2_fill_2 FILLER_36_780 ();
 sg13g2_fill_1 FILLER_36_789 ();
 sg13g2_fill_2 FILLER_36_819 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_fill_1 FILLER_36_862 ();
 sg13g2_fill_2 FILLER_36_893 ();
 sg13g2_fill_1 FILLER_36_895 ();
 sg13g2_fill_2 FILLER_36_904 ();
 sg13g2_fill_1 FILLER_36_906 ();
 sg13g2_fill_2 FILLER_36_971 ();
 sg13g2_fill_2 FILLER_36_986 ();
 sg13g2_fill_2 FILLER_36_1017 ();
 sg13g2_fill_1 FILLER_36_1053 ();
 sg13g2_decap_8 FILLER_36_1085 ();
 sg13g2_fill_2 FILLER_36_1092 ();
 sg13g2_fill_2 FILLER_36_1115 ();
 sg13g2_fill_1 FILLER_36_1117 ();
 sg13g2_fill_1 FILLER_36_1144 ();
 sg13g2_fill_2 FILLER_36_1189 ();
 sg13g2_fill_2 FILLER_36_1195 ();
 sg13g2_fill_2 FILLER_36_1201 ();
 sg13g2_fill_1 FILLER_36_1203 ();
 sg13g2_fill_2 FILLER_36_1266 ();
 sg13g2_fill_1 FILLER_36_1268 ();
 sg13g2_fill_1 FILLER_36_1307 ();
 sg13g2_fill_2 FILLER_36_1326 ();
 sg13g2_fill_1 FILLER_36_1332 ();
 sg13g2_fill_1 FILLER_36_1359 ();
 sg13g2_fill_1 FILLER_36_1364 ();
 sg13g2_fill_1 FILLER_36_1370 ();
 sg13g2_fill_1 FILLER_36_1397 ();
 sg13g2_fill_2 FILLER_36_1402 ();
 sg13g2_fill_2 FILLER_36_1444 ();
 sg13g2_decap_4 FILLER_36_1450 ();
 sg13g2_fill_1 FILLER_36_1454 ();
 sg13g2_fill_1 FILLER_36_1485 ();
 sg13g2_fill_2 FILLER_36_1527 ();
 sg13g2_fill_1 FILLER_36_1529 ();
 sg13g2_fill_2 FILLER_36_1549 ();
 sg13g2_fill_1 FILLER_36_1559 ();
 sg13g2_fill_1 FILLER_36_1564 ();
 sg13g2_fill_1 FILLER_36_1586 ();
 sg13g2_fill_2 FILLER_36_1613 ();
 sg13g2_fill_1 FILLER_36_1615 ();
 sg13g2_fill_1 FILLER_36_1648 ();
 sg13g2_fill_2 FILLER_36_1670 ();
 sg13g2_fill_2 FILLER_36_1676 ();
 sg13g2_fill_2 FILLER_36_1739 ();
 sg13g2_fill_1 FILLER_36_1741 ();
 sg13g2_fill_2 FILLER_36_1808 ();
 sg13g2_fill_1 FILLER_36_1815 ();
 sg13g2_fill_1 FILLER_36_1882 ();
 sg13g2_fill_1 FILLER_36_1887 ();
 sg13g2_fill_2 FILLER_36_1893 ();
 sg13g2_fill_2 FILLER_36_1979 ();
 sg13g2_fill_1 FILLER_36_1998 ();
 sg13g2_fill_2 FILLER_36_2030 ();
 sg13g2_fill_1 FILLER_36_2062 ();
 sg13g2_decap_8 FILLER_36_2085 ();
 sg13g2_decap_8 FILLER_36_2092 ();
 sg13g2_decap_8 FILLER_36_2099 ();
 sg13g2_decap_4 FILLER_36_2106 ();
 sg13g2_fill_1 FILLER_36_2110 ();
 sg13g2_fill_2 FILLER_36_2120 ();
 sg13g2_decap_4 FILLER_36_2148 ();
 sg13g2_fill_1 FILLER_36_2152 ();
 sg13g2_fill_2 FILLER_36_2172 ();
 sg13g2_decap_8 FILLER_36_2191 ();
 sg13g2_decap_8 FILLER_36_2198 ();
 sg13g2_decap_4 FILLER_36_2205 ();
 sg13g2_fill_2 FILLER_36_2209 ();
 sg13g2_fill_1 FILLER_36_2216 ();
 sg13g2_decap_4 FILLER_36_2226 ();
 sg13g2_fill_1 FILLER_36_2230 ();
 sg13g2_fill_2 FILLER_36_2238 ();
 sg13g2_fill_1 FILLER_36_2240 ();
 sg13g2_fill_2 FILLER_36_2275 ();
 sg13g2_decap_8 FILLER_36_2290 ();
 sg13g2_decap_8 FILLER_36_2297 ();
 sg13g2_decap_8 FILLER_36_2304 ();
 sg13g2_decap_4 FILLER_36_2311 ();
 sg13g2_fill_2 FILLER_36_2315 ();
 sg13g2_fill_2 FILLER_36_2327 ();
 sg13g2_fill_2 FILLER_36_2342 ();
 sg13g2_fill_1 FILLER_36_2344 ();
 sg13g2_decap_8 FILLER_36_2372 ();
 sg13g2_fill_2 FILLER_36_2379 ();
 sg13g2_fill_1 FILLER_36_2381 ();
 sg13g2_fill_2 FILLER_36_2400 ();
 sg13g2_fill_1 FILLER_36_2402 ();
 sg13g2_fill_2 FILLER_36_2411 ();
 sg13g2_fill_2 FILLER_36_2418 ();
 sg13g2_decap_4 FILLER_36_2435 ();
 sg13g2_fill_1 FILLER_36_2439 ();
 sg13g2_fill_1 FILLER_36_2448 ();
 sg13g2_decap_8 FILLER_36_2478 ();
 sg13g2_fill_1 FILLER_36_2485 ();
 sg13g2_decap_8 FILLER_36_2490 ();
 sg13g2_fill_2 FILLER_36_2497 ();
 sg13g2_decap_8 FILLER_36_2517 ();
 sg13g2_fill_2 FILLER_36_2524 ();
 sg13g2_fill_1 FILLER_36_2530 ();
 sg13g2_decap_4 FILLER_36_2548 ();
 sg13g2_fill_2 FILLER_36_2552 ();
 sg13g2_fill_1 FILLER_36_2559 ();
 sg13g2_decap_4 FILLER_36_2609 ();
 sg13g2_decap_8 FILLER_36_2662 ();
 sg13g2_fill_1 FILLER_36_2669 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_33 ();
 sg13g2_fill_2 FILLER_37_40 ();
 sg13g2_decap_8 FILLER_37_46 ();
 sg13g2_decap_4 FILLER_37_53 ();
 sg13g2_decap_8 FILLER_37_76 ();
 sg13g2_decap_4 FILLER_37_83 ();
 sg13g2_fill_2 FILLER_37_104 ();
 sg13g2_fill_1 FILLER_37_115 ();
 sg13g2_fill_2 FILLER_37_121 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_fill_2 FILLER_37_154 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_fill_1 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_200 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_decap_8 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_251 ();
 sg13g2_decap_4 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_298 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_411 ();
 sg13g2_decap_4 FILLER_37_418 ();
 sg13g2_fill_1 FILLER_37_422 ();
 sg13g2_fill_2 FILLER_37_436 ();
 sg13g2_fill_2 FILLER_37_452 ();
 sg13g2_fill_1 FILLER_37_537 ();
 sg13g2_fill_1 FILLER_37_641 ();
 sg13g2_fill_1 FILLER_37_650 ();
 sg13g2_fill_1 FILLER_37_681 ();
 sg13g2_fill_2 FILLER_37_737 ();
 sg13g2_fill_1 FILLER_37_773 ();
 sg13g2_fill_2 FILLER_37_779 ();
 sg13g2_fill_1 FILLER_37_807 ();
 sg13g2_decap_4 FILLER_37_857 ();
 sg13g2_decap_4 FILLER_37_865 ();
 sg13g2_fill_2 FILLER_37_869 ();
 sg13g2_decap_8 FILLER_37_879 ();
 sg13g2_decap_8 FILLER_37_929 ();
 sg13g2_fill_2 FILLER_37_936 ();
 sg13g2_fill_1 FILLER_37_938 ();
 sg13g2_decap_4 FILLER_37_953 ();
 sg13g2_fill_1 FILLER_37_957 ();
 sg13g2_decap_4 FILLER_37_961 ();
 sg13g2_fill_1 FILLER_37_965 ();
 sg13g2_fill_1 FILLER_37_1020 ();
 sg13g2_fill_1 FILLER_37_1118 ();
 sg13g2_fill_2 FILLER_37_1165 ();
 sg13g2_fill_1 FILLER_37_1173 ();
 sg13g2_fill_1 FILLER_37_1177 ();
 sg13g2_fill_1 FILLER_37_1183 ();
 sg13g2_fill_1 FILLER_37_1189 ();
 sg13g2_fill_2 FILLER_37_1195 ();
 sg13g2_fill_2 FILLER_37_1201 ();
 sg13g2_fill_1 FILLER_37_1207 ();
 sg13g2_fill_2 FILLER_37_1269 ();
 sg13g2_fill_1 FILLER_37_1346 ();
 sg13g2_fill_2 FILLER_37_1373 ();
 sg13g2_fill_1 FILLER_37_1375 ();
 sg13g2_fill_1 FILLER_37_1383 ();
 sg13g2_decap_8 FILLER_37_1449 ();
 sg13g2_fill_1 FILLER_37_1456 ();
 sg13g2_fill_2 FILLER_37_1462 ();
 sg13g2_fill_1 FILLER_37_1464 ();
 sg13g2_fill_1 FILLER_37_1473 ();
 sg13g2_fill_1 FILLER_37_1479 ();
 sg13g2_fill_1 FILLER_37_1484 ();
 sg13g2_fill_2 FILLER_37_1489 ();
 sg13g2_fill_2 FILLER_37_1529 ();
 sg13g2_fill_1 FILLER_37_1531 ();
 sg13g2_fill_1 FILLER_37_1558 ();
 sg13g2_fill_1 FILLER_37_1568 ();
 sg13g2_fill_1 FILLER_37_1577 ();
 sg13g2_fill_2 FILLER_37_1643 ();
 sg13g2_decap_8 FILLER_37_1649 ();
 sg13g2_fill_2 FILLER_37_1656 ();
 sg13g2_fill_1 FILLER_37_1658 ();
 sg13g2_fill_2 FILLER_37_1684 ();
 sg13g2_fill_1 FILLER_37_1707 ();
 sg13g2_decap_8 FILLER_37_1733 ();
 sg13g2_fill_2 FILLER_37_1740 ();
 sg13g2_fill_1 FILLER_37_1756 ();
 sg13g2_fill_2 FILLER_37_1803 ();
 sg13g2_fill_2 FILLER_37_1836 ();
 sg13g2_fill_1 FILLER_37_1846 ();
 sg13g2_fill_2 FILLER_37_1855 ();
 sg13g2_fill_1 FILLER_37_1874 ();
 sg13g2_fill_1 FILLER_37_1879 ();
 sg13g2_fill_1 FILLER_37_1885 ();
 sg13g2_fill_2 FILLER_37_1907 ();
 sg13g2_fill_1 FILLER_37_1919 ();
 sg13g2_fill_2 FILLER_37_1962 ();
 sg13g2_fill_1 FILLER_37_1974 ();
 sg13g2_fill_2 FILLER_37_1995 ();
 sg13g2_fill_1 FILLER_37_2046 ();
 sg13g2_fill_1 FILLER_37_2068 ();
 sg13g2_decap_4 FILLER_37_2073 ();
 sg13g2_fill_1 FILLER_37_2077 ();
 sg13g2_fill_1 FILLER_37_2116 ();
 sg13g2_decap_8 FILLER_37_2143 ();
 sg13g2_decap_4 FILLER_37_2150 ();
 sg13g2_fill_2 FILLER_37_2154 ();
 sg13g2_fill_2 FILLER_37_2169 ();
 sg13g2_fill_1 FILLER_37_2171 ();
 sg13g2_decap_4 FILLER_37_2198 ();
 sg13g2_fill_1 FILLER_37_2202 ();
 sg13g2_decap_8 FILLER_37_2206 ();
 sg13g2_decap_8 FILLER_37_2213 ();
 sg13g2_decap_8 FILLER_37_2220 ();
 sg13g2_decap_8 FILLER_37_2227 ();
 sg13g2_fill_1 FILLER_37_2259 ();
 sg13g2_fill_2 FILLER_37_2264 ();
 sg13g2_fill_1 FILLER_37_2272 ();
 sg13g2_decap_8 FILLER_37_2278 ();
 sg13g2_fill_1 FILLER_37_2285 ();
 sg13g2_decap_8 FILLER_37_2312 ();
 sg13g2_decap_8 FILLER_37_2319 ();
 sg13g2_decap_4 FILLER_37_2326 ();
 sg13g2_fill_1 FILLER_37_2341 ();
 sg13g2_decap_8 FILLER_37_2357 ();
 sg13g2_fill_2 FILLER_37_2372 ();
 sg13g2_fill_2 FILLER_37_2382 ();
 sg13g2_decap_4 FILLER_37_2397 ();
 sg13g2_fill_2 FILLER_37_2401 ();
 sg13g2_decap_4 FILLER_37_2408 ();
 sg13g2_fill_2 FILLER_37_2412 ();
 sg13g2_fill_1 FILLER_37_2422 ();
 sg13g2_fill_2 FILLER_37_2427 ();
 sg13g2_fill_1 FILLER_37_2435 ();
 sg13g2_fill_1 FILLER_37_2440 ();
 sg13g2_decap_8 FILLER_37_2451 ();
 sg13g2_decap_8 FILLER_37_2458 ();
 sg13g2_decap_8 FILLER_37_2465 ();
 sg13g2_decap_8 FILLER_37_2472 ();
 sg13g2_decap_8 FILLER_37_2479 ();
 sg13g2_decap_8 FILLER_37_2486 ();
 sg13g2_fill_2 FILLER_37_2493 ();
 sg13g2_fill_1 FILLER_37_2495 ();
 sg13g2_decap_4 FILLER_37_2520 ();
 sg13g2_fill_1 FILLER_37_2524 ();
 sg13g2_fill_2 FILLER_37_2530 ();
 sg13g2_fill_1 FILLER_37_2532 ();
 sg13g2_fill_1 FILLER_37_2555 ();
 sg13g2_fill_1 FILLER_37_2593 ();
 sg13g2_decap_8 FILLER_37_2604 ();
 sg13g2_decap_4 FILLER_37_2611 ();
 sg13g2_fill_2 FILLER_37_2615 ();
 sg13g2_fill_1 FILLER_37_2629 ();
 sg13g2_fill_2 FILLER_37_2634 ();
 sg13g2_fill_1 FILLER_37_2636 ();
 sg13g2_decap_8 FILLER_37_2663 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_13 ();
 sg13g2_fill_2 FILLER_38_20 ();
 sg13g2_decap_8 FILLER_38_26 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_135 ();
 sg13g2_decap_8 FILLER_38_142 ();
 sg13g2_decap_4 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_fill_2 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_309 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_decap_4 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_405 ();
 sg13g2_fill_2 FILLER_38_456 ();
 sg13g2_fill_1 FILLER_38_495 ();
 sg13g2_fill_1 FILLER_38_506 ();
 sg13g2_fill_1 FILLER_38_537 ();
 sg13g2_fill_1 FILLER_38_543 ();
 sg13g2_fill_2 FILLER_38_666 ();
 sg13g2_fill_2 FILLER_38_672 ();
 sg13g2_decap_8 FILLER_38_678 ();
 sg13g2_fill_2 FILLER_38_750 ();
 sg13g2_fill_2 FILLER_38_781 ();
 sg13g2_fill_2 FILLER_38_845 ();
 sg13g2_decap_4 FILLER_38_853 ();
 sg13g2_fill_1 FILLER_38_857 ();
 sg13g2_fill_2 FILLER_38_871 ();
 sg13g2_fill_1 FILLER_38_894 ();
 sg13g2_decap_4 FILLER_38_908 ();
 sg13g2_decap_8 FILLER_38_916 ();
 sg13g2_decap_8 FILLER_38_923 ();
 sg13g2_decap_8 FILLER_38_930 ();
 sg13g2_fill_2 FILLER_38_937 ();
 sg13g2_fill_1 FILLER_38_943 ();
 sg13g2_fill_2 FILLER_38_982 ();
 sg13g2_fill_1 FILLER_38_984 ();
 sg13g2_fill_1 FILLER_38_992 ();
 sg13g2_fill_2 FILLER_38_1023 ();
 sg13g2_fill_2 FILLER_38_1053 ();
 sg13g2_fill_1 FILLER_38_1063 ();
 sg13g2_fill_1 FILLER_38_1104 ();
 sg13g2_fill_1 FILLER_38_1132 ();
 sg13g2_fill_2 FILLER_38_1162 ();
 sg13g2_fill_1 FILLER_38_1169 ();
 sg13g2_fill_1 FILLER_38_1173 ();
 sg13g2_fill_2 FILLER_38_1234 ();
 sg13g2_fill_2 FILLER_38_1240 ();
 sg13g2_fill_1 FILLER_38_1282 ();
 sg13g2_fill_2 FILLER_38_1292 ();
 sg13g2_fill_2 FILLER_38_1301 ();
 sg13g2_fill_2 FILLER_38_1310 ();
 sg13g2_fill_2 FILLER_38_1318 ();
 sg13g2_fill_2 FILLER_38_1326 ();
 sg13g2_fill_1 FILLER_38_1337 ();
 sg13g2_decap_4 FILLER_38_1342 ();
 sg13g2_fill_1 FILLER_38_1346 ();
 sg13g2_fill_2 FILLER_38_1368 ();
 sg13g2_fill_1 FILLER_38_1375 ();
 sg13g2_fill_2 FILLER_38_1413 ();
 sg13g2_fill_1 FILLER_38_1415 ();
 sg13g2_fill_1 FILLER_38_1442 ();
 sg13g2_fill_1 FILLER_38_1473 ();
 sg13g2_fill_1 FILLER_38_1570 ();
 sg13g2_fill_1 FILLER_38_1586 ();
 sg13g2_fill_2 FILLER_38_1591 ();
 sg13g2_fill_1 FILLER_38_1606 ();
 sg13g2_fill_2 FILLER_38_1631 ();
 sg13g2_decap_8 FILLER_38_1637 ();
 sg13g2_decap_8 FILLER_38_1644 ();
 sg13g2_fill_2 FILLER_38_1651 ();
 sg13g2_fill_2 FILLER_38_1657 ();
 sg13g2_decap_4 FILLER_38_1676 ();
 sg13g2_decap_8 FILLER_38_1684 ();
 sg13g2_decap_4 FILLER_38_1691 ();
 sg13g2_fill_2 FILLER_38_1718 ();
 sg13g2_fill_1 FILLER_38_1720 ();
 sg13g2_decap_4 FILLER_38_1747 ();
 sg13g2_fill_1 FILLER_38_1757 ();
 sg13g2_fill_1 FILLER_38_1768 ();
 sg13g2_fill_2 FILLER_38_1775 ();
 sg13g2_fill_2 FILLER_38_1876 ();
 sg13g2_fill_2 FILLER_38_1889 ();
 sg13g2_fill_1 FILLER_38_1921 ();
 sg13g2_fill_1 FILLER_38_1925 ();
 sg13g2_fill_1 FILLER_38_1929 ();
 sg13g2_fill_2 FILLER_38_1959 ();
 sg13g2_fill_2 FILLER_38_2040 ();
 sg13g2_fill_1 FILLER_38_2068 ();
 sg13g2_fill_1 FILLER_38_2074 ();
 sg13g2_decap_8 FILLER_38_2148 ();
 sg13g2_fill_1 FILLER_38_2155 ();
 sg13g2_decap_8 FILLER_38_2195 ();
 sg13g2_fill_2 FILLER_38_2202 ();
 sg13g2_fill_1 FILLER_38_2204 ();
 sg13g2_decap_4 FILLER_38_2218 ();
 sg13g2_fill_1 FILLER_38_2226 ();
 sg13g2_fill_1 FILLER_38_2236 ();
 sg13g2_fill_2 FILLER_38_2241 ();
 sg13g2_decap_8 FILLER_38_2270 ();
 sg13g2_decap_8 FILLER_38_2277 ();
 sg13g2_fill_1 FILLER_38_2284 ();
 sg13g2_decap_8 FILLER_38_2297 ();
 sg13g2_decap_4 FILLER_38_2304 ();
 sg13g2_decap_8 FILLER_38_2313 ();
 sg13g2_fill_2 FILLER_38_2320 ();
 sg13g2_fill_1 FILLER_38_2322 ();
 sg13g2_fill_2 FILLER_38_2357 ();
 sg13g2_fill_2 FILLER_38_2367 ();
 sg13g2_fill_1 FILLER_38_2394 ();
 sg13g2_fill_2 FILLER_38_2408 ();
 sg13g2_decap_8 FILLER_38_2415 ();
 sg13g2_decap_8 FILLER_38_2452 ();
 sg13g2_decap_8 FILLER_38_2459 ();
 sg13g2_decap_4 FILLER_38_2466 ();
 sg13g2_fill_2 FILLER_38_2470 ();
 sg13g2_decap_4 FILLER_38_2476 ();
 sg13g2_fill_1 FILLER_38_2502 ();
 sg13g2_decap_4 FILLER_38_2547 ();
 sg13g2_fill_2 FILLER_38_2575 ();
 sg13g2_fill_1 FILLER_38_2585 ();
 sg13g2_fill_2 FILLER_38_2608 ();
 sg13g2_fill_1 FILLER_38_2610 ();
 sg13g2_fill_1 FILLER_38_2619 ();
 sg13g2_decap_8 FILLER_38_2634 ();
 sg13g2_fill_2 FILLER_38_2641 ();
 sg13g2_decap_8 FILLER_38_2655 ();
 sg13g2_decap_8 FILLER_38_2662 ();
 sg13g2_fill_1 FILLER_38_2669 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_fill_1 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_45 ();
 sg13g2_fill_2 FILLER_39_52 ();
 sg13g2_fill_1 FILLER_39_54 ();
 sg13g2_fill_1 FILLER_39_94 ();
 sg13g2_fill_1 FILLER_39_99 ();
 sg13g2_fill_2 FILLER_39_109 ();
 sg13g2_fill_1 FILLER_39_115 ();
 sg13g2_fill_1 FILLER_39_125 ();
 sg13g2_fill_2 FILLER_39_152 ();
 sg13g2_fill_1 FILLER_39_162 ();
 sg13g2_fill_2 FILLER_39_218 ();
 sg13g2_decap_8 FILLER_39_251 ();
 sg13g2_decap_8 FILLER_39_258 ();
 sg13g2_decap_8 FILLER_39_302 ();
 sg13g2_fill_1 FILLER_39_313 ();
 sg13g2_decap_8 FILLER_39_401 ();
 sg13g2_decap_8 FILLER_39_408 ();
 sg13g2_fill_2 FILLER_39_415 ();
 sg13g2_fill_1 FILLER_39_448 ();
 sg13g2_fill_1 FILLER_39_482 ();
 sg13g2_fill_2 FILLER_39_492 ();
 sg13g2_fill_1 FILLER_39_514 ();
 sg13g2_fill_2 FILLER_39_519 ();
 sg13g2_fill_1 FILLER_39_542 ();
 sg13g2_fill_2 FILLER_39_551 ();
 sg13g2_fill_1 FILLER_39_604 ();
 sg13g2_fill_1 FILLER_39_609 ();
 sg13g2_fill_1 FILLER_39_615 ();
 sg13g2_fill_1 FILLER_39_620 ();
 sg13g2_fill_1 FILLER_39_647 ();
 sg13g2_fill_2 FILLER_39_657 ();
 sg13g2_fill_1 FILLER_39_659 ();
 sg13g2_fill_2 FILLER_39_690 ();
 sg13g2_fill_1 FILLER_39_692 ();
 sg13g2_decap_4 FILLER_39_726 ();
 sg13g2_fill_1 FILLER_39_730 ();
 sg13g2_decap_8 FILLER_39_738 ();
 sg13g2_fill_2 FILLER_39_745 ();
 sg13g2_decap_8 FILLER_39_772 ();
 sg13g2_decap_4 FILLER_39_779 ();
 sg13g2_fill_2 FILLER_39_787 ();
 sg13g2_fill_1 FILLER_39_789 ();
 sg13g2_decap_8 FILLER_39_794 ();
 sg13g2_decap_8 FILLER_39_801 ();
 sg13g2_decap_4 FILLER_39_808 ();
 sg13g2_fill_2 FILLER_39_847 ();
 sg13g2_fill_1 FILLER_39_849 ();
 sg13g2_fill_2 FILLER_39_867 ();
 sg13g2_fill_2 FILLER_39_874 ();
 sg13g2_fill_1 FILLER_39_876 ();
 sg13g2_fill_2 FILLER_39_907 ();
 sg13g2_fill_2 FILLER_39_914 ();
 sg13g2_fill_1 FILLER_39_921 ();
 sg13g2_fill_1 FILLER_39_930 ();
 sg13g2_fill_2 FILLER_39_940 ();
 sg13g2_fill_1 FILLER_39_942 ();
 sg13g2_fill_2 FILLER_39_948 ();
 sg13g2_fill_1 FILLER_39_950 ();
 sg13g2_fill_1 FILLER_39_960 ();
 sg13g2_decap_8 FILLER_39_965 ();
 sg13g2_decap_4 FILLER_39_972 ();
 sg13g2_fill_2 FILLER_39_976 ();
 sg13g2_fill_2 FILLER_39_1004 ();
 sg13g2_decap_8 FILLER_39_1010 ();
 sg13g2_fill_2 FILLER_39_1017 ();
 sg13g2_fill_1 FILLER_39_1027 ();
 sg13g2_fill_2 FILLER_39_1039 ();
 sg13g2_fill_2 FILLER_39_1079 ();
 sg13g2_fill_2 FILLER_39_1117 ();
 sg13g2_fill_2 FILLER_39_1140 ();
 sg13g2_fill_2 FILLER_39_1155 ();
 sg13g2_fill_2 FILLER_39_1164 ();
 sg13g2_fill_1 FILLER_39_1187 ();
 sg13g2_fill_1 FILLER_39_1192 ();
 sg13g2_fill_1 FILLER_39_1222 ();
 sg13g2_fill_1 FILLER_39_1244 ();
 sg13g2_fill_1 FILLER_39_1265 ();
 sg13g2_fill_1 FILLER_39_1282 ();
 sg13g2_fill_1 FILLER_39_1287 ();
 sg13g2_fill_2 FILLER_39_1317 ();
 sg13g2_fill_1 FILLER_39_1326 ();
 sg13g2_fill_2 FILLER_39_1366 ();
 sg13g2_fill_1 FILLER_39_1389 ();
 sg13g2_decap_4 FILLER_39_1436 ();
 sg13g2_fill_1 FILLER_39_1444 ();
 sg13g2_fill_1 FILLER_39_1501 ();
 sg13g2_fill_1 FILLER_39_1510 ();
 sg13g2_fill_1 FILLER_39_1515 ();
 sg13g2_fill_1 FILLER_39_1521 ();
 sg13g2_fill_2 FILLER_39_1527 ();
 sg13g2_fill_1 FILLER_39_1559 ();
 sg13g2_fill_1 FILLER_39_1573 ();
 sg13g2_fill_1 FILLER_39_1581 ();
 sg13g2_fill_2 FILLER_39_1591 ();
 sg13g2_fill_1 FILLER_39_1593 ();
 sg13g2_decap_4 FILLER_39_1623 ();
 sg13g2_fill_1 FILLER_39_1627 ();
 sg13g2_fill_1 FILLER_39_1664 ();
 sg13g2_fill_1 FILLER_39_1696 ();
 sg13g2_fill_1 FILLER_39_1741 ();
 sg13g2_fill_2 FILLER_39_1746 ();
 sg13g2_fill_1 FILLER_39_1748 ();
 sg13g2_fill_1 FILLER_39_1809 ();
 sg13g2_fill_1 FILLER_39_1854 ();
 sg13g2_fill_2 FILLER_39_1910 ();
 sg13g2_fill_1 FILLER_39_1921 ();
 sg13g2_fill_1 FILLER_39_1948 ();
 sg13g2_fill_1 FILLER_39_2028 ();
 sg13g2_fill_1 FILLER_39_2034 ();
 sg13g2_fill_2 FILLER_39_2049 ();
 sg13g2_fill_2 FILLER_39_2055 ();
 sg13g2_decap_4 FILLER_39_2061 ();
 sg13g2_fill_1 FILLER_39_2065 ();
 sg13g2_decap_4 FILLER_39_2078 ();
 sg13g2_fill_1 FILLER_39_2112 ();
 sg13g2_fill_2 FILLER_39_2149 ();
 sg13g2_fill_1 FILLER_39_2182 ();
 sg13g2_fill_1 FILLER_39_2188 ();
 sg13g2_fill_1 FILLER_39_2194 ();
 sg13g2_fill_2 FILLER_39_2203 ();
 sg13g2_fill_1 FILLER_39_2213 ();
 sg13g2_decap_8 FILLER_39_2261 ();
 sg13g2_decap_8 FILLER_39_2268 ();
 sg13g2_fill_2 FILLER_39_2275 ();
 sg13g2_decap_8 FILLER_39_2295 ();
 sg13g2_decap_8 FILLER_39_2302 ();
 sg13g2_decap_4 FILLER_39_2309 ();
 sg13g2_fill_2 FILLER_39_2313 ();
 sg13g2_decap_8 FILLER_39_2333 ();
 sg13g2_fill_2 FILLER_39_2340 ();
 sg13g2_fill_1 FILLER_39_2342 ();
 sg13g2_fill_2 FILLER_39_2357 ();
 sg13g2_fill_1 FILLER_39_2359 ();
 sg13g2_decap_8 FILLER_39_2368 ();
 sg13g2_decap_8 FILLER_39_2375 ();
 sg13g2_fill_1 FILLER_39_2382 ();
 sg13g2_fill_1 FILLER_39_2401 ();
 sg13g2_decap_4 FILLER_39_2410 ();
 sg13g2_fill_1 FILLER_39_2414 ();
 sg13g2_fill_1 FILLER_39_2423 ();
 sg13g2_fill_2 FILLER_39_2429 ();
 sg13g2_fill_2 FILLER_39_2435 ();
 sg13g2_decap_8 FILLER_39_2442 ();
 sg13g2_decap_8 FILLER_39_2449 ();
 sg13g2_decap_8 FILLER_39_2456 ();
 sg13g2_decap_4 FILLER_39_2463 ();
 sg13g2_fill_2 FILLER_39_2467 ();
 sg13g2_decap_8 FILLER_39_2473 ();
 sg13g2_decap_8 FILLER_39_2480 ();
 sg13g2_decap_8 FILLER_39_2487 ();
 sg13g2_fill_1 FILLER_39_2494 ();
 sg13g2_fill_1 FILLER_39_2523 ();
 sg13g2_fill_2 FILLER_39_2528 ();
 sg13g2_fill_1 FILLER_39_2530 ();
 sg13g2_fill_2 FILLER_39_2536 ();
 sg13g2_decap_8 FILLER_39_2542 ();
 sg13g2_decap_8 FILLER_39_2553 ();
 sg13g2_decap_4 FILLER_39_2560 ();
 sg13g2_fill_1 FILLER_39_2564 ();
 sg13g2_fill_1 FILLER_39_2569 ();
 sg13g2_decap_8 FILLER_39_2575 ();
 sg13g2_fill_2 FILLER_39_2582 ();
 sg13g2_fill_1 FILLER_39_2592 ();
 sg13g2_fill_1 FILLER_39_2597 ();
 sg13g2_decap_8 FILLER_39_2624 ();
 sg13g2_fill_2 FILLER_39_2635 ();
 sg13g2_decap_8 FILLER_39_2663 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_9 ();
 sg13g2_fill_2 FILLER_40_49 ();
 sg13g2_fill_2 FILLER_40_60 ();
 sg13g2_fill_2 FILLER_40_75 ();
 sg13g2_fill_1 FILLER_40_99 ();
 sg13g2_decap_8 FILLER_40_109 ();
 sg13g2_fill_2 FILLER_40_116 ();
 sg13g2_fill_2 FILLER_40_144 ();
 sg13g2_fill_1 FILLER_40_146 ();
 sg13g2_fill_2 FILLER_40_173 ();
 sg13g2_fill_1 FILLER_40_201 ();
 sg13g2_fill_2 FILLER_40_254 ();
 sg13g2_fill_1 FILLER_40_287 ();
 sg13g2_fill_2 FILLER_40_309 ();
 sg13g2_fill_1 FILLER_40_362 ();
 sg13g2_fill_1 FILLER_40_401 ();
 sg13g2_decap_4 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_418 ();
 sg13g2_fill_1 FILLER_40_457 ();
 sg13g2_fill_2 FILLER_40_463 ();
 sg13g2_fill_2 FILLER_40_495 ();
 sg13g2_fill_1 FILLER_40_508 ();
 sg13g2_fill_2 FILLER_40_519 ();
 sg13g2_fill_1 FILLER_40_537 ();
 sg13g2_fill_1 FILLER_40_542 ();
 sg13g2_fill_1 FILLER_40_547 ();
 sg13g2_fill_1 FILLER_40_622 ();
 sg13g2_fill_1 FILLER_40_632 ();
 sg13g2_fill_1 FILLER_40_637 ();
 sg13g2_decap_4 FILLER_40_664 ();
 sg13g2_fill_1 FILLER_40_668 ();
 sg13g2_decap_8 FILLER_40_699 ();
 sg13g2_decap_4 FILLER_40_706 ();
 sg13g2_fill_1 FILLER_40_710 ();
 sg13g2_fill_1 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_772 ();
 sg13g2_decap_8 FILLER_40_779 ();
 sg13g2_decap_8 FILLER_40_786 ();
 sg13g2_decap_8 FILLER_40_793 ();
 sg13g2_decap_8 FILLER_40_800 ();
 sg13g2_fill_2 FILLER_40_807 ();
 sg13g2_fill_1 FILLER_40_809 ();
 sg13g2_fill_2 FILLER_40_852 ();
 sg13g2_fill_2 FILLER_40_936 ();
 sg13g2_fill_2 FILLER_40_955 ();
 sg13g2_fill_1 FILLER_40_966 ();
 sg13g2_fill_1 FILLER_40_972 ();
 sg13g2_fill_1 FILLER_40_977 ();
 sg13g2_fill_1 FILLER_40_986 ();
 sg13g2_fill_1 FILLER_40_991 ();
 sg13g2_decap_4 FILLER_40_997 ();
 sg13g2_fill_1 FILLER_40_1001 ();
 sg13g2_decap_4 FILLER_40_1010 ();
 sg13g2_fill_1 FILLER_40_1014 ();
 sg13g2_fill_2 FILLER_40_1110 ();
 sg13g2_fill_2 FILLER_40_1117 ();
 sg13g2_fill_1 FILLER_40_1122 ();
 sg13g2_fill_1 FILLER_40_1157 ();
 sg13g2_fill_1 FILLER_40_1165 ();
 sg13g2_fill_1 FILLER_40_1178 ();
 sg13g2_fill_2 FILLER_40_1209 ();
 sg13g2_fill_2 FILLER_40_1266 ();
 sg13g2_fill_2 FILLER_40_1286 ();
 sg13g2_fill_2 FILLER_40_1292 ();
 sg13g2_fill_1 FILLER_40_1376 ();
 sg13g2_decap_8 FILLER_40_1389 ();
 sg13g2_decap_4 FILLER_40_1396 ();
 sg13g2_fill_1 FILLER_40_1407 ();
 sg13g2_fill_2 FILLER_40_1412 ();
 sg13g2_fill_1 FILLER_40_1414 ();
 sg13g2_decap_8 FILLER_40_1441 ();
 sg13g2_fill_2 FILLER_40_1448 ();
 sg13g2_decap_4 FILLER_40_1458 ();
 sg13g2_fill_1 FILLER_40_1462 ();
 sg13g2_fill_2 FILLER_40_1478 ();
 sg13g2_fill_1 FILLER_40_1480 ();
 sg13g2_fill_2 FILLER_40_1485 ();
 sg13g2_decap_8 FILLER_40_1513 ();
 sg13g2_fill_2 FILLER_40_1520 ();
 sg13g2_fill_1 FILLER_40_1522 ();
 sg13g2_fill_2 FILLER_40_1539 ();
 sg13g2_fill_1 FILLER_40_1541 ();
 sg13g2_fill_2 FILLER_40_1547 ();
 sg13g2_fill_2 FILLER_40_1582 ();
 sg13g2_fill_1 FILLER_40_1584 ();
 sg13g2_fill_1 FILLER_40_1611 ();
 sg13g2_fill_2 FILLER_40_1618 ();
 sg13g2_fill_1 FILLER_40_1692 ();
 sg13g2_fill_1 FILLER_40_1697 ();
 sg13g2_fill_2 FILLER_40_1767 ();
 sg13g2_fill_1 FILLER_40_1778 ();
 sg13g2_fill_2 FILLER_40_1790 ();
 sg13g2_fill_2 FILLER_40_1803 ();
 sg13g2_fill_2 FILLER_40_1841 ();
 sg13g2_fill_1 FILLER_40_1877 ();
 sg13g2_fill_1 FILLER_40_1899 ();
 sg13g2_fill_2 FILLER_40_1911 ();
 sg13g2_fill_1 FILLER_40_1925 ();
 sg13g2_fill_1 FILLER_40_1929 ();
 sg13g2_fill_1 FILLER_40_2034 ();
 sg13g2_fill_2 FILLER_40_2039 ();
 sg13g2_fill_2 FILLER_40_2055 ();
 sg13g2_fill_2 FILLER_40_2069 ();
 sg13g2_fill_1 FILLER_40_2076 ();
 sg13g2_decap_8 FILLER_40_2139 ();
 sg13g2_decap_8 FILLER_40_2146 ();
 sg13g2_fill_1 FILLER_40_2153 ();
 sg13g2_decap_4 FILLER_40_2162 ();
 sg13g2_decap_4 FILLER_40_2198 ();
 sg13g2_fill_1 FILLER_40_2202 ();
 sg13g2_fill_2 FILLER_40_2219 ();
 sg13g2_fill_1 FILLER_40_2221 ();
 sg13g2_fill_1 FILLER_40_2227 ();
 sg13g2_fill_1 FILLER_40_2240 ();
 sg13g2_fill_2 FILLER_40_2245 ();
 sg13g2_decap_8 FILLER_40_2252 ();
 sg13g2_decap_8 FILLER_40_2259 ();
 sg13g2_decap_8 FILLER_40_2266 ();
 sg13g2_fill_2 FILLER_40_2273 ();
 sg13g2_fill_1 FILLER_40_2275 ();
 sg13g2_decap_4 FILLER_40_2288 ();
 sg13g2_fill_1 FILLER_40_2296 ();
 sg13g2_decap_8 FILLER_40_2301 ();
 sg13g2_decap_4 FILLER_40_2308 ();
 sg13g2_decap_8 FILLER_40_2316 ();
 sg13g2_fill_2 FILLER_40_2323 ();
 sg13g2_decap_8 FILLER_40_2346 ();
 sg13g2_decap_4 FILLER_40_2353 ();
 sg13g2_fill_1 FILLER_40_2357 ();
 sg13g2_decap_8 FILLER_40_2375 ();
 sg13g2_decap_8 FILLER_40_2382 ();
 sg13g2_decap_8 FILLER_40_2389 ();
 sg13g2_fill_2 FILLER_40_2396 ();
 sg13g2_fill_1 FILLER_40_2398 ();
 sg13g2_fill_2 FILLER_40_2404 ();
 sg13g2_fill_1 FILLER_40_2406 ();
 sg13g2_fill_1 FILLER_40_2412 ();
 sg13g2_decap_4 FILLER_40_2421 ();
 sg13g2_fill_1 FILLER_40_2425 ();
 sg13g2_fill_2 FILLER_40_2443 ();
 sg13g2_fill_1 FILLER_40_2445 ();
 sg13g2_decap_8 FILLER_40_2451 ();
 sg13g2_decap_8 FILLER_40_2458 ();
 sg13g2_decap_4 FILLER_40_2465 ();
 sg13g2_fill_1 FILLER_40_2469 ();
 sg13g2_decap_4 FILLER_40_2492 ();
 sg13g2_fill_1 FILLER_40_2496 ();
 sg13g2_fill_2 FILLER_40_2502 ();
 sg13g2_decap_4 FILLER_40_2514 ();
 sg13g2_fill_2 FILLER_40_2518 ();
 sg13g2_fill_2 FILLER_40_2525 ();
 sg13g2_fill_1 FILLER_40_2527 ();
 sg13g2_fill_1 FILLER_40_2538 ();
 sg13g2_fill_1 FILLER_40_2544 ();
 sg13g2_decap_8 FILLER_40_2549 ();
 sg13g2_fill_1 FILLER_40_2556 ();
 sg13g2_fill_2 FILLER_40_2572 ();
 sg13g2_decap_4 FILLER_40_2582 ();
 sg13g2_decap_4 FILLER_40_2607 ();
 sg13g2_fill_1 FILLER_40_2615 ();
 sg13g2_fill_2 FILLER_40_2622 ();
 sg13g2_decap_8 FILLER_40_2660 ();
 sg13g2_fill_2 FILLER_40_2667 ();
 sg13g2_fill_1 FILLER_40_2669 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_27 ();
 sg13g2_fill_2 FILLER_41_37 ();
 sg13g2_fill_1 FILLER_41_86 ();
 sg13g2_decap_4 FILLER_41_96 ();
 sg13g2_fill_2 FILLER_41_108 ();
 sg13g2_fill_1 FILLER_41_110 ();
 sg13g2_fill_2 FILLER_41_132 ();
 sg13g2_fill_2 FILLER_41_188 ();
 sg13g2_fill_2 FILLER_41_212 ();
 sg13g2_fill_1 FILLER_41_237 ();
 sg13g2_fill_1 FILLER_41_246 ();
 sg13g2_decap_4 FILLER_41_314 ();
 sg13g2_fill_1 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_362 ();
 sg13g2_fill_2 FILLER_41_394 ();
 sg13g2_fill_2 FILLER_41_417 ();
 sg13g2_fill_1 FILLER_41_419 ();
 sg13g2_fill_1 FILLER_41_434 ();
 sg13g2_fill_1 FILLER_41_440 ();
 sg13g2_fill_2 FILLER_41_462 ();
 sg13g2_fill_1 FILLER_41_464 ();
 sg13g2_fill_2 FILLER_41_469 ();
 sg13g2_fill_1 FILLER_41_471 ();
 sg13g2_fill_2 FILLER_41_493 ();
 sg13g2_fill_2 FILLER_41_523 ();
 sg13g2_fill_2 FILLER_41_545 ();
 sg13g2_fill_2 FILLER_41_551 ();
 sg13g2_fill_2 FILLER_41_571 ();
 sg13g2_fill_2 FILLER_41_584 ();
 sg13g2_fill_1 FILLER_41_606 ();
 sg13g2_fill_1 FILLER_41_611 ();
 sg13g2_decap_8 FILLER_41_669 ();
 sg13g2_fill_1 FILLER_41_676 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_4 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_799 ();
 sg13g2_decap_8 FILLER_41_806 ();
 sg13g2_decap_8 FILLER_41_813 ();
 sg13g2_decap_4 FILLER_41_820 ();
 sg13g2_fill_1 FILLER_41_858 ();
 sg13g2_fill_2 FILLER_41_914 ();
 sg13g2_decap_8 FILLER_41_942 ();
 sg13g2_fill_2 FILLER_41_949 ();
 sg13g2_fill_2 FILLER_41_983 ();
 sg13g2_fill_1 FILLER_41_985 ();
 sg13g2_fill_2 FILLER_41_994 ();
 sg13g2_fill_2 FILLER_41_1010 ();
 sg13g2_fill_2 FILLER_41_1038 ();
 sg13g2_fill_2 FILLER_41_1070 ();
 sg13g2_fill_2 FILLER_41_1077 ();
 sg13g2_fill_1 FILLER_41_1090 ();
 sg13g2_fill_2 FILLER_41_1104 ();
 sg13g2_fill_1 FILLER_41_1162 ();
 sg13g2_fill_2 FILLER_41_1206 ();
 sg13g2_fill_1 FILLER_41_1244 ();
 sg13g2_fill_1 FILLER_41_1266 ();
 sg13g2_fill_2 FILLER_41_1289 ();
 sg13g2_fill_1 FILLER_41_1291 ();
 sg13g2_fill_2 FILLER_41_1308 ();
 sg13g2_fill_2 FILLER_41_1325 ();
 sg13g2_fill_2 FILLER_41_1358 ();
 sg13g2_fill_2 FILLER_41_1364 ();
 sg13g2_fill_2 FILLER_41_1397 ();
 sg13g2_fill_1 FILLER_41_1429 ();
 sg13g2_fill_2 FILLER_41_1438 ();
 sg13g2_fill_2 FILLER_41_1447 ();
 sg13g2_fill_1 FILLER_41_1454 ();
 sg13g2_decap_4 FILLER_41_1460 ();
 sg13g2_fill_1 FILLER_41_1468 ();
 sg13g2_fill_2 FILLER_41_1473 ();
 sg13g2_decap_4 FILLER_41_1484 ();
 sg13g2_fill_2 FILLER_41_1488 ();
 sg13g2_decap_8 FILLER_41_1499 ();
 sg13g2_fill_1 FILLER_41_1532 ();
 sg13g2_decap_4 FILLER_41_1542 ();
 sg13g2_fill_1 FILLER_41_1558 ();
 sg13g2_fill_1 FILLER_41_1567 ();
 sg13g2_fill_2 FILLER_41_1600 ();
 sg13g2_fill_1 FILLER_41_1619 ();
 sg13g2_fill_2 FILLER_41_1625 ();
 sg13g2_fill_1 FILLER_41_1638 ();
 sg13g2_fill_1 FILLER_41_1642 ();
 sg13g2_fill_2 FILLER_41_1651 ();
 sg13g2_fill_1 FILLER_41_1700 ();
 sg13g2_fill_2 FILLER_41_1734 ();
 sg13g2_fill_1 FILLER_41_1736 ();
 sg13g2_fill_1 FILLER_41_1773 ();
 sg13g2_fill_1 FILLER_41_1779 ();
 sg13g2_fill_2 FILLER_41_1786 ();
 sg13g2_fill_1 FILLER_41_1866 ();
 sg13g2_fill_1 FILLER_41_1871 ();
 sg13g2_fill_1 FILLER_41_1903 ();
 sg13g2_fill_1 FILLER_41_1922 ();
 sg13g2_fill_1 FILLER_41_1930 ();
 sg13g2_fill_1 FILLER_41_1976 ();
 sg13g2_fill_2 FILLER_41_1984 ();
 sg13g2_fill_1 FILLER_41_2000 ();
 sg13g2_fill_1 FILLER_41_2010 ();
 sg13g2_fill_2 FILLER_41_2049 ();
 sg13g2_decap_4 FILLER_41_2077 ();
 sg13g2_fill_2 FILLER_41_2081 ();
 sg13g2_decap_8 FILLER_41_2087 ();
 sg13g2_decap_8 FILLER_41_2094 ();
 sg13g2_decap_8 FILLER_41_2101 ();
 sg13g2_decap_8 FILLER_41_2108 ();
 sg13g2_decap_4 FILLER_41_2115 ();
 sg13g2_fill_1 FILLER_41_2119 ();
 sg13g2_decap_8 FILLER_41_2128 ();
 sg13g2_decap_8 FILLER_41_2135 ();
 sg13g2_decap_8 FILLER_41_2142 ();
 sg13g2_decap_4 FILLER_41_2149 ();
 sg13g2_fill_1 FILLER_41_2176 ();
 sg13g2_fill_1 FILLER_41_2182 ();
 sg13g2_fill_2 FILLER_41_2187 ();
 sg13g2_decap_8 FILLER_41_2195 ();
 sg13g2_decap_4 FILLER_41_2202 ();
 sg13g2_fill_2 FILLER_41_2210 ();
 sg13g2_fill_1 FILLER_41_2212 ();
 sg13g2_fill_1 FILLER_41_2250 ();
 sg13g2_fill_2 FILLER_41_2255 ();
 sg13g2_fill_1 FILLER_41_2257 ();
 sg13g2_fill_2 FILLER_41_2280 ();
 sg13g2_fill_1 FILLER_41_2282 ();
 sg13g2_fill_2 FILLER_41_2307 ();
 sg13g2_fill_1 FILLER_41_2309 ();
 sg13g2_decap_4 FILLER_41_2323 ();
 sg13g2_fill_2 FILLER_41_2327 ();
 sg13g2_decap_4 FILLER_41_2334 ();
 sg13g2_fill_2 FILLER_41_2338 ();
 sg13g2_decap_4 FILLER_41_2344 ();
 sg13g2_fill_1 FILLER_41_2352 ();
 sg13g2_fill_2 FILLER_41_2357 ();
 sg13g2_fill_2 FILLER_41_2365 ();
 sg13g2_fill_2 FILLER_41_2371 ();
 sg13g2_fill_1 FILLER_41_2373 ();
 sg13g2_decap_8 FILLER_41_2378 ();
 sg13g2_decap_4 FILLER_41_2385 ();
 sg13g2_fill_1 FILLER_41_2389 ();
 sg13g2_fill_2 FILLER_41_2395 ();
 sg13g2_fill_1 FILLER_41_2397 ();
 sg13g2_decap_4 FILLER_41_2403 ();
 sg13g2_fill_2 FILLER_41_2407 ();
 sg13g2_fill_2 FILLER_41_2413 ();
 sg13g2_fill_1 FILLER_41_2415 ();
 sg13g2_fill_1 FILLER_41_2421 ();
 sg13g2_decap_8 FILLER_41_2459 ();
 sg13g2_decap_8 FILLER_41_2466 ();
 sg13g2_fill_2 FILLER_41_2473 ();
 sg13g2_decap_8 FILLER_41_2480 ();
 sg13g2_decap_8 FILLER_41_2487 ();
 sg13g2_fill_1 FILLER_41_2494 ();
 sg13g2_decap_8 FILLER_41_2500 ();
 sg13g2_decap_8 FILLER_41_2507 ();
 sg13g2_decap_4 FILLER_41_2514 ();
 sg13g2_fill_1 FILLER_41_2560 ();
 sg13g2_fill_2 FILLER_41_2600 ();
 sg13g2_fill_1 FILLER_41_2613 ();
 sg13g2_fill_2 FILLER_41_2625 ();
 sg13g2_fill_1 FILLER_41_2627 ();
 sg13g2_decap_8 FILLER_41_2633 ();
 sg13g2_fill_2 FILLER_41_2640 ();
 sg13g2_decap_8 FILLER_41_2646 ();
 sg13g2_decap_8 FILLER_41_2653 ();
 sg13g2_decap_8 FILLER_41_2660 ();
 sg13g2_fill_2 FILLER_41_2667 ();
 sg13g2_fill_1 FILLER_41_2669 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_2 ();
 sg13g2_fill_1 FILLER_42_40 ();
 sg13g2_fill_1 FILLER_42_99 ();
 sg13g2_fill_1 FILLER_42_104 ();
 sg13g2_decap_4 FILLER_42_109 ();
 sg13g2_fill_2 FILLER_42_118 ();
 sg13g2_decap_8 FILLER_42_129 ();
 sg13g2_fill_2 FILLER_42_136 ();
 sg13g2_fill_2 FILLER_42_142 ();
 sg13g2_fill_1 FILLER_42_144 ();
 sg13g2_fill_2 FILLER_42_176 ();
 sg13g2_fill_2 FILLER_42_198 ();
 sg13g2_fill_2 FILLER_42_241 ();
 sg13g2_fill_2 FILLER_42_289 ();
 sg13g2_fill_1 FILLER_42_296 ();
 sg13g2_fill_2 FILLER_42_354 ();
 sg13g2_decap_4 FILLER_42_477 ();
 sg13g2_fill_1 FILLER_42_481 ();
 sg13g2_fill_1 FILLER_42_485 ();
 sg13g2_fill_1 FILLER_42_504 ();
 sg13g2_fill_1 FILLER_42_516 ();
 sg13g2_fill_1 FILLER_42_550 ();
 sg13g2_fill_1 FILLER_42_573 ();
 sg13g2_fill_2 FILLER_42_581 ();
 sg13g2_fill_2 FILLER_42_604 ();
 sg13g2_fill_1 FILLER_42_606 ();
 sg13g2_fill_2 FILLER_42_621 ();
 sg13g2_fill_1 FILLER_42_623 ();
 sg13g2_fill_2 FILLER_42_628 ();
 sg13g2_decap_4 FILLER_42_634 ();
 sg13g2_fill_1 FILLER_42_642 ();
 sg13g2_fill_2 FILLER_42_651 ();
 sg13g2_fill_1 FILLER_42_662 ();
 sg13g2_fill_1 FILLER_42_667 ();
 sg13g2_fill_1 FILLER_42_687 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_fill_1 FILLER_42_730 ();
 sg13g2_fill_1 FILLER_42_768 ();
 sg13g2_decap_4 FILLER_42_816 ();
 sg13g2_fill_1 FILLER_42_868 ();
 sg13g2_decap_4 FILLER_42_873 ();
 sg13g2_decap_8 FILLER_42_882 ();
 sg13g2_fill_1 FILLER_42_889 ();
 sg13g2_fill_2 FILLER_42_898 ();
 sg13g2_fill_1 FILLER_42_900 ();
 sg13g2_fill_1 FILLER_42_913 ();
 sg13g2_fill_1 FILLER_42_940 ();
 sg13g2_fill_1 FILLER_42_972 ();
 sg13g2_fill_2 FILLER_42_1048 ();
 sg13g2_fill_1 FILLER_42_1084 ();
 sg13g2_fill_2 FILLER_42_1135 ();
 sg13g2_fill_1 FILLER_42_1161 ();
 sg13g2_fill_2 FILLER_42_1169 ();
 sg13g2_fill_2 FILLER_42_1174 ();
 sg13g2_fill_2 FILLER_42_1188 ();
 sg13g2_fill_2 FILLER_42_1194 ();
 sg13g2_fill_2 FILLER_42_1231 ();
 sg13g2_fill_1 FILLER_42_1242 ();
 sg13g2_decap_4 FILLER_42_1260 ();
 sg13g2_fill_2 FILLER_42_1264 ();
 sg13g2_fill_2 FILLER_42_1297 ();
 sg13g2_fill_1 FILLER_42_1367 ();
 sg13g2_fill_1 FILLER_42_1376 ();
 sg13g2_fill_2 FILLER_42_1385 ();
 sg13g2_fill_2 FILLER_42_1396 ();
 sg13g2_fill_1 FILLER_42_1413 ();
 sg13g2_fill_1 FILLER_42_1418 ();
 sg13g2_fill_1 FILLER_42_1424 ();
 sg13g2_decap_8 FILLER_42_1553 ();
 sg13g2_fill_1 FILLER_42_1560 ();
 sg13g2_fill_1 FILLER_42_1566 ();
 sg13g2_fill_2 FILLER_42_1576 ();
 sg13g2_fill_1 FILLER_42_1578 ();
 sg13g2_fill_2 FILLER_42_1634 ();
 sg13g2_fill_1 FILLER_42_1655 ();
 sg13g2_decap_4 FILLER_42_1673 ();
 sg13g2_fill_2 FILLER_42_1677 ();
 sg13g2_fill_2 FILLER_42_1687 ();
 sg13g2_fill_2 FILLER_42_1693 ();
 sg13g2_fill_1 FILLER_42_1695 ();
 sg13g2_fill_2 FILLER_42_1700 ();
 sg13g2_fill_1 FILLER_42_1702 ();
 sg13g2_fill_1 FILLER_42_1711 ();
 sg13g2_decap_4 FILLER_42_1721 ();
 sg13g2_fill_1 FILLER_42_1751 ();
 sg13g2_fill_1 FILLER_42_1755 ();
 sg13g2_fill_1 FILLER_42_1773 ();
 sg13g2_fill_2 FILLER_42_1778 ();
 sg13g2_fill_2 FILLER_42_1809 ();
 sg13g2_fill_2 FILLER_42_1824 ();
 sg13g2_fill_2 FILLER_42_1833 ();
 sg13g2_fill_1 FILLER_42_1849 ();
 sg13g2_fill_1 FILLER_42_1876 ();
 sg13g2_fill_1 FILLER_42_1888 ();
 sg13g2_decap_8 FILLER_42_1894 ();
 sg13g2_fill_1 FILLER_42_1933 ();
 sg13g2_fill_2 FILLER_42_1947 ();
 sg13g2_fill_2 FILLER_42_1989 ();
 sg13g2_fill_1 FILLER_42_1996 ();
 sg13g2_fill_1 FILLER_42_2010 ();
 sg13g2_fill_1 FILLER_42_2015 ();
 sg13g2_fill_1 FILLER_42_2021 ();
 sg13g2_fill_1 FILLER_42_2027 ();
 sg13g2_fill_2 FILLER_42_2032 ();
 sg13g2_decap_8 FILLER_42_2038 ();
 sg13g2_fill_2 FILLER_42_2045 ();
 sg13g2_decap_4 FILLER_42_2098 ();
 sg13g2_fill_1 FILLER_42_2102 ();
 sg13g2_decap_8 FILLER_42_2139 ();
 sg13g2_decap_4 FILLER_42_2146 ();
 sg13g2_fill_2 FILLER_42_2165 ();
 sg13g2_fill_1 FILLER_42_2167 ();
 sg13g2_fill_2 FILLER_42_2177 ();
 sg13g2_fill_1 FILLER_42_2179 ();
 sg13g2_decap_8 FILLER_42_2195 ();
 sg13g2_decap_4 FILLER_42_2202 ();
 sg13g2_fill_2 FILLER_42_2206 ();
 sg13g2_decap_8 FILLER_42_2212 ();
 sg13g2_decap_4 FILLER_42_2219 ();
 sg13g2_fill_2 FILLER_42_2255 ();
 sg13g2_fill_2 FILLER_42_2265 ();
 sg13g2_decap_4 FILLER_42_2272 ();
 sg13g2_fill_2 FILLER_42_2282 ();
 sg13g2_decap_4 FILLER_42_2290 ();
 sg13g2_fill_2 FILLER_42_2304 ();
 sg13g2_decap_4 FILLER_42_2321 ();
 sg13g2_decap_4 FILLER_42_2347 ();
 sg13g2_fill_1 FILLER_42_2351 ();
 sg13g2_decap_4 FILLER_42_2373 ();
 sg13g2_fill_2 FILLER_42_2377 ();
 sg13g2_decap_8 FILLER_42_2395 ();
 sg13g2_fill_2 FILLER_42_2402 ();
 sg13g2_decap_8 FILLER_42_2437 ();
 sg13g2_fill_1 FILLER_42_2444 ();
 sg13g2_fill_1 FILLER_42_2471 ();
 sg13g2_decap_8 FILLER_42_2485 ();
 sg13g2_decap_8 FILLER_42_2501 ();
 sg13g2_fill_2 FILLER_42_2508 ();
 sg13g2_fill_1 FILLER_42_2553 ();
 sg13g2_decap_4 FILLER_42_2561 ();
 sg13g2_decap_4 FILLER_42_2611 ();
 sg13g2_fill_2 FILLER_42_2615 ();
 sg13g2_decap_8 FILLER_42_2629 ();
 sg13g2_fill_2 FILLER_42_2636 ();
 sg13g2_decap_8 FILLER_42_2663 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_33 ();
 sg13g2_fill_1 FILLER_43_65 ();
 sg13g2_fill_2 FILLER_43_76 ();
 sg13g2_fill_2 FILLER_43_82 ();
 sg13g2_fill_1 FILLER_43_84 ();
 sg13g2_fill_1 FILLER_43_177 ();
 sg13g2_fill_1 FILLER_43_183 ();
 sg13g2_fill_1 FILLER_43_216 ();
 sg13g2_fill_1 FILLER_43_252 ();
 sg13g2_fill_1 FILLER_43_281 ();
 sg13g2_fill_1 FILLER_43_295 ();
 sg13g2_fill_1 FILLER_43_300 ();
 sg13g2_fill_1 FILLER_43_305 ();
 sg13g2_fill_1 FILLER_43_310 ();
 sg13g2_fill_1 FILLER_43_316 ();
 sg13g2_fill_1 FILLER_43_322 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_fill_1 FILLER_43_332 ();
 sg13g2_fill_1 FILLER_43_367 ();
 sg13g2_decap_8 FILLER_43_397 ();
 sg13g2_fill_1 FILLER_43_404 ();
 sg13g2_fill_2 FILLER_43_445 ();
 sg13g2_fill_1 FILLER_43_447 ();
 sg13g2_fill_1 FILLER_43_484 ();
 sg13g2_fill_1 FILLER_43_489 ();
 sg13g2_fill_1 FILLER_43_494 ();
 sg13g2_fill_2 FILLER_43_515 ();
 sg13g2_fill_2 FILLER_43_581 ();
 sg13g2_fill_1 FILLER_43_586 ();
 sg13g2_decap_8 FILLER_43_600 ();
 sg13g2_decap_8 FILLER_43_607 ();
 sg13g2_decap_8 FILLER_43_614 ();
 sg13g2_decap_4 FILLER_43_625 ();
 sg13g2_decap_4 FILLER_43_642 ();
 sg13g2_fill_1 FILLER_43_646 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_fill_2 FILLER_43_665 ();
 sg13g2_fill_2 FILLER_43_672 ();
 sg13g2_decap_4 FILLER_43_688 ();
 sg13g2_fill_1 FILLER_43_692 ();
 sg13g2_fill_1 FILLER_43_723 ();
 sg13g2_fill_2 FILLER_43_733 ();
 sg13g2_fill_2 FILLER_43_765 ();
 sg13g2_fill_2 FILLER_43_778 ();
 sg13g2_fill_1 FILLER_43_792 ();
 sg13g2_fill_2 FILLER_43_827 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_fill_2 FILLER_43_875 ();
 sg13g2_decap_4 FILLER_43_889 ();
 sg13g2_fill_2 FILLER_43_893 ();
 sg13g2_decap_8 FILLER_43_899 ();
 sg13g2_fill_1 FILLER_43_906 ();
 sg13g2_decap_4 FILLER_43_932 ();
 sg13g2_fill_1 FILLER_43_976 ();
 sg13g2_fill_1 FILLER_43_982 ();
 sg13g2_fill_1 FILLER_43_988 ();
 sg13g2_fill_1 FILLER_43_1015 ();
 sg13g2_fill_2 FILLER_43_1046 ();
 sg13g2_fill_2 FILLER_43_1068 ();
 sg13g2_fill_1 FILLER_43_1097 ();
 sg13g2_fill_1 FILLER_43_1130 ();
 sg13g2_fill_1 FILLER_43_1155 ();
 sg13g2_fill_1 FILLER_43_1221 ();
 sg13g2_fill_1 FILLER_43_1236 ();
 sg13g2_fill_1 FILLER_43_1255 ();
 sg13g2_decap_4 FILLER_43_1287 ();
 sg13g2_fill_1 FILLER_43_1291 ();
 sg13g2_decap_4 FILLER_43_1332 ();
 sg13g2_fill_1 FILLER_43_1336 ();
 sg13g2_fill_1 FILLER_43_1341 ();
 sg13g2_fill_2 FILLER_43_1389 ();
 sg13g2_fill_1 FILLER_43_1401 ();
 sg13g2_fill_1 FILLER_43_1439 ();
 sg13g2_fill_1 FILLER_43_1447 ();
 sg13g2_fill_1 FILLER_43_1458 ();
 sg13g2_decap_4 FILLER_43_1481 ();
 sg13g2_fill_2 FILLER_43_1485 ();
 sg13g2_decap_8 FILLER_43_1495 ();
 sg13g2_fill_2 FILLER_43_1502 ();
 sg13g2_decap_8 FILLER_43_1509 ();
 sg13g2_decap_4 FILLER_43_1520 ();
 sg13g2_fill_1 FILLER_43_1524 ();
 sg13g2_fill_1 FILLER_43_1556 ();
 sg13g2_fill_2 FILLER_43_1588 ();
 sg13g2_decap_4 FILLER_43_1594 ();
 sg13g2_fill_1 FILLER_43_1598 ();
 sg13g2_fill_1 FILLER_43_1623 ();
 sg13g2_fill_1 FILLER_43_1650 ();
 sg13g2_fill_1 FILLER_43_1664 ();
 sg13g2_fill_2 FILLER_43_1688 ();
 sg13g2_decap_8 FILLER_43_1725 ();
 sg13g2_fill_2 FILLER_43_1732 ();
 sg13g2_fill_1 FILLER_43_1742 ();
 sg13g2_fill_2 FILLER_43_1760 ();
 sg13g2_fill_2 FILLER_43_1795 ();
 sg13g2_fill_2 FILLER_43_1856 ();
 sg13g2_fill_2 FILLER_43_1882 ();
 sg13g2_fill_1 FILLER_43_1884 ();
 sg13g2_decap_4 FILLER_43_1919 ();
 sg13g2_fill_2 FILLER_43_1923 ();
 sg13g2_fill_1 FILLER_43_1946 ();
 sg13g2_fill_1 FILLER_43_1950 ();
 sg13g2_fill_2 FILLER_43_1954 ();
 sg13g2_decap_8 FILLER_43_1960 ();
 sg13g2_decap_4 FILLER_43_1967 ();
 sg13g2_fill_2 FILLER_43_1971 ();
 sg13g2_fill_2 FILLER_43_1977 ();
 sg13g2_fill_1 FILLER_43_1979 ();
 sg13g2_decap_8 FILLER_43_2043 ();
 sg13g2_decap_4 FILLER_43_2050 ();
 sg13g2_decap_8 FILLER_43_2096 ();
 sg13g2_fill_1 FILLER_43_2103 ();
 sg13g2_decap_8 FILLER_43_2130 ();
 sg13g2_decap_8 FILLER_43_2137 ();
 sg13g2_decap_4 FILLER_43_2144 ();
 sg13g2_fill_2 FILLER_43_2148 ();
 sg13g2_fill_2 FILLER_43_2154 ();
 sg13g2_fill_1 FILLER_43_2160 ();
 sg13g2_fill_1 FILLER_43_2169 ();
 sg13g2_fill_1 FILLER_43_2175 ();
 sg13g2_decap_8 FILLER_43_2202 ();
 sg13g2_fill_1 FILLER_43_2209 ();
 sg13g2_decap_8 FILLER_43_2214 ();
 sg13g2_fill_1 FILLER_43_2221 ();
 sg13g2_fill_1 FILLER_43_2230 ();
 sg13g2_fill_1 FILLER_43_2236 ();
 sg13g2_fill_1 FILLER_43_2252 ();
 sg13g2_decap_8 FILLER_43_2257 ();
 sg13g2_fill_2 FILLER_43_2264 ();
 sg13g2_decap_8 FILLER_43_2305 ();
 sg13g2_decap_4 FILLER_43_2312 ();
 sg13g2_fill_1 FILLER_43_2322 ();
 sg13g2_decap_8 FILLER_43_2327 ();
 sg13g2_fill_2 FILLER_43_2334 ();
 sg13g2_fill_1 FILLER_43_2336 ();
 sg13g2_fill_2 FILLER_43_2398 ();
 sg13g2_fill_1 FILLER_43_2400 ();
 sg13g2_fill_2 FILLER_43_2412 ();
 sg13g2_decap_8 FILLER_43_2419 ();
 sg13g2_decap_4 FILLER_43_2426 ();
 sg13g2_fill_2 FILLER_43_2438 ();
 sg13g2_fill_1 FILLER_43_2440 ();
 sg13g2_fill_1 FILLER_43_2449 ();
 sg13g2_fill_1 FILLER_43_2456 ();
 sg13g2_fill_2 FILLER_43_2463 ();
 sg13g2_decap_8 FILLER_43_2500 ();
 sg13g2_decap_8 FILLER_43_2507 ();
 sg13g2_decap_4 FILLER_43_2514 ();
 sg13g2_fill_1 FILLER_43_2548 ();
 sg13g2_fill_2 FILLER_43_2600 ();
 sg13g2_decap_4 FILLER_43_2607 ();
 sg13g2_decap_4 FILLER_43_2664 ();
 sg13g2_fill_2 FILLER_43_2668 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_decap_4 FILLER_44_32 ();
 sg13g2_fill_2 FILLER_44_36 ();
 sg13g2_fill_2 FILLER_44_47 ();
 sg13g2_fill_1 FILLER_44_49 ();
 sg13g2_fill_1 FILLER_44_54 ();
 sg13g2_decap_4 FILLER_44_80 ();
 sg13g2_decap_4 FILLER_44_88 ();
 sg13g2_decap_8 FILLER_44_96 ();
 sg13g2_fill_2 FILLER_44_107 ();
 sg13g2_decap_8 FILLER_44_143 ();
 sg13g2_fill_2 FILLER_44_150 ();
 sg13g2_fill_1 FILLER_44_152 ();
 sg13g2_decap_8 FILLER_44_157 ();
 sg13g2_fill_2 FILLER_44_202 ();
 sg13g2_fill_1 FILLER_44_208 ();
 sg13g2_decap_4 FILLER_44_282 ();
 sg13g2_fill_1 FILLER_44_286 ();
 sg13g2_decap_8 FILLER_44_291 ();
 sg13g2_decap_8 FILLER_44_298 ();
 sg13g2_decap_8 FILLER_44_305 ();
 sg13g2_fill_2 FILLER_44_312 ();
 sg13g2_decap_4 FILLER_44_318 ();
 sg13g2_fill_1 FILLER_44_322 ();
 sg13g2_fill_2 FILLER_44_331 ();
 sg13g2_fill_1 FILLER_44_333 ();
 sg13g2_fill_1 FILLER_44_338 ();
 sg13g2_fill_2 FILLER_44_366 ();
 sg13g2_fill_1 FILLER_44_378 ();
 sg13g2_fill_1 FILLER_44_383 ();
 sg13g2_fill_1 FILLER_44_398 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_fill_1 FILLER_44_459 ();
 sg13g2_fill_2 FILLER_44_481 ();
 sg13g2_fill_1 FILLER_44_483 ();
 sg13g2_fill_2 FILLER_44_489 ();
 sg13g2_fill_2 FILLER_44_526 ();
 sg13g2_fill_1 FILLER_44_528 ();
 sg13g2_fill_2 FILLER_44_534 ();
 sg13g2_fill_1 FILLER_44_536 ();
 sg13g2_fill_2 FILLER_44_580 ();
 sg13g2_fill_1 FILLER_44_586 ();
 sg13g2_decap_8 FILLER_44_596 ();
 sg13g2_fill_1 FILLER_44_626 ();
 sg13g2_fill_1 FILLER_44_631 ();
 sg13g2_fill_1 FILLER_44_658 ();
 sg13g2_fill_2 FILLER_44_663 ();
 sg13g2_fill_2 FILLER_44_673 ();
 sg13g2_decap_8 FILLER_44_691 ();
 sg13g2_decap_8 FILLER_44_698 ();
 sg13g2_decap_8 FILLER_44_705 ();
 sg13g2_fill_1 FILLER_44_712 ();
 sg13g2_fill_2 FILLER_44_717 ();
 sg13g2_fill_2 FILLER_44_740 ();
 sg13g2_fill_1 FILLER_44_755 ();
 sg13g2_fill_1 FILLER_44_764 ();
 sg13g2_fill_1 FILLER_44_769 ();
 sg13g2_fill_1 FILLER_44_775 ();
 sg13g2_fill_1 FILLER_44_797 ();
 sg13g2_fill_1 FILLER_44_803 ();
 sg13g2_fill_2 FILLER_44_830 ();
 sg13g2_decap_4 FILLER_44_865 ();
 sg13g2_fill_2 FILLER_44_869 ();
 sg13g2_decap_8 FILLER_44_906 ();
 sg13g2_decap_8 FILLER_44_913 ();
 sg13g2_decap_8 FILLER_44_920 ();
 sg13g2_fill_1 FILLER_44_927 ();
 sg13g2_fill_2 FILLER_44_951 ();
 sg13g2_fill_2 FILLER_44_1000 ();
 sg13g2_fill_1 FILLER_44_1005 ();
 sg13g2_fill_1 FILLER_44_1026 ();
 sg13g2_fill_1 FILLER_44_1047 ();
 sg13g2_fill_1 FILLER_44_1053 ();
 sg13g2_fill_1 FILLER_44_1059 ();
 sg13g2_fill_1 FILLER_44_1089 ();
 sg13g2_fill_1 FILLER_44_1100 ();
 sg13g2_fill_2 FILLER_44_1139 ();
 sg13g2_fill_1 FILLER_44_1187 ();
 sg13g2_fill_2 FILLER_44_1212 ();
 sg13g2_fill_1 FILLER_44_1261 ();
 sg13g2_decap_8 FILLER_44_1297 ();
 sg13g2_fill_1 FILLER_44_1304 ();
 sg13g2_fill_2 FILLER_44_1313 ();
 sg13g2_fill_2 FILLER_44_1330 ();
 sg13g2_fill_1 FILLER_44_1365 ();
 sg13g2_fill_1 FILLER_44_1377 ();
 sg13g2_fill_1 FILLER_44_1399 ();
 sg13g2_fill_1 FILLER_44_1447 ();
 sg13g2_fill_2 FILLER_44_1460 ();
 sg13g2_decap_8 FILLER_44_1488 ();
 sg13g2_decap_8 FILLER_44_1495 ();
 sg13g2_decap_8 FILLER_44_1502 ();
 sg13g2_fill_2 FILLER_44_1509 ();
 sg13g2_fill_1 FILLER_44_1524 ();
 sg13g2_fill_2 FILLER_44_1567 ();
 sg13g2_decap_4 FILLER_44_1599 ();
 sg13g2_fill_1 FILLER_44_1603 ();
 sg13g2_decap_8 FILLER_44_1609 ();
 sg13g2_decap_4 FILLER_44_1616 ();
 sg13g2_fill_1 FILLER_44_1658 ();
 sg13g2_fill_2 FILLER_44_1745 ();
 sg13g2_fill_1 FILLER_44_1751 ();
 sg13g2_fill_1 FILLER_44_1759 ();
 sg13g2_fill_2 FILLER_44_1779 ();
 sg13g2_fill_1 FILLER_44_1807 ();
 sg13g2_fill_2 FILLER_44_1821 ();
 sg13g2_fill_1 FILLER_44_1828 ();
 sg13g2_fill_2 FILLER_44_1833 ();
 sg13g2_fill_2 FILLER_44_1840 ();
 sg13g2_fill_2 FILLER_44_1846 ();
 sg13g2_fill_1 FILLER_44_1873 ();
 sg13g2_decap_4 FILLER_44_1954 ();
 sg13g2_fill_2 FILLER_44_1958 ();
 sg13g2_fill_2 FILLER_44_1964 ();
 sg13g2_fill_2 FILLER_44_1970 ();
 sg13g2_decap_4 FILLER_44_1977 ();
 sg13g2_fill_2 FILLER_44_1981 ();
 sg13g2_decap_4 FILLER_44_2030 ();
 sg13g2_decap_4 FILLER_44_2055 ();
 sg13g2_fill_2 FILLER_44_2059 ();
 sg13g2_decap_4 FILLER_44_2087 ();
 sg13g2_fill_1 FILLER_44_2091 ();
 sg13g2_fill_2 FILLER_44_2102 ();
 sg13g2_fill_1 FILLER_44_2104 ();
 sg13g2_decap_4 FILLER_44_2135 ();
 sg13g2_fill_2 FILLER_44_2139 ();
 sg13g2_decap_8 FILLER_44_2145 ();
 sg13g2_fill_2 FILLER_44_2152 ();
 sg13g2_fill_1 FILLER_44_2199 ();
 sg13g2_decap_8 FILLER_44_2215 ();
 sg13g2_fill_1 FILLER_44_2230 ();
 sg13g2_fill_2 FILLER_44_2266 ();
 sg13g2_fill_1 FILLER_44_2268 ();
 sg13g2_decap_4 FILLER_44_2273 ();
 sg13g2_fill_1 FILLER_44_2277 ();
 sg13g2_decap_8 FILLER_44_2283 ();
 sg13g2_decap_8 FILLER_44_2290 ();
 sg13g2_decap_8 FILLER_44_2297 ();
 sg13g2_fill_1 FILLER_44_2304 ();
 sg13g2_decap_8 FILLER_44_2309 ();
 sg13g2_decap_4 FILLER_44_2316 ();
 sg13g2_fill_1 FILLER_44_2320 ();
 sg13g2_fill_1 FILLER_44_2357 ();
 sg13g2_fill_2 FILLER_44_2364 ();
 sg13g2_decap_8 FILLER_44_2371 ();
 sg13g2_fill_2 FILLER_44_2378 ();
 sg13g2_fill_1 FILLER_44_2380 ();
 sg13g2_decap_8 FILLER_44_2393 ();
 sg13g2_decap_8 FILLER_44_2400 ();
 sg13g2_fill_2 FILLER_44_2411 ();
 sg13g2_fill_1 FILLER_44_2424 ();
 sg13g2_decap_4 FILLER_44_2435 ();
 sg13g2_fill_2 FILLER_44_2439 ();
 sg13g2_fill_2 FILLER_44_2445 ();
 sg13g2_decap_4 FILLER_44_2451 ();
 sg13g2_fill_2 FILLER_44_2455 ();
 sg13g2_decap_8 FILLER_44_2462 ();
 sg13g2_decap_4 FILLER_44_2469 ();
 sg13g2_fill_2 FILLER_44_2473 ();
 sg13g2_decap_8 FILLER_44_2486 ();
 sg13g2_fill_1 FILLER_44_2493 ();
 sg13g2_decap_8 FILLER_44_2532 ();
 sg13g2_fill_1 FILLER_44_2539 ();
 sg13g2_decap_4 FILLER_44_2545 ();
 sg13g2_fill_1 FILLER_44_2549 ();
 sg13g2_decap_4 FILLER_44_2555 ();
 sg13g2_fill_1 FILLER_44_2559 ();
 sg13g2_decap_8 FILLER_44_2586 ();
 sg13g2_decap_4 FILLER_44_2593 ();
 sg13g2_fill_2 FILLER_44_2597 ();
 sg13g2_fill_1 FILLER_44_2634 ();
 sg13g2_decap_8 FILLER_44_2656 ();
 sg13g2_decap_8 FILLER_44_2663 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_15 ();
 sg13g2_fill_2 FILLER_45_22 ();
 sg13g2_fill_1 FILLER_45_24 ();
 sg13g2_decap_8 FILLER_45_34 ();
 sg13g2_decap_4 FILLER_45_41 ();
 sg13g2_decap_4 FILLER_45_54 ();
 sg13g2_fill_1 FILLER_45_58 ();
 sg13g2_fill_2 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_69 ();
 sg13g2_fill_1 FILLER_45_71 ();
 sg13g2_decap_4 FILLER_45_77 ();
 sg13g2_fill_1 FILLER_45_81 ();
 sg13g2_fill_2 FILLER_45_107 ();
 sg13g2_fill_2 FILLER_45_140 ();
 sg13g2_fill_1 FILLER_45_142 ();
 sg13g2_decap_4 FILLER_45_164 ();
 sg13g2_fill_1 FILLER_45_172 ();
 sg13g2_fill_2 FILLER_45_207 ();
 sg13g2_fill_2 FILLER_45_238 ();
 sg13g2_fill_1 FILLER_45_244 ();
 sg13g2_fill_2 FILLER_45_271 ();
 sg13g2_fill_2 FILLER_45_277 ();
 sg13g2_fill_2 FILLER_45_284 ();
 sg13g2_decap_4 FILLER_45_290 ();
 sg13g2_fill_1 FILLER_45_294 ();
 sg13g2_decap_4 FILLER_45_308 ();
 sg13g2_fill_2 FILLER_45_312 ();
 sg13g2_decap_8 FILLER_45_318 ();
 sg13g2_decap_8 FILLER_45_325 ();
 sg13g2_decap_8 FILLER_45_332 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_decap_8 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_356 ();
 sg13g2_fill_1 FILLER_45_361 ();
 sg13g2_decap_8 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_373 ();
 sg13g2_fill_2 FILLER_45_390 ();
 sg13g2_decap_4 FILLER_45_396 ();
 sg13g2_fill_1 FILLER_45_412 ();
 sg13g2_fill_1 FILLER_45_458 ();
 sg13g2_fill_1 FILLER_45_463 ();
 sg13g2_fill_1 FILLER_45_621 ();
 sg13g2_fill_2 FILLER_45_653 ();
 sg13g2_fill_1 FILLER_45_673 ();
 sg13g2_fill_1 FILLER_45_677 ();
 sg13g2_decap_8 FILLER_45_690 ();
 sg13g2_fill_1 FILLER_45_836 ();
 sg13g2_fill_1 FILLER_45_841 ();
 sg13g2_fill_2 FILLER_45_857 ();
 sg13g2_fill_2 FILLER_45_885 ();
 sg13g2_fill_2 FILLER_45_912 ();
 sg13g2_fill_1 FILLER_45_914 ();
 sg13g2_fill_1 FILLER_45_928 ();
 sg13g2_fill_1 FILLER_45_963 ();
 sg13g2_fill_1 FILLER_45_968 ();
 sg13g2_fill_1 FILLER_45_973 ();
 sg13g2_fill_1 FILLER_45_1032 ();
 sg13g2_fill_2 FILLER_45_1041 ();
 sg13g2_fill_1 FILLER_45_1050 ();
 sg13g2_fill_2 FILLER_45_1071 ();
 sg13g2_fill_1 FILLER_45_1108 ();
 sg13g2_fill_1 FILLER_45_1112 ();
 sg13g2_fill_1 FILLER_45_1122 ();
 sg13g2_fill_2 FILLER_45_1224 ();
 sg13g2_fill_2 FILLER_45_1230 ();
 sg13g2_fill_1 FILLER_45_1242 ();
 sg13g2_decap_4 FILLER_45_1269 ();
 sg13g2_fill_2 FILLER_45_1286 ();
 sg13g2_fill_1 FILLER_45_1288 ();
 sg13g2_fill_1 FILLER_45_1294 ();
 sg13g2_decap_8 FILLER_45_1299 ();
 sg13g2_fill_2 FILLER_45_1318 ();
 sg13g2_fill_2 FILLER_45_1328 ();
 sg13g2_fill_1 FILLER_45_1330 ();
 sg13g2_decap_8 FILLER_45_1336 ();
 sg13g2_fill_1 FILLER_45_1343 ();
 sg13g2_fill_2 FILLER_45_1359 ();
 sg13g2_fill_2 FILLER_45_1406 ();
 sg13g2_fill_1 FILLER_45_1448 ();
 sg13g2_fill_1 FILLER_45_1464 ();
 sg13g2_fill_1 FILLER_45_1511 ();
 sg13g2_decap_4 FILLER_45_1551 ();
 sg13g2_fill_2 FILLER_45_1555 ();
 sg13g2_fill_1 FILLER_45_1570 ();
 sg13g2_fill_1 FILLER_45_1610 ();
 sg13g2_decap_4 FILLER_45_1615 ();
 sg13g2_decap_8 FILLER_45_1623 ();
 sg13g2_fill_2 FILLER_45_1630 ();
 sg13g2_fill_1 FILLER_45_1632 ();
 sg13g2_fill_1 FILLER_45_1705 ();
 sg13g2_fill_1 FILLER_45_1744 ();
 sg13g2_fill_2 FILLER_45_1793 ();
 sg13g2_fill_1 FILLER_45_1808 ();
 sg13g2_fill_2 FILLER_45_1832 ();
 sg13g2_fill_2 FILLER_45_1860 ();
 sg13g2_fill_1 FILLER_45_1888 ();
 sg13g2_fill_1 FILLER_45_1893 ();
 sg13g2_fill_2 FILLER_45_1946 ();
 sg13g2_fill_1 FILLER_45_1978 ();
 sg13g2_decap_8 FILLER_45_2013 ();
 sg13g2_decap_8 FILLER_45_2020 ();
 sg13g2_fill_1 FILLER_45_2061 ();
 sg13g2_decap_8 FILLER_45_2066 ();
 sg13g2_decap_8 FILLER_45_2081 ();
 sg13g2_decap_8 FILLER_45_2088 ();
 sg13g2_decap_4 FILLER_45_2095 ();
 sg13g2_fill_2 FILLER_45_2099 ();
 sg13g2_decap_8 FILLER_45_2111 ();
 sg13g2_decap_8 FILLER_45_2122 ();
 sg13g2_decap_8 FILLER_45_2129 ();
 sg13g2_decap_8 FILLER_45_2136 ();
 sg13g2_fill_2 FILLER_45_2143 ();
 sg13g2_fill_1 FILLER_45_2145 ();
 sg13g2_fill_2 FILLER_45_2151 ();
 sg13g2_fill_1 FILLER_45_2157 ();
 sg13g2_fill_2 FILLER_45_2163 ();
 sg13g2_fill_2 FILLER_45_2179 ();
 sg13g2_fill_1 FILLER_45_2181 ();
 sg13g2_fill_2 FILLER_45_2193 ();
 sg13g2_fill_1 FILLER_45_2195 ();
 sg13g2_fill_1 FILLER_45_2201 ();
 sg13g2_decap_4 FILLER_45_2213 ();
 sg13g2_decap_8 FILLER_45_2225 ();
 sg13g2_fill_1 FILLER_45_2232 ();
 sg13g2_fill_1 FILLER_45_2241 ();
 sg13g2_fill_1 FILLER_45_2249 ();
 sg13g2_fill_2 FILLER_45_2260 ();
 sg13g2_decap_4 FILLER_45_2272 ();
 sg13g2_decap_4 FILLER_45_2280 ();
 sg13g2_fill_2 FILLER_45_2284 ();
 sg13g2_decap_8 FILLER_45_2294 ();
 sg13g2_fill_2 FILLER_45_2301 ();
 sg13g2_fill_1 FILLER_45_2303 ();
 sg13g2_fill_1 FILLER_45_2328 ();
 sg13g2_decap_8 FILLER_45_2334 ();
 sg13g2_fill_2 FILLER_45_2341 ();
 sg13g2_decap_4 FILLER_45_2348 ();
 sg13g2_fill_1 FILLER_45_2363 ();
 sg13g2_fill_2 FILLER_45_2372 ();
 sg13g2_fill_2 FILLER_45_2383 ();
 sg13g2_decap_8 FILLER_45_2389 ();
 sg13g2_decap_8 FILLER_45_2396 ();
 sg13g2_decap_4 FILLER_45_2403 ();
 sg13g2_fill_1 FILLER_45_2407 ();
 sg13g2_fill_2 FILLER_45_2421 ();
 sg13g2_fill_1 FILLER_45_2434 ();
 sg13g2_fill_1 FILLER_45_2448 ();
 sg13g2_decap_4 FILLER_45_2457 ();
 sg13g2_fill_1 FILLER_45_2461 ();
 sg13g2_fill_1 FILLER_45_2476 ();
 sg13g2_fill_1 FILLER_45_2557 ();
 sg13g2_fill_2 FILLER_45_2564 ();
 sg13g2_decap_8 FILLER_45_2575 ();
 sg13g2_fill_1 FILLER_45_2582 ();
 sg13g2_fill_1 FILLER_45_2630 ();
 sg13g2_decap_8 FILLER_45_2661 ();
 sg13g2_fill_2 FILLER_45_2668 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_decap_4 FILLER_46_35 ();
 sg13g2_fill_2 FILLER_46_65 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_fill_2 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_137 ();
 sg13g2_decap_8 FILLER_46_144 ();
 sg13g2_decap_4 FILLER_46_151 ();
 sg13g2_fill_1 FILLER_46_228 ();
 sg13g2_decap_4 FILLER_46_243 ();
 sg13g2_decap_8 FILLER_46_255 ();
 sg13g2_fill_1 FILLER_46_305 ();
 sg13g2_fill_2 FILLER_46_354 ();
 sg13g2_fill_1 FILLER_46_356 ();
 sg13g2_decap_8 FILLER_46_362 ();
 sg13g2_fill_2 FILLER_46_369 ();
 sg13g2_fill_1 FILLER_46_406 ();
 sg13g2_fill_2 FILLER_46_417 ();
 sg13g2_fill_1 FILLER_46_445 ();
 sg13g2_fill_2 FILLER_46_450 ();
 sg13g2_fill_1 FILLER_46_452 ();
 sg13g2_fill_2 FILLER_46_462 ();
 sg13g2_decap_4 FILLER_46_485 ();
 sg13g2_fill_2 FILLER_46_510 ();
 sg13g2_fill_1 FILLER_46_512 ();
 sg13g2_fill_1 FILLER_46_550 ();
 sg13g2_fill_2 FILLER_46_577 ();
 sg13g2_fill_1 FILLER_46_579 ();
 sg13g2_decap_4 FILLER_46_605 ();
 sg13g2_fill_2 FILLER_46_613 ();
 sg13g2_fill_1 FILLER_46_623 ();
 sg13g2_decap_4 FILLER_46_671 ();
 sg13g2_fill_2 FILLER_46_707 ();
 sg13g2_fill_1 FILLER_46_709 ();
 sg13g2_fill_1 FILLER_46_749 ();
 sg13g2_fill_2 FILLER_46_793 ();
 sg13g2_fill_1 FILLER_46_835 ();
 sg13g2_fill_1 FILLER_46_846 ();
 sg13g2_fill_1 FILLER_46_854 ();
 sg13g2_fill_1 FILLER_46_886 ();
 sg13g2_fill_1 FILLER_46_897 ();
 sg13g2_fill_2 FILLER_46_907 ();
 sg13g2_fill_1 FILLER_46_909 ();
 sg13g2_decap_4 FILLER_46_940 ();
 sg13g2_fill_1 FILLER_46_944 ();
 sg13g2_fill_1 FILLER_46_949 ();
 sg13g2_decap_4 FILLER_46_954 ();
 sg13g2_fill_2 FILLER_46_958 ();
 sg13g2_fill_2 FILLER_46_964 ();
 sg13g2_fill_1 FILLER_46_978 ();
 sg13g2_fill_2 FILLER_46_1025 ();
 sg13g2_fill_2 FILLER_46_1056 ();
 sg13g2_fill_1 FILLER_46_1080 ();
 sg13g2_fill_1 FILLER_46_1099 ();
 sg13g2_fill_1 FILLER_46_1150 ();
 sg13g2_fill_1 FILLER_46_1157 ();
 sg13g2_fill_2 FILLER_46_1165 ();
 sg13g2_fill_1 FILLER_46_1270 ();
 sg13g2_fill_2 FILLER_46_1311 ();
 sg13g2_fill_2 FILLER_46_1325 ();
 sg13g2_fill_1 FILLER_46_1339 ();
 sg13g2_fill_1 FILLER_46_1344 ();
 sg13g2_fill_2 FILLER_46_1369 ();
 sg13g2_fill_1 FILLER_46_1385 ();
 sg13g2_fill_1 FILLER_46_1390 ();
 sg13g2_fill_1 FILLER_46_1395 ();
 sg13g2_fill_1 FILLER_46_1400 ();
 sg13g2_fill_2 FILLER_46_1477 ();
 sg13g2_decap_4 FILLER_46_1514 ();
 sg13g2_fill_1 FILLER_46_1518 ();
 sg13g2_decap_8 FILLER_46_1523 ();
 sg13g2_decap_8 FILLER_46_1530 ();
 sg13g2_fill_2 FILLER_46_1537 ();
 sg13g2_fill_2 FILLER_46_1543 ();
 sg13g2_fill_1 FILLER_46_1606 ();
 sg13g2_decap_8 FILLER_46_1638 ();
 sg13g2_fill_2 FILLER_46_1645 ();
 sg13g2_fill_1 FILLER_46_1647 ();
 sg13g2_fill_2 FILLER_46_1652 ();
 sg13g2_decap_8 FILLER_46_1687 ();
 sg13g2_decap_8 FILLER_46_1694 ();
 sg13g2_fill_1 FILLER_46_1701 ();
 sg13g2_fill_2 FILLER_46_1709 ();
 sg13g2_fill_2 FILLER_46_1715 ();
 sg13g2_fill_2 FILLER_46_1735 ();
 sg13g2_fill_1 FILLER_46_1745 ();
 sg13g2_fill_2 FILLER_46_1759 ();
 sg13g2_fill_1 FILLER_46_1764 ();
 sg13g2_fill_2 FILLER_46_1786 ();
 sg13g2_fill_2 FILLER_46_1800 ();
 sg13g2_fill_2 FILLER_46_1806 ();
 sg13g2_fill_2 FILLER_46_1819 ();
 sg13g2_fill_1 FILLER_46_1825 ();
 sg13g2_fill_1 FILLER_46_1851 ();
 sg13g2_fill_2 FILLER_46_1856 ();
 sg13g2_fill_1 FILLER_46_1880 ();
 sg13g2_fill_2 FILLER_46_1886 ();
 sg13g2_fill_1 FILLER_46_1907 ();
 sg13g2_fill_2 FILLER_46_1912 ();
 sg13g2_fill_2 FILLER_46_1949 ();
 sg13g2_fill_1 FILLER_46_1996 ();
 sg13g2_fill_2 FILLER_46_2009 ();
 sg13g2_fill_2 FILLER_46_2050 ();
 sg13g2_decap_4 FILLER_46_2066 ();
 sg13g2_fill_1 FILLER_46_2096 ();
 sg13g2_fill_1 FILLER_46_2102 ();
 sg13g2_fill_1 FILLER_46_2129 ();
 sg13g2_fill_1 FILLER_46_2135 ();
 sg13g2_fill_1 FILLER_46_2178 ();
 sg13g2_fill_1 FILLER_46_2210 ();
 sg13g2_fill_2 FILLER_46_2216 ();
 sg13g2_fill_2 FILLER_46_2222 ();
 sg13g2_fill_1 FILLER_46_2224 ();
 sg13g2_fill_2 FILLER_46_2229 ();
 sg13g2_fill_2 FILLER_46_2235 ();
 sg13g2_fill_1 FILLER_46_2237 ();
 sg13g2_fill_2 FILLER_46_2242 ();
 sg13g2_fill_1 FILLER_46_2244 ();
 sg13g2_fill_2 FILLER_46_2253 ();
 sg13g2_decap_4 FILLER_46_2265 ();
 sg13g2_fill_2 FILLER_46_2274 ();
 sg13g2_fill_1 FILLER_46_2276 ();
 sg13g2_decap_4 FILLER_46_2280 ();
 sg13g2_fill_1 FILLER_46_2288 ();
 sg13g2_decap_4 FILLER_46_2307 ();
 sg13g2_fill_1 FILLER_46_2323 ();
 sg13g2_decap_8 FILLER_46_2343 ();
 sg13g2_fill_1 FILLER_46_2359 ();
 sg13g2_fill_2 FILLER_46_2383 ();
 sg13g2_fill_1 FILLER_46_2397 ();
 sg13g2_fill_2 FILLER_46_2417 ();
 sg13g2_fill_1 FILLER_46_2419 ();
 sg13g2_fill_2 FILLER_46_2424 ();
 sg13g2_fill_2 FILLER_46_2436 ();
 sg13g2_fill_1 FILLER_46_2438 ();
 sg13g2_decap_8 FILLER_46_2459 ();
 sg13g2_fill_2 FILLER_46_2466 ();
 sg13g2_fill_1 FILLER_46_2468 ();
 sg13g2_fill_1 FILLER_46_2512 ();
 sg13g2_fill_1 FILLER_46_2524 ();
 sg13g2_fill_1 FILLER_46_2541 ();
 sg13g2_fill_2 FILLER_46_2547 ();
 sg13g2_fill_2 FILLER_46_2559 ();
 sg13g2_decap_4 FILLER_46_2575 ();
 sg13g2_fill_1 FILLER_46_2579 ();
 sg13g2_fill_2 FILLER_46_2588 ();
 sg13g2_fill_1 FILLER_46_2590 ();
 sg13g2_decap_4 FILLER_46_2596 ();
 sg13g2_fill_1 FILLER_46_2600 ();
 sg13g2_fill_2 FILLER_46_2622 ();
 sg13g2_fill_1 FILLER_46_2665 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_4 ();
 sg13g2_decap_4 FILLER_47_39 ();
 sg13g2_fill_2 FILLER_47_43 ();
 sg13g2_fill_2 FILLER_47_89 ();
 sg13g2_decap_8 FILLER_47_116 ();
 sg13g2_fill_1 FILLER_47_123 ();
 sg13g2_decap_8 FILLER_47_150 ();
 sg13g2_decap_8 FILLER_47_157 ();
 sg13g2_fill_2 FILLER_47_164 ();
 sg13g2_fill_1 FILLER_47_166 ();
 sg13g2_fill_1 FILLER_47_219 ();
 sg13g2_fill_1 FILLER_47_224 ();
 sg13g2_fill_2 FILLER_47_231 ();
 sg13g2_decap_4 FILLER_47_236 ();
 sg13g2_fill_2 FILLER_47_305 ();
 sg13g2_fill_1 FILLER_47_307 ();
 sg13g2_fill_1 FILLER_47_347 ();
 sg13g2_fill_2 FILLER_47_374 ();
 sg13g2_fill_2 FILLER_47_380 ();
 sg13g2_decap_8 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_47_415 ();
 sg13g2_fill_2 FILLER_47_422 ();
 sg13g2_fill_2 FILLER_47_462 ();
 sg13g2_fill_2 FILLER_47_478 ();
 sg13g2_fill_1 FILLER_47_480 ();
 sg13g2_fill_1 FILLER_47_511 ();
 sg13g2_fill_2 FILLER_47_517 ();
 sg13g2_fill_1 FILLER_47_519 ();
 sg13g2_fill_2 FILLER_47_550 ();
 sg13g2_fill_1 FILLER_47_591 ();
 sg13g2_fill_2 FILLER_47_596 ();
 sg13g2_fill_1 FILLER_47_602 ();
 sg13g2_fill_1 FILLER_47_634 ();
 sg13g2_fill_1 FILLER_47_643 ();
 sg13g2_decap_4 FILLER_47_668 ();
 sg13g2_fill_2 FILLER_47_672 ();
 sg13g2_fill_1 FILLER_47_700 ();
 sg13g2_fill_2 FILLER_47_744 ();
 sg13g2_fill_1 FILLER_47_759 ();
 sg13g2_fill_2 FILLER_47_776 ();
 sg13g2_fill_1 FILLER_47_787 ();
 sg13g2_fill_2 FILLER_47_818 ();
 sg13g2_fill_1 FILLER_47_833 ();
 sg13g2_fill_2 FILLER_47_839 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_fill_1 FILLER_47_896 ();
 sg13g2_fill_1 FILLER_47_954 ();
 sg13g2_fill_2 FILLER_47_976 ();
 sg13g2_fill_2 FILLER_47_1001 ();
 sg13g2_fill_1 FILLER_47_1011 ();
 sg13g2_fill_2 FILLER_47_1046 ();
 sg13g2_fill_1 FILLER_47_1129 ();
 sg13g2_fill_2 FILLER_47_1159 ();
 sg13g2_fill_2 FILLER_47_1231 ();
 sg13g2_fill_1 FILLER_47_1233 ();
 sg13g2_fill_1 FILLER_47_1243 ();
 sg13g2_fill_2 FILLER_47_1248 ();
 sg13g2_decap_8 FILLER_47_1258 ();
 sg13g2_decap_8 FILLER_47_1265 ();
 sg13g2_decap_4 FILLER_47_1272 ();
 sg13g2_fill_2 FILLER_47_1276 ();
 sg13g2_decap_4 FILLER_47_1282 ();
 sg13g2_fill_1 FILLER_47_1327 ();
 sg13g2_fill_1 FILLER_47_1370 ();
 sg13g2_fill_1 FILLER_47_1374 ();
 sg13g2_fill_1 FILLER_47_1430 ();
 sg13g2_fill_1 FILLER_47_1450 ();
 sg13g2_fill_1 FILLER_47_1492 ();
 sg13g2_decap_8 FILLER_47_1505 ();
 sg13g2_decap_8 FILLER_47_1512 ();
 sg13g2_decap_4 FILLER_47_1519 ();
 sg13g2_fill_2 FILLER_47_1523 ();
 sg13g2_fill_1 FILLER_47_1551 ();
 sg13g2_decap_8 FILLER_47_1624 ();
 sg13g2_decap_8 FILLER_47_1631 ();
 sg13g2_decap_8 FILLER_47_1638 ();
 sg13g2_decap_8 FILLER_47_1645 ();
 sg13g2_decap_8 FILLER_47_1652 ();
 sg13g2_decap_8 FILLER_47_1659 ();
 sg13g2_fill_2 FILLER_47_1666 ();
 sg13g2_decap_8 FILLER_47_1672 ();
 sg13g2_fill_1 FILLER_47_1692 ();
 sg13g2_fill_2 FILLER_47_1697 ();
 sg13g2_fill_1 FILLER_47_1699 ();
 sg13g2_fill_1 FILLER_47_1727 ();
 sg13g2_fill_1 FILLER_47_1809 ();
 sg13g2_fill_1 FILLER_47_1830 ();
 sg13g2_fill_1 FILLER_47_1836 ();
 sg13g2_fill_2 FILLER_47_1846 ();
 sg13g2_fill_1 FILLER_47_1900 ();
 sg13g2_fill_1 FILLER_47_1914 ();
 sg13g2_fill_1 FILLER_47_1935 ();
 sg13g2_fill_2 FILLER_47_2010 ();
 sg13g2_decap_4 FILLER_47_2016 ();
 sg13g2_fill_1 FILLER_47_2020 ();
 sg13g2_fill_1 FILLER_47_2029 ();
 sg13g2_fill_2 FILLER_47_2043 ();
 sg13g2_fill_1 FILLER_47_2050 ();
 sg13g2_fill_2 FILLER_47_2055 ();
 sg13g2_decap_8 FILLER_47_2088 ();
 sg13g2_fill_2 FILLER_47_2095 ();
 sg13g2_decap_4 FILLER_47_2107 ();
 sg13g2_fill_1 FILLER_47_2111 ();
 sg13g2_decap_8 FILLER_47_2116 ();
 sg13g2_decap_4 FILLER_47_2123 ();
 sg13g2_fill_2 FILLER_47_2127 ();
 sg13g2_decap_4 FILLER_47_2181 ();
 sg13g2_fill_1 FILLER_47_2189 ();
 sg13g2_decap_8 FILLER_47_2201 ();
 sg13g2_fill_2 FILLER_47_2208 ();
 sg13g2_fill_1 FILLER_47_2210 ();
 sg13g2_fill_1 FILLER_47_2231 ();
 sg13g2_fill_1 FILLER_47_2236 ();
 sg13g2_fill_2 FILLER_47_2242 ();
 sg13g2_fill_1 FILLER_47_2244 ();
 sg13g2_fill_2 FILLER_47_2250 ();
 sg13g2_decap_8 FILLER_47_2257 ();
 sg13g2_decap_8 FILLER_47_2264 ();
 sg13g2_decap_8 FILLER_47_2271 ();
 sg13g2_decap_4 FILLER_47_2278 ();
 sg13g2_fill_1 FILLER_47_2282 ();
 sg13g2_fill_1 FILLER_47_2292 ();
 sg13g2_fill_1 FILLER_47_2311 ();
 sg13g2_fill_2 FILLER_47_2317 ();
 sg13g2_fill_1 FILLER_47_2323 ();
 sg13g2_fill_1 FILLER_47_2338 ();
 sg13g2_decap_4 FILLER_47_2343 ();
 sg13g2_fill_1 FILLER_47_2353 ();
 sg13g2_decap_8 FILLER_47_2401 ();
 sg13g2_fill_1 FILLER_47_2408 ();
 sg13g2_fill_1 FILLER_47_2413 ();
 sg13g2_decap_4 FILLER_47_2418 ();
 sg13g2_decap_4 FILLER_47_2431 ();
 sg13g2_fill_1 FILLER_47_2435 ();
 sg13g2_decap_8 FILLER_47_2445 ();
 sg13g2_fill_1 FILLER_47_2452 ();
 sg13g2_fill_1 FILLER_47_2462 ();
 sg13g2_fill_2 FILLER_47_2468 ();
 sg13g2_fill_1 FILLER_47_2480 ();
 sg13g2_fill_1 FILLER_47_2487 ();
 sg13g2_fill_2 FILLER_47_2494 ();
 sg13g2_fill_2 FILLER_47_2502 ();
 sg13g2_fill_1 FILLER_47_2504 ();
 sg13g2_fill_1 FILLER_47_2510 ();
 sg13g2_fill_1 FILLER_47_2523 ();
 sg13g2_decap_4 FILLER_47_2536 ();
 sg13g2_fill_1 FILLER_47_2540 ();
 sg13g2_fill_2 FILLER_47_2554 ();
 sg13g2_fill_1 FILLER_47_2556 ();
 sg13g2_fill_1 FILLER_47_2577 ();
 sg13g2_decap_4 FILLER_47_2582 ();
 sg13g2_fill_1 FILLER_47_2586 ();
 sg13g2_decap_4 FILLER_47_2591 ();
 sg13g2_decap_4 FILLER_47_2613 ();
 sg13g2_fill_1 FILLER_47_2637 ();
 sg13g2_decap_8 FILLER_47_2659 ();
 sg13g2_decap_4 FILLER_47_2666 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_13 ();
 sg13g2_fill_1 FILLER_48_18 ();
 sg13g2_fill_1 FILLER_48_53 ();
 sg13g2_fill_2 FILLER_48_80 ();
 sg13g2_fill_2 FILLER_48_87 ();
 sg13g2_fill_1 FILLER_48_89 ();
 sg13g2_decap_4 FILLER_48_120 ();
 sg13g2_decap_8 FILLER_48_162 ();
 sg13g2_fill_1 FILLER_48_169 ();
 sg13g2_fill_1 FILLER_48_212 ();
 sg13g2_decap_4 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_272 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_fill_2 FILLER_48_347 ();
 sg13g2_fill_2 FILLER_48_380 ();
 sg13g2_fill_1 FILLER_48_382 ();
 sg13g2_decap_8 FILLER_48_409 ();
 sg13g2_decap_8 FILLER_48_429 ();
 sg13g2_fill_1 FILLER_48_484 ();
 sg13g2_fill_1 FILLER_48_535 ();
 sg13g2_fill_2 FILLER_48_560 ();
 sg13g2_fill_1 FILLER_48_566 ();
 sg13g2_fill_1 FILLER_48_572 ();
 sg13g2_fill_1 FILLER_48_577 ();
 sg13g2_fill_1 FILLER_48_582 ();
 sg13g2_fill_1 FILLER_48_609 ();
 sg13g2_fill_2 FILLER_48_632 ();
 sg13g2_fill_1 FILLER_48_649 ();
 sg13g2_fill_2 FILLER_48_720 ();
 sg13g2_fill_2 FILLER_48_753 ();
 sg13g2_fill_1 FILLER_48_768 ();
 sg13g2_fill_2 FILLER_48_829 ();
 sg13g2_fill_1 FILLER_48_862 ();
 sg13g2_fill_1 FILLER_48_873 ();
 sg13g2_fill_2 FILLER_48_878 ();
 sg13g2_fill_1 FILLER_48_889 ();
 sg13g2_fill_1 FILLER_48_898 ();
 sg13g2_fill_1 FILLER_48_908 ();
 sg13g2_fill_2 FILLER_48_921 ();
 sg13g2_fill_1 FILLER_48_953 ();
 sg13g2_fill_1 FILLER_48_959 ();
 sg13g2_fill_1 FILLER_48_965 ();
 sg13g2_fill_1 FILLER_48_974 ();
 sg13g2_fill_1 FILLER_48_1055 ();
 sg13g2_fill_2 FILLER_48_1150 ();
 sg13g2_fill_1 FILLER_48_1159 ();
 sg13g2_fill_1 FILLER_48_1205 ();
 sg13g2_fill_2 FILLER_48_1213 ();
 sg13g2_fill_2 FILLER_48_1253 ();
 sg13g2_decap_8 FILLER_48_1259 ();
 sg13g2_fill_1 FILLER_48_1266 ();
 sg13g2_fill_2 FILLER_48_1271 ();
 sg13g2_fill_1 FILLER_48_1289 ();
 sg13g2_fill_1 FILLER_48_1347 ();
 sg13g2_fill_1 FILLER_48_1366 ();
 sg13g2_fill_1 FILLER_48_1371 ();
 sg13g2_fill_1 FILLER_48_1427 ();
 sg13g2_fill_2 FILLER_48_1475 ();
 sg13g2_fill_2 FILLER_48_1529 ();
 sg13g2_fill_2 FILLER_48_1544 ();
 sg13g2_fill_2 FILLER_48_1583 ();
 sg13g2_fill_2 FILLER_48_1589 ();
 sg13g2_fill_2 FILLER_48_1605 ();
 sg13g2_fill_1 FILLER_48_1619 ();
 sg13g2_decap_8 FILLER_48_1651 ();
 sg13g2_fill_2 FILLER_48_1658 ();
 sg13g2_fill_2 FILLER_48_1728 ();
 sg13g2_fill_2 FILLER_48_1829 ();
 sg13g2_fill_2 FILLER_48_1840 ();
 sg13g2_fill_1 FILLER_48_1887 ();
 sg13g2_fill_1 FILLER_48_1891 ();
 sg13g2_fill_1 FILLER_48_1896 ();
 sg13g2_fill_2 FILLER_48_1943 ();
 sg13g2_fill_1 FILLER_48_1957 ();
 sg13g2_fill_2 FILLER_48_1969 ();
 sg13g2_fill_1 FILLER_48_1984 ();
 sg13g2_decap_8 FILLER_48_2019 ();
 sg13g2_fill_2 FILLER_48_2026 ();
 sg13g2_fill_2 FILLER_48_2037 ();
 sg13g2_fill_1 FILLER_48_2039 ();
 sg13g2_decap_8 FILLER_48_2077 ();
 sg13g2_decap_4 FILLER_48_2084 ();
 sg13g2_fill_2 FILLER_48_2088 ();
 sg13g2_decap_4 FILLER_48_2116 ();
 sg13g2_fill_2 FILLER_48_2120 ();
 sg13g2_fill_1 FILLER_48_2126 ();
 sg13g2_decap_8 FILLER_48_2146 ();
 sg13g2_fill_1 FILLER_48_2166 ();
 sg13g2_fill_1 FILLER_48_2173 ();
 sg13g2_fill_1 FILLER_48_2179 ();
 sg13g2_fill_1 FILLER_48_2193 ();
 sg13g2_fill_2 FILLER_48_2200 ();
 sg13g2_fill_1 FILLER_48_2206 ();
 sg13g2_fill_2 FILLER_48_2217 ();
 sg13g2_fill_2 FILLER_48_2223 ();
 sg13g2_fill_2 FILLER_48_2231 ();
 sg13g2_fill_2 FILLER_48_2237 ();
 sg13g2_decap_8 FILLER_48_2252 ();
 sg13g2_decap_8 FILLER_48_2259 ();
 sg13g2_fill_2 FILLER_48_2266 ();
 sg13g2_decap_4 FILLER_48_2286 ();
 sg13g2_decap_8 FILLER_48_2294 ();
 sg13g2_fill_2 FILLER_48_2301 ();
 sg13g2_fill_1 FILLER_48_2307 ();
 sg13g2_fill_2 FILLER_48_2312 ();
 sg13g2_fill_1 FILLER_48_2319 ();
 sg13g2_fill_2 FILLER_48_2324 ();
 sg13g2_fill_2 FILLER_48_2334 ();
 sg13g2_decap_4 FILLER_48_2342 ();
 sg13g2_fill_1 FILLER_48_2346 ();
 sg13g2_fill_2 FILLER_48_2350 ();
 sg13g2_fill_1 FILLER_48_2352 ();
 sg13g2_fill_1 FILLER_48_2369 ();
 sg13g2_fill_1 FILLER_48_2374 ();
 sg13g2_fill_1 FILLER_48_2380 ();
 sg13g2_fill_1 FILLER_48_2386 ();
 sg13g2_fill_1 FILLER_48_2400 ();
 sg13g2_fill_2 FILLER_48_2406 ();
 sg13g2_fill_1 FILLER_48_2408 ();
 sg13g2_decap_8 FILLER_48_2413 ();
 sg13g2_fill_1 FILLER_48_2420 ();
 sg13g2_fill_2 FILLER_48_2433 ();
 sg13g2_decap_8 FILLER_48_2440 ();
 sg13g2_decap_4 FILLER_48_2447 ();
 sg13g2_fill_2 FILLER_48_2451 ();
 sg13g2_fill_1 FILLER_48_2463 ();
 sg13g2_fill_2 FILLER_48_2468 ();
 sg13g2_fill_1 FILLER_48_2470 ();
 sg13g2_fill_1 FILLER_48_2488 ();
 sg13g2_fill_2 FILLER_48_2494 ();
 sg13g2_fill_1 FILLER_48_2496 ();
 sg13g2_decap_4 FILLER_48_2533 ();
 sg13g2_fill_1 FILLER_48_2537 ();
 sg13g2_fill_1 FILLER_48_2543 ();
 sg13g2_fill_2 FILLER_48_2549 ();
 sg13g2_fill_1 FILLER_48_2551 ();
 sg13g2_decap_8 FILLER_48_2558 ();
 sg13g2_fill_2 FILLER_48_2565 ();
 sg13g2_decap_8 FILLER_48_2593 ();
 sg13g2_decap_4 FILLER_48_2664 ();
 sg13g2_fill_2 FILLER_48_2668 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_28 ();
 sg13g2_decap_4 FILLER_49_41 ();
 sg13g2_fill_1 FILLER_49_45 ();
 sg13g2_fill_2 FILLER_49_59 ();
 sg13g2_fill_2 FILLER_49_65 ();
 sg13g2_fill_1 FILLER_49_67 ();
 sg13g2_decap_4 FILLER_49_72 ();
 sg13g2_fill_2 FILLER_49_123 ();
 sg13g2_fill_1 FILLER_49_125 ();
 sg13g2_fill_1 FILLER_49_135 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_decap_4 FILLER_49_228 ();
 sg13g2_fill_2 FILLER_49_236 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_285 ();
 sg13g2_decap_8 FILLER_49_292 ();
 sg13g2_decap_4 FILLER_49_299 ();
 sg13g2_fill_2 FILLER_49_312 ();
 sg13g2_fill_2 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_335 ();
 sg13g2_decap_4 FILLER_49_342 ();
 sg13g2_fill_1 FILLER_49_346 ();
 sg13g2_fill_1 FILLER_49_351 ();
 sg13g2_fill_1 FILLER_49_356 ();
 sg13g2_fill_2 FILLER_49_391 ();
 sg13g2_fill_1 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_419 ();
 sg13g2_fill_1 FILLER_49_426 ();
 sg13g2_fill_2 FILLER_49_457 ();
 sg13g2_fill_1 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_509 ();
 sg13g2_fill_1 FILLER_49_523 ();
 sg13g2_decap_4 FILLER_49_528 ();
 sg13g2_fill_1 FILLER_49_560 ();
 sg13g2_fill_2 FILLER_49_596 ();
 sg13g2_fill_1 FILLER_49_602 ();
 sg13g2_fill_2 FILLER_49_663 ();
 sg13g2_fill_1 FILLER_49_674 ();
 sg13g2_fill_1 FILLER_49_807 ();
 sg13g2_fill_1 FILLER_49_812 ();
 sg13g2_fill_2 FILLER_49_824 ();
 sg13g2_fill_1 FILLER_49_878 ();
 sg13g2_fill_1 FILLER_49_918 ();
 sg13g2_fill_1 FILLER_49_941 ();
 sg13g2_fill_1 FILLER_49_946 ();
 sg13g2_fill_1 FILLER_49_978 ();
 sg13g2_fill_1 FILLER_49_988 ();
 sg13g2_fill_1 FILLER_49_1018 ();
 sg13g2_fill_1 FILLER_49_1035 ();
 sg13g2_fill_1 FILLER_49_1070 ();
 sg13g2_fill_2 FILLER_49_1076 ();
 sg13g2_fill_1 FILLER_49_1104 ();
 sg13g2_fill_2 FILLER_49_1160 ();
 sg13g2_fill_2 FILLER_49_1255 ();
 sg13g2_fill_2 FILLER_49_1293 ();
 sg13g2_decap_8 FILLER_49_1318 ();
 sg13g2_fill_2 FILLER_49_1325 ();
 sg13g2_fill_1 FILLER_49_1331 ();
 sg13g2_fill_1 FILLER_49_1403 ();
 sg13g2_fill_1 FILLER_49_1450 ();
 sg13g2_fill_1 FILLER_49_1460 ();
 sg13g2_fill_2 FILLER_49_1475 ();
 sg13g2_decap_8 FILLER_49_1520 ();
 sg13g2_decap_4 FILLER_49_1527 ();
 sg13g2_fill_2 FILLER_49_1531 ();
 sg13g2_fill_1 FILLER_49_1563 ();
 sg13g2_fill_1 FILLER_49_1613 ();
 sg13g2_fill_2 FILLER_49_1618 ();
 sg13g2_fill_1 FILLER_49_1624 ();
 sg13g2_decap_4 FILLER_49_1651 ();
 sg13g2_fill_1 FILLER_49_1655 ();
 sg13g2_fill_2 FILLER_49_1690 ();
 sg13g2_fill_1 FILLER_49_1697 ();
 sg13g2_fill_2 FILLER_49_1746 ();
 sg13g2_fill_1 FILLER_49_1794 ();
 sg13g2_fill_1 FILLER_49_1816 ();
 sg13g2_fill_2 FILLER_49_1855 ();
 sg13g2_fill_2 FILLER_49_1882 ();
 sg13g2_fill_2 FILLER_49_1887 ();
 sg13g2_fill_1 FILLER_49_1952 ();
 sg13g2_fill_2 FILLER_49_1966 ();
 sg13g2_fill_1 FILLER_49_1976 ();
 sg13g2_fill_2 FILLER_49_2011 ();
 sg13g2_fill_1 FILLER_49_2026 ();
 sg13g2_fill_2 FILLER_49_2031 ();
 sg13g2_fill_1 FILLER_49_2033 ();
 sg13g2_decap_4 FILLER_49_2083 ();
 sg13g2_fill_1 FILLER_49_2087 ();
 sg13g2_decap_8 FILLER_49_2118 ();
 sg13g2_fill_2 FILLER_49_2125 ();
 sg13g2_fill_1 FILLER_49_2169 ();
 sg13g2_fill_2 FILLER_49_2175 ();
 sg13g2_fill_1 FILLER_49_2187 ();
 sg13g2_fill_1 FILLER_49_2192 ();
 sg13g2_fill_2 FILLER_49_2205 ();
 sg13g2_decap_8 FILLER_49_2215 ();
 sg13g2_fill_2 FILLER_49_2222 ();
 sg13g2_fill_1 FILLER_49_2224 ();
 sg13g2_decap_8 FILLER_49_2233 ();
 sg13g2_fill_2 FILLER_49_2240 ();
 sg13g2_fill_2 FILLER_49_2246 ();
 sg13g2_fill_2 FILLER_49_2256 ();
 sg13g2_decap_4 FILLER_49_2266 ();
 sg13g2_fill_2 FILLER_49_2276 ();
 sg13g2_fill_1 FILLER_49_2278 ();
 sg13g2_fill_2 FILLER_49_2309 ();
 sg13g2_fill_2 FILLER_49_2323 ();
 sg13g2_fill_1 FILLER_49_2343 ();
 sg13g2_fill_1 FILLER_49_2367 ();
 sg13g2_decap_8 FILLER_49_2383 ();
 sg13g2_fill_2 FILLER_49_2390 ();
 sg13g2_fill_1 FILLER_49_2398 ();
 sg13g2_fill_1 FILLER_49_2404 ();
 sg13g2_fill_1 FILLER_49_2411 ();
 sg13g2_fill_1 FILLER_49_2424 ();
 sg13g2_fill_1 FILLER_49_2456 ();
 sg13g2_fill_2 FILLER_49_2462 ();
 sg13g2_fill_2 FILLER_49_2469 ();
 sg13g2_fill_2 FILLER_49_2477 ();
 sg13g2_fill_1 FILLER_49_2479 ();
 sg13g2_fill_1 FILLER_49_2492 ();
 sg13g2_fill_1 FILLER_49_2502 ();
 sg13g2_decap_8 FILLER_49_2511 ();
 sg13g2_decap_8 FILLER_49_2518 ();
 sg13g2_fill_2 FILLER_49_2525 ();
 sg13g2_fill_1 FILLER_49_2527 ();
 sg13g2_fill_1 FILLER_49_2533 ();
 sg13g2_fill_2 FILLER_49_2539 ();
 sg13g2_decap_8 FILLER_49_2545 ();
 sg13g2_fill_1 FILLER_49_2558 ();
 sg13g2_decap_8 FILLER_49_2592 ();
 sg13g2_decap_4 FILLER_49_2599 ();
 sg13g2_fill_1 FILLER_49_2609 ();
 sg13g2_fill_1 FILLER_49_2618 ();
 sg13g2_fill_1 FILLER_49_2623 ();
 sg13g2_fill_2 FILLER_49_2629 ();
 sg13g2_decap_8 FILLER_49_2652 ();
 sg13g2_decap_8 FILLER_49_2659 ();
 sg13g2_decap_4 FILLER_49_2666 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_14 ();
 sg13g2_fill_2 FILLER_50_58 ();
 sg13g2_fill_1 FILLER_50_60 ();
 sg13g2_fill_1 FILLER_50_70 ();
 sg13g2_fill_1 FILLER_50_80 ();
 sg13g2_fill_2 FILLER_50_116 ();
 sg13g2_fill_1 FILLER_50_131 ();
 sg13g2_fill_1 FILLER_50_163 ();
 sg13g2_fill_1 FILLER_50_168 ();
 sg13g2_fill_1 FILLER_50_175 ();
 sg13g2_fill_2 FILLER_50_215 ();
 sg13g2_fill_2 FILLER_50_221 ();
 sg13g2_fill_2 FILLER_50_231 ();
 sg13g2_fill_1 FILLER_50_254 ();
 sg13g2_fill_2 FILLER_50_276 ();
 sg13g2_fill_1 FILLER_50_278 ();
 sg13g2_fill_2 FILLER_50_283 ();
 sg13g2_fill_1 FILLER_50_285 ();
 sg13g2_decap_4 FILLER_50_358 ();
 sg13g2_fill_1 FILLER_50_366 ();
 sg13g2_fill_1 FILLER_50_388 ();
 sg13g2_fill_2 FILLER_50_398 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_1 FILLER_50_440 ();
 sg13g2_fill_2 FILLER_50_445 ();
 sg13g2_fill_1 FILLER_50_454 ();
 sg13g2_fill_1 FILLER_50_459 ();
 sg13g2_decap_8 FILLER_50_471 ();
 sg13g2_decap_4 FILLER_50_478 ();
 sg13g2_fill_1 FILLER_50_482 ();
 sg13g2_decap_4 FILLER_50_487 ();
 sg13g2_fill_2 FILLER_50_491 ();
 sg13g2_decap_8 FILLER_50_497 ();
 sg13g2_decap_8 FILLER_50_504 ();
 sg13g2_decap_8 FILLER_50_511 ();
 sg13g2_decap_4 FILLER_50_518 ();
 sg13g2_fill_1 FILLER_50_522 ();
 sg13g2_decap_8 FILLER_50_526 ();
 sg13g2_decap_4 FILLER_50_533 ();
 sg13g2_decap_8 FILLER_50_544 ();
 sg13g2_decap_8 FILLER_50_551 ();
 sg13g2_decap_8 FILLER_50_558 ();
 sg13g2_fill_1 FILLER_50_565 ();
 sg13g2_decap_8 FILLER_50_570 ();
 sg13g2_decap_4 FILLER_50_577 ();
 sg13g2_fill_2 FILLER_50_607 ();
 sg13g2_fill_2 FILLER_50_623 ();
 sg13g2_fill_1 FILLER_50_636 ();
 sg13g2_fill_1 FILLER_50_681 ();
 sg13g2_fill_2 FILLER_50_705 ();
 sg13g2_fill_1 FILLER_50_737 ();
 sg13g2_fill_2 FILLER_50_833 ();
 sg13g2_fill_1 FILLER_50_909 ();
 sg13g2_decap_8 FILLER_50_935 ();
 sg13g2_decap_8 FILLER_50_942 ();
 sg13g2_decap_4 FILLER_50_949 ();
 sg13g2_fill_1 FILLER_50_953 ();
 sg13g2_fill_1 FILLER_50_958 ();
 sg13g2_fill_2 FILLER_50_993 ();
 sg13g2_fill_2 FILLER_50_999 ();
 sg13g2_fill_1 FILLER_50_1001 ();
 sg13g2_fill_1 FILLER_50_1026 ();
 sg13g2_fill_1 FILLER_50_1031 ();
 sg13g2_fill_2 FILLER_50_1066 ();
 sg13g2_fill_2 FILLER_50_1071 ();
 sg13g2_fill_1 FILLER_50_1098 ();
 sg13g2_fill_1 FILLER_50_1192 ();
 sg13g2_fill_1 FILLER_50_1204 ();
 sg13g2_fill_2 FILLER_50_1221 ();
 sg13g2_fill_2 FILLER_50_1252 ();
 sg13g2_fill_1 FILLER_50_1327 ();
 sg13g2_decap_8 FILLER_50_1332 ();
 sg13g2_decap_8 FILLER_50_1339 ();
 sg13g2_decap_4 FILLER_50_1363 ();
 sg13g2_fill_1 FILLER_50_1377 ();
 sg13g2_fill_2 FILLER_50_1486 ();
 sg13g2_decap_4 FILLER_50_1495 ();
 sg13g2_fill_1 FILLER_50_1499 ();
 sg13g2_decap_4 FILLER_50_1504 ();
 sg13g2_fill_2 FILLER_50_1516 ();
 sg13g2_fill_1 FILLER_50_1518 ();
 sg13g2_decap_8 FILLER_50_1523 ();
 sg13g2_decap_8 FILLER_50_1530 ();
 sg13g2_fill_2 FILLER_50_1537 ();
 sg13g2_fill_1 FILLER_50_1539 ();
 sg13g2_fill_2 FILLER_50_1552 ();
 sg13g2_fill_1 FILLER_50_1575 ();
 sg13g2_fill_2 FILLER_50_1605 ();
 sg13g2_fill_1 FILLER_50_1612 ();
 sg13g2_fill_2 FILLER_50_1650 ();
 sg13g2_decap_4 FILLER_50_1661 ();
 sg13g2_fill_1 FILLER_50_1665 ();
 sg13g2_fill_1 FILLER_50_1717 ();
 sg13g2_fill_1 FILLER_50_1799 ();
 sg13g2_fill_2 FILLER_50_1811 ();
 sg13g2_fill_2 FILLER_50_1827 ();
 sg13g2_fill_2 FILLER_50_1837 ();
 sg13g2_fill_1 FILLER_50_1844 ();
 sg13g2_fill_2 FILLER_50_1849 ();
 sg13g2_fill_2 FILLER_50_1869 ();
 sg13g2_fill_2 FILLER_50_1881 ();
 sg13g2_fill_1 FILLER_50_1888 ();
 sg13g2_fill_1 FILLER_50_1898 ();
 sg13g2_fill_1 FILLER_50_1913 ();
 sg13g2_fill_2 FILLER_50_1976 ();
 sg13g2_fill_1 FILLER_50_1982 ();
 sg13g2_fill_1 FILLER_50_1988 ();
 sg13g2_fill_2 FILLER_50_2002 ();
 sg13g2_fill_1 FILLER_50_2009 ();
 sg13g2_fill_1 FILLER_50_2062 ();
 sg13g2_decap_4 FILLER_50_2089 ();
 sg13g2_fill_2 FILLER_50_2097 ();
 sg13g2_decap_8 FILLER_50_2103 ();
 sg13g2_decap_8 FILLER_50_2110 ();
 sg13g2_fill_2 FILLER_50_2117 ();
 sg13g2_fill_1 FILLER_50_2119 ();
 sg13g2_fill_2 FILLER_50_2149 ();
 sg13g2_fill_1 FILLER_50_2151 ();
 sg13g2_fill_1 FILLER_50_2156 ();
 sg13g2_fill_2 FILLER_50_2163 ();
 sg13g2_fill_2 FILLER_50_2170 ();
 sg13g2_fill_2 FILLER_50_2194 ();
 sg13g2_decap_8 FILLER_50_2208 ();
 sg13g2_decap_8 FILLER_50_2215 ();
 sg13g2_decap_8 FILLER_50_2222 ();
 sg13g2_decap_8 FILLER_50_2229 ();
 sg13g2_decap_8 FILLER_50_2236 ();
 sg13g2_decap_4 FILLER_50_2243 ();
 sg13g2_fill_1 FILLER_50_2247 ();
 sg13g2_fill_1 FILLER_50_2252 ();
 sg13g2_decap_8 FILLER_50_2258 ();
 sg13g2_fill_1 FILLER_50_2282 ();
 sg13g2_fill_2 FILLER_50_2296 ();
 sg13g2_fill_1 FILLER_50_2303 ();
 sg13g2_decap_8 FILLER_50_2307 ();
 sg13g2_decap_4 FILLER_50_2314 ();
 sg13g2_fill_1 FILLER_50_2318 ();
 sg13g2_fill_1 FILLER_50_2328 ();
 sg13g2_fill_2 FILLER_50_2333 ();
 sg13g2_fill_1 FILLER_50_2349 ();
 sg13g2_fill_1 FILLER_50_2355 ();
 sg13g2_fill_1 FILLER_50_2376 ();
 sg13g2_fill_1 FILLER_50_2387 ();
 sg13g2_fill_1 FILLER_50_2398 ();
 sg13g2_fill_1 FILLER_50_2404 ();
 sg13g2_fill_1 FILLER_50_2414 ();
 sg13g2_fill_1 FILLER_50_2420 ();
 sg13g2_fill_2 FILLER_50_2428 ();
 sg13g2_fill_1 FILLER_50_2480 ();
 sg13g2_fill_2 FILLER_50_2486 ();
 sg13g2_fill_1 FILLER_50_2542 ();
 sg13g2_fill_2 FILLER_50_2558 ();
 sg13g2_fill_1 FILLER_50_2576 ();
 sg13g2_decap_8 FILLER_50_2595 ();
 sg13g2_decap_8 FILLER_50_2602 ();
 sg13g2_fill_2 FILLER_50_2609 ();
 sg13g2_fill_1 FILLER_50_2614 ();
 sg13g2_fill_2 FILLER_50_2620 ();
 sg13g2_fill_2 FILLER_50_2633 ();
 sg13g2_fill_1 FILLER_50_2635 ();
 sg13g2_decap_4 FILLER_50_2666 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_41 ();
 sg13g2_fill_1 FILLER_51_48 ();
 sg13g2_decap_8 FILLER_51_75 ();
 sg13g2_decap_4 FILLER_51_82 ();
 sg13g2_decap_4 FILLER_51_90 ();
 sg13g2_fill_2 FILLER_51_94 ();
 sg13g2_decap_8 FILLER_51_100 ();
 sg13g2_decap_8 FILLER_51_107 ();
 sg13g2_decap_4 FILLER_51_114 ();
 sg13g2_fill_2 FILLER_51_152 ();
 sg13g2_fill_2 FILLER_51_233 ();
 sg13g2_fill_1 FILLER_51_261 ();
 sg13g2_fill_1 FILLER_51_266 ();
 sg13g2_fill_2 FILLER_51_293 ();
 sg13g2_fill_1 FILLER_51_295 ();
 sg13g2_decap_4 FILLER_51_300 ();
 sg13g2_fill_1 FILLER_51_304 ();
 sg13g2_decap_8 FILLER_51_309 ();
 sg13g2_decap_8 FILLER_51_316 ();
 sg13g2_decap_8 FILLER_51_323 ();
 sg13g2_decap_8 FILLER_51_330 ();
 sg13g2_fill_2 FILLER_51_337 ();
 sg13g2_fill_1 FILLER_51_339 ();
 sg13g2_decap_4 FILLER_51_374 ();
 sg13g2_fill_2 FILLER_51_378 ();
 sg13g2_fill_2 FILLER_51_384 ();
 sg13g2_fill_2 FILLER_51_398 ();
 sg13g2_fill_1 FILLER_51_400 ();
 sg13g2_decap_8 FILLER_51_463 ();
 sg13g2_decap_8 FILLER_51_470 ();
 sg13g2_fill_2 FILLER_51_498 ();
 sg13g2_fill_1 FILLER_51_500 ();
 sg13g2_fill_2 FILLER_51_505 ();
 sg13g2_fill_1 FILLER_51_507 ();
 sg13g2_decap_8 FILLER_51_512 ();
 sg13g2_fill_1 FILLER_51_519 ();
 sg13g2_fill_2 FILLER_51_531 ();
 sg13g2_fill_2 FILLER_51_559 ();
 sg13g2_fill_1 FILLER_51_561 ();
 sg13g2_fill_2 FILLER_51_566 ();
 sg13g2_decap_4 FILLER_51_572 ();
 sg13g2_decap_8 FILLER_51_580 ();
 sg13g2_decap_4 FILLER_51_587 ();
 sg13g2_fill_2 FILLER_51_594 ();
 sg13g2_fill_1 FILLER_51_596 ();
 sg13g2_fill_2 FILLER_51_602 ();
 sg13g2_fill_1 FILLER_51_604 ();
 sg13g2_fill_1 FILLER_51_612 ();
 sg13g2_fill_1 FILLER_51_650 ();
 sg13g2_fill_2 FILLER_51_656 ();
 sg13g2_fill_1 FILLER_51_675 ();
 sg13g2_fill_2 FILLER_51_691 ();
 sg13g2_fill_1 FILLER_51_716 ();
 sg13g2_fill_1 FILLER_51_720 ();
 sg13g2_fill_1 FILLER_51_766 ();
 sg13g2_fill_2 FILLER_51_805 ();
 sg13g2_fill_1 FILLER_51_833 ();
 sg13g2_fill_2 FILLER_51_837 ();
 sg13g2_fill_1 FILLER_51_839 ();
 sg13g2_fill_1 FILLER_51_862 ();
 sg13g2_fill_1 FILLER_51_892 ();
 sg13g2_fill_2 FILLER_51_919 ();
 sg13g2_fill_2 FILLER_51_947 ();
 sg13g2_fill_2 FILLER_51_953 ();
 sg13g2_fill_1 FILLER_51_955 ();
 sg13g2_fill_1 FILLER_51_982 ();
 sg13g2_fill_1 FILLER_51_1015 ();
 sg13g2_fill_2 FILLER_51_1029 ();
 sg13g2_fill_1 FILLER_51_1038 ();
 sg13g2_fill_1 FILLER_51_1047 ();
 sg13g2_fill_2 FILLER_51_1123 ();
 sg13g2_fill_1 FILLER_51_1134 ();
 sg13g2_fill_1 FILLER_51_1182 ();
 sg13g2_fill_2 FILLER_51_1191 ();
 sg13g2_fill_2 FILLER_51_1202 ();
 sg13g2_fill_2 FILLER_51_1304 ();
 sg13g2_decap_8 FILLER_51_1318 ();
 sg13g2_decap_8 FILLER_51_1325 ();
 sg13g2_decap_8 FILLER_51_1332 ();
 sg13g2_decap_8 FILLER_51_1339 ();
 sg13g2_decap_8 FILLER_51_1346 ();
 sg13g2_decap_4 FILLER_51_1353 ();
 sg13g2_decap_4 FILLER_51_1362 ();
 sg13g2_fill_2 FILLER_51_1392 ();
 sg13g2_fill_1 FILLER_51_1403 ();
 sg13g2_fill_1 FILLER_51_1421 ();
 sg13g2_fill_1 FILLER_51_1430 ();
 sg13g2_decap_8 FILLER_51_1491 ();
 sg13g2_fill_2 FILLER_51_1498 ();
 sg13g2_fill_1 FILLER_51_1500 ();
 sg13g2_fill_2 FILLER_51_1539 ();
 sg13g2_fill_1 FILLER_51_1568 ();
 sg13g2_fill_2 FILLER_51_1583 ();
 sg13g2_fill_2 FILLER_51_1634 ();
 sg13g2_decap_8 FILLER_51_1640 ();
 sg13g2_decap_8 FILLER_51_1650 ();
 sg13g2_decap_8 FILLER_51_1657 ();
 sg13g2_decap_4 FILLER_51_1664 ();
 sg13g2_fill_1 FILLER_51_1668 ();
 sg13g2_fill_2 FILLER_51_1677 ();
 sg13g2_decap_8 FILLER_51_1687 ();
 sg13g2_fill_1 FILLER_51_1703 ();
 sg13g2_fill_2 FILLER_51_1720 ();
 sg13g2_fill_2 FILLER_51_1748 ();
 sg13g2_fill_1 FILLER_51_1775 ();
 sg13g2_fill_1 FILLER_51_1837 ();
 sg13g2_fill_1 FILLER_51_1870 ();
 sg13g2_fill_2 FILLER_51_1875 ();
 sg13g2_fill_1 FILLER_51_1922 ();
 sg13g2_fill_2 FILLER_51_1933 ();
 sg13g2_fill_1 FILLER_51_1967 ();
 sg13g2_fill_1 FILLER_51_1997 ();
 sg13g2_fill_1 FILLER_51_2013 ();
 sg13g2_fill_2 FILLER_51_2021 ();
 sg13g2_fill_2 FILLER_51_2083 ();
 sg13g2_fill_2 FILLER_51_2098 ();
 sg13g2_decap_8 FILLER_51_2111 ();
 sg13g2_decap_8 FILLER_51_2118 ();
 sg13g2_decap_8 FILLER_51_2125 ();
 sg13g2_decap_4 FILLER_51_2132 ();
 sg13g2_fill_2 FILLER_51_2156 ();
 sg13g2_fill_2 FILLER_51_2167 ();
 sg13g2_fill_2 FILLER_51_2182 ();
 sg13g2_decap_8 FILLER_51_2201 ();
 sg13g2_fill_2 FILLER_51_2208 ();
 sg13g2_fill_2 FILLER_51_2214 ();
 sg13g2_fill_1 FILLER_51_2216 ();
 sg13g2_decap_8 FILLER_51_2221 ();
 sg13g2_decap_4 FILLER_51_2228 ();
 sg13g2_fill_1 FILLER_51_2232 ();
 sg13g2_decap_4 FILLER_51_2264 ();
 sg13g2_fill_1 FILLER_51_2272 ();
 sg13g2_decap_4 FILLER_51_2278 ();
 sg13g2_decap_8 FILLER_51_2316 ();
 sg13g2_fill_2 FILLER_51_2323 ();
 sg13g2_decap_8 FILLER_51_2341 ();
 sg13g2_fill_1 FILLER_51_2348 ();
 sg13g2_fill_1 FILLER_51_2354 ();
 sg13g2_fill_2 FILLER_51_2359 ();
 sg13g2_fill_1 FILLER_51_2361 ();
 sg13g2_fill_1 FILLER_51_2366 ();
 sg13g2_fill_2 FILLER_51_2371 ();
 sg13g2_decap_4 FILLER_51_2378 ();
 sg13g2_decap_8 FILLER_51_2394 ();
 sg13g2_fill_2 FILLER_51_2401 ();
 sg13g2_fill_1 FILLER_51_2403 ();
 sg13g2_fill_2 FILLER_51_2409 ();
 sg13g2_fill_2 FILLER_51_2414 ();
 sg13g2_fill_2 FILLER_51_2442 ();
 sg13g2_decap_4 FILLER_51_2457 ();
 sg13g2_fill_1 FILLER_51_2461 ();
 sg13g2_fill_2 FILLER_51_2466 ();
 sg13g2_fill_1 FILLER_51_2468 ();
 sg13g2_fill_1 FILLER_51_2528 ();
 sg13g2_fill_1 FILLER_51_2569 ();
 sg13g2_decap_4 FILLER_51_2578 ();
 sg13g2_decap_8 FILLER_51_2587 ();
 sg13g2_decap_8 FILLER_51_2599 ();
 sg13g2_fill_2 FILLER_51_2606 ();
 sg13g2_fill_1 FILLER_51_2608 ();
 sg13g2_decap_4 FILLER_51_2614 ();
 sg13g2_fill_2 FILLER_51_2618 ();
 sg13g2_fill_1 FILLER_51_2626 ();
 sg13g2_decap_4 FILLER_51_2632 ();
 sg13g2_fill_2 FILLER_51_2636 ();
 sg13g2_decap_4 FILLER_51_2664 ();
 sg13g2_fill_2 FILLER_51_2668 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_13 ();
 sg13g2_fill_1 FILLER_52_19 ();
 sg13g2_fill_2 FILLER_52_25 ();
 sg13g2_fill_2 FILLER_52_48 ();
 sg13g2_fill_1 FILLER_52_59 ();
 sg13g2_fill_1 FILLER_52_64 ();
 sg13g2_fill_1 FILLER_52_70 ();
 sg13g2_decap_4 FILLER_52_75 ();
 sg13g2_fill_2 FILLER_52_79 ();
 sg13g2_fill_1 FILLER_52_129 ();
 sg13g2_decap_4 FILLER_52_138 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_decap_4 FILLER_52_148 ();
 sg13g2_fill_1 FILLER_52_152 ();
 sg13g2_fill_2 FILLER_52_183 ();
 sg13g2_fill_1 FILLER_52_204 ();
 sg13g2_fill_1 FILLER_52_210 ();
 sg13g2_decap_4 FILLER_52_267 ();
 sg13g2_fill_1 FILLER_52_275 ();
 sg13g2_fill_2 FILLER_52_280 ();
 sg13g2_fill_1 FILLER_52_282 ();
 sg13g2_fill_2 FILLER_52_335 ();
 sg13g2_fill_1 FILLER_52_337 ();
 sg13g2_fill_2 FILLER_52_368 ();
 sg13g2_fill_1 FILLER_52_370 ();
 sg13g2_fill_2 FILLER_52_388 ();
 sg13g2_fill_2 FILLER_52_395 ();
 sg13g2_decap_4 FILLER_52_432 ();
 sg13g2_decap_8 FILLER_52_452 ();
 sg13g2_decap_8 FILLER_52_459 ();
 sg13g2_fill_1 FILLER_52_466 ();
 sg13g2_fill_2 FILLER_52_480 ();
 sg13g2_fill_2 FILLER_52_530 ();
 sg13g2_fill_1 FILLER_52_532 ();
 sg13g2_fill_2 FILLER_52_585 ();
 sg13g2_fill_1 FILLER_52_640 ();
 sg13g2_fill_1 FILLER_52_695 ();
 sg13g2_fill_2 FILLER_52_722 ();
 sg13g2_fill_2 FILLER_52_755 ();
 sg13g2_fill_1 FILLER_52_777 ();
 sg13g2_fill_2 FILLER_52_818 ();
 sg13g2_fill_1 FILLER_52_833 ();
 sg13g2_decap_4 FILLER_52_844 ();
 sg13g2_fill_1 FILLER_52_852 ();
 sg13g2_decap_4 FILLER_52_876 ();
 sg13g2_fill_2 FILLER_52_915 ();
 sg13g2_fill_1 FILLER_52_917 ();
 sg13g2_fill_1 FILLER_52_923 ();
 sg13g2_decap_8 FILLER_52_933 ();
 sg13g2_decap_8 FILLER_52_940 ();
 sg13g2_decap_4 FILLER_52_947 ();
 sg13g2_decap_4 FILLER_52_976 ();
 sg13g2_fill_1 FILLER_52_980 ();
 sg13g2_fill_2 FILLER_52_997 ();
 sg13g2_fill_1 FILLER_52_1100 ();
 sg13g2_fill_1 FILLER_52_1121 ();
 sg13g2_fill_2 FILLER_52_1132 ();
 sg13g2_fill_1 FILLER_52_1142 ();
 sg13g2_fill_2 FILLER_52_1161 ();
 sg13g2_fill_2 FILLER_52_1193 ();
 sg13g2_fill_1 FILLER_52_1201 ();
 sg13g2_fill_2 FILLER_52_1207 ();
 sg13g2_fill_1 FILLER_52_1242 ();
 sg13g2_fill_2 FILLER_52_1325 ();
 sg13g2_fill_2 FILLER_52_1353 ();
 sg13g2_fill_1 FILLER_52_1355 ();
 sg13g2_fill_2 FILLER_52_1382 ();
 sg13g2_fill_1 FILLER_52_1384 ();
 sg13g2_fill_2 FILLER_52_1389 ();
 sg13g2_fill_1 FILLER_52_1396 ();
 sg13g2_decap_4 FILLER_52_1406 ();
 sg13g2_fill_1 FILLER_52_1410 ();
 sg13g2_fill_1 FILLER_52_1436 ();
 sg13g2_fill_1 FILLER_52_1471 ();
 sg13g2_fill_2 FILLER_52_1475 ();
 sg13g2_decap_4 FILLER_52_1483 ();
 sg13g2_fill_1 FILLER_52_1563 ();
 sg13g2_fill_1 FILLER_52_1596 ();
 sg13g2_fill_1 FILLER_52_1610 ();
 sg13g2_fill_2 FILLER_52_1678 ();
 sg13g2_fill_2 FILLER_52_1701 ();
 sg13g2_fill_2 FILLER_52_1743 ();
 sg13g2_fill_1 FILLER_52_1761 ();
 sg13g2_fill_1 FILLER_52_1823 ();
 sg13g2_fill_1 FILLER_52_1862 ();
 sg13g2_fill_2 FILLER_52_1889 ();
 sg13g2_fill_1 FILLER_52_1920 ();
 sg13g2_fill_1 FILLER_52_1957 ();
 sg13g2_fill_1 FILLER_52_1972 ();
 sg13g2_fill_1 FILLER_52_1989 ();
 sg13g2_fill_2 FILLER_52_1994 ();
 sg13g2_fill_2 FILLER_52_2000 ();
 sg13g2_fill_2 FILLER_52_2006 ();
 sg13g2_fill_1 FILLER_52_2012 ();
 sg13g2_fill_2 FILLER_52_2039 ();
 sg13g2_fill_2 FILLER_52_2051 ();
 sg13g2_fill_1 FILLER_52_2060 ();
 sg13g2_fill_2 FILLER_52_2076 ();
 sg13g2_fill_1 FILLER_52_2092 ();
 sg13g2_decap_4 FILLER_52_2129 ();
 sg13g2_fill_1 FILLER_52_2133 ();
 sg13g2_fill_1 FILLER_52_2139 ();
 sg13g2_fill_2 FILLER_52_2150 ();
 sg13g2_fill_2 FILLER_52_2156 ();
 sg13g2_decap_4 FILLER_52_2162 ();
 sg13g2_fill_2 FILLER_52_2166 ();
 sg13g2_fill_2 FILLER_52_2177 ();
 sg13g2_fill_1 FILLER_52_2179 ();
 sg13g2_decap_8 FILLER_52_2198 ();
 sg13g2_decap_4 FILLER_52_2205 ();
 sg13g2_fill_2 FILLER_52_2209 ();
 sg13g2_decap_4 FILLER_52_2216 ();
 sg13g2_fill_1 FILLER_52_2224 ();
 sg13g2_fill_1 FILLER_52_2245 ();
 sg13g2_fill_2 FILLER_52_2250 ();
 sg13g2_decap_8 FILLER_52_2256 ();
 sg13g2_decap_8 FILLER_52_2263 ();
 sg13g2_decap_8 FILLER_52_2270 ();
 sg13g2_decap_4 FILLER_52_2277 ();
 sg13g2_fill_2 FILLER_52_2309 ();
 sg13g2_fill_2 FILLER_52_2316 ();
 sg13g2_fill_1 FILLER_52_2318 ();
 sg13g2_fill_1 FILLER_52_2345 ();
 sg13g2_decap_4 FILLER_52_2351 ();
 sg13g2_fill_1 FILLER_52_2355 ();
 sg13g2_fill_2 FILLER_52_2366 ();
 sg13g2_decap_8 FILLER_52_2374 ();
 sg13g2_decap_8 FILLER_52_2381 ();
 sg13g2_fill_1 FILLER_52_2388 ();
 sg13g2_decap_8 FILLER_52_2397 ();
 sg13g2_fill_1 FILLER_52_2404 ();
 sg13g2_fill_1 FILLER_52_2413 ();
 sg13g2_decap_8 FILLER_52_2450 ();
 sg13g2_decap_4 FILLER_52_2462 ();
 sg13g2_fill_2 FILLER_52_2466 ();
 sg13g2_decap_8 FILLER_52_2473 ();
 sg13g2_fill_2 FILLER_52_2480 ();
 sg13g2_fill_1 FILLER_52_2482 ();
 sg13g2_decap_4 FILLER_52_2487 ();
 sg13g2_fill_1 FILLER_52_2491 ();
 sg13g2_decap_4 FILLER_52_2522 ();
 sg13g2_fill_2 FILLER_52_2544 ();
 sg13g2_fill_1 FILLER_52_2579 ();
 sg13g2_fill_1 FILLER_52_2586 ();
 sg13g2_fill_1 FILLER_52_2592 ();
 sg13g2_fill_2 FILLER_52_2619 ();
 sg13g2_fill_1 FILLER_52_2632 ();
 sg13g2_decap_8 FILLER_52_2659 ();
 sg13g2_decap_4 FILLER_52_2666 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_14 ();
 sg13g2_decap_4 FILLER_53_39 ();
 sg13g2_fill_1 FILLER_53_52 ();
 sg13g2_fill_2 FILLER_53_83 ();
 sg13g2_fill_1 FILLER_53_89 ();
 sg13g2_decap_4 FILLER_53_116 ();
 sg13g2_fill_2 FILLER_53_120 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_fill_2 FILLER_53_140 ();
 sg13g2_fill_1 FILLER_53_142 ();
 sg13g2_fill_2 FILLER_53_164 ();
 sg13g2_fill_1 FILLER_53_186 ();
 sg13g2_fill_2 FILLER_53_228 ();
 sg13g2_fill_1 FILLER_53_241 ();
 sg13g2_fill_1 FILLER_53_246 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_decap_4 FILLER_53_296 ();
 sg13g2_fill_1 FILLER_53_300 ();
 sg13g2_decap_4 FILLER_53_305 ();
 sg13g2_fill_2 FILLER_53_309 ();
 sg13g2_decap_8 FILLER_53_419 ();
 sg13g2_decap_4 FILLER_53_426 ();
 sg13g2_fill_2 FILLER_53_438 ();
 sg13g2_fill_1 FILLER_53_440 ();
 sg13g2_decap_4 FILLER_53_447 ();
 sg13g2_fill_2 FILLER_53_451 ();
 sg13g2_fill_1 FILLER_53_476 ();
 sg13g2_fill_2 FILLER_53_481 ();
 sg13g2_fill_1 FILLER_53_483 ();
 sg13g2_fill_1 FILLER_53_515 ();
 sg13g2_fill_2 FILLER_53_537 ();
 sg13g2_fill_1 FILLER_53_542 ();
 sg13g2_fill_2 FILLER_53_555 ();
 sg13g2_fill_2 FILLER_53_570 ();
 sg13g2_fill_1 FILLER_53_572 ();
 sg13g2_fill_1 FILLER_53_612 ();
 sg13g2_fill_1 FILLER_53_773 ();
 sg13g2_fill_2 FILLER_53_790 ();
 sg13g2_fill_1 FILLER_53_855 ();
 sg13g2_fill_2 FILLER_53_892 ();
 sg13g2_fill_2 FILLER_53_899 ();
 sg13g2_decap_8 FILLER_53_923 ();
 sg13g2_decap_8 FILLER_53_930 ();
 sg13g2_decap_4 FILLER_53_937 ();
 sg13g2_fill_1 FILLER_53_941 ();
 sg13g2_fill_2 FILLER_53_981 ();
 sg13g2_fill_1 FILLER_53_1053 ();
 sg13g2_fill_1 FILLER_53_1085 ();
 sg13g2_fill_1 FILLER_53_1112 ();
 sg13g2_fill_1 FILLER_53_1123 ();
 sg13g2_fill_1 FILLER_53_1155 ();
 sg13g2_fill_2 FILLER_53_1193 ();
 sg13g2_fill_2 FILLER_53_1218 ();
 sg13g2_fill_2 FILLER_53_1249 ();
 sg13g2_fill_2 FILLER_53_1259 ();
 sg13g2_fill_2 FILLER_53_1280 ();
 sg13g2_fill_2 FILLER_53_1311 ();
 sg13g2_fill_2 FILLER_53_1319 ();
 sg13g2_fill_2 FILLER_53_1354 ();
 sg13g2_fill_1 FILLER_53_1386 ();
 sg13g2_fill_2 FILLER_53_1392 ();
 sg13g2_fill_1 FILLER_53_1398 ();
 sg13g2_fill_2 FILLER_53_1492 ();
 sg13g2_fill_2 FILLER_53_1507 ();
 sg13g2_fill_1 FILLER_53_1519 ();
 sg13g2_fill_2 FILLER_53_1550 ();
 sg13g2_fill_2 FILLER_53_1561 ();
 sg13g2_fill_1 FILLER_53_1574 ();
 sg13g2_fill_1 FILLER_53_1616 ();
 sg13g2_fill_1 FILLER_53_1643 ();
 sg13g2_fill_1 FILLER_53_1676 ();
 sg13g2_fill_1 FILLER_53_1718 ();
 sg13g2_fill_1 FILLER_53_1728 ();
 sg13g2_fill_1 FILLER_53_1761 ();
 sg13g2_fill_2 FILLER_53_1774 ();
 sg13g2_fill_2 FILLER_53_1784 ();
 sg13g2_fill_2 FILLER_53_1794 ();
 sg13g2_fill_1 FILLER_53_1906 ();
 sg13g2_fill_1 FILLER_53_1972 ();
 sg13g2_decap_8 FILLER_53_2025 ();
 sg13g2_decap_4 FILLER_53_2036 ();
 sg13g2_fill_2 FILLER_53_2040 ();
 sg13g2_fill_1 FILLER_53_2052 ();
 sg13g2_fill_1 FILLER_53_2068 ();
 sg13g2_fill_2 FILLER_53_2082 ();
 sg13g2_fill_2 FILLER_53_2095 ();
 sg13g2_decap_4 FILLER_53_2135 ();
 sg13g2_decap_4 FILLER_53_2143 ();
 sg13g2_fill_1 FILLER_53_2147 ();
 sg13g2_fill_1 FILLER_53_2167 ();
 sg13g2_fill_1 FILLER_53_2172 ();
 sg13g2_decap_4 FILLER_53_2182 ();
 sg13g2_fill_1 FILLER_53_2186 ();
 sg13g2_decap_4 FILLER_53_2196 ();
 sg13g2_fill_1 FILLER_53_2200 ();
 sg13g2_fill_1 FILLER_53_2216 ();
 sg13g2_fill_2 FILLER_53_2227 ();
 sg13g2_fill_1 FILLER_53_2245 ();
 sg13g2_decap_8 FILLER_53_2267 ();
 sg13g2_decap_8 FILLER_53_2274 ();
 sg13g2_fill_2 FILLER_53_2281 ();
 sg13g2_fill_2 FILLER_53_2292 ();
 sg13g2_fill_2 FILLER_53_2298 ();
 sg13g2_fill_1 FILLER_53_2300 ();
 sg13g2_fill_1 FILLER_53_2315 ();
 sg13g2_fill_1 FILLER_53_2326 ();
 sg13g2_fill_2 FILLER_53_2338 ();
 sg13g2_decap_8 FILLER_53_2350 ();
 sg13g2_decap_8 FILLER_53_2357 ();
 sg13g2_fill_1 FILLER_53_2364 ();
 sg13g2_fill_1 FILLER_53_2369 ();
 sg13g2_decap_8 FILLER_53_2374 ();
 sg13g2_decap_8 FILLER_53_2381 ();
 sg13g2_decap_8 FILLER_53_2388 ();
 sg13g2_decap_8 FILLER_53_2395 ();
 sg13g2_decap_4 FILLER_53_2402 ();
 sg13g2_fill_1 FILLER_53_2406 ();
 sg13g2_fill_1 FILLER_53_2422 ();
 sg13g2_fill_2 FILLER_53_2428 ();
 sg13g2_fill_1 FILLER_53_2434 ();
 sg13g2_fill_2 FILLER_53_2440 ();
 sg13g2_decap_8 FILLER_53_2477 ();
 sg13g2_decap_8 FILLER_53_2484 ();
 sg13g2_decap_4 FILLER_53_2491 ();
 sg13g2_fill_2 FILLER_53_2495 ();
 sg13g2_fill_2 FILLER_53_2521 ();
 sg13g2_fill_1 FILLER_53_2523 ();
 sg13g2_fill_2 FILLER_53_2530 ();
 sg13g2_fill_1 FILLER_53_2543 ();
 sg13g2_fill_1 FILLER_53_2552 ();
 sg13g2_fill_1 FILLER_53_2566 ();
 sg13g2_fill_1 FILLER_53_2608 ();
 sg13g2_fill_2 FILLER_53_2667 ();
 sg13g2_fill_1 FILLER_53_2669 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_74 ();
 sg13g2_fill_2 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_decap_8 FILLER_54_122 ();
 sg13g2_fill_2 FILLER_54_129 ();
 sg13g2_fill_1 FILLER_54_131 ();
 sg13g2_fill_1 FILLER_54_167 ();
 sg13g2_fill_1 FILLER_54_196 ();
 sg13g2_fill_1 FILLER_54_214 ();
 sg13g2_fill_1 FILLER_54_223 ();
 sg13g2_fill_1 FILLER_54_269 ();
 sg13g2_decap_4 FILLER_54_318 ();
 sg13g2_fill_1 FILLER_54_327 ();
 sg13g2_fill_2 FILLER_54_332 ();
 sg13g2_fill_1 FILLER_54_338 ();
 sg13g2_fill_1 FILLER_54_368 ();
 sg13g2_fill_1 FILLER_54_389 ();
 sg13g2_fill_2 FILLER_54_395 ();
 sg13g2_fill_1 FILLER_54_397 ();
 sg13g2_fill_2 FILLER_54_428 ();
 sg13g2_fill_2 FILLER_54_461 ();
 sg13g2_fill_1 FILLER_54_463 ();
 sg13g2_fill_1 FILLER_54_530 ();
 sg13g2_fill_2 FILLER_54_561 ();
 sg13g2_fill_1 FILLER_54_563 ();
 sg13g2_fill_2 FILLER_54_569 ();
 sg13g2_fill_2 FILLER_54_576 ();
 sg13g2_fill_2 FILLER_54_664 ();
 sg13g2_fill_1 FILLER_54_696 ();
 sg13g2_fill_2 FILLER_54_711 ();
 sg13g2_fill_1 FILLER_54_742 ();
 sg13g2_fill_1 FILLER_54_791 ();
 sg13g2_fill_2 FILLER_54_830 ();
 sg13g2_fill_1 FILLER_54_984 ();
 sg13g2_fill_1 FILLER_54_1004 ();
 sg13g2_fill_1 FILLER_54_1009 ();
 sg13g2_fill_2 FILLER_54_1069 ();
 sg13g2_fill_1 FILLER_54_1075 ();
 sg13g2_fill_2 FILLER_54_1174 ();
 sg13g2_fill_1 FILLER_54_1192 ();
 sg13g2_fill_2 FILLER_54_1265 ();
 sg13g2_fill_1 FILLER_54_1275 ();
 sg13g2_fill_2 FILLER_54_1371 ();
 sg13g2_fill_1 FILLER_54_1373 ();
 sg13g2_fill_1 FILLER_54_1400 ();
 sg13g2_fill_1 FILLER_54_1440 ();
 sg13g2_fill_2 FILLER_54_1458 ();
 sg13g2_fill_1 FILLER_54_1470 ();
 sg13g2_fill_2 FILLER_54_1504 ();
 sg13g2_fill_1 FILLER_54_1575 ();
 sg13g2_fill_1 FILLER_54_1606 ();
 sg13g2_fill_2 FILLER_54_1656 ();
 sg13g2_fill_1 FILLER_54_1710 ();
 sg13g2_fill_2 FILLER_54_1766 ();
 sg13g2_fill_2 FILLER_54_1818 ();
 sg13g2_fill_2 FILLER_54_1838 ();
 sg13g2_fill_1 FILLER_54_1866 ();
 sg13g2_fill_2 FILLER_54_1910 ();
 sg13g2_fill_1 FILLER_54_1919 ();
 sg13g2_fill_1 FILLER_54_1928 ();
 sg13g2_fill_1 FILLER_54_1949 ();
 sg13g2_fill_1 FILLER_54_1968 ();
 sg13g2_decap_4 FILLER_54_2029 ();
 sg13g2_fill_1 FILLER_54_2038 ();
 sg13g2_fill_1 FILLER_54_2068 ();
 sg13g2_fill_2 FILLER_54_2073 ();
 sg13g2_fill_1 FILLER_54_2167 ();
 sg13g2_fill_1 FILLER_54_2173 ();
 sg13g2_fill_2 FILLER_54_2215 ();
 sg13g2_fill_1 FILLER_54_2217 ();
 sg13g2_fill_2 FILLER_54_2279 ();
 sg13g2_decap_4 FILLER_54_2286 ();
 sg13g2_fill_1 FILLER_54_2312 ();
 sg13g2_decap_8 FILLER_54_2370 ();
 sg13g2_decap_8 FILLER_54_2381 ();
 sg13g2_fill_1 FILLER_54_2413 ();
 sg13g2_fill_1 FILLER_54_2428 ();
 sg13g2_fill_2 FILLER_54_2433 ();
 sg13g2_fill_1 FILLER_54_2435 ();
 sg13g2_fill_1 FILLER_54_2442 ();
 sg13g2_fill_1 FILLER_54_2453 ();
 sg13g2_fill_1 FILLER_54_2464 ();
 sg13g2_decap_4 FILLER_54_2473 ();
 sg13g2_fill_1 FILLER_54_2477 ();
 sg13g2_decap_8 FILLER_54_2496 ();
 sg13g2_decap_4 FILLER_54_2503 ();
 sg13g2_fill_2 FILLER_54_2507 ();
 sg13g2_fill_2 FILLER_54_2540 ();
 sg13g2_fill_1 FILLER_54_2556 ();
 sg13g2_fill_1 FILLER_54_2602 ();
 sg13g2_fill_1 FILLER_54_2607 ();
 sg13g2_fill_1 FILLER_54_2614 ();
 sg13g2_decap_8 FILLER_54_2661 ();
 sg13g2_fill_2 FILLER_54_2668 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_34 ();
 sg13g2_fill_2 FILLER_55_39 ();
 sg13g2_fill_1 FILLER_55_41 ();
 sg13g2_fill_1 FILLER_55_50 ();
 sg13g2_fill_2 FILLER_55_60 ();
 sg13g2_fill_1 FILLER_55_62 ();
 sg13g2_decap_8 FILLER_55_115 ();
 sg13g2_fill_1 FILLER_55_122 ();
 sg13g2_fill_1 FILLER_55_162 ();
 sg13g2_fill_2 FILLER_55_210 ();
 sg13g2_fill_1 FILLER_55_238 ();
 sg13g2_fill_1 FILLER_55_294 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_309 ();
 sg13g2_decap_8 FILLER_55_319 ();
 sg13g2_fill_2 FILLER_55_326 ();
 sg13g2_fill_1 FILLER_55_328 ();
 sg13g2_fill_2 FILLER_55_333 ();
 sg13g2_decap_8 FILLER_55_339 ();
 sg13g2_fill_2 FILLER_55_377 ();
 sg13g2_fill_1 FILLER_55_403 ();
 sg13g2_fill_1 FILLER_55_476 ();
 sg13g2_fill_1 FILLER_55_483 ();
 sg13g2_fill_1 FILLER_55_505 ();
 sg13g2_fill_2 FILLER_55_518 ();
 sg13g2_fill_2 FILLER_55_568 ();
 sg13g2_fill_2 FILLER_55_616 ();
 sg13g2_fill_1 FILLER_55_633 ();
 sg13g2_fill_2 FILLER_55_673 ();
 sg13g2_fill_2 FILLER_55_683 ();
 sg13g2_fill_1 FILLER_55_693 ();
 sg13g2_fill_1 FILLER_55_698 ();
 sg13g2_fill_1 FILLER_55_709 ();
 sg13g2_fill_1 FILLER_55_804 ();
 sg13g2_fill_1 FILLER_55_809 ();
 sg13g2_fill_1 FILLER_55_849 ();
 sg13g2_decap_4 FILLER_55_854 ();
 sg13g2_fill_1 FILLER_55_858 ();
 sg13g2_fill_1 FILLER_55_875 ();
 sg13g2_fill_2 FILLER_55_900 ();
 sg13g2_fill_1 FILLER_55_906 ();
 sg13g2_fill_2 FILLER_55_946 ();
 sg13g2_fill_1 FILLER_55_963 ();
 sg13g2_fill_1 FILLER_55_992 ();
 sg13g2_fill_2 FILLER_55_1045 ();
 sg13g2_fill_1 FILLER_55_1052 ();
 sg13g2_fill_2 FILLER_55_1081 ();
 sg13g2_fill_1 FILLER_55_1087 ();
 sg13g2_fill_2 FILLER_55_1109 ();
 sg13g2_fill_2 FILLER_55_1170 ();
 sg13g2_fill_1 FILLER_55_1190 ();
 sg13g2_fill_2 FILLER_55_1222 ();
 sg13g2_fill_2 FILLER_55_1274 ();
 sg13g2_fill_1 FILLER_55_1286 ();
 sg13g2_fill_1 FILLER_55_1290 ();
 sg13g2_fill_2 FILLER_55_1327 ();
 sg13g2_fill_1 FILLER_55_1352 ();
 sg13g2_decap_8 FILLER_55_1366 ();
 sg13g2_decap_4 FILLER_55_1373 ();
 sg13g2_fill_1 FILLER_55_1377 ();
 sg13g2_fill_2 FILLER_55_1416 ();
 sg13g2_fill_2 FILLER_55_1426 ();
 sg13g2_fill_1 FILLER_55_1428 ();
 sg13g2_fill_2 FILLER_55_1455 ();
 sg13g2_fill_1 FILLER_55_1457 ();
 sg13g2_fill_1 FILLER_55_1603 ();
 sg13g2_fill_1 FILLER_55_1614 ();
 sg13g2_fill_1 FILLER_55_1641 ();
 sg13g2_fill_1 FILLER_55_1662 ();
 sg13g2_fill_1 FILLER_55_1698 ();
 sg13g2_fill_2 FILLER_55_1802 ();
 sg13g2_decap_8 FILLER_55_1862 ();
 sg13g2_fill_2 FILLER_55_1889 ();
 sg13g2_fill_2 FILLER_55_1964 ();
 sg13g2_fill_1 FILLER_55_1988 ();
 sg13g2_fill_1 FILLER_55_2015 ();
 sg13g2_fill_2 FILLER_55_2020 ();
 sg13g2_fill_1 FILLER_55_2078 ();
 sg13g2_fill_1 FILLER_55_2103 ();
 sg13g2_fill_1 FILLER_55_2128 ();
 sg13g2_fill_2 FILLER_55_2133 ();
 sg13g2_fill_1 FILLER_55_2156 ();
 sg13g2_fill_1 FILLER_55_2162 ();
 sg13g2_fill_2 FILLER_55_2167 ();
 sg13g2_fill_1 FILLER_55_2169 ();
 sg13g2_fill_2 FILLER_55_2179 ();
 sg13g2_fill_1 FILLER_55_2185 ();
 sg13g2_decap_4 FILLER_55_2198 ();
 sg13g2_fill_1 FILLER_55_2207 ();
 sg13g2_fill_1 FILLER_55_2212 ();
 sg13g2_fill_1 FILLER_55_2220 ();
 sg13g2_fill_1 FILLER_55_2226 ();
 sg13g2_fill_2 FILLER_55_2245 ();
 sg13g2_fill_1 FILLER_55_2247 ();
 sg13g2_fill_2 FILLER_55_2253 ();
 sg13g2_fill_1 FILLER_55_2255 ();
 sg13g2_fill_2 FILLER_55_2271 ();
 sg13g2_fill_1 FILLER_55_2313 ();
 sg13g2_fill_1 FILLER_55_2340 ();
 sg13g2_fill_2 FILLER_55_2349 ();
 sg13g2_fill_2 FILLER_55_2355 ();
 sg13g2_fill_2 FILLER_55_2367 ();
 sg13g2_fill_1 FILLER_55_2373 ();
 sg13g2_fill_1 FILLER_55_2405 ();
 sg13g2_fill_1 FILLER_55_2436 ();
 sg13g2_fill_1 FILLER_55_2442 ();
 sg13g2_fill_1 FILLER_55_2454 ();
 sg13g2_fill_1 FILLER_55_2469 ();
 sg13g2_fill_1 FILLER_55_2482 ();
 sg13g2_fill_1 FILLER_55_2535 ();
 sg13g2_fill_2 FILLER_55_2544 ();
 sg13g2_fill_1 FILLER_55_2565 ();
 sg13g2_fill_2 FILLER_55_2578 ();
 sg13g2_decap_8 FILLER_55_2585 ();
 sg13g2_decap_8 FILLER_55_2592 ();
 sg13g2_fill_1 FILLER_55_2599 ();
 sg13g2_fill_2 FILLER_55_2646 ();
 sg13g2_decap_8 FILLER_55_2652 ();
 sg13g2_decap_8 FILLER_55_2659 ();
 sg13g2_decap_4 FILLER_55_2666 ();
 sg13g2_fill_2 FILLER_56_35 ();
 sg13g2_fill_2 FILLER_56_46 ();
 sg13g2_fill_1 FILLER_56_48 ();
 sg13g2_fill_1 FILLER_56_80 ();
 sg13g2_fill_1 FILLER_56_85 ();
 sg13g2_fill_2 FILLER_56_112 ();
 sg13g2_fill_1 FILLER_56_118 ();
 sg13g2_decap_4 FILLER_56_154 ();
 sg13g2_fill_1 FILLER_56_158 ();
 sg13g2_decap_8 FILLER_56_163 ();
 sg13g2_fill_1 FILLER_56_170 ();
 sg13g2_fill_1 FILLER_56_197 ();
 sg13g2_fill_1 FILLER_56_204 ();
 sg13g2_fill_1 FILLER_56_282 ();
 sg13g2_fill_2 FILLER_56_287 ();
 sg13g2_fill_2 FILLER_56_293 ();
 sg13g2_fill_2 FILLER_56_299 ();
 sg13g2_fill_1 FILLER_56_305 ();
 sg13g2_decap_4 FILLER_56_332 ();
 sg13g2_fill_2 FILLER_56_336 ();
 sg13g2_fill_1 FILLER_56_364 ();
 sg13g2_fill_1 FILLER_56_369 ();
 sg13g2_fill_2 FILLER_56_507 ();
 sg13g2_fill_1 FILLER_56_509 ();
 sg13g2_fill_1 FILLER_56_534 ();
 sg13g2_fill_1 FILLER_56_574 ();
 sg13g2_fill_1 FILLER_56_604 ();
 sg13g2_fill_2 FILLER_56_616 ();
 sg13g2_fill_1 FILLER_56_671 ();
 sg13g2_fill_2 FILLER_56_679 ();
 sg13g2_fill_1 FILLER_56_690 ();
 sg13g2_fill_2 FILLER_56_695 ();
 sg13g2_fill_1 FILLER_56_710 ();
 sg13g2_fill_1 FILLER_56_748 ();
 sg13g2_fill_1 FILLER_56_775 ();
 sg13g2_fill_2 FILLER_56_829 ();
 sg13g2_decap_4 FILLER_56_835 ();
 sg13g2_fill_2 FILLER_56_839 ();
 sg13g2_decap_8 FILLER_56_870 ();
 sg13g2_fill_2 FILLER_56_877 ();
 sg13g2_fill_1 FILLER_56_879 ();
 sg13g2_fill_2 FILLER_56_884 ();
 sg13g2_decap_8 FILLER_56_890 ();
 sg13g2_fill_2 FILLER_56_902 ();
 sg13g2_fill_1 FILLER_56_904 ();
 sg13g2_fill_1 FILLER_56_956 ();
 sg13g2_fill_1 FILLER_56_977 ();
 sg13g2_fill_1 FILLER_56_995 ();
 sg13g2_fill_2 FILLER_56_1001 ();
 sg13g2_fill_1 FILLER_56_1077 ();
 sg13g2_fill_2 FILLER_56_1095 ();
 sg13g2_fill_1 FILLER_56_1104 ();
 sg13g2_fill_1 FILLER_56_1108 ();
 sg13g2_fill_2 FILLER_56_1136 ();
 sg13g2_fill_1 FILLER_56_1232 ();
 sg13g2_fill_2 FILLER_56_1262 ();
 sg13g2_decap_8 FILLER_56_1380 ();
 sg13g2_fill_2 FILLER_56_1387 ();
 sg13g2_fill_1 FILLER_56_1389 ();
 sg13g2_decap_4 FILLER_56_1398 ();
 sg13g2_fill_1 FILLER_56_1402 ();
 sg13g2_fill_2 FILLER_56_1438 ();
 sg13g2_fill_1 FILLER_56_1519 ();
 sg13g2_fill_2 FILLER_56_1525 ();
 sg13g2_fill_1 FILLER_56_1553 ();
 sg13g2_fill_1 FILLER_56_1558 ();
 sg13g2_fill_1 FILLER_56_1563 ();
 sg13g2_fill_1 FILLER_56_1572 ();
 sg13g2_fill_1 FILLER_56_1603 ();
 sg13g2_fill_2 FILLER_56_1665 ();
 sg13g2_fill_2 FILLER_56_1679 ();
 sg13g2_fill_2 FILLER_56_1693 ();
 sg13g2_fill_2 FILLER_56_1711 ();
 sg13g2_fill_2 FILLER_56_1724 ();
 sg13g2_fill_2 FILLER_56_1748 ();
 sg13g2_fill_1 FILLER_56_1795 ();
 sg13g2_fill_2 FILLER_56_1859 ();
 sg13g2_decap_8 FILLER_56_1871 ();
 sg13g2_decap_4 FILLER_56_1878 ();
 sg13g2_fill_1 FILLER_56_1882 ();
 sg13g2_fill_1 FILLER_56_1909 ();
 sg13g2_fill_1 FILLER_56_1915 ();
 sg13g2_fill_1 FILLER_56_1920 ();
 sg13g2_fill_2 FILLER_56_1925 ();
 sg13g2_fill_2 FILLER_56_1945 ();
 sg13g2_fill_2 FILLER_56_1954 ();
 sg13g2_fill_1 FILLER_56_1978 ();
 sg13g2_fill_1 FILLER_56_2017 ();
 sg13g2_decap_4 FILLER_56_2044 ();
 sg13g2_fill_1 FILLER_56_2053 ();
 sg13g2_fill_1 FILLER_56_2080 ();
 sg13g2_fill_1 FILLER_56_2107 ();
 sg13g2_fill_2 FILLER_56_2121 ();
 sg13g2_fill_2 FILLER_56_2142 ();
 sg13g2_decap_8 FILLER_56_2156 ();
 sg13g2_fill_1 FILLER_56_2163 ();
 sg13g2_fill_2 FILLER_56_2192 ();
 sg13g2_fill_1 FILLER_56_2194 ();
 sg13g2_decap_4 FILLER_56_2199 ();
 sg13g2_fill_1 FILLER_56_2207 ();
 sg13g2_fill_2 FILLER_56_2220 ();
 sg13g2_fill_2 FILLER_56_2226 ();
 sg13g2_fill_1 FILLER_56_2228 ();
 sg13g2_fill_2 FILLER_56_2233 ();
 sg13g2_fill_1 FILLER_56_2235 ();
 sg13g2_fill_2 FILLER_56_2257 ();
 sg13g2_fill_1 FILLER_56_2259 ();
 sg13g2_fill_2 FILLER_56_2302 ();
 sg13g2_fill_1 FILLER_56_2313 ();
 sg13g2_fill_1 FILLER_56_2341 ();
 sg13g2_fill_2 FILLER_56_2351 ();
 sg13g2_fill_1 FILLER_56_2362 ();
 sg13g2_fill_1 FILLER_56_2389 ();
 sg13g2_fill_1 FILLER_56_2411 ();
 sg13g2_fill_1 FILLER_56_2436 ();
 sg13g2_fill_1 FILLER_56_2442 ();
 sg13g2_fill_1 FILLER_56_2464 ();
 sg13g2_fill_1 FILLER_56_2538 ();
 sg13g2_fill_1 FILLER_56_2544 ();
 sg13g2_fill_1 FILLER_56_2557 ();
 sg13g2_fill_2 FILLER_56_2580 ();
 sg13g2_fill_1 FILLER_56_2582 ();
 sg13g2_decap_8 FILLER_56_2586 ();
 sg13g2_fill_2 FILLER_56_2593 ();
 sg13g2_decap_8 FILLER_56_2616 ();
 sg13g2_decap_8 FILLER_56_2623 ();
 sg13g2_decap_8 FILLER_56_2655 ();
 sg13g2_decap_8 FILLER_56_2662 ();
 sg13g2_fill_1 FILLER_56_2669 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_5 ();
 sg13g2_fill_1 FILLER_57_11 ();
 sg13g2_fill_1 FILLER_57_16 ();
 sg13g2_fill_1 FILLER_57_26 ();
 sg13g2_decap_4 FILLER_57_31 ();
 sg13g2_fill_1 FILLER_57_35 ();
 sg13g2_fill_1 FILLER_57_42 ();
 sg13g2_fill_1 FILLER_57_60 ();
 sg13g2_decap_4 FILLER_57_114 ();
 sg13g2_decap_4 FILLER_57_127 ();
 sg13g2_fill_1 FILLER_57_131 ();
 sg13g2_decap_4 FILLER_57_144 ();
 sg13g2_fill_1 FILLER_57_148 ();
 sg13g2_decap_4 FILLER_57_153 ();
 sg13g2_fill_2 FILLER_57_157 ();
 sg13g2_fill_2 FILLER_57_163 ();
 sg13g2_fill_2 FILLER_57_170 ();
 sg13g2_fill_1 FILLER_57_172 ();
 sg13g2_fill_1 FILLER_57_177 ();
 sg13g2_fill_1 FILLER_57_182 ();
 sg13g2_decap_4 FILLER_57_209 ();
 sg13g2_fill_1 FILLER_57_231 ();
 sg13g2_decap_4 FILLER_57_241 ();
 sg13g2_decap_4 FILLER_57_251 ();
 sg13g2_fill_1 FILLER_57_255 ();
 sg13g2_decap_8 FILLER_57_260 ();
 sg13g2_decap_4 FILLER_57_267 ();
 sg13g2_fill_1 FILLER_57_271 ();
 sg13g2_fill_2 FILLER_57_285 ();
 sg13g2_decap_8 FILLER_57_310 ();
 sg13g2_decap_8 FILLER_57_317 ();
 sg13g2_decap_4 FILLER_57_324 ();
 sg13g2_fill_2 FILLER_57_342 ();
 sg13g2_fill_1 FILLER_57_374 ();
 sg13g2_fill_1 FILLER_57_380 ();
 sg13g2_fill_2 FILLER_57_430 ();
 sg13g2_fill_1 FILLER_57_461 ();
 sg13g2_fill_1 FILLER_57_487 ();
 sg13g2_fill_1 FILLER_57_525 ();
 sg13g2_fill_2 FILLER_57_560 ();
 sg13g2_fill_1 FILLER_57_587 ();
 sg13g2_fill_1 FILLER_57_625 ();
 sg13g2_fill_2 FILLER_57_641 ();
 sg13g2_fill_2 FILLER_57_669 ();
 sg13g2_fill_1 FILLER_57_680 ();
 sg13g2_fill_1 FILLER_57_728 ();
 sg13g2_fill_2 FILLER_57_733 ();
 sg13g2_fill_2 FILLER_57_739 ();
 sg13g2_fill_2 FILLER_57_815 ();
 sg13g2_decap_8 FILLER_57_824 ();
 sg13g2_decap_4 FILLER_57_831 ();
 sg13g2_fill_2 FILLER_57_839 ();
 sg13g2_fill_1 FILLER_57_852 ();
 sg13g2_decap_8 FILLER_57_860 ();
 sg13g2_decap_8 FILLER_57_867 ();
 sg13g2_fill_1 FILLER_57_878 ();
 sg13g2_fill_2 FILLER_57_909 ();
 sg13g2_fill_1 FILLER_57_941 ();
 sg13g2_fill_1 FILLER_57_991 ();
 sg13g2_fill_1 FILLER_57_1095 ();
 sg13g2_fill_2 FILLER_57_1122 ();
 sg13g2_fill_2 FILLER_57_1208 ();
 sg13g2_fill_1 FILLER_57_1280 ();
 sg13g2_fill_2 FILLER_57_1327 ();
 sg13g2_fill_2 FILLER_57_1338 ();
 sg13g2_fill_2 FILLER_57_1344 ();
 sg13g2_decap_8 FILLER_57_1381 ();
 sg13g2_decap_4 FILLER_57_1388 ();
 sg13g2_fill_2 FILLER_57_1392 ();
 sg13g2_fill_2 FILLER_57_1402 ();
 sg13g2_fill_1 FILLER_57_1422 ();
 sg13g2_fill_1 FILLER_57_1437 ();
 sg13g2_fill_1 FILLER_57_1454 ();
 sg13g2_fill_2 FILLER_57_1480 ();
 sg13g2_fill_1 FILLER_57_1482 ();
 sg13g2_fill_2 FILLER_57_1513 ();
 sg13g2_fill_1 FILLER_57_1515 ();
 sg13g2_fill_1 FILLER_57_1554 ();
 sg13g2_fill_1 FILLER_57_1559 ();
 sg13g2_fill_2 FILLER_57_1570 ();
 sg13g2_fill_2 FILLER_57_1601 ();
 sg13g2_fill_2 FILLER_57_1634 ();
 sg13g2_fill_1 FILLER_57_1636 ();
 sg13g2_fill_2 FILLER_57_1648 ();
 sg13g2_fill_2 FILLER_57_1687 ();
 sg13g2_fill_1 FILLER_57_1703 ();
 sg13g2_fill_1 FILLER_57_1716 ();
 sg13g2_fill_1 FILLER_57_1734 ();
 sg13g2_fill_1 FILLER_57_1831 ();
 sg13g2_fill_1 FILLER_57_1837 ();
 sg13g2_fill_2 FILLER_57_1918 ();
 sg13g2_fill_1 FILLER_57_1926 ();
 sg13g2_fill_2 FILLER_57_2016 ();
 sg13g2_fill_2 FILLER_57_2031 ();
 sg13g2_fill_2 FILLER_57_2037 ();
 sg13g2_fill_1 FILLER_57_2039 ();
 sg13g2_fill_1 FILLER_57_2061 ();
 sg13g2_fill_2 FILLER_57_2076 ();
 sg13g2_fill_1 FILLER_57_2081 ();
 sg13g2_decap_4 FILLER_57_2168 ();
 sg13g2_fill_1 FILLER_57_2172 ();
 sg13g2_fill_1 FILLER_57_2178 ();
 sg13g2_fill_1 FILLER_57_2196 ();
 sg13g2_fill_2 FILLER_57_2212 ();
 sg13g2_fill_1 FILLER_57_2218 ();
 sg13g2_decap_4 FILLER_57_2249 ();
 sg13g2_fill_1 FILLER_57_2253 ();
 sg13g2_fill_1 FILLER_57_2324 ();
 sg13g2_fill_2 FILLER_57_2367 ();
 sg13g2_fill_1 FILLER_57_2369 ();
 sg13g2_decap_4 FILLER_57_2400 ();
 sg13g2_fill_1 FILLER_57_2404 ();
 sg13g2_decap_8 FILLER_57_2431 ();
 sg13g2_fill_2 FILLER_57_2449 ();
 sg13g2_fill_1 FILLER_57_2451 ();
 sg13g2_decap_4 FILLER_57_2455 ();
 sg13g2_fill_1 FILLER_57_2463 ();
 sg13g2_fill_2 FILLER_57_2489 ();
 sg13g2_fill_1 FILLER_57_2491 ();
 sg13g2_decap_8 FILLER_57_2502 ();
 sg13g2_decap_8 FILLER_57_2509 ();
 sg13g2_fill_2 FILLER_57_2516 ();
 sg13g2_fill_1 FILLER_57_2518 ();
 sg13g2_fill_1 FILLER_57_2526 ();
 sg13g2_decap_8 FILLER_57_2531 ();
 sg13g2_fill_2 FILLER_57_2538 ();
 sg13g2_fill_1 FILLER_57_2560 ();
 sg13g2_decap_8 FILLER_57_2590 ();
 sg13g2_fill_2 FILLER_57_2597 ();
 sg13g2_decap_8 FILLER_57_2620 ();
 sg13g2_decap_8 FILLER_57_2627 ();
 sg13g2_decap_4 FILLER_57_2634 ();
 sg13g2_decap_8 FILLER_57_2659 ();
 sg13g2_decap_4 FILLER_57_2666 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_10 ();
 sg13g2_fill_1 FILLER_58_20 ();
 sg13g2_fill_1 FILLER_58_29 ();
 sg13g2_fill_1 FILLER_58_56 ();
 sg13g2_fill_1 FILLER_58_109 ();
 sg13g2_fill_2 FILLER_58_118 ();
 sg13g2_fill_1 FILLER_58_124 ();
 sg13g2_fill_2 FILLER_58_129 ();
 sg13g2_decap_4 FILLER_58_136 ();
 sg13g2_decap_4 FILLER_58_158 ();
 sg13g2_fill_2 FILLER_58_162 ();
 sg13g2_decap_4 FILLER_58_177 ();
 sg13g2_fill_2 FILLER_58_186 ();
 sg13g2_fill_1 FILLER_58_188 ();
 sg13g2_fill_1 FILLER_58_193 ();
 sg13g2_decap_4 FILLER_58_208 ();
 sg13g2_fill_2 FILLER_58_217 ();
 sg13g2_fill_1 FILLER_58_219 ();
 sg13g2_fill_2 FILLER_58_275 ();
 sg13g2_fill_1 FILLER_58_290 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_fill_2 FILLER_58_329 ();
 sg13g2_fill_1 FILLER_58_331 ();
 sg13g2_fill_1 FILLER_58_481 ();
 sg13g2_fill_1 FILLER_58_493 ();
 sg13g2_fill_1 FILLER_58_498 ();
 sg13g2_fill_2 FILLER_58_505 ();
 sg13g2_fill_1 FILLER_58_629 ();
 sg13g2_fill_1 FILLER_58_639 ();
 sg13g2_fill_1 FILLER_58_671 ();
 sg13g2_fill_1 FILLER_58_706 ();
 sg13g2_fill_1 FILLER_58_729 ();
 sg13g2_fill_2 FILLER_58_734 ();
 sg13g2_fill_2 FILLER_58_862 ();
 sg13g2_fill_1 FILLER_58_981 ();
 sg13g2_fill_1 FILLER_58_991 ();
 sg13g2_fill_2 FILLER_58_1004 ();
 sg13g2_fill_2 FILLER_58_1024 ();
 sg13g2_fill_2 FILLER_58_1114 ();
 sg13g2_fill_1 FILLER_58_1163 ();
 sg13g2_fill_2 FILLER_58_1203 ();
 sg13g2_fill_2 FILLER_58_1229 ();
 sg13g2_fill_2 FILLER_58_1257 ();
 sg13g2_fill_2 FILLER_58_1280 ();
 sg13g2_fill_1 FILLER_58_1312 ();
 sg13g2_fill_1 FILLER_58_1317 ();
 sg13g2_fill_2 FILLER_58_1358 ();
 sg13g2_fill_2 FILLER_58_1379 ();
 sg13g2_fill_1 FILLER_58_1381 ();
 sg13g2_decap_8 FILLER_58_1388 ();
 sg13g2_decap_8 FILLER_58_1395 ();
 sg13g2_fill_2 FILLER_58_1402 ();
 sg13g2_fill_1 FILLER_58_1432 ();
 sg13g2_fill_1 FILLER_58_1442 ();
 sg13g2_fill_1 FILLER_58_1463 ();
 sg13g2_fill_2 FILLER_58_1507 ();
 sg13g2_decap_4 FILLER_58_1532 ();
 sg13g2_fill_1 FILLER_58_1536 ();
 sg13g2_fill_1 FILLER_58_1609 ();
 sg13g2_decap_4 FILLER_58_1636 ();
 sg13g2_fill_1 FILLER_58_1640 ();
 sg13g2_fill_2 FILLER_58_1671 ();
 sg13g2_fill_2 FILLER_58_1710 ();
 sg13g2_fill_2 FILLER_58_1724 ();
 sg13g2_fill_2 FILLER_58_1760 ();
 sg13g2_fill_2 FILLER_58_1775 ();
 sg13g2_fill_1 FILLER_58_1817 ();
 sg13g2_fill_2 FILLER_58_1889 ();
 sg13g2_fill_1 FILLER_58_1964 ();
 sg13g2_fill_2 FILLER_58_1969 ();
 sg13g2_fill_2 FILLER_58_1976 ();
 sg13g2_decap_4 FILLER_58_2004 ();
 sg13g2_fill_1 FILLER_58_2008 ();
 sg13g2_decap_4 FILLER_58_2022 ();
 sg13g2_fill_2 FILLER_58_2026 ();
 sg13g2_fill_2 FILLER_58_2036 ();
 sg13g2_fill_1 FILLER_58_2071 ();
 sg13g2_fill_1 FILLER_58_2078 ();
 sg13g2_fill_1 FILLER_58_2127 ();
 sg13g2_fill_2 FILLER_58_2154 ();
 sg13g2_fill_1 FILLER_58_2189 ();
 sg13g2_fill_1 FILLER_58_2205 ();
 sg13g2_fill_2 FILLER_58_2215 ();
 sg13g2_fill_1 FILLER_58_2226 ();
 sg13g2_fill_2 FILLER_58_2232 ();
 sg13g2_fill_1 FILLER_58_2273 ();
 sg13g2_fill_2 FILLER_58_2282 ();
 sg13g2_fill_1 FILLER_58_2284 ();
 sg13g2_fill_1 FILLER_58_2289 ();
 sg13g2_fill_1 FILLER_58_2304 ();
 sg13g2_fill_1 FILLER_58_2317 ();
 sg13g2_fill_2 FILLER_58_2342 ();
 sg13g2_fill_2 FILLER_58_2351 ();
 sg13g2_decap_4 FILLER_58_2371 ();
 sg13g2_fill_1 FILLER_58_2375 ();
 sg13g2_decap_8 FILLER_58_2407 ();
 sg13g2_decap_8 FILLER_58_2420 ();
 sg13g2_decap_4 FILLER_58_2427 ();
 sg13g2_fill_1 FILLER_58_2431 ();
 sg13g2_fill_1 FILLER_58_2476 ();
 sg13g2_decap_4 FILLER_58_2488 ();
 sg13g2_fill_1 FILLER_58_2496 ();
 sg13g2_fill_2 FILLER_58_2502 ();
 sg13g2_fill_2 FILLER_58_2525 ();
 sg13g2_fill_2 FILLER_58_2532 ();
 sg13g2_fill_1 FILLER_58_2534 ();
 sg13g2_fill_2 FILLER_58_2540 ();
 sg13g2_fill_2 FILLER_58_2547 ();
 sg13g2_decap_4 FILLER_58_2621 ();
 sg13g2_fill_1 FILLER_58_2636 ();
 sg13g2_decap_8 FILLER_58_2663 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_15 ();
 sg13g2_fill_1 FILLER_59_25 ();
 sg13g2_fill_1 FILLER_59_87 ();
 sg13g2_fill_1 FILLER_59_92 ();
 sg13g2_fill_2 FILLER_59_97 ();
 sg13g2_fill_2 FILLER_59_130 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_1 FILLER_59_187 ();
 sg13g2_fill_2 FILLER_59_217 ();
 sg13g2_fill_1 FILLER_59_219 ();
 sg13g2_fill_2 FILLER_59_224 ();
 sg13g2_fill_1 FILLER_59_273 ();
 sg13g2_fill_1 FILLER_59_279 ();
 sg13g2_fill_1 FILLER_59_333 ();
 sg13g2_fill_1 FILLER_59_351 ();
 sg13g2_fill_2 FILLER_59_405 ();
 sg13g2_fill_2 FILLER_59_480 ();
 sg13g2_fill_2 FILLER_59_485 ();
 sg13g2_fill_1 FILLER_59_515 ();
 sg13g2_fill_1 FILLER_59_563 ();
 sg13g2_fill_2 FILLER_59_569 ();
 sg13g2_fill_1 FILLER_59_579 ();
 sg13g2_fill_1 FILLER_59_600 ();
 sg13g2_fill_1 FILLER_59_623 ();
 sg13g2_fill_1 FILLER_59_628 ();
 sg13g2_fill_1 FILLER_59_641 ();
 sg13g2_fill_2 FILLER_59_653 ();
 sg13g2_fill_2 FILLER_59_670 ();
 sg13g2_fill_1 FILLER_59_676 ();
 sg13g2_fill_1 FILLER_59_682 ();
 sg13g2_fill_1 FILLER_59_688 ();
 sg13g2_fill_1 FILLER_59_767 ();
 sg13g2_fill_2 FILLER_59_779 ();
 sg13g2_fill_1 FILLER_59_818 ();
 sg13g2_fill_2 FILLER_59_849 ();
 sg13g2_fill_1 FILLER_59_851 ();
 sg13g2_fill_2 FILLER_59_895 ();
 sg13g2_fill_1 FILLER_59_961 ();
 sg13g2_fill_2 FILLER_59_1041 ();
 sg13g2_fill_1 FILLER_59_1047 ();
 sg13g2_fill_2 FILLER_59_1077 ();
 sg13g2_fill_2 FILLER_59_1096 ();
 sg13g2_fill_2 FILLER_59_1129 ();
 sg13g2_fill_1 FILLER_59_1144 ();
 sg13g2_fill_2 FILLER_59_1195 ();
 sg13g2_fill_1 FILLER_59_1204 ();
 sg13g2_fill_1 FILLER_59_1209 ();
 sg13g2_fill_1 FILLER_59_1271 ();
 sg13g2_fill_1 FILLER_59_1276 ();
 sg13g2_fill_1 FILLER_59_1281 ();
 sg13g2_fill_1 FILLER_59_1381 ();
 sg13g2_fill_1 FILLER_59_1385 ();
 sg13g2_fill_2 FILLER_59_1449 ();
 sg13g2_decap_8 FILLER_59_1519 ();
 sg13g2_decap_8 FILLER_59_1526 ();
 sg13g2_fill_1 FILLER_59_1533 ();
 sg13g2_decap_8 FILLER_59_1548 ();
 sg13g2_decap_4 FILLER_59_1555 ();
 sg13g2_fill_1 FILLER_59_1559 ();
 sg13g2_fill_2 FILLER_59_1592 ();
 sg13g2_fill_1 FILLER_59_1594 ();
 sg13g2_fill_2 FILLER_59_1598 ();
 sg13g2_decap_8 FILLER_59_1625 ();
 sg13g2_decap_4 FILLER_59_1632 ();
 sg13g2_fill_2 FILLER_59_1644 ();
 sg13g2_fill_1 FILLER_59_1646 ();
 sg13g2_fill_1 FILLER_59_1662 ();
 sg13g2_fill_2 FILLER_59_1764 ();
 sg13g2_fill_1 FILLER_59_1792 ();
 sg13g2_fill_2 FILLER_59_1804 ();
 sg13g2_fill_1 FILLER_59_1818 ();
 sg13g2_fill_2 FILLER_59_1828 ();
 sg13g2_fill_2 FILLER_59_1862 ();
 sg13g2_fill_1 FILLER_59_1922 ();
 sg13g2_fill_1 FILLER_59_1953 ();
 sg13g2_fill_1 FILLER_59_1959 ();
 sg13g2_fill_2 FILLER_59_1999 ();
 sg13g2_fill_2 FILLER_59_2005 ();
 sg13g2_fill_2 FILLER_59_2021 ();
 sg13g2_fill_1 FILLER_59_2023 ();
 sg13g2_fill_2 FILLER_59_2070 ();
 sg13g2_fill_1 FILLER_59_2107 ();
 sg13g2_fill_1 FILLER_59_2147 ();
 sg13g2_decap_8 FILLER_59_2226 ();
 sg13g2_decap_4 FILLER_59_2233 ();
 sg13g2_decap_8 FILLER_59_2263 ();
 sg13g2_decap_8 FILLER_59_2270 ();
 sg13g2_fill_2 FILLER_59_2277 ();
 sg13g2_fill_1 FILLER_59_2279 ();
 sg13g2_decap_8 FILLER_59_2284 ();
 sg13g2_fill_2 FILLER_59_2291 ();
 sg13g2_fill_1 FILLER_59_2293 ();
 sg13g2_fill_2 FILLER_59_2299 ();
 sg13g2_fill_1 FILLER_59_2306 ();
 sg13g2_fill_2 FILLER_59_2314 ();
 sg13g2_decap_4 FILLER_59_2342 ();
 sg13g2_decap_4 FILLER_59_2350 ();
 sg13g2_fill_2 FILLER_59_2358 ();
 sg13g2_fill_1 FILLER_59_2360 ();
 sg13g2_fill_2 FILLER_59_2366 ();
 sg13g2_fill_1 FILLER_59_2376 ();
 sg13g2_fill_2 FILLER_59_2404 ();
 sg13g2_fill_2 FILLER_59_2451 ();
 sg13g2_decap_8 FILLER_59_2457 ();
 sg13g2_fill_1 FILLER_59_2464 ();
 sg13g2_fill_2 FILLER_59_2538 ();
 sg13g2_decap_8 FILLER_59_2583 ();
 sg13g2_fill_1 FILLER_59_2590 ();
 sg13g2_fill_1 FILLER_59_2595 ();
 sg13g2_decap_8 FILLER_59_2626 ();
 sg13g2_decap_8 FILLER_59_2663 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_27 ();
 sg13g2_fill_2 FILLER_60_96 ();
 sg13g2_fill_1 FILLER_60_189 ();
 sg13g2_fill_2 FILLER_60_275 ();
 sg13g2_fill_2 FILLER_60_286 ();
 sg13g2_fill_2 FILLER_60_292 ();
 sg13g2_fill_1 FILLER_60_364 ();
 sg13g2_fill_1 FILLER_60_374 ();
 sg13g2_fill_1 FILLER_60_427 ();
 sg13g2_fill_2 FILLER_60_459 ();
 sg13g2_fill_1 FILLER_60_481 ();
 sg13g2_fill_2 FILLER_60_486 ();
 sg13g2_fill_2 FILLER_60_497 ();
 sg13g2_fill_2 FILLER_60_519 ();
 sg13g2_fill_1 FILLER_60_550 ();
 sg13g2_fill_1 FILLER_60_577 ();
 sg13g2_fill_2 FILLER_60_583 ();
 sg13g2_fill_1 FILLER_60_615 ();
 sg13g2_fill_2 FILLER_60_646 ();
 sg13g2_fill_2 FILLER_60_656 ();
 sg13g2_fill_2 FILLER_60_662 ();
 sg13g2_fill_2 FILLER_60_671 ();
 sg13g2_fill_1 FILLER_60_676 ();
 sg13g2_fill_1 FILLER_60_694 ();
 sg13g2_fill_1 FILLER_60_700 ();
 sg13g2_fill_1 FILLER_60_705 ();
 sg13g2_fill_1 FILLER_60_710 ();
 sg13g2_fill_2 FILLER_60_737 ();
 sg13g2_fill_1 FILLER_60_778 ();
 sg13g2_fill_2 FILLER_60_789 ();
 sg13g2_fill_1 FILLER_60_821 ();
 sg13g2_fill_2 FILLER_60_856 ();
 sg13g2_fill_1 FILLER_60_863 ();
 sg13g2_fill_2 FILLER_60_868 ();
 sg13g2_fill_1 FILLER_60_870 ();
 sg13g2_fill_2 FILLER_60_904 ();
 sg13g2_fill_1 FILLER_60_915 ();
 sg13g2_fill_1 FILLER_60_923 ();
 sg13g2_fill_1 FILLER_60_1000 ();
 sg13g2_fill_2 FILLER_60_1018 ();
 sg13g2_fill_2 FILLER_60_1053 ();
 sg13g2_fill_1 FILLER_60_1067 ();
 sg13g2_fill_2 FILLER_60_1072 ();
 sg13g2_fill_1 FILLER_60_1081 ();
 sg13g2_fill_1 FILLER_60_1104 ();
 sg13g2_fill_2 FILLER_60_1147 ();
 sg13g2_fill_2 FILLER_60_1156 ();
 sg13g2_fill_2 FILLER_60_1199 ();
 sg13g2_fill_2 FILLER_60_1205 ();
 sg13g2_fill_2 FILLER_60_1262 ();
 sg13g2_fill_2 FILLER_60_1302 ();
 sg13g2_fill_2 FILLER_60_1316 ();
 sg13g2_fill_1 FILLER_60_1327 ();
 sg13g2_fill_1 FILLER_60_1331 ();
 sg13g2_fill_2 FILLER_60_1340 ();
 sg13g2_fill_1 FILLER_60_1364 ();
 sg13g2_fill_1 FILLER_60_1448 ();
 sg13g2_fill_1 FILLER_60_1458 ();
 sg13g2_decap_8 FILLER_60_1490 ();
 sg13g2_fill_2 FILLER_60_1497 ();
 sg13g2_decap_8 FILLER_60_1503 ();
 sg13g2_decap_8 FILLER_60_1510 ();
 sg13g2_fill_1 FILLER_60_1517 ();
 sg13g2_decap_8 FILLER_60_1528 ();
 sg13g2_decap_4 FILLER_60_1535 ();
 sg13g2_fill_1 FILLER_60_1539 ();
 sg13g2_fill_1 FILLER_60_1599 ();
 sg13g2_fill_2 FILLER_60_1626 ();
 sg13g2_decap_8 FILLER_60_1633 ();
 sg13g2_decap_8 FILLER_60_1640 ();
 sg13g2_fill_1 FILLER_60_1673 ();
 sg13g2_fill_2 FILLER_60_1700 ();
 sg13g2_fill_1 FILLER_60_1710 ();
 sg13g2_fill_2 FILLER_60_1715 ();
 sg13g2_fill_1 FILLER_60_1717 ();
 sg13g2_fill_1 FILLER_60_1729 ();
 sg13g2_fill_2 FILLER_60_1792 ();
 sg13g2_fill_2 FILLER_60_1857 ();
 sg13g2_fill_2 FILLER_60_1868 ();
 sg13g2_fill_2 FILLER_60_1887 ();
 sg13g2_fill_2 FILLER_60_1902 ();
 sg13g2_fill_2 FILLER_60_1917 ();
 sg13g2_fill_1 FILLER_60_1938 ();
 sg13g2_fill_2 FILLER_60_1953 ();
 sg13g2_fill_2 FILLER_60_2052 ();
 sg13g2_fill_1 FILLER_60_2054 ();
 sg13g2_fill_1 FILLER_60_2094 ();
 sg13g2_fill_2 FILLER_60_2106 ();
 sg13g2_fill_1 FILLER_60_2132 ();
 sg13g2_fill_2 FILLER_60_2151 ();
 sg13g2_fill_1 FILLER_60_2156 ();
 sg13g2_fill_1 FILLER_60_2204 ();
 sg13g2_fill_1 FILLER_60_2213 ();
 sg13g2_fill_1 FILLER_60_2218 ();
 sg13g2_decap_8 FILLER_60_2229 ();
 sg13g2_decap_4 FILLER_60_2236 ();
 sg13g2_fill_1 FILLER_60_2240 ();
 sg13g2_fill_2 FILLER_60_2258 ();
 sg13g2_fill_2 FILLER_60_2270 ();
 sg13g2_fill_2 FILLER_60_2277 ();
 sg13g2_decap_8 FILLER_60_2284 ();
 sg13g2_fill_2 FILLER_60_2291 ();
 sg13g2_fill_1 FILLER_60_2293 ();
 sg13g2_decap_8 FILLER_60_2298 ();
 sg13g2_fill_2 FILLER_60_2312 ();
 sg13g2_fill_2 FILLER_60_2322 ();
 sg13g2_fill_1 FILLER_60_2331 ();
 sg13g2_fill_2 FILLER_60_2336 ();
 sg13g2_fill_2 FILLER_60_2377 ();
 sg13g2_fill_1 FILLER_60_2379 ();
 sg13g2_fill_2 FILLER_60_2405 ();
 sg13g2_fill_1 FILLER_60_2407 ();
 sg13g2_fill_1 FILLER_60_2434 ();
 sg13g2_decap_8 FILLER_60_2456 ();
 sg13g2_decap_4 FILLER_60_2468 ();
 sg13g2_fill_1 FILLER_60_2472 ();
 sg13g2_fill_1 FILLER_60_2503 ();
 sg13g2_fill_2 FILLER_60_2544 ();
 sg13g2_fill_1 FILLER_60_2559 ();
 sg13g2_fill_2 FILLER_60_2573 ();
 sg13g2_fill_1 FILLER_60_2580 ();
 sg13g2_decap_8 FILLER_60_2587 ();
 sg13g2_fill_2 FILLER_60_2594 ();
 sg13g2_decap_4 FILLER_60_2618 ();
 sg13g2_fill_1 FILLER_60_2633 ();
 sg13g2_decap_8 FILLER_60_2651 ();
 sg13g2_decap_8 FILLER_60_2658 ();
 sg13g2_decap_4 FILLER_60_2665 ();
 sg13g2_fill_1 FILLER_60_2669 ();
 sg13g2_fill_1 FILLER_61_50 ();
 sg13g2_fill_1 FILLER_61_85 ();
 sg13g2_fill_2 FILLER_61_103 ();
 sg13g2_fill_1 FILLER_61_144 ();
 sg13g2_fill_1 FILLER_61_223 ();
 sg13g2_fill_2 FILLER_61_233 ();
 sg13g2_fill_1 FILLER_61_251 ();
 sg13g2_fill_1 FILLER_61_256 ();
 sg13g2_fill_2 FILLER_61_288 ();
 sg13g2_fill_1 FILLER_61_298 ();
 sg13g2_fill_1 FILLER_61_308 ();
 sg13g2_fill_1 FILLER_61_313 ();
 sg13g2_fill_1 FILLER_61_318 ();
 sg13g2_fill_1 FILLER_61_345 ();
 sg13g2_fill_1 FILLER_61_354 ();
 sg13g2_fill_1 FILLER_61_432 ();
 sg13g2_fill_1 FILLER_61_473 ();
 sg13g2_fill_1 FILLER_61_563 ();
 sg13g2_fill_2 FILLER_61_589 ();
 sg13g2_fill_1 FILLER_61_600 ();
 sg13g2_fill_1 FILLER_61_605 ();
 sg13g2_fill_2 FILLER_61_610 ();
 sg13g2_fill_1 FILLER_61_667 ();
 sg13g2_fill_1 FILLER_61_672 ();
 sg13g2_fill_1 FILLER_61_694 ();
 sg13g2_fill_2 FILLER_61_699 ();
 sg13g2_fill_1 FILLER_61_711 ();
 sg13g2_fill_1 FILLER_61_732 ();
 sg13g2_fill_1 FILLER_61_782 ();
 sg13g2_fill_1 FILLER_61_825 ();
 sg13g2_fill_2 FILLER_61_835 ();
 sg13g2_fill_1 FILLER_61_837 ();
 sg13g2_fill_2 FILLER_61_857 ();
 sg13g2_fill_1 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_893 ();
 sg13g2_fill_1 FILLER_61_935 ();
 sg13g2_fill_1 FILLER_61_941 ();
 sg13g2_fill_2 FILLER_61_979 ();
 sg13g2_fill_2 FILLER_61_1011 ();
 sg13g2_fill_1 FILLER_61_1061 ();
 sg13g2_fill_1 FILLER_61_1080 ();
 sg13g2_fill_1 FILLER_61_1093 ();
 sg13g2_fill_1 FILLER_61_1109 ();
 sg13g2_fill_1 FILLER_61_1130 ();
 sg13g2_fill_1 FILLER_61_1203 ();
 sg13g2_fill_1 FILLER_61_1220 ();
 sg13g2_fill_1 FILLER_61_1305 ();
 sg13g2_fill_1 FILLER_61_1341 ();
 sg13g2_fill_2 FILLER_61_1352 ();
 sg13g2_fill_2 FILLER_61_1357 ();
 sg13g2_fill_2 FILLER_61_1376 ();
 sg13g2_fill_1 FILLER_61_1391 ();
 sg13g2_fill_1 FILLER_61_1397 ();
 sg13g2_fill_1 FILLER_61_1402 ();
 sg13g2_fill_1 FILLER_61_1407 ();
 sg13g2_fill_2 FILLER_61_1417 ();
 sg13g2_fill_1 FILLER_61_1454 ();
 sg13g2_decap_8 FILLER_61_1485 ();
 sg13g2_fill_2 FILLER_61_1492 ();
 sg13g2_fill_1 FILLER_61_1494 ();
 sg13g2_fill_2 FILLER_61_1523 ();
 sg13g2_fill_2 FILLER_61_1530 ();
 sg13g2_fill_1 FILLER_61_1532 ();
 sg13g2_decap_4 FILLER_61_1571 ();
 sg13g2_fill_2 FILLER_61_1575 ();
 sg13g2_fill_2 FILLER_61_1589 ();
 sg13g2_decap_8 FILLER_61_1632 ();
 sg13g2_decap_8 FILLER_61_1639 ();
 sg13g2_fill_2 FILLER_61_1689 ();
 sg13g2_fill_2 FILLER_61_1717 ();
 sg13g2_fill_1 FILLER_61_1784 ();
 sg13g2_fill_1 FILLER_61_1796 ();
 sg13g2_fill_2 FILLER_61_1843 ();
 sg13g2_fill_1 FILLER_61_1871 ();
 sg13g2_fill_2 FILLER_61_1924 ();
 sg13g2_fill_2 FILLER_61_1988 ();
 sg13g2_decap_8 FILLER_61_1998 ();
 sg13g2_fill_2 FILLER_61_2005 ();
 sg13g2_fill_1 FILLER_61_2007 ();
 sg13g2_fill_1 FILLER_61_2017 ();
 sg13g2_fill_1 FILLER_61_2026 ();
 sg13g2_fill_2 FILLER_61_2032 ();
 sg13g2_fill_1 FILLER_61_2034 ();
 sg13g2_fill_1 FILLER_61_2085 ();
 sg13g2_fill_2 FILLER_61_2101 ();
 sg13g2_fill_1 FILLER_61_2124 ();
 sg13g2_fill_1 FILLER_61_2134 ();
 sg13g2_fill_2 FILLER_61_2175 ();
 sg13g2_fill_2 FILLER_61_2187 ();
 sg13g2_fill_1 FILLER_61_2225 ();
 sg13g2_decap_8 FILLER_61_2234 ();
 sg13g2_fill_2 FILLER_61_2241 ();
 sg13g2_fill_1 FILLER_61_2247 ();
 sg13g2_fill_1 FILLER_61_2256 ();
 sg13g2_fill_1 FILLER_61_2266 ();
 sg13g2_decap_8 FILLER_61_2281 ();
 sg13g2_fill_1 FILLER_61_2293 ();
 sg13g2_decap_4 FILLER_61_2302 ();
 sg13g2_decap_4 FILLER_61_2315 ();
 sg13g2_fill_1 FILLER_61_2319 ();
 sg13g2_decap_4 FILLER_61_2328 ();
 sg13g2_fill_2 FILLER_61_2336 ();
 sg13g2_fill_1 FILLER_61_2346 ();
 sg13g2_fill_1 FILLER_61_2352 ();
 sg13g2_fill_1 FILLER_61_2358 ();
 sg13g2_fill_1 FILLER_61_2372 ();
 sg13g2_fill_2 FILLER_61_2378 ();
 sg13g2_decap_8 FILLER_61_2434 ();
 sg13g2_fill_2 FILLER_61_2441 ();
 sg13g2_decap_8 FILLER_61_2447 ();
 sg13g2_decap_4 FILLER_61_2466 ();
 sg13g2_fill_2 FILLER_61_2470 ();
 sg13g2_fill_2 FILLER_61_2477 ();
 sg13g2_decap_4 FILLER_61_2483 ();
 sg13g2_fill_2 FILLER_61_2491 ();
 sg13g2_fill_2 FILLER_61_2504 ();
 sg13g2_fill_2 FILLER_61_2510 ();
 sg13g2_decap_8 FILLER_61_2516 ();
 sg13g2_fill_2 FILLER_61_2523 ();
 sg13g2_decap_4 FILLER_61_2538 ();
 sg13g2_fill_1 FILLER_61_2542 ();
 sg13g2_fill_2 FILLER_61_2548 ();
 sg13g2_fill_1 FILLER_61_2550 ();
 sg13g2_decap_8 FILLER_61_2567 ();
 sg13g2_fill_1 FILLER_61_2584 ();
 sg13g2_decap_4 FILLER_61_2589 ();
 sg13g2_fill_1 FILLER_61_2593 ();
 sg13g2_decap_8 FILLER_61_2599 ();
 sg13g2_decap_4 FILLER_61_2606 ();
 sg13g2_fill_1 FILLER_61_2610 ();
 sg13g2_decap_4 FILLER_61_2624 ();
 sg13g2_fill_2 FILLER_61_2628 ();
 sg13g2_decap_8 FILLER_61_2636 ();
 sg13g2_decap_8 FILLER_61_2643 ();
 sg13g2_decap_8 FILLER_61_2650 ();
 sg13g2_decap_8 FILLER_61_2657 ();
 sg13g2_decap_4 FILLER_61_2664 ();
 sg13g2_fill_2 FILLER_61_2668 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_44 ();
 sg13g2_fill_1 FILLER_62_138 ();
 sg13g2_fill_1 FILLER_62_146 ();
 sg13g2_fill_1 FILLER_62_160 ();
 sg13g2_fill_2 FILLER_62_211 ();
 sg13g2_fill_1 FILLER_62_226 ();
 sg13g2_fill_1 FILLER_62_245 ();
 sg13g2_fill_1 FILLER_62_279 ();
 sg13g2_fill_1 FILLER_62_292 ();
 sg13g2_fill_2 FILLER_62_324 ();
 sg13g2_fill_2 FILLER_62_377 ();
 sg13g2_fill_2 FILLER_62_386 ();
 sg13g2_fill_1 FILLER_62_449 ();
 sg13g2_fill_2 FILLER_62_521 ();
 sg13g2_decap_4 FILLER_62_624 ();
 sg13g2_fill_1 FILLER_62_667 ();
 sg13g2_fill_1 FILLER_62_703 ();
 sg13g2_fill_2 FILLER_62_724 ();
 sg13g2_fill_1 FILLER_62_729 ();
 sg13g2_fill_1 FILLER_62_782 ();
 sg13g2_fill_1 FILLER_62_787 ();
 sg13g2_fill_2 FILLER_62_814 ();
 sg13g2_fill_1 FILLER_62_816 ();
 sg13g2_fill_2 FILLER_62_821 ();
 sg13g2_fill_1 FILLER_62_823 ();
 sg13g2_fill_2 FILLER_62_841 ();
 sg13g2_fill_1 FILLER_62_874 ();
 sg13g2_fill_1 FILLER_62_943 ();
 sg13g2_fill_2 FILLER_62_954 ();
 sg13g2_fill_1 FILLER_62_960 ();
 sg13g2_fill_1 FILLER_62_990 ();
 sg13g2_fill_2 FILLER_62_1007 ();
 sg13g2_fill_1 FILLER_62_1060 ();
 sg13g2_fill_2 FILLER_62_1132 ();
 sg13g2_fill_2 FILLER_62_1172 ();
 sg13g2_fill_1 FILLER_62_1187 ();
 sg13g2_fill_2 FILLER_62_1232 ();
 sg13g2_fill_2 FILLER_62_1314 ();
 sg13g2_fill_1 FILLER_62_1372 ();
 sg13g2_fill_2 FILLER_62_1416 ();
 sg13g2_fill_1 FILLER_62_1418 ();
 sg13g2_fill_1 FILLER_62_1424 ();
 sg13g2_fill_1 FILLER_62_1429 ();
 sg13g2_fill_2 FILLER_62_1434 ();
 sg13g2_decap_8 FILLER_62_1440 ();
 sg13g2_fill_1 FILLER_62_1447 ();
 sg13g2_decap_8 FILLER_62_1456 ();
 sg13g2_decap_4 FILLER_62_1463 ();
 sg13g2_decap_4 FILLER_62_1475 ();
 sg13g2_fill_1 FILLER_62_1479 ();
 sg13g2_decap_8 FILLER_62_1484 ();
 sg13g2_fill_1 FILLER_62_1491 ();
 sg13g2_fill_2 FILLER_62_1518 ();
 sg13g2_fill_2 FILLER_62_1553 ();
 sg13g2_fill_1 FILLER_62_1555 ();
 sg13g2_fill_2 FILLER_62_1632 ();
 sg13g2_decap_8 FILLER_62_1647 ();
 sg13g2_fill_2 FILLER_62_1654 ();
 sg13g2_fill_1 FILLER_62_1656 ();
 sg13g2_fill_2 FILLER_62_1666 ();
 sg13g2_fill_1 FILLER_62_1668 ();
 sg13g2_fill_2 FILLER_62_1673 ();
 sg13g2_decap_8 FILLER_62_1679 ();
 sg13g2_fill_1 FILLER_62_1686 ();
 sg13g2_fill_2 FILLER_62_1691 ();
 sg13g2_fill_1 FILLER_62_1693 ();
 sg13g2_fill_1 FILLER_62_1718 ();
 sg13g2_fill_1 FILLER_62_1723 ();
 sg13g2_fill_2 FILLER_62_1740 ();
 sg13g2_fill_1 FILLER_62_1742 ();
 sg13g2_fill_1 FILLER_62_1749 ();
 sg13g2_fill_2 FILLER_62_1758 ();
 sg13g2_fill_1 FILLER_62_1764 ();
 sg13g2_fill_2 FILLER_62_1769 ();
 sg13g2_fill_1 FILLER_62_1771 ();
 sg13g2_fill_2 FILLER_62_1793 ();
 sg13g2_fill_2 FILLER_62_1843 ();
 sg13g2_fill_1 FILLER_62_1875 ();
 sg13g2_fill_1 FILLER_62_1890 ();
 sg13g2_fill_2 FILLER_62_1895 ();
 sg13g2_fill_2 FILLER_62_1902 ();
 sg13g2_fill_1 FILLER_62_1904 ();
 sg13g2_fill_1 FILLER_62_1932 ();
 sg13g2_fill_1 FILLER_62_1941 ();
 sg13g2_fill_1 FILLER_62_1981 ();
 sg13g2_fill_1 FILLER_62_1986 ();
 sg13g2_fill_2 FILLER_62_1991 ();
 sg13g2_fill_2 FILLER_62_2014 ();
 sg13g2_fill_1 FILLER_62_2020 ();
 sg13g2_fill_2 FILLER_62_2030 ();
 sg13g2_fill_1 FILLER_62_2032 ();
 sg13g2_fill_2 FILLER_62_2049 ();
 sg13g2_fill_1 FILLER_62_2051 ();
 sg13g2_fill_2 FILLER_62_2056 ();
 sg13g2_decap_4 FILLER_62_2070 ();
 sg13g2_fill_2 FILLER_62_2077 ();
 sg13g2_fill_1 FILLER_62_2106 ();
 sg13g2_fill_2 FILLER_62_2141 ();
 sg13g2_fill_1 FILLER_62_2150 ();
 sg13g2_fill_1 FILLER_62_2227 ();
 sg13g2_fill_1 FILLER_62_2259 ();
 sg13g2_fill_2 FILLER_62_2268 ();
 sg13g2_fill_2 FILLER_62_2301 ();
 sg13g2_decap_8 FILLER_62_2338 ();
 sg13g2_decap_8 FILLER_62_2345 ();
 sg13g2_decap_4 FILLER_62_2352 ();
 sg13g2_fill_1 FILLER_62_2356 ();
 sg13g2_fill_1 FILLER_62_2397 ();
 sg13g2_fill_2 FILLER_62_2409 ();
 sg13g2_fill_1 FILLER_62_2417 ();
 sg13g2_fill_2 FILLER_62_2444 ();
 sg13g2_fill_2 FILLER_62_2467 ();
 sg13g2_fill_2 FILLER_62_2474 ();
 sg13g2_fill_1 FILLER_62_2476 ();
 sg13g2_fill_1 FILLER_62_2497 ();
 sg13g2_fill_2 FILLER_62_2523 ();
 sg13g2_fill_1 FILLER_62_2530 ();
 sg13g2_fill_2 FILLER_62_2536 ();
 sg13g2_decap_8 FILLER_62_2558 ();
 sg13g2_fill_1 FILLER_62_2565 ();
 sg13g2_decap_4 FILLER_62_2571 ();
 sg13g2_fill_1 FILLER_62_2575 ();
 sg13g2_fill_2 FILLER_62_2594 ();
 sg13g2_fill_1 FILLER_62_2596 ();
 sg13g2_fill_2 FILLER_62_2608 ();
 sg13g2_fill_1 FILLER_62_2610 ();
 sg13g2_fill_1 FILLER_62_2633 ();
 sg13g2_fill_2 FILLER_62_2639 ();
 sg13g2_fill_2 FILLER_62_2667 ();
 sg13g2_fill_1 FILLER_62_2669 ();
 sg13g2_fill_2 FILLER_63_40 ();
 sg13g2_fill_2 FILLER_63_45 ();
 sg13g2_fill_2 FILLER_63_73 ();
 sg13g2_fill_2 FILLER_63_80 ();
 sg13g2_fill_1 FILLER_63_107 ();
 sg13g2_fill_1 FILLER_63_115 ();
 sg13g2_fill_1 FILLER_63_158 ();
 sg13g2_fill_2 FILLER_63_181 ();
 sg13g2_fill_2 FILLER_63_217 ();
 sg13g2_fill_2 FILLER_63_223 ();
 sg13g2_fill_1 FILLER_63_251 ();
 sg13g2_fill_2 FILLER_63_257 ();
 sg13g2_fill_2 FILLER_63_289 ();
 sg13g2_fill_1 FILLER_63_333 ();
 sg13g2_fill_1 FILLER_63_379 ();
 sg13g2_fill_2 FILLER_63_392 ();
 sg13g2_fill_1 FILLER_63_412 ();
 sg13g2_fill_1 FILLER_63_482 ();
 sg13g2_fill_2 FILLER_63_528 ();
 sg13g2_fill_1 FILLER_63_530 ();
 sg13g2_fill_2 FILLER_63_606 ();
 sg13g2_fill_2 FILLER_63_634 ();
 sg13g2_fill_1 FILLER_63_636 ();
 sg13g2_fill_1 FILLER_63_646 ();
 sg13g2_fill_1 FILLER_63_673 ();
 sg13g2_fill_2 FILLER_63_700 ();
 sg13g2_fill_1 FILLER_63_731 ();
 sg13g2_fill_2 FILLER_63_739 ();
 sg13g2_fill_1 FILLER_63_767 ();
 sg13g2_fill_2 FILLER_63_776 ();
 sg13g2_fill_2 FILLER_63_786 ();
 sg13g2_fill_2 FILLER_63_861 ();
 sg13g2_fill_1 FILLER_63_863 ();
 sg13g2_fill_1 FILLER_63_946 ();
 sg13g2_fill_1 FILLER_63_964 ();
 sg13g2_fill_1 FILLER_63_1002 ();
 sg13g2_fill_2 FILLER_63_1015 ();
 sg13g2_fill_1 FILLER_63_1051 ();
 sg13g2_fill_2 FILLER_63_1091 ();
 sg13g2_fill_1 FILLER_63_1119 ();
 sg13g2_fill_1 FILLER_63_1154 ();
 sg13g2_fill_2 FILLER_63_1159 ();
 sg13g2_fill_2 FILLER_63_1177 ();
 sg13g2_fill_1 FILLER_63_1253 ();
 sg13g2_fill_1 FILLER_63_1275 ();
 sg13g2_fill_2 FILLER_63_1331 ();
 sg13g2_fill_2 FILLER_63_1405 ();
 sg13g2_decap_8 FILLER_63_1440 ();
 sg13g2_decap_8 FILLER_63_1447 ();
 sg13g2_fill_1 FILLER_63_1454 ();
 sg13g2_decap_8 FILLER_63_1459 ();
 sg13g2_decap_8 FILLER_63_1466 ();
 sg13g2_fill_2 FILLER_63_1473 ();
 sg13g2_fill_1 FILLER_63_1475 ();
 sg13g2_fill_1 FILLER_63_1480 ();
 sg13g2_fill_1 FILLER_63_1516 ();
 sg13g2_fill_1 FILLER_63_1544 ();
 sg13g2_fill_2 FILLER_63_1562 ();
 sg13g2_fill_1 FILLER_63_1611 ();
 sg13g2_decap_8 FILLER_63_1652 ();
 sg13g2_decap_8 FILLER_63_1659 ();
 sg13g2_fill_2 FILLER_63_1666 ();
 sg13g2_fill_2 FILLER_63_1698 ();
 sg13g2_fill_1 FILLER_63_1700 ();
 sg13g2_fill_2 FILLER_63_1758 ();
 sg13g2_fill_1 FILLER_63_1760 ();
 sg13g2_fill_1 FILLER_63_1770 ();
 sg13g2_fill_2 FILLER_63_1820 ();
 sg13g2_fill_2 FILLER_63_1855 ();
 sg13g2_fill_1 FILLER_63_1878 ();
 sg13g2_fill_2 FILLER_63_1938 ();
 sg13g2_fill_1 FILLER_63_1970 ();
 sg13g2_fill_1 FILLER_63_1975 ();
 sg13g2_fill_1 FILLER_63_2017 ();
 sg13g2_fill_1 FILLER_63_2023 ();
 sg13g2_fill_1 FILLER_63_2050 ();
 sg13g2_fill_2 FILLER_63_2085 ();
 sg13g2_fill_2 FILLER_63_2109 ();
 sg13g2_fill_1 FILLER_63_2126 ();
 sg13g2_fill_1 FILLER_63_2158 ();
 sg13g2_fill_2 FILLER_63_2276 ();
 sg13g2_fill_2 FILLER_63_2289 ();
 sg13g2_fill_2 FILLER_63_2295 ();
 sg13g2_fill_1 FILLER_63_2336 ();
 sg13g2_fill_1 FILLER_63_2363 ();
 sg13g2_fill_1 FILLER_63_2385 ();
 sg13g2_decap_4 FILLER_63_2521 ();
 sg13g2_fill_2 FILLER_63_2525 ();
 sg13g2_fill_1 FILLER_63_2564 ();
 sg13g2_fill_2 FILLER_63_2570 ();
 sg13g2_fill_2 FILLER_63_2577 ();
 sg13g2_fill_2 FILLER_63_2587 ();
 sg13g2_fill_1 FILLER_63_2589 ();
 sg13g2_decap_8 FILLER_63_2611 ();
 sg13g2_decap_4 FILLER_63_2618 ();
 sg13g2_fill_1 FILLER_63_2622 ();
 sg13g2_fill_1 FILLER_63_2629 ();
 sg13g2_fill_2 FILLER_63_2635 ();
 sg13g2_fill_1 FILLER_63_2663 ();
 sg13g2_fill_2 FILLER_63_2668 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_55 ();
 sg13g2_fill_1 FILLER_64_81 ();
 sg13g2_fill_2 FILLER_64_171 ();
 sg13g2_fill_1 FILLER_64_250 ();
 sg13g2_fill_2 FILLER_64_289 ();
 sg13g2_fill_1 FILLER_64_299 ();
 sg13g2_fill_1 FILLER_64_304 ();
 sg13g2_fill_2 FILLER_64_316 ();
 sg13g2_fill_1 FILLER_64_325 ();
 sg13g2_fill_2 FILLER_64_353 ();
 sg13g2_fill_2 FILLER_64_359 ();
 sg13g2_fill_2 FILLER_64_370 ();
 sg13g2_fill_1 FILLER_64_401 ();
 sg13g2_fill_1 FILLER_64_432 ();
 sg13g2_fill_1 FILLER_64_438 ();
 sg13g2_fill_1 FILLER_64_512 ();
 sg13g2_fill_2 FILLER_64_584 ();
 sg13g2_fill_1 FILLER_64_611 ();
 sg13g2_fill_2 FILLER_64_651 ();
 sg13g2_fill_1 FILLER_64_679 ();
 sg13g2_fill_2 FILLER_64_697 ();
 sg13g2_fill_2 FILLER_64_759 ();
 sg13g2_fill_2 FILLER_64_811 ();
 sg13g2_fill_2 FILLER_64_838 ();
 sg13g2_fill_1 FILLER_64_840 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_fill_2 FILLER_64_856 ();
 sg13g2_fill_2 FILLER_64_892 ();
 sg13g2_fill_1 FILLER_64_907 ();
 sg13g2_fill_2 FILLER_64_912 ();
 sg13g2_fill_2 FILLER_64_1014 ();
 sg13g2_fill_1 FILLER_64_1024 ();
 sg13g2_fill_1 FILLER_64_1062 ();
 sg13g2_fill_2 FILLER_64_1097 ();
 sg13g2_fill_2 FILLER_64_1117 ();
 sg13g2_fill_1 FILLER_64_1162 ();
 sg13g2_fill_1 FILLER_64_1221 ();
 sg13g2_fill_1 FILLER_64_1226 ();
 sg13g2_fill_2 FILLER_64_1235 ();
 sg13g2_fill_1 FILLER_64_1266 ();
 sg13g2_fill_1 FILLER_64_1291 ();
 sg13g2_fill_1 FILLER_64_1307 ();
 sg13g2_fill_1 FILLER_64_1319 ();
 sg13g2_fill_1 FILLER_64_1367 ();
 sg13g2_fill_1 FILLER_64_1412 ();
 sg13g2_fill_2 FILLER_64_1444 ();
 sg13g2_fill_1 FILLER_64_1476 ();
 sg13g2_fill_2 FILLER_64_1490 ();
 sg13g2_fill_1 FILLER_64_1496 ();
 sg13g2_decap_8 FILLER_64_1527 ();
 sg13g2_fill_2 FILLER_64_1534 ();
 sg13g2_fill_1 FILLER_64_1536 ();
 sg13g2_decap_8 FILLER_64_1542 ();
 sg13g2_fill_1 FILLER_64_1558 ();
 sg13g2_fill_1 FILLER_64_1563 ();
 sg13g2_fill_1 FILLER_64_1568 ();
 sg13g2_fill_1 FILLER_64_1573 ();
 sg13g2_fill_2 FILLER_64_1578 ();
 sg13g2_fill_1 FILLER_64_1584 ();
 sg13g2_fill_1 FILLER_64_1590 ();
 sg13g2_fill_1 FILLER_64_1631 ();
 sg13g2_decap_8 FILLER_64_1663 ();
 sg13g2_decap_8 FILLER_64_1670 ();
 sg13g2_fill_1 FILLER_64_1677 ();
 sg13g2_decap_4 FILLER_64_1687 ();
 sg13g2_fill_2 FILLER_64_1691 ();
 sg13g2_fill_1 FILLER_64_1718 ();
 sg13g2_fill_1 FILLER_64_1728 ();
 sg13g2_fill_1 FILLER_64_1734 ();
 sg13g2_fill_1 FILLER_64_1808 ();
 sg13g2_decap_8 FILLER_64_1867 ();
 sg13g2_fill_1 FILLER_64_1926 ();
 sg13g2_fill_1 FILLER_64_1930 ();
 sg13g2_fill_2 FILLER_64_1969 ();
 sg13g2_fill_1 FILLER_64_2058 ();
 sg13g2_fill_2 FILLER_64_2074 ();
 sg13g2_fill_1 FILLER_64_2097 ();
 sg13g2_fill_2 FILLER_64_2101 ();
 sg13g2_fill_2 FILLER_64_2108 ();
 sg13g2_fill_1 FILLER_64_2187 ();
 sg13g2_fill_2 FILLER_64_2226 ();
 sg13g2_fill_1 FILLER_64_2258 ();
 sg13g2_fill_2 FILLER_64_2264 ();
 sg13g2_decap_4 FILLER_64_2292 ();
 sg13g2_fill_1 FILLER_64_2296 ();
 sg13g2_fill_1 FILLER_64_2302 ();
 sg13g2_decap_8 FILLER_64_2309 ();
 sg13g2_fill_1 FILLER_64_2324 ();
 sg13g2_fill_1 FILLER_64_2332 ();
 sg13g2_decap_4 FILLER_64_2338 ();
 sg13g2_fill_2 FILLER_64_2346 ();
 sg13g2_decap_4 FILLER_64_2352 ();
 sg13g2_decap_8 FILLER_64_2377 ();
 sg13g2_decap_4 FILLER_64_2384 ();
 sg13g2_fill_1 FILLER_64_2460 ();
 sg13g2_fill_2 FILLER_64_2468 ();
 sg13g2_fill_1 FILLER_64_2470 ();
 sg13g2_fill_2 FILLER_64_2480 ();
 sg13g2_fill_1 FILLER_64_2499 ();
 sg13g2_decap_8 FILLER_64_2521 ();
 sg13g2_decap_4 FILLER_64_2528 ();
 sg13g2_fill_2 FILLER_64_2532 ();
 sg13g2_fill_1 FILLER_64_2583 ();
 sg13g2_fill_2 FILLER_64_2605 ();
 sg13g2_fill_1 FILLER_64_2628 ();
 sg13g2_decap_4 FILLER_64_2635 ();
 sg13g2_fill_1 FILLER_64_2639 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_13 ();
 sg13g2_fill_1 FILLER_65_66 ();
 sg13g2_fill_1 FILLER_65_108 ();
 sg13g2_fill_1 FILLER_65_123 ();
 sg13g2_fill_2 FILLER_65_159 ();
 sg13g2_fill_2 FILLER_65_204 ();
 sg13g2_fill_2 FILLER_65_236 ();
 sg13g2_fill_2 FILLER_65_253 ();
 sg13g2_fill_1 FILLER_65_289 ();
 sg13g2_fill_1 FILLER_65_312 ();
 sg13g2_fill_1 FILLER_65_332 ();
 sg13g2_fill_1 FILLER_65_337 ();
 sg13g2_fill_2 FILLER_65_342 ();
 sg13g2_fill_2 FILLER_65_360 ();
 sg13g2_fill_1 FILLER_65_456 ();
 sg13g2_fill_1 FILLER_65_488 ();
 sg13g2_fill_1 FILLER_65_630 ();
 sg13g2_decap_4 FILLER_65_635 ();
 sg13g2_fill_1 FILLER_65_644 ();
 sg13g2_decap_8 FILLER_65_649 ();
 sg13g2_fill_2 FILLER_65_656 ();
 sg13g2_fill_1 FILLER_65_658 ();
 sg13g2_decap_8 FILLER_65_664 ();
 sg13g2_fill_2 FILLER_65_671 ();
 sg13g2_fill_1 FILLER_65_673 ();
 sg13g2_fill_2 FILLER_65_692 ();
 sg13g2_fill_2 FILLER_65_713 ();
 sg13g2_fill_2 FILLER_65_780 ();
 sg13g2_fill_2 FILLER_65_799 ();
 sg13g2_decap_4 FILLER_65_810 ();
 sg13g2_fill_2 FILLER_65_835 ();
 sg13g2_decap_8 FILLER_65_846 ();
 sg13g2_fill_1 FILLER_65_853 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_fill_2 FILLER_65_981 ();
 sg13g2_fill_1 FILLER_65_1020 ();
 sg13g2_fill_1 FILLER_65_1052 ();
 sg13g2_fill_2 FILLER_65_1084 ();
 sg13g2_fill_1 FILLER_65_1097 ();
 sg13g2_fill_1 FILLER_65_1102 ();
 sg13g2_fill_1 FILLER_65_1161 ();
 sg13g2_fill_1 FILLER_65_1185 ();
 sg13g2_fill_2 FILLER_65_1195 ();
 sg13g2_fill_2 FILLER_65_1207 ();
 sg13g2_fill_1 FILLER_65_1243 ();
 sg13g2_fill_2 FILLER_65_1270 ();
 sg13g2_fill_2 FILLER_65_1310 ();
 sg13g2_decap_8 FILLER_65_1321 ();
 sg13g2_fill_1 FILLER_65_1356 ();
 sg13g2_fill_1 FILLER_65_1364 ();
 sg13g2_fill_1 FILLER_65_1370 ();
 sg13g2_fill_2 FILLER_65_1376 ();
 sg13g2_fill_1 FILLER_65_1417 ();
 sg13g2_fill_2 FILLER_65_1446 ();
 sg13g2_decap_4 FILLER_65_1452 ();
 sg13g2_fill_2 FILLER_65_1461 ();
 sg13g2_fill_1 FILLER_65_1463 ();
 sg13g2_fill_2 FILLER_65_1476 ();
 sg13g2_fill_2 FILLER_65_1492 ();
 sg13g2_fill_2 FILLER_65_1505 ();
 sg13g2_fill_1 FILLER_65_1520 ();
 sg13g2_fill_2 FILLER_65_1529 ();
 sg13g2_decap_8 FILLER_65_1536 ();
 sg13g2_fill_1 FILLER_65_1543 ();
 sg13g2_decap_8 FILLER_65_1548 ();
 sg13g2_decap_8 FILLER_65_1555 ();
 sg13g2_fill_1 FILLER_65_1562 ();
 sg13g2_fill_2 FILLER_65_1572 ();
 sg13g2_decap_4 FILLER_65_1663 ();
 sg13g2_decap_4 FILLER_65_1693 ();
 sg13g2_fill_1 FILLER_65_1727 ();
 sg13g2_fill_1 FILLER_65_1754 ();
 sg13g2_decap_8 FILLER_65_1760 ();
 sg13g2_fill_2 FILLER_65_1775 ();
 sg13g2_fill_2 FILLER_65_1783 ();
 sg13g2_fill_1 FILLER_65_1785 ();
 sg13g2_decap_4 FILLER_65_1819 ();
 sg13g2_fill_2 FILLER_65_1827 ();
 sg13g2_fill_2 FILLER_65_1888 ();
 sg13g2_fill_1 FILLER_65_1890 ();
 sg13g2_decap_4 FILLER_65_1903 ();
 sg13g2_fill_1 FILLER_65_1925 ();
 sg13g2_fill_2 FILLER_65_1944 ();
 sg13g2_fill_2 FILLER_65_1950 ();
 sg13g2_fill_2 FILLER_65_1967 ();
 sg13g2_fill_2 FILLER_65_1986 ();
 sg13g2_decap_4 FILLER_65_2017 ();
 sg13g2_fill_2 FILLER_65_2025 ();
 sg13g2_fill_1 FILLER_65_2027 ();
 sg13g2_fill_1 FILLER_65_2065 ();
 sg13g2_fill_1 FILLER_65_2092 ();
 sg13g2_fill_2 FILLER_65_2130 ();
 sg13g2_fill_2 FILLER_65_2153 ();
 sg13g2_fill_2 FILLER_65_2180 ();
 sg13g2_fill_2 FILLER_65_2192 ();
 sg13g2_fill_1 FILLER_65_2203 ();
 sg13g2_fill_1 FILLER_65_2294 ();
 sg13g2_decap_4 FILLER_65_2300 ();
 sg13g2_fill_2 FILLER_65_2304 ();
 sg13g2_decap_4 FILLER_65_2310 ();
 sg13g2_fill_1 FILLER_65_2314 ();
 sg13g2_fill_1 FILLER_65_2325 ();
 sg13g2_fill_2 FILLER_65_2334 ();
 sg13g2_fill_1 FILLER_65_2336 ();
 sg13g2_decap_4 FILLER_65_2341 ();
 sg13g2_decap_4 FILLER_65_2350 ();
 sg13g2_fill_1 FILLER_65_2375 ();
 sg13g2_fill_2 FILLER_65_2400 ();
 sg13g2_fill_1 FILLER_65_2402 ();
 sg13g2_decap_8 FILLER_65_2407 ();
 sg13g2_decap_4 FILLER_65_2414 ();
 sg13g2_fill_1 FILLER_65_2418 ();
 sg13g2_decap_8 FILLER_65_2426 ();
 sg13g2_decap_4 FILLER_65_2433 ();
 sg13g2_decap_8 FILLER_65_2461 ();
 sg13g2_fill_2 FILLER_65_2494 ();
 sg13g2_fill_1 FILLER_65_2506 ();
 sg13g2_fill_2 FILLER_65_2528 ();
 sg13g2_fill_2 FILLER_65_2539 ();
 sg13g2_fill_1 FILLER_65_2541 ();
 sg13g2_fill_2 FILLER_65_2562 ();
 sg13g2_decap_8 FILLER_65_2600 ();
 sg13g2_fill_1 FILLER_65_2607 ();
 sg13g2_decap_8 FILLER_65_2629 ();
 sg13g2_fill_1 FILLER_65_2636 ();
 sg13g2_fill_1 FILLER_65_2658 ();
 sg13g2_decap_8 FILLER_65_2663 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_110 ();
 sg13g2_fill_1 FILLER_66_116 ();
 sg13g2_fill_1 FILLER_66_121 ();
 sg13g2_fill_2 FILLER_66_143 ();
 sg13g2_fill_2 FILLER_66_187 ();
 sg13g2_fill_2 FILLER_66_348 ();
 sg13g2_fill_2 FILLER_66_376 ();
 sg13g2_fill_2 FILLER_66_390 ();
 sg13g2_fill_1 FILLER_66_403 ();
 sg13g2_fill_1 FILLER_66_420 ();
 sg13g2_fill_1 FILLER_66_449 ();
 sg13g2_fill_2 FILLER_66_457 ();
 sg13g2_fill_2 FILLER_66_467 ();
 sg13g2_fill_1 FILLER_66_473 ();
 sg13g2_fill_1 FILLER_66_507 ();
 sg13g2_fill_1 FILLER_66_557 ();
 sg13g2_fill_1 FILLER_66_565 ();
 sg13g2_fill_1 FILLER_66_572 ();
 sg13g2_fill_1 FILLER_66_611 ();
 sg13g2_fill_2 FILLER_66_625 ();
 sg13g2_fill_1 FILLER_66_666 ();
 sg13g2_fill_2 FILLER_66_677 ();
 sg13g2_fill_1 FILLER_66_686 ();
 sg13g2_fill_2 FILLER_66_704 ();
 sg13g2_fill_1 FILLER_66_718 ();
 sg13g2_fill_2 FILLER_66_728 ();
 sg13g2_fill_2 FILLER_66_734 ();
 sg13g2_fill_1 FILLER_66_739 ();
 sg13g2_fill_2 FILLER_66_764 ();
 sg13g2_fill_2 FILLER_66_771 ();
 sg13g2_fill_1 FILLER_66_781 ();
 sg13g2_fill_2 FILLER_66_816 ();
 sg13g2_decap_4 FILLER_66_848 ();
 sg13g2_fill_2 FILLER_66_861 ();
 sg13g2_fill_1 FILLER_66_870 ();
 sg13g2_fill_1 FILLER_66_875 ();
 sg13g2_fill_2 FILLER_66_961 ();
 sg13g2_fill_1 FILLER_66_994 ();
 sg13g2_fill_2 FILLER_66_1025 ();
 sg13g2_fill_2 FILLER_66_1037 ();
 sg13g2_fill_1 FILLER_66_1089 ();
 sg13g2_fill_2 FILLER_66_1146 ();
 sg13g2_fill_2 FILLER_66_1178 ();
 sg13g2_fill_1 FILLER_66_1283 ();
 sg13g2_fill_1 FILLER_66_1298 ();
 sg13g2_decap_4 FILLER_66_1329 ();
 sg13g2_fill_2 FILLER_66_1333 ();
 sg13g2_fill_2 FILLER_66_1356 ();
 sg13g2_fill_1 FILLER_66_1414 ();
 sg13g2_fill_2 FILLER_66_1441 ();
 sg13g2_fill_1 FILLER_66_1443 ();
 sg13g2_fill_2 FILLER_66_1474 ();
 sg13g2_fill_2 FILLER_66_1513 ();
 sg13g2_fill_1 FILLER_66_1541 ();
 sg13g2_fill_1 FILLER_66_1551 ();
 sg13g2_fill_1 FILLER_66_1556 ();
 sg13g2_fill_1 FILLER_66_1561 ();
 sg13g2_fill_2 FILLER_66_1566 ();
 sg13g2_fill_2 FILLER_66_1633 ();
 sg13g2_fill_1 FILLER_66_1642 ();
 sg13g2_fill_1 FILLER_66_1739 ();
 sg13g2_fill_2 FILLER_66_1745 ();
 sg13g2_fill_1 FILLER_66_1747 ();
 sg13g2_decap_8 FILLER_66_1784 ();
 sg13g2_decap_8 FILLER_66_1791 ();
 sg13g2_decap_4 FILLER_66_1798 ();
 sg13g2_fill_2 FILLER_66_1828 ();
 sg13g2_fill_1 FILLER_66_1830 ();
 sg13g2_fill_2 FILLER_66_1853 ();
 sg13g2_fill_2 FILLER_66_1869 ();
 sg13g2_fill_2 FILLER_66_1925 ();
 sg13g2_fill_2 FILLER_66_1959 ();
 sg13g2_decap_8 FILLER_66_2010 ();
 sg13g2_decap_8 FILLER_66_2017 ();
 sg13g2_decap_8 FILLER_66_2024 ();
 sg13g2_decap_8 FILLER_66_2031 ();
 sg13g2_decap_8 FILLER_66_2038 ();
 sg13g2_fill_1 FILLER_66_2049 ();
 sg13g2_fill_2 FILLER_66_2071 ();
 sg13g2_fill_2 FILLER_66_2093 ();
 sg13g2_fill_1 FILLER_66_2188 ();
 sg13g2_fill_2 FILLER_66_2196 ();
 sg13g2_fill_2 FILLER_66_2268 ();
 sg13g2_fill_2 FILLER_66_2274 ();
 sg13g2_fill_2 FILLER_66_2302 ();
 sg13g2_fill_1 FILLER_66_2304 ();
 sg13g2_decap_8 FILLER_66_2309 ();
 sg13g2_fill_1 FILLER_66_2316 ();
 sg13g2_decap_4 FILLER_66_2322 ();
 sg13g2_fill_2 FILLER_66_2326 ();
 sg13g2_fill_1 FILLER_66_2340 ();
 sg13g2_fill_2 FILLER_66_2345 ();
 sg13g2_fill_1 FILLER_66_2373 ();
 sg13g2_decap_8 FILLER_66_2395 ();
 sg13g2_decap_8 FILLER_66_2402 ();
 sg13g2_fill_2 FILLER_66_2409 ();
 sg13g2_fill_2 FILLER_66_2434 ();
 sg13g2_fill_1 FILLER_66_2446 ();
 sg13g2_decap_8 FILLER_66_2450 ();
 sg13g2_decap_8 FILLER_66_2513 ();
 sg13g2_decap_8 FILLER_66_2520 ();
 sg13g2_decap_4 FILLER_66_2527 ();
 sg13g2_fill_2 FILLER_66_2531 ();
 sg13g2_fill_2 FILLER_66_2567 ();
 sg13g2_fill_1 FILLER_66_2569 ();
 sg13g2_fill_1 FILLER_66_2607 ();
 sg13g2_decap_8 FILLER_66_2631 ();
 sg13g2_fill_1 FILLER_66_2638 ();
 sg13g2_decap_4 FILLER_66_2665 ();
 sg13g2_fill_1 FILLER_66_2669 ();
 sg13g2_fill_1 FILLER_67_33 ();
 sg13g2_fill_1 FILLER_67_153 ();
 sg13g2_fill_1 FILLER_67_180 ();
 sg13g2_fill_1 FILLER_67_259 ();
 sg13g2_fill_1 FILLER_67_273 ();
 sg13g2_fill_1 FILLER_67_279 ();
 sg13g2_fill_2 FILLER_67_351 ();
 sg13g2_fill_2 FILLER_67_374 ();
 sg13g2_fill_2 FILLER_67_384 ();
 sg13g2_fill_2 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_67_439 ();
 sg13g2_fill_2 FILLER_67_448 ();
 sg13g2_fill_1 FILLER_67_494 ();
 sg13g2_fill_1 FILLER_67_577 ();
 sg13g2_fill_1 FILLER_67_582 ();
 sg13g2_fill_2 FILLER_67_591 ();
 sg13g2_fill_1 FILLER_67_598 ();
 sg13g2_fill_1 FILLER_67_602 ();
 sg13g2_fill_2 FILLER_67_606 ();
 sg13g2_fill_2 FILLER_67_641 ();
 sg13g2_fill_1 FILLER_67_643 ();
 sg13g2_fill_2 FILLER_67_647 ();
 sg13g2_fill_1 FILLER_67_697 ();
 sg13g2_fill_2 FILLER_67_705 ();
 sg13g2_fill_1 FILLER_67_711 ();
 sg13g2_fill_2 FILLER_67_717 ();
 sg13g2_fill_1 FILLER_67_728 ();
 sg13g2_fill_1 FILLER_67_745 ();
 sg13g2_fill_2 FILLER_67_853 ();
 sg13g2_fill_1 FILLER_67_855 ();
 sg13g2_fill_2 FILLER_67_895 ();
 sg13g2_fill_2 FILLER_67_948 ();
 sg13g2_fill_2 FILLER_67_980 ();
 sg13g2_fill_2 FILLER_67_1021 ();
 sg13g2_fill_1 FILLER_67_1033 ();
 sg13g2_fill_1 FILLER_67_1066 ();
 sg13g2_fill_1 FILLER_67_1091 ();
 sg13g2_fill_1 FILLER_67_1119 ();
 sg13g2_fill_1 FILLER_67_1125 ();
 sg13g2_fill_1 FILLER_67_1203 ();
 sg13g2_fill_1 FILLER_67_1231 ();
 sg13g2_decap_4 FILLER_67_1313 ();
 sg13g2_fill_1 FILLER_67_1343 ();
 sg13g2_fill_1 FILLER_67_1349 ();
 sg13g2_fill_2 FILLER_67_1354 ();
 sg13g2_fill_1 FILLER_67_1363 ();
 sg13g2_fill_2 FILLER_67_1379 ();
 sg13g2_fill_2 FILLER_67_1415 ();
 sg13g2_fill_1 FILLER_67_1448 ();
 sg13g2_fill_1 FILLER_67_1480 ();
 sg13g2_fill_1 FILLER_67_1585 ();
 sg13g2_fill_2 FILLER_67_1590 ();
 sg13g2_fill_1 FILLER_67_1601 ();
 sg13g2_fill_2 FILLER_67_1606 ();
 sg13g2_fill_1 FILLER_67_1612 ();
 sg13g2_fill_2 FILLER_67_1626 ();
 sg13g2_decap_4 FILLER_67_1679 ();
 sg13g2_fill_1 FILLER_67_1688 ();
 sg13g2_fill_2 FILLER_67_1731 ();
 sg13g2_fill_2 FILLER_67_1770 ();
 sg13g2_decap_8 FILLER_67_1798 ();
 sg13g2_decap_8 FILLER_67_1808 ();
 sg13g2_fill_1 FILLER_67_1815 ();
 sg13g2_decap_8 FILLER_67_1822 ();
 sg13g2_fill_2 FILLER_67_1829 ();
 sg13g2_fill_1 FILLER_67_1831 ();
 sg13g2_decap_4 FILLER_67_1836 ();
 sg13g2_fill_1 FILLER_67_1866 ();
 sg13g2_fill_2 FILLER_67_1875 ();
 sg13g2_fill_2 FILLER_67_1917 ();
 sg13g2_fill_1 FILLER_67_1926 ();
 sg13g2_fill_2 FILLER_67_1935 ();
 sg13g2_fill_1 FILLER_67_1976 ();
 sg13g2_decap_8 FILLER_67_1984 ();
 sg13g2_fill_1 FILLER_67_1991 ();
 sg13g2_fill_1 FILLER_67_2023 ();
 sg13g2_decap_4 FILLER_67_2028 ();
 sg13g2_fill_1 FILLER_67_2032 ();
 sg13g2_fill_2 FILLER_67_2037 ();
 sg13g2_fill_1 FILLER_67_2039 ();
 sg13g2_fill_1 FILLER_67_2078 ();
 sg13g2_fill_1 FILLER_67_2090 ();
 sg13g2_fill_1 FILLER_67_2104 ();
 sg13g2_fill_1 FILLER_67_2123 ();
 sg13g2_fill_2 FILLER_67_2166 ();
 sg13g2_fill_2 FILLER_67_2193 ();
 sg13g2_fill_1 FILLER_67_2210 ();
 sg13g2_fill_1 FILLER_67_2223 ();
 sg13g2_fill_1 FILLER_67_2241 ();
 sg13g2_fill_2 FILLER_67_2251 ();
 sg13g2_decap_8 FILLER_67_2295 ();
 sg13g2_decap_8 FILLER_67_2302 ();
 sg13g2_decap_8 FILLER_67_2309 ();
 sg13g2_decap_4 FILLER_67_2316 ();
 sg13g2_fill_1 FILLER_67_2320 ();
 sg13g2_fill_2 FILLER_67_2328 ();
 sg13g2_decap_8 FILLER_67_2351 ();
 sg13g2_decap_8 FILLER_67_2358 ();
 sg13g2_fill_2 FILLER_67_2365 ();
 sg13g2_decap_8 FILLER_67_2375 ();
 sg13g2_decap_8 FILLER_67_2387 ();
 sg13g2_decap_4 FILLER_67_2394 ();
 sg13g2_fill_2 FILLER_67_2398 ();
 sg13g2_fill_1 FILLER_67_2406 ();
 sg13g2_decap_8 FILLER_67_2438 ();
 sg13g2_decap_8 FILLER_67_2445 ();
 sg13g2_fill_2 FILLER_67_2459 ();
 sg13g2_fill_1 FILLER_67_2503 ();
 sg13g2_fill_1 FILLER_67_2538 ();
 sg13g2_fill_2 FILLER_67_2548 ();
 sg13g2_decap_4 FILLER_67_2554 ();
 sg13g2_fill_2 FILLER_67_2558 ();
 sg13g2_decap_8 FILLER_67_2570 ();
 sg13g2_decap_4 FILLER_67_2577 ();
 sg13g2_fill_2 FILLER_67_2581 ();
 sg13g2_fill_1 FILLER_67_2633 ();
 sg13g2_decap_8 FILLER_67_2660 ();
 sg13g2_fill_2 FILLER_67_2667 ();
 sg13g2_fill_1 FILLER_67_2669 ();
 sg13g2_fill_1 FILLER_68_31 ();
 sg13g2_fill_1 FILLER_68_83 ();
 sg13g2_fill_2 FILLER_68_147 ();
 sg13g2_fill_1 FILLER_68_213 ();
 sg13g2_fill_1 FILLER_68_218 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_251 ();
 sg13g2_fill_1 FILLER_68_288 ();
 sg13g2_fill_2 FILLER_68_372 ();
 sg13g2_fill_2 FILLER_68_403 ();
 sg13g2_decap_8 FILLER_68_532 ();
 sg13g2_fill_1 FILLER_68_539 ();
 sg13g2_fill_1 FILLER_68_544 ();
 sg13g2_fill_2 FILLER_68_569 ();
 sg13g2_fill_1 FILLER_68_589 ();
 sg13g2_fill_1 FILLER_68_600 ();
 sg13g2_fill_2 FILLER_68_712 ();
 sg13g2_fill_1 FILLER_68_772 ();
 sg13g2_fill_2 FILLER_68_811 ();
 sg13g2_fill_1 FILLER_68_869 ();
 sg13g2_fill_2 FILLER_68_880 ();
 sg13g2_fill_1 FILLER_68_886 ();
 sg13g2_fill_1 FILLER_68_904 ();
 sg13g2_fill_1 FILLER_68_1049 ();
 sg13g2_fill_1 FILLER_68_1084 ();
 sg13g2_fill_1 FILLER_68_1095 ();
 sg13g2_fill_1 FILLER_68_1108 ();
 sg13g2_fill_2 FILLER_68_1142 ();
 sg13g2_fill_2 FILLER_68_1151 ();
 sg13g2_fill_2 FILLER_68_1158 ();
 sg13g2_fill_1 FILLER_68_1168 ();
 sg13g2_fill_1 FILLER_68_1179 ();
 sg13g2_fill_2 FILLER_68_1186 ();
 sg13g2_fill_2 FILLER_68_1215 ();
 sg13g2_fill_1 FILLER_68_1237 ();
 sg13g2_fill_2 FILLER_68_1286 ();
 sg13g2_fill_2 FILLER_68_1315 ();
 sg13g2_fill_2 FILLER_68_1452 ();
 sg13g2_fill_1 FILLER_68_1454 ();
 sg13g2_fill_1 FILLER_68_1476 ();
 sg13g2_fill_2 FILLER_68_1542 ();
 sg13g2_fill_1 FILLER_68_1544 ();
 sg13g2_fill_1 FILLER_68_1571 ();
 sg13g2_fill_1 FILLER_68_1576 ();
 sg13g2_fill_1 FILLER_68_1581 ();
 sg13g2_fill_2 FILLER_68_1587 ();
 sg13g2_decap_8 FILLER_68_1593 ();
 sg13g2_decap_4 FILLER_68_1600 ();
 sg13g2_fill_2 FILLER_68_1604 ();
 sg13g2_fill_1 FILLER_68_1702 ();
 sg13g2_fill_2 FILLER_68_1707 ();
 sg13g2_fill_1 FILLER_68_1751 ();
 sg13g2_fill_1 FILLER_68_1790 ();
 sg13g2_decap_4 FILLER_68_1795 ();
 sg13g2_fill_2 FILLER_68_1803 ();
 sg13g2_fill_2 FILLER_68_1819 ();
 sg13g2_decap_8 FILLER_68_1834 ();
 sg13g2_decap_8 FILLER_68_1841 ();
 sg13g2_decap_8 FILLER_68_1848 ();
 sg13g2_fill_2 FILLER_68_1855 ();
 sg13g2_fill_1 FILLER_68_1857 ();
 sg13g2_fill_1 FILLER_68_1871 ();
 sg13g2_fill_2 FILLER_68_1925 ();
 sg13g2_fill_1 FILLER_68_1959 ();
 sg13g2_fill_1 FILLER_68_1968 ();
 sg13g2_fill_1 FILLER_68_2032 ();
 sg13g2_fill_1 FILLER_68_2059 ();
 sg13g2_fill_2 FILLER_68_2069 ();
 sg13g2_fill_2 FILLER_68_2090 ();
 sg13g2_fill_2 FILLER_68_2112 ();
 sg13g2_fill_2 FILLER_68_2135 ();
 sg13g2_fill_2 FILLER_68_2155 ();
 sg13g2_fill_1 FILLER_68_2173 ();
 sg13g2_fill_1 FILLER_68_2191 ();
 sg13g2_fill_2 FILLER_68_2243 ();
 sg13g2_fill_1 FILLER_68_2274 ();
 sg13g2_decap_4 FILLER_68_2279 ();
 sg13g2_decap_8 FILLER_68_2288 ();
 sg13g2_decap_8 FILLER_68_2295 ();
 sg13g2_fill_2 FILLER_68_2302 ();
 sg13g2_fill_1 FILLER_68_2304 ();
 sg13g2_fill_1 FILLER_68_2309 ();
 sg13g2_fill_2 FILLER_68_2336 ();
 sg13g2_fill_1 FILLER_68_2338 ();
 sg13g2_fill_2 FILLER_68_2367 ();
 sg13g2_fill_2 FILLER_68_2380 ();
 sg13g2_fill_1 FILLER_68_2418 ();
 sg13g2_fill_2 FILLER_68_2423 ();
 sg13g2_fill_2 FILLER_68_2430 ();
 sg13g2_fill_1 FILLER_68_2432 ();
 sg13g2_fill_1 FILLER_68_2467 ();
 sg13g2_fill_2 FILLER_68_2480 ();
 sg13g2_fill_2 FILLER_68_2553 ();
 sg13g2_fill_2 FILLER_68_2560 ();
 sg13g2_decap_8 FILLER_68_2575 ();
 sg13g2_fill_2 FILLER_68_2582 ();
 sg13g2_decap_8 FILLER_68_2589 ();
 sg13g2_decap_8 FILLER_68_2600 ();
 sg13g2_decap_8 FILLER_68_2607 ();
 sg13g2_fill_1 FILLER_68_2614 ();
 sg13g2_decap_8 FILLER_68_2656 ();
 sg13g2_decap_8 FILLER_68_2663 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_63 ();
 sg13g2_fill_2 FILLER_69_69 ();
 sg13g2_fill_1 FILLER_69_161 ();
 sg13g2_fill_2 FILLER_69_205 ();
 sg13g2_fill_1 FILLER_69_216 ();
 sg13g2_fill_1 FILLER_69_221 ();
 sg13g2_fill_2 FILLER_69_323 ();
 sg13g2_fill_2 FILLER_69_363 ();
 sg13g2_fill_1 FILLER_69_400 ();
 sg13g2_fill_1 FILLER_69_432 ();
 sg13g2_fill_1 FILLER_69_465 ();
 sg13g2_fill_2 FILLER_69_508 ();
 sg13g2_decap_8 FILLER_69_518 ();
 sg13g2_decap_4 FILLER_69_525 ();
 sg13g2_decap_8 FILLER_69_533 ();
 sg13g2_decap_4 FILLER_69_540 ();
 sg13g2_fill_2 FILLER_69_573 ();
 sg13g2_fill_2 FILLER_69_606 ();
 sg13g2_decap_4 FILLER_69_625 ();
 sg13g2_fill_1 FILLER_69_679 ();
 sg13g2_fill_1 FILLER_69_695 ();
 sg13g2_fill_1 FILLER_69_711 ();
 sg13g2_fill_1 FILLER_69_748 ();
 sg13g2_fill_1 FILLER_69_780 ();
 sg13g2_fill_1 FILLER_69_792 ();
 sg13g2_fill_2 FILLER_69_816 ();
 sg13g2_fill_1 FILLER_69_827 ();
 sg13g2_fill_1 FILLER_69_832 ();
 sg13g2_fill_1 FILLER_69_859 ();
 sg13g2_fill_1 FILLER_69_935 ();
 sg13g2_fill_2 FILLER_69_966 ();
 sg13g2_fill_2 FILLER_69_972 ();
 sg13g2_fill_2 FILLER_69_1045 ();
 sg13g2_fill_1 FILLER_69_1103 ();
 sg13g2_fill_1 FILLER_69_1176 ();
 sg13g2_fill_2 FILLER_69_1207 ();
 sg13g2_fill_2 FILLER_69_1259 ();
 sg13g2_fill_1 FILLER_69_1327 ();
 sg13g2_fill_2 FILLER_69_1340 ();
 sg13g2_decap_8 FILLER_69_1454 ();
 sg13g2_fill_1 FILLER_69_1461 ();
 sg13g2_decap_8 FILLER_69_1465 ();
 sg13g2_decap_4 FILLER_69_1472 ();
 sg13g2_fill_2 FILLER_69_1476 ();
 sg13g2_fill_1 FILLER_69_1498 ();
 sg13g2_fill_1 FILLER_69_1507 ();
 sg13g2_fill_2 FILLER_69_1516 ();
 sg13g2_fill_1 FILLER_69_1542 ();
 sg13g2_fill_2 FILLER_69_1556 ();
 sg13g2_fill_1 FILLER_69_1558 ();
 sg13g2_decap_4 FILLER_69_1588 ();
 sg13g2_fill_1 FILLER_69_1592 ();
 sg13g2_fill_2 FILLER_69_1679 ();
 sg13g2_fill_1 FILLER_69_1718 ();
 sg13g2_fill_1 FILLER_69_1808 ();
 sg13g2_fill_2 FILLER_69_1835 ();
 sg13g2_fill_1 FILLER_69_1837 ();
 sg13g2_decap_4 FILLER_69_1842 ();
 sg13g2_fill_1 FILLER_69_1846 ();
 sg13g2_fill_2 FILLER_69_1852 ();
 sg13g2_fill_1 FILLER_69_1881 ();
 sg13g2_fill_1 FILLER_69_1936 ();
 sg13g2_fill_2 FILLER_69_1963 ();
 sg13g2_fill_2 FILLER_69_2002 ();
 sg13g2_fill_1 FILLER_69_2022 ();
 sg13g2_fill_1 FILLER_69_2028 ();
 sg13g2_fill_1 FILLER_69_2054 ();
 sg13g2_fill_1 FILLER_69_2088 ();
 sg13g2_fill_2 FILLER_69_2125 ();
 sg13g2_fill_1 FILLER_69_2140 ();
 sg13g2_fill_1 FILLER_69_2162 ();
 sg13g2_fill_1 FILLER_69_2171 ();
 sg13g2_fill_1 FILLER_69_2204 ();
 sg13g2_fill_1 FILLER_69_2218 ();
 sg13g2_fill_2 FILLER_69_2224 ();
 sg13g2_fill_2 FILLER_69_2277 ();
 sg13g2_fill_1 FILLER_69_2283 ();
 sg13g2_decap_4 FILLER_69_2291 ();
 sg13g2_fill_2 FILLER_69_2380 ();
 sg13g2_fill_1 FILLER_69_2382 ();
 sg13g2_decap_4 FILLER_69_2392 ();
 sg13g2_fill_1 FILLER_69_2396 ();
 sg13g2_decap_4 FILLER_69_2406 ();
 sg13g2_fill_1 FILLER_69_2410 ();
 sg13g2_fill_1 FILLER_69_2467 ();
 sg13g2_fill_1 FILLER_69_2473 ();
 sg13g2_fill_1 FILLER_69_2490 ();
 sg13g2_fill_1 FILLER_69_2539 ();
 sg13g2_fill_1 FILLER_69_2573 ();
 sg13g2_fill_2 FILLER_69_2587 ();
 sg13g2_fill_1 FILLER_69_2589 ();
 sg13g2_decap_4 FILLER_69_2594 ();
 sg13g2_fill_2 FILLER_69_2598 ();
 sg13g2_decap_4 FILLER_69_2606 ();
 sg13g2_fill_2 FILLER_69_2610 ();
 sg13g2_decap_4 FILLER_69_2630 ();
 sg13g2_fill_2 FILLER_69_2634 ();
 sg13g2_decap_4 FILLER_69_2666 ();
 sg13g2_fill_2 FILLER_70_50 ();
 sg13g2_fill_1 FILLER_70_89 ();
 sg13g2_fill_2 FILLER_70_115 ();
 sg13g2_fill_1 FILLER_70_163 ();
 sg13g2_fill_1 FILLER_70_204 ();
 sg13g2_fill_2 FILLER_70_240 ();
 sg13g2_fill_1 FILLER_70_254 ();
 sg13g2_fill_2 FILLER_70_286 ();
 sg13g2_fill_2 FILLER_70_345 ();
 sg13g2_fill_2 FILLER_70_360 ();
 sg13g2_fill_2 FILLER_70_405 ();
 sg13g2_fill_1 FILLER_70_463 ();
 sg13g2_decap_8 FILLER_70_541 ();
 sg13g2_decap_4 FILLER_70_548 ();
 sg13g2_fill_2 FILLER_70_552 ();
 sg13g2_fill_1 FILLER_70_599 ();
 sg13g2_fill_1 FILLER_70_629 ();
 sg13g2_fill_1 FILLER_70_651 ();
 sg13g2_fill_1 FILLER_70_663 ();
 sg13g2_fill_2 FILLER_70_674 ();
 sg13g2_fill_1 FILLER_70_768 ();
 sg13g2_fill_1 FILLER_70_785 ();
 sg13g2_fill_2 FILLER_70_798 ();
 sg13g2_fill_1 FILLER_70_800 ();
 sg13g2_fill_2 FILLER_70_820 ();
 sg13g2_fill_2 FILLER_70_855 ();
 sg13g2_fill_1 FILLER_70_872 ();
 sg13g2_fill_1 FILLER_70_878 ();
 sg13g2_fill_1 FILLER_70_895 ();
 sg13g2_decap_4 FILLER_70_949 ();
 sg13g2_decap_8 FILLER_70_958 ();
 sg13g2_decap_8 FILLER_70_965 ();
 sg13g2_fill_1 FILLER_70_972 ();
 sg13g2_fill_2 FILLER_70_999 ();
 sg13g2_fill_1 FILLER_70_1017 ();
 sg13g2_fill_2 FILLER_70_1027 ();
 sg13g2_fill_2 FILLER_70_1045 ();
 sg13g2_fill_1 FILLER_70_1055 ();
 sg13g2_fill_2 FILLER_70_1063 ();
 sg13g2_fill_1 FILLER_70_1083 ();
 sg13g2_fill_2 FILLER_70_1131 ();
 sg13g2_fill_2 FILLER_70_1192 ();
 sg13g2_fill_1 FILLER_70_1198 ();
 sg13g2_fill_2 FILLER_70_1231 ();
 sg13g2_fill_2 FILLER_70_1244 ();
 sg13g2_fill_2 FILLER_70_1269 ();
 sg13g2_fill_1 FILLER_70_1275 ();
 sg13g2_fill_1 FILLER_70_1290 ();
 sg13g2_decap_8 FILLER_70_1311 ();
 sg13g2_decap_8 FILLER_70_1318 ();
 sg13g2_decap_8 FILLER_70_1325 ();
 sg13g2_decap_4 FILLER_70_1332 ();
 sg13g2_fill_1 FILLER_70_1336 ();
 sg13g2_fill_2 FILLER_70_1378 ();
 sg13g2_decap_8 FILLER_70_1442 ();
 sg13g2_decap_8 FILLER_70_1449 ();
 sg13g2_fill_1 FILLER_70_1456 ();
 sg13g2_decap_4 FILLER_70_1466 ();
 sg13g2_fill_2 FILLER_70_1470 ();
 sg13g2_fill_2 FILLER_70_1476 ();
 sg13g2_decap_4 FILLER_70_1487 ();
 sg13g2_fill_1 FILLER_70_1504 ();
 sg13g2_decap_4 FILLER_70_1543 ();
 sg13g2_fill_2 FILLER_70_1547 ();
 sg13g2_fill_1 FILLER_70_1553 ();
 sg13g2_decap_4 FILLER_70_1575 ();
 sg13g2_fill_1 FILLER_70_1579 ();
 sg13g2_decap_8 FILLER_70_1589 ();
 sg13g2_decap_4 FILLER_70_1596 ();
 sg13g2_fill_1 FILLER_70_1600 ();
 sg13g2_decap_4 FILLER_70_1605 ();
 sg13g2_fill_2 FILLER_70_1609 ();
 sg13g2_fill_1 FILLER_70_1619 ();
 sg13g2_fill_1 FILLER_70_1628 ();
 sg13g2_fill_1 FILLER_70_1637 ();
 sg13g2_fill_2 FILLER_70_1682 ();
 sg13g2_fill_1 FILLER_70_1684 ();
 sg13g2_fill_1 FILLER_70_1722 ();
 sg13g2_fill_1 FILLER_70_1756 ();
 sg13g2_fill_2 FILLER_70_1796 ();
 sg13g2_fill_1 FILLER_70_1826 ();
 sg13g2_fill_1 FILLER_70_1831 ();
 sg13g2_fill_2 FILLER_70_1870 ();
 sg13g2_fill_1 FILLER_70_1888 ();
 sg13g2_fill_1 FILLER_70_1913 ();
 sg13g2_fill_2 FILLER_70_1935 ();
 sg13g2_fill_2 FILLER_70_1956 ();
 sg13g2_fill_1 FILLER_70_1986 ();
 sg13g2_fill_2 FILLER_70_2008 ();
 sg13g2_fill_2 FILLER_70_2019 ();
 sg13g2_fill_2 FILLER_70_2087 ();
 sg13g2_fill_2 FILLER_70_2115 ();
 sg13g2_fill_2 FILLER_70_2158 ();
 sg13g2_fill_1 FILLER_70_2171 ();
 sg13g2_fill_2 FILLER_70_2190 ();
 sg13g2_fill_2 FILLER_70_2200 ();
 sg13g2_fill_2 FILLER_70_2210 ();
 sg13g2_fill_2 FILLER_70_2246 ();
 sg13g2_fill_1 FILLER_70_2287 ();
 sg13g2_fill_1 FILLER_70_2314 ();
 sg13g2_fill_2 FILLER_70_2328 ();
 sg13g2_fill_2 FILLER_70_2352 ();
 sg13g2_fill_1 FILLER_70_2359 ();
 sg13g2_fill_2 FILLER_70_2376 ();
 sg13g2_fill_1 FILLER_70_2378 ();
 sg13g2_decap_8 FILLER_70_2394 ();
 sg13g2_decap_8 FILLER_70_2401 ();
 sg13g2_decap_8 FILLER_70_2408 ();
 sg13g2_fill_1 FILLER_70_2415 ();
 sg13g2_fill_1 FILLER_70_2460 ();
 sg13g2_fill_2 FILLER_70_2471 ();
 sg13g2_fill_2 FILLER_70_2517 ();
 sg13g2_fill_1 FILLER_70_2570 ();
 sg13g2_decap_4 FILLER_70_2578 ();
 sg13g2_fill_2 FILLER_70_2619 ();
 sg13g2_fill_1 FILLER_70_2621 ();
 sg13g2_decap_8 FILLER_70_2652 ();
 sg13g2_decap_8 FILLER_70_2659 ();
 sg13g2_decap_4 FILLER_70_2666 ();
 sg13g2_fill_2 FILLER_71_36 ();
 sg13g2_fill_1 FILLER_71_59 ();
 sg13g2_fill_2 FILLER_71_120 ();
 sg13g2_fill_1 FILLER_71_132 ();
 sg13g2_fill_1 FILLER_71_145 ();
 sg13g2_fill_2 FILLER_71_150 ();
 sg13g2_fill_2 FILLER_71_182 ();
 sg13g2_fill_1 FILLER_71_205 ();
 sg13g2_fill_2 FILLER_71_221 ();
 sg13g2_fill_2 FILLER_71_231 ();
 sg13g2_fill_1 FILLER_71_241 ();
 sg13g2_fill_1 FILLER_71_275 ();
 sg13g2_fill_2 FILLER_71_283 ();
 sg13g2_fill_2 FILLER_71_420 ();
 sg13g2_fill_1 FILLER_71_460 ();
 sg13g2_fill_1 FILLER_71_486 ();
 sg13g2_fill_1 FILLER_71_500 ();
 sg13g2_fill_2 FILLER_71_642 ();
 sg13g2_fill_1 FILLER_71_651 ();
 sg13g2_fill_2 FILLER_71_676 ();
 sg13g2_fill_1 FILLER_71_699 ();
 sg13g2_fill_1 FILLER_71_761 ();
 sg13g2_fill_1 FILLER_71_774 ();
 sg13g2_fill_2 FILLER_71_778 ();
 sg13g2_fill_1 FILLER_71_780 ();
 sg13g2_decap_4 FILLER_71_800 ();
 sg13g2_fill_2 FILLER_71_804 ();
 sg13g2_fill_1 FILLER_71_814 ();
 sg13g2_decap_4 FILLER_71_848 ();
 sg13g2_fill_1 FILLER_71_852 ();
 sg13g2_fill_2 FILLER_71_857 ();
 sg13g2_decap_4 FILLER_71_874 ();
 sg13g2_fill_2 FILLER_71_878 ();
 sg13g2_fill_2 FILLER_71_912 ();
 sg13g2_fill_2 FILLER_71_935 ();
 sg13g2_fill_1 FILLER_71_937 ();
 sg13g2_decap_4 FILLER_71_947 ();
 sg13g2_fill_2 FILLER_71_951 ();
 sg13g2_decap_8 FILLER_71_957 ();
 sg13g2_fill_2 FILLER_71_964 ();
 sg13g2_fill_1 FILLER_71_966 ();
 sg13g2_decap_8 FILLER_71_971 ();
 sg13g2_decap_4 FILLER_71_978 ();
 sg13g2_fill_2 FILLER_71_982 ();
 sg13g2_fill_2 FILLER_71_991 ();
 sg13g2_fill_1 FILLER_71_997 ();
 sg13g2_fill_1 FILLER_71_1043 ();
 sg13g2_fill_2 FILLER_71_1052 ();
 sg13g2_fill_1 FILLER_71_1104 ();
 sg13g2_fill_1 FILLER_71_1157 ();
 sg13g2_fill_2 FILLER_71_1168 ();
 sg13g2_fill_1 FILLER_71_1183 ();
 sg13g2_fill_2 FILLER_71_1217 ();
 sg13g2_fill_2 FILLER_71_1247 ();
 sg13g2_decap_8 FILLER_71_1305 ();
 sg13g2_decap_4 FILLER_71_1312 ();
 sg13g2_fill_1 FILLER_71_1316 ();
 sg13g2_decap_8 FILLER_71_1326 ();
 sg13g2_decap_8 FILLER_71_1333 ();
 sg13g2_decap_4 FILLER_71_1340 ();
 sg13g2_fill_1 FILLER_71_1344 ();
 sg13g2_fill_1 FILLER_71_1354 ();
 sg13g2_fill_1 FILLER_71_1359 ();
 sg13g2_fill_2 FILLER_71_1372 ();
 sg13g2_fill_1 FILLER_71_1427 ();
 sg13g2_decap_8 FILLER_71_1433 ();
 sg13g2_decap_4 FILLER_71_1440 ();
 sg13g2_fill_1 FILLER_71_1444 ();
 sg13g2_fill_1 FILLER_71_1505 ();
 sg13g2_fill_2 FILLER_71_1536 ();
 sg13g2_fill_1 FILLER_71_1538 ();
 sg13g2_decap_8 FILLER_71_1570 ();
 sg13g2_decap_4 FILLER_71_1607 ();
 sg13g2_decap_8 FILLER_71_1675 ();
 sg13g2_fill_2 FILLER_71_1682 ();
 sg13g2_fill_1 FILLER_71_1705 ();
 sg13g2_fill_1 FILLER_71_1721 ();
 sg13g2_fill_1 FILLER_71_1735 ();
 sg13g2_fill_1 FILLER_71_1756 ();
 sg13g2_fill_1 FILLER_71_1766 ();
 sg13g2_fill_1 FILLER_71_1801 ();
 sg13g2_fill_1 FILLER_71_1823 ();
 sg13g2_decap_4 FILLER_71_1859 ();
 sg13g2_fill_2 FILLER_71_1872 ();
 sg13g2_fill_1 FILLER_71_1874 ();
 sg13g2_fill_1 FILLER_71_1926 ();
 sg13g2_fill_1 FILLER_71_1952 ();
 sg13g2_fill_1 FILLER_71_1976 ();
 sg13g2_fill_1 FILLER_71_2126 ();
 sg13g2_fill_1 FILLER_71_2136 ();
 sg13g2_fill_2 FILLER_71_2180 ();
 sg13g2_fill_2 FILLER_71_2265 ();
 sg13g2_fill_2 FILLER_71_2327 ();
 sg13g2_fill_1 FILLER_71_2329 ();
 sg13g2_fill_1 FILLER_71_2335 ();
 sg13g2_fill_1 FILLER_71_2340 ();
 sg13g2_fill_1 FILLER_71_2360 ();
 sg13g2_fill_1 FILLER_71_2371 ();
 sg13g2_fill_2 FILLER_71_2388 ();
 sg13g2_fill_2 FILLER_71_2416 ();
 sg13g2_fill_1 FILLER_71_2467 ();
 sg13g2_fill_1 FILLER_71_2476 ();
 sg13g2_fill_1 FILLER_71_2535 ();
 sg13g2_fill_1 FILLER_71_2541 ();
 sg13g2_fill_2 FILLER_71_2610 ();
 sg13g2_fill_1 FILLER_71_2612 ();
 sg13g2_fill_1 FILLER_71_2618 ();
 sg13g2_decap_8 FILLER_71_2650 ();
 sg13g2_decap_8 FILLER_71_2657 ();
 sg13g2_decap_4 FILLER_71_2664 ();
 sg13g2_fill_2 FILLER_71_2668 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_45 ();
 sg13g2_fill_1 FILLER_72_60 ();
 sg13g2_fill_1 FILLER_72_87 ();
 sg13g2_fill_2 FILLER_72_135 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_fill_1 FILLER_72_180 ();
 sg13g2_fill_1 FILLER_72_207 ();
 sg13g2_fill_2 FILLER_72_250 ();
 sg13g2_fill_2 FILLER_72_277 ();
 sg13g2_fill_1 FILLER_72_305 ();
 sg13g2_fill_1 FILLER_72_383 ();
 sg13g2_fill_1 FILLER_72_407 ();
 sg13g2_fill_2 FILLER_72_464 ();
 sg13g2_fill_1 FILLER_72_500 ();
 sg13g2_fill_1 FILLER_72_505 ();
 sg13g2_fill_1 FILLER_72_515 ();
 sg13g2_fill_1 FILLER_72_520 ();
 sg13g2_fill_1 FILLER_72_672 ();
 sg13g2_fill_2 FILLER_72_711 ();
 sg13g2_fill_1 FILLER_72_739 ();
 sg13g2_fill_1 FILLER_72_747 ();
 sg13g2_fill_2 FILLER_72_777 ();
 sg13g2_fill_1 FILLER_72_779 ();
 sg13g2_fill_2 FILLER_72_888 ();
 sg13g2_fill_2 FILLER_72_894 ();
 sg13g2_decap_4 FILLER_72_900 ();
 sg13g2_fill_2 FILLER_72_904 ();
 sg13g2_fill_1 FILLER_72_920 ();
 sg13g2_fill_2 FILLER_72_929 ();
 sg13g2_fill_1 FILLER_72_987 ();
 sg13g2_fill_1 FILLER_72_992 ();
 sg13g2_fill_1 FILLER_72_997 ();
 sg13g2_fill_1 FILLER_72_1024 ();
 sg13g2_fill_1 FILLER_72_1030 ();
 sg13g2_fill_2 FILLER_72_1091 ();
 sg13g2_fill_1 FILLER_72_1135 ();
 sg13g2_fill_2 FILLER_72_1224 ();
 sg13g2_fill_1 FILLER_72_1313 ();
 sg13g2_fill_2 FILLER_72_1340 ();
 sg13g2_fill_1 FILLER_72_1368 ();
 sg13g2_fill_2 FILLER_72_1373 ();
 sg13g2_fill_2 FILLER_72_1417 ();
 sg13g2_fill_1 FILLER_72_1445 ();
 sg13g2_fill_1 FILLER_72_1476 ();
 sg13g2_fill_1 FILLER_72_1503 ();
 sg13g2_fill_1 FILLER_72_1508 ();
 sg13g2_decap_8 FILLER_72_1535 ();
 sg13g2_fill_2 FILLER_72_1542 ();
 sg13g2_fill_1 FILLER_72_1544 ();
 sg13g2_decap_4 FILLER_72_1571 ();
 sg13g2_fill_1 FILLER_72_1579 ();
 sg13g2_decap_4 FILLER_72_1602 ();
 sg13g2_fill_2 FILLER_72_1606 ();
 sg13g2_decap_4 FILLER_72_1612 ();
 sg13g2_fill_2 FILLER_72_1621 ();
 sg13g2_fill_1 FILLER_72_1623 ();
 sg13g2_decap_4 FILLER_72_1661 ();
 sg13g2_fill_2 FILLER_72_1693 ();
 sg13g2_fill_1 FILLER_72_1729 ();
 sg13g2_fill_2 FILLER_72_1792 ();
 sg13g2_fill_2 FILLER_72_1827 ();
 sg13g2_fill_1 FILLER_72_1829 ();
 sg13g2_decap_4 FILLER_72_1834 ();
 sg13g2_fill_2 FILLER_72_1842 ();
 sg13g2_fill_2 FILLER_72_1853 ();
 sg13g2_fill_1 FILLER_72_1885 ();
 sg13g2_fill_1 FILLER_72_1959 ();
 sg13g2_fill_1 FILLER_72_1990 ();
 sg13g2_fill_2 FILLER_72_1994 ();
 sg13g2_fill_1 FILLER_72_2079 ();
 sg13g2_fill_2 FILLER_72_2184 ();
 sg13g2_fill_1 FILLER_72_2193 ();
 sg13g2_fill_2 FILLER_72_2229 ();
 sg13g2_fill_2 FILLER_72_2239 ();
 sg13g2_fill_2 FILLER_72_2295 ();
 sg13g2_fill_1 FILLER_72_2308 ();
 sg13g2_fill_2 FILLER_72_2322 ();
 sg13g2_fill_1 FILLER_72_2328 ();
 sg13g2_fill_1 FILLER_72_2355 ();
 sg13g2_fill_1 FILLER_72_2367 ();
 sg13g2_fill_1 FILLER_72_2374 ();
 sg13g2_fill_1 FILLER_72_2463 ();
 sg13g2_fill_2 FILLER_72_2535 ();
 sg13g2_fill_2 FILLER_72_2546 ();
 sg13g2_fill_1 FILLER_72_2555 ();
 sg13g2_fill_2 FILLER_72_2585 ();
 sg13g2_fill_2 FILLER_72_2591 ();
 sg13g2_fill_2 FILLER_72_2612 ();
 sg13g2_fill_1 FILLER_72_2614 ();
 sg13g2_fill_2 FILLER_72_2635 ();
 sg13g2_decap_8 FILLER_72_2663 ();
 sg13g2_fill_1 FILLER_73_55 ();
 sg13g2_fill_2 FILLER_73_89 ();
 sg13g2_fill_2 FILLER_73_95 ();
 sg13g2_fill_1 FILLER_73_101 ();
 sg13g2_fill_1 FILLER_73_114 ();
 sg13g2_fill_2 FILLER_73_175 ();
 sg13g2_fill_2 FILLER_73_254 ();
 sg13g2_fill_2 FILLER_73_267 ();
 sg13g2_fill_2 FILLER_73_286 ();
 sg13g2_fill_2 FILLER_73_304 ();
 sg13g2_fill_2 FILLER_73_338 ();
 sg13g2_fill_2 FILLER_73_384 ();
 sg13g2_fill_2 FILLER_73_408 ();
 sg13g2_fill_1 FILLER_73_443 ();
 sg13g2_fill_2 FILLER_73_453 ();
 sg13g2_fill_2 FILLER_73_546 ();
 sg13g2_decap_4 FILLER_73_618 ();
 sg13g2_fill_1 FILLER_73_622 ();
 sg13g2_fill_1 FILLER_73_637 ();
 sg13g2_fill_1 FILLER_73_642 ();
 sg13g2_fill_1 FILLER_73_699 ();
 sg13g2_fill_1 FILLER_73_705 ();
 sg13g2_fill_1 FILLER_73_710 ();
 sg13g2_fill_2 FILLER_73_716 ();
 sg13g2_fill_2 FILLER_73_756 ();
 sg13g2_fill_2 FILLER_73_766 ();
 sg13g2_fill_2 FILLER_73_808 ();
 sg13g2_fill_2 FILLER_73_856 ();
 sg13g2_fill_1 FILLER_73_858 ();
 sg13g2_fill_1 FILLER_73_872 ();
 sg13g2_decap_8 FILLER_73_899 ();
 sg13g2_decap_4 FILLER_73_906 ();
 sg13g2_fill_2 FILLER_73_910 ();
 sg13g2_fill_2 FILLER_73_933 ();
 sg13g2_fill_1 FILLER_73_935 ();
 sg13g2_fill_1 FILLER_73_988 ();
 sg13g2_fill_2 FILLER_73_1071 ();
 sg13g2_fill_1 FILLER_73_1108 ();
 sg13g2_fill_2 FILLER_73_1139 ();
 sg13g2_fill_2 FILLER_73_1154 ();
 sg13g2_fill_1 FILLER_73_1161 ();
 sg13g2_fill_2 FILLER_73_1169 ();
 sg13g2_fill_1 FILLER_73_1176 ();
 sg13g2_fill_1 FILLER_73_1185 ();
 sg13g2_fill_2 FILLER_73_1200 ();
 sg13g2_fill_2 FILLER_73_1206 ();
 sg13g2_fill_1 FILLER_73_1248 ();
 sg13g2_fill_1 FILLER_73_1322 ();
 sg13g2_decap_8 FILLER_73_1327 ();
 sg13g2_decap_4 FILLER_73_1334 ();
 sg13g2_fill_1 FILLER_73_1338 ();
 sg13g2_decap_4 FILLER_73_1343 ();
 sg13g2_fill_2 FILLER_73_1355 ();
 sg13g2_decap_8 FILLER_73_1361 ();
 sg13g2_decap_4 FILLER_73_1407 ();
 sg13g2_fill_2 FILLER_73_1445 ();
 sg13g2_fill_1 FILLER_73_1447 ();
 sg13g2_fill_2 FILLER_73_1470 ();
 sg13g2_fill_1 FILLER_73_1472 ();
 sg13g2_fill_2 FILLER_73_1507 ();
 sg13g2_fill_2 FILLER_73_1514 ();
 sg13g2_fill_1 FILLER_73_1516 ();
 sg13g2_fill_1 FILLER_73_1538 ();
 sg13g2_decap_4 FILLER_73_1556 ();
 sg13g2_fill_1 FILLER_73_1560 ();
 sg13g2_decap_4 FILLER_73_1569 ();
 sg13g2_fill_1 FILLER_73_1590 ();
 sg13g2_fill_2 FILLER_73_1628 ();
 sg13g2_fill_1 FILLER_73_1646 ();
 sg13g2_decap_8 FILLER_73_1668 ();
 sg13g2_fill_2 FILLER_73_1675 ();
 sg13g2_fill_1 FILLER_73_1677 ();
 sg13g2_fill_1 FILLER_73_1744 ();
 sg13g2_fill_2 FILLER_73_1749 ();
 sg13g2_fill_1 FILLER_73_1756 ();
 sg13g2_decap_4 FILLER_73_1796 ();
 sg13g2_decap_8 FILLER_73_1830 ();
 sg13g2_decap_8 FILLER_73_1837 ();
 sg13g2_fill_2 FILLER_73_1844 ();
 sg13g2_fill_1 FILLER_73_1846 ();
 sg13g2_fill_2 FILLER_73_1865 ();
 sg13g2_fill_1 FILLER_73_1931 ();
 sg13g2_fill_1 FILLER_73_1937 ();
 sg13g2_fill_1 FILLER_73_1964 ();
 sg13g2_fill_2 FILLER_73_1970 ();
 sg13g2_fill_2 FILLER_73_1976 ();
 sg13g2_fill_1 FILLER_73_1978 ();
 sg13g2_fill_2 FILLER_73_1984 ();
 sg13g2_fill_1 FILLER_73_2023 ();
 sg13g2_fill_1 FILLER_73_2053 ();
 sg13g2_fill_2 FILLER_73_2120 ();
 sg13g2_fill_2 FILLER_73_2137 ();
 sg13g2_fill_1 FILLER_73_2175 ();
 sg13g2_fill_2 FILLER_73_2183 ();
 sg13g2_fill_2 FILLER_73_2193 ();
 sg13g2_fill_2 FILLER_73_2205 ();
 sg13g2_fill_1 FILLER_73_2229 ();
 sg13g2_fill_2 FILLER_73_2247 ();
 sg13g2_fill_1 FILLER_73_2253 ();
 sg13g2_fill_2 FILLER_73_2265 ();
 sg13g2_fill_2 FILLER_73_2329 ();
 sg13g2_fill_1 FILLER_73_2331 ();
 sg13g2_fill_2 FILLER_73_2369 ();
 sg13g2_fill_2 FILLER_73_2376 ();
 sg13g2_fill_1 FILLER_73_2382 ();
 sg13g2_fill_2 FILLER_73_2387 ();
 sg13g2_fill_1 FILLER_73_2389 ();
 sg13g2_fill_2 FILLER_73_2395 ();
 sg13g2_fill_1 FILLER_73_2397 ();
 sg13g2_fill_1 FILLER_73_2403 ();
 sg13g2_fill_1 FILLER_73_2415 ();
 sg13g2_fill_2 FILLER_73_2427 ();
 sg13g2_fill_2 FILLER_73_2472 ();
 sg13g2_fill_2 FILLER_73_2542 ();
 sg13g2_fill_1 FILLER_73_2555 ();
 sg13g2_fill_1 FILLER_73_2566 ();
 sg13g2_decap_8 FILLER_73_2576 ();
 sg13g2_decap_8 FILLER_73_2583 ();
 sg13g2_fill_2 FILLER_73_2590 ();
 sg13g2_fill_1 FILLER_73_2592 ();
 sg13g2_decap_4 FILLER_73_2614 ();
 sg13g2_decap_8 FILLER_73_2648 ();
 sg13g2_decap_8 FILLER_73_2655 ();
 sg13g2_decap_8 FILLER_73_2662 ();
 sg13g2_fill_1 FILLER_73_2669 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_22 ();
 sg13g2_fill_1 FILLER_74_88 ();
 sg13g2_fill_1 FILLER_74_184 ();
 sg13g2_fill_1 FILLER_74_194 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_fill_2 FILLER_74_220 ();
 sg13g2_fill_1 FILLER_74_241 ();
 sg13g2_fill_1 FILLER_74_250 ();
 sg13g2_fill_2 FILLER_74_340 ();
 sg13g2_fill_2 FILLER_74_355 ();
 sg13g2_fill_1 FILLER_74_373 ();
 sg13g2_fill_1 FILLER_74_382 ();
 sg13g2_fill_1 FILLER_74_386 ();
 sg13g2_fill_1 FILLER_74_404 ();
 sg13g2_fill_2 FILLER_74_408 ();
 sg13g2_fill_1 FILLER_74_515 ();
 sg13g2_fill_2 FILLER_74_521 ();
 sg13g2_decap_4 FILLER_74_527 ();
 sg13g2_decap_8 FILLER_74_535 ();
 sg13g2_decap_4 FILLER_74_542 ();
 sg13g2_fill_2 FILLER_74_546 ();
 sg13g2_decap_4 FILLER_74_553 ();
 sg13g2_fill_1 FILLER_74_557 ();
 sg13g2_fill_1 FILLER_74_562 ();
 sg13g2_fill_2 FILLER_74_580 ();
 sg13g2_fill_1 FILLER_74_586 ();
 sg13g2_decap_8 FILLER_74_617 ();
 sg13g2_decap_4 FILLER_74_624 ();
 sg13g2_fill_1 FILLER_74_674 ();
 sg13g2_fill_1 FILLER_74_679 ();
 sg13g2_fill_2 FILLER_74_749 ();
 sg13g2_fill_1 FILLER_74_751 ();
 sg13g2_fill_1 FILLER_74_778 ();
 sg13g2_fill_2 FILLER_74_796 ();
 sg13g2_fill_1 FILLER_74_798 ();
 sg13g2_fill_1 FILLER_74_825 ();
 sg13g2_fill_2 FILLER_74_830 ();
 sg13g2_fill_1 FILLER_74_832 ();
 sg13g2_fill_2 FILLER_74_838 ();
 sg13g2_fill_1 FILLER_74_840 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_fill_2 FILLER_74_852 ();
 sg13g2_fill_1 FILLER_74_854 ();
 sg13g2_fill_1 FILLER_74_889 ();
 sg13g2_fill_1 FILLER_74_894 ();
 sg13g2_fill_1 FILLER_74_903 ();
 sg13g2_fill_1 FILLER_74_930 ();
 sg13g2_fill_1 FILLER_74_940 ();
 sg13g2_fill_2 FILLER_74_962 ();
 sg13g2_fill_1 FILLER_74_964 ();
 sg13g2_fill_1 FILLER_74_970 ();
 sg13g2_fill_2 FILLER_74_975 ();
 sg13g2_fill_1 FILLER_74_989 ();
 sg13g2_fill_1 FILLER_74_995 ();
 sg13g2_fill_1 FILLER_74_1001 ();
 sg13g2_fill_2 FILLER_74_1006 ();
 sg13g2_fill_1 FILLER_74_1012 ();
 sg13g2_fill_2 FILLER_74_1050 ();
 sg13g2_fill_1 FILLER_74_1060 ();
 sg13g2_fill_1 FILLER_74_1095 ();
 sg13g2_fill_1 FILLER_74_1100 ();
 sg13g2_fill_1 FILLER_74_1105 ();
 sg13g2_fill_1 FILLER_74_1111 ();
 sg13g2_fill_1 FILLER_74_1116 ();
 sg13g2_fill_1 FILLER_74_1121 ();
 sg13g2_fill_2 FILLER_74_1126 ();
 sg13g2_fill_2 FILLER_74_1208 ();
 sg13g2_fill_2 FILLER_74_1248 ();
 sg13g2_fill_2 FILLER_74_1296 ();
 sg13g2_fill_1 FILLER_74_1298 ();
 sg13g2_fill_2 FILLER_74_1303 ();
 sg13g2_fill_2 FILLER_74_1309 ();
 sg13g2_fill_2 FILLER_74_1337 ();
 sg13g2_fill_1 FILLER_74_1339 ();
 sg13g2_decap_8 FILLER_74_1345 ();
 sg13g2_decap_8 FILLER_74_1352 ();
 sg13g2_decap_8 FILLER_74_1359 ();
 sg13g2_decap_8 FILLER_74_1366 ();
 sg13g2_decap_4 FILLER_74_1373 ();
 sg13g2_fill_1 FILLER_74_1377 ();
 sg13g2_fill_2 FILLER_74_1383 ();
 sg13g2_fill_1 FILLER_74_1410 ();
 sg13g2_fill_1 FILLER_74_1428 ();
 sg13g2_decap_4 FILLER_74_1459 ();
 sg13g2_fill_2 FILLER_74_1463 ();
 sg13g2_fill_2 FILLER_74_1490 ();
 sg13g2_fill_1 FILLER_74_1492 ();
 sg13g2_fill_2 FILLER_74_1514 ();
 sg13g2_fill_1 FILLER_74_1516 ();
 sg13g2_decap_8 FILLER_74_1525 ();
 sg13g2_fill_2 FILLER_74_1532 ();
 sg13g2_decap_8 FILLER_74_1543 ();
 sg13g2_decap_4 FILLER_74_1550 ();
 sg13g2_fill_1 FILLER_74_1585 ();
 sg13g2_decap_8 FILLER_74_1616 ();
 sg13g2_decap_4 FILLER_74_1623 ();
 sg13g2_fill_2 FILLER_74_1738 ();
 sg13g2_decap_4 FILLER_74_1802 ();
 sg13g2_fill_1 FILLER_74_1806 ();
 sg13g2_decap_8 FILLER_74_1824 ();
 sg13g2_decap_4 FILLER_74_1831 ();
 sg13g2_fill_1 FILLER_74_1835 ();
 sg13g2_fill_2 FILLER_74_1845 ();
 sg13g2_fill_1 FILLER_74_1847 ();
 sg13g2_fill_1 FILLER_74_1882 ();
 sg13g2_fill_1 FILLER_74_1909 ();
 sg13g2_fill_1 FILLER_74_1915 ();
 sg13g2_fill_2 FILLER_74_1921 ();
 sg13g2_decap_8 FILLER_74_1968 ();
 sg13g2_decap_8 FILLER_74_1984 ();
 sg13g2_decap_4 FILLER_74_1991 ();
 sg13g2_fill_2 FILLER_74_1995 ();
 sg13g2_fill_2 FILLER_74_2126 ();
 sg13g2_fill_1 FILLER_74_2216 ();
 sg13g2_fill_1 FILLER_74_2229 ();
 sg13g2_fill_1 FILLER_74_2265 ();
 sg13g2_fill_2 FILLER_74_2271 ();
 sg13g2_fill_2 FILLER_74_2328 ();
 sg13g2_fill_1 FILLER_74_2334 ();
 sg13g2_fill_2 FILLER_74_2343 ();
 sg13g2_decap_8 FILLER_74_2350 ();
 sg13g2_decap_8 FILLER_74_2357 ();
 sg13g2_decap_8 FILLER_74_2364 ();
 sg13g2_fill_1 FILLER_74_2371 ();
 sg13g2_decap_4 FILLER_74_2376 ();
 sg13g2_decap_4 FILLER_74_2396 ();
 sg13g2_fill_2 FILLER_74_2400 ();
 sg13g2_fill_1 FILLER_74_2411 ();
 sg13g2_fill_1 FILLER_74_2436 ();
 sg13g2_fill_2 FILLER_74_2450 ();
 sg13g2_fill_1 FILLER_74_2474 ();
 sg13g2_fill_2 FILLER_74_2500 ();
 sg13g2_fill_2 FILLER_74_2529 ();
 sg13g2_decap_8 FILLER_74_2561 ();
 sg13g2_decap_4 FILLER_74_2568 ();
 sg13g2_decap_8 FILLER_74_2619 ();
 sg13g2_decap_8 FILLER_74_2626 ();
 sg13g2_decap_8 FILLER_74_2633 ();
 sg13g2_decap_8 FILLER_74_2644 ();
 sg13g2_decap_8 FILLER_74_2651 ();
 sg13g2_decap_8 FILLER_74_2658 ();
 sg13g2_decap_4 FILLER_74_2665 ();
 sg13g2_fill_1 FILLER_74_2669 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_107 ();
 sg13g2_fill_1 FILLER_75_121 ();
 sg13g2_fill_1 FILLER_75_127 ();
 sg13g2_fill_2 FILLER_75_133 ();
 sg13g2_fill_2 FILLER_75_160 ();
 sg13g2_fill_1 FILLER_75_197 ();
 sg13g2_fill_2 FILLER_75_217 ();
 sg13g2_fill_2 FILLER_75_281 ();
 sg13g2_fill_2 FILLER_75_414 ();
 sg13g2_fill_2 FILLER_75_420 ();
 sg13g2_fill_2 FILLER_75_520 ();
 sg13g2_fill_1 FILLER_75_526 ();
 sg13g2_decap_8 FILLER_75_535 ();
 sg13g2_fill_2 FILLER_75_546 ();
 sg13g2_fill_1 FILLER_75_552 ();
 sg13g2_decap_4 FILLER_75_566 ();
 sg13g2_fill_2 FILLER_75_570 ();
 sg13g2_fill_1 FILLER_75_608 ();
 sg13g2_fill_2 FILLER_75_613 ();
 sg13g2_fill_2 FILLER_75_619 ();
 sg13g2_fill_1 FILLER_75_626 ();
 sg13g2_fill_1 FILLER_75_648 ();
 sg13g2_fill_2 FILLER_75_655 ();
 sg13g2_fill_1 FILLER_75_682 ();
 sg13g2_fill_1 FILLER_75_687 ();
 sg13g2_fill_1 FILLER_75_702 ();
 sg13g2_decap_8 FILLER_75_711 ();
 sg13g2_fill_1 FILLER_75_747 ();
 sg13g2_decap_8 FILLER_75_752 ();
 sg13g2_decap_4 FILLER_75_763 ();
 sg13g2_fill_1 FILLER_75_779 ();
 sg13g2_decap_8 FILLER_75_784 ();
 sg13g2_fill_2 FILLER_75_791 ();
 sg13g2_fill_1 FILLER_75_798 ();
 sg13g2_fill_2 FILLER_75_803 ();
 sg13g2_fill_1 FILLER_75_809 ();
 sg13g2_fill_2 FILLER_75_814 ();
 sg13g2_fill_1 FILLER_75_816 ();
 sg13g2_fill_2 FILLER_75_821 ();
 sg13g2_fill_1 FILLER_75_823 ();
 sg13g2_fill_1 FILLER_75_855 ();
 sg13g2_fill_2 FILLER_75_877 ();
 sg13g2_fill_2 FILLER_75_884 ();
 sg13g2_fill_1 FILLER_75_904 ();
 sg13g2_fill_1 FILLER_75_909 ();
 sg13g2_fill_2 FILLER_75_914 ();
 sg13g2_fill_2 FILLER_75_920 ();
 sg13g2_fill_2 FILLER_75_926 ();
 sg13g2_fill_2 FILLER_75_948 ();
 sg13g2_fill_1 FILLER_75_958 ();
 sg13g2_decap_8 FILLER_75_964 ();
 sg13g2_decap_8 FILLER_75_971 ();
 sg13g2_decap_4 FILLER_75_978 ();
 sg13g2_fill_2 FILLER_75_1003 ();
 sg13g2_fill_1 FILLER_75_1009 ();
 sg13g2_fill_1 FILLER_75_1014 ();
 sg13g2_fill_1 FILLER_75_1019 ();
 sg13g2_fill_1 FILLER_75_1039 ();
 sg13g2_fill_2 FILLER_75_1048 ();
 sg13g2_fill_1 FILLER_75_1081 ();
 sg13g2_fill_1 FILLER_75_1097 ();
 sg13g2_fill_1 FILLER_75_1111 ();
 sg13g2_fill_1 FILLER_75_1120 ();
 sg13g2_decap_8 FILLER_75_1126 ();
 sg13g2_fill_2 FILLER_75_1133 ();
 sg13g2_fill_1 FILLER_75_1135 ();
 sg13g2_fill_2 FILLER_75_1146 ();
 sg13g2_fill_1 FILLER_75_1169 ();
 sg13g2_fill_2 FILLER_75_1182 ();
 sg13g2_fill_2 FILLER_75_1197 ();
 sg13g2_fill_1 FILLER_75_1202 ();
 sg13g2_fill_1 FILLER_75_1215 ();
 sg13g2_fill_1 FILLER_75_1261 ();
 sg13g2_fill_1 FILLER_75_1266 ();
 sg13g2_decap_8 FILLER_75_1274 ();
 sg13g2_decap_8 FILLER_75_1281 ();
 sg13g2_decap_4 FILLER_75_1296 ();
 sg13g2_fill_1 FILLER_75_1300 ();
 sg13g2_fill_1 FILLER_75_1318 ();
 sg13g2_decap_8 FILLER_75_1323 ();
 sg13g2_fill_2 FILLER_75_1330 ();
 sg13g2_decap_8 FILLER_75_1341 ();
 sg13g2_fill_1 FILLER_75_1348 ();
 sg13g2_decap_4 FILLER_75_1379 ();
 sg13g2_fill_1 FILLER_75_1383 ();
 sg13g2_decap_8 FILLER_75_1388 ();
 sg13g2_decap_4 FILLER_75_1429 ();
 sg13g2_fill_1 FILLER_75_1433 ();
 sg13g2_decap_8 FILLER_75_1438 ();
 sg13g2_fill_2 FILLER_75_1445 ();
 sg13g2_fill_1 FILLER_75_1447 ();
 sg13g2_decap_4 FILLER_75_1465 ();
 sg13g2_fill_2 FILLER_75_1512 ();
 sg13g2_fill_1 FILLER_75_1535 ();
 sg13g2_fill_2 FILLER_75_1540 ();
 sg13g2_decap_8 FILLER_75_1546 ();
 sg13g2_decap_8 FILLER_75_1553 ();
 sg13g2_decap_4 FILLER_75_1560 ();
 sg13g2_fill_1 FILLER_75_1564 ();
 sg13g2_decap_4 FILLER_75_1572 ();
 sg13g2_fill_2 FILLER_75_1576 ();
 sg13g2_decap_8 FILLER_75_1582 ();
 sg13g2_fill_1 FILLER_75_1589 ();
 sg13g2_decap_4 FILLER_75_1611 ();
 sg13g2_decap_8 FILLER_75_1660 ();
 sg13g2_decap_8 FILLER_75_1667 ();
 sg13g2_decap_4 FILLER_75_1674 ();
 sg13g2_fill_2 FILLER_75_1678 ();
 sg13g2_fill_1 FILLER_75_1687 ();
 sg13g2_fill_2 FILLER_75_1736 ();
 sg13g2_fill_1 FILLER_75_1741 ();
 sg13g2_fill_1 FILLER_75_1755 ();
 sg13g2_fill_2 FILLER_75_1798 ();
 sg13g2_decap_8 FILLER_75_1804 ();
 sg13g2_fill_2 FILLER_75_1811 ();
 sg13g2_fill_1 FILLER_75_1813 ();
 sg13g2_decap_4 FILLER_75_1819 ();
 sg13g2_fill_2 FILLER_75_1823 ();
 sg13g2_decap_4 FILLER_75_1859 ();
 sg13g2_fill_2 FILLER_75_1875 ();
 sg13g2_fill_1 FILLER_75_1877 ();
 sg13g2_fill_2 FILLER_75_1896 ();
 sg13g2_decap_4 FILLER_75_1906 ();
 sg13g2_fill_2 FILLER_75_1910 ();
 sg13g2_decap_4 FILLER_75_1921 ();
 sg13g2_fill_1 FILLER_75_1925 ();
 sg13g2_fill_2 FILLER_75_1942 ();
 sg13g2_decap_8 FILLER_75_1958 ();
 sg13g2_decap_4 FILLER_75_1965 ();
 sg13g2_decap_4 FILLER_75_1999 ();
 sg13g2_fill_1 FILLER_75_2003 ();
 sg13g2_fill_1 FILLER_75_2039 ();
 sg13g2_fill_2 FILLER_75_2059 ();
 sg13g2_fill_1 FILLER_75_2074 ();
 sg13g2_fill_2 FILLER_75_2127 ();
 sg13g2_fill_2 FILLER_75_2135 ();
 sg13g2_fill_1 FILLER_75_2188 ();
 sg13g2_fill_1 FILLER_75_2194 ();
 sg13g2_fill_2 FILLER_75_2218 ();
 sg13g2_fill_1 FILLER_75_2241 ();
 sg13g2_fill_1 FILLER_75_2248 ();
 sg13g2_fill_1 FILLER_75_2300 ();
 sg13g2_fill_2 FILLER_75_2327 ();
 sg13g2_decap_8 FILLER_75_2351 ();
 sg13g2_fill_2 FILLER_75_2358 ();
 sg13g2_decap_4 FILLER_75_2364 ();
 sg13g2_fill_1 FILLER_75_2396 ();
 sg13g2_decap_4 FILLER_75_2438 ();
 sg13g2_fill_1 FILLER_75_2513 ();
 sg13g2_fill_2 FILLER_75_2531 ();
 sg13g2_decap_8 FILLER_75_2587 ();
 sg13g2_decap_4 FILLER_75_2600 ();
 sg13g2_decap_8 FILLER_75_2630 ();
 sg13g2_decap_8 FILLER_75_2637 ();
 sg13g2_decap_8 FILLER_75_2644 ();
 sg13g2_decap_8 FILLER_75_2651 ();
 sg13g2_decap_8 FILLER_75_2658 ();
 sg13g2_decap_4 FILLER_75_2665 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_51 ();
 sg13g2_fill_1 FILLER_76_78 ();
 sg13g2_fill_2 FILLER_76_108 ();
 sg13g2_fill_2 FILLER_76_179 ();
 sg13g2_fill_1 FILLER_76_209 ();
 sg13g2_fill_2 FILLER_76_216 ();
 sg13g2_fill_1 FILLER_76_250 ();
 sg13g2_fill_1 FILLER_76_291 ();
 sg13g2_fill_1 FILLER_76_303 ();
 sg13g2_fill_1 FILLER_76_320 ();
 sg13g2_fill_2 FILLER_76_351 ();
 sg13g2_fill_1 FILLER_76_407 ();
 sg13g2_fill_2 FILLER_76_445 ();
 sg13g2_fill_1 FILLER_76_471 ();
 sg13g2_fill_2 FILLER_76_495 ();
 sg13g2_fill_2 FILLER_76_506 ();
 sg13g2_fill_1 FILLER_76_512 ();
 sg13g2_fill_2 FILLER_76_580 ();
 sg13g2_fill_1 FILLER_76_582 ();
 sg13g2_fill_1 FILLER_76_592 ();
 sg13g2_fill_1 FILLER_76_598 ();
 sg13g2_fill_2 FILLER_76_633 ();
 sg13g2_fill_1 FILLER_76_668 ();
 sg13g2_fill_1 FILLER_76_673 ();
 sg13g2_fill_2 FILLER_76_678 ();
 sg13g2_fill_2 FILLER_76_685 ();
 sg13g2_fill_2 FILLER_76_693 ();
 sg13g2_fill_1 FILLER_76_695 ();
 sg13g2_fill_1 FILLER_76_705 ();
 sg13g2_fill_2 FILLER_76_715 ();
 sg13g2_fill_1 FILLER_76_717 ();
 sg13g2_decap_8 FILLER_76_743 ();
 sg13g2_decap_8 FILLER_76_750 ();
 sg13g2_decap_4 FILLER_76_757 ();
 sg13g2_decap_8 FILLER_76_779 ();
 sg13g2_fill_1 FILLER_76_808 ();
 sg13g2_fill_1 FILLER_76_813 ();
 sg13g2_fill_1 FILLER_76_839 ();
 sg13g2_decap_8 FILLER_76_844 ();
 sg13g2_fill_2 FILLER_76_851 ();
 sg13g2_fill_2 FILLER_76_897 ();
 sg13g2_fill_1 FILLER_76_899 ();
 sg13g2_fill_1 FILLER_76_909 ();
 sg13g2_fill_1 FILLER_76_931 ();
 sg13g2_fill_1 FILLER_76_942 ();
 sg13g2_decap_8 FILLER_76_965 ();
 sg13g2_decap_8 FILLER_76_972 ();
 sg13g2_fill_2 FILLER_76_979 ();
 sg13g2_fill_2 FILLER_76_986 ();
 sg13g2_fill_1 FILLER_76_988 ();
 sg13g2_fill_2 FILLER_76_1023 ();
 sg13g2_fill_1 FILLER_76_1035 ();
 sg13g2_fill_1 FILLER_76_1062 ();
 sg13g2_fill_2 FILLER_76_1112 ();
 sg13g2_fill_1 FILLER_76_1139 ();
 sg13g2_fill_1 FILLER_76_1144 ();
 sg13g2_fill_1 FILLER_76_1185 ();
 sg13g2_fill_1 FILLER_76_1255 ();
 sg13g2_fill_2 FILLER_76_1273 ();
 sg13g2_decap_8 FILLER_76_1318 ();
 sg13g2_decap_4 FILLER_76_1325 ();
 sg13g2_fill_2 FILLER_76_1329 ();
 sg13g2_decap_4 FILLER_76_1361 ();
 sg13g2_fill_1 FILLER_76_1365 ();
 sg13g2_fill_1 FILLER_76_1392 ();
 sg13g2_decap_8 FILLER_76_1423 ();
 sg13g2_decap_8 FILLER_76_1430 ();
 sg13g2_decap_4 FILLER_76_1437 ();
 sg13g2_fill_2 FILLER_76_1441 ();
 sg13g2_fill_1 FILLER_76_1478 ();
 sg13g2_fill_2 FILLER_76_1496 ();
 sg13g2_fill_1 FILLER_76_1498 ();
 sg13g2_fill_1 FILLER_76_1565 ();
 sg13g2_fill_2 FILLER_76_1578 ();
 sg13g2_fill_1 FILLER_76_1580 ();
 sg13g2_fill_1 FILLER_76_1609 ();
 sg13g2_fill_1 FILLER_76_1713 ();
 sg13g2_decap_4 FILLER_76_1830 ();
 sg13g2_fill_1 FILLER_76_1851 ();
 sg13g2_fill_2 FILLER_76_1861 ();
 sg13g2_fill_2 FILLER_76_1894 ();
 sg13g2_fill_1 FILLER_76_1896 ();
 sg13g2_fill_2 FILLER_76_1906 ();
 sg13g2_fill_2 FILLER_76_1912 ();
 sg13g2_fill_1 FILLER_76_1914 ();
 sg13g2_decap_8 FILLER_76_1945 ();
 sg13g2_fill_1 FILLER_76_1978 ();
 sg13g2_fill_2 FILLER_76_2000 ();
 sg13g2_fill_2 FILLER_76_2010 ();
 sg13g2_fill_1 FILLER_76_2012 ();
 sg13g2_fill_1 FILLER_76_2017 ();
 sg13g2_fill_1 FILLER_76_2065 ();
 sg13g2_fill_2 FILLER_76_2101 ();
 sg13g2_fill_1 FILLER_76_2136 ();
 sg13g2_fill_1 FILLER_76_2227 ();
 sg13g2_fill_1 FILLER_76_2235 ();
 sg13g2_fill_1 FILLER_76_2240 ();
 sg13g2_fill_1 FILLER_76_2273 ();
 sg13g2_fill_1 FILLER_76_2313 ();
 sg13g2_fill_2 FILLER_76_2345 ();
 sg13g2_decap_4 FILLER_76_2373 ();
 sg13g2_decap_4 FILLER_76_2385 ();
 sg13g2_fill_2 FILLER_76_2431 ();
 sg13g2_decap_8 FILLER_76_2438 ();
 sg13g2_decap_8 FILLER_76_2445 ();
 sg13g2_fill_2 FILLER_76_2470 ();
 sg13g2_fill_1 FILLER_76_2478 ();
 sg13g2_fill_1 FILLER_76_2535 ();
 sg13g2_fill_2 FILLER_76_2550 ();
 sg13g2_fill_1 FILLER_76_2552 ();
 sg13g2_fill_1 FILLER_76_2558 ();
 sg13g2_fill_1 FILLER_76_2567 ();
 sg13g2_fill_1 FILLER_76_2573 ();
 sg13g2_fill_2 FILLER_76_2579 ();
 sg13g2_decap_8 FILLER_76_2637 ();
 sg13g2_decap_8 FILLER_76_2644 ();
 sg13g2_decap_8 FILLER_76_2651 ();
 sg13g2_decap_8 FILLER_76_2658 ();
 sg13g2_decap_4 FILLER_76_2665 ();
 sg13g2_fill_1 FILLER_76_2669 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_24 ();
 sg13g2_fill_1 FILLER_77_95 ();
 sg13g2_fill_2 FILLER_77_122 ();
 sg13g2_fill_2 FILLER_77_136 ();
 sg13g2_fill_1 FILLER_77_146 ();
 sg13g2_fill_2 FILLER_77_158 ();
 sg13g2_fill_2 FILLER_77_168 ();
 sg13g2_fill_1 FILLER_77_226 ();
 sg13g2_fill_1 FILLER_77_269 ();
 sg13g2_fill_1 FILLER_77_334 ();
 sg13g2_fill_1 FILLER_77_405 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_fill_1 FILLER_77_484 ();
 sg13g2_fill_2 FILLER_77_499 ();
 sg13g2_fill_1 FILLER_77_581 ();
 sg13g2_fill_1 FILLER_77_638 ();
 sg13g2_fill_2 FILLER_77_646 ();
 sg13g2_fill_2 FILLER_77_700 ();
 sg13g2_fill_1 FILLER_77_702 ();
 sg13g2_decap_8 FILLER_77_734 ();
 sg13g2_decap_4 FILLER_77_741 ();
 sg13g2_fill_2 FILLER_77_745 ();
 sg13g2_fill_1 FILLER_77_773 ();
 sg13g2_fill_1 FILLER_77_779 ();
 sg13g2_fill_1 FILLER_77_785 ();
 sg13g2_fill_1 FILLER_77_816 ();
 sg13g2_fill_1 FILLER_77_821 ();
 sg13g2_fill_1 FILLER_77_826 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_fill_2 FILLER_77_866 ();
 sg13g2_fill_2 FILLER_77_899 ();
 sg13g2_fill_1 FILLER_77_985 ();
 sg13g2_fill_1 FILLER_77_991 ();
 sg13g2_fill_1 FILLER_77_1018 ();
 sg13g2_fill_2 FILLER_77_1070 ();
 sg13g2_fill_1 FILLER_77_1091 ();
 sg13g2_fill_2 FILLER_77_1173 ();
 sg13g2_fill_2 FILLER_77_1179 ();
 sg13g2_fill_1 FILLER_77_1207 ();
 sg13g2_fill_1 FILLER_77_1250 ();
 sg13g2_fill_1 FILLER_77_1338 ();
 sg13g2_fill_1 FILLER_77_1343 ();
 sg13g2_fill_1 FILLER_77_1370 ();
 sg13g2_fill_2 FILLER_77_1396 ();
 sg13g2_fill_1 FILLER_77_1398 ();
 sg13g2_fill_2 FILLER_77_1403 ();
 sg13g2_decap_8 FILLER_77_1426 ();
 sg13g2_decap_4 FILLER_77_1433 ();
 sg13g2_fill_2 FILLER_77_1437 ();
 sg13g2_fill_2 FILLER_77_1469 ();
 sg13g2_fill_2 FILLER_77_1480 ();
 sg13g2_fill_1 FILLER_77_1482 ();
 sg13g2_fill_1 FILLER_77_1514 ();
 sg13g2_fill_1 FILLER_77_1544 ();
 sg13g2_fill_1 FILLER_77_1549 ();
 sg13g2_decap_8 FILLER_77_1555 ();
 sg13g2_fill_2 FILLER_77_1566 ();
 sg13g2_fill_1 FILLER_77_1568 ();
 sg13g2_fill_2 FILLER_77_1573 ();
 sg13g2_fill_1 FILLER_77_1575 ();
 sg13g2_fill_2 FILLER_77_1602 ();
 sg13g2_fill_2 FILLER_77_1630 ();
 sg13g2_fill_2 FILLER_77_1661 ();
 sg13g2_fill_1 FILLER_77_1663 ();
 sg13g2_fill_2 FILLER_77_1685 ();
 sg13g2_fill_1 FILLER_77_1713 ();
 sg13g2_fill_2 FILLER_77_1761 ();
 sg13g2_fill_1 FILLER_77_1798 ();
 sg13g2_decap_4 FILLER_77_1875 ();
 sg13g2_fill_2 FILLER_77_1883 ();
 sg13g2_fill_2 FILLER_77_1889 ();
 sg13g2_decap_4 FILLER_77_1895 ();
 sg13g2_fill_1 FILLER_77_1925 ();
 sg13g2_fill_2 FILLER_77_1930 ();
 sg13g2_fill_1 FILLER_77_1932 ();
 sg13g2_fill_1 FILLER_77_1937 ();
 sg13g2_fill_1 FILLER_77_1964 ();
 sg13g2_fill_2 FILLER_77_1999 ();
 sg13g2_fill_1 FILLER_77_2005 ();
 sg13g2_fill_1 FILLER_77_2049 ();
 sg13g2_fill_2 FILLER_77_2058 ();
 sg13g2_fill_2 FILLER_77_2113 ();
 sg13g2_fill_1 FILLER_77_2140 ();
 sg13g2_fill_1 FILLER_77_2172 ();
 sg13g2_fill_1 FILLER_77_2244 ();
 sg13g2_fill_1 FILLER_77_2384 ();
 sg13g2_fill_1 FILLER_77_2409 ();
 sg13g2_decap_8 FILLER_77_2440 ();
 sg13g2_fill_2 FILLER_77_2447 ();
 sg13g2_fill_1 FILLER_77_2449 ();
 sg13g2_fill_1 FILLER_77_2471 ();
 sg13g2_fill_2 FILLER_77_2484 ();
 sg13g2_decap_4 FILLER_77_2542 ();
 sg13g2_fill_2 FILLER_77_2598 ();
 sg13g2_decap_8 FILLER_77_2605 ();
 sg13g2_decap_8 FILLER_77_2612 ();
 sg13g2_decap_8 FILLER_77_2619 ();
 sg13g2_decap_8 FILLER_77_2626 ();
 sg13g2_decap_8 FILLER_77_2633 ();
 sg13g2_decap_8 FILLER_77_2640 ();
 sg13g2_decap_8 FILLER_77_2647 ();
 sg13g2_decap_8 FILLER_77_2654 ();
 sg13g2_decap_8 FILLER_77_2661 ();
 sg13g2_fill_2 FILLER_77_2668 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_178 ();
 sg13g2_fill_1 FILLER_78_243 ();
 sg13g2_fill_1 FILLER_78_279 ();
 sg13g2_fill_1 FILLER_78_324 ();
 sg13g2_fill_1 FILLER_78_364 ();
 sg13g2_fill_1 FILLER_78_399 ();
 sg13g2_fill_2 FILLER_78_442 ();
 sg13g2_fill_2 FILLER_78_450 ();
 sg13g2_decap_4 FILLER_78_576 ();
 sg13g2_fill_2 FILLER_78_606 ();
 sg13g2_fill_1 FILLER_78_612 ();
 sg13g2_fill_2 FILLER_78_639 ();
 sg13g2_fill_2 FILLER_78_646 ();
 sg13g2_fill_1 FILLER_78_700 ();
 sg13g2_fill_2 FILLER_78_749 ();
 sg13g2_fill_1 FILLER_78_786 ();
 sg13g2_fill_1 FILLER_78_792 ();
 sg13g2_fill_1 FILLER_78_823 ();
 sg13g2_fill_1 FILLER_78_855 ();
 sg13g2_fill_2 FILLER_78_896 ();
 sg13g2_fill_1 FILLER_78_898 ();
 sg13g2_fill_1 FILLER_78_1012 ();
 sg13g2_fill_2 FILLER_78_1073 ();
 sg13g2_fill_2 FILLER_78_1084 ();
 sg13g2_fill_2 FILLER_78_1100 ();
 sg13g2_fill_1 FILLER_78_1180 ();
 sg13g2_fill_1 FILLER_78_1227 ();
 sg13g2_fill_1 FILLER_78_1233 ();
 sg13g2_fill_1 FILLER_78_1286 ();
 sg13g2_fill_1 FILLER_78_1313 ();
 sg13g2_fill_1 FILLER_78_1366 ();
 sg13g2_fill_1 FILLER_78_1389 ();
 sg13g2_fill_1 FILLER_78_1408 ();
 sg13g2_decap_4 FILLER_78_1439 ();
 sg13g2_fill_1 FILLER_78_1443 ();
 sg13g2_decap_4 FILLER_78_1517 ();
 sg13g2_fill_2 FILLER_78_1521 ();
 sg13g2_fill_1 FILLER_78_1527 ();
 sg13g2_fill_1 FILLER_78_1559 ();
 sg13g2_fill_2 FILLER_78_1595 ();
 sg13g2_fill_1 FILLER_78_1602 ();
 sg13g2_fill_1 FILLER_78_1629 ();
 sg13g2_fill_1 FILLER_78_1635 ();
 sg13g2_fill_1 FILLER_78_1662 ();
 sg13g2_fill_2 FILLER_78_1684 ();
 sg13g2_fill_1 FILLER_78_1790 ();
 sg13g2_fill_2 FILLER_78_1851 ();
 sg13g2_fill_1 FILLER_78_1884 ();
 sg13g2_fill_1 FILLER_78_1916 ();
 sg13g2_fill_2 FILLER_78_2023 ();
 sg13g2_fill_2 FILLER_78_2030 ();
 sg13g2_fill_1 FILLER_78_2088 ();
 sg13g2_fill_2 FILLER_78_2147 ();
 sg13g2_fill_1 FILLER_78_2157 ();
 sg13g2_fill_2 FILLER_78_2177 ();
 sg13g2_fill_1 FILLER_78_2199 ();
 sg13g2_fill_1 FILLER_78_2226 ();
 sg13g2_fill_1 FILLER_78_2247 ();
 sg13g2_fill_2 FILLER_78_2285 ();
 sg13g2_fill_1 FILLER_78_2292 ();
 sg13g2_fill_2 FILLER_78_2330 ();
 sg13g2_fill_1 FILLER_78_2411 ();
 sg13g2_fill_1 FILLER_78_2416 ();
 sg13g2_fill_1 FILLER_78_2422 ();
 sg13g2_fill_1 FILLER_78_2449 ();
 sg13g2_fill_2 FILLER_78_2480 ();
 sg13g2_fill_1 FILLER_78_2485 ();
 sg13g2_fill_2 FILLER_78_2489 ();
 sg13g2_fill_2 FILLER_78_2542 ();
 sg13g2_fill_1 FILLER_78_2544 ();
 sg13g2_decap_4 FILLER_78_2558 ();
 sg13g2_fill_1 FILLER_78_2588 ();
 sg13g2_decap_8 FILLER_78_2593 ();
 sg13g2_decap_8 FILLER_78_2600 ();
 sg13g2_decap_8 FILLER_78_2607 ();
 sg13g2_decap_8 FILLER_78_2614 ();
 sg13g2_decap_8 FILLER_78_2621 ();
 sg13g2_decap_8 FILLER_78_2628 ();
 sg13g2_decap_8 FILLER_78_2635 ();
 sg13g2_decap_8 FILLER_78_2642 ();
 sg13g2_decap_8 FILLER_78_2649 ();
 sg13g2_decap_8 FILLER_78_2656 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_101 ();
 sg13g2_fill_1 FILLER_79_172 ();
 sg13g2_fill_1 FILLER_79_199 ();
 sg13g2_fill_1 FILLER_79_231 ();
 sg13g2_fill_2 FILLER_79_311 ();
 sg13g2_fill_1 FILLER_79_330 ();
 sg13g2_fill_1 FILLER_79_376 ();
 sg13g2_fill_2 FILLER_79_429 ();
 sg13g2_fill_1 FILLER_79_465 ();
 sg13g2_fill_1 FILLER_79_491 ();
 sg13g2_fill_1 FILLER_79_576 ();
 sg13g2_fill_2 FILLER_79_590 ();
 sg13g2_fill_1 FILLER_79_592 ();
 sg13g2_fill_2 FILLER_79_597 ();
 sg13g2_fill_2 FILLER_79_603 ();
 sg13g2_fill_2 FILLER_79_609 ();
 sg13g2_fill_2 FILLER_79_616 ();
 sg13g2_fill_1 FILLER_79_618 ();
 sg13g2_fill_2 FILLER_79_623 ();
 sg13g2_fill_1 FILLER_79_625 ();
 sg13g2_decap_8 FILLER_79_630 ();
 sg13g2_decap_4 FILLER_79_667 ();
 sg13g2_fill_2 FILLER_79_731 ();
 sg13g2_decap_8 FILLER_79_737 ();
 sg13g2_fill_2 FILLER_79_744 ();
 sg13g2_fill_1 FILLER_79_776 ();
 sg13g2_fill_1 FILLER_79_781 ();
 sg13g2_fill_1 FILLER_79_808 ();
 sg13g2_fill_2 FILLER_79_852 ();
 sg13g2_decap_4 FILLER_79_888 ();
 sg13g2_fill_2 FILLER_79_892 ();
 sg13g2_decap_4 FILLER_79_898 ();
 sg13g2_fill_2 FILLER_79_902 ();
 sg13g2_fill_2 FILLER_79_929 ();
 sg13g2_fill_1 FILLER_79_931 ();
 sg13g2_fill_2 FILLER_79_936 ();
 sg13g2_fill_1 FILLER_79_964 ();
 sg13g2_fill_1 FILLER_79_969 ();
 sg13g2_fill_1 FILLER_79_974 ();
 sg13g2_fill_2 FILLER_79_1001 ();
 sg13g2_fill_2 FILLER_79_1012 ();
 sg13g2_fill_1 FILLER_79_1059 ();
 sg13g2_fill_2 FILLER_79_1067 ();
 sg13g2_fill_1 FILLER_79_1118 ();
 sg13g2_fill_2 FILLER_79_1144 ();
 sg13g2_fill_1 FILLER_79_1146 ();
 sg13g2_fill_1 FILLER_79_1190 ();
 sg13g2_fill_1 FILLER_79_1217 ();
 sg13g2_fill_1 FILLER_79_1221 ();
 sg13g2_fill_1 FILLER_79_1256 ();
 sg13g2_fill_2 FILLER_79_1267 ();
 sg13g2_fill_1 FILLER_79_1269 ();
 sg13g2_decap_8 FILLER_79_1330 ();
 sg13g2_decap_4 FILLER_79_1337 ();
 sg13g2_fill_2 FILLER_79_1341 ();
 sg13g2_fill_2 FILLER_79_1390 ();
 sg13g2_fill_1 FILLER_79_1397 ();
 sg13g2_decap_8 FILLER_79_1424 ();
 sg13g2_decap_8 FILLER_79_1431 ();
 sg13g2_fill_1 FILLER_79_1438 ();
 sg13g2_fill_1 FILLER_79_1504 ();
 sg13g2_fill_1 FILLER_79_1573 ();
 sg13g2_fill_1 FILLER_79_1630 ();
 sg13g2_decap_8 FILLER_79_1661 ();
 sg13g2_decap_8 FILLER_79_1668 ();
 sg13g2_decap_8 FILLER_79_1675 ();
 sg13g2_decap_4 FILLER_79_1682 ();
 sg13g2_fill_1 FILLER_79_1686 ();
 sg13g2_fill_1 FILLER_79_1705 ();
 sg13g2_fill_1 FILLER_79_1710 ();
 sg13g2_fill_2 FILLER_79_1728 ();
 sg13g2_decap_4 FILLER_79_1785 ();
 sg13g2_fill_1 FILLER_79_1789 ();
 sg13g2_decap_4 FILLER_79_1794 ();
 sg13g2_fill_1 FILLER_79_1824 ();
 sg13g2_fill_2 FILLER_79_1838 ();
 sg13g2_decap_8 FILLER_79_1871 ();
 sg13g2_fill_1 FILLER_79_1878 ();
 sg13g2_fill_2 FILLER_79_1909 ();
 sg13g2_fill_1 FILLER_79_1915 ();
 sg13g2_fill_1 FILLER_79_1920 ();
 sg13g2_decap_8 FILLER_79_1956 ();
 sg13g2_fill_1 FILLER_79_1963 ();
 sg13g2_fill_2 FILLER_79_1998 ();
 sg13g2_fill_1 FILLER_79_2048 ();
 sg13g2_fill_2 FILLER_79_2066 ();
 sg13g2_fill_2 FILLER_79_2072 ();
 sg13g2_fill_1 FILLER_79_2078 ();
 sg13g2_fill_2 FILLER_79_2083 ();
 sg13g2_fill_1 FILLER_79_2150 ();
 sg13g2_fill_2 FILLER_79_2155 ();
 sg13g2_fill_1 FILLER_79_2197 ();
 sg13g2_fill_1 FILLER_79_2214 ();
 sg13g2_fill_1 FILLER_79_2264 ();
 sg13g2_fill_1 FILLER_79_2274 ();
 sg13g2_fill_1 FILLER_79_2356 ();
 sg13g2_decap_4 FILLER_79_2386 ();
 sg13g2_fill_2 FILLER_79_2390 ();
 sg13g2_fill_1 FILLER_79_2397 ();
 sg13g2_fill_1 FILLER_79_2429 ();
 sg13g2_fill_1 FILLER_79_2456 ();
 sg13g2_decap_4 FILLER_79_2461 ();
 sg13g2_fill_2 FILLER_79_2465 ();
 sg13g2_fill_1 FILLER_79_2493 ();
 sg13g2_decap_8 FILLER_79_2533 ();
 sg13g2_fill_2 FILLER_79_2540 ();
 sg13g2_decap_8 FILLER_79_2568 ();
 sg13g2_decap_8 FILLER_79_2601 ();
 sg13g2_decap_8 FILLER_79_2608 ();
 sg13g2_decap_8 FILLER_79_2615 ();
 sg13g2_decap_8 FILLER_79_2622 ();
 sg13g2_decap_8 FILLER_79_2629 ();
 sg13g2_decap_8 FILLER_79_2636 ();
 sg13g2_decap_8 FILLER_79_2643 ();
 sg13g2_decap_8 FILLER_79_2650 ();
 sg13g2_decap_8 FILLER_79_2657 ();
 sg13g2_decap_4 FILLER_79_2664 ();
 sg13g2_fill_2 FILLER_79_2668 ();
 sg13g2_fill_1 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_96 ();
 sg13g2_fill_2 FILLER_80_192 ();
 sg13g2_fill_2 FILLER_80_303 ();
 sg13g2_fill_2 FILLER_80_404 ();
 sg13g2_fill_1 FILLER_80_468 ();
 sg13g2_fill_1 FILLER_80_517 ();
 sg13g2_fill_2 FILLER_80_552 ();
 sg13g2_fill_1 FILLER_80_561 ();
 sg13g2_decap_8 FILLER_80_580 ();
 sg13g2_fill_2 FILLER_80_587 ();
 sg13g2_fill_1 FILLER_80_589 ();
 sg13g2_decap_8 FILLER_80_629 ();
 sg13g2_decap_8 FILLER_80_636 ();
 sg13g2_fill_2 FILLER_80_643 ();
 sg13g2_decap_4 FILLER_80_649 ();
 sg13g2_fill_1 FILLER_80_653 ();
 sg13g2_decap_8 FILLER_80_658 ();
 sg13g2_decap_8 FILLER_80_665 ();
 sg13g2_decap_8 FILLER_80_672 ();
 sg13g2_decap_8 FILLER_80_687 ();
 sg13g2_decap_8 FILLER_80_694 ();
 sg13g2_fill_2 FILLER_80_701 ();
 sg13g2_fill_1 FILLER_80_703 ();
 sg13g2_fill_2 FILLER_80_717 ();
 sg13g2_decap_8 FILLER_80_723 ();
 sg13g2_decap_8 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_737 ();
 sg13g2_decap_4 FILLER_80_744 ();
 sg13g2_fill_2 FILLER_80_748 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_fill_2 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_792 ();
 sg13g2_fill_2 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_fill_1 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_852 ();
 sg13g2_decap_8 FILLER_80_859 ();
 sg13g2_decap_8 FILLER_80_866 ();
 sg13g2_fill_2 FILLER_80_873 ();
 sg13g2_fill_1 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_880 ();
 sg13g2_decap_8 FILLER_80_887 ();
 sg13g2_decap_8 FILLER_80_894 ();
 sg13g2_decap_8 FILLER_80_901 ();
 sg13g2_fill_2 FILLER_80_908 ();
 sg13g2_fill_1 FILLER_80_910 ();
 sg13g2_decap_8 FILLER_80_915 ();
 sg13g2_decap_8 FILLER_80_922 ();
 sg13g2_decap_4 FILLER_80_929 ();
 sg13g2_decap_4 FILLER_80_942 ();
 sg13g2_decap_8 FILLER_80_950 ();
 sg13g2_decap_8 FILLER_80_957 ();
 sg13g2_decap_8 FILLER_80_964 ();
 sg13g2_decap_8 FILLER_80_971 ();
 sg13g2_decap_4 FILLER_80_978 ();
 sg13g2_fill_1 FILLER_80_986 ();
 sg13g2_fill_2 FILLER_80_991 ();
 sg13g2_fill_2 FILLER_80_1042 ();
 sg13g2_decap_4 FILLER_80_1113 ();
 sg13g2_fill_1 FILLER_80_1117 ();
 sg13g2_decap_8 FILLER_80_1131 ();
 sg13g2_decap_8 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_decap_4 FILLER_80_1152 ();
 sg13g2_fill_2 FILLER_80_1173 ();
 sg13g2_fill_1 FILLER_80_1175 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_fill_1 FILLER_80_1194 ();
 sg13g2_fill_1 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1228 ();
 sg13g2_decap_4 FILLER_80_1256 ();
 sg13g2_fill_2 FILLER_80_1260 ();
 sg13g2_decap_8 FILLER_80_1274 ();
 sg13g2_decap_4 FILLER_80_1281 ();
 sg13g2_fill_2 FILLER_80_1285 ();
 sg13g2_fill_2 FILLER_80_1296 ();
 sg13g2_fill_1 FILLER_80_1302 ();
 sg13g2_decap_8 FILLER_80_1307 ();
 sg13g2_decap_8 FILLER_80_1314 ();
 sg13g2_decap_8 FILLER_80_1321 ();
 sg13g2_decap_8 FILLER_80_1328 ();
 sg13g2_decap_8 FILLER_80_1335 ();
 sg13g2_decap_4 FILLER_80_1342 ();
 sg13g2_fill_1 FILLER_80_1346 ();
 sg13g2_decap_4 FILLER_80_1355 ();
 sg13g2_fill_2 FILLER_80_1359 ();
 sg13g2_fill_2 FILLER_80_1379 ();
 sg13g2_fill_1 FILLER_80_1381 ();
 sg13g2_fill_1 FILLER_80_1386 ();
 sg13g2_decap_4 FILLER_80_1395 ();
 sg13g2_decap_8 FILLER_80_1429 ();
 sg13g2_decap_8 FILLER_80_1436 ();
 sg13g2_decap_4 FILLER_80_1443 ();
 sg13g2_fill_1 FILLER_80_1447 ();
 sg13g2_decap_8 FILLER_80_1452 ();
 sg13g2_decap_8 FILLER_80_1459 ();
 sg13g2_decap_4 FILLER_80_1466 ();
 sg13g2_decap_8 FILLER_80_1478 ();
 sg13g2_fill_2 FILLER_80_1485 ();
 sg13g2_decap_4 FILLER_80_1505 ();
 sg13g2_fill_1 FILLER_80_1509 ();
 sg13g2_decap_4 FILLER_80_1518 ();
 sg13g2_fill_2 FILLER_80_1522 ();
 sg13g2_decap_4 FILLER_80_1532 ();
 sg13g2_fill_2 FILLER_80_1536 ();
 sg13g2_decap_8 FILLER_80_1546 ();
 sg13g2_decap_8 FILLER_80_1553 ();
 sg13g2_decap_8 FILLER_80_1560 ();
 sg13g2_fill_2 FILLER_80_1567 ();
 sg13g2_fill_1 FILLER_80_1569 ();
 sg13g2_fill_1 FILLER_80_1587 ();
 sg13g2_decap_4 FILLER_80_1592 ();
 sg13g2_fill_2 FILLER_80_1596 ();
 sg13g2_decap_8 FILLER_80_1623 ();
 sg13g2_decap_4 FILLER_80_1634 ();
 sg13g2_fill_2 FILLER_80_1642 ();
 sg13g2_fill_1 FILLER_80_1644 ();
 sg13g2_decap_8 FILLER_80_1649 ();
 sg13g2_decap_8 FILLER_80_1656 ();
 sg13g2_decap_8 FILLER_80_1663 ();
 sg13g2_decap_8 FILLER_80_1670 ();
 sg13g2_decap_8 FILLER_80_1677 ();
 sg13g2_decap_8 FILLER_80_1684 ();
 sg13g2_decap_8 FILLER_80_1691 ();
 sg13g2_decap_8 FILLER_80_1698 ();
 sg13g2_fill_1 FILLER_80_1705 ();
 sg13g2_decap_8 FILLER_80_1710 ();
 sg13g2_decap_4 FILLER_80_1717 ();
 sg13g2_fill_1 FILLER_80_1721 ();
 sg13g2_fill_2 FILLER_80_1729 ();
 sg13g2_decap_8 FILLER_80_1782 ();
 sg13g2_decap_8 FILLER_80_1789 ();
 sg13g2_decap_8 FILLER_80_1796 ();
 sg13g2_decap_8 FILLER_80_1807 ();
 sg13g2_decap_8 FILLER_80_1814 ();
 sg13g2_decap_8 FILLER_80_1821 ();
 sg13g2_decap_8 FILLER_80_1828 ();
 sg13g2_decap_8 FILLER_80_1835 ();
 sg13g2_decap_4 FILLER_80_1842 ();
 sg13g2_fill_1 FILLER_80_1846 ();
 sg13g2_decap_4 FILLER_80_1855 ();
 sg13g2_decap_8 FILLER_80_1867 ();
 sg13g2_decap_8 FILLER_80_1874 ();
 sg13g2_decap_4 FILLER_80_1881 ();
 sg13g2_decap_8 FILLER_80_1889 ();
 sg13g2_fill_2 FILLER_80_1896 ();
 sg13g2_fill_1 FILLER_80_1898 ();
 sg13g2_decap_8 FILLER_80_1903 ();
 sg13g2_decap_8 FILLER_80_1910 ();
 sg13g2_decap_8 FILLER_80_1917 ();
 sg13g2_fill_2 FILLER_80_1924 ();
 sg13g2_fill_1 FILLER_80_1926 ();
 sg13g2_decap_8 FILLER_80_1931 ();
 sg13g2_decap_8 FILLER_80_1946 ();
 sg13g2_decap_8 FILLER_80_1953 ();
 sg13g2_decap_8 FILLER_80_1960 ();
 sg13g2_fill_2 FILLER_80_1967 ();
 sg13g2_fill_1 FILLER_80_1969 ();
 sg13g2_decap_8 FILLER_80_1978 ();
 sg13g2_fill_1 FILLER_80_1985 ();
 sg13g2_decap_8 FILLER_80_1990 ();
 sg13g2_decap_8 FILLER_80_1997 ();
 sg13g2_decap_8 FILLER_80_2004 ();
 sg13g2_fill_1 FILLER_80_2011 ();
 sg13g2_fill_2 FILLER_80_2020 ();
 sg13g2_fill_2 FILLER_80_2104 ();
 sg13g2_fill_2 FILLER_80_2148 ();
 sg13g2_fill_2 FILLER_80_2160 ();
 sg13g2_fill_2 FILLER_80_2189 ();
 sg13g2_fill_2 FILLER_80_2206 ();
 sg13g2_fill_2 FILLER_80_2216 ();
 sg13g2_fill_1 FILLER_80_2227 ();
 sg13g2_fill_2 FILLER_80_2270 ();
 sg13g2_fill_1 FILLER_80_2294 ();
 sg13g2_fill_2 FILLER_80_2299 ();
 sg13g2_fill_1 FILLER_80_2317 ();
 sg13g2_fill_1 FILLER_80_2323 ();
 sg13g2_fill_1 FILLER_80_2363 ();
 sg13g2_decap_8 FILLER_80_2396 ();
 sg13g2_decap_8 FILLER_80_2403 ();
 sg13g2_fill_1 FILLER_80_2410 ();
 sg13g2_decap_8 FILLER_80_2415 ();
 sg13g2_fill_1 FILLER_80_2422 ();
 sg13g2_fill_2 FILLER_80_2436 ();
 sg13g2_decap_8 FILLER_80_2442 ();
 sg13g2_decap_8 FILLER_80_2449 ();
 sg13g2_decap_8 FILLER_80_2456 ();
 sg13g2_fill_1 FILLER_80_2463 ();
 sg13g2_decap_4 FILLER_80_2506 ();
 sg13g2_decap_8 FILLER_80_2518 ();
 sg13g2_decap_8 FILLER_80_2525 ();
 sg13g2_decap_8 FILLER_80_2532 ();
 sg13g2_decap_8 FILLER_80_2539 ();
 sg13g2_decap_4 FILLER_80_2546 ();
 sg13g2_decap_8 FILLER_80_2554 ();
 sg13g2_decap_8 FILLER_80_2561 ();
 sg13g2_decap_8 FILLER_80_2568 ();
 sg13g2_decap_8 FILLER_80_2575 ();
 sg13g2_decap_8 FILLER_80_2586 ();
 sg13g2_decap_8 FILLER_80_2593 ();
 sg13g2_decap_8 FILLER_80_2600 ();
 sg13g2_decap_8 FILLER_80_2607 ();
 sg13g2_decap_8 FILLER_80_2614 ();
 sg13g2_decap_8 FILLER_80_2621 ();
 sg13g2_decap_8 FILLER_80_2628 ();
 sg13g2_decap_8 FILLER_80_2635 ();
 sg13g2_decap_8 FILLER_80_2642 ();
 sg13g2_decap_8 FILLER_80_2649 ();
 sg13g2_decap_8 FILLER_80_2656 ();
 sg13g2_decap_8 FILLER_80_2663 ();
endmodule
