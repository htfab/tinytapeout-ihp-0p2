module tt_um_hpretl_minilogix (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire _4601_;
 wire _4602_;
 wire _4603_;
 wire _4604_;
 wire _4605_;
 wire _4606_;
 wire _4607_;
 wire _4608_;
 wire _4609_;
 wire _4610_;
 wire _4611_;
 wire _4612_;
 wire _4613_;
 wire _4614_;
 wire _4615_;
 wire _4616_;
 wire _4617_;
 wire _4618_;
 wire _4619_;
 wire _4620_;
 wire _4621_;
 wire _4622_;
 wire _4623_;
 wire _4624_;
 wire _4625_;
 wire _4626_;
 wire _4627_;
 wire _4628_;
 wire _4629_;
 wire _4630_;
 wire _4631_;
 wire _4632_;
 wire _4633_;
 wire _4634_;
 wire _4635_;
 wire _4636_;
 wire _4637_;
 wire _4638_;
 wire _4639_;
 wire _4640_;
 wire _4641_;
 wire _4642_;
 wire _4643_;
 wire _4644_;
 wire _4645_;
 wire _4646_;
 wire _4647_;
 wire _4648_;
 wire _4649_;
 wire _4650_;
 wire _4651_;
 wire _4652_;
 wire _4653_;
 wire _4654_;
 wire _4655_;
 wire _4656_;
 wire _4657_;
 wire _4658_;
 wire _4659_;
 wire _4660_;
 wire _4661_;
 wire _4662_;
 wire _4663_;
 wire _4664_;
 wire _4665_;
 wire _4666_;
 wire _4667_;
 wire _4668_;
 wire _4669_;
 wire _4670_;
 wire _4671_;
 wire _4672_;
 wire _4673_;
 wire _4674_;
 wire _4675_;
 wire _4676_;
 wire _4677_;
 wire _4678_;
 wire _4679_;
 wire _4680_;
 wire _4681_;
 wire _4682_;
 wire _4683_;
 wire _4684_;
 wire _4685_;
 wire _4686_;
 wire _4687_;
 wire _4688_;
 wire _4689_;
 wire _4690_;
 wire _4691_;
 wire _4692_;
 wire _4693_;
 wire _4694_;
 wire _4695_;
 wire _4696_;
 wire _4697_;
 wire _4698_;
 wire _4699_;
 wire _4700_;
 wire _4701_;
 wire _4702_;
 wire _4703_;
 wire _4704_;
 wire _4705_;
 wire _4706_;
 wire _4707_;
 wire _4708_;
 wire _4709_;
 wire _4710_;
 wire _4711_;
 wire _4712_;
 wire _4713_;
 wire _4714_;
 wire _4715_;
 wire _4716_;
 wire _4717_;
 wire _4718_;
 wire _4719_;
 wire _4720_;
 wire _4721_;
 wire _4722_;
 wire _4723_;
 wire _4724_;
 wire _4725_;
 wire _4726_;
 wire _4727_;
 wire _4728_;
 wire _4729_;
 wire _4730_;
 wire _4731_;
 wire _4732_;
 wire _4733_;
 wire _4734_;
 wire _4735_;
 wire _4736_;
 wire _4737_;
 wire _4738_;
 wire _4739_;
 wire _4740_;
 wire _4741_;
 wire _4742_;
 wire _4743_;
 wire _4744_;
 wire _4745_;
 wire _4746_;
 wire _4747_;
 wire _4748_;
 wire _4749_;
 wire _4750_;
 wire _4751_;
 wire _4752_;
 wire _4753_;
 wire _4754_;
 wire _4755_;
 wire _4756_;
 wire _4757_;
 wire _4758_;
 wire _4759_;
 wire _4760_;
 wire _4761_;
 wire _4762_;
 wire _4763_;
 wire _4764_;
 wire _4765_;
 wire _4766_;
 wire _4767_;
 wire _4768_;
 wire _4769_;
 wire _4770_;
 wire _4771_;
 wire _4772_;
 wire _4773_;
 wire _4774_;
 wire _4775_;
 wire _4776_;
 wire _4777_;
 wire _4778_;
 wire _4779_;
 wire _4780_;
 wire _4781_;
 wire _4782_;
 wire _4783_;
 wire _4784_;
 wire _4785_;
 wire _4786_;
 wire _4787_;
 wire _4788_;
 wire _4789_;
 wire _4790_;
 wire _4791_;
 wire _4792_;
 wire _4793_;
 wire _4794_;
 wire _4795_;
 wire _4796_;
 wire _4797_;
 wire _4798_;
 wire _4799_;
 wire _4800_;
 wire _4801_;
 wire _4802_;
 wire _4803_;
 wire _4804_;
 wire _4805_;
 wire _4806_;
 wire _4807_;
 wire _4808_;
 wire _4809_;
 wire _4810_;
 wire _4811_;
 wire _4812_;
 wire _4813_;
 wire _4814_;
 wire _4815_;
 wire _4816_;
 wire _4817_;
 wire _4818_;
 wire _4819_;
 wire _4820_;
 wire _4821_;
 wire _4822_;
 wire _4823_;
 wire _4824_;
 wire _4825_;
 wire _4826_;
 wire _4827_;
 wire _4828_;
 wire _4829_;
 wire _4830_;
 wire _4831_;
 wire _4832_;
 wire _4833_;
 wire _4834_;
 wire _4835_;
 wire _4836_;
 wire _4837_;
 wire _4838_;
 wire _4839_;
 wire _4840_;
 wire _4841_;
 wire _4842_;
 wire _4843_;
 wire _4844_;
 wire _4845_;
 wire _4846_;
 wire _4847_;
 wire _4848_;
 wire _4849_;
 wire _4850_;
 wire _4851_;
 wire _4852_;
 wire _4853_;
 wire _4854_;
 wire _4855_;
 wire _4856_;
 wire _4857_;
 wire _4858_;
 wire _4859_;
 wire _4860_;
 wire _4861_;
 wire _4862_;
 wire _4863_;
 wire _4864_;
 wire _4865_;
 wire _4866_;
 wire _4867_;
 wire _4868_;
 wire _4869_;
 wire _4870_;
 wire _4871_;
 wire _4872_;
 wire _4873_;
 wire _4874_;
 wire _4875_;
 wire _4876_;
 wire _4877_;
 wire _4878_;
 wire _4879_;
 wire _4880_;
 wire _4881_;
 wire _4882_;
 wire _4883_;
 wire _4884_;
 wire _4885_;
 wire _4886_;
 wire _4887_;
 wire _4888_;
 wire _4889_;
 wire _4890_;
 wire _4891_;
 wire _4892_;
 wire _4893_;
 wire _4894_;
 wire _4895_;
 wire _4896_;
 wire _4897_;
 wire _4898_;
 wire _4899_;
 wire _4900_;
 wire _4901_;
 wire _4902_;
 wire _4903_;
 wire _4904_;
 wire _4905_;
 wire _4906_;
 wire _4907_;
 wire _4908_;
 wire _4909_;
 wire _4910_;
 wire _4911_;
 wire _4912_;
 wire _4913_;
 wire _4914_;
 wire _4915_;
 wire _4916_;
 wire _4917_;
 wire _4918_;
 wire _4919_;
 wire _4920_;
 wire _4921_;
 wire _4922_;
 wire _4923_;
 wire _4924_;
 wire _4925_;
 wire _4926_;
 wire _4927_;
 wire _4928_;
 wire _4929_;
 wire _4930_;
 wire _4931_;
 wire _4932_;
 wire _4933_;
 wire _4934_;
 wire _4935_;
 wire _4936_;
 wire _4937_;
 wire _4938_;
 wire _4939_;
 wire _4940_;
 wire _4941_;
 wire _4942_;
 wire _4943_;
 wire _4944_;
 wire _4945_;
 wire _4946_;
 wire _4947_;
 wire _4948_;
 wire _4949_;
 wire _4950_;
 wire _4951_;
 wire _4952_;
 wire _4953_;
 wire _4954_;
 wire _4955_;
 wire _4956_;
 wire _4957_;
 wire _4958_;
 wire _4959_;
 wire _4960_;
 wire _4961_;
 wire _4962_;
 wire _4963_;
 wire _4964_;
 wire _4965_;
 wire _4966_;
 wire _4967_;
 wire _4968_;
 wire _4969_;
 wire _4970_;
 wire _4971_;
 wire _4972_;
 wire _4973_;
 wire _4974_;
 wire _4975_;
 wire _4976_;
 wire _4977_;
 wire _4978_;
 wire _4979_;
 wire _4980_;
 wire _4981_;
 wire _4982_;
 wire _4983_;
 wire _4984_;
 wire _4985_;
 wire _4986_;
 wire _4987_;
 wire _4988_;
 wire _4989_;
 wire _4990_;
 wire _4991_;
 wire _4992_;
 wire _4993_;
 wire _4994_;
 wire _4995_;
 wire _4996_;
 wire _4997_;
 wire _4998_;
 wire _4999_;
 wire _5000_;
 wire _5001_;
 wire _5002_;
 wire _5003_;
 wire _5004_;
 wire _5005_;
 wire _5006_;
 wire _5007_;
 wire _5008_;
 wire _5009_;
 wire _5010_;
 wire _5011_;
 wire _5012_;
 wire _5013_;
 wire _5014_;
 wire _5015_;
 wire _5016_;
 wire _5017_;
 wire _5018_;
 wire _5019_;
 wire _5020_;
 wire _5021_;
 wire _5022_;
 wire _5023_;
 wire _5024_;
 wire _5025_;
 wire _5026_;
 wire _5027_;
 wire _5028_;
 wire _5029_;
 wire _5030_;
 wire _5031_;
 wire _5032_;
 wire _5033_;
 wire _5034_;
 wire _5035_;
 wire _5036_;
 wire _5037_;
 wire _5038_;
 wire _5039_;
 wire _5040_;
 wire _5041_;
 wire _5042_;
 wire _5043_;
 wire _5044_;
 wire _5045_;
 wire _5046_;
 wire _5047_;
 wire _5048_;
 wire _5049_;
 wire _5050_;
 wire _5051_;
 wire _5052_;
 wire _5053_;
 wire _5054_;
 wire _5055_;
 wire _5056_;
 wire _5057_;
 wire _5058_;
 wire _5059_;
 wire _5060_;
 wire _5061_;
 wire _5062_;
 wire _5063_;
 wire _5064_;
 wire _5065_;
 wire _5066_;
 wire _5067_;
 wire _5068_;
 wire _5069_;
 wire _5070_;
 wire _5071_;
 wire _5072_;
 wire _5073_;
 wire _5074_;
 wire _5075_;
 wire _5076_;
 wire _5077_;
 wire _5078_;
 wire _5079_;
 wire _5080_;
 wire _5081_;
 wire _5082_;
 wire _5083_;
 wire _5084_;
 wire _5085_;
 wire _5086_;
 wire _5087_;
 wire _5088_;
 wire _5089_;
 wire _5090_;
 wire _5091_;
 wire _5092_;
 wire _5093_;
 wire _5094_;
 wire _5095_;
 wire _5096_;
 wire _5097_;
 wire _5098_;
 wire _5099_;
 wire _5100_;
 wire _5101_;
 wire _5102_;
 wire _5103_;
 wire _5104_;
 wire _5105_;
 wire _5106_;
 wire _5107_;
 wire _5108_;
 wire _5109_;
 wire _5110_;
 wire _5111_;
 wire _5112_;
 wire _5113_;
 wire _5114_;
 wire _5115_;
 wire _5116_;
 wire _5117_;
 wire _5118_;
 wire _5119_;
 wire _5120_;
 wire _5121_;
 wire _5122_;
 wire _5123_;
 wire _5124_;
 wire _5125_;
 wire _5126_;
 wire _5127_;
 wire _5128_;
 wire _5129_;
 wire _5130_;
 wire _5131_;
 wire _5132_;
 wire _5133_;
 wire _5134_;
 wire _5135_;
 wire _5136_;
 wire _5137_;
 wire _5138_;
 wire _5139_;
 wire _5140_;
 wire _5141_;
 wire _5142_;
 wire _5143_;
 wire _5144_;
 wire _5145_;
 wire _5146_;
 wire _5147_;
 wire _5148_;
 wire _5149_;
 wire _5150_;
 wire _5151_;
 wire _5152_;
 wire _5153_;
 wire _5154_;
 wire _5155_;
 wire _5156_;
 wire _5157_;
 wire _5158_;
 wire _5159_;
 wire _5160_;
 wire _5161_;
 wire _5162_;
 wire _5163_;
 wire _5164_;
 wire _5165_;
 wire _5166_;
 wire _5167_;
 wire _5168_;
 wire _5169_;
 wire _5170_;
 wire _5171_;
 wire _5172_;
 wire _5173_;
 wire _5174_;
 wire _5175_;
 wire _5176_;
 wire _5177_;
 wire _5178_;
 wire _5179_;
 wire _5180_;
 wire _5181_;
 wire _5182_;
 wire _5183_;
 wire _5184_;
 wire _5185_;
 wire _5186_;
 wire _5187_;
 wire _5188_;
 wire _5189_;
 wire _5190_;
 wire _5191_;
 wire _5192_;
 wire _5193_;
 wire _5194_;
 wire _5195_;
 wire _5196_;
 wire _5197_;
 wire _5198_;
 wire _5199_;
 wire _5200_;
 wire _5201_;
 wire _5202_;
 wire _5203_;
 wire _5204_;
 wire _5205_;
 wire _5206_;
 wire _5207_;
 wire _5208_;
 wire _5209_;
 wire _5210_;
 wire _5211_;
 wire _5212_;
 wire _5213_;
 wire _5214_;
 wire _5215_;
 wire _5216_;
 wire _5217_;
 wire _5218_;
 wire _5219_;
 wire _5220_;
 wire _5221_;
 wire _5222_;
 wire _5223_;
 wire _5224_;
 wire _5225_;
 wire _5226_;
 wire _5227_;
 wire _5228_;
 wire _5229_;
 wire _5230_;
 wire _5231_;
 wire _5232_;
 wire _5233_;
 wire _5234_;
 wire _5235_;
 wire _5236_;
 wire _5237_;
 wire _5238_;
 wire _5239_;
 wire _5240_;
 wire _5241_;
 wire _5242_;
 wire _5243_;
 wire _5244_;
 wire _5245_;
 wire _5246_;
 wire _5247_;
 wire _5248_;
 wire _5249_;
 wire _5250_;
 wire _5251_;
 wire _5252_;
 wire _5253_;
 wire _5254_;
 wire _5255_;
 wire _5256_;
 wire _5257_;
 wire _5258_;
 wire _5259_;
 wire _5260_;
 wire _5261_;
 wire _5262_;
 wire _5263_;
 wire _5264_;
 wire _5265_;
 wire _5266_;
 wire _5267_;
 wire _5268_;
 wire _5269_;
 wire _5270_;
 wire _5271_;
 wire _5272_;
 wire _5273_;
 wire _5274_;
 wire _5275_;
 wire _5276_;
 wire _5277_;
 wire _5278_;
 wire _5279_;
 wire _5280_;
 wire _5281_;
 wire _5282_;
 wire _5283_;
 wire _5284_;
 wire _5285_;
 wire _5286_;
 wire _5287_;
 wire _5288_;
 wire _5289_;
 wire _5290_;
 wire _5291_;
 wire _5292_;
 wire _5293_;
 wire _5294_;
 wire _5295_;
 wire _5296_;
 wire _5297_;
 wire _5298_;
 wire _5299_;
 wire _5300_;
 wire _5301_;
 wire _5302_;
 wire _5303_;
 wire _5304_;
 wire _5305_;
 wire _5306_;
 wire _5307_;
 wire _5308_;
 wire _5309_;
 wire _5310_;
 wire _5311_;
 wire _5312_;
 wire _5313_;
 wire _5314_;
 wire _5315_;
 wire _5316_;
 wire _5317_;
 wire _5318_;
 wire _5319_;
 wire _5320_;
 wire _5321_;
 wire _5322_;
 wire _5323_;
 wire _5324_;
 wire _5325_;
 wire _5326_;
 wire _5327_;
 wire _5328_;
 wire _5329_;
 wire _5330_;
 wire _5331_;
 wire _5332_;
 wire _5333_;
 wire _5334_;
 wire _5335_;
 wire _5336_;
 wire _5337_;
 wire _5338_;
 wire _5339_;
 wire _5340_;
 wire _5341_;
 wire _5342_;
 wire _5343_;
 wire _5344_;
 wire _5345_;
 wire _5346_;
 wire _5347_;
 wire _5348_;
 wire _5349_;
 wire _5350_;
 wire _5351_;
 wire _5352_;
 wire _5353_;
 wire _5354_;
 wire _5355_;
 wire _5356_;
 wire _5357_;
 wire _5358_;
 wire _5359_;
 wire _5360_;
 wire _5361_;
 wire _5362_;
 wire _5363_;
 wire _5364_;
 wire _5365_;
 wire _5366_;
 wire _5367_;
 wire _5368_;
 wire _5369_;
 wire _5370_;
 wire _5371_;
 wire _5372_;
 wire _5373_;
 wire _5374_;
 wire _5375_;
 wire _5376_;
 wire _5377_;
 wire _5378_;
 wire _5379_;
 wire _5380_;
 wire _5381_;
 wire _5382_;
 wire _5383_;
 wire _5384_;
 wire _5385_;
 wire _5386_;
 wire _5387_;
 wire _5388_;
 wire _5389_;
 wire _5390_;
 wire _5391_;
 wire _5392_;
 wire _5393_;
 wire _5394_;
 wire _5395_;
 wire _5396_;
 wire _5397_;
 wire _5398_;
 wire _5399_;
 wire _5400_;
 wire _5401_;
 wire _5402_;
 wire _5403_;
 wire _5404_;
 wire _5405_;
 wire _5406_;
 wire _5407_;
 wire _5408_;
 wire _5409_;
 wire _5410_;
 wire _5411_;
 wire _5412_;
 wire _5413_;
 wire _5414_;
 wire _5415_;
 wire _5416_;
 wire _5417_;
 wire _5418_;
 wire _5419_;
 wire _5420_;
 wire _5421_;
 wire _5422_;
 wire _5423_;
 wire _5424_;
 wire _5425_;
 wire _5426_;
 wire _5427_;
 wire _5428_;
 wire _5429_;
 wire _5430_;
 wire _5431_;
 wire _5432_;
 wire _5433_;
 wire _5434_;
 wire _5435_;
 wire _5436_;
 wire _5437_;
 wire _5438_;
 wire _5439_;
 wire _5440_;
 wire _5441_;
 wire _5442_;
 wire _5443_;
 wire _5444_;
 wire _5445_;
 wire _5446_;
 wire _5447_;
 wire _5448_;
 wire _5449_;
 wire _5450_;
 wire _5451_;
 wire _5452_;
 wire _5453_;
 wire _5454_;
 wire _5455_;
 wire _5456_;
 wire _5457_;
 wire _5458_;
 wire _5459_;
 wire _5460_;
 wire _5461_;
 wire _5462_;
 wire _5463_;
 wire _5464_;
 wire _5465_;
 wire _5466_;
 wire _5467_;
 wire _5468_;
 wire _5469_;
 wire _5470_;
 wire _5471_;
 wire _5472_;
 wire _5473_;
 wire _5474_;
 wire _5475_;
 wire _5476_;
 wire _5477_;
 wire _5478_;
 wire _5479_;
 wire _5480_;
 wire _5481_;
 wire _5482_;
 wire _5483_;
 wire _5484_;
 wire _5485_;
 wire _5486_;
 wire _5487_;
 wire _5488_;
 wire _5489_;
 wire _5490_;
 wire _5491_;
 wire _5492_;
 wire _5493_;
 wire _5494_;
 wire _5495_;
 wire _5496_;
 wire _5497_;
 wire _5498_;
 wire _5499_;
 wire _5500_;
 wire _5501_;
 wire _5502_;
 wire _5503_;
 wire _5504_;
 wire _5505_;
 wire _5506_;
 wire _5507_;
 wire _5508_;
 wire _5509_;
 wire _5510_;
 wire _5511_;
 wire _5512_;
 wire _5513_;
 wire _5514_;
 wire _5515_;
 wire _5516_;
 wire _5517_;
 wire _5518_;
 wire _5519_;
 wire _5520_;
 wire _5521_;
 wire _5522_;
 wire _5523_;
 wire _5524_;
 wire _5525_;
 wire _5526_;
 wire _5527_;
 wire _5528_;
 wire _5529_;
 wire _5530_;
 wire _5531_;
 wire _5532_;
 wire _5533_;
 wire _5534_;
 wire _5535_;
 wire _5536_;
 wire _5537_;
 wire _5538_;
 wire _5539_;
 wire _5540_;
 wire _5541_;
 wire _5542_;
 wire _5543_;
 wire _5544_;
 wire _5545_;
 wire _5546_;
 wire _5547_;
 wire _5548_;
 wire _5549_;
 wire _5550_;
 wire _5551_;
 wire _5552_;
 wire _5553_;
 wire _5554_;
 wire _5555_;
 wire _5556_;
 wire _5557_;
 wire _5558_;
 wire _5559_;
 wire _5560_;
 wire _5561_;
 wire _5562_;
 wire _5563_;
 wire _5564_;
 wire _5565_;
 wire _5566_;
 wire _5567_;
 wire _5568_;
 wire _5569_;
 wire _5570_;
 wire _5571_;
 wire _5572_;
 wire _5573_;
 wire _5574_;
 wire _5575_;
 wire _5576_;
 wire _5577_;
 wire _5578_;
 wire _5579_;
 wire _5580_;
 wire _5581_;
 wire _5582_;
 wire _5583_;
 wire _5584_;
 wire _5585_;
 wire _5586_;
 wire _5587_;
 wire _5588_;
 wire _5589_;
 wire _5590_;
 wire _5591_;
 wire _5592_;
 wire _5593_;
 wire _5594_;
 wire _5595_;
 wire _5596_;
 wire _5597_;
 wire _5598_;
 wire _5599_;
 wire _5600_;
 wire _5601_;
 wire _5602_;
 wire _5603_;
 wire _5604_;
 wire _5605_;
 wire _5606_;
 wire _5607_;
 wire _5608_;
 wire _5609_;
 wire _5610_;
 wire _5611_;
 wire _5612_;
 wire _5613_;
 wire _5614_;
 wire _5615_;
 wire _5616_;
 wire _5617_;
 wire _5618_;
 wire _5619_;
 wire _5620_;
 wire _5621_;
 wire _5622_;
 wire _5623_;
 wire _5624_;
 wire _5625_;
 wire _5626_;
 wire _5627_;
 wire _5628_;
 wire _5629_;
 wire _5630_;
 wire _5631_;
 wire _5632_;
 wire _5633_;
 wire _5634_;
 wire _5635_;
 wire _5636_;
 wire _5637_;
 wire _5638_;
 wire _5639_;
 wire _5640_;
 wire _5641_;
 wire _5642_;
 wire _5643_;
 wire _5644_;
 wire _5645_;
 wire _5646_;
 wire _5647_;
 wire _5648_;
 wire _5649_;
 wire _5650_;
 wire _5651_;
 wire _5652_;
 wire _5653_;
 wire _5654_;
 wire _5655_;
 wire _5656_;
 wire _5657_;
 wire _5658_;
 wire _5659_;
 wire _5660_;
 wire _5661_;
 wire _5662_;
 wire _5663_;
 wire _5664_;
 wire _5665_;
 wire _5666_;
 wire _5667_;
 wire _5668_;
 wire _5669_;
 wire _5670_;
 wire _5671_;
 wire _5672_;
 wire _5673_;
 wire _5674_;
 wire _5675_;
 wire _5676_;
 wire _5677_;
 wire _5678_;
 wire _5679_;
 wire _5680_;
 wire _5681_;
 wire _5682_;
 wire _5683_;
 wire _5684_;
 wire _5685_;
 wire _5686_;
 wire _5687_;
 wire _5688_;
 wire _5689_;
 wire _5690_;
 wire _5691_;
 wire _5692_;
 wire _5693_;
 wire _5694_;
 wire _5695_;
 wire _5696_;
 wire _5697_;
 wire _5698_;
 wire _5699_;
 wire _5700_;
 wire _5701_;
 wire _5702_;
 wire _5703_;
 wire _5704_;
 wire _5705_;
 wire _5706_;
 wire _5707_;
 wire _5708_;
 wire _5709_;
 wire _5710_;
 wire _5711_;
 wire _5712_;
 wire _5713_;
 wire _5714_;
 wire _5715_;
 wire _5716_;
 wire _5717_;
 wire _5718_;
 wire _5719_;
 wire _5720_;
 wire _5721_;
 wire _5722_;
 wire _5723_;
 wire _5724_;
 wire _5725_;
 wire _5726_;
 wire _5727_;
 wire _5728_;
 wire _5729_;
 wire _5730_;
 wire _5731_;
 wire _5732_;
 wire _5733_;
 wire _5734_;
 wire _5735_;
 wire _5736_;
 wire _5737_;
 wire _5738_;
 wire _5739_;
 wire _5740_;
 wire _5741_;
 wire _5742_;
 wire _5743_;
 wire _5744_;
 wire _5745_;
 wire _5746_;
 wire _5747_;
 wire _5748_;
 wire _5749_;
 wire _5750_;
 wire _5751_;
 wire _5752_;
 wire _5753_;
 wire _5754_;
 wire _5755_;
 wire _5756_;
 wire _5757_;
 wire _5758_;
 wire _5759_;
 wire _5760_;
 wire _5761_;
 wire _5762_;
 wire _5763_;
 wire _5764_;
 wire _5765_;
 wire _5766_;
 wire _5767_;
 wire _5768_;
 wire _5769_;
 wire _5770_;
 wire _5771_;
 wire _5772_;
 wire _5773_;
 wire _5774_;
 wire _5775_;
 wire _5776_;
 wire _5777_;
 wire _5778_;
 wire _5779_;
 wire _5780_;
 wire _5781_;
 wire _5782_;
 wire _5783_;
 wire _5784_;
 wire _5785_;
 wire _5786_;
 wire _5787_;
 wire _5788_;
 wire _5789_;
 wire _5790_;
 wire _5791_;
 wire _5792_;
 wire _5793_;
 wire _5794_;
 wire _5795_;
 wire _5796_;
 wire _5797_;
 wire _5798_;
 wire _5799_;
 wire _5800_;
 wire _5801_;
 wire _5802_;
 wire _5803_;
 wire _5804_;
 wire _5805_;
 wire _5806_;
 wire _5807_;
 wire _5808_;
 wire _5809_;
 wire _5810_;
 wire _5811_;
 wire _5812_;
 wire _5813_;
 wire _5814_;
 wire _5815_;
 wire _5816_;
 wire _5817_;
 wire _5818_;
 wire _5819_;
 wire _5820_;
 wire _5821_;
 wire _5822_;
 wire _5823_;
 wire _5824_;
 wire _5825_;
 wire _5826_;
 wire _5827_;
 wire _5828_;
 wire _5829_;
 wire _5830_;
 wire _5831_;
 wire _5832_;
 wire _5833_;
 wire _5834_;
 wire _5835_;
 wire _5836_;
 wire _5837_;
 wire _5838_;
 wire _5839_;
 wire _5840_;
 wire _5841_;
 wire _5842_;
 wire _5843_;
 wire _5844_;
 wire _5845_;
 wire _5846_;
 wire _5847_;
 wire _5848_;
 wire _5849_;
 wire _5850_;
 wire _5851_;
 wire _5852_;
 wire _5853_;
 wire _5854_;
 wire _5855_;
 wire _5856_;
 wire _5857_;
 wire _5858_;
 wire _5859_;
 wire _5860_;
 wire _5861_;
 wire _5862_;
 wire _5863_;
 wire _5864_;
 wire _5865_;
 wire _5866_;
 wire _5867_;
 wire _5868_;
 wire _5869_;
 wire _5870_;
 wire _5871_;
 wire _5872_;
 wire _5873_;
 wire _5874_;
 wire _5875_;
 wire _5876_;
 wire _5877_;
 wire _5878_;
 wire _5879_;
 wire _5880_;
 wire _5881_;
 wire _5882_;
 wire _5883_;
 wire _5884_;
 wire _5885_;
 wire _5886_;
 wire _5887_;
 wire _5888_;
 wire _5889_;
 wire _5890_;
 wire _5891_;
 wire _5892_;
 wire _5893_;
 wire _5894_;
 wire _5895_;
 wire _5896_;
 wire _5897_;
 wire _5898_;
 wire _5899_;
 wire _5900_;
 wire _5901_;
 wire _5902_;
 wire _5903_;
 wire _5904_;
 wire _5905_;
 wire _5906_;
 wire _5907_;
 wire _5908_;
 wire _5909_;
 wire _5910_;
 wire _5911_;
 wire _5912_;
 wire _5913_;
 wire _5914_;
 wire _5915_;
 wire _5916_;
 wire _5917_;
 wire _5918_;
 wire _5919_;
 wire _5920_;
 wire _5921_;
 wire _5922_;
 wire _5923_;
 wire _5924_;
 wire _5925_;
 wire _5926_;
 wire _5927_;
 wire _5928_;
 wire _5929_;
 wire _5930_;
 wire _5931_;
 wire _5932_;
 wire _5933_;
 wire _5934_;
 wire _5935_;
 wire _5936_;
 wire _5937_;
 wire _5938_;
 wire _5939_;
 wire _5940_;
 wire _5941_;
 wire _5942_;
 wire _5943_;
 wire _5944_;
 wire _5945_;
 wire _5946_;
 wire _5947_;
 wire _5948_;
 wire _5949_;
 wire _5950_;
 wire _5951_;
 wire _5952_;
 wire _5953_;
 wire _5954_;
 wire _5955_;
 wire _5956_;
 wire _5957_;
 wire _5958_;
 wire _5959_;
 wire _5960_;
 wire _5961_;
 wire _5962_;
 wire _5963_;
 wire _5964_;
 wire _5965_;
 wire _5966_;
 wire _5967_;
 wire _5968_;
 wire _5969_;
 wire _5970_;
 wire _5971_;
 wire _5972_;
 wire _5973_;
 wire _5974_;
 wire _5975_;
 wire _5976_;
 wire _5977_;
 wire _5978_;
 wire _5979_;
 wire _5980_;
 wire _5981_;
 wire _5982_;
 wire _5983_;
 wire _5984_;
 wire _5985_;
 wire _5986_;
 wire _5987_;
 wire _5988_;
 wire _5989_;
 wire _5990_;
 wire _5991_;
 wire _5992_;
 wire clknet_0_clk;
 wire net787;
 wire \logix.feedback_r[0] ;
 wire \logix.feedback_r[1] ;
 wire \logix.feedback_r[2] ;
 wire \logix.feedback_r[3] ;
 wire \logix.feedback_r[4] ;
 wire \logix.feedback_r[5] ;
 wire \logix.feedback_r[6] ;
 wire \logix.feedback_r[7] ;
 wire \logix.input_sel_cfg_w[0] ;
 wire \logix.input_sel_cfg_w[1] ;
 wire \logix.input_sel_cfg_w[2] ;
 wire \logix.input_sel_cfg_w[3] ;
 wire \logix.input_sel_cfg_w[4] ;
 wire \logix.input_sel_cfg_w[5] ;
 wire \logix.input_sel_cfg_w[6] ;
 wire \logix.input_sel_cfg_w[7] ;
 wire \logix.ram_r[0] ;
 wire \logix.ram_r[1000] ;
 wire \logix.ram_r[1001] ;
 wire \logix.ram_r[1002] ;
 wire \logix.ram_r[1003] ;
 wire \logix.ram_r[1004] ;
 wire \logix.ram_r[1005] ;
 wire \logix.ram_r[1006] ;
 wire \logix.ram_r[1007] ;
 wire \logix.ram_r[1008] ;
 wire \logix.ram_r[1009] ;
 wire \logix.ram_r[100] ;
 wire \logix.ram_r[1010] ;
 wire \logix.ram_r[1011] ;
 wire \logix.ram_r[1012] ;
 wire \logix.ram_r[1013] ;
 wire \logix.ram_r[1014] ;
 wire \logix.ram_r[1015] ;
 wire \logix.ram_r[1016] ;
 wire \logix.ram_r[1017] ;
 wire \logix.ram_r[1018] ;
 wire \logix.ram_r[1019] ;
 wire \logix.ram_r[101] ;
 wire \logix.ram_r[1020] ;
 wire \logix.ram_r[1021] ;
 wire \logix.ram_r[1022] ;
 wire \logix.ram_r[1023] ;
 wire \logix.ram_r[1024] ;
 wire \logix.ram_r[1025] ;
 wire \logix.ram_r[1026] ;
 wire \logix.ram_r[1027] ;
 wire \logix.ram_r[1028] ;
 wire \logix.ram_r[1029] ;
 wire \logix.ram_r[102] ;
 wire \logix.ram_r[1030] ;
 wire \logix.ram_r[1031] ;
 wire \logix.ram_r[1032] ;
 wire \logix.ram_r[1033] ;
 wire \logix.ram_r[1034] ;
 wire \logix.ram_r[1035] ;
 wire \logix.ram_r[1036] ;
 wire \logix.ram_r[1037] ;
 wire \logix.ram_r[1038] ;
 wire \logix.ram_r[1039] ;
 wire \logix.ram_r[103] ;
 wire \logix.ram_r[1040] ;
 wire \logix.ram_r[1041] ;
 wire \logix.ram_r[1042] ;
 wire \logix.ram_r[1043] ;
 wire \logix.ram_r[1044] ;
 wire \logix.ram_r[1045] ;
 wire \logix.ram_r[1046] ;
 wire \logix.ram_r[1047] ;
 wire \logix.ram_r[1048] ;
 wire \logix.ram_r[1049] ;
 wire \logix.ram_r[104] ;
 wire \logix.ram_r[1050] ;
 wire \logix.ram_r[1051] ;
 wire \logix.ram_r[1052] ;
 wire \logix.ram_r[1053] ;
 wire \logix.ram_r[1054] ;
 wire \logix.ram_r[1055] ;
 wire \logix.ram_r[1056] ;
 wire \logix.ram_r[1057] ;
 wire \logix.ram_r[1058] ;
 wire \logix.ram_r[1059] ;
 wire \logix.ram_r[105] ;
 wire \logix.ram_r[1060] ;
 wire \logix.ram_r[1061] ;
 wire \logix.ram_r[1062] ;
 wire \logix.ram_r[1063] ;
 wire \logix.ram_r[1064] ;
 wire \logix.ram_r[1065] ;
 wire \logix.ram_r[1066] ;
 wire \logix.ram_r[1067] ;
 wire \logix.ram_r[1068] ;
 wire \logix.ram_r[1069] ;
 wire \logix.ram_r[106] ;
 wire \logix.ram_r[1070] ;
 wire \logix.ram_r[1071] ;
 wire \logix.ram_r[1072] ;
 wire \logix.ram_r[1073] ;
 wire \logix.ram_r[1074] ;
 wire \logix.ram_r[1075] ;
 wire \logix.ram_r[1076] ;
 wire \logix.ram_r[1077] ;
 wire \logix.ram_r[1078] ;
 wire \logix.ram_r[1079] ;
 wire \logix.ram_r[107] ;
 wire \logix.ram_r[1080] ;
 wire \logix.ram_r[1081] ;
 wire \logix.ram_r[1082] ;
 wire \logix.ram_r[1083] ;
 wire \logix.ram_r[1084] ;
 wire \logix.ram_r[1085] ;
 wire \logix.ram_r[1086] ;
 wire \logix.ram_r[1087] ;
 wire \logix.ram_r[1088] ;
 wire \logix.ram_r[1089] ;
 wire \logix.ram_r[108] ;
 wire \logix.ram_r[1090] ;
 wire \logix.ram_r[1091] ;
 wire \logix.ram_r[1092] ;
 wire \logix.ram_r[1093] ;
 wire \logix.ram_r[1094] ;
 wire \logix.ram_r[1095] ;
 wire \logix.ram_r[1096] ;
 wire \logix.ram_r[1097] ;
 wire \logix.ram_r[1098] ;
 wire \logix.ram_r[1099] ;
 wire \logix.ram_r[109] ;
 wire \logix.ram_r[10] ;
 wire \logix.ram_r[1100] ;
 wire \logix.ram_r[1101] ;
 wire \logix.ram_r[1102] ;
 wire \logix.ram_r[1103] ;
 wire \logix.ram_r[1104] ;
 wire \logix.ram_r[1105] ;
 wire \logix.ram_r[1106] ;
 wire \logix.ram_r[1107] ;
 wire \logix.ram_r[1108] ;
 wire \logix.ram_r[1109] ;
 wire \logix.ram_r[110] ;
 wire \logix.ram_r[1110] ;
 wire \logix.ram_r[1111] ;
 wire \logix.ram_r[1112] ;
 wire \logix.ram_r[1113] ;
 wire \logix.ram_r[1114] ;
 wire \logix.ram_r[1115] ;
 wire \logix.ram_r[1116] ;
 wire \logix.ram_r[1117] ;
 wire \logix.ram_r[1118] ;
 wire \logix.ram_r[1119] ;
 wire \logix.ram_r[111] ;
 wire \logix.ram_r[1120] ;
 wire \logix.ram_r[1121] ;
 wire \logix.ram_r[1122] ;
 wire \logix.ram_r[1123] ;
 wire \logix.ram_r[1124] ;
 wire \logix.ram_r[1125] ;
 wire \logix.ram_r[1126] ;
 wire \logix.ram_r[1127] ;
 wire \logix.ram_r[1128] ;
 wire \logix.ram_r[1129] ;
 wire \logix.ram_r[112] ;
 wire \logix.ram_r[1130] ;
 wire \logix.ram_r[1131] ;
 wire \logix.ram_r[1132] ;
 wire \logix.ram_r[1133] ;
 wire \logix.ram_r[1134] ;
 wire \logix.ram_r[1135] ;
 wire \logix.ram_r[1136] ;
 wire \logix.ram_r[1137] ;
 wire \logix.ram_r[1138] ;
 wire \logix.ram_r[1139] ;
 wire \logix.ram_r[113] ;
 wire \logix.ram_r[1140] ;
 wire \logix.ram_r[1141] ;
 wire \logix.ram_r[1142] ;
 wire \logix.ram_r[1143] ;
 wire \logix.ram_r[1144] ;
 wire \logix.ram_r[1145] ;
 wire \logix.ram_r[1146] ;
 wire \logix.ram_r[1147] ;
 wire \logix.ram_r[1148] ;
 wire \logix.ram_r[1149] ;
 wire \logix.ram_r[114] ;
 wire \logix.ram_r[1150] ;
 wire \logix.ram_r[1151] ;
 wire \logix.ram_r[1152] ;
 wire \logix.ram_r[1153] ;
 wire \logix.ram_r[1154] ;
 wire \logix.ram_r[1155] ;
 wire \logix.ram_r[1156] ;
 wire \logix.ram_r[1157] ;
 wire \logix.ram_r[1158] ;
 wire \logix.ram_r[1159] ;
 wire \logix.ram_r[115] ;
 wire \logix.ram_r[1160] ;
 wire \logix.ram_r[1161] ;
 wire \logix.ram_r[1162] ;
 wire \logix.ram_r[1163] ;
 wire \logix.ram_r[1164] ;
 wire \logix.ram_r[1165] ;
 wire \logix.ram_r[1166] ;
 wire \logix.ram_r[1167] ;
 wire \logix.ram_r[1168] ;
 wire \logix.ram_r[1169] ;
 wire \logix.ram_r[116] ;
 wire \logix.ram_r[1170] ;
 wire \logix.ram_r[1171] ;
 wire \logix.ram_r[1172] ;
 wire \logix.ram_r[1173] ;
 wire \logix.ram_r[1174] ;
 wire \logix.ram_r[1175] ;
 wire \logix.ram_r[1176] ;
 wire \logix.ram_r[1177] ;
 wire \logix.ram_r[1178] ;
 wire \logix.ram_r[1179] ;
 wire \logix.ram_r[117] ;
 wire \logix.ram_r[1180] ;
 wire \logix.ram_r[1181] ;
 wire \logix.ram_r[1182] ;
 wire \logix.ram_r[1183] ;
 wire \logix.ram_r[1184] ;
 wire \logix.ram_r[1185] ;
 wire \logix.ram_r[1186] ;
 wire \logix.ram_r[1187] ;
 wire \logix.ram_r[1188] ;
 wire \logix.ram_r[1189] ;
 wire \logix.ram_r[118] ;
 wire \logix.ram_r[1190] ;
 wire \logix.ram_r[1191] ;
 wire \logix.ram_r[1192] ;
 wire \logix.ram_r[1193] ;
 wire \logix.ram_r[1194] ;
 wire \logix.ram_r[1195] ;
 wire \logix.ram_r[1196] ;
 wire \logix.ram_r[1197] ;
 wire \logix.ram_r[1198] ;
 wire \logix.ram_r[1199] ;
 wire \logix.ram_r[119] ;
 wire \logix.ram_r[11] ;
 wire \logix.ram_r[1200] ;
 wire \logix.ram_r[1201] ;
 wire \logix.ram_r[1202] ;
 wire \logix.ram_r[1203] ;
 wire \logix.ram_r[1204] ;
 wire \logix.ram_r[1205] ;
 wire \logix.ram_r[1206] ;
 wire \logix.ram_r[1207] ;
 wire \logix.ram_r[1208] ;
 wire \logix.ram_r[1209] ;
 wire \logix.ram_r[120] ;
 wire \logix.ram_r[1210] ;
 wire \logix.ram_r[1211] ;
 wire \logix.ram_r[1212] ;
 wire \logix.ram_r[1213] ;
 wire \logix.ram_r[1214] ;
 wire \logix.ram_r[1215] ;
 wire \logix.ram_r[1216] ;
 wire \logix.ram_r[1217] ;
 wire \logix.ram_r[1218] ;
 wire \logix.ram_r[1219] ;
 wire \logix.ram_r[121] ;
 wire \logix.ram_r[1220] ;
 wire \logix.ram_r[1221] ;
 wire \logix.ram_r[1222] ;
 wire \logix.ram_r[1223] ;
 wire \logix.ram_r[1224] ;
 wire \logix.ram_r[1225] ;
 wire \logix.ram_r[1226] ;
 wire \logix.ram_r[1227] ;
 wire \logix.ram_r[1228] ;
 wire \logix.ram_r[1229] ;
 wire \logix.ram_r[122] ;
 wire \logix.ram_r[1230] ;
 wire \logix.ram_r[1231] ;
 wire \logix.ram_r[1232] ;
 wire \logix.ram_r[1233] ;
 wire \logix.ram_r[1234] ;
 wire \logix.ram_r[1235] ;
 wire \logix.ram_r[1236] ;
 wire \logix.ram_r[1237] ;
 wire \logix.ram_r[1238] ;
 wire \logix.ram_r[1239] ;
 wire \logix.ram_r[123] ;
 wire \logix.ram_r[1240] ;
 wire \logix.ram_r[1241] ;
 wire \logix.ram_r[1242] ;
 wire \logix.ram_r[1243] ;
 wire \logix.ram_r[1244] ;
 wire \logix.ram_r[1245] ;
 wire \logix.ram_r[1246] ;
 wire \logix.ram_r[1247] ;
 wire \logix.ram_r[1248] ;
 wire \logix.ram_r[1249] ;
 wire \logix.ram_r[124] ;
 wire \logix.ram_r[1250] ;
 wire \logix.ram_r[1251] ;
 wire \logix.ram_r[1252] ;
 wire \logix.ram_r[1253] ;
 wire \logix.ram_r[1254] ;
 wire \logix.ram_r[1255] ;
 wire \logix.ram_r[1256] ;
 wire \logix.ram_r[1257] ;
 wire \logix.ram_r[1258] ;
 wire \logix.ram_r[1259] ;
 wire \logix.ram_r[125] ;
 wire \logix.ram_r[1260] ;
 wire \logix.ram_r[1261] ;
 wire \logix.ram_r[1262] ;
 wire \logix.ram_r[1263] ;
 wire \logix.ram_r[1264] ;
 wire \logix.ram_r[1265] ;
 wire \logix.ram_r[1266] ;
 wire \logix.ram_r[1267] ;
 wire \logix.ram_r[1268] ;
 wire \logix.ram_r[1269] ;
 wire \logix.ram_r[126] ;
 wire \logix.ram_r[1270] ;
 wire \logix.ram_r[1271] ;
 wire \logix.ram_r[1272] ;
 wire \logix.ram_r[1273] ;
 wire \logix.ram_r[1274] ;
 wire \logix.ram_r[1275] ;
 wire \logix.ram_r[1276] ;
 wire \logix.ram_r[1277] ;
 wire \logix.ram_r[1278] ;
 wire \logix.ram_r[1279] ;
 wire \logix.ram_r[127] ;
 wire \logix.ram_r[1280] ;
 wire \logix.ram_r[1281] ;
 wire \logix.ram_r[1282] ;
 wire \logix.ram_r[1283] ;
 wire \logix.ram_r[1284] ;
 wire \logix.ram_r[1285] ;
 wire \logix.ram_r[1286] ;
 wire \logix.ram_r[1287] ;
 wire \logix.ram_r[1288] ;
 wire \logix.ram_r[1289] ;
 wire \logix.ram_r[128] ;
 wire \logix.ram_r[1290] ;
 wire \logix.ram_r[1291] ;
 wire \logix.ram_r[1292] ;
 wire \logix.ram_r[1293] ;
 wire \logix.ram_r[1294] ;
 wire \logix.ram_r[1295] ;
 wire \logix.ram_r[1296] ;
 wire \logix.ram_r[1297] ;
 wire \logix.ram_r[1298] ;
 wire \logix.ram_r[1299] ;
 wire \logix.ram_r[129] ;
 wire \logix.ram_r[12] ;
 wire \logix.ram_r[1300] ;
 wire \logix.ram_r[1301] ;
 wire \logix.ram_r[1302] ;
 wire \logix.ram_r[1303] ;
 wire \logix.ram_r[1304] ;
 wire \logix.ram_r[1305] ;
 wire \logix.ram_r[1306] ;
 wire \logix.ram_r[1307] ;
 wire \logix.ram_r[1308] ;
 wire \logix.ram_r[1309] ;
 wire \logix.ram_r[130] ;
 wire \logix.ram_r[1310] ;
 wire \logix.ram_r[1311] ;
 wire \logix.ram_r[1312] ;
 wire \logix.ram_r[1313] ;
 wire \logix.ram_r[1314] ;
 wire \logix.ram_r[1315] ;
 wire \logix.ram_r[1316] ;
 wire \logix.ram_r[1317] ;
 wire \logix.ram_r[1318] ;
 wire \logix.ram_r[1319] ;
 wire \logix.ram_r[131] ;
 wire \logix.ram_r[1320] ;
 wire \logix.ram_r[1321] ;
 wire \logix.ram_r[1322] ;
 wire \logix.ram_r[1323] ;
 wire \logix.ram_r[1324] ;
 wire \logix.ram_r[1325] ;
 wire \logix.ram_r[1326] ;
 wire \logix.ram_r[1327] ;
 wire \logix.ram_r[1328] ;
 wire \logix.ram_r[1329] ;
 wire \logix.ram_r[132] ;
 wire \logix.ram_r[1330] ;
 wire \logix.ram_r[1331] ;
 wire \logix.ram_r[1332] ;
 wire \logix.ram_r[1333] ;
 wire \logix.ram_r[1334] ;
 wire \logix.ram_r[1335] ;
 wire \logix.ram_r[1336] ;
 wire \logix.ram_r[1337] ;
 wire \logix.ram_r[1338] ;
 wire \logix.ram_r[1339] ;
 wire \logix.ram_r[133] ;
 wire \logix.ram_r[1340] ;
 wire \logix.ram_r[1341] ;
 wire \logix.ram_r[1342] ;
 wire \logix.ram_r[1343] ;
 wire \logix.ram_r[1344] ;
 wire \logix.ram_r[1345] ;
 wire \logix.ram_r[1346] ;
 wire \logix.ram_r[1347] ;
 wire \logix.ram_r[1348] ;
 wire \logix.ram_r[1349] ;
 wire \logix.ram_r[134] ;
 wire \logix.ram_r[1350] ;
 wire \logix.ram_r[1351] ;
 wire \logix.ram_r[1352] ;
 wire \logix.ram_r[1353] ;
 wire \logix.ram_r[1354] ;
 wire \logix.ram_r[1355] ;
 wire \logix.ram_r[1356] ;
 wire \logix.ram_r[1357] ;
 wire \logix.ram_r[1358] ;
 wire \logix.ram_r[1359] ;
 wire \logix.ram_r[135] ;
 wire \logix.ram_r[1360] ;
 wire \logix.ram_r[1361] ;
 wire \logix.ram_r[1362] ;
 wire \logix.ram_r[1363] ;
 wire \logix.ram_r[1364] ;
 wire \logix.ram_r[1365] ;
 wire \logix.ram_r[1366] ;
 wire \logix.ram_r[1367] ;
 wire \logix.ram_r[1368] ;
 wire \logix.ram_r[1369] ;
 wire \logix.ram_r[136] ;
 wire \logix.ram_r[1370] ;
 wire \logix.ram_r[1371] ;
 wire \logix.ram_r[1372] ;
 wire \logix.ram_r[1373] ;
 wire \logix.ram_r[1374] ;
 wire \logix.ram_r[1375] ;
 wire \logix.ram_r[1376] ;
 wire \logix.ram_r[1377] ;
 wire \logix.ram_r[1378] ;
 wire \logix.ram_r[1379] ;
 wire \logix.ram_r[137] ;
 wire \logix.ram_r[1380] ;
 wire \logix.ram_r[1381] ;
 wire \logix.ram_r[1382] ;
 wire \logix.ram_r[1383] ;
 wire \logix.ram_r[1384] ;
 wire \logix.ram_r[1385] ;
 wire \logix.ram_r[1386] ;
 wire \logix.ram_r[1387] ;
 wire \logix.ram_r[1388] ;
 wire \logix.ram_r[1389] ;
 wire \logix.ram_r[138] ;
 wire \logix.ram_r[1390] ;
 wire \logix.ram_r[1391] ;
 wire \logix.ram_r[1392] ;
 wire \logix.ram_r[1393] ;
 wire \logix.ram_r[1394] ;
 wire \logix.ram_r[1395] ;
 wire \logix.ram_r[1396] ;
 wire \logix.ram_r[1397] ;
 wire \logix.ram_r[1398] ;
 wire \logix.ram_r[1399] ;
 wire \logix.ram_r[139] ;
 wire \logix.ram_r[13] ;
 wire \logix.ram_r[1400] ;
 wire \logix.ram_r[1401] ;
 wire \logix.ram_r[1402] ;
 wire \logix.ram_r[1403] ;
 wire \logix.ram_r[1404] ;
 wire \logix.ram_r[1405] ;
 wire \logix.ram_r[1406] ;
 wire \logix.ram_r[1407] ;
 wire \logix.ram_r[1408] ;
 wire \logix.ram_r[1409] ;
 wire \logix.ram_r[140] ;
 wire \logix.ram_r[1410] ;
 wire \logix.ram_r[1411] ;
 wire \logix.ram_r[1412] ;
 wire \logix.ram_r[1413] ;
 wire \logix.ram_r[1414] ;
 wire \logix.ram_r[1415] ;
 wire \logix.ram_r[1416] ;
 wire \logix.ram_r[1417] ;
 wire \logix.ram_r[1418] ;
 wire \logix.ram_r[1419] ;
 wire \logix.ram_r[141] ;
 wire \logix.ram_r[1420] ;
 wire \logix.ram_r[1421] ;
 wire \logix.ram_r[1422] ;
 wire \logix.ram_r[1423] ;
 wire \logix.ram_r[1424] ;
 wire \logix.ram_r[1425] ;
 wire \logix.ram_r[1426] ;
 wire \logix.ram_r[1427] ;
 wire \logix.ram_r[1428] ;
 wire \logix.ram_r[1429] ;
 wire \logix.ram_r[142] ;
 wire \logix.ram_r[1430] ;
 wire \logix.ram_r[1431] ;
 wire \logix.ram_r[1432] ;
 wire \logix.ram_r[1433] ;
 wire \logix.ram_r[1434] ;
 wire \logix.ram_r[1435] ;
 wire \logix.ram_r[1436] ;
 wire \logix.ram_r[1437] ;
 wire \logix.ram_r[1438] ;
 wire \logix.ram_r[1439] ;
 wire \logix.ram_r[143] ;
 wire \logix.ram_r[1440] ;
 wire \logix.ram_r[1441] ;
 wire \logix.ram_r[1442] ;
 wire \logix.ram_r[1443] ;
 wire \logix.ram_r[1444] ;
 wire \logix.ram_r[1445] ;
 wire \logix.ram_r[1446] ;
 wire \logix.ram_r[1447] ;
 wire \logix.ram_r[1448] ;
 wire \logix.ram_r[1449] ;
 wire \logix.ram_r[144] ;
 wire \logix.ram_r[1450] ;
 wire \logix.ram_r[1451] ;
 wire \logix.ram_r[1452] ;
 wire \logix.ram_r[1453] ;
 wire \logix.ram_r[1454] ;
 wire \logix.ram_r[1455] ;
 wire \logix.ram_r[1456] ;
 wire \logix.ram_r[1457] ;
 wire \logix.ram_r[1458] ;
 wire \logix.ram_r[1459] ;
 wire \logix.ram_r[145] ;
 wire \logix.ram_r[1460] ;
 wire \logix.ram_r[1461] ;
 wire \logix.ram_r[1462] ;
 wire \logix.ram_r[1463] ;
 wire \logix.ram_r[1464] ;
 wire \logix.ram_r[1465] ;
 wire \logix.ram_r[1466] ;
 wire \logix.ram_r[1467] ;
 wire \logix.ram_r[1468] ;
 wire \logix.ram_r[1469] ;
 wire \logix.ram_r[146] ;
 wire \logix.ram_r[1470] ;
 wire \logix.ram_r[1471] ;
 wire \logix.ram_r[1472] ;
 wire \logix.ram_r[1473] ;
 wire \logix.ram_r[1474] ;
 wire \logix.ram_r[1475] ;
 wire \logix.ram_r[1476] ;
 wire \logix.ram_r[1477] ;
 wire \logix.ram_r[1478] ;
 wire \logix.ram_r[1479] ;
 wire \logix.ram_r[147] ;
 wire \logix.ram_r[1480] ;
 wire \logix.ram_r[1481] ;
 wire \logix.ram_r[1482] ;
 wire \logix.ram_r[1483] ;
 wire \logix.ram_r[1484] ;
 wire \logix.ram_r[1485] ;
 wire \logix.ram_r[1486] ;
 wire \logix.ram_r[1487] ;
 wire \logix.ram_r[1488] ;
 wire \logix.ram_r[1489] ;
 wire \logix.ram_r[148] ;
 wire \logix.ram_r[1490] ;
 wire \logix.ram_r[1491] ;
 wire \logix.ram_r[1492] ;
 wire \logix.ram_r[1493] ;
 wire \logix.ram_r[1494] ;
 wire \logix.ram_r[1495] ;
 wire \logix.ram_r[1496] ;
 wire \logix.ram_r[1497] ;
 wire \logix.ram_r[1498] ;
 wire \logix.ram_r[1499] ;
 wire \logix.ram_r[149] ;
 wire \logix.ram_r[14] ;
 wire \logix.ram_r[1500] ;
 wire \logix.ram_r[1501] ;
 wire \logix.ram_r[1502] ;
 wire \logix.ram_r[1503] ;
 wire \logix.ram_r[1504] ;
 wire \logix.ram_r[1505] ;
 wire \logix.ram_r[1506] ;
 wire \logix.ram_r[1507] ;
 wire \logix.ram_r[1508] ;
 wire \logix.ram_r[1509] ;
 wire \logix.ram_r[150] ;
 wire \logix.ram_r[1510] ;
 wire \logix.ram_r[1511] ;
 wire \logix.ram_r[1512] ;
 wire \logix.ram_r[1513] ;
 wire \logix.ram_r[1514] ;
 wire \logix.ram_r[1515] ;
 wire \logix.ram_r[1516] ;
 wire \logix.ram_r[1517] ;
 wire \logix.ram_r[1518] ;
 wire \logix.ram_r[1519] ;
 wire \logix.ram_r[151] ;
 wire \logix.ram_r[1520] ;
 wire \logix.ram_r[1521] ;
 wire \logix.ram_r[1522] ;
 wire \logix.ram_r[1523] ;
 wire \logix.ram_r[1524] ;
 wire \logix.ram_r[1525] ;
 wire \logix.ram_r[1526] ;
 wire \logix.ram_r[1527] ;
 wire \logix.ram_r[1528] ;
 wire \logix.ram_r[1529] ;
 wire \logix.ram_r[152] ;
 wire \logix.ram_r[1530] ;
 wire \logix.ram_r[1531] ;
 wire \logix.ram_r[1532] ;
 wire \logix.ram_r[1533] ;
 wire \logix.ram_r[1534] ;
 wire \logix.ram_r[1535] ;
 wire \logix.ram_r[1536] ;
 wire \logix.ram_r[1537] ;
 wire \logix.ram_r[1538] ;
 wire \logix.ram_r[1539] ;
 wire \logix.ram_r[153] ;
 wire \logix.ram_r[1540] ;
 wire \logix.ram_r[1541] ;
 wire \logix.ram_r[1542] ;
 wire \logix.ram_r[1543] ;
 wire \logix.ram_r[1544] ;
 wire \logix.ram_r[1545] ;
 wire \logix.ram_r[1546] ;
 wire \logix.ram_r[1547] ;
 wire \logix.ram_r[1548] ;
 wire \logix.ram_r[1549] ;
 wire \logix.ram_r[154] ;
 wire \logix.ram_r[1550] ;
 wire \logix.ram_r[1551] ;
 wire \logix.ram_r[1552] ;
 wire \logix.ram_r[1553] ;
 wire \logix.ram_r[1554] ;
 wire \logix.ram_r[1555] ;
 wire \logix.ram_r[1556] ;
 wire \logix.ram_r[1557] ;
 wire \logix.ram_r[1558] ;
 wire \logix.ram_r[1559] ;
 wire \logix.ram_r[155] ;
 wire \logix.ram_r[1560] ;
 wire \logix.ram_r[1561] ;
 wire \logix.ram_r[1562] ;
 wire \logix.ram_r[1563] ;
 wire \logix.ram_r[1564] ;
 wire \logix.ram_r[1565] ;
 wire \logix.ram_r[1566] ;
 wire \logix.ram_r[1567] ;
 wire \logix.ram_r[1568] ;
 wire \logix.ram_r[1569] ;
 wire \logix.ram_r[156] ;
 wire \logix.ram_r[1570] ;
 wire \logix.ram_r[1571] ;
 wire \logix.ram_r[1572] ;
 wire \logix.ram_r[1573] ;
 wire \logix.ram_r[1574] ;
 wire \logix.ram_r[1575] ;
 wire \logix.ram_r[1576] ;
 wire \logix.ram_r[1577] ;
 wire \logix.ram_r[1578] ;
 wire \logix.ram_r[1579] ;
 wire \logix.ram_r[157] ;
 wire \logix.ram_r[1580] ;
 wire \logix.ram_r[1581] ;
 wire \logix.ram_r[1582] ;
 wire \logix.ram_r[1583] ;
 wire \logix.ram_r[1584] ;
 wire \logix.ram_r[1585] ;
 wire \logix.ram_r[1586] ;
 wire \logix.ram_r[1587] ;
 wire \logix.ram_r[1588] ;
 wire \logix.ram_r[1589] ;
 wire \logix.ram_r[158] ;
 wire \logix.ram_r[1590] ;
 wire \logix.ram_r[1591] ;
 wire \logix.ram_r[1592] ;
 wire \logix.ram_r[1593] ;
 wire \logix.ram_r[1594] ;
 wire \logix.ram_r[1595] ;
 wire \logix.ram_r[1596] ;
 wire \logix.ram_r[1597] ;
 wire \logix.ram_r[1598] ;
 wire \logix.ram_r[1599] ;
 wire \logix.ram_r[159] ;
 wire \logix.ram_r[15] ;
 wire \logix.ram_r[1600] ;
 wire \logix.ram_r[1601] ;
 wire \logix.ram_r[1602] ;
 wire \logix.ram_r[1603] ;
 wire \logix.ram_r[1604] ;
 wire \logix.ram_r[1605] ;
 wire \logix.ram_r[1606] ;
 wire \logix.ram_r[1607] ;
 wire \logix.ram_r[1608] ;
 wire \logix.ram_r[1609] ;
 wire \logix.ram_r[160] ;
 wire \logix.ram_r[1610] ;
 wire \logix.ram_r[1611] ;
 wire \logix.ram_r[1612] ;
 wire \logix.ram_r[1613] ;
 wire \logix.ram_r[1614] ;
 wire \logix.ram_r[1615] ;
 wire \logix.ram_r[1616] ;
 wire \logix.ram_r[1617] ;
 wire \logix.ram_r[1618] ;
 wire \logix.ram_r[1619] ;
 wire \logix.ram_r[161] ;
 wire \logix.ram_r[1620] ;
 wire \logix.ram_r[1621] ;
 wire \logix.ram_r[1622] ;
 wire \logix.ram_r[1623] ;
 wire \logix.ram_r[1624] ;
 wire \logix.ram_r[1625] ;
 wire \logix.ram_r[1626] ;
 wire \logix.ram_r[1627] ;
 wire \logix.ram_r[1628] ;
 wire \logix.ram_r[1629] ;
 wire \logix.ram_r[162] ;
 wire \logix.ram_r[1630] ;
 wire \logix.ram_r[1631] ;
 wire \logix.ram_r[1632] ;
 wire \logix.ram_r[1633] ;
 wire \logix.ram_r[1634] ;
 wire \logix.ram_r[1635] ;
 wire \logix.ram_r[1636] ;
 wire \logix.ram_r[1637] ;
 wire \logix.ram_r[1638] ;
 wire \logix.ram_r[1639] ;
 wire \logix.ram_r[163] ;
 wire \logix.ram_r[1640] ;
 wire \logix.ram_r[1641] ;
 wire \logix.ram_r[1642] ;
 wire \logix.ram_r[1643] ;
 wire \logix.ram_r[1644] ;
 wire \logix.ram_r[1645] ;
 wire \logix.ram_r[1646] ;
 wire \logix.ram_r[1647] ;
 wire \logix.ram_r[1648] ;
 wire \logix.ram_r[1649] ;
 wire \logix.ram_r[164] ;
 wire \logix.ram_r[1650] ;
 wire \logix.ram_r[1651] ;
 wire \logix.ram_r[1652] ;
 wire \logix.ram_r[1653] ;
 wire \logix.ram_r[1654] ;
 wire \logix.ram_r[1655] ;
 wire \logix.ram_r[1656] ;
 wire \logix.ram_r[1657] ;
 wire \logix.ram_r[1658] ;
 wire \logix.ram_r[1659] ;
 wire \logix.ram_r[165] ;
 wire \logix.ram_r[1660] ;
 wire \logix.ram_r[1661] ;
 wire \logix.ram_r[1662] ;
 wire \logix.ram_r[1663] ;
 wire \logix.ram_r[1664] ;
 wire \logix.ram_r[1665] ;
 wire \logix.ram_r[1666] ;
 wire \logix.ram_r[1667] ;
 wire \logix.ram_r[1668] ;
 wire \logix.ram_r[1669] ;
 wire \logix.ram_r[166] ;
 wire \logix.ram_r[1670] ;
 wire \logix.ram_r[1671] ;
 wire \logix.ram_r[1672] ;
 wire \logix.ram_r[1673] ;
 wire \logix.ram_r[1674] ;
 wire \logix.ram_r[1675] ;
 wire \logix.ram_r[1676] ;
 wire \logix.ram_r[1677] ;
 wire \logix.ram_r[1678] ;
 wire \logix.ram_r[1679] ;
 wire \logix.ram_r[167] ;
 wire \logix.ram_r[1680] ;
 wire \logix.ram_r[1681] ;
 wire \logix.ram_r[1682] ;
 wire \logix.ram_r[1683] ;
 wire \logix.ram_r[1684] ;
 wire \logix.ram_r[1685] ;
 wire \logix.ram_r[1686] ;
 wire \logix.ram_r[1687] ;
 wire \logix.ram_r[1688] ;
 wire \logix.ram_r[1689] ;
 wire \logix.ram_r[168] ;
 wire \logix.ram_r[1690] ;
 wire \logix.ram_r[1691] ;
 wire \logix.ram_r[1692] ;
 wire \logix.ram_r[1693] ;
 wire \logix.ram_r[1694] ;
 wire \logix.ram_r[1695] ;
 wire \logix.ram_r[1696] ;
 wire \logix.ram_r[1697] ;
 wire \logix.ram_r[1698] ;
 wire \logix.ram_r[1699] ;
 wire \logix.ram_r[169] ;
 wire \logix.ram_r[16] ;
 wire \logix.ram_r[1700] ;
 wire \logix.ram_r[1701] ;
 wire \logix.ram_r[1702] ;
 wire \logix.ram_r[1703] ;
 wire \logix.ram_r[1704] ;
 wire \logix.ram_r[1705] ;
 wire \logix.ram_r[1706] ;
 wire \logix.ram_r[1707] ;
 wire \logix.ram_r[1708] ;
 wire \logix.ram_r[1709] ;
 wire \logix.ram_r[170] ;
 wire \logix.ram_r[1710] ;
 wire \logix.ram_r[1711] ;
 wire \logix.ram_r[1712] ;
 wire \logix.ram_r[1713] ;
 wire \logix.ram_r[1714] ;
 wire \logix.ram_r[1715] ;
 wire \logix.ram_r[1716] ;
 wire \logix.ram_r[1717] ;
 wire \logix.ram_r[1718] ;
 wire \logix.ram_r[1719] ;
 wire \logix.ram_r[171] ;
 wire \logix.ram_r[1720] ;
 wire \logix.ram_r[1721] ;
 wire \logix.ram_r[1722] ;
 wire \logix.ram_r[1723] ;
 wire \logix.ram_r[1724] ;
 wire \logix.ram_r[1725] ;
 wire \logix.ram_r[1726] ;
 wire \logix.ram_r[1727] ;
 wire \logix.ram_r[1728] ;
 wire \logix.ram_r[1729] ;
 wire \logix.ram_r[172] ;
 wire \logix.ram_r[1730] ;
 wire \logix.ram_r[1731] ;
 wire \logix.ram_r[1732] ;
 wire \logix.ram_r[1733] ;
 wire \logix.ram_r[1734] ;
 wire \logix.ram_r[1735] ;
 wire \logix.ram_r[1736] ;
 wire \logix.ram_r[1737] ;
 wire \logix.ram_r[1738] ;
 wire \logix.ram_r[1739] ;
 wire \logix.ram_r[173] ;
 wire \logix.ram_r[1740] ;
 wire \logix.ram_r[1741] ;
 wire \logix.ram_r[1742] ;
 wire \logix.ram_r[1743] ;
 wire \logix.ram_r[1744] ;
 wire \logix.ram_r[1745] ;
 wire \logix.ram_r[1746] ;
 wire \logix.ram_r[1747] ;
 wire \logix.ram_r[1748] ;
 wire \logix.ram_r[1749] ;
 wire \logix.ram_r[174] ;
 wire \logix.ram_r[1750] ;
 wire \logix.ram_r[1751] ;
 wire \logix.ram_r[1752] ;
 wire \logix.ram_r[1753] ;
 wire \logix.ram_r[1754] ;
 wire \logix.ram_r[1755] ;
 wire \logix.ram_r[1756] ;
 wire \logix.ram_r[1757] ;
 wire \logix.ram_r[1758] ;
 wire \logix.ram_r[1759] ;
 wire \logix.ram_r[175] ;
 wire \logix.ram_r[1760] ;
 wire \logix.ram_r[1761] ;
 wire \logix.ram_r[1762] ;
 wire \logix.ram_r[1763] ;
 wire \logix.ram_r[1764] ;
 wire \logix.ram_r[1765] ;
 wire \logix.ram_r[1766] ;
 wire \logix.ram_r[1767] ;
 wire \logix.ram_r[1768] ;
 wire \logix.ram_r[1769] ;
 wire \logix.ram_r[176] ;
 wire \logix.ram_r[1770] ;
 wire \logix.ram_r[1771] ;
 wire \logix.ram_r[1772] ;
 wire \logix.ram_r[1773] ;
 wire \logix.ram_r[1774] ;
 wire \logix.ram_r[1775] ;
 wire \logix.ram_r[1776] ;
 wire \logix.ram_r[1777] ;
 wire \logix.ram_r[1778] ;
 wire \logix.ram_r[1779] ;
 wire \logix.ram_r[177] ;
 wire \logix.ram_r[1780] ;
 wire \logix.ram_r[1781] ;
 wire \logix.ram_r[1782] ;
 wire \logix.ram_r[1783] ;
 wire \logix.ram_r[1784] ;
 wire \logix.ram_r[1785] ;
 wire \logix.ram_r[1786] ;
 wire \logix.ram_r[1787] ;
 wire \logix.ram_r[1788] ;
 wire \logix.ram_r[1789] ;
 wire \logix.ram_r[178] ;
 wire \logix.ram_r[1790] ;
 wire \logix.ram_r[1791] ;
 wire \logix.ram_r[1792] ;
 wire \logix.ram_r[1793] ;
 wire \logix.ram_r[1794] ;
 wire \logix.ram_r[1795] ;
 wire \logix.ram_r[1796] ;
 wire \logix.ram_r[1797] ;
 wire \logix.ram_r[1798] ;
 wire \logix.ram_r[1799] ;
 wire \logix.ram_r[179] ;
 wire \logix.ram_r[17] ;
 wire \logix.ram_r[1800] ;
 wire \logix.ram_r[1801] ;
 wire \logix.ram_r[1802] ;
 wire \logix.ram_r[1803] ;
 wire \logix.ram_r[1804] ;
 wire \logix.ram_r[1805] ;
 wire \logix.ram_r[1806] ;
 wire \logix.ram_r[1807] ;
 wire \logix.ram_r[1808] ;
 wire \logix.ram_r[1809] ;
 wire \logix.ram_r[180] ;
 wire \logix.ram_r[1810] ;
 wire \logix.ram_r[1811] ;
 wire \logix.ram_r[1812] ;
 wire \logix.ram_r[1813] ;
 wire \logix.ram_r[1814] ;
 wire \logix.ram_r[1815] ;
 wire \logix.ram_r[1816] ;
 wire \logix.ram_r[1817] ;
 wire \logix.ram_r[1818] ;
 wire \logix.ram_r[1819] ;
 wire \logix.ram_r[181] ;
 wire \logix.ram_r[1820] ;
 wire \logix.ram_r[1821] ;
 wire \logix.ram_r[1822] ;
 wire \logix.ram_r[1823] ;
 wire \logix.ram_r[1824] ;
 wire \logix.ram_r[1825] ;
 wire \logix.ram_r[1826] ;
 wire \logix.ram_r[1827] ;
 wire \logix.ram_r[1828] ;
 wire \logix.ram_r[1829] ;
 wire \logix.ram_r[182] ;
 wire \logix.ram_r[1830] ;
 wire \logix.ram_r[1831] ;
 wire \logix.ram_r[1832] ;
 wire \logix.ram_r[1833] ;
 wire \logix.ram_r[1834] ;
 wire \logix.ram_r[1835] ;
 wire \logix.ram_r[1836] ;
 wire \logix.ram_r[1837] ;
 wire \logix.ram_r[1838] ;
 wire \logix.ram_r[1839] ;
 wire \logix.ram_r[183] ;
 wire \logix.ram_r[1840] ;
 wire \logix.ram_r[1841] ;
 wire \logix.ram_r[1842] ;
 wire \logix.ram_r[1843] ;
 wire \logix.ram_r[1844] ;
 wire \logix.ram_r[1845] ;
 wire \logix.ram_r[1846] ;
 wire \logix.ram_r[1847] ;
 wire \logix.ram_r[1848] ;
 wire \logix.ram_r[1849] ;
 wire \logix.ram_r[184] ;
 wire \logix.ram_r[1850] ;
 wire \logix.ram_r[1851] ;
 wire \logix.ram_r[1852] ;
 wire \logix.ram_r[1853] ;
 wire \logix.ram_r[1854] ;
 wire \logix.ram_r[1855] ;
 wire \logix.ram_r[1856] ;
 wire \logix.ram_r[1857] ;
 wire \logix.ram_r[1858] ;
 wire \logix.ram_r[1859] ;
 wire \logix.ram_r[185] ;
 wire \logix.ram_r[1860] ;
 wire \logix.ram_r[1861] ;
 wire \logix.ram_r[1862] ;
 wire \logix.ram_r[1863] ;
 wire \logix.ram_r[1864] ;
 wire \logix.ram_r[1865] ;
 wire \logix.ram_r[1866] ;
 wire \logix.ram_r[1867] ;
 wire \logix.ram_r[1868] ;
 wire \logix.ram_r[1869] ;
 wire \logix.ram_r[186] ;
 wire \logix.ram_r[1870] ;
 wire \logix.ram_r[1871] ;
 wire \logix.ram_r[1872] ;
 wire \logix.ram_r[1873] ;
 wire \logix.ram_r[1874] ;
 wire \logix.ram_r[1875] ;
 wire \logix.ram_r[1876] ;
 wire \logix.ram_r[1877] ;
 wire \logix.ram_r[1878] ;
 wire \logix.ram_r[1879] ;
 wire \logix.ram_r[187] ;
 wire \logix.ram_r[1880] ;
 wire \logix.ram_r[1881] ;
 wire \logix.ram_r[1882] ;
 wire \logix.ram_r[1883] ;
 wire \logix.ram_r[1884] ;
 wire \logix.ram_r[1885] ;
 wire \logix.ram_r[1886] ;
 wire \logix.ram_r[1887] ;
 wire \logix.ram_r[1888] ;
 wire \logix.ram_r[1889] ;
 wire \logix.ram_r[188] ;
 wire \logix.ram_r[1890] ;
 wire \logix.ram_r[1891] ;
 wire \logix.ram_r[1892] ;
 wire \logix.ram_r[1893] ;
 wire \logix.ram_r[1894] ;
 wire \logix.ram_r[1895] ;
 wire \logix.ram_r[1896] ;
 wire \logix.ram_r[1897] ;
 wire \logix.ram_r[1898] ;
 wire \logix.ram_r[1899] ;
 wire \logix.ram_r[189] ;
 wire \logix.ram_r[18] ;
 wire \logix.ram_r[1900] ;
 wire \logix.ram_r[1901] ;
 wire \logix.ram_r[1902] ;
 wire \logix.ram_r[1903] ;
 wire \logix.ram_r[1904] ;
 wire \logix.ram_r[1905] ;
 wire \logix.ram_r[1906] ;
 wire \logix.ram_r[1907] ;
 wire \logix.ram_r[1908] ;
 wire \logix.ram_r[1909] ;
 wire \logix.ram_r[190] ;
 wire \logix.ram_r[1910] ;
 wire \logix.ram_r[1911] ;
 wire \logix.ram_r[1912] ;
 wire \logix.ram_r[1913] ;
 wire \logix.ram_r[1914] ;
 wire \logix.ram_r[1915] ;
 wire \logix.ram_r[1916] ;
 wire \logix.ram_r[1917] ;
 wire \logix.ram_r[1918] ;
 wire \logix.ram_r[1919] ;
 wire \logix.ram_r[191] ;
 wire \logix.ram_r[1920] ;
 wire \logix.ram_r[1921] ;
 wire \logix.ram_r[1922] ;
 wire \logix.ram_r[1923] ;
 wire \logix.ram_r[1924] ;
 wire \logix.ram_r[1925] ;
 wire \logix.ram_r[1926] ;
 wire \logix.ram_r[1927] ;
 wire \logix.ram_r[1928] ;
 wire \logix.ram_r[1929] ;
 wire \logix.ram_r[192] ;
 wire \logix.ram_r[1930] ;
 wire \logix.ram_r[1931] ;
 wire \logix.ram_r[1932] ;
 wire \logix.ram_r[1933] ;
 wire \logix.ram_r[1934] ;
 wire \logix.ram_r[1935] ;
 wire \logix.ram_r[1936] ;
 wire \logix.ram_r[1937] ;
 wire \logix.ram_r[1938] ;
 wire \logix.ram_r[1939] ;
 wire \logix.ram_r[193] ;
 wire \logix.ram_r[1940] ;
 wire \logix.ram_r[1941] ;
 wire \logix.ram_r[1942] ;
 wire \logix.ram_r[1943] ;
 wire \logix.ram_r[1944] ;
 wire \logix.ram_r[1945] ;
 wire \logix.ram_r[1946] ;
 wire \logix.ram_r[1947] ;
 wire \logix.ram_r[1948] ;
 wire \logix.ram_r[1949] ;
 wire \logix.ram_r[194] ;
 wire \logix.ram_r[1950] ;
 wire \logix.ram_r[1951] ;
 wire \logix.ram_r[1952] ;
 wire \logix.ram_r[1953] ;
 wire \logix.ram_r[1954] ;
 wire \logix.ram_r[1955] ;
 wire \logix.ram_r[1956] ;
 wire \logix.ram_r[1957] ;
 wire \logix.ram_r[1958] ;
 wire \logix.ram_r[1959] ;
 wire \logix.ram_r[195] ;
 wire \logix.ram_r[1960] ;
 wire \logix.ram_r[1961] ;
 wire \logix.ram_r[1962] ;
 wire \logix.ram_r[1963] ;
 wire \logix.ram_r[1964] ;
 wire \logix.ram_r[1965] ;
 wire \logix.ram_r[1966] ;
 wire \logix.ram_r[1967] ;
 wire \logix.ram_r[1968] ;
 wire \logix.ram_r[1969] ;
 wire \logix.ram_r[196] ;
 wire \logix.ram_r[1970] ;
 wire \logix.ram_r[1971] ;
 wire \logix.ram_r[1972] ;
 wire \logix.ram_r[1973] ;
 wire \logix.ram_r[1974] ;
 wire \logix.ram_r[1975] ;
 wire \logix.ram_r[1976] ;
 wire \logix.ram_r[1977] ;
 wire \logix.ram_r[1978] ;
 wire \logix.ram_r[1979] ;
 wire \logix.ram_r[197] ;
 wire \logix.ram_r[1980] ;
 wire \logix.ram_r[1981] ;
 wire \logix.ram_r[1982] ;
 wire \logix.ram_r[1983] ;
 wire \logix.ram_r[1984] ;
 wire \logix.ram_r[1985] ;
 wire \logix.ram_r[1986] ;
 wire \logix.ram_r[1987] ;
 wire \logix.ram_r[1988] ;
 wire \logix.ram_r[1989] ;
 wire \logix.ram_r[198] ;
 wire \logix.ram_r[1990] ;
 wire \logix.ram_r[1991] ;
 wire \logix.ram_r[1992] ;
 wire \logix.ram_r[1993] ;
 wire \logix.ram_r[1994] ;
 wire \logix.ram_r[1995] ;
 wire \logix.ram_r[1996] ;
 wire \logix.ram_r[1997] ;
 wire \logix.ram_r[1998] ;
 wire \logix.ram_r[1999] ;
 wire \logix.ram_r[199] ;
 wire \logix.ram_r[19] ;
 wire \logix.ram_r[1] ;
 wire \logix.ram_r[2000] ;
 wire \logix.ram_r[2001] ;
 wire \logix.ram_r[2002] ;
 wire \logix.ram_r[2003] ;
 wire \logix.ram_r[2004] ;
 wire \logix.ram_r[2005] ;
 wire \logix.ram_r[2006] ;
 wire \logix.ram_r[2007] ;
 wire \logix.ram_r[2008] ;
 wire \logix.ram_r[2009] ;
 wire \logix.ram_r[200] ;
 wire \logix.ram_r[2010] ;
 wire \logix.ram_r[2011] ;
 wire \logix.ram_r[2012] ;
 wire \logix.ram_r[2013] ;
 wire \logix.ram_r[2014] ;
 wire \logix.ram_r[2015] ;
 wire \logix.ram_r[2016] ;
 wire \logix.ram_r[2017] ;
 wire \logix.ram_r[2018] ;
 wire \logix.ram_r[2019] ;
 wire \logix.ram_r[201] ;
 wire \logix.ram_r[2020] ;
 wire \logix.ram_r[2021] ;
 wire \logix.ram_r[2022] ;
 wire \logix.ram_r[2023] ;
 wire \logix.ram_r[2024] ;
 wire \logix.ram_r[2025] ;
 wire \logix.ram_r[2026] ;
 wire \logix.ram_r[2027] ;
 wire \logix.ram_r[2028] ;
 wire \logix.ram_r[2029] ;
 wire \logix.ram_r[202] ;
 wire \logix.ram_r[2030] ;
 wire \logix.ram_r[2031] ;
 wire \logix.ram_r[2032] ;
 wire \logix.ram_r[2033] ;
 wire \logix.ram_r[2034] ;
 wire \logix.ram_r[2035] ;
 wire \logix.ram_r[2036] ;
 wire \logix.ram_r[2037] ;
 wire \logix.ram_r[2038] ;
 wire \logix.ram_r[2039] ;
 wire \logix.ram_r[203] ;
 wire \logix.ram_r[2040] ;
 wire \logix.ram_r[2041] ;
 wire \logix.ram_r[2042] ;
 wire \logix.ram_r[2043] ;
 wire \logix.ram_r[2044] ;
 wire \logix.ram_r[2045] ;
 wire \logix.ram_r[2046] ;
 wire \logix.ram_r[2047] ;
 wire \logix.ram_r[204] ;
 wire \logix.ram_r[205] ;
 wire \logix.ram_r[206] ;
 wire \logix.ram_r[207] ;
 wire \logix.ram_r[208] ;
 wire \logix.ram_r[209] ;
 wire \logix.ram_r[20] ;
 wire \logix.ram_r[210] ;
 wire \logix.ram_r[211] ;
 wire \logix.ram_r[212] ;
 wire \logix.ram_r[213] ;
 wire \logix.ram_r[214] ;
 wire \logix.ram_r[215] ;
 wire \logix.ram_r[216] ;
 wire \logix.ram_r[217] ;
 wire \logix.ram_r[218] ;
 wire \logix.ram_r[219] ;
 wire \logix.ram_r[21] ;
 wire \logix.ram_r[220] ;
 wire \logix.ram_r[221] ;
 wire \logix.ram_r[222] ;
 wire \logix.ram_r[223] ;
 wire \logix.ram_r[224] ;
 wire \logix.ram_r[225] ;
 wire \logix.ram_r[226] ;
 wire \logix.ram_r[227] ;
 wire \logix.ram_r[228] ;
 wire \logix.ram_r[229] ;
 wire \logix.ram_r[22] ;
 wire \logix.ram_r[230] ;
 wire \logix.ram_r[231] ;
 wire \logix.ram_r[232] ;
 wire \logix.ram_r[233] ;
 wire \logix.ram_r[234] ;
 wire \logix.ram_r[235] ;
 wire \logix.ram_r[236] ;
 wire \logix.ram_r[237] ;
 wire \logix.ram_r[238] ;
 wire \logix.ram_r[239] ;
 wire \logix.ram_r[23] ;
 wire \logix.ram_r[240] ;
 wire \logix.ram_r[241] ;
 wire \logix.ram_r[242] ;
 wire \logix.ram_r[243] ;
 wire \logix.ram_r[244] ;
 wire \logix.ram_r[245] ;
 wire \logix.ram_r[246] ;
 wire \logix.ram_r[247] ;
 wire \logix.ram_r[248] ;
 wire \logix.ram_r[249] ;
 wire \logix.ram_r[24] ;
 wire \logix.ram_r[250] ;
 wire \logix.ram_r[251] ;
 wire \logix.ram_r[252] ;
 wire \logix.ram_r[253] ;
 wire \logix.ram_r[254] ;
 wire \logix.ram_r[255] ;
 wire \logix.ram_r[256] ;
 wire \logix.ram_r[257] ;
 wire \logix.ram_r[258] ;
 wire \logix.ram_r[259] ;
 wire \logix.ram_r[25] ;
 wire \logix.ram_r[260] ;
 wire \logix.ram_r[261] ;
 wire \logix.ram_r[262] ;
 wire \logix.ram_r[263] ;
 wire \logix.ram_r[264] ;
 wire \logix.ram_r[265] ;
 wire \logix.ram_r[266] ;
 wire \logix.ram_r[267] ;
 wire \logix.ram_r[268] ;
 wire \logix.ram_r[269] ;
 wire \logix.ram_r[26] ;
 wire \logix.ram_r[270] ;
 wire \logix.ram_r[271] ;
 wire \logix.ram_r[272] ;
 wire \logix.ram_r[273] ;
 wire \logix.ram_r[274] ;
 wire \logix.ram_r[275] ;
 wire \logix.ram_r[276] ;
 wire \logix.ram_r[277] ;
 wire \logix.ram_r[278] ;
 wire \logix.ram_r[279] ;
 wire \logix.ram_r[27] ;
 wire \logix.ram_r[280] ;
 wire \logix.ram_r[281] ;
 wire \logix.ram_r[282] ;
 wire \logix.ram_r[283] ;
 wire \logix.ram_r[284] ;
 wire \logix.ram_r[285] ;
 wire \logix.ram_r[286] ;
 wire \logix.ram_r[287] ;
 wire \logix.ram_r[288] ;
 wire \logix.ram_r[289] ;
 wire \logix.ram_r[28] ;
 wire \logix.ram_r[290] ;
 wire \logix.ram_r[291] ;
 wire \logix.ram_r[292] ;
 wire \logix.ram_r[293] ;
 wire \logix.ram_r[294] ;
 wire \logix.ram_r[295] ;
 wire \logix.ram_r[296] ;
 wire \logix.ram_r[297] ;
 wire \logix.ram_r[298] ;
 wire \logix.ram_r[299] ;
 wire \logix.ram_r[29] ;
 wire \logix.ram_r[2] ;
 wire \logix.ram_r[300] ;
 wire \logix.ram_r[301] ;
 wire \logix.ram_r[302] ;
 wire \logix.ram_r[303] ;
 wire \logix.ram_r[304] ;
 wire \logix.ram_r[305] ;
 wire \logix.ram_r[306] ;
 wire \logix.ram_r[307] ;
 wire \logix.ram_r[308] ;
 wire \logix.ram_r[309] ;
 wire \logix.ram_r[30] ;
 wire \logix.ram_r[310] ;
 wire \logix.ram_r[311] ;
 wire \logix.ram_r[312] ;
 wire \logix.ram_r[313] ;
 wire \logix.ram_r[314] ;
 wire \logix.ram_r[315] ;
 wire \logix.ram_r[316] ;
 wire \logix.ram_r[317] ;
 wire \logix.ram_r[318] ;
 wire \logix.ram_r[319] ;
 wire \logix.ram_r[31] ;
 wire \logix.ram_r[320] ;
 wire \logix.ram_r[321] ;
 wire \logix.ram_r[322] ;
 wire \logix.ram_r[323] ;
 wire \logix.ram_r[324] ;
 wire \logix.ram_r[325] ;
 wire \logix.ram_r[326] ;
 wire \logix.ram_r[327] ;
 wire \logix.ram_r[328] ;
 wire \logix.ram_r[329] ;
 wire \logix.ram_r[32] ;
 wire \logix.ram_r[330] ;
 wire \logix.ram_r[331] ;
 wire \logix.ram_r[332] ;
 wire \logix.ram_r[333] ;
 wire \logix.ram_r[334] ;
 wire \logix.ram_r[335] ;
 wire \logix.ram_r[336] ;
 wire \logix.ram_r[337] ;
 wire \logix.ram_r[338] ;
 wire \logix.ram_r[339] ;
 wire \logix.ram_r[33] ;
 wire \logix.ram_r[340] ;
 wire \logix.ram_r[341] ;
 wire \logix.ram_r[342] ;
 wire \logix.ram_r[343] ;
 wire \logix.ram_r[344] ;
 wire \logix.ram_r[345] ;
 wire \logix.ram_r[346] ;
 wire \logix.ram_r[347] ;
 wire \logix.ram_r[348] ;
 wire \logix.ram_r[349] ;
 wire \logix.ram_r[34] ;
 wire \logix.ram_r[350] ;
 wire \logix.ram_r[351] ;
 wire \logix.ram_r[352] ;
 wire \logix.ram_r[353] ;
 wire \logix.ram_r[354] ;
 wire \logix.ram_r[355] ;
 wire \logix.ram_r[356] ;
 wire \logix.ram_r[357] ;
 wire \logix.ram_r[358] ;
 wire \logix.ram_r[359] ;
 wire \logix.ram_r[35] ;
 wire \logix.ram_r[360] ;
 wire \logix.ram_r[361] ;
 wire \logix.ram_r[362] ;
 wire \logix.ram_r[363] ;
 wire \logix.ram_r[364] ;
 wire \logix.ram_r[365] ;
 wire \logix.ram_r[366] ;
 wire \logix.ram_r[367] ;
 wire \logix.ram_r[368] ;
 wire \logix.ram_r[369] ;
 wire \logix.ram_r[36] ;
 wire \logix.ram_r[370] ;
 wire \logix.ram_r[371] ;
 wire \logix.ram_r[372] ;
 wire \logix.ram_r[373] ;
 wire \logix.ram_r[374] ;
 wire \logix.ram_r[375] ;
 wire \logix.ram_r[376] ;
 wire \logix.ram_r[377] ;
 wire \logix.ram_r[378] ;
 wire \logix.ram_r[379] ;
 wire \logix.ram_r[37] ;
 wire \logix.ram_r[380] ;
 wire \logix.ram_r[381] ;
 wire \logix.ram_r[382] ;
 wire \logix.ram_r[383] ;
 wire \logix.ram_r[384] ;
 wire \logix.ram_r[385] ;
 wire \logix.ram_r[386] ;
 wire \logix.ram_r[387] ;
 wire \logix.ram_r[388] ;
 wire \logix.ram_r[389] ;
 wire \logix.ram_r[38] ;
 wire \logix.ram_r[390] ;
 wire \logix.ram_r[391] ;
 wire \logix.ram_r[392] ;
 wire \logix.ram_r[393] ;
 wire \logix.ram_r[394] ;
 wire \logix.ram_r[395] ;
 wire \logix.ram_r[396] ;
 wire \logix.ram_r[397] ;
 wire \logix.ram_r[398] ;
 wire \logix.ram_r[399] ;
 wire \logix.ram_r[39] ;
 wire \logix.ram_r[3] ;
 wire \logix.ram_r[400] ;
 wire \logix.ram_r[401] ;
 wire \logix.ram_r[402] ;
 wire \logix.ram_r[403] ;
 wire \logix.ram_r[404] ;
 wire \logix.ram_r[405] ;
 wire \logix.ram_r[406] ;
 wire \logix.ram_r[407] ;
 wire \logix.ram_r[408] ;
 wire \logix.ram_r[409] ;
 wire \logix.ram_r[40] ;
 wire \logix.ram_r[410] ;
 wire \logix.ram_r[411] ;
 wire \logix.ram_r[412] ;
 wire \logix.ram_r[413] ;
 wire \logix.ram_r[414] ;
 wire \logix.ram_r[415] ;
 wire \logix.ram_r[416] ;
 wire \logix.ram_r[417] ;
 wire \logix.ram_r[418] ;
 wire \logix.ram_r[419] ;
 wire \logix.ram_r[41] ;
 wire \logix.ram_r[420] ;
 wire \logix.ram_r[421] ;
 wire \logix.ram_r[422] ;
 wire \logix.ram_r[423] ;
 wire \logix.ram_r[424] ;
 wire \logix.ram_r[425] ;
 wire \logix.ram_r[426] ;
 wire \logix.ram_r[427] ;
 wire \logix.ram_r[428] ;
 wire \logix.ram_r[429] ;
 wire \logix.ram_r[42] ;
 wire \logix.ram_r[430] ;
 wire \logix.ram_r[431] ;
 wire \logix.ram_r[432] ;
 wire \logix.ram_r[433] ;
 wire \logix.ram_r[434] ;
 wire \logix.ram_r[435] ;
 wire \logix.ram_r[436] ;
 wire \logix.ram_r[437] ;
 wire \logix.ram_r[438] ;
 wire \logix.ram_r[439] ;
 wire \logix.ram_r[43] ;
 wire \logix.ram_r[440] ;
 wire \logix.ram_r[441] ;
 wire \logix.ram_r[442] ;
 wire \logix.ram_r[443] ;
 wire \logix.ram_r[444] ;
 wire \logix.ram_r[445] ;
 wire \logix.ram_r[446] ;
 wire \logix.ram_r[447] ;
 wire \logix.ram_r[448] ;
 wire \logix.ram_r[449] ;
 wire \logix.ram_r[44] ;
 wire \logix.ram_r[450] ;
 wire \logix.ram_r[451] ;
 wire \logix.ram_r[452] ;
 wire \logix.ram_r[453] ;
 wire \logix.ram_r[454] ;
 wire \logix.ram_r[455] ;
 wire \logix.ram_r[456] ;
 wire \logix.ram_r[457] ;
 wire \logix.ram_r[458] ;
 wire \logix.ram_r[459] ;
 wire \logix.ram_r[45] ;
 wire \logix.ram_r[460] ;
 wire \logix.ram_r[461] ;
 wire \logix.ram_r[462] ;
 wire \logix.ram_r[463] ;
 wire \logix.ram_r[464] ;
 wire \logix.ram_r[465] ;
 wire \logix.ram_r[466] ;
 wire \logix.ram_r[467] ;
 wire \logix.ram_r[468] ;
 wire \logix.ram_r[469] ;
 wire \logix.ram_r[46] ;
 wire \logix.ram_r[470] ;
 wire \logix.ram_r[471] ;
 wire \logix.ram_r[472] ;
 wire \logix.ram_r[473] ;
 wire \logix.ram_r[474] ;
 wire \logix.ram_r[475] ;
 wire \logix.ram_r[476] ;
 wire \logix.ram_r[477] ;
 wire \logix.ram_r[478] ;
 wire \logix.ram_r[479] ;
 wire \logix.ram_r[47] ;
 wire \logix.ram_r[480] ;
 wire \logix.ram_r[481] ;
 wire \logix.ram_r[482] ;
 wire \logix.ram_r[483] ;
 wire \logix.ram_r[484] ;
 wire \logix.ram_r[485] ;
 wire \logix.ram_r[486] ;
 wire \logix.ram_r[487] ;
 wire \logix.ram_r[488] ;
 wire \logix.ram_r[489] ;
 wire \logix.ram_r[48] ;
 wire \logix.ram_r[490] ;
 wire \logix.ram_r[491] ;
 wire \logix.ram_r[492] ;
 wire \logix.ram_r[493] ;
 wire \logix.ram_r[494] ;
 wire \logix.ram_r[495] ;
 wire \logix.ram_r[496] ;
 wire \logix.ram_r[497] ;
 wire \logix.ram_r[498] ;
 wire \logix.ram_r[499] ;
 wire \logix.ram_r[49] ;
 wire \logix.ram_r[4] ;
 wire \logix.ram_r[500] ;
 wire \logix.ram_r[501] ;
 wire \logix.ram_r[502] ;
 wire \logix.ram_r[503] ;
 wire \logix.ram_r[504] ;
 wire \logix.ram_r[505] ;
 wire \logix.ram_r[506] ;
 wire \logix.ram_r[507] ;
 wire \logix.ram_r[508] ;
 wire \logix.ram_r[509] ;
 wire \logix.ram_r[50] ;
 wire \logix.ram_r[510] ;
 wire \logix.ram_r[511] ;
 wire \logix.ram_r[512] ;
 wire \logix.ram_r[513] ;
 wire \logix.ram_r[514] ;
 wire \logix.ram_r[515] ;
 wire \logix.ram_r[516] ;
 wire \logix.ram_r[517] ;
 wire \logix.ram_r[518] ;
 wire \logix.ram_r[519] ;
 wire \logix.ram_r[51] ;
 wire \logix.ram_r[520] ;
 wire \logix.ram_r[521] ;
 wire \logix.ram_r[522] ;
 wire \logix.ram_r[523] ;
 wire \logix.ram_r[524] ;
 wire \logix.ram_r[525] ;
 wire \logix.ram_r[526] ;
 wire \logix.ram_r[527] ;
 wire \logix.ram_r[528] ;
 wire \logix.ram_r[529] ;
 wire \logix.ram_r[52] ;
 wire \logix.ram_r[530] ;
 wire \logix.ram_r[531] ;
 wire \logix.ram_r[532] ;
 wire \logix.ram_r[533] ;
 wire \logix.ram_r[534] ;
 wire \logix.ram_r[535] ;
 wire \logix.ram_r[536] ;
 wire \logix.ram_r[537] ;
 wire \logix.ram_r[538] ;
 wire \logix.ram_r[539] ;
 wire \logix.ram_r[53] ;
 wire \logix.ram_r[540] ;
 wire \logix.ram_r[541] ;
 wire \logix.ram_r[542] ;
 wire \logix.ram_r[543] ;
 wire \logix.ram_r[544] ;
 wire \logix.ram_r[545] ;
 wire \logix.ram_r[546] ;
 wire \logix.ram_r[547] ;
 wire \logix.ram_r[548] ;
 wire \logix.ram_r[549] ;
 wire \logix.ram_r[54] ;
 wire \logix.ram_r[550] ;
 wire \logix.ram_r[551] ;
 wire \logix.ram_r[552] ;
 wire \logix.ram_r[553] ;
 wire \logix.ram_r[554] ;
 wire \logix.ram_r[555] ;
 wire \logix.ram_r[556] ;
 wire \logix.ram_r[557] ;
 wire \logix.ram_r[558] ;
 wire \logix.ram_r[559] ;
 wire \logix.ram_r[55] ;
 wire \logix.ram_r[560] ;
 wire \logix.ram_r[561] ;
 wire \logix.ram_r[562] ;
 wire \logix.ram_r[563] ;
 wire \logix.ram_r[564] ;
 wire \logix.ram_r[565] ;
 wire \logix.ram_r[566] ;
 wire \logix.ram_r[567] ;
 wire \logix.ram_r[568] ;
 wire \logix.ram_r[569] ;
 wire \logix.ram_r[56] ;
 wire \logix.ram_r[570] ;
 wire \logix.ram_r[571] ;
 wire \logix.ram_r[572] ;
 wire \logix.ram_r[573] ;
 wire \logix.ram_r[574] ;
 wire \logix.ram_r[575] ;
 wire \logix.ram_r[576] ;
 wire \logix.ram_r[577] ;
 wire \logix.ram_r[578] ;
 wire \logix.ram_r[579] ;
 wire \logix.ram_r[57] ;
 wire \logix.ram_r[580] ;
 wire \logix.ram_r[581] ;
 wire \logix.ram_r[582] ;
 wire \logix.ram_r[583] ;
 wire \logix.ram_r[584] ;
 wire \logix.ram_r[585] ;
 wire \logix.ram_r[586] ;
 wire \logix.ram_r[587] ;
 wire \logix.ram_r[588] ;
 wire \logix.ram_r[589] ;
 wire \logix.ram_r[58] ;
 wire \logix.ram_r[590] ;
 wire \logix.ram_r[591] ;
 wire \logix.ram_r[592] ;
 wire \logix.ram_r[593] ;
 wire \logix.ram_r[594] ;
 wire \logix.ram_r[595] ;
 wire \logix.ram_r[596] ;
 wire \logix.ram_r[597] ;
 wire \logix.ram_r[598] ;
 wire \logix.ram_r[599] ;
 wire \logix.ram_r[59] ;
 wire \logix.ram_r[5] ;
 wire \logix.ram_r[600] ;
 wire \logix.ram_r[601] ;
 wire \logix.ram_r[602] ;
 wire \logix.ram_r[603] ;
 wire \logix.ram_r[604] ;
 wire \logix.ram_r[605] ;
 wire \logix.ram_r[606] ;
 wire \logix.ram_r[607] ;
 wire \logix.ram_r[608] ;
 wire \logix.ram_r[609] ;
 wire \logix.ram_r[60] ;
 wire \logix.ram_r[610] ;
 wire \logix.ram_r[611] ;
 wire \logix.ram_r[612] ;
 wire \logix.ram_r[613] ;
 wire \logix.ram_r[614] ;
 wire \logix.ram_r[615] ;
 wire \logix.ram_r[616] ;
 wire \logix.ram_r[617] ;
 wire \logix.ram_r[618] ;
 wire \logix.ram_r[619] ;
 wire \logix.ram_r[61] ;
 wire \logix.ram_r[620] ;
 wire \logix.ram_r[621] ;
 wire \logix.ram_r[622] ;
 wire \logix.ram_r[623] ;
 wire \logix.ram_r[624] ;
 wire \logix.ram_r[625] ;
 wire \logix.ram_r[626] ;
 wire \logix.ram_r[627] ;
 wire \logix.ram_r[628] ;
 wire \logix.ram_r[629] ;
 wire \logix.ram_r[62] ;
 wire \logix.ram_r[630] ;
 wire \logix.ram_r[631] ;
 wire \logix.ram_r[632] ;
 wire \logix.ram_r[633] ;
 wire \logix.ram_r[634] ;
 wire \logix.ram_r[635] ;
 wire \logix.ram_r[636] ;
 wire \logix.ram_r[637] ;
 wire \logix.ram_r[638] ;
 wire \logix.ram_r[639] ;
 wire \logix.ram_r[63] ;
 wire \logix.ram_r[640] ;
 wire \logix.ram_r[641] ;
 wire \logix.ram_r[642] ;
 wire \logix.ram_r[643] ;
 wire \logix.ram_r[644] ;
 wire \logix.ram_r[645] ;
 wire \logix.ram_r[646] ;
 wire \logix.ram_r[647] ;
 wire \logix.ram_r[648] ;
 wire \logix.ram_r[649] ;
 wire \logix.ram_r[64] ;
 wire \logix.ram_r[650] ;
 wire \logix.ram_r[651] ;
 wire \logix.ram_r[652] ;
 wire \logix.ram_r[653] ;
 wire \logix.ram_r[654] ;
 wire \logix.ram_r[655] ;
 wire \logix.ram_r[656] ;
 wire \logix.ram_r[657] ;
 wire \logix.ram_r[658] ;
 wire \logix.ram_r[659] ;
 wire \logix.ram_r[65] ;
 wire \logix.ram_r[660] ;
 wire \logix.ram_r[661] ;
 wire \logix.ram_r[662] ;
 wire \logix.ram_r[663] ;
 wire \logix.ram_r[664] ;
 wire \logix.ram_r[665] ;
 wire \logix.ram_r[666] ;
 wire \logix.ram_r[667] ;
 wire \logix.ram_r[668] ;
 wire \logix.ram_r[669] ;
 wire \logix.ram_r[66] ;
 wire \logix.ram_r[670] ;
 wire \logix.ram_r[671] ;
 wire \logix.ram_r[672] ;
 wire \logix.ram_r[673] ;
 wire \logix.ram_r[674] ;
 wire \logix.ram_r[675] ;
 wire \logix.ram_r[676] ;
 wire \logix.ram_r[677] ;
 wire \logix.ram_r[678] ;
 wire \logix.ram_r[679] ;
 wire \logix.ram_r[67] ;
 wire \logix.ram_r[680] ;
 wire \logix.ram_r[681] ;
 wire \logix.ram_r[682] ;
 wire \logix.ram_r[683] ;
 wire \logix.ram_r[684] ;
 wire \logix.ram_r[685] ;
 wire \logix.ram_r[686] ;
 wire \logix.ram_r[687] ;
 wire \logix.ram_r[688] ;
 wire \logix.ram_r[689] ;
 wire \logix.ram_r[68] ;
 wire \logix.ram_r[690] ;
 wire \logix.ram_r[691] ;
 wire \logix.ram_r[692] ;
 wire \logix.ram_r[693] ;
 wire \logix.ram_r[694] ;
 wire \logix.ram_r[695] ;
 wire \logix.ram_r[696] ;
 wire \logix.ram_r[697] ;
 wire \logix.ram_r[698] ;
 wire \logix.ram_r[699] ;
 wire \logix.ram_r[69] ;
 wire \logix.ram_r[6] ;
 wire \logix.ram_r[700] ;
 wire \logix.ram_r[701] ;
 wire \logix.ram_r[702] ;
 wire \logix.ram_r[703] ;
 wire \logix.ram_r[704] ;
 wire \logix.ram_r[705] ;
 wire \logix.ram_r[706] ;
 wire \logix.ram_r[707] ;
 wire \logix.ram_r[708] ;
 wire \logix.ram_r[709] ;
 wire \logix.ram_r[70] ;
 wire \logix.ram_r[710] ;
 wire \logix.ram_r[711] ;
 wire \logix.ram_r[712] ;
 wire \logix.ram_r[713] ;
 wire \logix.ram_r[714] ;
 wire \logix.ram_r[715] ;
 wire \logix.ram_r[716] ;
 wire \logix.ram_r[717] ;
 wire \logix.ram_r[718] ;
 wire \logix.ram_r[719] ;
 wire \logix.ram_r[71] ;
 wire \logix.ram_r[720] ;
 wire \logix.ram_r[721] ;
 wire \logix.ram_r[722] ;
 wire \logix.ram_r[723] ;
 wire \logix.ram_r[724] ;
 wire \logix.ram_r[725] ;
 wire \logix.ram_r[726] ;
 wire \logix.ram_r[727] ;
 wire \logix.ram_r[728] ;
 wire \logix.ram_r[729] ;
 wire \logix.ram_r[72] ;
 wire \logix.ram_r[730] ;
 wire \logix.ram_r[731] ;
 wire \logix.ram_r[732] ;
 wire \logix.ram_r[733] ;
 wire \logix.ram_r[734] ;
 wire \logix.ram_r[735] ;
 wire \logix.ram_r[736] ;
 wire \logix.ram_r[737] ;
 wire \logix.ram_r[738] ;
 wire \logix.ram_r[739] ;
 wire \logix.ram_r[73] ;
 wire \logix.ram_r[740] ;
 wire \logix.ram_r[741] ;
 wire \logix.ram_r[742] ;
 wire \logix.ram_r[743] ;
 wire \logix.ram_r[744] ;
 wire \logix.ram_r[745] ;
 wire \logix.ram_r[746] ;
 wire \logix.ram_r[747] ;
 wire \logix.ram_r[748] ;
 wire \logix.ram_r[749] ;
 wire \logix.ram_r[74] ;
 wire \logix.ram_r[750] ;
 wire \logix.ram_r[751] ;
 wire \logix.ram_r[752] ;
 wire \logix.ram_r[753] ;
 wire \logix.ram_r[754] ;
 wire \logix.ram_r[755] ;
 wire \logix.ram_r[756] ;
 wire \logix.ram_r[757] ;
 wire \logix.ram_r[758] ;
 wire \logix.ram_r[759] ;
 wire \logix.ram_r[75] ;
 wire \logix.ram_r[760] ;
 wire \logix.ram_r[761] ;
 wire \logix.ram_r[762] ;
 wire \logix.ram_r[763] ;
 wire \logix.ram_r[764] ;
 wire \logix.ram_r[765] ;
 wire \logix.ram_r[766] ;
 wire \logix.ram_r[767] ;
 wire \logix.ram_r[768] ;
 wire \logix.ram_r[769] ;
 wire \logix.ram_r[76] ;
 wire \logix.ram_r[770] ;
 wire \logix.ram_r[771] ;
 wire \logix.ram_r[772] ;
 wire \logix.ram_r[773] ;
 wire \logix.ram_r[774] ;
 wire \logix.ram_r[775] ;
 wire \logix.ram_r[776] ;
 wire \logix.ram_r[777] ;
 wire \logix.ram_r[778] ;
 wire \logix.ram_r[779] ;
 wire \logix.ram_r[77] ;
 wire \logix.ram_r[780] ;
 wire \logix.ram_r[781] ;
 wire \logix.ram_r[782] ;
 wire \logix.ram_r[783] ;
 wire \logix.ram_r[784] ;
 wire \logix.ram_r[785] ;
 wire \logix.ram_r[786] ;
 wire \logix.ram_r[787] ;
 wire \logix.ram_r[788] ;
 wire \logix.ram_r[789] ;
 wire \logix.ram_r[78] ;
 wire \logix.ram_r[790] ;
 wire \logix.ram_r[791] ;
 wire \logix.ram_r[792] ;
 wire \logix.ram_r[793] ;
 wire \logix.ram_r[794] ;
 wire \logix.ram_r[795] ;
 wire \logix.ram_r[796] ;
 wire \logix.ram_r[797] ;
 wire \logix.ram_r[798] ;
 wire \logix.ram_r[799] ;
 wire \logix.ram_r[79] ;
 wire \logix.ram_r[7] ;
 wire \logix.ram_r[800] ;
 wire \logix.ram_r[801] ;
 wire \logix.ram_r[802] ;
 wire \logix.ram_r[803] ;
 wire \logix.ram_r[804] ;
 wire \logix.ram_r[805] ;
 wire \logix.ram_r[806] ;
 wire \logix.ram_r[807] ;
 wire \logix.ram_r[808] ;
 wire \logix.ram_r[809] ;
 wire \logix.ram_r[80] ;
 wire \logix.ram_r[810] ;
 wire \logix.ram_r[811] ;
 wire \logix.ram_r[812] ;
 wire \logix.ram_r[813] ;
 wire \logix.ram_r[814] ;
 wire \logix.ram_r[815] ;
 wire \logix.ram_r[816] ;
 wire \logix.ram_r[817] ;
 wire \logix.ram_r[818] ;
 wire \logix.ram_r[819] ;
 wire \logix.ram_r[81] ;
 wire \logix.ram_r[820] ;
 wire \logix.ram_r[821] ;
 wire \logix.ram_r[822] ;
 wire \logix.ram_r[823] ;
 wire \logix.ram_r[824] ;
 wire \logix.ram_r[825] ;
 wire \logix.ram_r[826] ;
 wire \logix.ram_r[827] ;
 wire \logix.ram_r[828] ;
 wire \logix.ram_r[829] ;
 wire \logix.ram_r[82] ;
 wire \logix.ram_r[830] ;
 wire \logix.ram_r[831] ;
 wire \logix.ram_r[832] ;
 wire \logix.ram_r[833] ;
 wire \logix.ram_r[834] ;
 wire \logix.ram_r[835] ;
 wire \logix.ram_r[836] ;
 wire \logix.ram_r[837] ;
 wire \logix.ram_r[838] ;
 wire \logix.ram_r[839] ;
 wire \logix.ram_r[83] ;
 wire \logix.ram_r[840] ;
 wire \logix.ram_r[841] ;
 wire \logix.ram_r[842] ;
 wire \logix.ram_r[843] ;
 wire \logix.ram_r[844] ;
 wire \logix.ram_r[845] ;
 wire \logix.ram_r[846] ;
 wire \logix.ram_r[847] ;
 wire \logix.ram_r[848] ;
 wire \logix.ram_r[849] ;
 wire \logix.ram_r[84] ;
 wire \logix.ram_r[850] ;
 wire \logix.ram_r[851] ;
 wire \logix.ram_r[852] ;
 wire \logix.ram_r[853] ;
 wire \logix.ram_r[854] ;
 wire \logix.ram_r[855] ;
 wire \logix.ram_r[856] ;
 wire \logix.ram_r[857] ;
 wire \logix.ram_r[858] ;
 wire \logix.ram_r[859] ;
 wire \logix.ram_r[85] ;
 wire \logix.ram_r[860] ;
 wire \logix.ram_r[861] ;
 wire \logix.ram_r[862] ;
 wire \logix.ram_r[863] ;
 wire \logix.ram_r[864] ;
 wire \logix.ram_r[865] ;
 wire \logix.ram_r[866] ;
 wire \logix.ram_r[867] ;
 wire \logix.ram_r[868] ;
 wire \logix.ram_r[869] ;
 wire \logix.ram_r[86] ;
 wire \logix.ram_r[870] ;
 wire \logix.ram_r[871] ;
 wire \logix.ram_r[872] ;
 wire \logix.ram_r[873] ;
 wire \logix.ram_r[874] ;
 wire \logix.ram_r[875] ;
 wire \logix.ram_r[876] ;
 wire \logix.ram_r[877] ;
 wire \logix.ram_r[878] ;
 wire \logix.ram_r[879] ;
 wire \logix.ram_r[87] ;
 wire \logix.ram_r[880] ;
 wire \logix.ram_r[881] ;
 wire \logix.ram_r[882] ;
 wire \logix.ram_r[883] ;
 wire \logix.ram_r[884] ;
 wire \logix.ram_r[885] ;
 wire \logix.ram_r[886] ;
 wire \logix.ram_r[887] ;
 wire \logix.ram_r[888] ;
 wire \logix.ram_r[889] ;
 wire \logix.ram_r[88] ;
 wire \logix.ram_r[890] ;
 wire \logix.ram_r[891] ;
 wire \logix.ram_r[892] ;
 wire \logix.ram_r[893] ;
 wire \logix.ram_r[894] ;
 wire \logix.ram_r[895] ;
 wire \logix.ram_r[896] ;
 wire \logix.ram_r[897] ;
 wire \logix.ram_r[898] ;
 wire \logix.ram_r[899] ;
 wire \logix.ram_r[89] ;
 wire \logix.ram_r[8] ;
 wire \logix.ram_r[900] ;
 wire \logix.ram_r[901] ;
 wire \logix.ram_r[902] ;
 wire \logix.ram_r[903] ;
 wire \logix.ram_r[904] ;
 wire \logix.ram_r[905] ;
 wire \logix.ram_r[906] ;
 wire \logix.ram_r[907] ;
 wire \logix.ram_r[908] ;
 wire \logix.ram_r[909] ;
 wire \logix.ram_r[90] ;
 wire \logix.ram_r[910] ;
 wire \logix.ram_r[911] ;
 wire \logix.ram_r[912] ;
 wire \logix.ram_r[913] ;
 wire \logix.ram_r[914] ;
 wire \logix.ram_r[915] ;
 wire \logix.ram_r[916] ;
 wire \logix.ram_r[917] ;
 wire \logix.ram_r[918] ;
 wire \logix.ram_r[919] ;
 wire \logix.ram_r[91] ;
 wire \logix.ram_r[920] ;
 wire \logix.ram_r[921] ;
 wire \logix.ram_r[922] ;
 wire \logix.ram_r[923] ;
 wire \logix.ram_r[924] ;
 wire \logix.ram_r[925] ;
 wire \logix.ram_r[926] ;
 wire \logix.ram_r[927] ;
 wire \logix.ram_r[928] ;
 wire \logix.ram_r[929] ;
 wire \logix.ram_r[92] ;
 wire \logix.ram_r[930] ;
 wire \logix.ram_r[931] ;
 wire \logix.ram_r[932] ;
 wire \logix.ram_r[933] ;
 wire \logix.ram_r[934] ;
 wire \logix.ram_r[935] ;
 wire \logix.ram_r[936] ;
 wire \logix.ram_r[937] ;
 wire \logix.ram_r[938] ;
 wire \logix.ram_r[939] ;
 wire \logix.ram_r[93] ;
 wire \logix.ram_r[940] ;
 wire \logix.ram_r[941] ;
 wire \logix.ram_r[942] ;
 wire \logix.ram_r[943] ;
 wire \logix.ram_r[944] ;
 wire \logix.ram_r[945] ;
 wire \logix.ram_r[946] ;
 wire \logix.ram_r[947] ;
 wire \logix.ram_r[948] ;
 wire \logix.ram_r[949] ;
 wire \logix.ram_r[94] ;
 wire \logix.ram_r[950] ;
 wire \logix.ram_r[951] ;
 wire \logix.ram_r[952] ;
 wire \logix.ram_r[953] ;
 wire \logix.ram_r[954] ;
 wire \logix.ram_r[955] ;
 wire \logix.ram_r[956] ;
 wire \logix.ram_r[957] ;
 wire \logix.ram_r[958] ;
 wire \logix.ram_r[959] ;
 wire \logix.ram_r[95] ;
 wire \logix.ram_r[960] ;
 wire \logix.ram_r[961] ;
 wire \logix.ram_r[962] ;
 wire \logix.ram_r[963] ;
 wire \logix.ram_r[964] ;
 wire \logix.ram_r[965] ;
 wire \logix.ram_r[966] ;
 wire \logix.ram_r[967] ;
 wire \logix.ram_r[968] ;
 wire \logix.ram_r[969] ;
 wire \logix.ram_r[96] ;
 wire \logix.ram_r[970] ;
 wire \logix.ram_r[971] ;
 wire \logix.ram_r[972] ;
 wire \logix.ram_r[973] ;
 wire \logix.ram_r[974] ;
 wire \logix.ram_r[975] ;
 wire \logix.ram_r[976] ;
 wire \logix.ram_r[977] ;
 wire \logix.ram_r[978] ;
 wire \logix.ram_r[979] ;
 wire \logix.ram_r[97] ;
 wire \logix.ram_r[980] ;
 wire \logix.ram_r[981] ;
 wire \logix.ram_r[982] ;
 wire \logix.ram_r[983] ;
 wire \logix.ram_r[984] ;
 wire \logix.ram_r[985] ;
 wire \logix.ram_r[986] ;
 wire \logix.ram_r[987] ;
 wire \logix.ram_r[988] ;
 wire \logix.ram_r[989] ;
 wire \logix.ram_r[98] ;
 wire \logix.ram_r[990] ;
 wire \logix.ram_r[991] ;
 wire \logix.ram_r[992] ;
 wire \logix.ram_r[993] ;
 wire \logix.ram_r[994] ;
 wire \logix.ram_r[995] ;
 wire \logix.ram_r[996] ;
 wire \logix.ram_r[997] ;
 wire \logix.ram_r[998] ;
 wire \logix.ram_r[999] ;
 wire \logix.ram_r[99] ;
 wire \logix.ram_r[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sg13g2_buf_2 _5995_ (.A(uio_in[0]),
    .X(_2063_));
 sg13g2_buf_2 _5996_ (.A(_2063_),
    .X(_2064_));
 sg13g2_buf_1 _5997_ (.A(_2064_),
    .X(_2065_));
 sg13g2_buf_1 _5998_ (.A(net413),
    .X(_2066_));
 sg13g2_mux2_1 _5999_ (.A0(\logix.ram_r[0] ),
    .A1(net10),
    .S(net412),
    .X(_0007_));
 sg13g2_mux2_1 _6000_ (.A0(\logix.ram_r[1000] ),
    .A1(\logix.ram_r[999] ),
    .S(net412),
    .X(_0008_));
 sg13g2_mux2_1 _6001_ (.A0(\logix.ram_r[1001] ),
    .A1(\logix.ram_r[1000] ),
    .S(net412),
    .X(_0009_));
 sg13g2_mux2_1 _6002_ (.A0(\logix.ram_r[1002] ),
    .A1(\logix.ram_r[1001] ),
    .S(net412),
    .X(_0010_));
 sg13g2_mux2_1 _6003_ (.A0(\logix.ram_r[1003] ),
    .A1(\logix.ram_r[1002] ),
    .S(net412),
    .X(_0011_));
 sg13g2_mux2_1 _6004_ (.A0(\logix.ram_r[1004] ),
    .A1(\logix.ram_r[1003] ),
    .S(net412),
    .X(_0012_));
 sg13g2_mux2_1 _6005_ (.A0(\logix.ram_r[1005] ),
    .A1(\logix.ram_r[1004] ),
    .S(net412),
    .X(_0013_));
 sg13g2_mux2_1 _6006_ (.A0(\logix.ram_r[1006] ),
    .A1(\logix.ram_r[1005] ),
    .S(_2066_),
    .X(_0014_));
 sg13g2_mux2_1 _6007_ (.A0(\logix.ram_r[1007] ),
    .A1(\logix.ram_r[1006] ),
    .S(net412),
    .X(_0015_));
 sg13g2_mux2_1 _6008_ (.A0(\logix.ram_r[1008] ),
    .A1(\logix.ram_r[1007] ),
    .S(_2066_),
    .X(_0016_));
 sg13g2_buf_1 _6009_ (.A(net413),
    .X(_2067_));
 sg13g2_mux2_1 _6010_ (.A0(\logix.ram_r[1009] ),
    .A1(\logix.ram_r[1008] ),
    .S(net411),
    .X(_0017_));
 sg13g2_mux2_1 _6011_ (.A0(\logix.ram_r[100] ),
    .A1(\logix.ram_r[99] ),
    .S(_2067_),
    .X(_0018_));
 sg13g2_mux2_1 _6012_ (.A0(\logix.ram_r[1010] ),
    .A1(\logix.ram_r[1009] ),
    .S(net411),
    .X(_0019_));
 sg13g2_mux2_1 _6013_ (.A0(\logix.ram_r[1011] ),
    .A1(\logix.ram_r[1010] ),
    .S(net411),
    .X(_0020_));
 sg13g2_mux2_1 _6014_ (.A0(\logix.ram_r[1012] ),
    .A1(\logix.ram_r[1011] ),
    .S(net411),
    .X(_0021_));
 sg13g2_mux2_1 _6015_ (.A0(\logix.ram_r[1013] ),
    .A1(\logix.ram_r[1012] ),
    .S(_2067_),
    .X(_0022_));
 sg13g2_mux2_1 _6016_ (.A0(\logix.ram_r[1014] ),
    .A1(\logix.ram_r[1013] ),
    .S(net411),
    .X(_0023_));
 sg13g2_mux2_1 _6017_ (.A0(\logix.ram_r[1015] ),
    .A1(\logix.ram_r[1014] ),
    .S(net411),
    .X(_0024_));
 sg13g2_mux2_1 _6018_ (.A0(\logix.ram_r[1016] ),
    .A1(\logix.ram_r[1015] ),
    .S(net411),
    .X(_0025_));
 sg13g2_mux2_1 _6019_ (.A0(\logix.ram_r[1017] ),
    .A1(\logix.ram_r[1016] ),
    .S(net411),
    .X(_0026_));
 sg13g2_buf_1 _6020_ (.A(net413),
    .X(_2068_));
 sg13g2_mux2_1 _6021_ (.A0(\logix.ram_r[1018] ),
    .A1(\logix.ram_r[1017] ),
    .S(net410),
    .X(_0027_));
 sg13g2_mux2_1 _6022_ (.A0(\logix.ram_r[1019] ),
    .A1(\logix.ram_r[1018] ),
    .S(net410),
    .X(_0028_));
 sg13g2_mux2_1 _6023_ (.A0(\logix.ram_r[101] ),
    .A1(\logix.ram_r[100] ),
    .S(net410),
    .X(_0029_));
 sg13g2_mux2_1 _6024_ (.A0(\logix.ram_r[1020] ),
    .A1(\logix.ram_r[1019] ),
    .S(net410),
    .X(_0030_));
 sg13g2_mux2_1 _6025_ (.A0(\logix.ram_r[1021] ),
    .A1(\logix.ram_r[1020] ),
    .S(net410),
    .X(_0031_));
 sg13g2_mux2_1 _6026_ (.A0(\logix.ram_r[1022] ),
    .A1(\logix.ram_r[1021] ),
    .S(net410),
    .X(_0032_));
 sg13g2_mux2_1 _6027_ (.A0(\logix.ram_r[1023] ),
    .A1(\logix.ram_r[1022] ),
    .S(net410),
    .X(_0033_));
 sg13g2_mux2_1 _6028_ (.A0(\logix.ram_r[1024] ),
    .A1(\logix.ram_r[1023] ),
    .S(net410),
    .X(_0034_));
 sg13g2_mux2_1 _6029_ (.A0(\logix.ram_r[1025] ),
    .A1(\logix.ram_r[1024] ),
    .S(_2068_),
    .X(_0035_));
 sg13g2_mux2_1 _6030_ (.A0(\logix.ram_r[1026] ),
    .A1(\logix.ram_r[1025] ),
    .S(_2068_),
    .X(_0036_));
 sg13g2_buf_1 _6031_ (.A(_2065_),
    .X(_2069_));
 sg13g2_mux2_1 _6032_ (.A0(\logix.ram_r[1027] ),
    .A1(\logix.ram_r[1026] ),
    .S(net409),
    .X(_0037_));
 sg13g2_mux2_1 _6033_ (.A0(\logix.ram_r[1028] ),
    .A1(\logix.ram_r[1027] ),
    .S(net409),
    .X(_0038_));
 sg13g2_mux2_1 _6034_ (.A0(\logix.ram_r[1029] ),
    .A1(\logix.ram_r[1028] ),
    .S(net409),
    .X(_0039_));
 sg13g2_mux2_1 _6035_ (.A0(\logix.ram_r[102] ),
    .A1(\logix.ram_r[101] ),
    .S(_2069_),
    .X(_0040_));
 sg13g2_mux2_1 _6036_ (.A0(\logix.ram_r[1030] ),
    .A1(\logix.ram_r[1029] ),
    .S(_2069_),
    .X(_0041_));
 sg13g2_mux2_1 _6037_ (.A0(\logix.ram_r[1031] ),
    .A1(\logix.ram_r[1030] ),
    .S(net409),
    .X(_0042_));
 sg13g2_mux2_1 _6038_ (.A0(\logix.ram_r[1032] ),
    .A1(\logix.ram_r[1031] ),
    .S(net409),
    .X(_0043_));
 sg13g2_mux2_1 _6039_ (.A0(\logix.ram_r[1033] ),
    .A1(\logix.ram_r[1032] ),
    .S(net409),
    .X(_0044_));
 sg13g2_mux2_1 _6040_ (.A0(\logix.ram_r[1034] ),
    .A1(\logix.ram_r[1033] ),
    .S(net409),
    .X(_0045_));
 sg13g2_mux2_1 _6041_ (.A0(\logix.ram_r[1035] ),
    .A1(\logix.ram_r[1034] ),
    .S(net409),
    .X(_0046_));
 sg13g2_buf_2 _6042_ (.A(_2064_),
    .X(_2070_));
 sg13g2_buf_1 _6043_ (.A(_2070_),
    .X(_2071_));
 sg13g2_buf_2 _6044_ (.A(_2071_),
    .X(_2072_));
 sg13g2_mux2_1 _6045_ (.A0(\logix.ram_r[1036] ),
    .A1(\logix.ram_r[1035] ),
    .S(net221),
    .X(_0047_));
 sg13g2_mux2_1 _6046_ (.A0(\logix.ram_r[1037] ),
    .A1(\logix.ram_r[1036] ),
    .S(net221),
    .X(_0048_));
 sg13g2_mux2_1 _6047_ (.A0(\logix.ram_r[1038] ),
    .A1(\logix.ram_r[1037] ),
    .S(net221),
    .X(_0049_));
 sg13g2_mux2_1 _6048_ (.A0(\logix.ram_r[1039] ),
    .A1(\logix.ram_r[1038] ),
    .S(net221),
    .X(_0050_));
 sg13g2_mux2_1 _6049_ (.A0(\logix.ram_r[103] ),
    .A1(\logix.ram_r[102] ),
    .S(net221),
    .X(_0051_));
 sg13g2_mux2_1 _6050_ (.A0(\logix.ram_r[1040] ),
    .A1(\logix.ram_r[1039] ),
    .S(_2072_),
    .X(_0052_));
 sg13g2_mux2_1 _6051_ (.A0(\logix.ram_r[1041] ),
    .A1(\logix.ram_r[1040] ),
    .S(_2072_),
    .X(_0053_));
 sg13g2_mux2_1 _6052_ (.A0(\logix.ram_r[1042] ),
    .A1(\logix.ram_r[1041] ),
    .S(net221),
    .X(_0054_));
 sg13g2_mux2_1 _6053_ (.A0(\logix.ram_r[1043] ),
    .A1(\logix.ram_r[1042] ),
    .S(net221),
    .X(_0055_));
 sg13g2_mux2_1 _6054_ (.A0(\logix.ram_r[1044] ),
    .A1(\logix.ram_r[1043] ),
    .S(net221),
    .X(_0056_));
 sg13g2_buf_2 _6055_ (.A(_2071_),
    .X(_2073_));
 sg13g2_mux2_1 _6056_ (.A0(\logix.ram_r[1045] ),
    .A1(\logix.ram_r[1044] ),
    .S(net220),
    .X(_0057_));
 sg13g2_mux2_1 _6057_ (.A0(\logix.ram_r[1046] ),
    .A1(\logix.ram_r[1045] ),
    .S(net220),
    .X(_0058_));
 sg13g2_mux2_1 _6058_ (.A0(\logix.ram_r[1047] ),
    .A1(\logix.ram_r[1046] ),
    .S(net220),
    .X(_0059_));
 sg13g2_mux2_1 _6059_ (.A0(\logix.ram_r[1048] ),
    .A1(\logix.ram_r[1047] ),
    .S(net220),
    .X(_0060_));
 sg13g2_mux2_1 _6060_ (.A0(\logix.ram_r[1049] ),
    .A1(\logix.ram_r[1048] ),
    .S(net220),
    .X(_0061_));
 sg13g2_mux2_1 _6061_ (.A0(\logix.ram_r[104] ),
    .A1(\logix.ram_r[103] ),
    .S(net220),
    .X(_0062_));
 sg13g2_mux2_1 _6062_ (.A0(\logix.ram_r[1050] ),
    .A1(\logix.ram_r[1049] ),
    .S(net220),
    .X(_0063_));
 sg13g2_mux2_1 _6063_ (.A0(\logix.ram_r[1051] ),
    .A1(\logix.ram_r[1050] ),
    .S(net220),
    .X(_0064_));
 sg13g2_mux2_1 _6064_ (.A0(\logix.ram_r[1052] ),
    .A1(\logix.ram_r[1051] ),
    .S(_2073_),
    .X(_0065_));
 sg13g2_mux2_1 _6065_ (.A0(\logix.ram_r[1053] ),
    .A1(\logix.ram_r[1052] ),
    .S(_2073_),
    .X(_0066_));
 sg13g2_buf_2 _6066_ (.A(_2071_),
    .X(_2074_));
 sg13g2_mux2_1 _6067_ (.A0(\logix.ram_r[1054] ),
    .A1(\logix.ram_r[1053] ),
    .S(net219),
    .X(_0067_));
 sg13g2_mux2_1 _6068_ (.A0(\logix.ram_r[1055] ),
    .A1(\logix.ram_r[1054] ),
    .S(net219),
    .X(_0068_));
 sg13g2_mux2_1 _6069_ (.A0(\logix.ram_r[1056] ),
    .A1(\logix.ram_r[1055] ),
    .S(net219),
    .X(_0069_));
 sg13g2_mux2_1 _6070_ (.A0(\logix.ram_r[1057] ),
    .A1(\logix.ram_r[1056] ),
    .S(net219),
    .X(_0070_));
 sg13g2_mux2_1 _6071_ (.A0(\logix.ram_r[1058] ),
    .A1(\logix.ram_r[1057] ),
    .S(net219),
    .X(_0071_));
 sg13g2_mux2_1 _6072_ (.A0(\logix.ram_r[1059] ),
    .A1(\logix.ram_r[1058] ),
    .S(net219),
    .X(_0072_));
 sg13g2_mux2_1 _6073_ (.A0(\logix.ram_r[105] ),
    .A1(\logix.ram_r[104] ),
    .S(net219),
    .X(_0073_));
 sg13g2_mux2_1 _6074_ (.A0(\logix.ram_r[1060] ),
    .A1(\logix.ram_r[1059] ),
    .S(_2074_),
    .X(_0074_));
 sg13g2_mux2_1 _6075_ (.A0(\logix.ram_r[1061] ),
    .A1(\logix.ram_r[1060] ),
    .S(_2074_),
    .X(_0075_));
 sg13g2_mux2_1 _6076_ (.A0(\logix.ram_r[1062] ),
    .A1(\logix.ram_r[1061] ),
    .S(net219),
    .X(_0076_));
 sg13g2_buf_2 _6077_ (.A(_2071_),
    .X(_2075_));
 sg13g2_mux2_1 _6078_ (.A0(\logix.ram_r[1063] ),
    .A1(\logix.ram_r[1062] ),
    .S(net218),
    .X(_0077_));
 sg13g2_mux2_1 _6079_ (.A0(\logix.ram_r[1064] ),
    .A1(\logix.ram_r[1063] ),
    .S(net218),
    .X(_0078_));
 sg13g2_mux2_1 _6080_ (.A0(\logix.ram_r[1065] ),
    .A1(\logix.ram_r[1064] ),
    .S(_2075_),
    .X(_0079_));
 sg13g2_mux2_1 _6081_ (.A0(\logix.ram_r[1066] ),
    .A1(\logix.ram_r[1065] ),
    .S(net218),
    .X(_0080_));
 sg13g2_mux2_1 _6082_ (.A0(\logix.ram_r[1067] ),
    .A1(\logix.ram_r[1066] ),
    .S(_2075_),
    .X(_0081_));
 sg13g2_mux2_1 _6083_ (.A0(\logix.ram_r[1068] ),
    .A1(\logix.ram_r[1067] ),
    .S(net218),
    .X(_0082_));
 sg13g2_mux2_1 _6084_ (.A0(\logix.ram_r[1069] ),
    .A1(\logix.ram_r[1068] ),
    .S(net218),
    .X(_0083_));
 sg13g2_mux2_1 _6085_ (.A0(\logix.ram_r[106] ),
    .A1(\logix.ram_r[105] ),
    .S(net218),
    .X(_0084_));
 sg13g2_mux2_1 _6086_ (.A0(\logix.ram_r[1070] ),
    .A1(\logix.ram_r[1069] ),
    .S(net218),
    .X(_0085_));
 sg13g2_mux2_1 _6087_ (.A0(\logix.ram_r[1071] ),
    .A1(\logix.ram_r[1070] ),
    .S(net218),
    .X(_0086_));
 sg13g2_buf_2 _6088_ (.A(_2071_),
    .X(_2076_));
 sg13g2_mux2_1 _6089_ (.A0(\logix.ram_r[1072] ),
    .A1(\logix.ram_r[1071] ),
    .S(net217),
    .X(_0087_));
 sg13g2_mux2_1 _6090_ (.A0(\logix.ram_r[1073] ),
    .A1(\logix.ram_r[1072] ),
    .S(_2076_),
    .X(_0088_));
 sg13g2_mux2_1 _6091_ (.A0(\logix.ram_r[1074] ),
    .A1(\logix.ram_r[1073] ),
    .S(net217),
    .X(_0089_));
 sg13g2_mux2_1 _6092_ (.A0(\logix.ram_r[1075] ),
    .A1(\logix.ram_r[1074] ),
    .S(net217),
    .X(_0090_));
 sg13g2_mux2_1 _6093_ (.A0(\logix.ram_r[1076] ),
    .A1(\logix.ram_r[1075] ),
    .S(_2076_),
    .X(_0091_));
 sg13g2_mux2_1 _6094_ (.A0(\logix.ram_r[1077] ),
    .A1(\logix.ram_r[1076] ),
    .S(net217),
    .X(_0092_));
 sg13g2_mux2_1 _6095_ (.A0(\logix.ram_r[1078] ),
    .A1(\logix.ram_r[1077] ),
    .S(net217),
    .X(_0093_));
 sg13g2_mux2_1 _6096_ (.A0(\logix.ram_r[1079] ),
    .A1(\logix.ram_r[1078] ),
    .S(net217),
    .X(_0094_));
 sg13g2_mux2_1 _6097_ (.A0(\logix.ram_r[107] ),
    .A1(\logix.ram_r[106] ),
    .S(net217),
    .X(_0095_));
 sg13g2_mux2_1 _6098_ (.A0(\logix.ram_r[1080] ),
    .A1(\logix.ram_r[1079] ),
    .S(net217),
    .X(_0096_));
 sg13g2_buf_2 _6099_ (.A(_2071_),
    .X(_2077_));
 sg13g2_mux2_1 _6100_ (.A0(\logix.ram_r[1081] ),
    .A1(\logix.ram_r[1080] ),
    .S(_2077_),
    .X(_0097_));
 sg13g2_mux2_1 _6101_ (.A0(\logix.ram_r[1082] ),
    .A1(\logix.ram_r[1081] ),
    .S(net216),
    .X(_0098_));
 sg13g2_mux2_1 _6102_ (.A0(\logix.ram_r[1083] ),
    .A1(\logix.ram_r[1082] ),
    .S(net216),
    .X(_0099_));
 sg13g2_mux2_1 _6103_ (.A0(\logix.ram_r[1084] ),
    .A1(\logix.ram_r[1083] ),
    .S(_2077_),
    .X(_0100_));
 sg13g2_mux2_1 _6104_ (.A0(\logix.ram_r[1085] ),
    .A1(\logix.ram_r[1084] ),
    .S(net216),
    .X(_0101_));
 sg13g2_mux2_1 _6105_ (.A0(\logix.ram_r[1086] ),
    .A1(\logix.ram_r[1085] ),
    .S(net216),
    .X(_0102_));
 sg13g2_mux2_1 _6106_ (.A0(\logix.ram_r[1087] ),
    .A1(\logix.ram_r[1086] ),
    .S(net216),
    .X(_0103_));
 sg13g2_mux2_1 _6107_ (.A0(\logix.ram_r[1088] ),
    .A1(\logix.ram_r[1087] ),
    .S(net216),
    .X(_0104_));
 sg13g2_mux2_1 _6108_ (.A0(\logix.ram_r[1089] ),
    .A1(\logix.ram_r[1088] ),
    .S(net216),
    .X(_0105_));
 sg13g2_mux2_1 _6109_ (.A0(\logix.ram_r[108] ),
    .A1(\logix.ram_r[107] ),
    .S(net216),
    .X(_0106_));
 sg13g2_buf_2 _6110_ (.A(_2071_),
    .X(_2078_));
 sg13g2_mux2_1 _6111_ (.A0(\logix.ram_r[1090] ),
    .A1(\logix.ram_r[1089] ),
    .S(net215),
    .X(_0107_));
 sg13g2_mux2_1 _6112_ (.A0(\logix.ram_r[1091] ),
    .A1(\logix.ram_r[1090] ),
    .S(net215),
    .X(_0108_));
 sg13g2_mux2_1 _6113_ (.A0(\logix.ram_r[1092] ),
    .A1(\logix.ram_r[1091] ),
    .S(net215),
    .X(_0109_));
 sg13g2_mux2_1 _6114_ (.A0(\logix.ram_r[1093] ),
    .A1(\logix.ram_r[1092] ),
    .S(net215),
    .X(_0110_));
 sg13g2_mux2_1 _6115_ (.A0(\logix.ram_r[1094] ),
    .A1(\logix.ram_r[1093] ),
    .S(net215),
    .X(_0111_));
 sg13g2_mux2_1 _6116_ (.A0(\logix.ram_r[1095] ),
    .A1(\logix.ram_r[1094] ),
    .S(net215),
    .X(_0112_));
 sg13g2_mux2_1 _6117_ (.A0(\logix.ram_r[1096] ),
    .A1(\logix.ram_r[1095] ),
    .S(net215),
    .X(_0113_));
 sg13g2_mux2_1 _6118_ (.A0(\logix.ram_r[1097] ),
    .A1(\logix.ram_r[1096] ),
    .S(_2078_),
    .X(_0114_));
 sg13g2_mux2_1 _6119_ (.A0(\logix.ram_r[1098] ),
    .A1(\logix.ram_r[1097] ),
    .S(_2078_),
    .X(_0115_));
 sg13g2_mux2_1 _6120_ (.A0(\logix.ram_r[1099] ),
    .A1(\logix.ram_r[1098] ),
    .S(net215),
    .X(_0116_));
 sg13g2_buf_1 _6121_ (.A(_2070_),
    .X(_2079_));
 sg13g2_buf_2 _6122_ (.A(_2079_),
    .X(_2080_));
 sg13g2_mux2_1 _6123_ (.A0(\logix.ram_r[109] ),
    .A1(\logix.ram_r[108] ),
    .S(_2080_),
    .X(_0117_));
 sg13g2_mux2_1 _6124_ (.A0(\logix.ram_r[10] ),
    .A1(\logix.ram_r[9] ),
    .S(_2080_),
    .X(_0118_));
 sg13g2_mux2_1 _6125_ (.A0(\logix.ram_r[1100] ),
    .A1(\logix.ram_r[1099] ),
    .S(net214),
    .X(_0119_));
 sg13g2_mux2_1 _6126_ (.A0(\logix.ram_r[1101] ),
    .A1(\logix.ram_r[1100] ),
    .S(net214),
    .X(_0120_));
 sg13g2_mux2_1 _6127_ (.A0(\logix.ram_r[1102] ),
    .A1(\logix.ram_r[1101] ),
    .S(net214),
    .X(_0121_));
 sg13g2_mux2_1 _6128_ (.A0(\logix.ram_r[1103] ),
    .A1(\logix.ram_r[1102] ),
    .S(net214),
    .X(_0122_));
 sg13g2_mux2_1 _6129_ (.A0(\logix.ram_r[1104] ),
    .A1(\logix.ram_r[1103] ),
    .S(net214),
    .X(_0123_));
 sg13g2_mux2_1 _6130_ (.A0(\logix.ram_r[1105] ),
    .A1(\logix.ram_r[1104] ),
    .S(net214),
    .X(_0124_));
 sg13g2_mux2_1 _6131_ (.A0(\logix.ram_r[1106] ),
    .A1(\logix.ram_r[1105] ),
    .S(net214),
    .X(_0125_));
 sg13g2_mux2_1 _6132_ (.A0(\logix.ram_r[1107] ),
    .A1(\logix.ram_r[1106] ),
    .S(net214),
    .X(_0126_));
 sg13g2_buf_2 _6133_ (.A(_2079_),
    .X(_2081_));
 sg13g2_mux2_1 _6134_ (.A0(\logix.ram_r[1108] ),
    .A1(\logix.ram_r[1107] ),
    .S(net213),
    .X(_0127_));
 sg13g2_mux2_1 _6135_ (.A0(\logix.ram_r[1109] ),
    .A1(\logix.ram_r[1108] ),
    .S(net213),
    .X(_0128_));
 sg13g2_mux2_1 _6136_ (.A0(\logix.ram_r[110] ),
    .A1(\logix.ram_r[109] ),
    .S(_2081_),
    .X(_0129_));
 sg13g2_mux2_1 _6137_ (.A0(\logix.ram_r[1110] ),
    .A1(\logix.ram_r[1109] ),
    .S(net213),
    .X(_0130_));
 sg13g2_mux2_1 _6138_ (.A0(\logix.ram_r[1111] ),
    .A1(\logix.ram_r[1110] ),
    .S(net213),
    .X(_0131_));
 sg13g2_mux2_1 _6139_ (.A0(\logix.ram_r[1112] ),
    .A1(\logix.ram_r[1111] ),
    .S(net213),
    .X(_0132_));
 sg13g2_mux2_1 _6140_ (.A0(\logix.ram_r[1113] ),
    .A1(\logix.ram_r[1112] ),
    .S(net213),
    .X(_0133_));
 sg13g2_mux2_1 _6141_ (.A0(\logix.ram_r[1114] ),
    .A1(\logix.ram_r[1113] ),
    .S(_2081_),
    .X(_0134_));
 sg13g2_mux2_1 _6142_ (.A0(\logix.ram_r[1115] ),
    .A1(\logix.ram_r[1114] ),
    .S(net213),
    .X(_0135_));
 sg13g2_mux2_1 _6143_ (.A0(\logix.ram_r[1116] ),
    .A1(\logix.ram_r[1115] ),
    .S(net213),
    .X(_0136_));
 sg13g2_buf_2 _6144_ (.A(_2079_),
    .X(_2082_));
 sg13g2_mux2_1 _6145_ (.A0(\logix.ram_r[1117] ),
    .A1(\logix.ram_r[1116] ),
    .S(net212),
    .X(_0137_));
 sg13g2_mux2_1 _6146_ (.A0(\logix.ram_r[1118] ),
    .A1(\logix.ram_r[1117] ),
    .S(net212),
    .X(_0138_));
 sg13g2_mux2_1 _6147_ (.A0(\logix.ram_r[1119] ),
    .A1(\logix.ram_r[1118] ),
    .S(net212),
    .X(_0139_));
 sg13g2_mux2_1 _6148_ (.A0(\logix.ram_r[111] ),
    .A1(\logix.ram_r[110] ),
    .S(_2082_),
    .X(_0140_));
 sg13g2_mux2_1 _6149_ (.A0(\logix.ram_r[1120] ),
    .A1(\logix.ram_r[1119] ),
    .S(net212),
    .X(_0141_));
 sg13g2_mux2_1 _6150_ (.A0(\logix.ram_r[1121] ),
    .A1(\logix.ram_r[1120] ),
    .S(net212),
    .X(_0142_));
 sg13g2_mux2_1 _6151_ (.A0(\logix.ram_r[1122] ),
    .A1(\logix.ram_r[1121] ),
    .S(net212),
    .X(_0143_));
 sg13g2_mux2_1 _6152_ (.A0(\logix.ram_r[1123] ),
    .A1(\logix.ram_r[1122] ),
    .S(net212),
    .X(_0144_));
 sg13g2_mux2_1 _6153_ (.A0(\logix.ram_r[1124] ),
    .A1(\logix.ram_r[1123] ),
    .S(net212),
    .X(_0145_));
 sg13g2_mux2_1 _6154_ (.A0(\logix.ram_r[1125] ),
    .A1(\logix.ram_r[1124] ),
    .S(_2082_),
    .X(_0146_));
 sg13g2_buf_2 _6155_ (.A(_2079_),
    .X(_2083_));
 sg13g2_mux2_1 _6156_ (.A0(\logix.ram_r[1126] ),
    .A1(\logix.ram_r[1125] ),
    .S(net211),
    .X(_0147_));
 sg13g2_mux2_1 _6157_ (.A0(\logix.ram_r[1127] ),
    .A1(\logix.ram_r[1126] ),
    .S(net211),
    .X(_0148_));
 sg13g2_mux2_1 _6158_ (.A0(\logix.ram_r[1128] ),
    .A1(\logix.ram_r[1127] ),
    .S(net211),
    .X(_0149_));
 sg13g2_mux2_1 _6159_ (.A0(\logix.ram_r[1129] ),
    .A1(\logix.ram_r[1128] ),
    .S(net211),
    .X(_0150_));
 sg13g2_mux2_1 _6160_ (.A0(\logix.ram_r[112] ),
    .A1(\logix.ram_r[111] ),
    .S(_2083_),
    .X(_0151_));
 sg13g2_mux2_1 _6161_ (.A0(\logix.ram_r[1130] ),
    .A1(\logix.ram_r[1129] ),
    .S(net211),
    .X(_0152_));
 sg13g2_mux2_1 _6162_ (.A0(\logix.ram_r[1131] ),
    .A1(\logix.ram_r[1130] ),
    .S(net211),
    .X(_0153_));
 sg13g2_mux2_1 _6163_ (.A0(\logix.ram_r[1132] ),
    .A1(\logix.ram_r[1131] ),
    .S(net211),
    .X(_0154_));
 sg13g2_mux2_1 _6164_ (.A0(\logix.ram_r[1133] ),
    .A1(\logix.ram_r[1132] ),
    .S(_2083_),
    .X(_0155_));
 sg13g2_mux2_1 _6165_ (.A0(\logix.ram_r[1134] ),
    .A1(\logix.ram_r[1133] ),
    .S(net211),
    .X(_0156_));
 sg13g2_buf_2 _6166_ (.A(_2079_),
    .X(_2084_));
 sg13g2_mux2_1 _6167_ (.A0(\logix.ram_r[1135] ),
    .A1(\logix.ram_r[1134] ),
    .S(net210),
    .X(_0157_));
 sg13g2_mux2_1 _6168_ (.A0(\logix.ram_r[1136] ),
    .A1(\logix.ram_r[1135] ),
    .S(net210),
    .X(_0158_));
 sg13g2_mux2_1 _6169_ (.A0(\logix.ram_r[1137] ),
    .A1(\logix.ram_r[1136] ),
    .S(net210),
    .X(_0159_));
 sg13g2_mux2_1 _6170_ (.A0(\logix.ram_r[1138] ),
    .A1(\logix.ram_r[1137] ),
    .S(net210),
    .X(_0160_));
 sg13g2_mux2_1 _6171_ (.A0(\logix.ram_r[1139] ),
    .A1(\logix.ram_r[1138] ),
    .S(net210),
    .X(_0161_));
 sg13g2_mux2_1 _6172_ (.A0(\logix.ram_r[113] ),
    .A1(\logix.ram_r[112] ),
    .S(_2084_),
    .X(_0162_));
 sg13g2_mux2_1 _6173_ (.A0(\logix.ram_r[1140] ),
    .A1(\logix.ram_r[1139] ),
    .S(net210),
    .X(_0163_));
 sg13g2_mux2_1 _6174_ (.A0(\logix.ram_r[1141] ),
    .A1(\logix.ram_r[1140] ),
    .S(_2084_),
    .X(_0164_));
 sg13g2_mux2_1 _6175_ (.A0(\logix.ram_r[1142] ),
    .A1(\logix.ram_r[1141] ),
    .S(net210),
    .X(_0165_));
 sg13g2_mux2_1 _6176_ (.A0(\logix.ram_r[1143] ),
    .A1(\logix.ram_r[1142] ),
    .S(net210),
    .X(_0166_));
 sg13g2_buf_2 _6177_ (.A(_2079_),
    .X(_2085_));
 sg13g2_mux2_1 _6178_ (.A0(\logix.ram_r[1144] ),
    .A1(\logix.ram_r[1143] ),
    .S(net209),
    .X(_0167_));
 sg13g2_mux2_1 _6179_ (.A0(\logix.ram_r[1145] ),
    .A1(\logix.ram_r[1144] ),
    .S(net209),
    .X(_0168_));
 sg13g2_mux2_1 _6180_ (.A0(\logix.ram_r[1146] ),
    .A1(\logix.ram_r[1145] ),
    .S(net209),
    .X(_0169_));
 sg13g2_mux2_1 _6181_ (.A0(\logix.ram_r[1147] ),
    .A1(\logix.ram_r[1146] ),
    .S(net209),
    .X(_0170_));
 sg13g2_mux2_1 _6182_ (.A0(\logix.ram_r[1148] ),
    .A1(\logix.ram_r[1147] ),
    .S(net209),
    .X(_0171_));
 sg13g2_mux2_1 _6183_ (.A0(\logix.ram_r[1149] ),
    .A1(\logix.ram_r[1148] ),
    .S(_2085_),
    .X(_0172_));
 sg13g2_mux2_1 _6184_ (.A0(\logix.ram_r[114] ),
    .A1(\logix.ram_r[113] ),
    .S(_2085_),
    .X(_0173_));
 sg13g2_mux2_1 _6185_ (.A0(\logix.ram_r[1150] ),
    .A1(\logix.ram_r[1149] ),
    .S(net209),
    .X(_0174_));
 sg13g2_mux2_1 _6186_ (.A0(\logix.ram_r[1151] ),
    .A1(\logix.ram_r[1150] ),
    .S(net209),
    .X(_0175_));
 sg13g2_mux2_1 _6187_ (.A0(\logix.ram_r[1152] ),
    .A1(\logix.ram_r[1151] ),
    .S(net209),
    .X(_0176_));
 sg13g2_buf_2 _6188_ (.A(_2079_),
    .X(_2086_));
 sg13g2_mux2_1 _6189_ (.A0(\logix.ram_r[1153] ),
    .A1(\logix.ram_r[1152] ),
    .S(net208),
    .X(_0177_));
 sg13g2_mux2_1 _6190_ (.A0(\logix.ram_r[1154] ),
    .A1(\logix.ram_r[1153] ),
    .S(net208),
    .X(_0178_));
 sg13g2_mux2_1 _6191_ (.A0(\logix.ram_r[1155] ),
    .A1(\logix.ram_r[1154] ),
    .S(net208),
    .X(_0179_));
 sg13g2_mux2_1 _6192_ (.A0(\logix.ram_r[1156] ),
    .A1(\logix.ram_r[1155] ),
    .S(net208),
    .X(_0180_));
 sg13g2_mux2_1 _6193_ (.A0(\logix.ram_r[1157] ),
    .A1(\logix.ram_r[1156] ),
    .S(net208),
    .X(_0181_));
 sg13g2_mux2_1 _6194_ (.A0(\logix.ram_r[1158] ),
    .A1(\logix.ram_r[1157] ),
    .S(net208),
    .X(_0182_));
 sg13g2_mux2_1 _6195_ (.A0(\logix.ram_r[1159] ),
    .A1(\logix.ram_r[1158] ),
    .S(net208),
    .X(_0183_));
 sg13g2_mux2_1 _6196_ (.A0(\logix.ram_r[115] ),
    .A1(\logix.ram_r[114] ),
    .S(_2086_),
    .X(_0184_));
 sg13g2_mux2_1 _6197_ (.A0(\logix.ram_r[1160] ),
    .A1(\logix.ram_r[1159] ),
    .S(_2086_),
    .X(_0185_));
 sg13g2_mux2_1 _6198_ (.A0(\logix.ram_r[1161] ),
    .A1(\logix.ram_r[1160] ),
    .S(net208),
    .X(_0186_));
 sg13g2_buf_2 _6199_ (.A(_2063_),
    .X(_2087_));
 sg13g2_buf_1 _6200_ (.A(_2087_),
    .X(_2088_));
 sg13g2_buf_2 _6201_ (.A(_2088_),
    .X(_2089_));
 sg13g2_mux2_1 _6202_ (.A0(\logix.ram_r[1162] ),
    .A1(\logix.ram_r[1161] ),
    .S(net408),
    .X(_0187_));
 sg13g2_mux2_1 _6203_ (.A0(\logix.ram_r[1163] ),
    .A1(\logix.ram_r[1162] ),
    .S(net408),
    .X(_0188_));
 sg13g2_mux2_1 _6204_ (.A0(\logix.ram_r[1164] ),
    .A1(\logix.ram_r[1163] ),
    .S(net408),
    .X(_0189_));
 sg13g2_mux2_1 _6205_ (.A0(\logix.ram_r[1165] ),
    .A1(\logix.ram_r[1164] ),
    .S(net408),
    .X(_0190_));
 sg13g2_mux2_1 _6206_ (.A0(\logix.ram_r[1166] ),
    .A1(\logix.ram_r[1165] ),
    .S(_2089_),
    .X(_0191_));
 sg13g2_mux2_1 _6207_ (.A0(\logix.ram_r[1167] ),
    .A1(\logix.ram_r[1166] ),
    .S(net408),
    .X(_0192_));
 sg13g2_mux2_1 _6208_ (.A0(\logix.ram_r[1168] ),
    .A1(\logix.ram_r[1167] ),
    .S(net408),
    .X(_0193_));
 sg13g2_mux2_1 _6209_ (.A0(\logix.ram_r[1169] ),
    .A1(\logix.ram_r[1168] ),
    .S(net408),
    .X(_0194_));
 sg13g2_mux2_1 _6210_ (.A0(\logix.ram_r[116] ),
    .A1(\logix.ram_r[115] ),
    .S(_2089_),
    .X(_0195_));
 sg13g2_mux2_1 _6211_ (.A0(\logix.ram_r[1170] ),
    .A1(\logix.ram_r[1169] ),
    .S(net408),
    .X(_0196_));
 sg13g2_buf_1 _6212_ (.A(_2088_),
    .X(_2090_));
 sg13g2_mux2_1 _6213_ (.A0(\logix.ram_r[1171] ),
    .A1(\logix.ram_r[1170] ),
    .S(net407),
    .X(_0197_));
 sg13g2_mux2_1 _6214_ (.A0(\logix.ram_r[1172] ),
    .A1(\logix.ram_r[1171] ),
    .S(net407),
    .X(_0198_));
 sg13g2_mux2_1 _6215_ (.A0(\logix.ram_r[1173] ),
    .A1(\logix.ram_r[1172] ),
    .S(net407),
    .X(_0199_));
 sg13g2_mux2_1 _6216_ (.A0(\logix.ram_r[1174] ),
    .A1(\logix.ram_r[1173] ),
    .S(net407),
    .X(_0200_));
 sg13g2_mux2_1 _6217_ (.A0(\logix.ram_r[1175] ),
    .A1(\logix.ram_r[1174] ),
    .S(net407),
    .X(_0201_));
 sg13g2_mux2_1 _6218_ (.A0(\logix.ram_r[1176] ),
    .A1(\logix.ram_r[1175] ),
    .S(_2090_),
    .X(_0202_));
 sg13g2_mux2_1 _6219_ (.A0(\logix.ram_r[1177] ),
    .A1(\logix.ram_r[1176] ),
    .S(net407),
    .X(_0203_));
 sg13g2_mux2_1 _6220_ (.A0(\logix.ram_r[1178] ),
    .A1(\logix.ram_r[1177] ),
    .S(net407),
    .X(_0204_));
 sg13g2_mux2_1 _6221_ (.A0(\logix.ram_r[1179] ),
    .A1(\logix.ram_r[1178] ),
    .S(net407),
    .X(_0205_));
 sg13g2_mux2_1 _6222_ (.A0(\logix.ram_r[117] ),
    .A1(\logix.ram_r[116] ),
    .S(_2090_),
    .X(_0206_));
 sg13g2_buf_1 _6223_ (.A(_2088_),
    .X(_2091_));
 sg13g2_mux2_1 _6224_ (.A0(\logix.ram_r[1180] ),
    .A1(\logix.ram_r[1179] ),
    .S(_2091_),
    .X(_0207_));
 sg13g2_mux2_1 _6225_ (.A0(\logix.ram_r[1181] ),
    .A1(\logix.ram_r[1180] ),
    .S(_2091_),
    .X(_0208_));
 sg13g2_mux2_1 _6226_ (.A0(\logix.ram_r[1182] ),
    .A1(\logix.ram_r[1181] ),
    .S(net406),
    .X(_0209_));
 sg13g2_mux2_1 _6227_ (.A0(\logix.ram_r[1183] ),
    .A1(\logix.ram_r[1182] ),
    .S(net406),
    .X(_0210_));
 sg13g2_mux2_1 _6228_ (.A0(\logix.ram_r[1184] ),
    .A1(\logix.ram_r[1183] ),
    .S(net406),
    .X(_0211_));
 sg13g2_mux2_1 _6229_ (.A0(\logix.ram_r[1185] ),
    .A1(\logix.ram_r[1184] ),
    .S(net406),
    .X(_0212_));
 sg13g2_mux2_1 _6230_ (.A0(\logix.ram_r[1186] ),
    .A1(\logix.ram_r[1185] ),
    .S(net406),
    .X(_0213_));
 sg13g2_mux2_1 _6231_ (.A0(\logix.ram_r[1187] ),
    .A1(\logix.ram_r[1186] ),
    .S(net406),
    .X(_0214_));
 sg13g2_mux2_1 _6232_ (.A0(\logix.ram_r[1188] ),
    .A1(\logix.ram_r[1187] ),
    .S(net406),
    .X(_0215_));
 sg13g2_mux2_1 _6233_ (.A0(\logix.ram_r[1189] ),
    .A1(\logix.ram_r[1188] ),
    .S(net406),
    .X(_0216_));
 sg13g2_buf_1 _6234_ (.A(_2088_),
    .X(_2092_));
 sg13g2_mux2_1 _6235_ (.A0(\logix.ram_r[118] ),
    .A1(\logix.ram_r[117] ),
    .S(_2092_),
    .X(_0217_));
 sg13g2_mux2_1 _6236_ (.A0(\logix.ram_r[1190] ),
    .A1(\logix.ram_r[1189] ),
    .S(net405),
    .X(_0218_));
 sg13g2_mux2_1 _6237_ (.A0(\logix.ram_r[1191] ),
    .A1(\logix.ram_r[1190] ),
    .S(net405),
    .X(_0219_));
 sg13g2_mux2_1 _6238_ (.A0(\logix.ram_r[1192] ),
    .A1(\logix.ram_r[1191] ),
    .S(_2092_),
    .X(_0220_));
 sg13g2_mux2_1 _6239_ (.A0(\logix.ram_r[1193] ),
    .A1(\logix.ram_r[1192] ),
    .S(net405),
    .X(_0221_));
 sg13g2_mux2_1 _6240_ (.A0(\logix.ram_r[1194] ),
    .A1(\logix.ram_r[1193] ),
    .S(net405),
    .X(_0222_));
 sg13g2_mux2_1 _6241_ (.A0(\logix.ram_r[1195] ),
    .A1(\logix.ram_r[1194] ),
    .S(net405),
    .X(_0223_));
 sg13g2_mux2_1 _6242_ (.A0(\logix.ram_r[1196] ),
    .A1(\logix.ram_r[1195] ),
    .S(net405),
    .X(_0224_));
 sg13g2_mux2_1 _6243_ (.A0(\logix.ram_r[1197] ),
    .A1(\logix.ram_r[1196] ),
    .S(net405),
    .X(_0225_));
 sg13g2_mux2_1 _6244_ (.A0(\logix.ram_r[1198] ),
    .A1(\logix.ram_r[1197] ),
    .S(net405),
    .X(_0226_));
 sg13g2_buf_2 _6245_ (.A(_2088_),
    .X(_2093_));
 sg13g2_mux2_1 _6246_ (.A0(\logix.ram_r[1199] ),
    .A1(\logix.ram_r[1198] ),
    .S(net404),
    .X(_0227_));
 sg13g2_mux2_1 _6247_ (.A0(\logix.ram_r[119] ),
    .A1(\logix.ram_r[118] ),
    .S(net404),
    .X(_0228_));
 sg13g2_mux2_1 _6248_ (.A0(\logix.ram_r[11] ),
    .A1(\logix.ram_r[10] ),
    .S(_2093_),
    .X(_0229_));
 sg13g2_mux2_1 _6249_ (.A0(\logix.ram_r[1200] ),
    .A1(\logix.ram_r[1199] ),
    .S(net404),
    .X(_0230_));
 sg13g2_mux2_1 _6250_ (.A0(\logix.ram_r[1201] ),
    .A1(\logix.ram_r[1200] ),
    .S(net404),
    .X(_0231_));
 sg13g2_mux2_1 _6251_ (.A0(\logix.ram_r[1202] ),
    .A1(\logix.ram_r[1201] ),
    .S(net404),
    .X(_0232_));
 sg13g2_mux2_1 _6252_ (.A0(\logix.ram_r[1203] ),
    .A1(\logix.ram_r[1202] ),
    .S(net404),
    .X(_0233_));
 sg13g2_mux2_1 _6253_ (.A0(\logix.ram_r[1204] ),
    .A1(\logix.ram_r[1203] ),
    .S(net404),
    .X(_0234_));
 sg13g2_mux2_1 _6254_ (.A0(\logix.ram_r[1205] ),
    .A1(\logix.ram_r[1204] ),
    .S(net404),
    .X(_0235_));
 sg13g2_mux2_1 _6255_ (.A0(\logix.ram_r[1206] ),
    .A1(\logix.ram_r[1205] ),
    .S(_2093_),
    .X(_0236_));
 sg13g2_buf_2 _6256_ (.A(_2088_),
    .X(_2094_));
 sg13g2_mux2_1 _6257_ (.A0(\logix.ram_r[1207] ),
    .A1(\logix.ram_r[1206] ),
    .S(net403),
    .X(_0237_));
 sg13g2_mux2_1 _6258_ (.A0(\logix.ram_r[1208] ),
    .A1(\logix.ram_r[1207] ),
    .S(net403),
    .X(_0238_));
 sg13g2_mux2_1 _6259_ (.A0(\logix.ram_r[1209] ),
    .A1(\logix.ram_r[1208] ),
    .S(net403),
    .X(_0239_));
 sg13g2_mux2_1 _6260_ (.A0(\logix.ram_r[120] ),
    .A1(\logix.ram_r[119] ),
    .S(net403),
    .X(_0240_));
 sg13g2_mux2_1 _6261_ (.A0(\logix.ram_r[1210] ),
    .A1(\logix.ram_r[1209] ),
    .S(net403),
    .X(_0241_));
 sg13g2_mux2_1 _6262_ (.A0(\logix.ram_r[1211] ),
    .A1(\logix.ram_r[1210] ),
    .S(net403),
    .X(_0242_));
 sg13g2_mux2_1 _6263_ (.A0(\logix.ram_r[1212] ),
    .A1(\logix.ram_r[1211] ),
    .S(net403),
    .X(_0243_));
 sg13g2_mux2_1 _6264_ (.A0(\logix.ram_r[1213] ),
    .A1(\logix.ram_r[1212] ),
    .S(net403),
    .X(_0244_));
 sg13g2_mux2_1 _6265_ (.A0(\logix.ram_r[1214] ),
    .A1(\logix.ram_r[1213] ),
    .S(_2094_),
    .X(_0245_));
 sg13g2_mux2_1 _6266_ (.A0(\logix.ram_r[1215] ),
    .A1(\logix.ram_r[1214] ),
    .S(_2094_),
    .X(_0246_));
 sg13g2_buf_2 _6267_ (.A(_2088_),
    .X(_2095_));
 sg13g2_mux2_1 _6268_ (.A0(\logix.ram_r[1216] ),
    .A1(\logix.ram_r[1215] ),
    .S(_2095_),
    .X(_0247_));
 sg13g2_mux2_1 _6269_ (.A0(\logix.ram_r[1217] ),
    .A1(\logix.ram_r[1216] ),
    .S(net402),
    .X(_0248_));
 sg13g2_mux2_1 _6270_ (.A0(\logix.ram_r[1218] ),
    .A1(\logix.ram_r[1217] ),
    .S(net402),
    .X(_0249_));
 sg13g2_mux2_1 _6271_ (.A0(\logix.ram_r[1219] ),
    .A1(\logix.ram_r[1218] ),
    .S(net402),
    .X(_0250_));
 sg13g2_mux2_1 _6272_ (.A0(\logix.ram_r[121] ),
    .A1(\logix.ram_r[120] ),
    .S(_2095_),
    .X(_0251_));
 sg13g2_mux2_1 _6273_ (.A0(\logix.ram_r[1220] ),
    .A1(\logix.ram_r[1219] ),
    .S(net402),
    .X(_0252_));
 sg13g2_mux2_1 _6274_ (.A0(\logix.ram_r[1221] ),
    .A1(\logix.ram_r[1220] ),
    .S(net402),
    .X(_0253_));
 sg13g2_mux2_1 _6275_ (.A0(\logix.ram_r[1222] ),
    .A1(\logix.ram_r[1221] ),
    .S(net402),
    .X(_0254_));
 sg13g2_mux2_1 _6276_ (.A0(\logix.ram_r[1223] ),
    .A1(\logix.ram_r[1222] ),
    .S(net402),
    .X(_0255_));
 sg13g2_mux2_1 _6277_ (.A0(\logix.ram_r[1224] ),
    .A1(\logix.ram_r[1223] ),
    .S(net402),
    .X(_0256_));
 sg13g2_buf_1 _6278_ (.A(_2087_),
    .X(_2096_));
 sg13g2_buf_2 _6279_ (.A(_2096_),
    .X(_2097_));
 sg13g2_mux2_1 _6280_ (.A0(\logix.ram_r[1225] ),
    .A1(\logix.ram_r[1224] ),
    .S(net401),
    .X(_0257_));
 sg13g2_mux2_1 _6281_ (.A0(\logix.ram_r[1226] ),
    .A1(\logix.ram_r[1225] ),
    .S(net401),
    .X(_0258_));
 sg13g2_mux2_1 _6282_ (.A0(\logix.ram_r[1227] ),
    .A1(\logix.ram_r[1226] ),
    .S(net401),
    .X(_0259_));
 sg13g2_mux2_1 _6283_ (.A0(\logix.ram_r[1228] ),
    .A1(\logix.ram_r[1227] ),
    .S(net401),
    .X(_0260_));
 sg13g2_mux2_1 _6284_ (.A0(\logix.ram_r[1229] ),
    .A1(\logix.ram_r[1228] ),
    .S(_2097_),
    .X(_0261_));
 sg13g2_mux2_1 _6285_ (.A0(\logix.ram_r[122] ),
    .A1(\logix.ram_r[121] ),
    .S(_2097_),
    .X(_0262_));
 sg13g2_mux2_1 _6286_ (.A0(\logix.ram_r[1230] ),
    .A1(\logix.ram_r[1229] ),
    .S(net401),
    .X(_0263_));
 sg13g2_mux2_1 _6287_ (.A0(\logix.ram_r[1231] ),
    .A1(\logix.ram_r[1230] ),
    .S(net401),
    .X(_0264_));
 sg13g2_mux2_1 _6288_ (.A0(\logix.ram_r[1232] ),
    .A1(\logix.ram_r[1231] ),
    .S(net401),
    .X(_0265_));
 sg13g2_mux2_1 _6289_ (.A0(\logix.ram_r[1233] ),
    .A1(\logix.ram_r[1232] ),
    .S(net401),
    .X(_0266_));
 sg13g2_buf_2 _6290_ (.A(_2096_),
    .X(_2098_));
 sg13g2_mux2_1 _6291_ (.A0(\logix.ram_r[1234] ),
    .A1(\logix.ram_r[1233] ),
    .S(net400),
    .X(_0267_));
 sg13g2_mux2_1 _6292_ (.A0(\logix.ram_r[1235] ),
    .A1(\logix.ram_r[1234] ),
    .S(net400),
    .X(_0268_));
 sg13g2_mux2_1 _6293_ (.A0(\logix.ram_r[1236] ),
    .A1(\logix.ram_r[1235] ),
    .S(net400),
    .X(_0269_));
 sg13g2_mux2_1 _6294_ (.A0(\logix.ram_r[1237] ),
    .A1(\logix.ram_r[1236] ),
    .S(_2098_),
    .X(_0270_));
 sg13g2_mux2_1 _6295_ (.A0(\logix.ram_r[1238] ),
    .A1(\logix.ram_r[1237] ),
    .S(net400),
    .X(_0271_));
 sg13g2_mux2_1 _6296_ (.A0(\logix.ram_r[1239] ),
    .A1(\logix.ram_r[1238] ),
    .S(net400),
    .X(_0272_));
 sg13g2_mux2_1 _6297_ (.A0(\logix.ram_r[123] ),
    .A1(\logix.ram_r[122] ),
    .S(_2098_),
    .X(_0273_));
 sg13g2_mux2_1 _6298_ (.A0(\logix.ram_r[1240] ),
    .A1(\logix.ram_r[1239] ),
    .S(net400),
    .X(_0274_));
 sg13g2_mux2_1 _6299_ (.A0(\logix.ram_r[1241] ),
    .A1(\logix.ram_r[1240] ),
    .S(net400),
    .X(_0275_));
 sg13g2_mux2_1 _6300_ (.A0(\logix.ram_r[1242] ),
    .A1(\logix.ram_r[1241] ),
    .S(net400),
    .X(_0276_));
 sg13g2_buf_2 _6301_ (.A(_2096_),
    .X(_2099_));
 sg13g2_mux2_1 _6302_ (.A0(\logix.ram_r[1243] ),
    .A1(\logix.ram_r[1242] ),
    .S(net399),
    .X(_0277_));
 sg13g2_mux2_1 _6303_ (.A0(\logix.ram_r[1244] ),
    .A1(\logix.ram_r[1243] ),
    .S(net399),
    .X(_0278_));
 sg13g2_mux2_1 _6304_ (.A0(\logix.ram_r[1245] ),
    .A1(\logix.ram_r[1244] ),
    .S(net399),
    .X(_0279_));
 sg13g2_mux2_1 _6305_ (.A0(\logix.ram_r[1246] ),
    .A1(\logix.ram_r[1245] ),
    .S(_2099_),
    .X(_0280_));
 sg13g2_mux2_1 _6306_ (.A0(\logix.ram_r[1247] ),
    .A1(\logix.ram_r[1246] ),
    .S(_2099_),
    .X(_0281_));
 sg13g2_mux2_1 _6307_ (.A0(\logix.ram_r[1248] ),
    .A1(\logix.ram_r[1247] ),
    .S(net399),
    .X(_0282_));
 sg13g2_mux2_1 _6308_ (.A0(\logix.ram_r[1249] ),
    .A1(\logix.ram_r[1248] ),
    .S(net399),
    .X(_0283_));
 sg13g2_mux2_1 _6309_ (.A0(\logix.ram_r[124] ),
    .A1(\logix.ram_r[123] ),
    .S(net399),
    .X(_0284_));
 sg13g2_mux2_1 _6310_ (.A0(\logix.ram_r[1250] ),
    .A1(\logix.ram_r[1249] ),
    .S(net399),
    .X(_0285_));
 sg13g2_mux2_1 _6311_ (.A0(\logix.ram_r[1251] ),
    .A1(\logix.ram_r[1250] ),
    .S(net399),
    .X(_0286_));
 sg13g2_buf_1 _6312_ (.A(_2096_),
    .X(_2100_));
 sg13g2_mux2_1 _6313_ (.A0(\logix.ram_r[1252] ),
    .A1(\logix.ram_r[1251] ),
    .S(net398),
    .X(_0287_));
 sg13g2_mux2_1 _6314_ (.A0(\logix.ram_r[1253] ),
    .A1(\logix.ram_r[1252] ),
    .S(net398),
    .X(_0288_));
 sg13g2_mux2_1 _6315_ (.A0(\logix.ram_r[1254] ),
    .A1(\logix.ram_r[1253] ),
    .S(net398),
    .X(_0289_));
 sg13g2_mux2_1 _6316_ (.A0(\logix.ram_r[1255] ),
    .A1(\logix.ram_r[1254] ),
    .S(net398),
    .X(_0290_));
 sg13g2_mux2_1 _6317_ (.A0(\logix.ram_r[1256] ),
    .A1(\logix.ram_r[1255] ),
    .S(net398),
    .X(_0291_));
 sg13g2_mux2_1 _6318_ (.A0(\logix.ram_r[1257] ),
    .A1(\logix.ram_r[1256] ),
    .S(net398),
    .X(_0292_));
 sg13g2_mux2_1 _6319_ (.A0(\logix.ram_r[1258] ),
    .A1(\logix.ram_r[1257] ),
    .S(net398),
    .X(_0293_));
 sg13g2_mux2_1 _6320_ (.A0(\logix.ram_r[1259] ),
    .A1(\logix.ram_r[1258] ),
    .S(_2100_),
    .X(_0294_));
 sg13g2_mux2_1 _6321_ (.A0(\logix.ram_r[125] ),
    .A1(\logix.ram_r[124] ),
    .S(net398),
    .X(_0295_));
 sg13g2_mux2_1 _6322_ (.A0(\logix.ram_r[1260] ),
    .A1(\logix.ram_r[1259] ),
    .S(_2100_),
    .X(_0296_));
 sg13g2_buf_1 _6323_ (.A(_2096_),
    .X(_2101_));
 sg13g2_mux2_1 _6324_ (.A0(\logix.ram_r[1261] ),
    .A1(\logix.ram_r[1260] ),
    .S(net397),
    .X(_0297_));
 sg13g2_mux2_1 _6325_ (.A0(\logix.ram_r[1262] ),
    .A1(\logix.ram_r[1261] ),
    .S(net397),
    .X(_0298_));
 sg13g2_mux2_1 _6326_ (.A0(\logix.ram_r[1263] ),
    .A1(\logix.ram_r[1262] ),
    .S(net397),
    .X(_0299_));
 sg13g2_mux2_1 _6327_ (.A0(\logix.ram_r[1264] ),
    .A1(\logix.ram_r[1263] ),
    .S(net397),
    .X(_0300_));
 sg13g2_mux2_1 _6328_ (.A0(\logix.ram_r[1265] ),
    .A1(\logix.ram_r[1264] ),
    .S(net397),
    .X(_0301_));
 sg13g2_mux2_1 _6329_ (.A0(\logix.ram_r[1266] ),
    .A1(\logix.ram_r[1265] ),
    .S(net397),
    .X(_0302_));
 sg13g2_mux2_1 _6330_ (.A0(\logix.ram_r[1267] ),
    .A1(\logix.ram_r[1266] ),
    .S(net397),
    .X(_0303_));
 sg13g2_mux2_1 _6331_ (.A0(\logix.ram_r[1268] ),
    .A1(\logix.ram_r[1267] ),
    .S(_2101_),
    .X(_0304_));
 sg13g2_mux2_1 _6332_ (.A0(\logix.ram_r[1269] ),
    .A1(\logix.ram_r[1268] ),
    .S(_2101_),
    .X(_0305_));
 sg13g2_mux2_1 _6333_ (.A0(\logix.ram_r[126] ),
    .A1(\logix.ram_r[125] ),
    .S(net397),
    .X(_0306_));
 sg13g2_buf_1 _6334_ (.A(_2096_),
    .X(_2102_));
 sg13g2_mux2_1 _6335_ (.A0(\logix.ram_r[1270] ),
    .A1(\logix.ram_r[1269] ),
    .S(_2102_),
    .X(_0307_));
 sg13g2_mux2_1 _6336_ (.A0(\logix.ram_r[1271] ),
    .A1(\logix.ram_r[1270] ),
    .S(net396),
    .X(_0308_));
 sg13g2_mux2_1 _6337_ (.A0(\logix.ram_r[1272] ),
    .A1(\logix.ram_r[1271] ),
    .S(net396),
    .X(_0309_));
 sg13g2_mux2_1 _6338_ (.A0(\logix.ram_r[1273] ),
    .A1(\logix.ram_r[1272] ),
    .S(net396),
    .X(_0310_));
 sg13g2_mux2_1 _6339_ (.A0(\logix.ram_r[1274] ),
    .A1(\logix.ram_r[1273] ),
    .S(net396),
    .X(_0311_));
 sg13g2_mux2_1 _6340_ (.A0(\logix.ram_r[1275] ),
    .A1(\logix.ram_r[1274] ),
    .S(net396),
    .X(_0312_));
 sg13g2_mux2_1 _6341_ (.A0(\logix.ram_r[1276] ),
    .A1(\logix.ram_r[1275] ),
    .S(net396),
    .X(_0313_));
 sg13g2_mux2_1 _6342_ (.A0(\logix.ram_r[1277] ),
    .A1(\logix.ram_r[1276] ),
    .S(net396),
    .X(_0314_));
 sg13g2_mux2_1 _6343_ (.A0(\logix.ram_r[1278] ),
    .A1(\logix.ram_r[1277] ),
    .S(_2102_),
    .X(_0315_));
 sg13g2_mux2_1 _6344_ (.A0(\logix.ram_r[1279] ),
    .A1(\logix.ram_r[1278] ),
    .S(net396),
    .X(_0316_));
 sg13g2_buf_2 _6345_ (.A(_2096_),
    .X(_2103_));
 sg13g2_mux2_1 _6346_ (.A0(\logix.ram_r[127] ),
    .A1(\logix.ram_r[126] ),
    .S(_2103_),
    .X(_0317_));
 sg13g2_mux2_1 _6347_ (.A0(\logix.ram_r[1280] ),
    .A1(\logix.ram_r[1279] ),
    .S(_2103_),
    .X(_0318_));
 sg13g2_mux2_1 _6348_ (.A0(\logix.ram_r[1281] ),
    .A1(\logix.ram_r[1280] ),
    .S(net395),
    .X(_0319_));
 sg13g2_mux2_1 _6349_ (.A0(\logix.ram_r[1282] ),
    .A1(\logix.ram_r[1281] ),
    .S(net395),
    .X(_0320_));
 sg13g2_mux2_1 _6350_ (.A0(\logix.ram_r[1283] ),
    .A1(\logix.ram_r[1282] ),
    .S(net395),
    .X(_0321_));
 sg13g2_mux2_1 _6351_ (.A0(\logix.ram_r[1284] ),
    .A1(\logix.ram_r[1283] ),
    .S(net395),
    .X(_0322_));
 sg13g2_mux2_1 _6352_ (.A0(\logix.ram_r[1285] ),
    .A1(\logix.ram_r[1284] ),
    .S(net395),
    .X(_0323_));
 sg13g2_mux2_1 _6353_ (.A0(\logix.ram_r[1286] ),
    .A1(\logix.ram_r[1285] ),
    .S(net395),
    .X(_0324_));
 sg13g2_mux2_1 _6354_ (.A0(\logix.ram_r[1287] ),
    .A1(\logix.ram_r[1286] ),
    .S(net395),
    .X(_0325_));
 sg13g2_mux2_1 _6355_ (.A0(\logix.ram_r[1288] ),
    .A1(\logix.ram_r[1287] ),
    .S(net395),
    .X(_0326_));
 sg13g2_buf_1 _6356_ (.A(_2087_),
    .X(_2104_));
 sg13g2_buf_1 _6357_ (.A(_2104_),
    .X(_2105_));
 sg13g2_mux2_1 _6358_ (.A0(\logix.ram_r[1289] ),
    .A1(\logix.ram_r[1288] ),
    .S(net394),
    .X(_0327_));
 sg13g2_mux2_1 _6359_ (.A0(\logix.ram_r[128] ),
    .A1(\logix.ram_r[127] ),
    .S(_2105_),
    .X(_0328_));
 sg13g2_mux2_1 _6360_ (.A0(\logix.ram_r[1290] ),
    .A1(\logix.ram_r[1289] ),
    .S(net394),
    .X(_0329_));
 sg13g2_mux2_1 _6361_ (.A0(\logix.ram_r[1291] ),
    .A1(\logix.ram_r[1290] ),
    .S(net394),
    .X(_0330_));
 sg13g2_mux2_1 _6362_ (.A0(\logix.ram_r[1292] ),
    .A1(\logix.ram_r[1291] ),
    .S(net394),
    .X(_0331_));
 sg13g2_mux2_1 _6363_ (.A0(\logix.ram_r[1293] ),
    .A1(\logix.ram_r[1292] ),
    .S(net394),
    .X(_0332_));
 sg13g2_mux2_1 _6364_ (.A0(\logix.ram_r[1294] ),
    .A1(\logix.ram_r[1293] ),
    .S(net394),
    .X(_0333_));
 sg13g2_mux2_1 _6365_ (.A0(\logix.ram_r[1295] ),
    .A1(\logix.ram_r[1294] ),
    .S(net394),
    .X(_0334_));
 sg13g2_mux2_1 _6366_ (.A0(\logix.ram_r[1296] ),
    .A1(\logix.ram_r[1295] ),
    .S(net394),
    .X(_0335_));
 sg13g2_mux2_1 _6367_ (.A0(\logix.ram_r[1297] ),
    .A1(\logix.ram_r[1296] ),
    .S(_2105_),
    .X(_0336_));
 sg13g2_buf_1 _6368_ (.A(_2104_),
    .X(_2106_));
 sg13g2_mux2_1 _6369_ (.A0(\logix.ram_r[1298] ),
    .A1(\logix.ram_r[1297] ),
    .S(net393),
    .X(_0337_));
 sg13g2_mux2_1 _6370_ (.A0(\logix.ram_r[1299] ),
    .A1(\logix.ram_r[1298] ),
    .S(net393),
    .X(_0338_));
 sg13g2_mux2_1 _6371_ (.A0(\logix.ram_r[129] ),
    .A1(\logix.ram_r[128] ),
    .S(_2106_),
    .X(_0339_));
 sg13g2_mux2_1 _6372_ (.A0(\logix.ram_r[12] ),
    .A1(\logix.ram_r[11] ),
    .S(_2106_),
    .X(_0340_));
 sg13g2_mux2_1 _6373_ (.A0(\logix.ram_r[1300] ),
    .A1(\logix.ram_r[1299] ),
    .S(net393),
    .X(_0341_));
 sg13g2_mux2_1 _6374_ (.A0(\logix.ram_r[1301] ),
    .A1(\logix.ram_r[1300] ),
    .S(net393),
    .X(_0342_));
 sg13g2_mux2_1 _6375_ (.A0(\logix.ram_r[1302] ),
    .A1(\logix.ram_r[1301] ),
    .S(net393),
    .X(_0343_));
 sg13g2_mux2_1 _6376_ (.A0(\logix.ram_r[1303] ),
    .A1(\logix.ram_r[1302] ),
    .S(net393),
    .X(_0344_));
 sg13g2_mux2_1 _6377_ (.A0(\logix.ram_r[1304] ),
    .A1(\logix.ram_r[1303] ),
    .S(net393),
    .X(_0345_));
 sg13g2_mux2_1 _6378_ (.A0(\logix.ram_r[1305] ),
    .A1(\logix.ram_r[1304] ),
    .S(net393),
    .X(_0346_));
 sg13g2_buf_1 _6379_ (.A(_2104_),
    .X(_2107_));
 sg13g2_mux2_1 _6380_ (.A0(\logix.ram_r[1306] ),
    .A1(\logix.ram_r[1305] ),
    .S(net392),
    .X(_0347_));
 sg13g2_mux2_1 _6381_ (.A0(\logix.ram_r[1307] ),
    .A1(\logix.ram_r[1306] ),
    .S(net392),
    .X(_0348_));
 sg13g2_mux2_1 _6382_ (.A0(\logix.ram_r[1308] ),
    .A1(\logix.ram_r[1307] ),
    .S(net392),
    .X(_0349_));
 sg13g2_mux2_1 _6383_ (.A0(\logix.ram_r[1309] ),
    .A1(\logix.ram_r[1308] ),
    .S(net392),
    .X(_0350_));
 sg13g2_mux2_1 _6384_ (.A0(\logix.ram_r[130] ),
    .A1(\logix.ram_r[129] ),
    .S(_2107_),
    .X(_0351_));
 sg13g2_mux2_1 _6385_ (.A0(\logix.ram_r[1310] ),
    .A1(\logix.ram_r[1309] ),
    .S(net392),
    .X(_0352_));
 sg13g2_mux2_1 _6386_ (.A0(\logix.ram_r[1311] ),
    .A1(\logix.ram_r[1310] ),
    .S(net392),
    .X(_0353_));
 sg13g2_mux2_1 _6387_ (.A0(\logix.ram_r[1312] ),
    .A1(\logix.ram_r[1311] ),
    .S(net392),
    .X(_0354_));
 sg13g2_mux2_1 _6388_ (.A0(\logix.ram_r[1313] ),
    .A1(\logix.ram_r[1312] ),
    .S(_2107_),
    .X(_0355_));
 sg13g2_mux2_1 _6389_ (.A0(\logix.ram_r[1314] ),
    .A1(\logix.ram_r[1313] ),
    .S(net392),
    .X(_0356_));
 sg13g2_buf_1 _6390_ (.A(_2104_),
    .X(_2108_));
 sg13g2_mux2_1 _6391_ (.A0(\logix.ram_r[1315] ),
    .A1(\logix.ram_r[1314] ),
    .S(net391),
    .X(_0357_));
 sg13g2_mux2_1 _6392_ (.A0(\logix.ram_r[1316] ),
    .A1(\logix.ram_r[1315] ),
    .S(net391),
    .X(_0358_));
 sg13g2_mux2_1 _6393_ (.A0(\logix.ram_r[1317] ),
    .A1(\logix.ram_r[1316] ),
    .S(net391),
    .X(_0359_));
 sg13g2_mux2_1 _6394_ (.A0(\logix.ram_r[1318] ),
    .A1(\logix.ram_r[1317] ),
    .S(_2108_),
    .X(_0360_));
 sg13g2_mux2_1 _6395_ (.A0(\logix.ram_r[1319] ),
    .A1(\logix.ram_r[1318] ),
    .S(net391),
    .X(_0361_));
 sg13g2_mux2_1 _6396_ (.A0(\logix.ram_r[131] ),
    .A1(\logix.ram_r[130] ),
    .S(_2108_),
    .X(_0362_));
 sg13g2_mux2_1 _6397_ (.A0(\logix.ram_r[1320] ),
    .A1(\logix.ram_r[1319] ),
    .S(net391),
    .X(_0363_));
 sg13g2_mux2_1 _6398_ (.A0(\logix.ram_r[1321] ),
    .A1(\logix.ram_r[1320] ),
    .S(net391),
    .X(_0364_));
 sg13g2_mux2_1 _6399_ (.A0(\logix.ram_r[1322] ),
    .A1(\logix.ram_r[1321] ),
    .S(net391),
    .X(_0365_));
 sg13g2_mux2_1 _6400_ (.A0(\logix.ram_r[1323] ),
    .A1(\logix.ram_r[1322] ),
    .S(net391),
    .X(_0366_));
 sg13g2_buf_1 _6401_ (.A(_2104_),
    .X(_2109_));
 sg13g2_mux2_1 _6402_ (.A0(\logix.ram_r[1324] ),
    .A1(\logix.ram_r[1323] ),
    .S(net390),
    .X(_0367_));
 sg13g2_mux2_1 _6403_ (.A0(\logix.ram_r[1325] ),
    .A1(\logix.ram_r[1324] ),
    .S(net390),
    .X(_0368_));
 sg13g2_mux2_1 _6404_ (.A0(\logix.ram_r[1326] ),
    .A1(\logix.ram_r[1325] ),
    .S(net390),
    .X(_0369_));
 sg13g2_mux2_1 _6405_ (.A0(\logix.ram_r[1327] ),
    .A1(\logix.ram_r[1326] ),
    .S(net390),
    .X(_0370_));
 sg13g2_mux2_1 _6406_ (.A0(\logix.ram_r[1328] ),
    .A1(\logix.ram_r[1327] ),
    .S(_2109_),
    .X(_0371_));
 sg13g2_mux2_1 _6407_ (.A0(\logix.ram_r[1329] ),
    .A1(\logix.ram_r[1328] ),
    .S(net390),
    .X(_0372_));
 sg13g2_mux2_1 _6408_ (.A0(\logix.ram_r[132] ),
    .A1(\logix.ram_r[131] ),
    .S(_2109_),
    .X(_0373_));
 sg13g2_mux2_1 _6409_ (.A0(\logix.ram_r[1330] ),
    .A1(\logix.ram_r[1329] ),
    .S(net390),
    .X(_0374_));
 sg13g2_mux2_1 _6410_ (.A0(\logix.ram_r[1331] ),
    .A1(\logix.ram_r[1330] ),
    .S(net390),
    .X(_0375_));
 sg13g2_mux2_1 _6411_ (.A0(\logix.ram_r[1332] ),
    .A1(\logix.ram_r[1331] ),
    .S(net390),
    .X(_0376_));
 sg13g2_buf_1 _6412_ (.A(_2104_),
    .X(_2110_));
 sg13g2_mux2_1 _6413_ (.A0(\logix.ram_r[1333] ),
    .A1(\logix.ram_r[1332] ),
    .S(net389),
    .X(_0377_));
 sg13g2_mux2_1 _6414_ (.A0(\logix.ram_r[1334] ),
    .A1(\logix.ram_r[1333] ),
    .S(net389),
    .X(_0378_));
 sg13g2_mux2_1 _6415_ (.A0(\logix.ram_r[1335] ),
    .A1(\logix.ram_r[1334] ),
    .S(_2110_),
    .X(_0379_));
 sg13g2_mux2_1 _6416_ (.A0(\logix.ram_r[1336] ),
    .A1(\logix.ram_r[1335] ),
    .S(net389),
    .X(_0380_));
 sg13g2_mux2_1 _6417_ (.A0(\logix.ram_r[1337] ),
    .A1(\logix.ram_r[1336] ),
    .S(net389),
    .X(_0381_));
 sg13g2_mux2_1 _6418_ (.A0(\logix.ram_r[1338] ),
    .A1(\logix.ram_r[1337] ),
    .S(net389),
    .X(_0382_));
 sg13g2_mux2_1 _6419_ (.A0(\logix.ram_r[1339] ),
    .A1(\logix.ram_r[1338] ),
    .S(net389),
    .X(_0383_));
 sg13g2_mux2_1 _6420_ (.A0(\logix.ram_r[133] ),
    .A1(\logix.ram_r[132] ),
    .S(_2110_),
    .X(_0384_));
 sg13g2_mux2_1 _6421_ (.A0(\logix.ram_r[1340] ),
    .A1(\logix.ram_r[1339] ),
    .S(net389),
    .X(_0385_));
 sg13g2_mux2_1 _6422_ (.A0(\logix.ram_r[1341] ),
    .A1(\logix.ram_r[1340] ),
    .S(net389),
    .X(_0386_));
 sg13g2_buf_1 _6423_ (.A(_2104_),
    .X(_2111_));
 sg13g2_mux2_1 _6424_ (.A0(\logix.ram_r[1342] ),
    .A1(\logix.ram_r[1341] ),
    .S(net388),
    .X(_0387_));
 sg13g2_mux2_1 _6425_ (.A0(\logix.ram_r[1343] ),
    .A1(\logix.ram_r[1342] ),
    .S(net388),
    .X(_0388_));
 sg13g2_mux2_1 _6426_ (.A0(\logix.ram_r[1344] ),
    .A1(\logix.ram_r[1343] ),
    .S(net388),
    .X(_0389_));
 sg13g2_mux2_1 _6427_ (.A0(\logix.ram_r[1345] ),
    .A1(\logix.ram_r[1344] ),
    .S(net388),
    .X(_0390_));
 sg13g2_mux2_1 _6428_ (.A0(\logix.ram_r[1346] ),
    .A1(\logix.ram_r[1345] ),
    .S(net388),
    .X(_0391_));
 sg13g2_mux2_1 _6429_ (.A0(\logix.ram_r[1347] ),
    .A1(\logix.ram_r[1346] ),
    .S(net388),
    .X(_0392_));
 sg13g2_mux2_1 _6430_ (.A0(\logix.ram_r[1348] ),
    .A1(\logix.ram_r[1347] ),
    .S(net388),
    .X(_0393_));
 sg13g2_mux2_1 _6431_ (.A0(\logix.ram_r[1349] ),
    .A1(\logix.ram_r[1348] ),
    .S(_2111_),
    .X(_0394_));
 sg13g2_mux2_1 _6432_ (.A0(\logix.ram_r[134] ),
    .A1(\logix.ram_r[133] ),
    .S(net388),
    .X(_0395_));
 sg13g2_mux2_1 _6433_ (.A0(\logix.ram_r[1350] ),
    .A1(\logix.ram_r[1349] ),
    .S(_2111_),
    .X(_0396_));
 sg13g2_buf_1 _6434_ (.A(_2087_),
    .X(_2112_));
 sg13g2_buf_1 _6435_ (.A(_2112_),
    .X(_2113_));
 sg13g2_mux2_1 _6436_ (.A0(\logix.ram_r[1351] ),
    .A1(\logix.ram_r[1350] ),
    .S(net387),
    .X(_0397_));
 sg13g2_mux2_1 _6437_ (.A0(\logix.ram_r[1352] ),
    .A1(\logix.ram_r[1351] ),
    .S(net387),
    .X(_0398_));
 sg13g2_mux2_1 _6438_ (.A0(\logix.ram_r[1353] ),
    .A1(\logix.ram_r[1352] ),
    .S(net387),
    .X(_0399_));
 sg13g2_mux2_1 _6439_ (.A0(\logix.ram_r[1354] ),
    .A1(\logix.ram_r[1353] ),
    .S(net387),
    .X(_0400_));
 sg13g2_mux2_1 _6440_ (.A0(\logix.ram_r[1355] ),
    .A1(\logix.ram_r[1354] ),
    .S(net387),
    .X(_0401_));
 sg13g2_mux2_1 _6441_ (.A0(\logix.ram_r[1356] ),
    .A1(\logix.ram_r[1355] ),
    .S(net387),
    .X(_0402_));
 sg13g2_mux2_1 _6442_ (.A0(\logix.ram_r[1357] ),
    .A1(\logix.ram_r[1356] ),
    .S(net387),
    .X(_0403_));
 sg13g2_mux2_1 _6443_ (.A0(\logix.ram_r[1358] ),
    .A1(\logix.ram_r[1357] ),
    .S(net387),
    .X(_0404_));
 sg13g2_mux2_1 _6444_ (.A0(\logix.ram_r[1359] ),
    .A1(\logix.ram_r[1358] ),
    .S(_2113_),
    .X(_0405_));
 sg13g2_mux2_1 _6445_ (.A0(\logix.ram_r[135] ),
    .A1(\logix.ram_r[134] ),
    .S(_2113_),
    .X(_0406_));
 sg13g2_buf_1 _6446_ (.A(_2112_),
    .X(_2114_));
 sg13g2_mux2_1 _6447_ (.A0(\logix.ram_r[1360] ),
    .A1(\logix.ram_r[1359] ),
    .S(_2114_),
    .X(_0407_));
 sg13g2_mux2_1 _6448_ (.A0(\logix.ram_r[1361] ),
    .A1(\logix.ram_r[1360] ),
    .S(net386),
    .X(_0408_));
 sg13g2_mux2_1 _6449_ (.A0(\logix.ram_r[1362] ),
    .A1(\logix.ram_r[1361] ),
    .S(net386),
    .X(_0409_));
 sg13g2_mux2_1 _6450_ (.A0(\logix.ram_r[1363] ),
    .A1(\logix.ram_r[1362] ),
    .S(net386),
    .X(_0410_));
 sg13g2_mux2_1 _6451_ (.A0(\logix.ram_r[1364] ),
    .A1(\logix.ram_r[1363] ),
    .S(net386),
    .X(_0411_));
 sg13g2_mux2_1 _6452_ (.A0(\logix.ram_r[1365] ),
    .A1(\logix.ram_r[1364] ),
    .S(net386),
    .X(_0412_));
 sg13g2_mux2_1 _6453_ (.A0(\logix.ram_r[1366] ),
    .A1(\logix.ram_r[1365] ),
    .S(net386),
    .X(_0413_));
 sg13g2_mux2_1 _6454_ (.A0(\logix.ram_r[1367] ),
    .A1(\logix.ram_r[1366] ),
    .S(net386),
    .X(_0414_));
 sg13g2_mux2_1 _6455_ (.A0(\logix.ram_r[1368] ),
    .A1(\logix.ram_r[1367] ),
    .S(_2114_),
    .X(_0415_));
 sg13g2_mux2_1 _6456_ (.A0(\logix.ram_r[1369] ),
    .A1(\logix.ram_r[1368] ),
    .S(net386),
    .X(_0416_));
 sg13g2_buf_1 _6457_ (.A(_2112_),
    .X(_2115_));
 sg13g2_mux2_1 _6458_ (.A0(\logix.ram_r[136] ),
    .A1(\logix.ram_r[135] ),
    .S(_2115_),
    .X(_0417_));
 sg13g2_mux2_1 _6459_ (.A0(\logix.ram_r[1370] ),
    .A1(\logix.ram_r[1369] ),
    .S(_2115_),
    .X(_0418_));
 sg13g2_mux2_1 _6460_ (.A0(\logix.ram_r[1371] ),
    .A1(\logix.ram_r[1370] ),
    .S(net385),
    .X(_0419_));
 sg13g2_mux2_1 _6461_ (.A0(\logix.ram_r[1372] ),
    .A1(\logix.ram_r[1371] ),
    .S(net385),
    .X(_0420_));
 sg13g2_mux2_1 _6462_ (.A0(\logix.ram_r[1373] ),
    .A1(\logix.ram_r[1372] ),
    .S(net385),
    .X(_0421_));
 sg13g2_mux2_1 _6463_ (.A0(\logix.ram_r[1374] ),
    .A1(\logix.ram_r[1373] ),
    .S(net385),
    .X(_0422_));
 sg13g2_mux2_1 _6464_ (.A0(\logix.ram_r[1375] ),
    .A1(\logix.ram_r[1374] ),
    .S(net385),
    .X(_0423_));
 sg13g2_mux2_1 _6465_ (.A0(\logix.ram_r[1376] ),
    .A1(\logix.ram_r[1375] ),
    .S(net385),
    .X(_0424_));
 sg13g2_mux2_1 _6466_ (.A0(\logix.ram_r[1377] ),
    .A1(\logix.ram_r[1376] ),
    .S(net385),
    .X(_0425_));
 sg13g2_mux2_1 _6467_ (.A0(\logix.ram_r[1378] ),
    .A1(\logix.ram_r[1377] ),
    .S(net385),
    .X(_0426_));
 sg13g2_buf_1 _6468_ (.A(_2112_),
    .X(_2116_));
 sg13g2_mux2_1 _6469_ (.A0(\logix.ram_r[1379] ),
    .A1(\logix.ram_r[1378] ),
    .S(net384),
    .X(_0427_));
 sg13g2_mux2_1 _6470_ (.A0(\logix.ram_r[137] ),
    .A1(\logix.ram_r[136] ),
    .S(_2116_),
    .X(_0428_));
 sg13g2_mux2_1 _6471_ (.A0(\logix.ram_r[1380] ),
    .A1(\logix.ram_r[1379] ),
    .S(net384),
    .X(_0429_));
 sg13g2_mux2_1 _6472_ (.A0(\logix.ram_r[1381] ),
    .A1(\logix.ram_r[1380] ),
    .S(net384),
    .X(_0430_));
 sg13g2_mux2_1 _6473_ (.A0(\logix.ram_r[1382] ),
    .A1(\logix.ram_r[1381] ),
    .S(_2116_),
    .X(_0431_));
 sg13g2_mux2_1 _6474_ (.A0(\logix.ram_r[1383] ),
    .A1(\logix.ram_r[1382] ),
    .S(net384),
    .X(_0432_));
 sg13g2_mux2_1 _6475_ (.A0(\logix.ram_r[1384] ),
    .A1(\logix.ram_r[1383] ),
    .S(net384),
    .X(_0433_));
 sg13g2_mux2_1 _6476_ (.A0(\logix.ram_r[1385] ),
    .A1(\logix.ram_r[1384] ),
    .S(net384),
    .X(_0434_));
 sg13g2_mux2_1 _6477_ (.A0(\logix.ram_r[1386] ),
    .A1(\logix.ram_r[1385] ),
    .S(net384),
    .X(_0435_));
 sg13g2_mux2_1 _6478_ (.A0(\logix.ram_r[1387] ),
    .A1(\logix.ram_r[1386] ),
    .S(net384),
    .X(_0436_));
 sg13g2_buf_2 _6479_ (.A(_2112_),
    .X(_2117_));
 sg13g2_mux2_1 _6480_ (.A0(\logix.ram_r[1388] ),
    .A1(\logix.ram_r[1387] ),
    .S(net383),
    .X(_0437_));
 sg13g2_mux2_1 _6481_ (.A0(\logix.ram_r[1389] ),
    .A1(\logix.ram_r[1388] ),
    .S(net383),
    .X(_0438_));
 sg13g2_mux2_1 _6482_ (.A0(\logix.ram_r[138] ),
    .A1(\logix.ram_r[137] ),
    .S(_2117_),
    .X(_0439_));
 sg13g2_mux2_1 _6483_ (.A0(\logix.ram_r[1390] ),
    .A1(\logix.ram_r[1389] ),
    .S(net383),
    .X(_0440_));
 sg13g2_mux2_1 _6484_ (.A0(\logix.ram_r[1391] ),
    .A1(\logix.ram_r[1390] ),
    .S(net383),
    .X(_0441_));
 sg13g2_mux2_1 _6485_ (.A0(\logix.ram_r[1392] ),
    .A1(\logix.ram_r[1391] ),
    .S(_2117_),
    .X(_0442_));
 sg13g2_mux2_1 _6486_ (.A0(\logix.ram_r[1393] ),
    .A1(\logix.ram_r[1392] ),
    .S(net383),
    .X(_0443_));
 sg13g2_mux2_1 _6487_ (.A0(\logix.ram_r[1394] ),
    .A1(\logix.ram_r[1393] ),
    .S(net383),
    .X(_0444_));
 sg13g2_mux2_1 _6488_ (.A0(\logix.ram_r[1395] ),
    .A1(\logix.ram_r[1394] ),
    .S(net383),
    .X(_0445_));
 sg13g2_mux2_1 _6489_ (.A0(\logix.ram_r[1396] ),
    .A1(\logix.ram_r[1395] ),
    .S(net383),
    .X(_0446_));
 sg13g2_buf_2 _6490_ (.A(_2112_),
    .X(_2118_));
 sg13g2_mux2_1 _6491_ (.A0(\logix.ram_r[1397] ),
    .A1(\logix.ram_r[1396] ),
    .S(net382),
    .X(_0447_));
 sg13g2_mux2_1 _6492_ (.A0(\logix.ram_r[1398] ),
    .A1(\logix.ram_r[1397] ),
    .S(net382),
    .X(_0448_));
 sg13g2_mux2_1 _6493_ (.A0(\logix.ram_r[1399] ),
    .A1(\logix.ram_r[1398] ),
    .S(net382),
    .X(_0449_));
 sg13g2_mux2_1 _6494_ (.A0(\logix.ram_r[139] ),
    .A1(\logix.ram_r[138] ),
    .S(_2118_),
    .X(_0450_));
 sg13g2_mux2_1 _6495_ (.A0(\logix.ram_r[13] ),
    .A1(\logix.ram_r[12] ),
    .S(_2118_),
    .X(_0451_));
 sg13g2_mux2_1 _6496_ (.A0(\logix.ram_r[1400] ),
    .A1(\logix.ram_r[1399] ),
    .S(net382),
    .X(_0452_));
 sg13g2_mux2_1 _6497_ (.A0(\logix.ram_r[1401] ),
    .A1(\logix.ram_r[1400] ),
    .S(net382),
    .X(_0453_));
 sg13g2_mux2_1 _6498_ (.A0(\logix.ram_r[1402] ),
    .A1(\logix.ram_r[1401] ),
    .S(net382),
    .X(_0454_));
 sg13g2_mux2_1 _6499_ (.A0(\logix.ram_r[1403] ),
    .A1(\logix.ram_r[1402] ),
    .S(net382),
    .X(_0455_));
 sg13g2_mux2_1 _6500_ (.A0(\logix.ram_r[1404] ),
    .A1(\logix.ram_r[1403] ),
    .S(net382),
    .X(_0456_));
 sg13g2_buf_2 _6501_ (.A(_2112_),
    .X(_2119_));
 sg13g2_mux2_1 _6502_ (.A0(\logix.ram_r[1405] ),
    .A1(\logix.ram_r[1404] ),
    .S(net381),
    .X(_0457_));
 sg13g2_mux2_1 _6503_ (.A0(\logix.ram_r[1406] ),
    .A1(\logix.ram_r[1405] ),
    .S(net381),
    .X(_0458_));
 sg13g2_mux2_1 _6504_ (.A0(\logix.ram_r[1407] ),
    .A1(\logix.ram_r[1406] ),
    .S(net381),
    .X(_0459_));
 sg13g2_mux2_1 _6505_ (.A0(\logix.ram_r[1408] ),
    .A1(\logix.ram_r[1407] ),
    .S(net381),
    .X(_0460_));
 sg13g2_mux2_1 _6506_ (.A0(\logix.ram_r[1409] ),
    .A1(\logix.ram_r[1408] ),
    .S(_2119_),
    .X(_0461_));
 sg13g2_mux2_1 _6507_ (.A0(\logix.ram_r[140] ),
    .A1(\logix.ram_r[139] ),
    .S(net381),
    .X(_0462_));
 sg13g2_mux2_1 _6508_ (.A0(\logix.ram_r[1410] ),
    .A1(\logix.ram_r[1409] ),
    .S(net381),
    .X(_0463_));
 sg13g2_mux2_1 _6509_ (.A0(\logix.ram_r[1411] ),
    .A1(\logix.ram_r[1410] ),
    .S(net381),
    .X(_0464_));
 sg13g2_mux2_1 _6510_ (.A0(\logix.ram_r[1412] ),
    .A1(\logix.ram_r[1411] ),
    .S(net381),
    .X(_0465_));
 sg13g2_mux2_1 _6511_ (.A0(\logix.ram_r[1413] ),
    .A1(\logix.ram_r[1412] ),
    .S(_2119_),
    .X(_0466_));
 sg13g2_buf_1 _6512_ (.A(_2087_),
    .X(_2120_));
 sg13g2_buf_2 _6513_ (.A(_2120_),
    .X(_2121_));
 sg13g2_mux2_1 _6514_ (.A0(\logix.ram_r[1414] ),
    .A1(\logix.ram_r[1413] ),
    .S(net380),
    .X(_0467_));
 sg13g2_mux2_1 _6515_ (.A0(\logix.ram_r[1415] ),
    .A1(\logix.ram_r[1414] ),
    .S(net380),
    .X(_0468_));
 sg13g2_mux2_1 _6516_ (.A0(\logix.ram_r[1416] ),
    .A1(\logix.ram_r[1415] ),
    .S(net380),
    .X(_0469_));
 sg13g2_mux2_1 _6517_ (.A0(\logix.ram_r[1417] ),
    .A1(\logix.ram_r[1416] ),
    .S(net380),
    .X(_0470_));
 sg13g2_mux2_1 _6518_ (.A0(\logix.ram_r[1418] ),
    .A1(\logix.ram_r[1417] ),
    .S(net380),
    .X(_0471_));
 sg13g2_mux2_1 _6519_ (.A0(\logix.ram_r[1419] ),
    .A1(\logix.ram_r[1418] ),
    .S(net380),
    .X(_0472_));
 sg13g2_mux2_1 _6520_ (.A0(\logix.ram_r[141] ),
    .A1(\logix.ram_r[140] ),
    .S(_2121_),
    .X(_0473_));
 sg13g2_mux2_1 _6521_ (.A0(\logix.ram_r[1420] ),
    .A1(\logix.ram_r[1419] ),
    .S(net380),
    .X(_0474_));
 sg13g2_mux2_1 _6522_ (.A0(\logix.ram_r[1421] ),
    .A1(\logix.ram_r[1420] ),
    .S(_2121_),
    .X(_0475_));
 sg13g2_mux2_1 _6523_ (.A0(\logix.ram_r[1422] ),
    .A1(\logix.ram_r[1421] ),
    .S(net380),
    .X(_0476_));
 sg13g2_buf_1 _6524_ (.A(_2120_),
    .X(_2122_));
 sg13g2_mux2_1 _6525_ (.A0(\logix.ram_r[1423] ),
    .A1(\logix.ram_r[1422] ),
    .S(_2122_),
    .X(_0477_));
 sg13g2_mux2_1 _6526_ (.A0(\logix.ram_r[1424] ),
    .A1(\logix.ram_r[1423] ),
    .S(net379),
    .X(_0478_));
 sg13g2_mux2_1 _6527_ (.A0(\logix.ram_r[1425] ),
    .A1(\logix.ram_r[1424] ),
    .S(net379),
    .X(_0479_));
 sg13g2_mux2_1 _6528_ (.A0(\logix.ram_r[1426] ),
    .A1(\logix.ram_r[1425] ),
    .S(net379),
    .X(_0480_));
 sg13g2_mux2_1 _6529_ (.A0(\logix.ram_r[1427] ),
    .A1(\logix.ram_r[1426] ),
    .S(net379),
    .X(_0481_));
 sg13g2_mux2_1 _6530_ (.A0(\logix.ram_r[1428] ),
    .A1(\logix.ram_r[1427] ),
    .S(net379),
    .X(_0482_));
 sg13g2_mux2_1 _6531_ (.A0(\logix.ram_r[1429] ),
    .A1(\logix.ram_r[1428] ),
    .S(net379),
    .X(_0483_));
 sg13g2_mux2_1 _6532_ (.A0(\logix.ram_r[142] ),
    .A1(\logix.ram_r[141] ),
    .S(_2122_),
    .X(_0484_));
 sg13g2_mux2_1 _6533_ (.A0(\logix.ram_r[1430] ),
    .A1(\logix.ram_r[1429] ),
    .S(net379),
    .X(_0485_));
 sg13g2_mux2_1 _6534_ (.A0(\logix.ram_r[1431] ),
    .A1(\logix.ram_r[1430] ),
    .S(net379),
    .X(_0486_));
 sg13g2_buf_2 _6535_ (.A(_2120_),
    .X(_2123_));
 sg13g2_mux2_1 _6536_ (.A0(\logix.ram_r[1432] ),
    .A1(\logix.ram_r[1431] ),
    .S(net378),
    .X(_0487_));
 sg13g2_mux2_1 _6537_ (.A0(\logix.ram_r[1433] ),
    .A1(\logix.ram_r[1432] ),
    .S(net378),
    .X(_0488_));
 sg13g2_mux2_1 _6538_ (.A0(\logix.ram_r[1434] ),
    .A1(\logix.ram_r[1433] ),
    .S(net378),
    .X(_0489_));
 sg13g2_mux2_1 _6539_ (.A0(\logix.ram_r[1435] ),
    .A1(\logix.ram_r[1434] ),
    .S(net378),
    .X(_0490_));
 sg13g2_mux2_1 _6540_ (.A0(\logix.ram_r[1436] ),
    .A1(\logix.ram_r[1435] ),
    .S(net378),
    .X(_0491_));
 sg13g2_mux2_1 _6541_ (.A0(\logix.ram_r[1437] ),
    .A1(\logix.ram_r[1436] ),
    .S(_2123_),
    .X(_0492_));
 sg13g2_mux2_1 _6542_ (.A0(\logix.ram_r[1438] ),
    .A1(\logix.ram_r[1437] ),
    .S(net378),
    .X(_0493_));
 sg13g2_mux2_1 _6543_ (.A0(\logix.ram_r[1439] ),
    .A1(\logix.ram_r[1438] ),
    .S(net378),
    .X(_0494_));
 sg13g2_mux2_1 _6544_ (.A0(\logix.ram_r[143] ),
    .A1(\logix.ram_r[142] ),
    .S(_2123_),
    .X(_0495_));
 sg13g2_mux2_1 _6545_ (.A0(\logix.ram_r[1440] ),
    .A1(\logix.ram_r[1439] ),
    .S(net378),
    .X(_0496_));
 sg13g2_buf_1 _6546_ (.A(_2120_),
    .X(_2124_));
 sg13g2_mux2_1 _6547_ (.A0(\logix.ram_r[1441] ),
    .A1(\logix.ram_r[1440] ),
    .S(net377),
    .X(_0497_));
 sg13g2_mux2_1 _6548_ (.A0(\logix.ram_r[1442] ),
    .A1(\logix.ram_r[1441] ),
    .S(net377),
    .X(_0498_));
 sg13g2_mux2_1 _6549_ (.A0(\logix.ram_r[1443] ),
    .A1(\logix.ram_r[1442] ),
    .S(net377),
    .X(_0499_));
 sg13g2_mux2_1 _6550_ (.A0(\logix.ram_r[1444] ),
    .A1(\logix.ram_r[1443] ),
    .S(net377),
    .X(_0500_));
 sg13g2_mux2_1 _6551_ (.A0(\logix.ram_r[1445] ),
    .A1(\logix.ram_r[1444] ),
    .S(_2124_),
    .X(_0501_));
 sg13g2_mux2_1 _6552_ (.A0(\logix.ram_r[1446] ),
    .A1(\logix.ram_r[1445] ),
    .S(net377),
    .X(_0502_));
 sg13g2_mux2_1 _6553_ (.A0(\logix.ram_r[1447] ),
    .A1(\logix.ram_r[1446] ),
    .S(net377),
    .X(_0503_));
 sg13g2_mux2_1 _6554_ (.A0(\logix.ram_r[1448] ),
    .A1(\logix.ram_r[1447] ),
    .S(net377),
    .X(_0504_));
 sg13g2_mux2_1 _6555_ (.A0(\logix.ram_r[1449] ),
    .A1(\logix.ram_r[1448] ),
    .S(net377),
    .X(_0505_));
 sg13g2_mux2_1 _6556_ (.A0(\logix.ram_r[144] ),
    .A1(\logix.ram_r[143] ),
    .S(_2124_),
    .X(_0506_));
 sg13g2_buf_1 _6557_ (.A(_2120_),
    .X(_2125_));
 sg13g2_mux2_1 _6558_ (.A0(\logix.ram_r[1450] ),
    .A1(\logix.ram_r[1449] ),
    .S(net376),
    .X(_0507_));
 sg13g2_mux2_1 _6559_ (.A0(\logix.ram_r[1451] ),
    .A1(\logix.ram_r[1450] ),
    .S(net376),
    .X(_0508_));
 sg13g2_mux2_1 _6560_ (.A0(\logix.ram_r[1452] ),
    .A1(\logix.ram_r[1451] ),
    .S(net376),
    .X(_0509_));
 sg13g2_mux2_1 _6561_ (.A0(\logix.ram_r[1453] ),
    .A1(\logix.ram_r[1452] ),
    .S(net376),
    .X(_0510_));
 sg13g2_mux2_1 _6562_ (.A0(\logix.ram_r[1454] ),
    .A1(\logix.ram_r[1453] ),
    .S(net376),
    .X(_0511_));
 sg13g2_mux2_1 _6563_ (.A0(\logix.ram_r[1455] ),
    .A1(\logix.ram_r[1454] ),
    .S(_2125_),
    .X(_0512_));
 sg13g2_mux2_1 _6564_ (.A0(\logix.ram_r[1456] ),
    .A1(\logix.ram_r[1455] ),
    .S(_2125_),
    .X(_0513_));
 sg13g2_mux2_1 _6565_ (.A0(\logix.ram_r[1457] ),
    .A1(\logix.ram_r[1456] ),
    .S(net376),
    .X(_0514_));
 sg13g2_mux2_1 _6566_ (.A0(\logix.ram_r[1458] ),
    .A1(\logix.ram_r[1457] ),
    .S(net376),
    .X(_0515_));
 sg13g2_mux2_1 _6567_ (.A0(\logix.ram_r[1459] ),
    .A1(\logix.ram_r[1458] ),
    .S(net376),
    .X(_0516_));
 sg13g2_buf_1 _6568_ (.A(_2120_),
    .X(_2126_));
 sg13g2_mux2_1 _6569_ (.A0(\logix.ram_r[145] ),
    .A1(\logix.ram_r[144] ),
    .S(_2126_),
    .X(_0517_));
 sg13g2_mux2_1 _6570_ (.A0(\logix.ram_r[1460] ),
    .A1(\logix.ram_r[1459] ),
    .S(net375),
    .X(_0518_));
 sg13g2_mux2_1 _6571_ (.A0(\logix.ram_r[1461] ),
    .A1(\logix.ram_r[1460] ),
    .S(net375),
    .X(_0519_));
 sg13g2_mux2_1 _6572_ (.A0(\logix.ram_r[1462] ),
    .A1(\logix.ram_r[1461] ),
    .S(net375),
    .X(_0520_));
 sg13g2_mux2_1 _6573_ (.A0(\logix.ram_r[1463] ),
    .A1(\logix.ram_r[1462] ),
    .S(_2126_),
    .X(_0521_));
 sg13g2_mux2_1 _6574_ (.A0(\logix.ram_r[1464] ),
    .A1(\logix.ram_r[1463] ),
    .S(net375),
    .X(_0522_));
 sg13g2_mux2_1 _6575_ (.A0(\logix.ram_r[1465] ),
    .A1(\logix.ram_r[1464] ),
    .S(net375),
    .X(_0523_));
 sg13g2_mux2_1 _6576_ (.A0(\logix.ram_r[1466] ),
    .A1(\logix.ram_r[1465] ),
    .S(net375),
    .X(_0524_));
 sg13g2_mux2_1 _6577_ (.A0(\logix.ram_r[1467] ),
    .A1(\logix.ram_r[1466] ),
    .S(net375),
    .X(_0525_));
 sg13g2_mux2_1 _6578_ (.A0(\logix.ram_r[1468] ),
    .A1(\logix.ram_r[1467] ),
    .S(net375),
    .X(_0526_));
 sg13g2_buf_2 _6579_ (.A(_2120_),
    .X(_2127_));
 sg13g2_mux2_1 _6580_ (.A0(\logix.ram_r[1469] ),
    .A1(\logix.ram_r[1468] ),
    .S(net374),
    .X(_0527_));
 sg13g2_mux2_1 _6581_ (.A0(\logix.ram_r[146] ),
    .A1(\logix.ram_r[145] ),
    .S(_2127_),
    .X(_0528_));
 sg13g2_mux2_1 _6582_ (.A0(\logix.ram_r[1470] ),
    .A1(\logix.ram_r[1469] ),
    .S(net374),
    .X(_0529_));
 sg13g2_mux2_1 _6583_ (.A0(\logix.ram_r[1471] ),
    .A1(\logix.ram_r[1470] ),
    .S(net374),
    .X(_0530_));
 sg13g2_mux2_1 _6584_ (.A0(\logix.ram_r[1472] ),
    .A1(\logix.ram_r[1471] ),
    .S(net374),
    .X(_0531_));
 sg13g2_mux2_1 _6585_ (.A0(\logix.ram_r[1473] ),
    .A1(\logix.ram_r[1472] ),
    .S(net374),
    .X(_0532_));
 sg13g2_mux2_1 _6586_ (.A0(\logix.ram_r[1474] ),
    .A1(\logix.ram_r[1473] ),
    .S(net374),
    .X(_0533_));
 sg13g2_mux2_1 _6587_ (.A0(\logix.ram_r[1475] ),
    .A1(\logix.ram_r[1474] ),
    .S(net374),
    .X(_0534_));
 sg13g2_mux2_1 _6588_ (.A0(\logix.ram_r[1476] ),
    .A1(\logix.ram_r[1475] ),
    .S(_2127_),
    .X(_0535_));
 sg13g2_mux2_1 _6589_ (.A0(\logix.ram_r[1477] ),
    .A1(\logix.ram_r[1476] ),
    .S(net374),
    .X(_0536_));
 sg13g2_buf_1 _6590_ (.A(_2087_),
    .X(_2128_));
 sg13g2_buf_1 _6591_ (.A(_2128_),
    .X(_2129_));
 sg13g2_mux2_1 _6592_ (.A0(\logix.ram_r[1478] ),
    .A1(\logix.ram_r[1477] ),
    .S(net373),
    .X(_0537_));
 sg13g2_mux2_1 _6593_ (.A0(\logix.ram_r[1479] ),
    .A1(\logix.ram_r[1478] ),
    .S(net373),
    .X(_0538_));
 sg13g2_mux2_1 _6594_ (.A0(\logix.ram_r[147] ),
    .A1(\logix.ram_r[146] ),
    .S(_2129_),
    .X(_0539_));
 sg13g2_mux2_1 _6595_ (.A0(\logix.ram_r[1480] ),
    .A1(\logix.ram_r[1479] ),
    .S(net373),
    .X(_0540_));
 sg13g2_mux2_1 _6596_ (.A0(\logix.ram_r[1481] ),
    .A1(\logix.ram_r[1480] ),
    .S(net373),
    .X(_0541_));
 sg13g2_mux2_1 _6597_ (.A0(\logix.ram_r[1482] ),
    .A1(\logix.ram_r[1481] ),
    .S(net373),
    .X(_0542_));
 sg13g2_mux2_1 _6598_ (.A0(\logix.ram_r[1483] ),
    .A1(\logix.ram_r[1482] ),
    .S(net373),
    .X(_0543_));
 sg13g2_mux2_1 _6599_ (.A0(\logix.ram_r[1484] ),
    .A1(\logix.ram_r[1483] ),
    .S(net373),
    .X(_0544_));
 sg13g2_mux2_1 _6600_ (.A0(\logix.ram_r[1485] ),
    .A1(\logix.ram_r[1484] ),
    .S(net373),
    .X(_0545_));
 sg13g2_mux2_1 _6601_ (.A0(\logix.ram_r[1486] ),
    .A1(\logix.ram_r[1485] ),
    .S(_2129_),
    .X(_0546_));
 sg13g2_buf_2 _6602_ (.A(_2128_),
    .X(_2130_));
 sg13g2_mux2_1 _6603_ (.A0(\logix.ram_r[1487] ),
    .A1(\logix.ram_r[1486] ),
    .S(net372),
    .X(_0547_));
 sg13g2_mux2_1 _6604_ (.A0(\logix.ram_r[1488] ),
    .A1(\logix.ram_r[1487] ),
    .S(net372),
    .X(_0548_));
 sg13g2_mux2_1 _6605_ (.A0(\logix.ram_r[1489] ),
    .A1(\logix.ram_r[1488] ),
    .S(net372),
    .X(_0549_));
 sg13g2_mux2_1 _6606_ (.A0(\logix.ram_r[148] ),
    .A1(\logix.ram_r[147] ),
    .S(_2130_),
    .X(_0550_));
 sg13g2_mux2_1 _6607_ (.A0(\logix.ram_r[1490] ),
    .A1(\logix.ram_r[1489] ),
    .S(net372),
    .X(_0551_));
 sg13g2_mux2_1 _6608_ (.A0(\logix.ram_r[1491] ),
    .A1(\logix.ram_r[1490] ),
    .S(net372),
    .X(_0552_));
 sg13g2_mux2_1 _6609_ (.A0(\logix.ram_r[1492] ),
    .A1(\logix.ram_r[1491] ),
    .S(net372),
    .X(_0553_));
 sg13g2_mux2_1 _6610_ (.A0(\logix.ram_r[1493] ),
    .A1(\logix.ram_r[1492] ),
    .S(net372),
    .X(_0554_));
 sg13g2_mux2_1 _6611_ (.A0(\logix.ram_r[1494] ),
    .A1(\logix.ram_r[1493] ),
    .S(net372),
    .X(_0555_));
 sg13g2_mux2_1 _6612_ (.A0(\logix.ram_r[1495] ),
    .A1(\logix.ram_r[1494] ),
    .S(_2130_),
    .X(_0556_));
 sg13g2_buf_2 _6613_ (.A(_2128_),
    .X(_2131_));
 sg13g2_mux2_1 _6614_ (.A0(\logix.ram_r[1496] ),
    .A1(\logix.ram_r[1495] ),
    .S(net371),
    .X(_0557_));
 sg13g2_mux2_1 _6615_ (.A0(\logix.ram_r[1497] ),
    .A1(\logix.ram_r[1496] ),
    .S(net371),
    .X(_0558_));
 sg13g2_mux2_1 _6616_ (.A0(\logix.ram_r[1498] ),
    .A1(\logix.ram_r[1497] ),
    .S(net371),
    .X(_0559_));
 sg13g2_mux2_1 _6617_ (.A0(\logix.ram_r[1499] ),
    .A1(\logix.ram_r[1498] ),
    .S(net371),
    .X(_0560_));
 sg13g2_mux2_1 _6618_ (.A0(\logix.ram_r[149] ),
    .A1(\logix.ram_r[148] ),
    .S(net371),
    .X(_0561_));
 sg13g2_mux2_1 _6619_ (.A0(\logix.ram_r[14] ),
    .A1(\logix.ram_r[13] ),
    .S(net371),
    .X(_0562_));
 sg13g2_mux2_1 _6620_ (.A0(\logix.ram_r[1500] ),
    .A1(\logix.ram_r[1499] ),
    .S(net371),
    .X(_0563_));
 sg13g2_mux2_1 _6621_ (.A0(\logix.ram_r[1501] ),
    .A1(\logix.ram_r[1500] ),
    .S(net371),
    .X(_0564_));
 sg13g2_mux2_1 _6622_ (.A0(\logix.ram_r[1502] ),
    .A1(\logix.ram_r[1501] ),
    .S(_2131_),
    .X(_0565_));
 sg13g2_mux2_1 _6623_ (.A0(\logix.ram_r[1503] ),
    .A1(\logix.ram_r[1502] ),
    .S(_2131_),
    .X(_0566_));
 sg13g2_buf_2 _6624_ (.A(_2128_),
    .X(_2132_));
 sg13g2_mux2_1 _6625_ (.A0(\logix.ram_r[1504] ),
    .A1(\logix.ram_r[1503] ),
    .S(net370),
    .X(_0567_));
 sg13g2_mux2_1 _6626_ (.A0(\logix.ram_r[1505] ),
    .A1(\logix.ram_r[1504] ),
    .S(net370),
    .X(_0568_));
 sg13g2_mux2_1 _6627_ (.A0(\logix.ram_r[1506] ),
    .A1(\logix.ram_r[1505] ),
    .S(net370),
    .X(_0569_));
 sg13g2_mux2_1 _6628_ (.A0(\logix.ram_r[1507] ),
    .A1(\logix.ram_r[1506] ),
    .S(net370),
    .X(_0570_));
 sg13g2_mux2_1 _6629_ (.A0(\logix.ram_r[1508] ),
    .A1(\logix.ram_r[1507] ),
    .S(net370),
    .X(_0571_));
 sg13g2_mux2_1 _6630_ (.A0(\logix.ram_r[1509] ),
    .A1(\logix.ram_r[1508] ),
    .S(net370),
    .X(_0572_));
 sg13g2_mux2_1 _6631_ (.A0(\logix.ram_r[150] ),
    .A1(\logix.ram_r[149] ),
    .S(_2132_),
    .X(_0573_));
 sg13g2_mux2_1 _6632_ (.A0(\logix.ram_r[1510] ),
    .A1(\logix.ram_r[1509] ),
    .S(net370),
    .X(_0574_));
 sg13g2_mux2_1 _6633_ (.A0(\logix.ram_r[1511] ),
    .A1(\logix.ram_r[1510] ),
    .S(_2132_),
    .X(_0575_));
 sg13g2_mux2_1 _6634_ (.A0(\logix.ram_r[1512] ),
    .A1(\logix.ram_r[1511] ),
    .S(net370),
    .X(_0576_));
 sg13g2_buf_1 _6635_ (.A(_2128_),
    .X(_2133_));
 sg13g2_mux2_1 _6636_ (.A0(\logix.ram_r[1513] ),
    .A1(\logix.ram_r[1512] ),
    .S(net369),
    .X(_0577_));
 sg13g2_mux2_1 _6637_ (.A0(\logix.ram_r[1514] ),
    .A1(\logix.ram_r[1513] ),
    .S(net369),
    .X(_0578_));
 sg13g2_mux2_1 _6638_ (.A0(\logix.ram_r[1515] ),
    .A1(\logix.ram_r[1514] ),
    .S(net369),
    .X(_0579_));
 sg13g2_mux2_1 _6639_ (.A0(\logix.ram_r[1516] ),
    .A1(\logix.ram_r[1515] ),
    .S(net369),
    .X(_0580_));
 sg13g2_mux2_1 _6640_ (.A0(\logix.ram_r[1517] ),
    .A1(\logix.ram_r[1516] ),
    .S(net369),
    .X(_0581_));
 sg13g2_mux2_1 _6641_ (.A0(\logix.ram_r[1518] ),
    .A1(\logix.ram_r[1517] ),
    .S(_2133_),
    .X(_0582_));
 sg13g2_mux2_1 _6642_ (.A0(\logix.ram_r[1519] ),
    .A1(\logix.ram_r[1518] ),
    .S(net369),
    .X(_0583_));
 sg13g2_mux2_1 _6643_ (.A0(\logix.ram_r[151] ),
    .A1(\logix.ram_r[150] ),
    .S(_2133_),
    .X(_0584_));
 sg13g2_mux2_1 _6644_ (.A0(\logix.ram_r[1520] ),
    .A1(\logix.ram_r[1519] ),
    .S(net369),
    .X(_0585_));
 sg13g2_mux2_1 _6645_ (.A0(\logix.ram_r[1521] ),
    .A1(\logix.ram_r[1520] ),
    .S(net369),
    .X(_0586_));
 sg13g2_buf_1 _6646_ (.A(_2128_),
    .X(_2134_));
 sg13g2_mux2_1 _6647_ (.A0(\logix.ram_r[1522] ),
    .A1(\logix.ram_r[1521] ),
    .S(net368),
    .X(_0587_));
 sg13g2_mux2_1 _6648_ (.A0(\logix.ram_r[1523] ),
    .A1(\logix.ram_r[1522] ),
    .S(net368),
    .X(_0588_));
 sg13g2_mux2_1 _6649_ (.A0(\logix.ram_r[1524] ),
    .A1(\logix.ram_r[1523] ),
    .S(net368),
    .X(_0589_));
 sg13g2_mux2_1 _6650_ (.A0(\logix.ram_r[1525] ),
    .A1(\logix.ram_r[1524] ),
    .S(net368),
    .X(_0590_));
 sg13g2_mux2_1 _6651_ (.A0(\logix.ram_r[1526] ),
    .A1(\logix.ram_r[1525] ),
    .S(net368),
    .X(_0591_));
 sg13g2_mux2_1 _6652_ (.A0(\logix.ram_r[1527] ),
    .A1(\logix.ram_r[1526] ),
    .S(net368),
    .X(_0592_));
 sg13g2_mux2_1 _6653_ (.A0(\logix.ram_r[1528] ),
    .A1(\logix.ram_r[1527] ),
    .S(net368),
    .X(_0593_));
 sg13g2_mux2_1 _6654_ (.A0(\logix.ram_r[1529] ),
    .A1(\logix.ram_r[1528] ),
    .S(_2134_),
    .X(_0594_));
 sg13g2_mux2_1 _6655_ (.A0(\logix.ram_r[152] ),
    .A1(\logix.ram_r[151] ),
    .S(_2134_),
    .X(_0595_));
 sg13g2_mux2_1 _6656_ (.A0(\logix.ram_r[1530] ),
    .A1(\logix.ram_r[1529] ),
    .S(net368),
    .X(_0596_));
 sg13g2_buf_2 _6657_ (.A(_2128_),
    .X(_2135_));
 sg13g2_mux2_1 _6658_ (.A0(\logix.ram_r[1531] ),
    .A1(\logix.ram_r[1530] ),
    .S(net367),
    .X(_0597_));
 sg13g2_mux2_1 _6659_ (.A0(\logix.ram_r[1532] ),
    .A1(\logix.ram_r[1531] ),
    .S(net367),
    .X(_0598_));
 sg13g2_mux2_1 _6660_ (.A0(\logix.ram_r[1533] ),
    .A1(\logix.ram_r[1532] ),
    .S(net367),
    .X(_0599_));
 sg13g2_mux2_1 _6661_ (.A0(\logix.ram_r[1534] ),
    .A1(\logix.ram_r[1533] ),
    .S(_2135_),
    .X(_0600_));
 sg13g2_mux2_1 _6662_ (.A0(\logix.ram_r[1535] ),
    .A1(\logix.ram_r[1534] ),
    .S(_2135_),
    .X(_0601_));
 sg13g2_mux2_1 _6663_ (.A0(\logix.ram_r[1536] ),
    .A1(\logix.ram_r[1535] ),
    .S(net367),
    .X(_0602_));
 sg13g2_mux2_1 _6664_ (.A0(\logix.ram_r[1537] ),
    .A1(\logix.ram_r[1536] ),
    .S(net367),
    .X(_0603_));
 sg13g2_mux2_1 _6665_ (.A0(\logix.ram_r[1538] ),
    .A1(\logix.ram_r[1537] ),
    .S(net367),
    .X(_0604_));
 sg13g2_mux2_1 _6666_ (.A0(\logix.ram_r[1539] ),
    .A1(\logix.ram_r[1538] ),
    .S(net367),
    .X(_0605_));
 sg13g2_mux2_1 _6667_ (.A0(\logix.ram_r[153] ),
    .A1(\logix.ram_r[152] ),
    .S(net367),
    .X(_0606_));
 sg13g2_buf_1 _6668_ (.A(_2087_),
    .X(_2136_));
 sg13g2_buf_2 _6669_ (.A(_2136_),
    .X(_2137_));
 sg13g2_mux2_1 _6670_ (.A0(\logix.ram_r[1540] ),
    .A1(\logix.ram_r[1539] ),
    .S(net366),
    .X(_0607_));
 sg13g2_mux2_1 _6671_ (.A0(\logix.ram_r[1541] ),
    .A1(\logix.ram_r[1540] ),
    .S(net366),
    .X(_0608_));
 sg13g2_mux2_1 _6672_ (.A0(\logix.ram_r[1542] ),
    .A1(\logix.ram_r[1541] ),
    .S(net366),
    .X(_0609_));
 sg13g2_mux2_1 _6673_ (.A0(\logix.ram_r[1543] ),
    .A1(\logix.ram_r[1542] ),
    .S(net366),
    .X(_0610_));
 sg13g2_mux2_1 _6674_ (.A0(\logix.ram_r[1544] ),
    .A1(\logix.ram_r[1543] ),
    .S(net366),
    .X(_0611_));
 sg13g2_mux2_1 _6675_ (.A0(\logix.ram_r[1545] ),
    .A1(\logix.ram_r[1544] ),
    .S(_2137_),
    .X(_0612_));
 sg13g2_mux2_1 _6676_ (.A0(\logix.ram_r[1546] ),
    .A1(\logix.ram_r[1545] ),
    .S(_2137_),
    .X(_0613_));
 sg13g2_mux2_1 _6677_ (.A0(\logix.ram_r[1547] ),
    .A1(\logix.ram_r[1546] ),
    .S(net366),
    .X(_0614_));
 sg13g2_mux2_1 _6678_ (.A0(\logix.ram_r[1548] ),
    .A1(\logix.ram_r[1547] ),
    .S(net366),
    .X(_0615_));
 sg13g2_mux2_1 _6679_ (.A0(\logix.ram_r[1549] ),
    .A1(\logix.ram_r[1548] ),
    .S(net366),
    .X(_0616_));
 sg13g2_buf_2 _6680_ (.A(_2136_),
    .X(_2138_));
 sg13g2_mux2_1 _6681_ (.A0(\logix.ram_r[154] ),
    .A1(\logix.ram_r[153] ),
    .S(_2138_),
    .X(_0617_));
 sg13g2_mux2_1 _6682_ (.A0(\logix.ram_r[1550] ),
    .A1(\logix.ram_r[1549] ),
    .S(net365),
    .X(_0618_));
 sg13g2_mux2_1 _6683_ (.A0(\logix.ram_r[1551] ),
    .A1(\logix.ram_r[1550] ),
    .S(net365),
    .X(_0619_));
 sg13g2_mux2_1 _6684_ (.A0(\logix.ram_r[1552] ),
    .A1(\logix.ram_r[1551] ),
    .S(_2138_),
    .X(_0620_));
 sg13g2_mux2_1 _6685_ (.A0(\logix.ram_r[1553] ),
    .A1(\logix.ram_r[1552] ),
    .S(net365),
    .X(_0621_));
 sg13g2_mux2_1 _6686_ (.A0(\logix.ram_r[1554] ),
    .A1(\logix.ram_r[1553] ),
    .S(net365),
    .X(_0622_));
 sg13g2_mux2_1 _6687_ (.A0(\logix.ram_r[1555] ),
    .A1(\logix.ram_r[1554] ),
    .S(net365),
    .X(_0623_));
 sg13g2_mux2_1 _6688_ (.A0(\logix.ram_r[1556] ),
    .A1(\logix.ram_r[1555] ),
    .S(net365),
    .X(_0624_));
 sg13g2_mux2_1 _6689_ (.A0(\logix.ram_r[1557] ),
    .A1(\logix.ram_r[1556] ),
    .S(net365),
    .X(_0625_));
 sg13g2_mux2_1 _6690_ (.A0(\logix.ram_r[1558] ),
    .A1(\logix.ram_r[1557] ),
    .S(net365),
    .X(_0626_));
 sg13g2_buf_1 _6691_ (.A(_2136_),
    .X(_2139_));
 sg13g2_mux2_1 _6692_ (.A0(\logix.ram_r[1559] ),
    .A1(\logix.ram_r[1558] ),
    .S(net364),
    .X(_0627_));
 sg13g2_mux2_1 _6693_ (.A0(\logix.ram_r[155] ),
    .A1(\logix.ram_r[154] ),
    .S(_2139_),
    .X(_0628_));
 sg13g2_mux2_1 _6694_ (.A0(\logix.ram_r[1560] ),
    .A1(\logix.ram_r[1559] ),
    .S(net364),
    .X(_0629_));
 sg13g2_mux2_1 _6695_ (.A0(\logix.ram_r[1561] ),
    .A1(\logix.ram_r[1560] ),
    .S(net364),
    .X(_0630_));
 sg13g2_mux2_1 _6696_ (.A0(\logix.ram_r[1562] ),
    .A1(\logix.ram_r[1561] ),
    .S(net364),
    .X(_0631_));
 sg13g2_mux2_1 _6697_ (.A0(\logix.ram_r[1563] ),
    .A1(\logix.ram_r[1562] ),
    .S(net364),
    .X(_0632_));
 sg13g2_mux2_1 _6698_ (.A0(\logix.ram_r[1564] ),
    .A1(\logix.ram_r[1563] ),
    .S(_2139_),
    .X(_0633_));
 sg13g2_mux2_1 _6699_ (.A0(\logix.ram_r[1565] ),
    .A1(\logix.ram_r[1564] ),
    .S(net364),
    .X(_0634_));
 sg13g2_mux2_1 _6700_ (.A0(\logix.ram_r[1566] ),
    .A1(\logix.ram_r[1565] ),
    .S(net364),
    .X(_0635_));
 sg13g2_mux2_1 _6701_ (.A0(\logix.ram_r[1567] ),
    .A1(\logix.ram_r[1566] ),
    .S(net364),
    .X(_0636_));
 sg13g2_buf_1 _6702_ (.A(_2136_),
    .X(_2140_));
 sg13g2_mux2_1 _6703_ (.A0(\logix.ram_r[1568] ),
    .A1(\logix.ram_r[1567] ),
    .S(net363),
    .X(_0637_));
 sg13g2_mux2_1 _6704_ (.A0(\logix.ram_r[1569] ),
    .A1(\logix.ram_r[1568] ),
    .S(net363),
    .X(_0638_));
 sg13g2_mux2_1 _6705_ (.A0(\logix.ram_r[156] ),
    .A1(\logix.ram_r[155] ),
    .S(_2140_),
    .X(_0639_));
 sg13g2_mux2_1 _6706_ (.A0(\logix.ram_r[1570] ),
    .A1(\logix.ram_r[1569] ),
    .S(net363),
    .X(_0640_));
 sg13g2_mux2_1 _6707_ (.A0(\logix.ram_r[1571] ),
    .A1(\logix.ram_r[1570] ),
    .S(net363),
    .X(_0641_));
 sg13g2_mux2_1 _6708_ (.A0(\logix.ram_r[1572] ),
    .A1(\logix.ram_r[1571] ),
    .S(net363),
    .X(_0642_));
 sg13g2_mux2_1 _6709_ (.A0(\logix.ram_r[1573] ),
    .A1(\logix.ram_r[1572] ),
    .S(net363),
    .X(_0643_));
 sg13g2_mux2_1 _6710_ (.A0(\logix.ram_r[1574] ),
    .A1(\logix.ram_r[1573] ),
    .S(_2140_),
    .X(_0644_));
 sg13g2_mux2_1 _6711_ (.A0(\logix.ram_r[1575] ),
    .A1(\logix.ram_r[1574] ),
    .S(net363),
    .X(_0645_));
 sg13g2_mux2_1 _6712_ (.A0(\logix.ram_r[1576] ),
    .A1(\logix.ram_r[1575] ),
    .S(net363),
    .X(_0646_));
 sg13g2_buf_1 _6713_ (.A(_2136_),
    .X(_2141_));
 sg13g2_mux2_1 _6714_ (.A0(\logix.ram_r[1577] ),
    .A1(\logix.ram_r[1576] ),
    .S(net362),
    .X(_0647_));
 sg13g2_mux2_1 _6715_ (.A0(\logix.ram_r[1578] ),
    .A1(\logix.ram_r[1577] ),
    .S(net362),
    .X(_0648_));
 sg13g2_mux2_1 _6716_ (.A0(\logix.ram_r[1579] ),
    .A1(\logix.ram_r[1578] ),
    .S(_2141_),
    .X(_0649_));
 sg13g2_mux2_1 _6717_ (.A0(\logix.ram_r[157] ),
    .A1(\logix.ram_r[156] ),
    .S(net362),
    .X(_0650_));
 sg13g2_mux2_1 _6718_ (.A0(\logix.ram_r[1580] ),
    .A1(\logix.ram_r[1579] ),
    .S(net362),
    .X(_0651_));
 sg13g2_mux2_1 _6719_ (.A0(\logix.ram_r[1581] ),
    .A1(\logix.ram_r[1580] ),
    .S(net362),
    .X(_0652_));
 sg13g2_mux2_1 _6720_ (.A0(\logix.ram_r[1582] ),
    .A1(\logix.ram_r[1581] ),
    .S(net362),
    .X(_0653_));
 sg13g2_mux2_1 _6721_ (.A0(\logix.ram_r[1583] ),
    .A1(\logix.ram_r[1582] ),
    .S(net362),
    .X(_0654_));
 sg13g2_mux2_1 _6722_ (.A0(\logix.ram_r[1584] ),
    .A1(\logix.ram_r[1583] ),
    .S(_2141_),
    .X(_0655_));
 sg13g2_mux2_1 _6723_ (.A0(\logix.ram_r[1585] ),
    .A1(\logix.ram_r[1584] ),
    .S(net362),
    .X(_0656_));
 sg13g2_buf_2 _6724_ (.A(_2136_),
    .X(_2142_));
 sg13g2_mux2_1 _6725_ (.A0(\logix.ram_r[1586] ),
    .A1(\logix.ram_r[1585] ),
    .S(net361),
    .X(_0657_));
 sg13g2_mux2_1 _6726_ (.A0(\logix.ram_r[1587] ),
    .A1(\logix.ram_r[1586] ),
    .S(net361),
    .X(_0658_));
 sg13g2_mux2_1 _6727_ (.A0(\logix.ram_r[1588] ),
    .A1(\logix.ram_r[1587] ),
    .S(net361),
    .X(_0659_));
 sg13g2_mux2_1 _6728_ (.A0(\logix.ram_r[1589] ),
    .A1(\logix.ram_r[1588] ),
    .S(net361),
    .X(_0660_));
 sg13g2_mux2_1 _6729_ (.A0(\logix.ram_r[158] ),
    .A1(\logix.ram_r[157] ),
    .S(net361),
    .X(_0661_));
 sg13g2_mux2_1 _6730_ (.A0(\logix.ram_r[1590] ),
    .A1(\logix.ram_r[1589] ),
    .S(net361),
    .X(_0662_));
 sg13g2_mux2_1 _6731_ (.A0(\logix.ram_r[1591] ),
    .A1(\logix.ram_r[1590] ),
    .S(net361),
    .X(_0663_));
 sg13g2_mux2_1 _6732_ (.A0(\logix.ram_r[1592] ),
    .A1(\logix.ram_r[1591] ),
    .S(net361),
    .X(_0664_));
 sg13g2_mux2_1 _6733_ (.A0(\logix.ram_r[1593] ),
    .A1(\logix.ram_r[1592] ),
    .S(_2142_),
    .X(_0665_));
 sg13g2_mux2_1 _6734_ (.A0(\logix.ram_r[1594] ),
    .A1(\logix.ram_r[1593] ),
    .S(_2142_),
    .X(_0666_));
 sg13g2_buf_2 _6735_ (.A(_2136_),
    .X(_2143_));
 sg13g2_mux2_1 _6736_ (.A0(\logix.ram_r[1595] ),
    .A1(\logix.ram_r[1594] ),
    .S(net360),
    .X(_0667_));
 sg13g2_mux2_1 _6737_ (.A0(\logix.ram_r[1596] ),
    .A1(\logix.ram_r[1595] ),
    .S(net360),
    .X(_0668_));
 sg13g2_mux2_1 _6738_ (.A0(\logix.ram_r[1597] ),
    .A1(\logix.ram_r[1596] ),
    .S(net360),
    .X(_0669_));
 sg13g2_mux2_1 _6739_ (.A0(\logix.ram_r[1598] ),
    .A1(\logix.ram_r[1597] ),
    .S(net360),
    .X(_0670_));
 sg13g2_mux2_1 _6740_ (.A0(\logix.ram_r[1599] ),
    .A1(\logix.ram_r[1598] ),
    .S(net360),
    .X(_0671_));
 sg13g2_mux2_1 _6741_ (.A0(\logix.ram_r[159] ),
    .A1(\logix.ram_r[158] ),
    .S(_2143_),
    .X(_0672_));
 sg13g2_mux2_1 _6742_ (.A0(\logix.ram_r[15] ),
    .A1(\logix.ram_r[14] ),
    .S(_2143_),
    .X(_0673_));
 sg13g2_mux2_1 _6743_ (.A0(\logix.ram_r[1600] ),
    .A1(\logix.ram_r[1599] ),
    .S(net360),
    .X(_0674_));
 sg13g2_mux2_1 _6744_ (.A0(\logix.ram_r[1601] ),
    .A1(\logix.ram_r[1600] ),
    .S(net360),
    .X(_0675_));
 sg13g2_mux2_1 _6745_ (.A0(\logix.ram_r[1602] ),
    .A1(\logix.ram_r[1601] ),
    .S(net360),
    .X(_0676_));
 sg13g2_buf_2 _6746_ (.A(_2063_),
    .X(_2144_));
 sg13g2_buf_1 _6747_ (.A(_2144_),
    .X(_2145_));
 sg13g2_buf_2 _6748_ (.A(_2145_),
    .X(_2146_));
 sg13g2_mux2_1 _6749_ (.A0(\logix.ram_r[1603] ),
    .A1(\logix.ram_r[1602] ),
    .S(net359),
    .X(_0677_));
 sg13g2_mux2_1 _6750_ (.A0(\logix.ram_r[1604] ),
    .A1(\logix.ram_r[1603] ),
    .S(net359),
    .X(_0678_));
 sg13g2_mux2_1 _6751_ (.A0(\logix.ram_r[1605] ),
    .A1(\logix.ram_r[1604] ),
    .S(net359),
    .X(_0679_));
 sg13g2_mux2_1 _6752_ (.A0(\logix.ram_r[1606] ),
    .A1(\logix.ram_r[1605] ),
    .S(net359),
    .X(_0680_));
 sg13g2_mux2_1 _6753_ (.A0(\logix.ram_r[1607] ),
    .A1(\logix.ram_r[1606] ),
    .S(net359),
    .X(_0681_));
 sg13g2_mux2_1 _6754_ (.A0(\logix.ram_r[1608] ),
    .A1(\logix.ram_r[1607] ),
    .S(_2146_),
    .X(_0682_));
 sg13g2_mux2_1 _6755_ (.A0(\logix.ram_r[1609] ),
    .A1(\logix.ram_r[1608] ),
    .S(net359),
    .X(_0683_));
 sg13g2_mux2_1 _6756_ (.A0(\logix.ram_r[160] ),
    .A1(\logix.ram_r[159] ),
    .S(net359),
    .X(_0684_));
 sg13g2_mux2_1 _6757_ (.A0(\logix.ram_r[1610] ),
    .A1(\logix.ram_r[1609] ),
    .S(_2146_),
    .X(_0685_));
 sg13g2_mux2_1 _6758_ (.A0(\logix.ram_r[1611] ),
    .A1(\logix.ram_r[1610] ),
    .S(net359),
    .X(_0686_));
 sg13g2_buf_1 _6759_ (.A(_2145_),
    .X(_2147_));
 sg13g2_mux2_1 _6760_ (.A0(\logix.ram_r[1612] ),
    .A1(\logix.ram_r[1611] ),
    .S(net358),
    .X(_0687_));
 sg13g2_mux2_1 _6761_ (.A0(\logix.ram_r[1613] ),
    .A1(\logix.ram_r[1612] ),
    .S(net358),
    .X(_0688_));
 sg13g2_mux2_1 _6762_ (.A0(\logix.ram_r[1614] ),
    .A1(\logix.ram_r[1613] ),
    .S(net358),
    .X(_0689_));
 sg13g2_mux2_1 _6763_ (.A0(\logix.ram_r[1615] ),
    .A1(\logix.ram_r[1614] ),
    .S(net358),
    .X(_0690_));
 sg13g2_mux2_1 _6764_ (.A0(\logix.ram_r[1616] ),
    .A1(\logix.ram_r[1615] ),
    .S(net358),
    .X(_0691_));
 sg13g2_mux2_1 _6765_ (.A0(\logix.ram_r[1617] ),
    .A1(\logix.ram_r[1616] ),
    .S(_2147_),
    .X(_0692_));
 sg13g2_mux2_1 _6766_ (.A0(\logix.ram_r[1618] ),
    .A1(\logix.ram_r[1617] ),
    .S(net358),
    .X(_0693_));
 sg13g2_mux2_1 _6767_ (.A0(\logix.ram_r[1619] ),
    .A1(\logix.ram_r[1618] ),
    .S(net358),
    .X(_0694_));
 sg13g2_mux2_1 _6768_ (.A0(\logix.ram_r[161] ),
    .A1(\logix.ram_r[160] ),
    .S(net358),
    .X(_0695_));
 sg13g2_mux2_1 _6769_ (.A0(\logix.ram_r[1620] ),
    .A1(\logix.ram_r[1619] ),
    .S(_2147_),
    .X(_0696_));
 sg13g2_buf_1 _6770_ (.A(_2145_),
    .X(_2148_));
 sg13g2_mux2_1 _6771_ (.A0(\logix.ram_r[1621] ),
    .A1(\logix.ram_r[1620] ),
    .S(net357),
    .X(_0697_));
 sg13g2_mux2_1 _6772_ (.A0(\logix.ram_r[1622] ),
    .A1(\logix.ram_r[1621] ),
    .S(net357),
    .X(_0698_));
 sg13g2_mux2_1 _6773_ (.A0(\logix.ram_r[1623] ),
    .A1(\logix.ram_r[1622] ),
    .S(net357),
    .X(_0699_));
 sg13g2_mux2_1 _6774_ (.A0(\logix.ram_r[1624] ),
    .A1(\logix.ram_r[1623] ),
    .S(_2148_),
    .X(_0700_));
 sg13g2_mux2_1 _6775_ (.A0(\logix.ram_r[1625] ),
    .A1(\logix.ram_r[1624] ),
    .S(net357),
    .X(_0701_));
 sg13g2_mux2_1 _6776_ (.A0(\logix.ram_r[1626] ),
    .A1(\logix.ram_r[1625] ),
    .S(net357),
    .X(_0702_));
 sg13g2_mux2_1 _6777_ (.A0(\logix.ram_r[1627] ),
    .A1(\logix.ram_r[1626] ),
    .S(_2148_),
    .X(_0703_));
 sg13g2_mux2_1 _6778_ (.A0(\logix.ram_r[1628] ),
    .A1(\logix.ram_r[1627] ),
    .S(net357),
    .X(_0704_));
 sg13g2_mux2_1 _6779_ (.A0(\logix.ram_r[1629] ),
    .A1(\logix.ram_r[1628] ),
    .S(net357),
    .X(_0705_));
 sg13g2_mux2_1 _6780_ (.A0(\logix.ram_r[162] ),
    .A1(\logix.ram_r[161] ),
    .S(net357),
    .X(_0706_));
 sg13g2_buf_1 _6781_ (.A(_2145_),
    .X(_2149_));
 sg13g2_mux2_1 _6782_ (.A0(\logix.ram_r[1630] ),
    .A1(\logix.ram_r[1629] ),
    .S(net356),
    .X(_0707_));
 sg13g2_mux2_1 _6783_ (.A0(\logix.ram_r[1631] ),
    .A1(\logix.ram_r[1630] ),
    .S(_2149_),
    .X(_0708_));
 sg13g2_mux2_1 _6784_ (.A0(\logix.ram_r[1632] ),
    .A1(\logix.ram_r[1631] ),
    .S(net356),
    .X(_0709_));
 sg13g2_mux2_1 _6785_ (.A0(\logix.ram_r[1633] ),
    .A1(\logix.ram_r[1632] ),
    .S(net356),
    .X(_0710_));
 sg13g2_mux2_1 _6786_ (.A0(\logix.ram_r[1634] ),
    .A1(\logix.ram_r[1633] ),
    .S(_2149_),
    .X(_0711_));
 sg13g2_mux2_1 _6787_ (.A0(\logix.ram_r[1635] ),
    .A1(\logix.ram_r[1634] ),
    .S(net356),
    .X(_0712_));
 sg13g2_mux2_1 _6788_ (.A0(\logix.ram_r[1636] ),
    .A1(\logix.ram_r[1635] ),
    .S(net356),
    .X(_0713_));
 sg13g2_mux2_1 _6789_ (.A0(\logix.ram_r[1637] ),
    .A1(\logix.ram_r[1636] ),
    .S(net356),
    .X(_0714_));
 sg13g2_mux2_1 _6790_ (.A0(\logix.ram_r[1638] ),
    .A1(\logix.ram_r[1637] ),
    .S(net356),
    .X(_0715_));
 sg13g2_mux2_1 _6791_ (.A0(\logix.ram_r[1639] ),
    .A1(\logix.ram_r[1638] ),
    .S(net356),
    .X(_0716_));
 sg13g2_buf_1 _6792_ (.A(_2145_),
    .X(_2150_));
 sg13g2_mux2_1 _6793_ (.A0(\logix.ram_r[163] ),
    .A1(\logix.ram_r[162] ),
    .S(net355),
    .X(_0717_));
 sg13g2_mux2_1 _6794_ (.A0(\logix.ram_r[1640] ),
    .A1(\logix.ram_r[1639] ),
    .S(net355),
    .X(_0718_));
 sg13g2_mux2_1 _6795_ (.A0(\logix.ram_r[1641] ),
    .A1(\logix.ram_r[1640] ),
    .S(_2150_),
    .X(_0719_));
 sg13g2_mux2_1 _6796_ (.A0(\logix.ram_r[1642] ),
    .A1(\logix.ram_r[1641] ),
    .S(_2150_),
    .X(_0720_));
 sg13g2_mux2_1 _6797_ (.A0(\logix.ram_r[1643] ),
    .A1(\logix.ram_r[1642] ),
    .S(net355),
    .X(_0721_));
 sg13g2_mux2_1 _6798_ (.A0(\logix.ram_r[1644] ),
    .A1(\logix.ram_r[1643] ),
    .S(net355),
    .X(_0722_));
 sg13g2_mux2_1 _6799_ (.A0(\logix.ram_r[1645] ),
    .A1(\logix.ram_r[1644] ),
    .S(net355),
    .X(_0723_));
 sg13g2_mux2_1 _6800_ (.A0(\logix.ram_r[1646] ),
    .A1(\logix.ram_r[1645] ),
    .S(net355),
    .X(_0724_));
 sg13g2_mux2_1 _6801_ (.A0(\logix.ram_r[1647] ),
    .A1(\logix.ram_r[1646] ),
    .S(net355),
    .X(_0725_));
 sg13g2_mux2_1 _6802_ (.A0(\logix.ram_r[1648] ),
    .A1(\logix.ram_r[1647] ),
    .S(net355),
    .X(_0726_));
 sg13g2_buf_1 _6803_ (.A(_2145_),
    .X(_2151_));
 sg13g2_mux2_1 _6804_ (.A0(\logix.ram_r[1649] ),
    .A1(\logix.ram_r[1648] ),
    .S(net354),
    .X(_0727_));
 sg13g2_mux2_1 _6805_ (.A0(\logix.ram_r[164] ),
    .A1(\logix.ram_r[163] ),
    .S(_2151_),
    .X(_0728_));
 sg13g2_mux2_1 _6806_ (.A0(\logix.ram_r[1650] ),
    .A1(\logix.ram_r[1649] ),
    .S(net354),
    .X(_0729_));
 sg13g2_mux2_1 _6807_ (.A0(\logix.ram_r[1651] ),
    .A1(\logix.ram_r[1650] ),
    .S(net354),
    .X(_0730_));
 sg13g2_mux2_1 _6808_ (.A0(\logix.ram_r[1652] ),
    .A1(\logix.ram_r[1651] ),
    .S(net354),
    .X(_0731_));
 sg13g2_mux2_1 _6809_ (.A0(\logix.ram_r[1653] ),
    .A1(\logix.ram_r[1652] ),
    .S(net354),
    .X(_0732_));
 sg13g2_mux2_1 _6810_ (.A0(\logix.ram_r[1654] ),
    .A1(\logix.ram_r[1653] ),
    .S(net354),
    .X(_0733_));
 sg13g2_mux2_1 _6811_ (.A0(\logix.ram_r[1655] ),
    .A1(\logix.ram_r[1654] ),
    .S(net354),
    .X(_0734_));
 sg13g2_mux2_1 _6812_ (.A0(\logix.ram_r[1656] ),
    .A1(\logix.ram_r[1655] ),
    .S(net354),
    .X(_0735_));
 sg13g2_mux2_1 _6813_ (.A0(\logix.ram_r[1657] ),
    .A1(\logix.ram_r[1656] ),
    .S(_2151_),
    .X(_0736_));
 sg13g2_buf_1 _6814_ (.A(_2145_),
    .X(_2152_));
 sg13g2_mux2_1 _6815_ (.A0(\logix.ram_r[1658] ),
    .A1(\logix.ram_r[1657] ),
    .S(net353),
    .X(_0737_));
 sg13g2_mux2_1 _6816_ (.A0(\logix.ram_r[1659] ),
    .A1(\logix.ram_r[1658] ),
    .S(net353),
    .X(_0738_));
 sg13g2_mux2_1 _6817_ (.A0(\logix.ram_r[165] ),
    .A1(\logix.ram_r[164] ),
    .S(net353),
    .X(_0739_));
 sg13g2_mux2_1 _6818_ (.A0(\logix.ram_r[1660] ),
    .A1(\logix.ram_r[1659] ),
    .S(net353),
    .X(_0740_));
 sg13g2_mux2_1 _6819_ (.A0(\logix.ram_r[1661] ),
    .A1(\logix.ram_r[1660] ),
    .S(net353),
    .X(_0741_));
 sg13g2_mux2_1 _6820_ (.A0(\logix.ram_r[1662] ),
    .A1(\logix.ram_r[1661] ),
    .S(net353),
    .X(_0742_));
 sg13g2_mux2_1 _6821_ (.A0(\logix.ram_r[1663] ),
    .A1(\logix.ram_r[1662] ),
    .S(net353),
    .X(_0743_));
 sg13g2_mux2_1 _6822_ (.A0(\logix.ram_r[1664] ),
    .A1(\logix.ram_r[1663] ),
    .S(_2152_),
    .X(_0744_));
 sg13g2_mux2_1 _6823_ (.A0(\logix.ram_r[1665] ),
    .A1(\logix.ram_r[1664] ),
    .S(_2152_),
    .X(_0745_));
 sg13g2_mux2_1 _6824_ (.A0(\logix.ram_r[1666] ),
    .A1(\logix.ram_r[1665] ),
    .S(net353),
    .X(_0746_));
 sg13g2_buf_1 _6825_ (.A(_2144_),
    .X(_2153_));
 sg13g2_buf_1 _6826_ (.A(_2153_),
    .X(_2154_));
 sg13g2_mux2_1 _6827_ (.A0(\logix.ram_r[1667] ),
    .A1(\logix.ram_r[1666] ),
    .S(net352),
    .X(_0747_));
 sg13g2_mux2_1 _6828_ (.A0(\logix.ram_r[1668] ),
    .A1(\logix.ram_r[1667] ),
    .S(net352),
    .X(_0748_));
 sg13g2_mux2_1 _6829_ (.A0(\logix.ram_r[1669] ),
    .A1(\logix.ram_r[1668] ),
    .S(net352),
    .X(_0749_));
 sg13g2_mux2_1 _6830_ (.A0(\logix.ram_r[166] ),
    .A1(\logix.ram_r[165] ),
    .S(net352),
    .X(_0750_));
 sg13g2_mux2_1 _6831_ (.A0(\logix.ram_r[1670] ),
    .A1(\logix.ram_r[1669] ),
    .S(net352),
    .X(_0751_));
 sg13g2_mux2_1 _6832_ (.A0(\logix.ram_r[1671] ),
    .A1(\logix.ram_r[1670] ),
    .S(net352),
    .X(_0752_));
 sg13g2_mux2_1 _6833_ (.A0(\logix.ram_r[1672] ),
    .A1(\logix.ram_r[1671] ),
    .S(net352),
    .X(_0753_));
 sg13g2_mux2_1 _6834_ (.A0(\logix.ram_r[1673] ),
    .A1(\logix.ram_r[1672] ),
    .S(_2154_),
    .X(_0754_));
 sg13g2_mux2_1 _6835_ (.A0(\logix.ram_r[1674] ),
    .A1(\logix.ram_r[1673] ),
    .S(_2154_),
    .X(_0755_));
 sg13g2_mux2_1 _6836_ (.A0(\logix.ram_r[1675] ),
    .A1(\logix.ram_r[1674] ),
    .S(net352),
    .X(_0756_));
 sg13g2_buf_1 _6837_ (.A(_2153_),
    .X(_2155_));
 sg13g2_mux2_1 _6838_ (.A0(\logix.ram_r[1676] ),
    .A1(\logix.ram_r[1675] ),
    .S(net351),
    .X(_0757_));
 sg13g2_mux2_1 _6839_ (.A0(\logix.ram_r[1677] ),
    .A1(\logix.ram_r[1676] ),
    .S(net351),
    .X(_0758_));
 sg13g2_mux2_1 _6840_ (.A0(\logix.ram_r[1678] ),
    .A1(\logix.ram_r[1677] ),
    .S(_2155_),
    .X(_0759_));
 sg13g2_mux2_1 _6841_ (.A0(\logix.ram_r[1679] ),
    .A1(\logix.ram_r[1678] ),
    .S(net351),
    .X(_0760_));
 sg13g2_mux2_1 _6842_ (.A0(\logix.ram_r[167] ),
    .A1(\logix.ram_r[166] ),
    .S(net351),
    .X(_0761_));
 sg13g2_mux2_1 _6843_ (.A0(\logix.ram_r[1680] ),
    .A1(\logix.ram_r[1679] ),
    .S(net351),
    .X(_0762_));
 sg13g2_mux2_1 _6844_ (.A0(\logix.ram_r[1681] ),
    .A1(\logix.ram_r[1680] ),
    .S(net351),
    .X(_0763_));
 sg13g2_mux2_1 _6845_ (.A0(\logix.ram_r[1682] ),
    .A1(\logix.ram_r[1681] ),
    .S(net351),
    .X(_0764_));
 sg13g2_mux2_1 _6846_ (.A0(\logix.ram_r[1683] ),
    .A1(\logix.ram_r[1682] ),
    .S(net351),
    .X(_0765_));
 sg13g2_mux2_1 _6847_ (.A0(\logix.ram_r[1684] ),
    .A1(\logix.ram_r[1683] ),
    .S(_2155_),
    .X(_0766_));
 sg13g2_buf_1 _6848_ (.A(_2153_),
    .X(_2156_));
 sg13g2_mux2_1 _6849_ (.A0(\logix.ram_r[1685] ),
    .A1(\logix.ram_r[1684] ),
    .S(net350),
    .X(_0767_));
 sg13g2_mux2_1 _6850_ (.A0(\logix.ram_r[1686] ),
    .A1(\logix.ram_r[1685] ),
    .S(_2156_),
    .X(_0768_));
 sg13g2_mux2_1 _6851_ (.A0(\logix.ram_r[1687] ),
    .A1(\logix.ram_r[1686] ),
    .S(net350),
    .X(_0769_));
 sg13g2_mux2_1 _6852_ (.A0(\logix.ram_r[1688] ),
    .A1(\logix.ram_r[1687] ),
    .S(net350),
    .X(_0770_));
 sg13g2_mux2_1 _6853_ (.A0(\logix.ram_r[1689] ),
    .A1(\logix.ram_r[1688] ),
    .S(net350),
    .X(_0771_));
 sg13g2_mux2_1 _6854_ (.A0(\logix.ram_r[168] ),
    .A1(\logix.ram_r[167] ),
    .S(net350),
    .X(_0772_));
 sg13g2_mux2_1 _6855_ (.A0(\logix.ram_r[1690] ),
    .A1(\logix.ram_r[1689] ),
    .S(_2156_),
    .X(_0773_));
 sg13g2_mux2_1 _6856_ (.A0(\logix.ram_r[1691] ),
    .A1(\logix.ram_r[1690] ),
    .S(net350),
    .X(_0774_));
 sg13g2_mux2_1 _6857_ (.A0(\logix.ram_r[1692] ),
    .A1(\logix.ram_r[1691] ),
    .S(net350),
    .X(_0775_));
 sg13g2_mux2_1 _6858_ (.A0(\logix.ram_r[1693] ),
    .A1(\logix.ram_r[1692] ),
    .S(net350),
    .X(_0776_));
 sg13g2_buf_1 _6859_ (.A(_2153_),
    .X(_2157_));
 sg13g2_mux2_1 _6860_ (.A0(\logix.ram_r[1694] ),
    .A1(\logix.ram_r[1693] ),
    .S(_2157_),
    .X(_0777_));
 sg13g2_mux2_1 _6861_ (.A0(\logix.ram_r[1695] ),
    .A1(\logix.ram_r[1694] ),
    .S(net349),
    .X(_0778_));
 sg13g2_mux2_1 _6862_ (.A0(\logix.ram_r[1696] ),
    .A1(\logix.ram_r[1695] ),
    .S(net349),
    .X(_0779_));
 sg13g2_mux2_1 _6863_ (.A0(\logix.ram_r[1697] ),
    .A1(\logix.ram_r[1696] ),
    .S(net349),
    .X(_0780_));
 sg13g2_mux2_1 _6864_ (.A0(\logix.ram_r[1698] ),
    .A1(\logix.ram_r[1697] ),
    .S(net349),
    .X(_0781_));
 sg13g2_mux2_1 _6865_ (.A0(\logix.ram_r[1699] ),
    .A1(\logix.ram_r[1698] ),
    .S(net349),
    .X(_0782_));
 sg13g2_mux2_1 _6866_ (.A0(\logix.ram_r[169] ),
    .A1(\logix.ram_r[168] ),
    .S(net349),
    .X(_0783_));
 sg13g2_mux2_1 _6867_ (.A0(\logix.ram_r[16] ),
    .A1(\logix.ram_r[15] ),
    .S(_2157_),
    .X(_0784_));
 sg13g2_mux2_1 _6868_ (.A0(\logix.ram_r[1700] ),
    .A1(\logix.ram_r[1699] ),
    .S(net349),
    .X(_0785_));
 sg13g2_mux2_1 _6869_ (.A0(\logix.ram_r[1701] ),
    .A1(\logix.ram_r[1700] ),
    .S(net349),
    .X(_0786_));
 sg13g2_buf_1 _6870_ (.A(_2153_),
    .X(_2158_));
 sg13g2_mux2_1 _6871_ (.A0(\logix.ram_r[1702] ),
    .A1(\logix.ram_r[1701] ),
    .S(net348),
    .X(_0787_));
 sg13g2_mux2_1 _6872_ (.A0(\logix.ram_r[1703] ),
    .A1(\logix.ram_r[1702] ),
    .S(_2158_),
    .X(_0788_));
 sg13g2_mux2_1 _6873_ (.A0(\logix.ram_r[1704] ),
    .A1(\logix.ram_r[1703] ),
    .S(net348),
    .X(_0789_));
 sg13g2_mux2_1 _6874_ (.A0(\logix.ram_r[1705] ),
    .A1(\logix.ram_r[1704] ),
    .S(_2158_),
    .X(_0790_));
 sg13g2_mux2_1 _6875_ (.A0(\logix.ram_r[1706] ),
    .A1(\logix.ram_r[1705] ),
    .S(net348),
    .X(_0791_));
 sg13g2_mux2_1 _6876_ (.A0(\logix.ram_r[1707] ),
    .A1(\logix.ram_r[1706] ),
    .S(net348),
    .X(_0792_));
 sg13g2_mux2_1 _6877_ (.A0(\logix.ram_r[1708] ),
    .A1(\logix.ram_r[1707] ),
    .S(net348),
    .X(_0793_));
 sg13g2_mux2_1 _6878_ (.A0(\logix.ram_r[1709] ),
    .A1(\logix.ram_r[1708] ),
    .S(net348),
    .X(_0794_));
 sg13g2_mux2_1 _6879_ (.A0(\logix.ram_r[170] ),
    .A1(\logix.ram_r[169] ),
    .S(net348),
    .X(_0795_));
 sg13g2_mux2_1 _6880_ (.A0(\logix.ram_r[1710] ),
    .A1(\logix.ram_r[1709] ),
    .S(net348),
    .X(_0796_));
 sg13g2_buf_1 _6881_ (.A(_2153_),
    .X(_2159_));
 sg13g2_mux2_1 _6882_ (.A0(\logix.ram_r[1711] ),
    .A1(\logix.ram_r[1710] ),
    .S(net347),
    .X(_0797_));
 sg13g2_mux2_1 _6883_ (.A0(\logix.ram_r[1712] ),
    .A1(\logix.ram_r[1711] ),
    .S(net347),
    .X(_0798_));
 sg13g2_mux2_1 _6884_ (.A0(\logix.ram_r[1713] ),
    .A1(\logix.ram_r[1712] ),
    .S(net347),
    .X(_0799_));
 sg13g2_mux2_1 _6885_ (.A0(\logix.ram_r[1714] ),
    .A1(\logix.ram_r[1713] ),
    .S(_2159_),
    .X(_0800_));
 sg13g2_mux2_1 _6886_ (.A0(\logix.ram_r[1715] ),
    .A1(\logix.ram_r[1714] ),
    .S(net347),
    .X(_0801_));
 sg13g2_mux2_1 _6887_ (.A0(\logix.ram_r[1716] ),
    .A1(\logix.ram_r[1715] ),
    .S(net347),
    .X(_0802_));
 sg13g2_mux2_1 _6888_ (.A0(\logix.ram_r[1717] ),
    .A1(\logix.ram_r[1716] ),
    .S(net347),
    .X(_0803_));
 sg13g2_mux2_1 _6889_ (.A0(\logix.ram_r[1718] ),
    .A1(\logix.ram_r[1717] ),
    .S(net347),
    .X(_0804_));
 sg13g2_mux2_1 _6890_ (.A0(\logix.ram_r[1719] ),
    .A1(\logix.ram_r[1718] ),
    .S(net347),
    .X(_0805_));
 sg13g2_mux2_1 _6891_ (.A0(\logix.ram_r[171] ),
    .A1(\logix.ram_r[170] ),
    .S(_2159_),
    .X(_0806_));
 sg13g2_buf_1 _6892_ (.A(_2153_),
    .X(_2160_));
 sg13g2_mux2_1 _6893_ (.A0(\logix.ram_r[1720] ),
    .A1(\logix.ram_r[1719] ),
    .S(_2160_),
    .X(_0807_));
 sg13g2_mux2_1 _6894_ (.A0(\logix.ram_r[1721] ),
    .A1(\logix.ram_r[1720] ),
    .S(net346),
    .X(_0808_));
 sg13g2_mux2_1 _6895_ (.A0(\logix.ram_r[1722] ),
    .A1(\logix.ram_r[1721] ),
    .S(_2160_),
    .X(_0809_));
 sg13g2_mux2_1 _6896_ (.A0(\logix.ram_r[1723] ),
    .A1(\logix.ram_r[1722] ),
    .S(net346),
    .X(_0810_));
 sg13g2_mux2_1 _6897_ (.A0(\logix.ram_r[1724] ),
    .A1(\logix.ram_r[1723] ),
    .S(net346),
    .X(_0811_));
 sg13g2_mux2_1 _6898_ (.A0(\logix.ram_r[1725] ),
    .A1(\logix.ram_r[1724] ),
    .S(net346),
    .X(_0812_));
 sg13g2_mux2_1 _6899_ (.A0(\logix.ram_r[1726] ),
    .A1(\logix.ram_r[1725] ),
    .S(net346),
    .X(_0813_));
 sg13g2_mux2_1 _6900_ (.A0(\logix.ram_r[1727] ),
    .A1(\logix.ram_r[1726] ),
    .S(net346),
    .X(_0814_));
 sg13g2_mux2_1 _6901_ (.A0(\logix.ram_r[1728] ),
    .A1(\logix.ram_r[1727] ),
    .S(net346),
    .X(_0815_));
 sg13g2_mux2_1 _6902_ (.A0(\logix.ram_r[1729] ),
    .A1(\logix.ram_r[1728] ),
    .S(net346),
    .X(_0816_));
 sg13g2_buf_1 _6903_ (.A(_2144_),
    .X(_2161_));
 sg13g2_buf_1 _6904_ (.A(_2161_),
    .X(_2162_));
 sg13g2_mux2_1 _6905_ (.A0(\logix.ram_r[172] ),
    .A1(\logix.ram_r[171] ),
    .S(net345),
    .X(_0817_));
 sg13g2_mux2_1 _6906_ (.A0(\logix.ram_r[1730] ),
    .A1(\logix.ram_r[1729] ),
    .S(net345),
    .X(_0818_));
 sg13g2_mux2_1 _6907_ (.A0(\logix.ram_r[1731] ),
    .A1(\logix.ram_r[1730] ),
    .S(net345),
    .X(_0819_));
 sg13g2_mux2_1 _6908_ (.A0(\logix.ram_r[1732] ),
    .A1(\logix.ram_r[1731] ),
    .S(net345),
    .X(_0820_));
 sg13g2_mux2_1 _6909_ (.A0(\logix.ram_r[1733] ),
    .A1(\logix.ram_r[1732] ),
    .S(net345),
    .X(_0821_));
 sg13g2_mux2_1 _6910_ (.A0(\logix.ram_r[1734] ),
    .A1(\logix.ram_r[1733] ),
    .S(net345),
    .X(_0822_));
 sg13g2_mux2_1 _6911_ (.A0(\logix.ram_r[1735] ),
    .A1(\logix.ram_r[1734] ),
    .S(_2162_),
    .X(_0823_));
 sg13g2_mux2_1 _6912_ (.A0(\logix.ram_r[1736] ),
    .A1(\logix.ram_r[1735] ),
    .S(net345),
    .X(_0824_));
 sg13g2_mux2_1 _6913_ (.A0(\logix.ram_r[1737] ),
    .A1(\logix.ram_r[1736] ),
    .S(net345),
    .X(_0825_));
 sg13g2_mux2_1 _6914_ (.A0(\logix.ram_r[1738] ),
    .A1(\logix.ram_r[1737] ),
    .S(_2162_),
    .X(_0826_));
 sg13g2_buf_1 _6915_ (.A(_2161_),
    .X(_2163_));
 sg13g2_mux2_1 _6916_ (.A0(\logix.ram_r[1739] ),
    .A1(\logix.ram_r[1738] ),
    .S(_2163_),
    .X(_0827_));
 sg13g2_mux2_1 _6917_ (.A0(\logix.ram_r[173] ),
    .A1(\logix.ram_r[172] ),
    .S(net344),
    .X(_0828_));
 sg13g2_mux2_1 _6918_ (.A0(\logix.ram_r[1740] ),
    .A1(\logix.ram_r[1739] ),
    .S(net344),
    .X(_0829_));
 sg13g2_mux2_1 _6919_ (.A0(\logix.ram_r[1741] ),
    .A1(\logix.ram_r[1740] ),
    .S(net344),
    .X(_0830_));
 sg13g2_mux2_1 _6920_ (.A0(\logix.ram_r[1742] ),
    .A1(\logix.ram_r[1741] ),
    .S(net344),
    .X(_0831_));
 sg13g2_mux2_1 _6921_ (.A0(\logix.ram_r[1743] ),
    .A1(\logix.ram_r[1742] ),
    .S(net344),
    .X(_0832_));
 sg13g2_mux2_1 _6922_ (.A0(\logix.ram_r[1744] ),
    .A1(\logix.ram_r[1743] ),
    .S(net344),
    .X(_0833_));
 sg13g2_mux2_1 _6923_ (.A0(\logix.ram_r[1745] ),
    .A1(\logix.ram_r[1744] ),
    .S(net344),
    .X(_0834_));
 sg13g2_mux2_1 _6924_ (.A0(\logix.ram_r[1746] ),
    .A1(\logix.ram_r[1745] ),
    .S(net344),
    .X(_0835_));
 sg13g2_mux2_1 _6925_ (.A0(\logix.ram_r[1747] ),
    .A1(\logix.ram_r[1746] ),
    .S(_2163_),
    .X(_0836_));
 sg13g2_buf_1 _6926_ (.A(_2161_),
    .X(_2164_));
 sg13g2_mux2_1 _6927_ (.A0(\logix.ram_r[1748] ),
    .A1(\logix.ram_r[1747] ),
    .S(net343),
    .X(_0837_));
 sg13g2_mux2_1 _6928_ (.A0(\logix.ram_r[1749] ),
    .A1(\logix.ram_r[1748] ),
    .S(net343),
    .X(_0838_));
 sg13g2_mux2_1 _6929_ (.A0(\logix.ram_r[174] ),
    .A1(\logix.ram_r[173] ),
    .S(net343),
    .X(_0839_));
 sg13g2_mux2_1 _6930_ (.A0(\logix.ram_r[1750] ),
    .A1(\logix.ram_r[1749] ),
    .S(net343),
    .X(_0840_));
 sg13g2_mux2_1 _6931_ (.A0(\logix.ram_r[1751] ),
    .A1(\logix.ram_r[1750] ),
    .S(_2164_),
    .X(_0841_));
 sg13g2_mux2_1 _6932_ (.A0(\logix.ram_r[1752] ),
    .A1(\logix.ram_r[1751] ),
    .S(net343),
    .X(_0842_));
 sg13g2_mux2_1 _6933_ (.A0(\logix.ram_r[1753] ),
    .A1(\logix.ram_r[1752] ),
    .S(_2164_),
    .X(_0843_));
 sg13g2_mux2_1 _6934_ (.A0(\logix.ram_r[1754] ),
    .A1(\logix.ram_r[1753] ),
    .S(net343),
    .X(_0844_));
 sg13g2_mux2_1 _6935_ (.A0(\logix.ram_r[1755] ),
    .A1(\logix.ram_r[1754] ),
    .S(net343),
    .X(_0845_));
 sg13g2_mux2_1 _6936_ (.A0(\logix.ram_r[1756] ),
    .A1(\logix.ram_r[1755] ),
    .S(net343),
    .X(_0846_));
 sg13g2_buf_1 _6937_ (.A(_2161_),
    .X(_2165_));
 sg13g2_mux2_1 _6938_ (.A0(\logix.ram_r[1757] ),
    .A1(\logix.ram_r[1756] ),
    .S(_2165_),
    .X(_0847_));
 sg13g2_mux2_1 _6939_ (.A0(\logix.ram_r[1758] ),
    .A1(\logix.ram_r[1757] ),
    .S(net342),
    .X(_0848_));
 sg13g2_mux2_1 _6940_ (.A0(\logix.ram_r[1759] ),
    .A1(\logix.ram_r[1758] ),
    .S(net342),
    .X(_0849_));
 sg13g2_mux2_1 _6941_ (.A0(\logix.ram_r[175] ),
    .A1(\logix.ram_r[174] ),
    .S(_2165_),
    .X(_0850_));
 sg13g2_mux2_1 _6942_ (.A0(\logix.ram_r[1760] ),
    .A1(\logix.ram_r[1759] ),
    .S(net342),
    .X(_0851_));
 sg13g2_mux2_1 _6943_ (.A0(\logix.ram_r[1761] ),
    .A1(\logix.ram_r[1760] ),
    .S(net342),
    .X(_0852_));
 sg13g2_mux2_1 _6944_ (.A0(\logix.ram_r[1762] ),
    .A1(\logix.ram_r[1761] ),
    .S(net342),
    .X(_0853_));
 sg13g2_mux2_1 _6945_ (.A0(\logix.ram_r[1763] ),
    .A1(\logix.ram_r[1762] ),
    .S(net342),
    .X(_0854_));
 sg13g2_mux2_1 _6946_ (.A0(\logix.ram_r[1764] ),
    .A1(\logix.ram_r[1763] ),
    .S(net342),
    .X(_0855_));
 sg13g2_mux2_1 _6947_ (.A0(\logix.ram_r[1765] ),
    .A1(\logix.ram_r[1764] ),
    .S(net342),
    .X(_0856_));
 sg13g2_buf_1 _6948_ (.A(_2161_),
    .X(_2166_));
 sg13g2_mux2_1 _6949_ (.A0(\logix.ram_r[1766] ),
    .A1(\logix.ram_r[1765] ),
    .S(net341),
    .X(_0857_));
 sg13g2_mux2_1 _6950_ (.A0(\logix.ram_r[1767] ),
    .A1(\logix.ram_r[1766] ),
    .S(net341),
    .X(_0858_));
 sg13g2_mux2_1 _6951_ (.A0(\logix.ram_r[1768] ),
    .A1(\logix.ram_r[1767] ),
    .S(_2166_),
    .X(_0859_));
 sg13g2_mux2_1 _6952_ (.A0(\logix.ram_r[1769] ),
    .A1(\logix.ram_r[1768] ),
    .S(net341),
    .X(_0860_));
 sg13g2_mux2_1 _6953_ (.A0(\logix.ram_r[176] ),
    .A1(\logix.ram_r[175] ),
    .S(_2166_),
    .X(_0861_));
 sg13g2_mux2_1 _6954_ (.A0(\logix.ram_r[1770] ),
    .A1(\logix.ram_r[1769] ),
    .S(net341),
    .X(_0862_));
 sg13g2_mux2_1 _6955_ (.A0(\logix.ram_r[1771] ),
    .A1(\logix.ram_r[1770] ),
    .S(net341),
    .X(_0863_));
 sg13g2_mux2_1 _6956_ (.A0(\logix.ram_r[1772] ),
    .A1(\logix.ram_r[1771] ),
    .S(net341),
    .X(_0864_));
 sg13g2_mux2_1 _6957_ (.A0(\logix.ram_r[1773] ),
    .A1(\logix.ram_r[1772] ),
    .S(net341),
    .X(_0865_));
 sg13g2_mux2_1 _6958_ (.A0(\logix.ram_r[1774] ),
    .A1(\logix.ram_r[1773] ),
    .S(net341),
    .X(_0866_));
 sg13g2_buf_1 _6959_ (.A(_2161_),
    .X(_2167_));
 sg13g2_mux2_1 _6960_ (.A0(\logix.ram_r[1775] ),
    .A1(\logix.ram_r[1774] ),
    .S(net340),
    .X(_0867_));
 sg13g2_mux2_1 _6961_ (.A0(\logix.ram_r[1776] ),
    .A1(\logix.ram_r[1775] ),
    .S(net340),
    .X(_0868_));
 sg13g2_mux2_1 _6962_ (.A0(\logix.ram_r[1777] ),
    .A1(\logix.ram_r[1776] ),
    .S(net340),
    .X(_0869_));
 sg13g2_mux2_1 _6963_ (.A0(\logix.ram_r[1778] ),
    .A1(\logix.ram_r[1777] ),
    .S(net340),
    .X(_0870_));
 sg13g2_mux2_1 _6964_ (.A0(\logix.ram_r[1779] ),
    .A1(\logix.ram_r[1778] ),
    .S(net340),
    .X(_0871_));
 sg13g2_mux2_1 _6965_ (.A0(\logix.ram_r[177] ),
    .A1(\logix.ram_r[176] ),
    .S(_2167_),
    .X(_0872_));
 sg13g2_mux2_1 _6966_ (.A0(\logix.ram_r[1780] ),
    .A1(\logix.ram_r[1779] ),
    .S(net340),
    .X(_0873_));
 sg13g2_mux2_1 _6967_ (.A0(\logix.ram_r[1781] ),
    .A1(\logix.ram_r[1780] ),
    .S(net340),
    .X(_0874_));
 sg13g2_mux2_1 _6968_ (.A0(\logix.ram_r[1782] ),
    .A1(\logix.ram_r[1781] ),
    .S(net340),
    .X(_0875_));
 sg13g2_mux2_1 _6969_ (.A0(\logix.ram_r[1783] ),
    .A1(\logix.ram_r[1782] ),
    .S(_2167_),
    .X(_0876_));
 sg13g2_buf_1 _6970_ (.A(_2161_),
    .X(_2168_));
 sg13g2_mux2_1 _6971_ (.A0(\logix.ram_r[1784] ),
    .A1(\logix.ram_r[1783] ),
    .S(net339),
    .X(_0877_));
 sg13g2_mux2_1 _6972_ (.A0(\logix.ram_r[1785] ),
    .A1(\logix.ram_r[1784] ),
    .S(net339),
    .X(_0878_));
 sg13g2_mux2_1 _6973_ (.A0(\logix.ram_r[1786] ),
    .A1(\logix.ram_r[1785] ),
    .S(net339),
    .X(_0879_));
 sg13g2_mux2_1 _6974_ (.A0(\logix.ram_r[1787] ),
    .A1(\logix.ram_r[1786] ),
    .S(net339),
    .X(_0880_));
 sg13g2_mux2_1 _6975_ (.A0(\logix.ram_r[1788] ),
    .A1(\logix.ram_r[1787] ),
    .S(net339),
    .X(_0881_));
 sg13g2_mux2_1 _6976_ (.A0(\logix.ram_r[1789] ),
    .A1(\logix.ram_r[1788] ),
    .S(net339),
    .X(_0882_));
 sg13g2_mux2_1 _6977_ (.A0(\logix.ram_r[178] ),
    .A1(\logix.ram_r[177] ),
    .S(_2168_),
    .X(_0883_));
 sg13g2_mux2_1 _6978_ (.A0(\logix.ram_r[1790] ),
    .A1(\logix.ram_r[1789] ),
    .S(net339),
    .X(_0884_));
 sg13g2_mux2_1 _6979_ (.A0(\logix.ram_r[1791] ),
    .A1(\logix.ram_r[1790] ),
    .S(_2168_),
    .X(_0885_));
 sg13g2_mux2_1 _6980_ (.A0(\logix.ram_r[1792] ),
    .A1(\logix.ram_r[1791] ),
    .S(net339),
    .X(_0886_));
 sg13g2_buf_1 _6981_ (.A(_2144_),
    .X(_2169_));
 sg13g2_buf_1 _6982_ (.A(_2169_),
    .X(_2170_));
 sg13g2_mux2_1 _6983_ (.A0(\logix.ram_r[1793] ),
    .A1(\logix.ram_r[1792] ),
    .S(net338),
    .X(_0887_));
 sg13g2_mux2_1 _6984_ (.A0(\logix.ram_r[1794] ),
    .A1(\logix.ram_r[1793] ),
    .S(net338),
    .X(_0888_));
 sg13g2_mux2_1 _6985_ (.A0(\logix.ram_r[1795] ),
    .A1(\logix.ram_r[1794] ),
    .S(net338),
    .X(_0889_));
 sg13g2_mux2_1 _6986_ (.A0(\logix.ram_r[1796] ),
    .A1(\logix.ram_r[1795] ),
    .S(net338),
    .X(_0890_));
 sg13g2_mux2_1 _6987_ (.A0(\logix.ram_r[1797] ),
    .A1(\logix.ram_r[1796] ),
    .S(net338),
    .X(_0891_));
 sg13g2_mux2_1 _6988_ (.A0(\logix.ram_r[1798] ),
    .A1(\logix.ram_r[1797] ),
    .S(net338),
    .X(_0892_));
 sg13g2_mux2_1 _6989_ (.A0(\logix.ram_r[1799] ),
    .A1(\logix.ram_r[1798] ),
    .S(net338),
    .X(_0893_));
 sg13g2_mux2_1 _6990_ (.A0(\logix.ram_r[179] ),
    .A1(\logix.ram_r[178] ),
    .S(_2170_),
    .X(_0894_));
 sg13g2_mux2_1 _6991_ (.A0(\logix.ram_r[17] ),
    .A1(\logix.ram_r[16] ),
    .S(_2170_),
    .X(_0895_));
 sg13g2_mux2_1 _6992_ (.A0(\logix.ram_r[1800] ),
    .A1(\logix.ram_r[1799] ),
    .S(net338),
    .X(_0896_));
 sg13g2_buf_2 _6993_ (.A(_2169_),
    .X(_2171_));
 sg13g2_mux2_1 _6994_ (.A0(\logix.ram_r[1801] ),
    .A1(\logix.ram_r[1800] ),
    .S(net337),
    .X(_0897_));
 sg13g2_mux2_1 _6995_ (.A0(\logix.ram_r[1802] ),
    .A1(\logix.ram_r[1801] ),
    .S(net337),
    .X(_0898_));
 sg13g2_mux2_1 _6996_ (.A0(\logix.ram_r[1803] ),
    .A1(\logix.ram_r[1802] ),
    .S(net337),
    .X(_0899_));
 sg13g2_mux2_1 _6997_ (.A0(\logix.ram_r[1804] ),
    .A1(\logix.ram_r[1803] ),
    .S(net337),
    .X(_0900_));
 sg13g2_mux2_1 _6998_ (.A0(\logix.ram_r[1805] ),
    .A1(\logix.ram_r[1804] ),
    .S(_2171_),
    .X(_0901_));
 sg13g2_mux2_1 _6999_ (.A0(\logix.ram_r[1806] ),
    .A1(\logix.ram_r[1805] ),
    .S(net337),
    .X(_0902_));
 sg13g2_mux2_1 _7000_ (.A0(\logix.ram_r[1807] ),
    .A1(\logix.ram_r[1806] ),
    .S(net337),
    .X(_0903_));
 sg13g2_mux2_1 _7001_ (.A0(\logix.ram_r[1808] ),
    .A1(\logix.ram_r[1807] ),
    .S(net337),
    .X(_0904_));
 sg13g2_mux2_1 _7002_ (.A0(\logix.ram_r[1809] ),
    .A1(\logix.ram_r[1808] ),
    .S(net337),
    .X(_0905_));
 sg13g2_mux2_1 _7003_ (.A0(\logix.ram_r[180] ),
    .A1(\logix.ram_r[179] ),
    .S(_2171_),
    .X(_0906_));
 sg13g2_buf_1 _7004_ (.A(_2169_),
    .X(_2172_));
 sg13g2_mux2_1 _7005_ (.A0(\logix.ram_r[1810] ),
    .A1(\logix.ram_r[1809] ),
    .S(_2172_),
    .X(_0907_));
 sg13g2_mux2_1 _7006_ (.A0(\logix.ram_r[1811] ),
    .A1(\logix.ram_r[1810] ),
    .S(net336),
    .X(_0908_));
 sg13g2_mux2_1 _7007_ (.A0(\logix.ram_r[1812] ),
    .A1(\logix.ram_r[1811] ),
    .S(net336),
    .X(_0909_));
 sg13g2_mux2_1 _7008_ (.A0(\logix.ram_r[1813] ),
    .A1(\logix.ram_r[1812] ),
    .S(net336),
    .X(_0910_));
 sg13g2_mux2_1 _7009_ (.A0(\logix.ram_r[1814] ),
    .A1(\logix.ram_r[1813] ),
    .S(_2172_),
    .X(_0911_));
 sg13g2_mux2_1 _7010_ (.A0(\logix.ram_r[1815] ),
    .A1(\logix.ram_r[1814] ),
    .S(net336),
    .X(_0912_));
 sg13g2_mux2_1 _7011_ (.A0(\logix.ram_r[1816] ),
    .A1(\logix.ram_r[1815] ),
    .S(net336),
    .X(_0913_));
 sg13g2_mux2_1 _7012_ (.A0(\logix.ram_r[1817] ),
    .A1(\logix.ram_r[1816] ),
    .S(net336),
    .X(_0914_));
 sg13g2_mux2_1 _7013_ (.A0(\logix.ram_r[1818] ),
    .A1(\logix.ram_r[1817] ),
    .S(net336),
    .X(_0915_));
 sg13g2_mux2_1 _7014_ (.A0(\logix.ram_r[1819] ),
    .A1(\logix.ram_r[1818] ),
    .S(net336),
    .X(_0916_));
 sg13g2_buf_1 _7015_ (.A(_2169_),
    .X(_2173_));
 sg13g2_mux2_1 _7016_ (.A0(\logix.ram_r[181] ),
    .A1(\logix.ram_r[180] ),
    .S(net335),
    .X(_0917_));
 sg13g2_mux2_1 _7017_ (.A0(\logix.ram_r[1820] ),
    .A1(\logix.ram_r[1819] ),
    .S(net335),
    .X(_0918_));
 sg13g2_mux2_1 _7018_ (.A0(\logix.ram_r[1821] ),
    .A1(\logix.ram_r[1820] ),
    .S(net335),
    .X(_0919_));
 sg13g2_mux2_1 _7019_ (.A0(\logix.ram_r[1822] ),
    .A1(\logix.ram_r[1821] ),
    .S(net335),
    .X(_0920_));
 sg13g2_mux2_1 _7020_ (.A0(\logix.ram_r[1823] ),
    .A1(\logix.ram_r[1822] ),
    .S(net335),
    .X(_0921_));
 sg13g2_mux2_1 _7021_ (.A0(\logix.ram_r[1824] ),
    .A1(\logix.ram_r[1823] ),
    .S(net335),
    .X(_0922_));
 sg13g2_mux2_1 _7022_ (.A0(\logix.ram_r[1825] ),
    .A1(\logix.ram_r[1824] ),
    .S(_2173_),
    .X(_0923_));
 sg13g2_mux2_1 _7023_ (.A0(\logix.ram_r[1826] ),
    .A1(\logix.ram_r[1825] ),
    .S(net335),
    .X(_0924_));
 sg13g2_mux2_1 _7024_ (.A0(\logix.ram_r[1827] ),
    .A1(\logix.ram_r[1826] ),
    .S(_2173_),
    .X(_0925_));
 sg13g2_mux2_1 _7025_ (.A0(\logix.ram_r[1828] ),
    .A1(\logix.ram_r[1827] ),
    .S(net335),
    .X(_0926_));
 sg13g2_buf_1 _7026_ (.A(_2169_),
    .X(_2174_));
 sg13g2_mux2_1 _7027_ (.A0(\logix.ram_r[1829] ),
    .A1(\logix.ram_r[1828] ),
    .S(_2174_),
    .X(_0927_));
 sg13g2_mux2_1 _7028_ (.A0(\logix.ram_r[182] ),
    .A1(\logix.ram_r[181] ),
    .S(net334),
    .X(_0928_));
 sg13g2_mux2_1 _7029_ (.A0(\logix.ram_r[1830] ),
    .A1(\logix.ram_r[1829] ),
    .S(net334),
    .X(_0929_));
 sg13g2_mux2_1 _7030_ (.A0(\logix.ram_r[1831] ),
    .A1(\logix.ram_r[1830] ),
    .S(net334),
    .X(_0930_));
 sg13g2_mux2_1 _7031_ (.A0(\logix.ram_r[1832] ),
    .A1(\logix.ram_r[1831] ),
    .S(net334),
    .X(_0931_));
 sg13g2_mux2_1 _7032_ (.A0(\logix.ram_r[1833] ),
    .A1(\logix.ram_r[1832] ),
    .S(net334),
    .X(_0932_));
 sg13g2_mux2_1 _7033_ (.A0(\logix.ram_r[1834] ),
    .A1(\logix.ram_r[1833] ),
    .S(net334),
    .X(_0933_));
 sg13g2_mux2_1 _7034_ (.A0(\logix.ram_r[1835] ),
    .A1(\logix.ram_r[1834] ),
    .S(net334),
    .X(_0934_));
 sg13g2_mux2_1 _7035_ (.A0(\logix.ram_r[1836] ),
    .A1(\logix.ram_r[1835] ),
    .S(net334),
    .X(_0935_));
 sg13g2_mux2_1 _7036_ (.A0(\logix.ram_r[1837] ),
    .A1(\logix.ram_r[1836] ),
    .S(_2174_),
    .X(_0936_));
 sg13g2_buf_1 _7037_ (.A(_2169_),
    .X(_2175_));
 sg13g2_mux2_1 _7038_ (.A0(\logix.ram_r[1838] ),
    .A1(\logix.ram_r[1837] ),
    .S(net333),
    .X(_0937_));
 sg13g2_mux2_1 _7039_ (.A0(\logix.ram_r[1839] ),
    .A1(\logix.ram_r[1838] ),
    .S(net333),
    .X(_0938_));
 sg13g2_mux2_1 _7040_ (.A0(\logix.ram_r[183] ),
    .A1(\logix.ram_r[182] ),
    .S(net333),
    .X(_0939_));
 sg13g2_mux2_1 _7041_ (.A0(\logix.ram_r[1840] ),
    .A1(\logix.ram_r[1839] ),
    .S(net333),
    .X(_0940_));
 sg13g2_mux2_1 _7042_ (.A0(\logix.ram_r[1841] ),
    .A1(\logix.ram_r[1840] ),
    .S(_2175_),
    .X(_0941_));
 sg13g2_mux2_1 _7043_ (.A0(\logix.ram_r[1842] ),
    .A1(\logix.ram_r[1841] ),
    .S(net333),
    .X(_0942_));
 sg13g2_mux2_1 _7044_ (.A0(\logix.ram_r[1843] ),
    .A1(\logix.ram_r[1842] ),
    .S(net333),
    .X(_0943_));
 sg13g2_mux2_1 _7045_ (.A0(\logix.ram_r[1844] ),
    .A1(\logix.ram_r[1843] ),
    .S(net333),
    .X(_0944_));
 sg13g2_mux2_1 _7046_ (.A0(\logix.ram_r[1845] ),
    .A1(\logix.ram_r[1844] ),
    .S(_2175_),
    .X(_0945_));
 sg13g2_mux2_1 _7047_ (.A0(\logix.ram_r[1846] ),
    .A1(\logix.ram_r[1845] ),
    .S(net333),
    .X(_0946_));
 sg13g2_buf_1 _7048_ (.A(_2169_),
    .X(_2176_));
 sg13g2_mux2_1 _7049_ (.A0(\logix.ram_r[1847] ),
    .A1(\logix.ram_r[1846] ),
    .S(net332),
    .X(_0947_));
 sg13g2_mux2_1 _7050_ (.A0(\logix.ram_r[1848] ),
    .A1(\logix.ram_r[1847] ),
    .S(net332),
    .X(_0948_));
 sg13g2_mux2_1 _7051_ (.A0(\logix.ram_r[1849] ),
    .A1(\logix.ram_r[1848] ),
    .S(net332),
    .X(_0949_));
 sg13g2_mux2_1 _7052_ (.A0(\logix.ram_r[184] ),
    .A1(\logix.ram_r[183] ),
    .S(net332),
    .X(_0950_));
 sg13g2_mux2_1 _7053_ (.A0(\logix.ram_r[1850] ),
    .A1(\logix.ram_r[1849] ),
    .S(net332),
    .X(_0951_));
 sg13g2_mux2_1 _7054_ (.A0(\logix.ram_r[1851] ),
    .A1(\logix.ram_r[1850] ),
    .S(_2176_),
    .X(_0952_));
 sg13g2_mux2_1 _7055_ (.A0(\logix.ram_r[1852] ),
    .A1(\logix.ram_r[1851] ),
    .S(_2176_),
    .X(_0953_));
 sg13g2_mux2_1 _7056_ (.A0(\logix.ram_r[1853] ),
    .A1(\logix.ram_r[1852] ),
    .S(net332),
    .X(_0954_));
 sg13g2_mux2_1 _7057_ (.A0(\logix.ram_r[1854] ),
    .A1(\logix.ram_r[1853] ),
    .S(net332),
    .X(_0955_));
 sg13g2_mux2_1 _7058_ (.A0(\logix.ram_r[1855] ),
    .A1(\logix.ram_r[1854] ),
    .S(net332),
    .X(_0956_));
 sg13g2_buf_1 _7059_ (.A(_2144_),
    .X(_2177_));
 sg13g2_buf_2 _7060_ (.A(_2177_),
    .X(_2178_));
 sg13g2_mux2_1 _7061_ (.A0(\logix.ram_r[1856] ),
    .A1(\logix.ram_r[1855] ),
    .S(net331),
    .X(_0957_));
 sg13g2_mux2_1 _7062_ (.A0(\logix.ram_r[1857] ),
    .A1(\logix.ram_r[1856] ),
    .S(net331),
    .X(_0958_));
 sg13g2_mux2_1 _7063_ (.A0(\logix.ram_r[1858] ),
    .A1(\logix.ram_r[1857] ),
    .S(net331),
    .X(_0959_));
 sg13g2_mux2_1 _7064_ (.A0(\logix.ram_r[1859] ),
    .A1(\logix.ram_r[1858] ),
    .S(net331),
    .X(_0960_));
 sg13g2_mux2_1 _7065_ (.A0(\logix.ram_r[185] ),
    .A1(\logix.ram_r[184] ),
    .S(_2178_),
    .X(_0961_));
 sg13g2_mux2_1 _7066_ (.A0(\logix.ram_r[1860] ),
    .A1(\logix.ram_r[1859] ),
    .S(net331),
    .X(_0962_));
 sg13g2_mux2_1 _7067_ (.A0(\logix.ram_r[1861] ),
    .A1(\logix.ram_r[1860] ),
    .S(net331),
    .X(_0963_));
 sg13g2_mux2_1 _7068_ (.A0(\logix.ram_r[1862] ),
    .A1(\logix.ram_r[1861] ),
    .S(net331),
    .X(_0964_));
 sg13g2_mux2_1 _7069_ (.A0(\logix.ram_r[1863] ),
    .A1(\logix.ram_r[1862] ),
    .S(net331),
    .X(_0965_));
 sg13g2_mux2_1 _7070_ (.A0(\logix.ram_r[1864] ),
    .A1(\logix.ram_r[1863] ),
    .S(_2178_),
    .X(_0966_));
 sg13g2_buf_1 _7071_ (.A(_2177_),
    .X(_2179_));
 sg13g2_mux2_1 _7072_ (.A0(\logix.ram_r[1865] ),
    .A1(\logix.ram_r[1864] ),
    .S(net330),
    .X(_0967_));
 sg13g2_mux2_1 _7073_ (.A0(\logix.ram_r[1866] ),
    .A1(\logix.ram_r[1865] ),
    .S(net330),
    .X(_0968_));
 sg13g2_mux2_1 _7074_ (.A0(\logix.ram_r[1867] ),
    .A1(\logix.ram_r[1866] ),
    .S(net330),
    .X(_0969_));
 sg13g2_mux2_1 _7075_ (.A0(\logix.ram_r[1868] ),
    .A1(\logix.ram_r[1867] ),
    .S(_2179_),
    .X(_0970_));
 sg13g2_mux2_1 _7076_ (.A0(\logix.ram_r[1869] ),
    .A1(\logix.ram_r[1868] ),
    .S(net330),
    .X(_0971_));
 sg13g2_mux2_1 _7077_ (.A0(\logix.ram_r[186] ),
    .A1(\logix.ram_r[185] ),
    .S(_2179_),
    .X(_0972_));
 sg13g2_mux2_1 _7078_ (.A0(\logix.ram_r[1870] ),
    .A1(\logix.ram_r[1869] ),
    .S(net330),
    .X(_0973_));
 sg13g2_mux2_1 _7079_ (.A0(\logix.ram_r[1871] ),
    .A1(\logix.ram_r[1870] ),
    .S(net330),
    .X(_0974_));
 sg13g2_mux2_1 _7080_ (.A0(\logix.ram_r[1872] ),
    .A1(\logix.ram_r[1871] ),
    .S(net330),
    .X(_0975_));
 sg13g2_mux2_1 _7081_ (.A0(\logix.ram_r[1873] ),
    .A1(\logix.ram_r[1872] ),
    .S(net330),
    .X(_0976_));
 sg13g2_buf_1 _7082_ (.A(_2177_),
    .X(_2180_));
 sg13g2_mux2_1 _7083_ (.A0(\logix.ram_r[1874] ),
    .A1(\logix.ram_r[1873] ),
    .S(net329),
    .X(_0977_));
 sg13g2_mux2_1 _7084_ (.A0(\logix.ram_r[1875] ),
    .A1(\logix.ram_r[1874] ),
    .S(net329),
    .X(_0978_));
 sg13g2_mux2_1 _7085_ (.A0(\logix.ram_r[1876] ),
    .A1(\logix.ram_r[1875] ),
    .S(_2180_),
    .X(_0979_));
 sg13g2_mux2_1 _7086_ (.A0(\logix.ram_r[1877] ),
    .A1(\logix.ram_r[1876] ),
    .S(net329),
    .X(_0980_));
 sg13g2_mux2_1 _7087_ (.A0(\logix.ram_r[1878] ),
    .A1(\logix.ram_r[1877] ),
    .S(net329),
    .X(_0981_));
 sg13g2_mux2_1 _7088_ (.A0(\logix.ram_r[1879] ),
    .A1(\logix.ram_r[1878] ),
    .S(net329),
    .X(_0982_));
 sg13g2_mux2_1 _7089_ (.A0(\logix.ram_r[187] ),
    .A1(\logix.ram_r[186] ),
    .S(_2180_),
    .X(_0983_));
 sg13g2_mux2_1 _7090_ (.A0(\logix.ram_r[1880] ),
    .A1(\logix.ram_r[1879] ),
    .S(net329),
    .X(_0984_));
 sg13g2_mux2_1 _7091_ (.A0(\logix.ram_r[1881] ),
    .A1(\logix.ram_r[1880] ),
    .S(net329),
    .X(_0985_));
 sg13g2_mux2_1 _7092_ (.A0(\logix.ram_r[1882] ),
    .A1(\logix.ram_r[1881] ),
    .S(net329),
    .X(_0986_));
 sg13g2_buf_1 _7093_ (.A(_2177_),
    .X(_2181_));
 sg13g2_mux2_1 _7094_ (.A0(\logix.ram_r[1883] ),
    .A1(\logix.ram_r[1882] ),
    .S(net328),
    .X(_0987_));
 sg13g2_mux2_1 _7095_ (.A0(\logix.ram_r[1884] ),
    .A1(\logix.ram_r[1883] ),
    .S(_2181_),
    .X(_0988_));
 sg13g2_mux2_1 _7096_ (.A0(\logix.ram_r[1885] ),
    .A1(\logix.ram_r[1884] ),
    .S(net328),
    .X(_0989_));
 sg13g2_mux2_1 _7097_ (.A0(\logix.ram_r[1886] ),
    .A1(\logix.ram_r[1885] ),
    .S(net328),
    .X(_0990_));
 sg13g2_mux2_1 _7098_ (.A0(\logix.ram_r[1887] ),
    .A1(\logix.ram_r[1886] ),
    .S(net328),
    .X(_0991_));
 sg13g2_mux2_1 _7099_ (.A0(\logix.ram_r[1888] ),
    .A1(\logix.ram_r[1887] ),
    .S(net328),
    .X(_0992_));
 sg13g2_mux2_1 _7100_ (.A0(\logix.ram_r[1889] ),
    .A1(\logix.ram_r[1888] ),
    .S(net328),
    .X(_0993_));
 sg13g2_mux2_1 _7101_ (.A0(\logix.ram_r[188] ),
    .A1(\logix.ram_r[187] ),
    .S(_2181_),
    .X(_0994_));
 sg13g2_mux2_1 _7102_ (.A0(\logix.ram_r[1890] ),
    .A1(\logix.ram_r[1889] ),
    .S(net328),
    .X(_0995_));
 sg13g2_mux2_1 _7103_ (.A0(\logix.ram_r[1891] ),
    .A1(\logix.ram_r[1890] ),
    .S(net328),
    .X(_0996_));
 sg13g2_buf_1 _7104_ (.A(_2177_),
    .X(_2182_));
 sg13g2_mux2_1 _7105_ (.A0(\logix.ram_r[1892] ),
    .A1(\logix.ram_r[1891] ),
    .S(net327),
    .X(_0997_));
 sg13g2_mux2_1 _7106_ (.A0(\logix.ram_r[1893] ),
    .A1(\logix.ram_r[1892] ),
    .S(net327),
    .X(_0998_));
 sg13g2_mux2_1 _7107_ (.A0(\logix.ram_r[1894] ),
    .A1(\logix.ram_r[1893] ),
    .S(net327),
    .X(_0999_));
 sg13g2_mux2_1 _7108_ (.A0(\logix.ram_r[1895] ),
    .A1(\logix.ram_r[1894] ),
    .S(net327),
    .X(_1000_));
 sg13g2_mux2_1 _7109_ (.A0(\logix.ram_r[1896] ),
    .A1(\logix.ram_r[1895] ),
    .S(net327),
    .X(_1001_));
 sg13g2_mux2_1 _7110_ (.A0(\logix.ram_r[1897] ),
    .A1(\logix.ram_r[1896] ),
    .S(_2182_),
    .X(_1002_));
 sg13g2_mux2_1 _7111_ (.A0(\logix.ram_r[1898] ),
    .A1(\logix.ram_r[1897] ),
    .S(net327),
    .X(_1003_));
 sg13g2_mux2_1 _7112_ (.A0(\logix.ram_r[1899] ),
    .A1(\logix.ram_r[1898] ),
    .S(net327),
    .X(_1004_));
 sg13g2_mux2_1 _7113_ (.A0(\logix.ram_r[189] ),
    .A1(\logix.ram_r[188] ),
    .S(net327),
    .X(_1005_));
 sg13g2_mux2_1 _7114_ (.A0(\logix.ram_r[18] ),
    .A1(\logix.ram_r[17] ),
    .S(_2182_),
    .X(_1006_));
 sg13g2_buf_1 _7115_ (.A(_2177_),
    .X(_2183_));
 sg13g2_mux2_1 _7116_ (.A0(\logix.ram_r[1900] ),
    .A1(\logix.ram_r[1899] ),
    .S(net326),
    .X(_1007_));
 sg13g2_mux2_1 _7117_ (.A0(\logix.ram_r[1901] ),
    .A1(\logix.ram_r[1900] ),
    .S(net326),
    .X(_1008_));
 sg13g2_mux2_1 _7118_ (.A0(\logix.ram_r[1902] ),
    .A1(\logix.ram_r[1901] ),
    .S(net326),
    .X(_1009_));
 sg13g2_mux2_1 _7119_ (.A0(\logix.ram_r[1903] ),
    .A1(\logix.ram_r[1902] ),
    .S(net326),
    .X(_1010_));
 sg13g2_mux2_1 _7120_ (.A0(\logix.ram_r[1904] ),
    .A1(\logix.ram_r[1903] ),
    .S(net326),
    .X(_1011_));
 sg13g2_mux2_1 _7121_ (.A0(\logix.ram_r[1905] ),
    .A1(\logix.ram_r[1904] ),
    .S(net326),
    .X(_1012_));
 sg13g2_mux2_1 _7122_ (.A0(\logix.ram_r[1906] ),
    .A1(\logix.ram_r[1905] ),
    .S(net326),
    .X(_1013_));
 sg13g2_mux2_1 _7123_ (.A0(\logix.ram_r[1907] ),
    .A1(\logix.ram_r[1906] ),
    .S(_2183_),
    .X(_1014_));
 sg13g2_mux2_1 _7124_ (.A0(\logix.ram_r[1908] ),
    .A1(\logix.ram_r[1907] ),
    .S(_2183_),
    .X(_1015_));
 sg13g2_mux2_1 _7125_ (.A0(\logix.ram_r[1909] ),
    .A1(\logix.ram_r[1908] ),
    .S(net326),
    .X(_1016_));
 sg13g2_buf_1 _7126_ (.A(_2177_),
    .X(_2184_));
 sg13g2_mux2_1 _7127_ (.A0(\logix.ram_r[190] ),
    .A1(\logix.ram_r[189] ),
    .S(_2184_),
    .X(_1017_));
 sg13g2_mux2_1 _7128_ (.A0(\logix.ram_r[1910] ),
    .A1(\logix.ram_r[1909] ),
    .S(net325),
    .X(_1018_));
 sg13g2_mux2_1 _7129_ (.A0(\logix.ram_r[1911] ),
    .A1(\logix.ram_r[1910] ),
    .S(net325),
    .X(_1019_));
 sg13g2_mux2_1 _7130_ (.A0(\logix.ram_r[1912] ),
    .A1(\logix.ram_r[1911] ),
    .S(net325),
    .X(_1020_));
 sg13g2_mux2_1 _7131_ (.A0(\logix.ram_r[1913] ),
    .A1(\logix.ram_r[1912] ),
    .S(net325),
    .X(_1021_));
 sg13g2_mux2_1 _7132_ (.A0(\logix.ram_r[1914] ),
    .A1(\logix.ram_r[1913] ),
    .S(net325),
    .X(_1022_));
 sg13g2_mux2_1 _7133_ (.A0(\logix.ram_r[1915] ),
    .A1(\logix.ram_r[1914] ),
    .S(net325),
    .X(_1023_));
 sg13g2_mux2_1 _7134_ (.A0(\logix.ram_r[1916] ),
    .A1(\logix.ram_r[1915] ),
    .S(_2184_),
    .X(_1024_));
 sg13g2_mux2_1 _7135_ (.A0(\logix.ram_r[1917] ),
    .A1(\logix.ram_r[1916] ),
    .S(net325),
    .X(_1025_));
 sg13g2_mux2_1 _7136_ (.A0(\logix.ram_r[1918] ),
    .A1(\logix.ram_r[1917] ),
    .S(net325),
    .X(_1026_));
 sg13g2_buf_1 _7137_ (.A(_2144_),
    .X(_2185_));
 sg13g2_buf_1 _7138_ (.A(_2185_),
    .X(_2186_));
 sg13g2_mux2_1 _7139_ (.A0(\logix.ram_r[1919] ),
    .A1(\logix.ram_r[1918] ),
    .S(_2186_),
    .X(_1027_));
 sg13g2_mux2_1 _7140_ (.A0(\logix.ram_r[191] ),
    .A1(\logix.ram_r[190] ),
    .S(_2186_),
    .X(_1028_));
 sg13g2_mux2_1 _7141_ (.A0(\logix.ram_r[1920] ),
    .A1(\logix.ram_r[1919] ),
    .S(net324),
    .X(_1029_));
 sg13g2_mux2_1 _7142_ (.A0(\logix.ram_r[1921] ),
    .A1(\logix.ram_r[1920] ),
    .S(net324),
    .X(_1030_));
 sg13g2_mux2_1 _7143_ (.A0(\logix.ram_r[1922] ),
    .A1(\logix.ram_r[1921] ),
    .S(net324),
    .X(_1031_));
 sg13g2_mux2_1 _7144_ (.A0(\logix.ram_r[1923] ),
    .A1(\logix.ram_r[1922] ),
    .S(net324),
    .X(_1032_));
 sg13g2_mux2_1 _7145_ (.A0(\logix.ram_r[1924] ),
    .A1(\logix.ram_r[1923] ),
    .S(net324),
    .X(_1033_));
 sg13g2_mux2_1 _7146_ (.A0(\logix.ram_r[1925] ),
    .A1(\logix.ram_r[1924] ),
    .S(net324),
    .X(_1034_));
 sg13g2_mux2_1 _7147_ (.A0(\logix.ram_r[1926] ),
    .A1(\logix.ram_r[1925] ),
    .S(net324),
    .X(_1035_));
 sg13g2_mux2_1 _7148_ (.A0(\logix.ram_r[1927] ),
    .A1(\logix.ram_r[1926] ),
    .S(net324),
    .X(_1036_));
 sg13g2_buf_2 _7149_ (.A(_2185_),
    .X(_2187_));
 sg13g2_mux2_1 _7150_ (.A0(\logix.ram_r[1928] ),
    .A1(\logix.ram_r[1927] ),
    .S(net323),
    .X(_1037_));
 sg13g2_mux2_1 _7151_ (.A0(\logix.ram_r[1929] ),
    .A1(\logix.ram_r[1928] ),
    .S(_2187_),
    .X(_1038_));
 sg13g2_mux2_1 _7152_ (.A0(\logix.ram_r[192] ),
    .A1(\logix.ram_r[191] ),
    .S(net323),
    .X(_1039_));
 sg13g2_mux2_1 _7153_ (.A0(\logix.ram_r[1930] ),
    .A1(\logix.ram_r[1929] ),
    .S(net323),
    .X(_1040_));
 sg13g2_mux2_1 _7154_ (.A0(\logix.ram_r[1931] ),
    .A1(\logix.ram_r[1930] ),
    .S(net323),
    .X(_1041_));
 sg13g2_mux2_1 _7155_ (.A0(\logix.ram_r[1932] ),
    .A1(\logix.ram_r[1931] ),
    .S(net323),
    .X(_1042_));
 sg13g2_mux2_1 _7156_ (.A0(\logix.ram_r[1933] ),
    .A1(\logix.ram_r[1932] ),
    .S(net323),
    .X(_1043_));
 sg13g2_mux2_1 _7157_ (.A0(\logix.ram_r[1934] ),
    .A1(\logix.ram_r[1933] ),
    .S(net323),
    .X(_1044_));
 sg13g2_mux2_1 _7158_ (.A0(\logix.ram_r[1935] ),
    .A1(\logix.ram_r[1934] ),
    .S(_2187_),
    .X(_1045_));
 sg13g2_mux2_1 _7159_ (.A0(\logix.ram_r[1936] ),
    .A1(\logix.ram_r[1935] ),
    .S(net323),
    .X(_1046_));
 sg13g2_buf_1 _7160_ (.A(_2185_),
    .X(_2188_));
 sg13g2_mux2_1 _7161_ (.A0(\logix.ram_r[1937] ),
    .A1(\logix.ram_r[1936] ),
    .S(net322),
    .X(_1047_));
 sg13g2_mux2_1 _7162_ (.A0(\logix.ram_r[1938] ),
    .A1(\logix.ram_r[1937] ),
    .S(net322),
    .X(_1048_));
 sg13g2_mux2_1 _7163_ (.A0(\logix.ram_r[1939] ),
    .A1(\logix.ram_r[1938] ),
    .S(net322),
    .X(_1049_));
 sg13g2_mux2_1 _7164_ (.A0(\logix.ram_r[193] ),
    .A1(\logix.ram_r[192] ),
    .S(_2188_),
    .X(_1050_));
 sg13g2_mux2_1 _7165_ (.A0(\logix.ram_r[1940] ),
    .A1(\logix.ram_r[1939] ),
    .S(net322),
    .X(_1051_));
 sg13g2_mux2_1 _7166_ (.A0(\logix.ram_r[1941] ),
    .A1(\logix.ram_r[1940] ),
    .S(net322),
    .X(_1052_));
 sg13g2_mux2_1 _7167_ (.A0(\logix.ram_r[1942] ),
    .A1(\logix.ram_r[1941] ),
    .S(net322),
    .X(_1053_));
 sg13g2_mux2_1 _7168_ (.A0(\logix.ram_r[1943] ),
    .A1(\logix.ram_r[1942] ),
    .S(net322),
    .X(_1054_));
 sg13g2_mux2_1 _7169_ (.A0(\logix.ram_r[1944] ),
    .A1(\logix.ram_r[1943] ),
    .S(net322),
    .X(_1055_));
 sg13g2_mux2_1 _7170_ (.A0(\logix.ram_r[1945] ),
    .A1(\logix.ram_r[1944] ),
    .S(_2188_),
    .X(_1056_));
 sg13g2_buf_1 _7171_ (.A(_2185_),
    .X(_2189_));
 sg13g2_mux2_1 _7172_ (.A0(\logix.ram_r[1946] ),
    .A1(\logix.ram_r[1945] ),
    .S(net321),
    .X(_1057_));
 sg13g2_mux2_1 _7173_ (.A0(\logix.ram_r[1947] ),
    .A1(\logix.ram_r[1946] ),
    .S(net321),
    .X(_1058_));
 sg13g2_mux2_1 _7174_ (.A0(\logix.ram_r[1948] ),
    .A1(\logix.ram_r[1947] ),
    .S(net321),
    .X(_1059_));
 sg13g2_mux2_1 _7175_ (.A0(\logix.ram_r[1949] ),
    .A1(\logix.ram_r[1948] ),
    .S(net321),
    .X(_1060_));
 sg13g2_mux2_1 _7176_ (.A0(\logix.ram_r[194] ),
    .A1(\logix.ram_r[193] ),
    .S(net321),
    .X(_1061_));
 sg13g2_mux2_1 _7177_ (.A0(\logix.ram_r[1950] ),
    .A1(\logix.ram_r[1949] ),
    .S(_2189_),
    .X(_1062_));
 sg13g2_mux2_1 _7178_ (.A0(\logix.ram_r[1951] ),
    .A1(\logix.ram_r[1950] ),
    .S(_2189_),
    .X(_1063_));
 sg13g2_mux2_1 _7179_ (.A0(\logix.ram_r[1952] ),
    .A1(\logix.ram_r[1951] ),
    .S(net321),
    .X(_1064_));
 sg13g2_mux2_1 _7180_ (.A0(\logix.ram_r[1953] ),
    .A1(\logix.ram_r[1952] ),
    .S(net321),
    .X(_1065_));
 sg13g2_mux2_1 _7181_ (.A0(\logix.ram_r[1954] ),
    .A1(\logix.ram_r[1953] ),
    .S(net321),
    .X(_1066_));
 sg13g2_buf_1 _7182_ (.A(_2185_),
    .X(_2190_));
 sg13g2_mux2_1 _7183_ (.A0(\logix.ram_r[1955] ),
    .A1(\logix.ram_r[1954] ),
    .S(net320),
    .X(_1067_));
 sg13g2_mux2_1 _7184_ (.A0(\logix.ram_r[1956] ),
    .A1(\logix.ram_r[1955] ),
    .S(net320),
    .X(_1068_));
 sg13g2_mux2_1 _7185_ (.A0(\logix.ram_r[1957] ),
    .A1(\logix.ram_r[1956] ),
    .S(net320),
    .X(_1069_));
 sg13g2_mux2_1 _7186_ (.A0(\logix.ram_r[1958] ),
    .A1(\logix.ram_r[1957] ),
    .S(net320),
    .X(_1070_));
 sg13g2_mux2_1 _7187_ (.A0(\logix.ram_r[1959] ),
    .A1(\logix.ram_r[1958] ),
    .S(net320),
    .X(_1071_));
 sg13g2_mux2_1 _7188_ (.A0(\logix.ram_r[195] ),
    .A1(\logix.ram_r[194] ),
    .S(_2190_),
    .X(_1072_));
 sg13g2_mux2_1 _7189_ (.A0(\logix.ram_r[1960] ),
    .A1(\logix.ram_r[1959] ),
    .S(_2190_),
    .X(_1073_));
 sg13g2_mux2_1 _7190_ (.A0(\logix.ram_r[1961] ),
    .A1(\logix.ram_r[1960] ),
    .S(net320),
    .X(_1074_));
 sg13g2_mux2_1 _7191_ (.A0(\logix.ram_r[1962] ),
    .A1(\logix.ram_r[1961] ),
    .S(net320),
    .X(_1075_));
 sg13g2_mux2_1 _7192_ (.A0(\logix.ram_r[1963] ),
    .A1(\logix.ram_r[1962] ),
    .S(net320),
    .X(_1076_));
 sg13g2_buf_1 _7193_ (.A(_2185_),
    .X(_2191_));
 sg13g2_mux2_1 _7194_ (.A0(\logix.ram_r[1964] ),
    .A1(\logix.ram_r[1963] ),
    .S(net319),
    .X(_1077_));
 sg13g2_mux2_1 _7195_ (.A0(\logix.ram_r[1965] ),
    .A1(\logix.ram_r[1964] ),
    .S(net319),
    .X(_1078_));
 sg13g2_mux2_1 _7196_ (.A0(\logix.ram_r[1966] ),
    .A1(\logix.ram_r[1965] ),
    .S(net319),
    .X(_1079_));
 sg13g2_mux2_1 _7197_ (.A0(\logix.ram_r[1967] ),
    .A1(\logix.ram_r[1966] ),
    .S(net319),
    .X(_1080_));
 sg13g2_mux2_1 _7198_ (.A0(\logix.ram_r[1968] ),
    .A1(\logix.ram_r[1967] ),
    .S(net319),
    .X(_1081_));
 sg13g2_mux2_1 _7199_ (.A0(\logix.ram_r[1969] ),
    .A1(\logix.ram_r[1968] ),
    .S(_2191_),
    .X(_1082_));
 sg13g2_mux2_1 _7200_ (.A0(\logix.ram_r[196] ),
    .A1(\logix.ram_r[195] ),
    .S(_2191_),
    .X(_1083_));
 sg13g2_mux2_1 _7201_ (.A0(\logix.ram_r[1970] ),
    .A1(\logix.ram_r[1969] ),
    .S(net319),
    .X(_1084_));
 sg13g2_mux2_1 _7202_ (.A0(\logix.ram_r[1971] ),
    .A1(\logix.ram_r[1970] ),
    .S(net319),
    .X(_1085_));
 sg13g2_mux2_1 _7203_ (.A0(\logix.ram_r[1972] ),
    .A1(\logix.ram_r[1971] ),
    .S(net319),
    .X(_1086_));
 sg13g2_buf_1 _7204_ (.A(_2185_),
    .X(_2192_));
 sg13g2_mux2_1 _7205_ (.A0(\logix.ram_r[1973] ),
    .A1(\logix.ram_r[1972] ),
    .S(net318),
    .X(_1087_));
 sg13g2_mux2_1 _7206_ (.A0(\logix.ram_r[1974] ),
    .A1(\logix.ram_r[1973] ),
    .S(net318),
    .X(_1088_));
 sg13g2_mux2_1 _7207_ (.A0(\logix.ram_r[1975] ),
    .A1(\logix.ram_r[1974] ),
    .S(net318),
    .X(_1089_));
 sg13g2_mux2_1 _7208_ (.A0(\logix.ram_r[1976] ),
    .A1(\logix.ram_r[1975] ),
    .S(_2192_),
    .X(_1090_));
 sg13g2_mux2_1 _7209_ (.A0(\logix.ram_r[1977] ),
    .A1(\logix.ram_r[1976] ),
    .S(net318),
    .X(_1091_));
 sg13g2_mux2_1 _7210_ (.A0(\logix.ram_r[1978] ),
    .A1(\logix.ram_r[1977] ),
    .S(net318),
    .X(_1092_));
 sg13g2_mux2_1 _7211_ (.A0(\logix.ram_r[1979] ),
    .A1(\logix.ram_r[1978] ),
    .S(net318),
    .X(_1093_));
 sg13g2_mux2_1 _7212_ (.A0(\logix.ram_r[197] ),
    .A1(\logix.ram_r[196] ),
    .S(_2192_),
    .X(_1094_));
 sg13g2_mux2_1 _7213_ (.A0(\logix.ram_r[1980] ),
    .A1(\logix.ram_r[1979] ),
    .S(net318),
    .X(_1095_));
 sg13g2_mux2_1 _7214_ (.A0(\logix.ram_r[1981] ),
    .A1(\logix.ram_r[1980] ),
    .S(net318),
    .X(_1096_));
 sg13g2_buf_1 _7215_ (.A(_2144_),
    .X(_2193_));
 sg13g2_buf_1 _7216_ (.A(_2193_),
    .X(_2194_));
 sg13g2_mux2_1 _7217_ (.A0(\logix.ram_r[1982] ),
    .A1(\logix.ram_r[1981] ),
    .S(net317),
    .X(_1097_));
 sg13g2_mux2_1 _7218_ (.A0(\logix.ram_r[1983] ),
    .A1(\logix.ram_r[1982] ),
    .S(net317),
    .X(_1098_));
 sg13g2_mux2_1 _7219_ (.A0(\logix.ram_r[1984] ),
    .A1(\logix.ram_r[1983] ),
    .S(_2194_),
    .X(_1099_));
 sg13g2_mux2_1 _7220_ (.A0(\logix.ram_r[1985] ),
    .A1(\logix.ram_r[1984] ),
    .S(_2194_),
    .X(_1100_));
 sg13g2_mux2_1 _7221_ (.A0(\logix.ram_r[1986] ),
    .A1(\logix.ram_r[1985] ),
    .S(net317),
    .X(_1101_));
 sg13g2_mux2_1 _7222_ (.A0(\logix.ram_r[1987] ),
    .A1(\logix.ram_r[1986] ),
    .S(net317),
    .X(_1102_));
 sg13g2_mux2_1 _7223_ (.A0(\logix.ram_r[1988] ),
    .A1(\logix.ram_r[1987] ),
    .S(net317),
    .X(_1103_));
 sg13g2_mux2_1 _7224_ (.A0(\logix.ram_r[1989] ),
    .A1(\logix.ram_r[1988] ),
    .S(net317),
    .X(_1104_));
 sg13g2_mux2_1 _7225_ (.A0(\logix.ram_r[198] ),
    .A1(\logix.ram_r[197] ),
    .S(net317),
    .X(_1105_));
 sg13g2_mux2_1 _7226_ (.A0(\logix.ram_r[1990] ),
    .A1(\logix.ram_r[1989] ),
    .S(net317),
    .X(_1106_));
 sg13g2_buf_1 _7227_ (.A(_2193_),
    .X(_2195_));
 sg13g2_mux2_1 _7228_ (.A0(\logix.ram_r[1991] ),
    .A1(\logix.ram_r[1990] ),
    .S(_2195_),
    .X(_1107_));
 sg13g2_mux2_1 _7229_ (.A0(\logix.ram_r[1992] ),
    .A1(\logix.ram_r[1991] ),
    .S(net316),
    .X(_1108_));
 sg13g2_mux2_1 _7230_ (.A0(\logix.ram_r[1993] ),
    .A1(\logix.ram_r[1992] ),
    .S(net316),
    .X(_1109_));
 sg13g2_mux2_1 _7231_ (.A0(\logix.ram_r[1994] ),
    .A1(\logix.ram_r[1993] ),
    .S(net316),
    .X(_1110_));
 sg13g2_mux2_1 _7232_ (.A0(\logix.ram_r[1995] ),
    .A1(\logix.ram_r[1994] ),
    .S(net316),
    .X(_1111_));
 sg13g2_mux2_1 _7233_ (.A0(\logix.ram_r[1996] ),
    .A1(\logix.ram_r[1995] ),
    .S(net316),
    .X(_1112_));
 sg13g2_mux2_1 _7234_ (.A0(\logix.ram_r[1997] ),
    .A1(\logix.ram_r[1996] ),
    .S(net316),
    .X(_1113_));
 sg13g2_mux2_1 _7235_ (.A0(\logix.ram_r[1998] ),
    .A1(\logix.ram_r[1997] ),
    .S(net316),
    .X(_1114_));
 sg13g2_mux2_1 _7236_ (.A0(\logix.ram_r[1999] ),
    .A1(\logix.ram_r[1998] ),
    .S(_2195_),
    .X(_1115_));
 sg13g2_mux2_1 _7237_ (.A0(\logix.ram_r[199] ),
    .A1(\logix.ram_r[198] ),
    .S(net316),
    .X(_1116_));
 sg13g2_buf_2 _7238_ (.A(_2193_),
    .X(_2196_));
 sg13g2_mux2_1 _7239_ (.A0(\logix.ram_r[19] ),
    .A1(\logix.ram_r[18] ),
    .S(_2196_),
    .X(_1117_));
 sg13g2_mux2_1 _7240_ (.A0(\logix.ram_r[1] ),
    .A1(\logix.ram_r[0] ),
    .S(_2196_),
    .X(_1118_));
 sg13g2_mux2_1 _7241_ (.A0(\logix.ram_r[2000] ),
    .A1(\logix.ram_r[1999] ),
    .S(net315),
    .X(_1119_));
 sg13g2_mux2_1 _7242_ (.A0(\logix.ram_r[2001] ),
    .A1(\logix.ram_r[2000] ),
    .S(net315),
    .X(_1120_));
 sg13g2_mux2_1 _7243_ (.A0(\logix.ram_r[2002] ),
    .A1(\logix.ram_r[2001] ),
    .S(net315),
    .X(_1121_));
 sg13g2_mux2_1 _7244_ (.A0(\logix.ram_r[2003] ),
    .A1(\logix.ram_r[2002] ),
    .S(net315),
    .X(_1122_));
 sg13g2_mux2_1 _7245_ (.A0(\logix.ram_r[2004] ),
    .A1(\logix.ram_r[2003] ),
    .S(net315),
    .X(_1123_));
 sg13g2_mux2_1 _7246_ (.A0(\logix.ram_r[2005] ),
    .A1(\logix.ram_r[2004] ),
    .S(net315),
    .X(_1124_));
 sg13g2_mux2_1 _7247_ (.A0(\logix.ram_r[2006] ),
    .A1(\logix.ram_r[2005] ),
    .S(net315),
    .X(_1125_));
 sg13g2_mux2_1 _7248_ (.A0(\logix.ram_r[2007] ),
    .A1(\logix.ram_r[2006] ),
    .S(net315),
    .X(_1126_));
 sg13g2_buf_1 _7249_ (.A(_2193_),
    .X(_2197_));
 sg13g2_mux2_1 _7250_ (.A0(\logix.ram_r[2008] ),
    .A1(\logix.ram_r[2007] ),
    .S(net314),
    .X(_1127_));
 sg13g2_mux2_1 _7251_ (.A0(\logix.ram_r[2009] ),
    .A1(\logix.ram_r[2008] ),
    .S(net314),
    .X(_1128_));
 sg13g2_mux2_1 _7252_ (.A0(\logix.ram_r[200] ),
    .A1(\logix.ram_r[199] ),
    .S(net314),
    .X(_1129_));
 sg13g2_mux2_1 _7253_ (.A0(\logix.ram_r[2010] ),
    .A1(\logix.ram_r[2009] ),
    .S(net314),
    .X(_1130_));
 sg13g2_mux2_1 _7254_ (.A0(\logix.ram_r[2011] ),
    .A1(\logix.ram_r[2010] ),
    .S(net314),
    .X(_1131_));
 sg13g2_mux2_1 _7255_ (.A0(\logix.ram_r[2012] ),
    .A1(\logix.ram_r[2011] ),
    .S(net314),
    .X(_1132_));
 sg13g2_mux2_1 _7256_ (.A0(\logix.ram_r[2013] ),
    .A1(\logix.ram_r[2012] ),
    .S(net314),
    .X(_1133_));
 sg13g2_mux2_1 _7257_ (.A0(\logix.ram_r[2014] ),
    .A1(\logix.ram_r[2013] ),
    .S(_2197_),
    .X(_1134_));
 sg13g2_mux2_1 _7258_ (.A0(\logix.ram_r[2015] ),
    .A1(\logix.ram_r[2014] ),
    .S(_2197_),
    .X(_1135_));
 sg13g2_mux2_1 _7259_ (.A0(\logix.ram_r[2016] ),
    .A1(\logix.ram_r[2015] ),
    .S(net314),
    .X(_1136_));
 sg13g2_buf_1 _7260_ (.A(_2193_),
    .X(_2198_));
 sg13g2_mux2_1 _7261_ (.A0(\logix.ram_r[2017] ),
    .A1(\logix.ram_r[2016] ),
    .S(net313),
    .X(_1137_));
 sg13g2_mux2_1 _7262_ (.A0(\logix.ram_r[2018] ),
    .A1(\logix.ram_r[2017] ),
    .S(net313),
    .X(_1138_));
 sg13g2_mux2_1 _7263_ (.A0(\logix.ram_r[2019] ),
    .A1(\logix.ram_r[2018] ),
    .S(net313),
    .X(_1139_));
 sg13g2_mux2_1 _7264_ (.A0(\logix.ram_r[201] ),
    .A1(\logix.ram_r[200] ),
    .S(net313),
    .X(_1140_));
 sg13g2_mux2_1 _7265_ (.A0(\logix.ram_r[2020] ),
    .A1(\logix.ram_r[2019] ),
    .S(net313),
    .X(_1141_));
 sg13g2_mux2_1 _7266_ (.A0(\logix.ram_r[2021] ),
    .A1(\logix.ram_r[2020] ),
    .S(net313),
    .X(_1142_));
 sg13g2_mux2_1 _7267_ (.A0(\logix.ram_r[2022] ),
    .A1(\logix.ram_r[2021] ),
    .S(_2198_),
    .X(_1143_));
 sg13g2_mux2_1 _7268_ (.A0(\logix.ram_r[2023] ),
    .A1(\logix.ram_r[2022] ),
    .S(_2198_),
    .X(_1144_));
 sg13g2_mux2_1 _7269_ (.A0(\logix.ram_r[2024] ),
    .A1(\logix.ram_r[2023] ),
    .S(net313),
    .X(_1145_));
 sg13g2_mux2_1 _7270_ (.A0(\logix.ram_r[2025] ),
    .A1(\logix.ram_r[2024] ),
    .S(net313),
    .X(_1146_));
 sg13g2_buf_1 _7271_ (.A(_2193_),
    .X(_2199_));
 sg13g2_mux2_1 _7272_ (.A0(\logix.ram_r[2026] ),
    .A1(\logix.ram_r[2025] ),
    .S(net312),
    .X(_1147_));
 sg13g2_mux2_1 _7273_ (.A0(\logix.ram_r[2027] ),
    .A1(\logix.ram_r[2026] ),
    .S(net312),
    .X(_1148_));
 sg13g2_mux2_1 _7274_ (.A0(\logix.ram_r[2028] ),
    .A1(\logix.ram_r[2027] ),
    .S(net312),
    .X(_1149_));
 sg13g2_mux2_1 _7275_ (.A0(\logix.ram_r[2029] ),
    .A1(\logix.ram_r[2028] ),
    .S(net312),
    .X(_1150_));
 sg13g2_mux2_1 _7276_ (.A0(\logix.ram_r[202] ),
    .A1(\logix.ram_r[201] ),
    .S(_2199_),
    .X(_1151_));
 sg13g2_mux2_1 _7277_ (.A0(\logix.ram_r[2030] ),
    .A1(\logix.ram_r[2029] ),
    .S(_2199_),
    .X(_1152_));
 sg13g2_mux2_1 _7278_ (.A0(\logix.ram_r[2031] ),
    .A1(\logix.ram_r[2030] ),
    .S(net312),
    .X(_1153_));
 sg13g2_mux2_1 _7279_ (.A0(\logix.ram_r[2032] ),
    .A1(\logix.ram_r[2031] ),
    .S(net312),
    .X(_1154_));
 sg13g2_mux2_1 _7280_ (.A0(\logix.ram_r[2033] ),
    .A1(\logix.ram_r[2032] ),
    .S(net312),
    .X(_1155_));
 sg13g2_mux2_1 _7281_ (.A0(\logix.ram_r[2034] ),
    .A1(\logix.ram_r[2033] ),
    .S(net312),
    .X(_1156_));
 sg13g2_buf_1 _7282_ (.A(_2193_),
    .X(_2200_));
 sg13g2_mux2_1 _7283_ (.A0(\logix.ram_r[2035] ),
    .A1(\logix.ram_r[2034] ),
    .S(net311),
    .X(_1157_));
 sg13g2_mux2_1 _7284_ (.A0(\logix.ram_r[2036] ),
    .A1(\logix.ram_r[2035] ),
    .S(net311),
    .X(_1158_));
 sg13g2_mux2_1 _7285_ (.A0(\logix.ram_r[2037] ),
    .A1(\logix.ram_r[2036] ),
    .S(net311),
    .X(_1159_));
 sg13g2_mux2_1 _7286_ (.A0(\logix.ram_r[2038] ),
    .A1(\logix.ram_r[2037] ),
    .S(net311),
    .X(_1160_));
 sg13g2_mux2_1 _7287_ (.A0(\logix.ram_r[2039] ),
    .A1(\logix.ram_r[2038] ),
    .S(_2200_),
    .X(_1161_));
 sg13g2_mux2_1 _7288_ (.A0(\logix.ram_r[203] ),
    .A1(\logix.ram_r[202] ),
    .S(_2200_),
    .X(_1162_));
 sg13g2_mux2_1 _7289_ (.A0(\logix.ram_r[2040] ),
    .A1(\logix.ram_r[2039] ),
    .S(net311),
    .X(_1163_));
 sg13g2_mux2_1 _7290_ (.A0(\logix.ram_r[2041] ),
    .A1(\logix.ram_r[2040] ),
    .S(net311),
    .X(_1164_));
 sg13g2_mux2_1 _7291_ (.A0(\logix.ram_r[2042] ),
    .A1(\logix.ram_r[2041] ),
    .S(net311),
    .X(_1165_));
 sg13g2_mux2_1 _7292_ (.A0(\logix.ram_r[2043] ),
    .A1(\logix.ram_r[2042] ),
    .S(net311),
    .X(_1166_));
 sg13g2_buf_2 _7293_ (.A(_2063_),
    .X(_2201_));
 sg13g2_buf_1 _7294_ (.A(_2201_),
    .X(_2202_));
 sg13g2_buf_1 _7295_ (.A(_2202_),
    .X(_2203_));
 sg13g2_mux2_1 _7296_ (.A0(\logix.ram_r[2044] ),
    .A1(\logix.ram_r[2043] ),
    .S(net310),
    .X(_1167_));
 sg13g2_mux2_1 _7297_ (.A0(\logix.ram_r[2045] ),
    .A1(\logix.ram_r[2044] ),
    .S(net310),
    .X(_1168_));
 sg13g2_mux2_1 _7298_ (.A0(\logix.ram_r[2046] ),
    .A1(\logix.ram_r[2045] ),
    .S(net310),
    .X(_1169_));
 sg13g2_mux2_1 _7299_ (.A0(\logix.ram_r[2047] ),
    .A1(\logix.ram_r[2046] ),
    .S(net310),
    .X(_1170_));
 sg13g2_buf_8 _7300_ (.A(\logix.input_sel_cfg_w[0] ),
    .X(_2204_));
 sg13g2_mux2_1 _7301_ (.A0(_2204_),
    .A1(\logix.ram_r[2047] ),
    .S(net310),
    .X(_1171_));
 sg13g2_buf_8 _7302_ (.A(\logix.input_sel_cfg_w[1] ),
    .X(_2205_));
 sg13g2_mux2_1 _7303_ (.A0(_2205_),
    .A1(_2204_),
    .S(net310),
    .X(_1172_));
 sg13g2_mux2_1 _7304_ (.A0(\logix.ram_r[204] ),
    .A1(\logix.ram_r[203] ),
    .S(_2203_),
    .X(_1173_));
 sg13g2_buf_8 _7305_ (.A(\logix.input_sel_cfg_w[2] ),
    .X(_2206_));
 sg13g2_mux2_1 _7306_ (.A0(_2206_),
    .A1(_2205_),
    .S(net310),
    .X(_1174_));
 sg13g2_buf_8 _7307_ (.A(\logix.input_sel_cfg_w[3] ),
    .X(_2207_));
 sg13g2_mux2_1 _7308_ (.A0(_2207_),
    .A1(_2206_),
    .S(net310),
    .X(_1175_));
 sg13g2_buf_1 _7309_ (.A(\logix.input_sel_cfg_w[4] ),
    .X(_2208_));
 sg13g2_mux2_1 _7310_ (.A0(_2208_),
    .A1(_2207_),
    .S(_2203_),
    .X(_1176_));
 sg13g2_buf_1 _7311_ (.A(\logix.input_sel_cfg_w[5] ),
    .X(_2209_));
 sg13g2_buf_2 _7312_ (.A(_2202_),
    .X(_2210_));
 sg13g2_mux2_1 _7313_ (.A0(_2209_),
    .A1(_2208_),
    .S(net309),
    .X(_1177_));
 sg13g2_buf_1 _7314_ (.A(\logix.input_sel_cfg_w[6] ),
    .X(_2211_));
 sg13g2_mux2_1 _7315_ (.A0(_2211_),
    .A1(_2209_),
    .S(net309),
    .X(_1178_));
 sg13g2_buf_1 _7316_ (.A(\logix.input_sel_cfg_w[7] ),
    .X(_2212_));
 sg13g2_mux2_1 _7317_ (.A0(_2212_),
    .A1(_2211_),
    .S(_2210_),
    .X(_1179_));
 sg13g2_mux2_1 _7318_ (.A0(\logix.ram_r[205] ),
    .A1(\logix.ram_r[204] ),
    .S(net309),
    .X(_1180_));
 sg13g2_mux2_1 _7319_ (.A0(\logix.ram_r[206] ),
    .A1(\logix.ram_r[205] ),
    .S(net309),
    .X(_1181_));
 sg13g2_mux2_1 _7320_ (.A0(\logix.ram_r[207] ),
    .A1(\logix.ram_r[206] ),
    .S(net309),
    .X(_1182_));
 sg13g2_mux2_1 _7321_ (.A0(\logix.ram_r[208] ),
    .A1(\logix.ram_r[207] ),
    .S(net309),
    .X(_1183_));
 sg13g2_mux2_1 _7322_ (.A0(\logix.ram_r[209] ),
    .A1(\logix.ram_r[208] ),
    .S(net309),
    .X(_1184_));
 sg13g2_mux2_1 _7323_ (.A0(\logix.ram_r[20] ),
    .A1(\logix.ram_r[19] ),
    .S(_2210_),
    .X(_1185_));
 sg13g2_mux2_1 _7324_ (.A0(\logix.ram_r[210] ),
    .A1(\logix.ram_r[209] ),
    .S(net309),
    .X(_1186_));
 sg13g2_buf_1 _7325_ (.A(_2202_),
    .X(_2213_));
 sg13g2_mux2_1 _7326_ (.A0(\logix.ram_r[211] ),
    .A1(\logix.ram_r[210] ),
    .S(net308),
    .X(_1187_));
 sg13g2_mux2_1 _7327_ (.A0(\logix.ram_r[212] ),
    .A1(\logix.ram_r[211] ),
    .S(net308),
    .X(_1188_));
 sg13g2_mux2_1 _7328_ (.A0(\logix.ram_r[213] ),
    .A1(\logix.ram_r[212] ),
    .S(net308),
    .X(_1189_));
 sg13g2_mux2_1 _7329_ (.A0(\logix.ram_r[214] ),
    .A1(\logix.ram_r[213] ),
    .S(net308),
    .X(_1190_));
 sg13g2_mux2_1 _7330_ (.A0(\logix.ram_r[215] ),
    .A1(\logix.ram_r[214] ),
    .S(_2213_),
    .X(_1191_));
 sg13g2_mux2_1 _7331_ (.A0(\logix.ram_r[216] ),
    .A1(\logix.ram_r[215] ),
    .S(net308),
    .X(_1192_));
 sg13g2_mux2_1 _7332_ (.A0(\logix.ram_r[217] ),
    .A1(\logix.ram_r[216] ),
    .S(net308),
    .X(_1193_));
 sg13g2_mux2_1 _7333_ (.A0(\logix.ram_r[218] ),
    .A1(\logix.ram_r[217] ),
    .S(net308),
    .X(_1194_));
 sg13g2_mux2_1 _7334_ (.A0(\logix.ram_r[219] ),
    .A1(\logix.ram_r[218] ),
    .S(net308),
    .X(_1195_));
 sg13g2_mux2_1 _7335_ (.A0(\logix.ram_r[21] ),
    .A1(\logix.ram_r[20] ),
    .S(_2213_),
    .X(_1196_));
 sg13g2_buf_1 _7336_ (.A(_2202_),
    .X(_2214_));
 sg13g2_mux2_1 _7337_ (.A0(\logix.ram_r[220] ),
    .A1(\logix.ram_r[219] ),
    .S(net307),
    .X(_1197_));
 sg13g2_mux2_1 _7338_ (.A0(\logix.ram_r[221] ),
    .A1(\logix.ram_r[220] ),
    .S(net307),
    .X(_1198_));
 sg13g2_mux2_1 _7339_ (.A0(\logix.ram_r[222] ),
    .A1(\logix.ram_r[221] ),
    .S(_2214_),
    .X(_1199_));
 sg13g2_mux2_1 _7340_ (.A0(\logix.ram_r[223] ),
    .A1(\logix.ram_r[222] ),
    .S(_2214_),
    .X(_1200_));
 sg13g2_mux2_1 _7341_ (.A0(\logix.ram_r[224] ),
    .A1(\logix.ram_r[223] ),
    .S(net307),
    .X(_1201_));
 sg13g2_mux2_1 _7342_ (.A0(\logix.ram_r[225] ),
    .A1(\logix.ram_r[224] ),
    .S(net307),
    .X(_1202_));
 sg13g2_mux2_1 _7343_ (.A0(\logix.ram_r[226] ),
    .A1(\logix.ram_r[225] ),
    .S(net307),
    .X(_1203_));
 sg13g2_mux2_1 _7344_ (.A0(\logix.ram_r[227] ),
    .A1(\logix.ram_r[226] ),
    .S(net307),
    .X(_1204_));
 sg13g2_mux2_1 _7345_ (.A0(\logix.ram_r[228] ),
    .A1(\logix.ram_r[227] ),
    .S(net307),
    .X(_1205_));
 sg13g2_mux2_1 _7346_ (.A0(\logix.ram_r[229] ),
    .A1(\logix.ram_r[228] ),
    .S(net307),
    .X(_1206_));
 sg13g2_buf_1 _7347_ (.A(_2202_),
    .X(_2215_));
 sg13g2_mux2_1 _7348_ (.A0(\logix.ram_r[22] ),
    .A1(\logix.ram_r[21] ),
    .S(_2215_),
    .X(_1207_));
 sg13g2_mux2_1 _7349_ (.A0(\logix.ram_r[230] ),
    .A1(\logix.ram_r[229] ),
    .S(net306),
    .X(_1208_));
 sg13g2_mux2_1 _7350_ (.A0(\logix.ram_r[231] ),
    .A1(\logix.ram_r[230] ),
    .S(_2215_),
    .X(_1209_));
 sg13g2_mux2_1 _7351_ (.A0(\logix.ram_r[232] ),
    .A1(\logix.ram_r[231] ),
    .S(net306),
    .X(_1210_));
 sg13g2_mux2_1 _7352_ (.A0(\logix.ram_r[233] ),
    .A1(\logix.ram_r[232] ),
    .S(net306),
    .X(_1211_));
 sg13g2_mux2_1 _7353_ (.A0(\logix.ram_r[234] ),
    .A1(\logix.ram_r[233] ),
    .S(net306),
    .X(_1212_));
 sg13g2_mux2_1 _7354_ (.A0(\logix.ram_r[235] ),
    .A1(\logix.ram_r[234] ),
    .S(net306),
    .X(_1213_));
 sg13g2_mux2_1 _7355_ (.A0(\logix.ram_r[236] ),
    .A1(\logix.ram_r[235] ),
    .S(net306),
    .X(_1214_));
 sg13g2_mux2_1 _7356_ (.A0(\logix.ram_r[237] ),
    .A1(\logix.ram_r[236] ),
    .S(net306),
    .X(_1215_));
 sg13g2_mux2_1 _7357_ (.A0(\logix.ram_r[238] ),
    .A1(\logix.ram_r[237] ),
    .S(net306),
    .X(_1216_));
 sg13g2_buf_1 _7358_ (.A(_2202_),
    .X(_2216_));
 sg13g2_mux2_1 _7359_ (.A0(\logix.ram_r[239] ),
    .A1(\logix.ram_r[238] ),
    .S(_2216_),
    .X(_1217_));
 sg13g2_mux2_1 _7360_ (.A0(\logix.ram_r[23] ),
    .A1(\logix.ram_r[22] ),
    .S(_2216_),
    .X(_1218_));
 sg13g2_mux2_1 _7361_ (.A0(\logix.ram_r[240] ),
    .A1(\logix.ram_r[239] ),
    .S(net305),
    .X(_1219_));
 sg13g2_mux2_1 _7362_ (.A0(\logix.ram_r[241] ),
    .A1(\logix.ram_r[240] ),
    .S(net305),
    .X(_1220_));
 sg13g2_mux2_1 _7363_ (.A0(\logix.ram_r[242] ),
    .A1(\logix.ram_r[241] ),
    .S(net305),
    .X(_1221_));
 sg13g2_mux2_1 _7364_ (.A0(\logix.ram_r[243] ),
    .A1(\logix.ram_r[242] ),
    .S(net305),
    .X(_1222_));
 sg13g2_mux2_1 _7365_ (.A0(\logix.ram_r[244] ),
    .A1(\logix.ram_r[243] ),
    .S(net305),
    .X(_1223_));
 sg13g2_mux2_1 _7366_ (.A0(\logix.ram_r[245] ),
    .A1(\logix.ram_r[244] ),
    .S(net305),
    .X(_1224_));
 sg13g2_mux2_1 _7367_ (.A0(\logix.ram_r[246] ),
    .A1(\logix.ram_r[245] ),
    .S(net305),
    .X(_1225_));
 sg13g2_mux2_1 _7368_ (.A0(\logix.ram_r[247] ),
    .A1(\logix.ram_r[246] ),
    .S(net305),
    .X(_1226_));
 sg13g2_buf_1 _7369_ (.A(_2202_),
    .X(_2217_));
 sg13g2_mux2_1 _7370_ (.A0(\logix.ram_r[248] ),
    .A1(\logix.ram_r[247] ),
    .S(net304),
    .X(_1227_));
 sg13g2_mux2_1 _7371_ (.A0(\logix.ram_r[249] ),
    .A1(\logix.ram_r[248] ),
    .S(net304),
    .X(_1228_));
 sg13g2_mux2_1 _7372_ (.A0(\logix.ram_r[24] ),
    .A1(\logix.ram_r[23] ),
    .S(_2217_),
    .X(_1229_));
 sg13g2_mux2_1 _7373_ (.A0(\logix.ram_r[250] ),
    .A1(\logix.ram_r[249] ),
    .S(net304),
    .X(_1230_));
 sg13g2_mux2_1 _7374_ (.A0(\logix.ram_r[251] ),
    .A1(\logix.ram_r[250] ),
    .S(net304),
    .X(_1231_));
 sg13g2_mux2_1 _7375_ (.A0(\logix.ram_r[252] ),
    .A1(\logix.ram_r[251] ),
    .S(net304),
    .X(_1232_));
 sg13g2_mux2_1 _7376_ (.A0(\logix.ram_r[253] ),
    .A1(\logix.ram_r[252] ),
    .S(net304),
    .X(_1233_));
 sg13g2_mux2_1 _7377_ (.A0(\logix.ram_r[254] ),
    .A1(\logix.ram_r[253] ),
    .S(net304),
    .X(_1234_));
 sg13g2_mux2_1 _7378_ (.A0(\logix.ram_r[255] ),
    .A1(\logix.ram_r[254] ),
    .S(net304),
    .X(_1235_));
 sg13g2_mux2_1 _7379_ (.A0(\logix.ram_r[256] ),
    .A1(\logix.ram_r[255] ),
    .S(_2217_),
    .X(_1236_));
 sg13g2_buf_1 _7380_ (.A(_2201_),
    .X(_2218_));
 sg13g2_buf_1 _7381_ (.A(_2218_),
    .X(_2219_));
 sg13g2_mux2_1 _7382_ (.A0(\logix.ram_r[257] ),
    .A1(\logix.ram_r[256] ),
    .S(net303),
    .X(_1237_));
 sg13g2_mux2_1 _7383_ (.A0(\logix.ram_r[258] ),
    .A1(\logix.ram_r[257] ),
    .S(net303),
    .X(_1238_));
 sg13g2_mux2_1 _7384_ (.A0(\logix.ram_r[259] ),
    .A1(\logix.ram_r[258] ),
    .S(net303),
    .X(_1239_));
 sg13g2_mux2_1 _7385_ (.A0(\logix.ram_r[25] ),
    .A1(\logix.ram_r[24] ),
    .S(net303),
    .X(_1240_));
 sg13g2_mux2_1 _7386_ (.A0(\logix.ram_r[260] ),
    .A1(\logix.ram_r[259] ),
    .S(net303),
    .X(_1241_));
 sg13g2_mux2_1 _7387_ (.A0(\logix.ram_r[261] ),
    .A1(\logix.ram_r[260] ),
    .S(net303),
    .X(_1242_));
 sg13g2_mux2_1 _7388_ (.A0(\logix.ram_r[262] ),
    .A1(\logix.ram_r[261] ),
    .S(_2219_),
    .X(_1243_));
 sg13g2_mux2_1 _7389_ (.A0(\logix.ram_r[263] ),
    .A1(\logix.ram_r[262] ),
    .S(_2219_),
    .X(_1244_));
 sg13g2_mux2_1 _7390_ (.A0(\logix.ram_r[264] ),
    .A1(\logix.ram_r[263] ),
    .S(net303),
    .X(_1245_));
 sg13g2_mux2_1 _7391_ (.A0(\logix.ram_r[265] ),
    .A1(\logix.ram_r[264] ),
    .S(net303),
    .X(_1246_));
 sg13g2_buf_1 _7392_ (.A(_2218_),
    .X(_2220_));
 sg13g2_mux2_1 _7393_ (.A0(\logix.ram_r[266] ),
    .A1(\logix.ram_r[265] ),
    .S(net302),
    .X(_1247_));
 sg13g2_mux2_1 _7394_ (.A0(\logix.ram_r[267] ),
    .A1(\logix.ram_r[266] ),
    .S(net302),
    .X(_1248_));
 sg13g2_mux2_1 _7395_ (.A0(\logix.ram_r[268] ),
    .A1(\logix.ram_r[267] ),
    .S(_2220_),
    .X(_1249_));
 sg13g2_mux2_1 _7396_ (.A0(\logix.ram_r[269] ),
    .A1(\logix.ram_r[268] ),
    .S(net302),
    .X(_1250_));
 sg13g2_mux2_1 _7397_ (.A0(\logix.ram_r[26] ),
    .A1(\logix.ram_r[25] ),
    .S(net302),
    .X(_1251_));
 sg13g2_mux2_1 _7398_ (.A0(\logix.ram_r[270] ),
    .A1(\logix.ram_r[269] ),
    .S(net302),
    .X(_1252_));
 sg13g2_mux2_1 _7399_ (.A0(\logix.ram_r[271] ),
    .A1(\logix.ram_r[270] ),
    .S(net302),
    .X(_1253_));
 sg13g2_mux2_1 _7400_ (.A0(\logix.ram_r[272] ),
    .A1(\logix.ram_r[271] ),
    .S(net302),
    .X(_1254_));
 sg13g2_mux2_1 _7401_ (.A0(\logix.ram_r[273] ),
    .A1(\logix.ram_r[272] ),
    .S(net302),
    .X(_1255_));
 sg13g2_mux2_1 _7402_ (.A0(\logix.ram_r[274] ),
    .A1(\logix.ram_r[273] ),
    .S(_2220_),
    .X(_1256_));
 sg13g2_buf_1 _7403_ (.A(_2218_),
    .X(_2221_));
 sg13g2_mux2_1 _7404_ (.A0(\logix.ram_r[275] ),
    .A1(\logix.ram_r[274] ),
    .S(net301),
    .X(_1257_));
 sg13g2_mux2_1 _7405_ (.A0(\logix.ram_r[276] ),
    .A1(\logix.ram_r[275] ),
    .S(net301),
    .X(_1258_));
 sg13g2_mux2_1 _7406_ (.A0(\logix.ram_r[277] ),
    .A1(\logix.ram_r[276] ),
    .S(net301),
    .X(_1259_));
 sg13g2_mux2_1 _7407_ (.A0(\logix.ram_r[278] ),
    .A1(\logix.ram_r[277] ),
    .S(_2221_),
    .X(_1260_));
 sg13g2_mux2_1 _7408_ (.A0(\logix.ram_r[279] ),
    .A1(\logix.ram_r[278] ),
    .S(_2221_),
    .X(_1261_));
 sg13g2_mux2_1 _7409_ (.A0(\logix.ram_r[27] ),
    .A1(\logix.ram_r[26] ),
    .S(net301),
    .X(_1262_));
 sg13g2_mux2_1 _7410_ (.A0(\logix.ram_r[280] ),
    .A1(\logix.ram_r[279] ),
    .S(net301),
    .X(_1263_));
 sg13g2_mux2_1 _7411_ (.A0(\logix.ram_r[281] ),
    .A1(\logix.ram_r[280] ),
    .S(net301),
    .X(_1264_));
 sg13g2_mux2_1 _7412_ (.A0(\logix.ram_r[282] ),
    .A1(\logix.ram_r[281] ),
    .S(net301),
    .X(_1265_));
 sg13g2_mux2_1 _7413_ (.A0(\logix.ram_r[283] ),
    .A1(\logix.ram_r[282] ),
    .S(net301),
    .X(_1266_));
 sg13g2_buf_1 _7414_ (.A(_2218_),
    .X(_2222_));
 sg13g2_mux2_1 _7415_ (.A0(\logix.ram_r[284] ),
    .A1(\logix.ram_r[283] ),
    .S(_2222_),
    .X(_1267_));
 sg13g2_mux2_1 _7416_ (.A0(\logix.ram_r[285] ),
    .A1(\logix.ram_r[284] ),
    .S(net300),
    .X(_1268_));
 sg13g2_mux2_1 _7417_ (.A0(\logix.ram_r[286] ),
    .A1(\logix.ram_r[285] ),
    .S(net300),
    .X(_1269_));
 sg13g2_mux2_1 _7418_ (.A0(\logix.ram_r[287] ),
    .A1(\logix.ram_r[286] ),
    .S(net300),
    .X(_1270_));
 sg13g2_mux2_1 _7419_ (.A0(\logix.ram_r[288] ),
    .A1(\logix.ram_r[287] ),
    .S(net300),
    .X(_1271_));
 sg13g2_mux2_1 _7420_ (.A0(\logix.ram_r[289] ),
    .A1(\logix.ram_r[288] ),
    .S(net300),
    .X(_1272_));
 sg13g2_mux2_1 _7421_ (.A0(\logix.ram_r[28] ),
    .A1(\logix.ram_r[27] ),
    .S(net300),
    .X(_1273_));
 sg13g2_mux2_1 _7422_ (.A0(\logix.ram_r[290] ),
    .A1(\logix.ram_r[289] ),
    .S(net300),
    .X(_1274_));
 sg13g2_mux2_1 _7423_ (.A0(\logix.ram_r[291] ),
    .A1(\logix.ram_r[290] ),
    .S(net300),
    .X(_1275_));
 sg13g2_mux2_1 _7424_ (.A0(\logix.ram_r[292] ),
    .A1(\logix.ram_r[291] ),
    .S(_2222_),
    .X(_1276_));
 sg13g2_buf_1 _7425_ (.A(_2218_),
    .X(_2223_));
 sg13g2_mux2_1 _7426_ (.A0(\logix.ram_r[293] ),
    .A1(\logix.ram_r[292] ),
    .S(net299),
    .X(_1277_));
 sg13g2_mux2_1 _7427_ (.A0(\logix.ram_r[294] ),
    .A1(\logix.ram_r[293] ),
    .S(net299),
    .X(_1278_));
 sg13g2_mux2_1 _7428_ (.A0(\logix.ram_r[295] ),
    .A1(\logix.ram_r[294] ),
    .S(net299),
    .X(_1279_));
 sg13g2_mux2_1 _7429_ (.A0(\logix.ram_r[296] ),
    .A1(\logix.ram_r[295] ),
    .S(net299),
    .X(_1280_));
 sg13g2_mux2_1 _7430_ (.A0(\logix.ram_r[297] ),
    .A1(\logix.ram_r[296] ),
    .S(net299),
    .X(_1281_));
 sg13g2_mux2_1 _7431_ (.A0(\logix.ram_r[298] ),
    .A1(\logix.ram_r[297] ),
    .S(net299),
    .X(_1282_));
 sg13g2_mux2_1 _7432_ (.A0(\logix.ram_r[299] ),
    .A1(\logix.ram_r[298] ),
    .S(_2223_),
    .X(_1283_));
 sg13g2_mux2_1 _7433_ (.A0(\logix.ram_r[29] ),
    .A1(\logix.ram_r[28] ),
    .S(net299),
    .X(_1284_));
 sg13g2_mux2_1 _7434_ (.A0(\logix.ram_r[2] ),
    .A1(\logix.ram_r[1] ),
    .S(net299),
    .X(_1285_));
 sg13g2_mux2_1 _7435_ (.A0(\logix.ram_r[300] ),
    .A1(\logix.ram_r[299] ),
    .S(_2223_),
    .X(_1286_));
 sg13g2_buf_1 _7436_ (.A(_2218_),
    .X(_2224_));
 sg13g2_mux2_1 _7437_ (.A0(\logix.ram_r[301] ),
    .A1(\logix.ram_r[300] ),
    .S(net298),
    .X(_1287_));
 sg13g2_mux2_1 _7438_ (.A0(\logix.ram_r[302] ),
    .A1(\logix.ram_r[301] ),
    .S(net298),
    .X(_1288_));
 sg13g2_mux2_1 _7439_ (.A0(\logix.ram_r[303] ),
    .A1(\logix.ram_r[302] ),
    .S(net298),
    .X(_1289_));
 sg13g2_mux2_1 _7440_ (.A0(\logix.ram_r[304] ),
    .A1(\logix.ram_r[303] ),
    .S(net298),
    .X(_1290_));
 sg13g2_mux2_1 _7441_ (.A0(\logix.ram_r[305] ),
    .A1(\logix.ram_r[304] ),
    .S(net298),
    .X(_1291_));
 sg13g2_mux2_1 _7442_ (.A0(\logix.ram_r[306] ),
    .A1(\logix.ram_r[305] ),
    .S(net298),
    .X(_1292_));
 sg13g2_mux2_1 _7443_ (.A0(\logix.ram_r[307] ),
    .A1(\logix.ram_r[306] ),
    .S(net298),
    .X(_1293_));
 sg13g2_mux2_1 _7444_ (.A0(\logix.ram_r[308] ),
    .A1(\logix.ram_r[307] ),
    .S(_2224_),
    .X(_1294_));
 sg13g2_mux2_1 _7445_ (.A0(\logix.ram_r[309] ),
    .A1(\logix.ram_r[308] ),
    .S(_2224_),
    .X(_1295_));
 sg13g2_mux2_1 _7446_ (.A0(\logix.ram_r[30] ),
    .A1(\logix.ram_r[29] ),
    .S(net298),
    .X(_1296_));
 sg13g2_buf_1 _7447_ (.A(_2218_),
    .X(_2225_));
 sg13g2_mux2_1 _7448_ (.A0(\logix.ram_r[310] ),
    .A1(\logix.ram_r[309] ),
    .S(net297),
    .X(_1297_));
 sg13g2_mux2_1 _7449_ (.A0(\logix.ram_r[311] ),
    .A1(\logix.ram_r[310] ),
    .S(net297),
    .X(_1298_));
 sg13g2_mux2_1 _7450_ (.A0(\logix.ram_r[312] ),
    .A1(\logix.ram_r[311] ),
    .S(net297),
    .X(_1299_));
 sg13g2_mux2_1 _7451_ (.A0(\logix.ram_r[313] ),
    .A1(\logix.ram_r[312] ),
    .S(net297),
    .X(_1300_));
 sg13g2_mux2_1 _7452_ (.A0(\logix.ram_r[314] ),
    .A1(\logix.ram_r[313] ),
    .S(_2225_),
    .X(_1301_));
 sg13g2_mux2_1 _7453_ (.A0(\logix.ram_r[315] ),
    .A1(\logix.ram_r[314] ),
    .S(net297),
    .X(_1302_));
 sg13g2_mux2_1 _7454_ (.A0(\logix.ram_r[316] ),
    .A1(\logix.ram_r[315] ),
    .S(net297),
    .X(_1303_));
 sg13g2_mux2_1 _7455_ (.A0(\logix.ram_r[317] ),
    .A1(\logix.ram_r[316] ),
    .S(_2225_),
    .X(_1304_));
 sg13g2_mux2_1 _7456_ (.A0(\logix.ram_r[318] ),
    .A1(\logix.ram_r[317] ),
    .S(net297),
    .X(_1305_));
 sg13g2_mux2_1 _7457_ (.A0(\logix.ram_r[319] ),
    .A1(\logix.ram_r[318] ),
    .S(net297),
    .X(_1306_));
 sg13g2_buf_1 _7458_ (.A(_2201_),
    .X(_2226_));
 sg13g2_buf_1 _7459_ (.A(_2226_),
    .X(_2227_));
 sg13g2_mux2_1 _7460_ (.A0(\logix.ram_r[31] ),
    .A1(\logix.ram_r[30] ),
    .S(net296),
    .X(_1307_));
 sg13g2_mux2_1 _7461_ (.A0(\logix.ram_r[320] ),
    .A1(\logix.ram_r[319] ),
    .S(net296),
    .X(_1308_));
 sg13g2_mux2_1 _7462_ (.A0(\logix.ram_r[321] ),
    .A1(\logix.ram_r[320] ),
    .S(net296),
    .X(_1309_));
 sg13g2_mux2_1 _7463_ (.A0(\logix.ram_r[322] ),
    .A1(\logix.ram_r[321] ),
    .S(net296),
    .X(_1310_));
 sg13g2_mux2_1 _7464_ (.A0(\logix.ram_r[323] ),
    .A1(\logix.ram_r[322] ),
    .S(net296),
    .X(_1311_));
 sg13g2_mux2_1 _7465_ (.A0(\logix.ram_r[324] ),
    .A1(\logix.ram_r[323] ),
    .S(net296),
    .X(_1312_));
 sg13g2_mux2_1 _7466_ (.A0(\logix.ram_r[325] ),
    .A1(\logix.ram_r[324] ),
    .S(_2227_),
    .X(_1313_));
 sg13g2_mux2_1 _7467_ (.A0(\logix.ram_r[326] ),
    .A1(\logix.ram_r[325] ),
    .S(net296),
    .X(_1314_));
 sg13g2_mux2_1 _7468_ (.A0(\logix.ram_r[327] ),
    .A1(\logix.ram_r[326] ),
    .S(net296),
    .X(_1315_));
 sg13g2_mux2_1 _7469_ (.A0(\logix.ram_r[328] ),
    .A1(\logix.ram_r[327] ),
    .S(_2227_),
    .X(_1316_));
 sg13g2_buf_1 _7470_ (.A(_2226_),
    .X(_2228_));
 sg13g2_mux2_1 _7471_ (.A0(\logix.ram_r[329] ),
    .A1(\logix.ram_r[328] ),
    .S(_2228_),
    .X(_1317_));
 sg13g2_mux2_1 _7472_ (.A0(\logix.ram_r[32] ),
    .A1(\logix.ram_r[31] ),
    .S(net295),
    .X(_1318_));
 sg13g2_mux2_1 _7473_ (.A0(\logix.ram_r[330] ),
    .A1(\logix.ram_r[329] ),
    .S(net295),
    .X(_1319_));
 sg13g2_mux2_1 _7474_ (.A0(\logix.ram_r[331] ),
    .A1(\logix.ram_r[330] ),
    .S(net295),
    .X(_1320_));
 sg13g2_mux2_1 _7475_ (.A0(\logix.ram_r[332] ),
    .A1(\logix.ram_r[331] ),
    .S(net295),
    .X(_1321_));
 sg13g2_mux2_1 _7476_ (.A0(\logix.ram_r[333] ),
    .A1(\logix.ram_r[332] ),
    .S(net295),
    .X(_1322_));
 sg13g2_mux2_1 _7477_ (.A0(\logix.ram_r[334] ),
    .A1(\logix.ram_r[333] ),
    .S(net295),
    .X(_1323_));
 sg13g2_mux2_1 _7478_ (.A0(\logix.ram_r[335] ),
    .A1(\logix.ram_r[334] ),
    .S(net295),
    .X(_1324_));
 sg13g2_mux2_1 _7479_ (.A0(\logix.ram_r[336] ),
    .A1(\logix.ram_r[335] ),
    .S(_2228_),
    .X(_1325_));
 sg13g2_mux2_1 _7480_ (.A0(\logix.ram_r[337] ),
    .A1(\logix.ram_r[336] ),
    .S(net295),
    .X(_1326_));
 sg13g2_buf_1 _7481_ (.A(_2226_),
    .X(_2229_));
 sg13g2_mux2_1 _7482_ (.A0(\logix.ram_r[338] ),
    .A1(\logix.ram_r[337] ),
    .S(net294),
    .X(_1327_));
 sg13g2_mux2_1 _7483_ (.A0(\logix.ram_r[339] ),
    .A1(\logix.ram_r[338] ),
    .S(net294),
    .X(_1328_));
 sg13g2_mux2_1 _7484_ (.A0(\logix.ram_r[33] ),
    .A1(\logix.ram_r[32] ),
    .S(net294),
    .X(_1329_));
 sg13g2_mux2_1 _7485_ (.A0(\logix.ram_r[340] ),
    .A1(\logix.ram_r[339] ),
    .S(net294),
    .X(_1330_));
 sg13g2_mux2_1 _7486_ (.A0(\logix.ram_r[341] ),
    .A1(\logix.ram_r[340] ),
    .S(net294),
    .X(_1331_));
 sg13g2_mux2_1 _7487_ (.A0(\logix.ram_r[342] ),
    .A1(\logix.ram_r[341] ),
    .S(net294),
    .X(_1332_));
 sg13g2_mux2_1 _7488_ (.A0(\logix.ram_r[343] ),
    .A1(\logix.ram_r[342] ),
    .S(net294),
    .X(_1333_));
 sg13g2_mux2_1 _7489_ (.A0(\logix.ram_r[344] ),
    .A1(\logix.ram_r[343] ),
    .S(_2229_),
    .X(_1334_));
 sg13g2_mux2_1 _7490_ (.A0(\logix.ram_r[345] ),
    .A1(\logix.ram_r[344] ),
    .S(_2229_),
    .X(_1335_));
 sg13g2_mux2_1 _7491_ (.A0(\logix.ram_r[346] ),
    .A1(\logix.ram_r[345] ),
    .S(net294),
    .X(_1336_));
 sg13g2_buf_1 _7492_ (.A(_2226_),
    .X(_2230_));
 sg13g2_mux2_1 _7493_ (.A0(\logix.ram_r[347] ),
    .A1(\logix.ram_r[346] ),
    .S(net293),
    .X(_1337_));
 sg13g2_mux2_1 _7494_ (.A0(\logix.ram_r[348] ),
    .A1(\logix.ram_r[347] ),
    .S(net293),
    .X(_1338_));
 sg13g2_mux2_1 _7495_ (.A0(\logix.ram_r[349] ),
    .A1(\logix.ram_r[348] ),
    .S(net293),
    .X(_1339_));
 sg13g2_mux2_1 _7496_ (.A0(\logix.ram_r[34] ),
    .A1(\logix.ram_r[33] ),
    .S(net293),
    .X(_1340_));
 sg13g2_mux2_1 _7497_ (.A0(\logix.ram_r[350] ),
    .A1(\logix.ram_r[349] ),
    .S(_2230_),
    .X(_1341_));
 sg13g2_mux2_1 _7498_ (.A0(\logix.ram_r[351] ),
    .A1(\logix.ram_r[350] ),
    .S(net293),
    .X(_1342_));
 sg13g2_mux2_1 _7499_ (.A0(\logix.ram_r[352] ),
    .A1(\logix.ram_r[351] ),
    .S(net293),
    .X(_1343_));
 sg13g2_mux2_1 _7500_ (.A0(\logix.ram_r[353] ),
    .A1(\logix.ram_r[352] ),
    .S(net293),
    .X(_1344_));
 sg13g2_mux2_1 _7501_ (.A0(\logix.ram_r[354] ),
    .A1(\logix.ram_r[353] ),
    .S(_2230_),
    .X(_1345_));
 sg13g2_mux2_1 _7502_ (.A0(\logix.ram_r[355] ),
    .A1(\logix.ram_r[354] ),
    .S(net293),
    .X(_1346_));
 sg13g2_buf_1 _7503_ (.A(_2226_),
    .X(_2231_));
 sg13g2_mux2_1 _7504_ (.A0(\logix.ram_r[356] ),
    .A1(\logix.ram_r[355] ),
    .S(net292),
    .X(_1347_));
 sg13g2_mux2_1 _7505_ (.A0(\logix.ram_r[357] ),
    .A1(\logix.ram_r[356] ),
    .S(net292),
    .X(_1348_));
 sg13g2_mux2_1 _7506_ (.A0(\logix.ram_r[358] ),
    .A1(\logix.ram_r[357] ),
    .S(net292),
    .X(_1349_));
 sg13g2_mux2_1 _7507_ (.A0(\logix.ram_r[359] ),
    .A1(\logix.ram_r[358] ),
    .S(net292),
    .X(_1350_));
 sg13g2_mux2_1 _7508_ (.A0(\logix.ram_r[35] ),
    .A1(\logix.ram_r[34] ),
    .S(_2231_),
    .X(_1351_));
 sg13g2_mux2_1 _7509_ (.A0(\logix.ram_r[360] ),
    .A1(\logix.ram_r[359] ),
    .S(net292),
    .X(_1352_));
 sg13g2_mux2_1 _7510_ (.A0(\logix.ram_r[361] ),
    .A1(\logix.ram_r[360] ),
    .S(net292),
    .X(_1353_));
 sg13g2_mux2_1 _7511_ (.A0(\logix.ram_r[362] ),
    .A1(\logix.ram_r[361] ),
    .S(net292),
    .X(_1354_));
 sg13g2_mux2_1 _7512_ (.A0(\logix.ram_r[363] ),
    .A1(\logix.ram_r[362] ),
    .S(net292),
    .X(_1355_));
 sg13g2_mux2_1 _7513_ (.A0(\logix.ram_r[364] ),
    .A1(\logix.ram_r[363] ),
    .S(_2231_),
    .X(_1356_));
 sg13g2_buf_1 _7514_ (.A(_2226_),
    .X(_2232_));
 sg13g2_mux2_1 _7515_ (.A0(\logix.ram_r[365] ),
    .A1(\logix.ram_r[364] ),
    .S(net291),
    .X(_1357_));
 sg13g2_mux2_1 _7516_ (.A0(\logix.ram_r[366] ),
    .A1(\logix.ram_r[365] ),
    .S(net291),
    .X(_1358_));
 sg13g2_mux2_1 _7517_ (.A0(\logix.ram_r[367] ),
    .A1(\logix.ram_r[366] ),
    .S(net291),
    .X(_1359_));
 sg13g2_mux2_1 _7518_ (.A0(\logix.ram_r[368] ),
    .A1(\logix.ram_r[367] ),
    .S(net291),
    .X(_1360_));
 sg13g2_mux2_1 _7519_ (.A0(\logix.ram_r[369] ),
    .A1(\logix.ram_r[368] ),
    .S(_2232_),
    .X(_1361_));
 sg13g2_mux2_1 _7520_ (.A0(\logix.ram_r[36] ),
    .A1(\logix.ram_r[35] ),
    .S(_2232_),
    .X(_1362_));
 sg13g2_mux2_1 _7521_ (.A0(\logix.ram_r[370] ),
    .A1(\logix.ram_r[369] ),
    .S(net291),
    .X(_1363_));
 sg13g2_mux2_1 _7522_ (.A0(\logix.ram_r[371] ),
    .A1(\logix.ram_r[370] ),
    .S(net291),
    .X(_1364_));
 sg13g2_mux2_1 _7523_ (.A0(\logix.ram_r[372] ),
    .A1(\logix.ram_r[371] ),
    .S(net291),
    .X(_1365_));
 sg13g2_mux2_1 _7524_ (.A0(\logix.ram_r[373] ),
    .A1(\logix.ram_r[372] ),
    .S(net291),
    .X(_1366_));
 sg13g2_buf_1 _7525_ (.A(_2226_),
    .X(_2233_));
 sg13g2_mux2_1 _7526_ (.A0(\logix.ram_r[374] ),
    .A1(\logix.ram_r[373] ),
    .S(net290),
    .X(_1367_));
 sg13g2_mux2_1 _7527_ (.A0(\logix.ram_r[375] ),
    .A1(\logix.ram_r[374] ),
    .S(net290),
    .X(_1368_));
 sg13g2_mux2_1 _7528_ (.A0(\logix.ram_r[376] ),
    .A1(\logix.ram_r[375] ),
    .S(net290),
    .X(_1369_));
 sg13g2_mux2_1 _7529_ (.A0(\logix.ram_r[377] ),
    .A1(\logix.ram_r[376] ),
    .S(net290),
    .X(_1370_));
 sg13g2_mux2_1 _7530_ (.A0(\logix.ram_r[378] ),
    .A1(\logix.ram_r[377] ),
    .S(net290),
    .X(_1371_));
 sg13g2_mux2_1 _7531_ (.A0(\logix.ram_r[379] ),
    .A1(\logix.ram_r[378] ),
    .S(_2233_),
    .X(_1372_));
 sg13g2_mux2_1 _7532_ (.A0(\logix.ram_r[37] ),
    .A1(\logix.ram_r[36] ),
    .S(net290),
    .X(_1373_));
 sg13g2_mux2_1 _7533_ (.A0(\logix.ram_r[380] ),
    .A1(\logix.ram_r[379] ),
    .S(_2233_),
    .X(_1374_));
 sg13g2_mux2_1 _7534_ (.A0(\logix.ram_r[381] ),
    .A1(\logix.ram_r[380] ),
    .S(net290),
    .X(_1375_));
 sg13g2_mux2_1 _7535_ (.A0(\logix.ram_r[382] ),
    .A1(\logix.ram_r[381] ),
    .S(net290),
    .X(_1376_));
 sg13g2_buf_1 _7536_ (.A(_2201_),
    .X(_2234_));
 sg13g2_buf_1 _7537_ (.A(_2234_),
    .X(_2235_));
 sg13g2_mux2_1 _7538_ (.A0(\logix.ram_r[383] ),
    .A1(\logix.ram_r[382] ),
    .S(_2235_),
    .X(_1377_));
 sg13g2_mux2_1 _7539_ (.A0(\logix.ram_r[384] ),
    .A1(\logix.ram_r[383] ),
    .S(net289),
    .X(_1378_));
 sg13g2_mux2_1 _7540_ (.A0(\logix.ram_r[385] ),
    .A1(\logix.ram_r[384] ),
    .S(net289),
    .X(_1379_));
 sg13g2_mux2_1 _7541_ (.A0(\logix.ram_r[386] ),
    .A1(\logix.ram_r[385] ),
    .S(net289),
    .X(_1380_));
 sg13g2_mux2_1 _7542_ (.A0(\logix.ram_r[387] ),
    .A1(\logix.ram_r[386] ),
    .S(net289),
    .X(_1381_));
 sg13g2_mux2_1 _7543_ (.A0(\logix.ram_r[388] ),
    .A1(\logix.ram_r[387] ),
    .S(net289),
    .X(_1382_));
 sg13g2_mux2_1 _7544_ (.A0(\logix.ram_r[389] ),
    .A1(\logix.ram_r[388] ),
    .S(net289),
    .X(_1383_));
 sg13g2_mux2_1 _7545_ (.A0(\logix.ram_r[38] ),
    .A1(\logix.ram_r[37] ),
    .S(_2235_),
    .X(_1384_));
 sg13g2_mux2_1 _7546_ (.A0(\logix.ram_r[390] ),
    .A1(\logix.ram_r[389] ),
    .S(net289),
    .X(_1385_));
 sg13g2_mux2_1 _7547_ (.A0(\logix.ram_r[391] ),
    .A1(\logix.ram_r[390] ),
    .S(net289),
    .X(_1386_));
 sg13g2_buf_1 _7548_ (.A(_2234_),
    .X(_2236_));
 sg13g2_mux2_1 _7549_ (.A0(\logix.ram_r[392] ),
    .A1(\logix.ram_r[391] ),
    .S(net288),
    .X(_1387_));
 sg13g2_mux2_1 _7550_ (.A0(\logix.ram_r[393] ),
    .A1(\logix.ram_r[392] ),
    .S(net288),
    .X(_1388_));
 sg13g2_mux2_1 _7551_ (.A0(\logix.ram_r[394] ),
    .A1(\logix.ram_r[393] ),
    .S(net288),
    .X(_1389_));
 sg13g2_mux2_1 _7552_ (.A0(\logix.ram_r[395] ),
    .A1(\logix.ram_r[394] ),
    .S(net288),
    .X(_1390_));
 sg13g2_mux2_1 _7553_ (.A0(\logix.ram_r[396] ),
    .A1(\logix.ram_r[395] ),
    .S(net288),
    .X(_1391_));
 sg13g2_mux2_1 _7554_ (.A0(\logix.ram_r[397] ),
    .A1(\logix.ram_r[396] ),
    .S(net288),
    .X(_1392_));
 sg13g2_mux2_1 _7555_ (.A0(\logix.ram_r[398] ),
    .A1(\logix.ram_r[397] ),
    .S(net288),
    .X(_1393_));
 sg13g2_mux2_1 _7556_ (.A0(\logix.ram_r[399] ),
    .A1(\logix.ram_r[398] ),
    .S(net288),
    .X(_1394_));
 sg13g2_mux2_1 _7557_ (.A0(\logix.ram_r[39] ),
    .A1(\logix.ram_r[38] ),
    .S(_2236_),
    .X(_1395_));
 sg13g2_mux2_1 _7558_ (.A0(\logix.ram_r[3] ),
    .A1(\logix.ram_r[2] ),
    .S(_2236_),
    .X(_1396_));
 sg13g2_buf_1 _7559_ (.A(_2234_),
    .X(_2237_));
 sg13g2_mux2_1 _7560_ (.A0(\logix.ram_r[400] ),
    .A1(\logix.ram_r[399] ),
    .S(_2237_),
    .X(_1397_));
 sg13g2_mux2_1 _7561_ (.A0(\logix.ram_r[401] ),
    .A1(\logix.ram_r[400] ),
    .S(net287),
    .X(_1398_));
 sg13g2_mux2_1 _7562_ (.A0(\logix.ram_r[402] ),
    .A1(\logix.ram_r[401] ),
    .S(net287),
    .X(_1399_));
 sg13g2_mux2_1 _7563_ (.A0(\logix.ram_r[403] ),
    .A1(\logix.ram_r[402] ),
    .S(net287),
    .X(_1400_));
 sg13g2_mux2_1 _7564_ (.A0(\logix.ram_r[404] ),
    .A1(\logix.ram_r[403] ),
    .S(net287),
    .X(_1401_));
 sg13g2_mux2_1 _7565_ (.A0(\logix.ram_r[405] ),
    .A1(\logix.ram_r[404] ),
    .S(net287),
    .X(_1402_));
 sg13g2_mux2_1 _7566_ (.A0(\logix.ram_r[406] ),
    .A1(\logix.ram_r[405] ),
    .S(net287),
    .X(_1403_));
 sg13g2_mux2_1 _7567_ (.A0(\logix.ram_r[407] ),
    .A1(\logix.ram_r[406] ),
    .S(net287),
    .X(_1404_));
 sg13g2_mux2_1 _7568_ (.A0(\logix.ram_r[408] ),
    .A1(\logix.ram_r[407] ),
    .S(_2237_),
    .X(_1405_));
 sg13g2_mux2_1 _7569_ (.A0(\logix.ram_r[409] ),
    .A1(\logix.ram_r[408] ),
    .S(net287),
    .X(_1406_));
 sg13g2_buf_1 _7570_ (.A(_2234_),
    .X(_2238_));
 sg13g2_mux2_1 _7571_ (.A0(\logix.ram_r[40] ),
    .A1(\logix.ram_r[39] ),
    .S(_2238_),
    .X(_1407_));
 sg13g2_mux2_1 _7572_ (.A0(\logix.ram_r[410] ),
    .A1(\logix.ram_r[409] ),
    .S(_2238_),
    .X(_1408_));
 sg13g2_mux2_1 _7573_ (.A0(\logix.ram_r[411] ),
    .A1(\logix.ram_r[410] ),
    .S(net286),
    .X(_1409_));
 sg13g2_mux2_1 _7574_ (.A0(\logix.ram_r[412] ),
    .A1(\logix.ram_r[411] ),
    .S(net286),
    .X(_1410_));
 sg13g2_mux2_1 _7575_ (.A0(\logix.ram_r[413] ),
    .A1(\logix.ram_r[412] ),
    .S(net286),
    .X(_1411_));
 sg13g2_mux2_1 _7576_ (.A0(\logix.ram_r[414] ),
    .A1(\logix.ram_r[413] ),
    .S(net286),
    .X(_1412_));
 sg13g2_mux2_1 _7577_ (.A0(\logix.ram_r[415] ),
    .A1(\logix.ram_r[414] ),
    .S(net286),
    .X(_1413_));
 sg13g2_mux2_1 _7578_ (.A0(\logix.ram_r[416] ),
    .A1(\logix.ram_r[415] ),
    .S(net286),
    .X(_1414_));
 sg13g2_mux2_1 _7579_ (.A0(\logix.ram_r[417] ),
    .A1(\logix.ram_r[416] ),
    .S(net286),
    .X(_1415_));
 sg13g2_mux2_1 _7580_ (.A0(\logix.ram_r[418] ),
    .A1(\logix.ram_r[417] ),
    .S(net286),
    .X(_1416_));
 sg13g2_buf_1 _7581_ (.A(_2234_),
    .X(_2239_));
 sg13g2_mux2_1 _7582_ (.A0(\logix.ram_r[419] ),
    .A1(\logix.ram_r[418] ),
    .S(net285),
    .X(_1417_));
 sg13g2_mux2_1 _7583_ (.A0(\logix.ram_r[41] ),
    .A1(\logix.ram_r[40] ),
    .S(_2239_),
    .X(_1418_));
 sg13g2_mux2_1 _7584_ (.A0(\logix.ram_r[420] ),
    .A1(\logix.ram_r[419] ),
    .S(net285),
    .X(_1419_));
 sg13g2_mux2_1 _7585_ (.A0(\logix.ram_r[421] ),
    .A1(\logix.ram_r[420] ),
    .S(_2239_),
    .X(_1420_));
 sg13g2_mux2_1 _7586_ (.A0(\logix.ram_r[422] ),
    .A1(\logix.ram_r[421] ),
    .S(net285),
    .X(_1421_));
 sg13g2_mux2_1 _7587_ (.A0(\logix.ram_r[423] ),
    .A1(\logix.ram_r[422] ),
    .S(net285),
    .X(_1422_));
 sg13g2_mux2_1 _7588_ (.A0(\logix.ram_r[424] ),
    .A1(\logix.ram_r[423] ),
    .S(net285),
    .X(_1423_));
 sg13g2_mux2_1 _7589_ (.A0(\logix.ram_r[425] ),
    .A1(\logix.ram_r[424] ),
    .S(net285),
    .X(_1424_));
 sg13g2_mux2_1 _7590_ (.A0(\logix.ram_r[426] ),
    .A1(\logix.ram_r[425] ),
    .S(net285),
    .X(_1425_));
 sg13g2_mux2_1 _7591_ (.A0(\logix.ram_r[427] ),
    .A1(\logix.ram_r[426] ),
    .S(net285),
    .X(_1426_));
 sg13g2_buf_1 _7592_ (.A(_2234_),
    .X(_2240_));
 sg13g2_mux2_1 _7593_ (.A0(\logix.ram_r[428] ),
    .A1(\logix.ram_r[427] ),
    .S(net284),
    .X(_1427_));
 sg13g2_mux2_1 _7594_ (.A0(\logix.ram_r[429] ),
    .A1(\logix.ram_r[428] ),
    .S(net284),
    .X(_1428_));
 sg13g2_mux2_1 _7595_ (.A0(\logix.ram_r[42] ),
    .A1(\logix.ram_r[41] ),
    .S(_2240_),
    .X(_1429_));
 sg13g2_mux2_1 _7596_ (.A0(\logix.ram_r[430] ),
    .A1(\logix.ram_r[429] ),
    .S(net284),
    .X(_1430_));
 sg13g2_mux2_1 _7597_ (.A0(\logix.ram_r[431] ),
    .A1(\logix.ram_r[430] ),
    .S(net284),
    .X(_1431_));
 sg13g2_mux2_1 _7598_ (.A0(\logix.ram_r[432] ),
    .A1(\logix.ram_r[431] ),
    .S(net284),
    .X(_1432_));
 sg13g2_mux2_1 _7599_ (.A0(\logix.ram_r[433] ),
    .A1(\logix.ram_r[432] ),
    .S(net284),
    .X(_1433_));
 sg13g2_mux2_1 _7600_ (.A0(\logix.ram_r[434] ),
    .A1(\logix.ram_r[433] ),
    .S(net284),
    .X(_1434_));
 sg13g2_mux2_1 _7601_ (.A0(\logix.ram_r[435] ),
    .A1(\logix.ram_r[434] ),
    .S(net284),
    .X(_1435_));
 sg13g2_mux2_1 _7602_ (.A0(\logix.ram_r[436] ),
    .A1(\logix.ram_r[435] ),
    .S(_2240_),
    .X(_1436_));
 sg13g2_buf_1 _7603_ (.A(_2234_),
    .X(_2241_));
 sg13g2_mux2_1 _7604_ (.A0(\logix.ram_r[437] ),
    .A1(\logix.ram_r[436] ),
    .S(net283),
    .X(_1437_));
 sg13g2_mux2_1 _7605_ (.A0(\logix.ram_r[438] ),
    .A1(\logix.ram_r[437] ),
    .S(net283),
    .X(_1438_));
 sg13g2_mux2_1 _7606_ (.A0(\logix.ram_r[439] ),
    .A1(\logix.ram_r[438] ),
    .S(net283),
    .X(_1439_));
 sg13g2_mux2_1 _7607_ (.A0(\logix.ram_r[43] ),
    .A1(\logix.ram_r[42] ),
    .S(_2241_),
    .X(_1440_));
 sg13g2_mux2_1 _7608_ (.A0(\logix.ram_r[440] ),
    .A1(\logix.ram_r[439] ),
    .S(net283),
    .X(_1441_));
 sg13g2_mux2_1 _7609_ (.A0(\logix.ram_r[441] ),
    .A1(\logix.ram_r[440] ),
    .S(net283),
    .X(_1442_));
 sg13g2_mux2_1 _7610_ (.A0(\logix.ram_r[442] ),
    .A1(\logix.ram_r[441] ),
    .S(net283),
    .X(_1443_));
 sg13g2_mux2_1 _7611_ (.A0(\logix.ram_r[443] ),
    .A1(\logix.ram_r[442] ),
    .S(net283),
    .X(_1444_));
 sg13g2_mux2_1 _7612_ (.A0(\logix.ram_r[444] ),
    .A1(\logix.ram_r[443] ),
    .S(net283),
    .X(_1445_));
 sg13g2_mux2_1 _7613_ (.A0(\logix.ram_r[445] ),
    .A1(\logix.ram_r[444] ),
    .S(_2241_),
    .X(_1446_));
 sg13g2_buf_1 _7614_ (.A(_2201_),
    .X(_2242_));
 sg13g2_buf_1 _7615_ (.A(_2242_),
    .X(_2243_));
 sg13g2_mux2_1 _7616_ (.A0(\logix.ram_r[446] ),
    .A1(\logix.ram_r[445] ),
    .S(net282),
    .X(_1447_));
 sg13g2_mux2_1 _7617_ (.A0(\logix.ram_r[447] ),
    .A1(\logix.ram_r[446] ),
    .S(net282),
    .X(_1448_));
 sg13g2_mux2_1 _7618_ (.A0(\logix.ram_r[448] ),
    .A1(\logix.ram_r[447] ),
    .S(net282),
    .X(_1449_));
 sg13g2_mux2_1 _7619_ (.A0(\logix.ram_r[449] ),
    .A1(\logix.ram_r[448] ),
    .S(net282),
    .X(_1450_));
 sg13g2_mux2_1 _7620_ (.A0(\logix.ram_r[44] ),
    .A1(\logix.ram_r[43] ),
    .S(net282),
    .X(_1451_));
 sg13g2_mux2_1 _7621_ (.A0(\logix.ram_r[450] ),
    .A1(\logix.ram_r[449] ),
    .S(net282),
    .X(_1452_));
 sg13g2_mux2_1 _7622_ (.A0(\logix.ram_r[451] ),
    .A1(\logix.ram_r[450] ),
    .S(net282),
    .X(_1453_));
 sg13g2_mux2_1 _7623_ (.A0(\logix.ram_r[452] ),
    .A1(\logix.ram_r[451] ),
    .S(net282),
    .X(_1454_));
 sg13g2_mux2_1 _7624_ (.A0(\logix.ram_r[453] ),
    .A1(\logix.ram_r[452] ),
    .S(_2243_),
    .X(_1455_));
 sg13g2_mux2_1 _7625_ (.A0(\logix.ram_r[454] ),
    .A1(\logix.ram_r[453] ),
    .S(_2243_),
    .X(_1456_));
 sg13g2_buf_1 _7626_ (.A(_2242_),
    .X(_2244_));
 sg13g2_mux2_1 _7627_ (.A0(\logix.ram_r[455] ),
    .A1(\logix.ram_r[454] ),
    .S(net281),
    .X(_1457_));
 sg13g2_mux2_1 _7628_ (.A0(\logix.ram_r[456] ),
    .A1(\logix.ram_r[455] ),
    .S(net281),
    .X(_1458_));
 sg13g2_mux2_1 _7629_ (.A0(\logix.ram_r[457] ),
    .A1(\logix.ram_r[456] ),
    .S(net281),
    .X(_1459_));
 sg13g2_mux2_1 _7630_ (.A0(\logix.ram_r[458] ),
    .A1(\logix.ram_r[457] ),
    .S(_2244_),
    .X(_1460_));
 sg13g2_mux2_1 _7631_ (.A0(\logix.ram_r[459] ),
    .A1(\logix.ram_r[458] ),
    .S(_2244_),
    .X(_1461_));
 sg13g2_mux2_1 _7632_ (.A0(\logix.ram_r[45] ),
    .A1(\logix.ram_r[44] ),
    .S(net281),
    .X(_1462_));
 sg13g2_mux2_1 _7633_ (.A0(\logix.ram_r[460] ),
    .A1(\logix.ram_r[459] ),
    .S(net281),
    .X(_1463_));
 sg13g2_mux2_1 _7634_ (.A0(\logix.ram_r[461] ),
    .A1(\logix.ram_r[460] ),
    .S(net281),
    .X(_1464_));
 sg13g2_mux2_1 _7635_ (.A0(\logix.ram_r[462] ),
    .A1(\logix.ram_r[461] ),
    .S(net281),
    .X(_1465_));
 sg13g2_mux2_1 _7636_ (.A0(\logix.ram_r[463] ),
    .A1(\logix.ram_r[462] ),
    .S(net281),
    .X(_1466_));
 sg13g2_buf_1 _7637_ (.A(_2242_),
    .X(_2245_));
 sg13g2_mux2_1 _7638_ (.A0(\logix.ram_r[464] ),
    .A1(\logix.ram_r[463] ),
    .S(_2245_),
    .X(_1467_));
 sg13g2_mux2_1 _7639_ (.A0(\logix.ram_r[465] ),
    .A1(\logix.ram_r[464] ),
    .S(net280),
    .X(_1468_));
 sg13g2_mux2_1 _7640_ (.A0(\logix.ram_r[466] ),
    .A1(\logix.ram_r[465] ),
    .S(net280),
    .X(_1469_));
 sg13g2_mux2_1 _7641_ (.A0(\logix.ram_r[467] ),
    .A1(\logix.ram_r[466] ),
    .S(net280),
    .X(_1470_));
 sg13g2_mux2_1 _7642_ (.A0(\logix.ram_r[468] ),
    .A1(\logix.ram_r[467] ),
    .S(net280),
    .X(_1471_));
 sg13g2_mux2_1 _7643_ (.A0(\logix.ram_r[469] ),
    .A1(\logix.ram_r[468] ),
    .S(net280),
    .X(_1472_));
 sg13g2_mux2_1 _7644_ (.A0(\logix.ram_r[46] ),
    .A1(\logix.ram_r[45] ),
    .S(_2245_),
    .X(_1473_));
 sg13g2_mux2_1 _7645_ (.A0(\logix.ram_r[470] ),
    .A1(\logix.ram_r[469] ),
    .S(net280),
    .X(_1474_));
 sg13g2_mux2_1 _7646_ (.A0(\logix.ram_r[471] ),
    .A1(\logix.ram_r[470] ),
    .S(net280),
    .X(_1475_));
 sg13g2_mux2_1 _7647_ (.A0(\logix.ram_r[472] ),
    .A1(\logix.ram_r[471] ),
    .S(net280),
    .X(_1476_));
 sg13g2_buf_1 _7648_ (.A(_2242_),
    .X(_2246_));
 sg13g2_mux2_1 _7649_ (.A0(\logix.ram_r[473] ),
    .A1(\logix.ram_r[472] ),
    .S(net279),
    .X(_1477_));
 sg13g2_mux2_1 _7650_ (.A0(\logix.ram_r[474] ),
    .A1(\logix.ram_r[473] ),
    .S(net279),
    .X(_1478_));
 sg13g2_mux2_1 _7651_ (.A0(\logix.ram_r[475] ),
    .A1(\logix.ram_r[474] ),
    .S(net279),
    .X(_1479_));
 sg13g2_mux2_1 _7652_ (.A0(\logix.ram_r[476] ),
    .A1(\logix.ram_r[475] ),
    .S(net279),
    .X(_1480_));
 sg13g2_mux2_1 _7653_ (.A0(\logix.ram_r[477] ),
    .A1(\logix.ram_r[476] ),
    .S(net279),
    .X(_1481_));
 sg13g2_mux2_1 _7654_ (.A0(\logix.ram_r[478] ),
    .A1(\logix.ram_r[477] ),
    .S(_2246_),
    .X(_1482_));
 sg13g2_mux2_1 _7655_ (.A0(\logix.ram_r[479] ),
    .A1(\logix.ram_r[478] ),
    .S(net279),
    .X(_1483_));
 sg13g2_mux2_1 _7656_ (.A0(\logix.ram_r[47] ),
    .A1(\logix.ram_r[46] ),
    .S(_2246_),
    .X(_1484_));
 sg13g2_mux2_1 _7657_ (.A0(\logix.ram_r[480] ),
    .A1(\logix.ram_r[479] ),
    .S(net279),
    .X(_1485_));
 sg13g2_mux2_1 _7658_ (.A0(\logix.ram_r[481] ),
    .A1(\logix.ram_r[480] ),
    .S(net279),
    .X(_1486_));
 sg13g2_buf_1 _7659_ (.A(_2242_),
    .X(_2247_));
 sg13g2_mux2_1 _7660_ (.A0(\logix.ram_r[482] ),
    .A1(\logix.ram_r[481] ),
    .S(net278),
    .X(_1487_));
 sg13g2_mux2_1 _7661_ (.A0(\logix.ram_r[483] ),
    .A1(\logix.ram_r[482] ),
    .S(net278),
    .X(_1488_));
 sg13g2_mux2_1 _7662_ (.A0(\logix.ram_r[484] ),
    .A1(\logix.ram_r[483] ),
    .S(net278),
    .X(_1489_));
 sg13g2_mux2_1 _7663_ (.A0(\logix.ram_r[485] ),
    .A1(\logix.ram_r[484] ),
    .S(net278),
    .X(_1490_));
 sg13g2_mux2_1 _7664_ (.A0(\logix.ram_r[486] ),
    .A1(\logix.ram_r[485] ),
    .S(net278),
    .X(_1491_));
 sg13g2_mux2_1 _7665_ (.A0(\logix.ram_r[487] ),
    .A1(\logix.ram_r[486] ),
    .S(_2247_),
    .X(_1492_));
 sg13g2_mux2_1 _7666_ (.A0(\logix.ram_r[488] ),
    .A1(\logix.ram_r[487] ),
    .S(net278),
    .X(_1493_));
 sg13g2_mux2_1 _7667_ (.A0(\logix.ram_r[489] ),
    .A1(\logix.ram_r[488] ),
    .S(net278),
    .X(_1494_));
 sg13g2_mux2_1 _7668_ (.A0(\logix.ram_r[48] ),
    .A1(\logix.ram_r[47] ),
    .S(_2247_),
    .X(_1495_));
 sg13g2_mux2_1 _7669_ (.A0(\logix.ram_r[490] ),
    .A1(\logix.ram_r[489] ),
    .S(net278),
    .X(_1496_));
 sg13g2_buf_1 _7670_ (.A(_2242_),
    .X(_2248_));
 sg13g2_mux2_1 _7671_ (.A0(\logix.ram_r[491] ),
    .A1(\logix.ram_r[490] ),
    .S(net277),
    .X(_1497_));
 sg13g2_mux2_1 _7672_ (.A0(\logix.ram_r[492] ),
    .A1(\logix.ram_r[491] ),
    .S(net277),
    .X(_1498_));
 sg13g2_mux2_1 _7673_ (.A0(\logix.ram_r[493] ),
    .A1(\logix.ram_r[492] ),
    .S(net277),
    .X(_1499_));
 sg13g2_mux2_1 _7674_ (.A0(\logix.ram_r[494] ),
    .A1(\logix.ram_r[493] ),
    .S(net277),
    .X(_1500_));
 sg13g2_mux2_1 _7675_ (.A0(\logix.ram_r[495] ),
    .A1(\logix.ram_r[494] ),
    .S(net277),
    .X(_1501_));
 sg13g2_mux2_1 _7676_ (.A0(\logix.ram_r[496] ),
    .A1(\logix.ram_r[495] ),
    .S(net277),
    .X(_1502_));
 sg13g2_mux2_1 _7677_ (.A0(\logix.ram_r[497] ),
    .A1(\logix.ram_r[496] ),
    .S(net277),
    .X(_1503_));
 sg13g2_mux2_1 _7678_ (.A0(\logix.ram_r[498] ),
    .A1(\logix.ram_r[497] ),
    .S(_2248_),
    .X(_1504_));
 sg13g2_mux2_1 _7679_ (.A0(\logix.ram_r[499] ),
    .A1(\logix.ram_r[498] ),
    .S(net277),
    .X(_1505_));
 sg13g2_mux2_1 _7680_ (.A0(\logix.ram_r[49] ),
    .A1(\logix.ram_r[48] ),
    .S(_2248_),
    .X(_1506_));
 sg13g2_buf_1 _7681_ (.A(_2242_),
    .X(_2249_));
 sg13g2_mux2_1 _7682_ (.A0(\logix.ram_r[4] ),
    .A1(\logix.ram_r[3] ),
    .S(_2249_),
    .X(_1507_));
 sg13g2_mux2_1 _7683_ (.A0(\logix.ram_r[500] ),
    .A1(\logix.ram_r[499] ),
    .S(net276),
    .X(_1508_));
 sg13g2_mux2_1 _7684_ (.A0(\logix.ram_r[501] ),
    .A1(\logix.ram_r[500] ),
    .S(_2249_),
    .X(_1509_));
 sg13g2_mux2_1 _7685_ (.A0(\logix.ram_r[502] ),
    .A1(\logix.ram_r[501] ),
    .S(net276),
    .X(_1510_));
 sg13g2_mux2_1 _7686_ (.A0(\logix.ram_r[503] ),
    .A1(\logix.ram_r[502] ),
    .S(net276),
    .X(_1511_));
 sg13g2_mux2_1 _7687_ (.A0(\logix.ram_r[504] ),
    .A1(\logix.ram_r[503] ),
    .S(net276),
    .X(_1512_));
 sg13g2_mux2_1 _7688_ (.A0(\logix.ram_r[505] ),
    .A1(\logix.ram_r[504] ),
    .S(net276),
    .X(_1513_));
 sg13g2_mux2_1 _7689_ (.A0(\logix.ram_r[506] ),
    .A1(\logix.ram_r[505] ),
    .S(net276),
    .X(_1514_));
 sg13g2_mux2_1 _7690_ (.A0(\logix.ram_r[507] ),
    .A1(\logix.ram_r[506] ),
    .S(net276),
    .X(_1515_));
 sg13g2_mux2_1 _7691_ (.A0(\logix.ram_r[508] ),
    .A1(\logix.ram_r[507] ),
    .S(net276),
    .X(_1516_));
 sg13g2_buf_1 _7692_ (.A(_2201_),
    .X(_2250_));
 sg13g2_buf_1 _7693_ (.A(_2250_),
    .X(_2251_));
 sg13g2_mux2_1 _7694_ (.A0(\logix.ram_r[509] ),
    .A1(\logix.ram_r[508] ),
    .S(net275),
    .X(_1517_));
 sg13g2_mux2_1 _7695_ (.A0(\logix.ram_r[50] ),
    .A1(\logix.ram_r[49] ),
    .S(_2251_),
    .X(_1518_));
 sg13g2_mux2_1 _7696_ (.A0(\logix.ram_r[510] ),
    .A1(\logix.ram_r[509] ),
    .S(net275),
    .X(_1519_));
 sg13g2_mux2_1 _7697_ (.A0(\logix.ram_r[511] ),
    .A1(\logix.ram_r[510] ),
    .S(net275),
    .X(_1520_));
 sg13g2_mux2_1 _7698_ (.A0(\logix.ram_r[512] ),
    .A1(\logix.ram_r[511] ),
    .S(net275),
    .X(_1521_));
 sg13g2_mux2_1 _7699_ (.A0(\logix.ram_r[513] ),
    .A1(\logix.ram_r[512] ),
    .S(net275),
    .X(_1522_));
 sg13g2_mux2_1 _7700_ (.A0(\logix.ram_r[514] ),
    .A1(\logix.ram_r[513] ),
    .S(net275),
    .X(_1523_));
 sg13g2_mux2_1 _7701_ (.A0(\logix.ram_r[515] ),
    .A1(\logix.ram_r[514] ),
    .S(net275),
    .X(_1524_));
 sg13g2_mux2_1 _7702_ (.A0(\logix.ram_r[516] ),
    .A1(\logix.ram_r[515] ),
    .S(_2251_),
    .X(_1525_));
 sg13g2_mux2_1 _7703_ (.A0(\logix.ram_r[517] ),
    .A1(\logix.ram_r[516] ),
    .S(net275),
    .X(_1526_));
 sg13g2_buf_1 _7704_ (.A(_2250_),
    .X(_2252_));
 sg13g2_mux2_1 _7705_ (.A0(\logix.ram_r[518] ),
    .A1(\logix.ram_r[517] ),
    .S(net274),
    .X(_1527_));
 sg13g2_mux2_1 _7706_ (.A0(\logix.ram_r[519] ),
    .A1(\logix.ram_r[518] ),
    .S(net274),
    .X(_1528_));
 sg13g2_mux2_1 _7707_ (.A0(\logix.ram_r[51] ),
    .A1(\logix.ram_r[50] ),
    .S(_2252_),
    .X(_1529_));
 sg13g2_mux2_1 _7708_ (.A0(\logix.ram_r[520] ),
    .A1(\logix.ram_r[519] ),
    .S(net274),
    .X(_1530_));
 sg13g2_mux2_1 _7709_ (.A0(\logix.ram_r[521] ),
    .A1(\logix.ram_r[520] ),
    .S(net274),
    .X(_1531_));
 sg13g2_mux2_1 _7710_ (.A0(\logix.ram_r[522] ),
    .A1(\logix.ram_r[521] ),
    .S(_2252_),
    .X(_1532_));
 sg13g2_mux2_1 _7711_ (.A0(\logix.ram_r[523] ),
    .A1(\logix.ram_r[522] ),
    .S(net274),
    .X(_1533_));
 sg13g2_mux2_1 _7712_ (.A0(\logix.ram_r[524] ),
    .A1(\logix.ram_r[523] ),
    .S(net274),
    .X(_1534_));
 sg13g2_mux2_1 _7713_ (.A0(\logix.ram_r[525] ),
    .A1(\logix.ram_r[524] ),
    .S(net274),
    .X(_1535_));
 sg13g2_mux2_1 _7714_ (.A0(\logix.ram_r[526] ),
    .A1(\logix.ram_r[525] ),
    .S(net274),
    .X(_1536_));
 sg13g2_buf_1 _7715_ (.A(_2250_),
    .X(_2253_));
 sg13g2_mux2_1 _7716_ (.A0(\logix.ram_r[527] ),
    .A1(\logix.ram_r[526] ),
    .S(net273),
    .X(_1537_));
 sg13g2_mux2_1 _7717_ (.A0(\logix.ram_r[528] ),
    .A1(\logix.ram_r[527] ),
    .S(net273),
    .X(_1538_));
 sg13g2_mux2_1 _7718_ (.A0(\logix.ram_r[529] ),
    .A1(\logix.ram_r[528] ),
    .S(net273),
    .X(_1539_));
 sg13g2_mux2_1 _7719_ (.A0(\logix.ram_r[52] ),
    .A1(\logix.ram_r[51] ),
    .S(_2253_),
    .X(_1540_));
 sg13g2_mux2_1 _7720_ (.A0(\logix.ram_r[530] ),
    .A1(\logix.ram_r[529] ),
    .S(net273),
    .X(_1541_));
 sg13g2_mux2_1 _7721_ (.A0(\logix.ram_r[531] ),
    .A1(\logix.ram_r[530] ),
    .S(net273),
    .X(_1542_));
 sg13g2_mux2_1 _7722_ (.A0(\logix.ram_r[532] ),
    .A1(\logix.ram_r[531] ),
    .S(net273),
    .X(_1543_));
 sg13g2_mux2_1 _7723_ (.A0(\logix.ram_r[533] ),
    .A1(\logix.ram_r[532] ),
    .S(net273),
    .X(_1544_));
 sg13g2_mux2_1 _7724_ (.A0(\logix.ram_r[534] ),
    .A1(\logix.ram_r[533] ),
    .S(net273),
    .X(_1545_));
 sg13g2_mux2_1 _7725_ (.A0(\logix.ram_r[535] ),
    .A1(\logix.ram_r[534] ),
    .S(_2253_),
    .X(_1546_));
 sg13g2_buf_1 _7726_ (.A(_2250_),
    .X(_2254_));
 sg13g2_mux2_1 _7727_ (.A0(\logix.ram_r[536] ),
    .A1(\logix.ram_r[535] ),
    .S(net272),
    .X(_1547_));
 sg13g2_mux2_1 _7728_ (.A0(\logix.ram_r[537] ),
    .A1(\logix.ram_r[536] ),
    .S(net272),
    .X(_1548_));
 sg13g2_mux2_1 _7729_ (.A0(\logix.ram_r[538] ),
    .A1(\logix.ram_r[537] ),
    .S(net272),
    .X(_1549_));
 sg13g2_mux2_1 _7730_ (.A0(\logix.ram_r[539] ),
    .A1(\logix.ram_r[538] ),
    .S(net272),
    .X(_1550_));
 sg13g2_mux2_1 _7731_ (.A0(\logix.ram_r[53] ),
    .A1(\logix.ram_r[52] ),
    .S(_2254_),
    .X(_1551_));
 sg13g2_mux2_1 _7732_ (.A0(\logix.ram_r[540] ),
    .A1(\logix.ram_r[539] ),
    .S(_2254_),
    .X(_1552_));
 sg13g2_mux2_1 _7733_ (.A0(\logix.ram_r[541] ),
    .A1(\logix.ram_r[540] ),
    .S(net272),
    .X(_1553_));
 sg13g2_mux2_1 _7734_ (.A0(\logix.ram_r[542] ),
    .A1(\logix.ram_r[541] ),
    .S(net272),
    .X(_1554_));
 sg13g2_mux2_1 _7735_ (.A0(\logix.ram_r[543] ),
    .A1(\logix.ram_r[542] ),
    .S(net272),
    .X(_1555_));
 sg13g2_mux2_1 _7736_ (.A0(\logix.ram_r[544] ),
    .A1(\logix.ram_r[543] ),
    .S(net272),
    .X(_1556_));
 sg13g2_buf_1 _7737_ (.A(_2250_),
    .X(_2255_));
 sg13g2_mux2_1 _7738_ (.A0(\logix.ram_r[545] ),
    .A1(\logix.ram_r[544] ),
    .S(net271),
    .X(_1557_));
 sg13g2_mux2_1 _7739_ (.A0(\logix.ram_r[546] ),
    .A1(\logix.ram_r[545] ),
    .S(net271),
    .X(_1558_));
 sg13g2_mux2_1 _7740_ (.A0(\logix.ram_r[547] ),
    .A1(\logix.ram_r[546] ),
    .S(net271),
    .X(_1559_));
 sg13g2_mux2_1 _7741_ (.A0(\logix.ram_r[548] ),
    .A1(\logix.ram_r[547] ),
    .S(net271),
    .X(_1560_));
 sg13g2_mux2_1 _7742_ (.A0(\logix.ram_r[549] ),
    .A1(\logix.ram_r[548] ),
    .S(net271),
    .X(_1561_));
 sg13g2_mux2_1 _7743_ (.A0(\logix.ram_r[54] ),
    .A1(\logix.ram_r[53] ),
    .S(net271),
    .X(_1562_));
 sg13g2_mux2_1 _7744_ (.A0(\logix.ram_r[550] ),
    .A1(\logix.ram_r[549] ),
    .S(net271),
    .X(_1563_));
 sg13g2_mux2_1 _7745_ (.A0(\logix.ram_r[551] ),
    .A1(\logix.ram_r[550] ),
    .S(net271),
    .X(_1564_));
 sg13g2_mux2_1 _7746_ (.A0(\logix.ram_r[552] ),
    .A1(\logix.ram_r[551] ),
    .S(_2255_),
    .X(_1565_));
 sg13g2_mux2_1 _7747_ (.A0(\logix.ram_r[553] ),
    .A1(\logix.ram_r[552] ),
    .S(_2255_),
    .X(_1566_));
 sg13g2_buf_1 _7748_ (.A(_2250_),
    .X(_2256_));
 sg13g2_mux2_1 _7749_ (.A0(\logix.ram_r[554] ),
    .A1(\logix.ram_r[553] ),
    .S(net270),
    .X(_1567_));
 sg13g2_mux2_1 _7750_ (.A0(\logix.ram_r[555] ),
    .A1(\logix.ram_r[554] ),
    .S(net270),
    .X(_1568_));
 sg13g2_mux2_1 _7751_ (.A0(\logix.ram_r[556] ),
    .A1(\logix.ram_r[555] ),
    .S(net270),
    .X(_1569_));
 sg13g2_mux2_1 _7752_ (.A0(\logix.ram_r[557] ),
    .A1(\logix.ram_r[556] ),
    .S(net270),
    .X(_1570_));
 sg13g2_mux2_1 _7753_ (.A0(\logix.ram_r[558] ),
    .A1(\logix.ram_r[557] ),
    .S(net270),
    .X(_1571_));
 sg13g2_mux2_1 _7754_ (.A0(\logix.ram_r[559] ),
    .A1(\logix.ram_r[558] ),
    .S(net270),
    .X(_1572_));
 sg13g2_mux2_1 _7755_ (.A0(\logix.ram_r[55] ),
    .A1(\logix.ram_r[54] ),
    .S(_2256_),
    .X(_1573_));
 sg13g2_mux2_1 _7756_ (.A0(\logix.ram_r[560] ),
    .A1(\logix.ram_r[559] ),
    .S(net270),
    .X(_1574_));
 sg13g2_mux2_1 _7757_ (.A0(\logix.ram_r[561] ),
    .A1(\logix.ram_r[560] ),
    .S(net270),
    .X(_1575_));
 sg13g2_mux2_1 _7758_ (.A0(\logix.ram_r[562] ),
    .A1(\logix.ram_r[561] ),
    .S(_2256_),
    .X(_1576_));
 sg13g2_buf_1 _7759_ (.A(_2250_),
    .X(_2257_));
 sg13g2_mux2_1 _7760_ (.A0(\logix.ram_r[563] ),
    .A1(\logix.ram_r[562] ),
    .S(net269),
    .X(_1577_));
 sg13g2_mux2_1 _7761_ (.A0(\logix.ram_r[564] ),
    .A1(\logix.ram_r[563] ),
    .S(net269),
    .X(_1578_));
 sg13g2_mux2_1 _7762_ (.A0(\logix.ram_r[565] ),
    .A1(\logix.ram_r[564] ),
    .S(_2257_),
    .X(_1579_));
 sg13g2_mux2_1 _7763_ (.A0(\logix.ram_r[566] ),
    .A1(\logix.ram_r[565] ),
    .S(net269),
    .X(_1580_));
 sg13g2_mux2_1 _7764_ (.A0(\logix.ram_r[567] ),
    .A1(\logix.ram_r[566] ),
    .S(net269),
    .X(_1581_));
 sg13g2_mux2_1 _7765_ (.A0(\logix.ram_r[568] ),
    .A1(\logix.ram_r[567] ),
    .S(net269),
    .X(_1582_));
 sg13g2_mux2_1 _7766_ (.A0(\logix.ram_r[569] ),
    .A1(\logix.ram_r[568] ),
    .S(net269),
    .X(_1583_));
 sg13g2_mux2_1 _7767_ (.A0(\logix.ram_r[56] ),
    .A1(\logix.ram_r[55] ),
    .S(net269),
    .X(_1584_));
 sg13g2_mux2_1 _7768_ (.A0(\logix.ram_r[570] ),
    .A1(\logix.ram_r[569] ),
    .S(net269),
    .X(_1585_));
 sg13g2_mux2_1 _7769_ (.A0(\logix.ram_r[571] ),
    .A1(\logix.ram_r[570] ),
    .S(_2257_),
    .X(_1586_));
 sg13g2_buf_1 _7770_ (.A(_2201_),
    .X(_2258_));
 sg13g2_buf_1 _7771_ (.A(_2258_),
    .X(_2259_));
 sg13g2_mux2_1 _7772_ (.A0(\logix.ram_r[572] ),
    .A1(\logix.ram_r[571] ),
    .S(net268),
    .X(_1587_));
 sg13g2_mux2_1 _7773_ (.A0(\logix.ram_r[573] ),
    .A1(\logix.ram_r[572] ),
    .S(net268),
    .X(_1588_));
 sg13g2_mux2_1 _7774_ (.A0(\logix.ram_r[574] ),
    .A1(\logix.ram_r[573] ),
    .S(net268),
    .X(_1589_));
 sg13g2_mux2_1 _7775_ (.A0(\logix.ram_r[575] ),
    .A1(\logix.ram_r[574] ),
    .S(net268),
    .X(_1590_));
 sg13g2_mux2_1 _7776_ (.A0(\logix.ram_r[576] ),
    .A1(\logix.ram_r[575] ),
    .S(net268),
    .X(_1591_));
 sg13g2_mux2_1 _7777_ (.A0(\logix.ram_r[577] ),
    .A1(\logix.ram_r[576] ),
    .S(net268),
    .X(_1592_));
 sg13g2_mux2_1 _7778_ (.A0(\logix.ram_r[578] ),
    .A1(\logix.ram_r[577] ),
    .S(_2259_),
    .X(_1593_));
 sg13g2_mux2_1 _7779_ (.A0(\logix.ram_r[579] ),
    .A1(\logix.ram_r[578] ),
    .S(net268),
    .X(_1594_));
 sg13g2_mux2_1 _7780_ (.A0(\logix.ram_r[57] ),
    .A1(\logix.ram_r[56] ),
    .S(_2259_),
    .X(_1595_));
 sg13g2_mux2_1 _7781_ (.A0(\logix.ram_r[580] ),
    .A1(\logix.ram_r[579] ),
    .S(net268),
    .X(_1596_));
 sg13g2_buf_1 _7782_ (.A(_2258_),
    .X(_2260_));
 sg13g2_mux2_1 _7783_ (.A0(\logix.ram_r[581] ),
    .A1(\logix.ram_r[580] ),
    .S(net267),
    .X(_1597_));
 sg13g2_mux2_1 _7784_ (.A0(\logix.ram_r[582] ),
    .A1(\logix.ram_r[581] ),
    .S(net267),
    .X(_1598_));
 sg13g2_mux2_1 _7785_ (.A0(\logix.ram_r[583] ),
    .A1(\logix.ram_r[582] ),
    .S(net267),
    .X(_1599_));
 sg13g2_mux2_1 _7786_ (.A0(\logix.ram_r[584] ),
    .A1(\logix.ram_r[583] ),
    .S(net267),
    .X(_1600_));
 sg13g2_mux2_1 _7787_ (.A0(\logix.ram_r[585] ),
    .A1(\logix.ram_r[584] ),
    .S(_2260_),
    .X(_1601_));
 sg13g2_mux2_1 _7788_ (.A0(\logix.ram_r[586] ),
    .A1(\logix.ram_r[585] ),
    .S(_2260_),
    .X(_1602_));
 sg13g2_mux2_1 _7789_ (.A0(\logix.ram_r[587] ),
    .A1(\logix.ram_r[586] ),
    .S(net267),
    .X(_1603_));
 sg13g2_mux2_1 _7790_ (.A0(\logix.ram_r[588] ),
    .A1(\logix.ram_r[587] ),
    .S(net267),
    .X(_1604_));
 sg13g2_mux2_1 _7791_ (.A0(\logix.ram_r[589] ),
    .A1(\logix.ram_r[588] ),
    .S(net267),
    .X(_1605_));
 sg13g2_mux2_1 _7792_ (.A0(\logix.ram_r[58] ),
    .A1(\logix.ram_r[57] ),
    .S(net267),
    .X(_1606_));
 sg13g2_buf_1 _7793_ (.A(_2258_),
    .X(_2261_));
 sg13g2_mux2_1 _7794_ (.A0(\logix.ram_r[590] ),
    .A1(\logix.ram_r[589] ),
    .S(net266),
    .X(_1607_));
 sg13g2_mux2_1 _7795_ (.A0(\logix.ram_r[591] ),
    .A1(\logix.ram_r[590] ),
    .S(net266),
    .X(_1608_));
 sg13g2_mux2_1 _7796_ (.A0(\logix.ram_r[592] ),
    .A1(\logix.ram_r[591] ),
    .S(net266),
    .X(_1609_));
 sg13g2_mux2_1 _7797_ (.A0(\logix.ram_r[593] ),
    .A1(\logix.ram_r[592] ),
    .S(net266),
    .X(_1610_));
 sg13g2_mux2_1 _7798_ (.A0(\logix.ram_r[594] ),
    .A1(\logix.ram_r[593] ),
    .S(_2261_),
    .X(_1611_));
 sg13g2_mux2_1 _7799_ (.A0(\logix.ram_r[595] ),
    .A1(\logix.ram_r[594] ),
    .S(net266),
    .X(_1612_));
 sg13g2_mux2_1 _7800_ (.A0(\logix.ram_r[596] ),
    .A1(\logix.ram_r[595] ),
    .S(net266),
    .X(_1613_));
 sg13g2_mux2_1 _7801_ (.A0(\logix.ram_r[597] ),
    .A1(\logix.ram_r[596] ),
    .S(net266),
    .X(_1614_));
 sg13g2_mux2_1 _7802_ (.A0(\logix.ram_r[598] ),
    .A1(\logix.ram_r[597] ),
    .S(net266),
    .X(_1615_));
 sg13g2_mux2_1 _7803_ (.A0(\logix.ram_r[599] ),
    .A1(\logix.ram_r[598] ),
    .S(_2261_),
    .X(_1616_));
 sg13g2_buf_1 _7804_ (.A(_2258_),
    .X(_2262_));
 sg13g2_mux2_1 _7805_ (.A0(\logix.ram_r[59] ),
    .A1(\logix.ram_r[58] ),
    .S(net265),
    .X(_1617_));
 sg13g2_mux2_1 _7806_ (.A0(\logix.ram_r[5] ),
    .A1(\logix.ram_r[4] ),
    .S(net265),
    .X(_1618_));
 sg13g2_mux2_1 _7807_ (.A0(\logix.ram_r[600] ),
    .A1(\logix.ram_r[599] ),
    .S(net265),
    .X(_1619_));
 sg13g2_mux2_1 _7808_ (.A0(\logix.ram_r[601] ),
    .A1(\logix.ram_r[600] ),
    .S(net265),
    .X(_1620_));
 sg13g2_mux2_1 _7809_ (.A0(\logix.ram_r[602] ),
    .A1(\logix.ram_r[601] ),
    .S(net265),
    .X(_1621_));
 sg13g2_mux2_1 _7810_ (.A0(\logix.ram_r[603] ),
    .A1(\logix.ram_r[602] ),
    .S(net265),
    .X(_1622_));
 sg13g2_mux2_1 _7811_ (.A0(\logix.ram_r[604] ),
    .A1(\logix.ram_r[603] ),
    .S(net265),
    .X(_1623_));
 sg13g2_mux2_1 _7812_ (.A0(\logix.ram_r[605] ),
    .A1(\logix.ram_r[604] ),
    .S(net265),
    .X(_1624_));
 sg13g2_mux2_1 _7813_ (.A0(\logix.ram_r[606] ),
    .A1(\logix.ram_r[605] ),
    .S(_2262_),
    .X(_1625_));
 sg13g2_mux2_1 _7814_ (.A0(\logix.ram_r[607] ),
    .A1(\logix.ram_r[606] ),
    .S(_2262_),
    .X(_1626_));
 sg13g2_buf_1 _7815_ (.A(_2258_),
    .X(_2263_));
 sg13g2_mux2_1 _7816_ (.A0(\logix.ram_r[608] ),
    .A1(\logix.ram_r[607] ),
    .S(net264),
    .X(_1627_));
 sg13g2_mux2_1 _7817_ (.A0(\logix.ram_r[609] ),
    .A1(\logix.ram_r[608] ),
    .S(net264),
    .X(_1628_));
 sg13g2_mux2_1 _7818_ (.A0(\logix.ram_r[60] ),
    .A1(\logix.ram_r[59] ),
    .S(_2263_),
    .X(_1629_));
 sg13g2_mux2_1 _7819_ (.A0(\logix.ram_r[610] ),
    .A1(\logix.ram_r[609] ),
    .S(_2263_),
    .X(_1630_));
 sg13g2_mux2_1 _7820_ (.A0(\logix.ram_r[611] ),
    .A1(\logix.ram_r[610] ),
    .S(net264),
    .X(_1631_));
 sg13g2_mux2_1 _7821_ (.A0(\logix.ram_r[612] ),
    .A1(\logix.ram_r[611] ),
    .S(net264),
    .X(_1632_));
 sg13g2_mux2_1 _7822_ (.A0(\logix.ram_r[613] ),
    .A1(\logix.ram_r[612] ),
    .S(net264),
    .X(_1633_));
 sg13g2_mux2_1 _7823_ (.A0(\logix.ram_r[614] ),
    .A1(\logix.ram_r[613] ),
    .S(net264),
    .X(_1634_));
 sg13g2_mux2_1 _7824_ (.A0(\logix.ram_r[615] ),
    .A1(\logix.ram_r[614] ),
    .S(net264),
    .X(_1635_));
 sg13g2_mux2_1 _7825_ (.A0(\logix.ram_r[616] ),
    .A1(\logix.ram_r[615] ),
    .S(net264),
    .X(_1636_));
 sg13g2_buf_1 _7826_ (.A(_2258_),
    .X(_2264_));
 sg13g2_mux2_1 _7827_ (.A0(\logix.ram_r[617] ),
    .A1(\logix.ram_r[616] ),
    .S(net263),
    .X(_1637_));
 sg13g2_mux2_1 _7828_ (.A0(\logix.ram_r[618] ),
    .A1(\logix.ram_r[617] ),
    .S(net263),
    .X(_1638_));
 sg13g2_mux2_1 _7829_ (.A0(\logix.ram_r[619] ),
    .A1(\logix.ram_r[618] ),
    .S(net263),
    .X(_1639_));
 sg13g2_mux2_1 _7830_ (.A0(\logix.ram_r[61] ),
    .A1(\logix.ram_r[60] ),
    .S(_2264_),
    .X(_1640_));
 sg13g2_mux2_1 _7831_ (.A0(\logix.ram_r[620] ),
    .A1(\logix.ram_r[619] ),
    .S(net263),
    .X(_1641_));
 sg13g2_mux2_1 _7832_ (.A0(\logix.ram_r[621] ),
    .A1(\logix.ram_r[620] ),
    .S(net263),
    .X(_1642_));
 sg13g2_mux2_1 _7833_ (.A0(\logix.ram_r[622] ),
    .A1(\logix.ram_r[621] ),
    .S(net263),
    .X(_1643_));
 sg13g2_mux2_1 _7834_ (.A0(\logix.ram_r[623] ),
    .A1(\logix.ram_r[622] ),
    .S(net263),
    .X(_1644_));
 sg13g2_mux2_1 _7835_ (.A0(\logix.ram_r[624] ),
    .A1(\logix.ram_r[623] ),
    .S(net263),
    .X(_1645_));
 sg13g2_mux2_1 _7836_ (.A0(\logix.ram_r[625] ),
    .A1(\logix.ram_r[624] ),
    .S(_2264_),
    .X(_1646_));
 sg13g2_buf_1 _7837_ (.A(_2258_),
    .X(_2265_));
 sg13g2_mux2_1 _7838_ (.A0(\logix.ram_r[626] ),
    .A1(\logix.ram_r[625] ),
    .S(net262),
    .X(_1647_));
 sg13g2_mux2_1 _7839_ (.A0(\logix.ram_r[627] ),
    .A1(\logix.ram_r[626] ),
    .S(net262),
    .X(_1648_));
 sg13g2_mux2_1 _7840_ (.A0(\logix.ram_r[628] ),
    .A1(\logix.ram_r[627] ),
    .S(net262),
    .X(_1649_));
 sg13g2_mux2_1 _7841_ (.A0(\logix.ram_r[629] ),
    .A1(\logix.ram_r[628] ),
    .S(net262),
    .X(_1650_));
 sg13g2_mux2_1 _7842_ (.A0(\logix.ram_r[62] ),
    .A1(\logix.ram_r[61] ),
    .S(_2265_),
    .X(_1651_));
 sg13g2_mux2_1 _7843_ (.A0(\logix.ram_r[630] ),
    .A1(\logix.ram_r[629] ),
    .S(net262),
    .X(_1652_));
 sg13g2_mux2_1 _7844_ (.A0(\logix.ram_r[631] ),
    .A1(\logix.ram_r[630] ),
    .S(net262),
    .X(_1653_));
 sg13g2_mux2_1 _7845_ (.A0(\logix.ram_r[632] ),
    .A1(\logix.ram_r[631] ),
    .S(_2265_),
    .X(_1654_));
 sg13g2_mux2_1 _7846_ (.A0(\logix.ram_r[633] ),
    .A1(\logix.ram_r[632] ),
    .S(net262),
    .X(_1655_));
 sg13g2_mux2_1 _7847_ (.A0(\logix.ram_r[634] ),
    .A1(\logix.ram_r[633] ),
    .S(net262),
    .X(_1656_));
 sg13g2_buf_1 _7848_ (.A(_2064_),
    .X(_2266_));
 sg13g2_buf_1 _7849_ (.A(_2266_),
    .X(_2267_));
 sg13g2_mux2_1 _7850_ (.A0(\logix.ram_r[635] ),
    .A1(\logix.ram_r[634] ),
    .S(net261),
    .X(_1657_));
 sg13g2_mux2_1 _7851_ (.A0(\logix.ram_r[636] ),
    .A1(\logix.ram_r[635] ),
    .S(net261),
    .X(_1658_));
 sg13g2_mux2_1 _7852_ (.A0(\logix.ram_r[637] ),
    .A1(\logix.ram_r[636] ),
    .S(_2267_),
    .X(_1659_));
 sg13g2_mux2_1 _7853_ (.A0(\logix.ram_r[638] ),
    .A1(\logix.ram_r[637] ),
    .S(net261),
    .X(_1660_));
 sg13g2_mux2_1 _7854_ (.A0(\logix.ram_r[639] ),
    .A1(\logix.ram_r[638] ),
    .S(_2267_),
    .X(_1661_));
 sg13g2_mux2_1 _7855_ (.A0(\logix.ram_r[63] ),
    .A1(\logix.ram_r[62] ),
    .S(net261),
    .X(_1662_));
 sg13g2_mux2_1 _7856_ (.A0(\logix.ram_r[640] ),
    .A1(\logix.ram_r[639] ),
    .S(net261),
    .X(_1663_));
 sg13g2_mux2_1 _7857_ (.A0(\logix.ram_r[641] ),
    .A1(\logix.ram_r[640] ),
    .S(net261),
    .X(_1664_));
 sg13g2_mux2_1 _7858_ (.A0(\logix.ram_r[642] ),
    .A1(\logix.ram_r[641] ),
    .S(net261),
    .X(_1665_));
 sg13g2_mux2_1 _7859_ (.A0(\logix.ram_r[643] ),
    .A1(\logix.ram_r[642] ),
    .S(net261),
    .X(_1666_));
 sg13g2_buf_1 _7860_ (.A(_2266_),
    .X(_2268_));
 sg13g2_mux2_1 _7861_ (.A0(\logix.ram_r[644] ),
    .A1(\logix.ram_r[643] ),
    .S(_2268_),
    .X(_1667_));
 sg13g2_mux2_1 _7862_ (.A0(\logix.ram_r[645] ),
    .A1(\logix.ram_r[644] ),
    .S(net260),
    .X(_1668_));
 sg13g2_mux2_1 _7863_ (.A0(\logix.ram_r[646] ),
    .A1(\logix.ram_r[645] ),
    .S(net260),
    .X(_1669_));
 sg13g2_mux2_1 _7864_ (.A0(\logix.ram_r[647] ),
    .A1(\logix.ram_r[646] ),
    .S(net260),
    .X(_1670_));
 sg13g2_mux2_1 _7865_ (.A0(\logix.ram_r[648] ),
    .A1(\logix.ram_r[647] ),
    .S(net260),
    .X(_1671_));
 sg13g2_mux2_1 _7866_ (.A0(\logix.ram_r[649] ),
    .A1(\logix.ram_r[648] ),
    .S(net260),
    .X(_1672_));
 sg13g2_mux2_1 _7867_ (.A0(\logix.ram_r[64] ),
    .A1(\logix.ram_r[63] ),
    .S(_2268_),
    .X(_1673_));
 sg13g2_mux2_1 _7868_ (.A0(\logix.ram_r[650] ),
    .A1(\logix.ram_r[649] ),
    .S(net260),
    .X(_1674_));
 sg13g2_mux2_1 _7869_ (.A0(\logix.ram_r[651] ),
    .A1(\logix.ram_r[650] ),
    .S(net260),
    .X(_1675_));
 sg13g2_mux2_1 _7870_ (.A0(\logix.ram_r[652] ),
    .A1(\logix.ram_r[651] ),
    .S(net260),
    .X(_1676_));
 sg13g2_buf_1 _7871_ (.A(_2266_),
    .X(_2269_));
 sg13g2_mux2_1 _7872_ (.A0(\logix.ram_r[653] ),
    .A1(\logix.ram_r[652] ),
    .S(net259),
    .X(_1677_));
 sg13g2_mux2_1 _7873_ (.A0(\logix.ram_r[654] ),
    .A1(\logix.ram_r[653] ),
    .S(net259),
    .X(_1678_));
 sg13g2_mux2_1 _7874_ (.A0(\logix.ram_r[655] ),
    .A1(\logix.ram_r[654] ),
    .S(net259),
    .X(_1679_));
 sg13g2_mux2_1 _7875_ (.A0(\logix.ram_r[656] ),
    .A1(\logix.ram_r[655] ),
    .S(_2269_),
    .X(_1680_));
 sg13g2_mux2_1 _7876_ (.A0(\logix.ram_r[657] ),
    .A1(\logix.ram_r[656] ),
    .S(net259),
    .X(_1681_));
 sg13g2_mux2_1 _7877_ (.A0(\logix.ram_r[658] ),
    .A1(\logix.ram_r[657] ),
    .S(net259),
    .X(_1682_));
 sg13g2_mux2_1 _7878_ (.A0(\logix.ram_r[659] ),
    .A1(\logix.ram_r[658] ),
    .S(net259),
    .X(_1683_));
 sg13g2_mux2_1 _7879_ (.A0(\logix.ram_r[65] ),
    .A1(\logix.ram_r[64] ),
    .S(_2269_),
    .X(_1684_));
 sg13g2_mux2_1 _7880_ (.A0(\logix.ram_r[660] ),
    .A1(\logix.ram_r[659] ),
    .S(net259),
    .X(_1685_));
 sg13g2_mux2_1 _7881_ (.A0(\logix.ram_r[661] ),
    .A1(\logix.ram_r[660] ),
    .S(net259),
    .X(_1686_));
 sg13g2_buf_1 _7882_ (.A(_2266_),
    .X(_2270_));
 sg13g2_mux2_1 _7883_ (.A0(\logix.ram_r[662] ),
    .A1(\logix.ram_r[661] ),
    .S(net258),
    .X(_1687_));
 sg13g2_mux2_1 _7884_ (.A0(\logix.ram_r[663] ),
    .A1(\logix.ram_r[662] ),
    .S(net258),
    .X(_1688_));
 sg13g2_mux2_1 _7885_ (.A0(\logix.ram_r[664] ),
    .A1(\logix.ram_r[663] ),
    .S(_2270_),
    .X(_1689_));
 sg13g2_mux2_1 _7886_ (.A0(\logix.ram_r[665] ),
    .A1(\logix.ram_r[664] ),
    .S(net258),
    .X(_1690_));
 sg13g2_mux2_1 _7887_ (.A0(\logix.ram_r[666] ),
    .A1(\logix.ram_r[665] ),
    .S(net258),
    .X(_1691_));
 sg13g2_mux2_1 _7888_ (.A0(\logix.ram_r[667] ),
    .A1(\logix.ram_r[666] ),
    .S(net258),
    .X(_1692_));
 sg13g2_mux2_1 _7889_ (.A0(\logix.ram_r[668] ),
    .A1(\logix.ram_r[667] ),
    .S(_2270_),
    .X(_1693_));
 sg13g2_mux2_1 _7890_ (.A0(\logix.ram_r[669] ),
    .A1(\logix.ram_r[668] ),
    .S(net258),
    .X(_1694_));
 sg13g2_mux2_1 _7891_ (.A0(\logix.ram_r[66] ),
    .A1(\logix.ram_r[65] ),
    .S(net258),
    .X(_1695_));
 sg13g2_mux2_1 _7892_ (.A0(\logix.ram_r[670] ),
    .A1(\logix.ram_r[669] ),
    .S(net258),
    .X(_1696_));
 sg13g2_buf_1 _7893_ (.A(_2266_),
    .X(_2271_));
 sg13g2_mux2_1 _7894_ (.A0(\logix.ram_r[671] ),
    .A1(\logix.ram_r[670] ),
    .S(net257),
    .X(_1697_));
 sg13g2_mux2_1 _7895_ (.A0(\logix.ram_r[672] ),
    .A1(\logix.ram_r[671] ),
    .S(net257),
    .X(_1698_));
 sg13g2_mux2_1 _7896_ (.A0(\logix.ram_r[673] ),
    .A1(\logix.ram_r[672] ),
    .S(_2271_),
    .X(_1699_));
 sg13g2_mux2_1 _7897_ (.A0(\logix.ram_r[674] ),
    .A1(\logix.ram_r[673] ),
    .S(_2271_),
    .X(_1700_));
 sg13g2_mux2_1 _7898_ (.A0(\logix.ram_r[675] ),
    .A1(\logix.ram_r[674] ),
    .S(net257),
    .X(_1701_));
 sg13g2_mux2_1 _7899_ (.A0(\logix.ram_r[676] ),
    .A1(\logix.ram_r[675] ),
    .S(net257),
    .X(_1702_));
 sg13g2_mux2_1 _7900_ (.A0(\logix.ram_r[677] ),
    .A1(\logix.ram_r[676] ),
    .S(net257),
    .X(_1703_));
 sg13g2_mux2_1 _7901_ (.A0(\logix.ram_r[678] ),
    .A1(\logix.ram_r[677] ),
    .S(net257),
    .X(_1704_));
 sg13g2_mux2_1 _7902_ (.A0(\logix.ram_r[679] ),
    .A1(\logix.ram_r[678] ),
    .S(net257),
    .X(_1705_));
 sg13g2_mux2_1 _7903_ (.A0(\logix.ram_r[67] ),
    .A1(\logix.ram_r[66] ),
    .S(net257),
    .X(_1706_));
 sg13g2_buf_1 _7904_ (.A(_2266_),
    .X(_2272_));
 sg13g2_mux2_1 _7905_ (.A0(\logix.ram_r[680] ),
    .A1(\logix.ram_r[679] ),
    .S(net256),
    .X(_1707_));
 sg13g2_mux2_1 _7906_ (.A0(\logix.ram_r[681] ),
    .A1(\logix.ram_r[680] ),
    .S(_2272_),
    .X(_1708_));
 sg13g2_mux2_1 _7907_ (.A0(\logix.ram_r[682] ),
    .A1(\logix.ram_r[681] ),
    .S(net256),
    .X(_1709_));
 sg13g2_mux2_1 _7908_ (.A0(\logix.ram_r[683] ),
    .A1(\logix.ram_r[682] ),
    .S(net256),
    .X(_1710_));
 sg13g2_mux2_1 _7909_ (.A0(\logix.ram_r[684] ),
    .A1(\logix.ram_r[683] ),
    .S(net256),
    .X(_1711_));
 sg13g2_mux2_1 _7910_ (.A0(\logix.ram_r[685] ),
    .A1(\logix.ram_r[684] ),
    .S(net256),
    .X(_1712_));
 sg13g2_mux2_1 _7911_ (.A0(\logix.ram_r[686] ),
    .A1(\logix.ram_r[685] ),
    .S(net256),
    .X(_1713_));
 sg13g2_mux2_1 _7912_ (.A0(\logix.ram_r[687] ),
    .A1(\logix.ram_r[686] ),
    .S(net256),
    .X(_1714_));
 sg13g2_mux2_1 _7913_ (.A0(\logix.ram_r[688] ),
    .A1(\logix.ram_r[687] ),
    .S(net256),
    .X(_1715_));
 sg13g2_mux2_1 _7914_ (.A0(\logix.ram_r[689] ),
    .A1(\logix.ram_r[688] ),
    .S(_2272_),
    .X(_1716_));
 sg13g2_buf_1 _7915_ (.A(_2266_),
    .X(_2273_));
 sg13g2_mux2_1 _7916_ (.A0(\logix.ram_r[68] ),
    .A1(\logix.ram_r[67] ),
    .S(_2273_),
    .X(_1717_));
 sg13g2_mux2_1 _7917_ (.A0(\logix.ram_r[690] ),
    .A1(\logix.ram_r[689] ),
    .S(_2273_),
    .X(_1718_));
 sg13g2_mux2_1 _7918_ (.A0(\logix.ram_r[691] ),
    .A1(\logix.ram_r[690] ),
    .S(net255),
    .X(_1719_));
 sg13g2_mux2_1 _7919_ (.A0(\logix.ram_r[692] ),
    .A1(\logix.ram_r[691] ),
    .S(net255),
    .X(_1720_));
 sg13g2_mux2_1 _7920_ (.A0(\logix.ram_r[693] ),
    .A1(\logix.ram_r[692] ),
    .S(net255),
    .X(_1721_));
 sg13g2_mux2_1 _7921_ (.A0(\logix.ram_r[694] ),
    .A1(\logix.ram_r[693] ),
    .S(net255),
    .X(_1722_));
 sg13g2_mux2_1 _7922_ (.A0(\logix.ram_r[695] ),
    .A1(\logix.ram_r[694] ),
    .S(net255),
    .X(_1723_));
 sg13g2_mux2_1 _7923_ (.A0(\logix.ram_r[696] ),
    .A1(\logix.ram_r[695] ),
    .S(net255),
    .X(_1724_));
 sg13g2_mux2_1 _7924_ (.A0(\logix.ram_r[697] ),
    .A1(\logix.ram_r[696] ),
    .S(net255),
    .X(_1725_));
 sg13g2_mux2_1 _7925_ (.A0(\logix.ram_r[698] ),
    .A1(\logix.ram_r[697] ),
    .S(net255),
    .X(_1726_));
 sg13g2_buf_1 _7926_ (.A(_2064_),
    .X(_2274_));
 sg13g2_buf_1 _7927_ (.A(_2274_),
    .X(_2275_));
 sg13g2_mux2_1 _7928_ (.A0(\logix.ram_r[699] ),
    .A1(\logix.ram_r[698] ),
    .S(_2275_),
    .X(_1727_));
 sg13g2_mux2_1 _7929_ (.A0(\logix.ram_r[69] ),
    .A1(\logix.ram_r[68] ),
    .S(net254),
    .X(_1728_));
 sg13g2_mux2_1 _7930_ (.A0(\logix.ram_r[6] ),
    .A1(\logix.ram_r[5] ),
    .S(_2275_),
    .X(_1729_));
 sg13g2_mux2_1 _7931_ (.A0(\logix.ram_r[700] ),
    .A1(\logix.ram_r[699] ),
    .S(net254),
    .X(_1730_));
 sg13g2_mux2_1 _7932_ (.A0(\logix.ram_r[701] ),
    .A1(\logix.ram_r[700] ),
    .S(net254),
    .X(_1731_));
 sg13g2_mux2_1 _7933_ (.A0(\logix.ram_r[702] ),
    .A1(\logix.ram_r[701] ),
    .S(net254),
    .X(_1732_));
 sg13g2_mux2_1 _7934_ (.A0(\logix.ram_r[703] ),
    .A1(\logix.ram_r[702] ),
    .S(net254),
    .X(_1733_));
 sg13g2_mux2_1 _7935_ (.A0(\logix.ram_r[704] ),
    .A1(\logix.ram_r[703] ),
    .S(net254),
    .X(_1734_));
 sg13g2_mux2_1 _7936_ (.A0(\logix.ram_r[705] ),
    .A1(\logix.ram_r[704] ),
    .S(net254),
    .X(_1735_));
 sg13g2_mux2_1 _7937_ (.A0(\logix.ram_r[706] ),
    .A1(\logix.ram_r[705] ),
    .S(net254),
    .X(_1736_));
 sg13g2_buf_1 _7938_ (.A(_2274_),
    .X(_2276_));
 sg13g2_mux2_1 _7939_ (.A0(\logix.ram_r[707] ),
    .A1(\logix.ram_r[706] ),
    .S(net253),
    .X(_1737_));
 sg13g2_mux2_1 _7940_ (.A0(\logix.ram_r[708] ),
    .A1(\logix.ram_r[707] ),
    .S(net253),
    .X(_1738_));
 sg13g2_mux2_1 _7941_ (.A0(\logix.ram_r[709] ),
    .A1(\logix.ram_r[708] ),
    .S(net253),
    .X(_1739_));
 sg13g2_mux2_1 _7942_ (.A0(\logix.ram_r[70] ),
    .A1(\logix.ram_r[69] ),
    .S(_2276_),
    .X(_1740_));
 sg13g2_mux2_1 _7943_ (.A0(\logix.ram_r[710] ),
    .A1(\logix.ram_r[709] ),
    .S(net253),
    .X(_1741_));
 sg13g2_mux2_1 _7944_ (.A0(\logix.ram_r[711] ),
    .A1(\logix.ram_r[710] ),
    .S(_2276_),
    .X(_1742_));
 sg13g2_mux2_1 _7945_ (.A0(\logix.ram_r[712] ),
    .A1(\logix.ram_r[711] ),
    .S(net253),
    .X(_1743_));
 sg13g2_mux2_1 _7946_ (.A0(\logix.ram_r[713] ),
    .A1(\logix.ram_r[712] ),
    .S(net253),
    .X(_1744_));
 sg13g2_mux2_1 _7947_ (.A0(\logix.ram_r[714] ),
    .A1(\logix.ram_r[713] ),
    .S(net253),
    .X(_1745_));
 sg13g2_mux2_1 _7948_ (.A0(\logix.ram_r[715] ),
    .A1(\logix.ram_r[714] ),
    .S(net253),
    .X(_1746_));
 sg13g2_buf_1 _7949_ (.A(_2274_),
    .X(_2277_));
 sg13g2_mux2_1 _7950_ (.A0(\logix.ram_r[716] ),
    .A1(\logix.ram_r[715] ),
    .S(net252),
    .X(_1747_));
 sg13g2_mux2_1 _7951_ (.A0(\logix.ram_r[717] ),
    .A1(\logix.ram_r[716] ),
    .S(net252),
    .X(_1748_));
 sg13g2_mux2_1 _7952_ (.A0(\logix.ram_r[718] ),
    .A1(\logix.ram_r[717] ),
    .S(net252),
    .X(_1749_));
 sg13g2_mux2_1 _7953_ (.A0(\logix.ram_r[719] ),
    .A1(\logix.ram_r[718] ),
    .S(_2277_),
    .X(_1750_));
 sg13g2_mux2_1 _7954_ (.A0(\logix.ram_r[71] ),
    .A1(\logix.ram_r[70] ),
    .S(_2277_),
    .X(_1751_));
 sg13g2_mux2_1 _7955_ (.A0(\logix.ram_r[720] ),
    .A1(\logix.ram_r[719] ),
    .S(net252),
    .X(_1752_));
 sg13g2_mux2_1 _7956_ (.A0(\logix.ram_r[721] ),
    .A1(\logix.ram_r[720] ),
    .S(net252),
    .X(_1753_));
 sg13g2_mux2_1 _7957_ (.A0(\logix.ram_r[722] ),
    .A1(\logix.ram_r[721] ),
    .S(net252),
    .X(_1754_));
 sg13g2_mux2_1 _7958_ (.A0(\logix.ram_r[723] ),
    .A1(\logix.ram_r[722] ),
    .S(net252),
    .X(_1755_));
 sg13g2_mux2_1 _7959_ (.A0(\logix.ram_r[724] ),
    .A1(\logix.ram_r[723] ),
    .S(net252),
    .X(_1756_));
 sg13g2_buf_1 _7960_ (.A(_2274_),
    .X(_2278_));
 sg13g2_mux2_1 _7961_ (.A0(\logix.ram_r[725] ),
    .A1(\logix.ram_r[724] ),
    .S(net251),
    .X(_1757_));
 sg13g2_mux2_1 _7962_ (.A0(\logix.ram_r[726] ),
    .A1(\logix.ram_r[725] ),
    .S(net251),
    .X(_1758_));
 sg13g2_mux2_1 _7963_ (.A0(\logix.ram_r[727] ),
    .A1(\logix.ram_r[726] ),
    .S(_2278_),
    .X(_1759_));
 sg13g2_mux2_1 _7964_ (.A0(\logix.ram_r[728] ),
    .A1(\logix.ram_r[727] ),
    .S(_2278_),
    .X(_1760_));
 sg13g2_mux2_1 _7965_ (.A0(\logix.ram_r[729] ),
    .A1(\logix.ram_r[728] ),
    .S(net251),
    .X(_1761_));
 sg13g2_mux2_1 _7966_ (.A0(\logix.ram_r[72] ),
    .A1(\logix.ram_r[71] ),
    .S(net251),
    .X(_1762_));
 sg13g2_mux2_1 _7967_ (.A0(\logix.ram_r[730] ),
    .A1(\logix.ram_r[729] ),
    .S(net251),
    .X(_1763_));
 sg13g2_mux2_1 _7968_ (.A0(\logix.ram_r[731] ),
    .A1(\logix.ram_r[730] ),
    .S(net251),
    .X(_1764_));
 sg13g2_mux2_1 _7969_ (.A0(\logix.ram_r[732] ),
    .A1(\logix.ram_r[731] ),
    .S(net251),
    .X(_1765_));
 sg13g2_mux2_1 _7970_ (.A0(\logix.ram_r[733] ),
    .A1(\logix.ram_r[732] ),
    .S(net251),
    .X(_1766_));
 sg13g2_buf_1 _7971_ (.A(_2274_),
    .X(_2279_));
 sg13g2_mux2_1 _7972_ (.A0(\logix.ram_r[734] ),
    .A1(\logix.ram_r[733] ),
    .S(net250),
    .X(_1767_));
 sg13g2_mux2_1 _7973_ (.A0(\logix.ram_r[735] ),
    .A1(\logix.ram_r[734] ),
    .S(net250),
    .X(_1768_));
 sg13g2_mux2_1 _7974_ (.A0(\logix.ram_r[736] ),
    .A1(\logix.ram_r[735] ),
    .S(net250),
    .X(_1769_));
 sg13g2_mux2_1 _7975_ (.A0(\logix.ram_r[737] ),
    .A1(\logix.ram_r[736] ),
    .S(net250),
    .X(_1770_));
 sg13g2_mux2_1 _7976_ (.A0(\logix.ram_r[738] ),
    .A1(\logix.ram_r[737] ),
    .S(_2279_),
    .X(_1771_));
 sg13g2_mux2_1 _7977_ (.A0(\logix.ram_r[739] ),
    .A1(\logix.ram_r[738] ),
    .S(net250),
    .X(_1772_));
 sg13g2_mux2_1 _7978_ (.A0(\logix.ram_r[73] ),
    .A1(\logix.ram_r[72] ),
    .S(_2279_),
    .X(_1773_));
 sg13g2_mux2_1 _7979_ (.A0(\logix.ram_r[740] ),
    .A1(\logix.ram_r[739] ),
    .S(net250),
    .X(_1774_));
 sg13g2_mux2_1 _7980_ (.A0(\logix.ram_r[741] ),
    .A1(\logix.ram_r[740] ),
    .S(net250),
    .X(_1775_));
 sg13g2_mux2_1 _7981_ (.A0(\logix.ram_r[742] ),
    .A1(\logix.ram_r[741] ),
    .S(net250),
    .X(_1776_));
 sg13g2_buf_1 _7982_ (.A(_2274_),
    .X(_2280_));
 sg13g2_mux2_1 _7983_ (.A0(\logix.ram_r[743] ),
    .A1(\logix.ram_r[742] ),
    .S(net249),
    .X(_1777_));
 sg13g2_mux2_1 _7984_ (.A0(\logix.ram_r[744] ),
    .A1(\logix.ram_r[743] ),
    .S(net249),
    .X(_1778_));
 sg13g2_mux2_1 _7985_ (.A0(\logix.ram_r[745] ),
    .A1(\logix.ram_r[744] ),
    .S(net249),
    .X(_1779_));
 sg13g2_mux2_1 _7986_ (.A0(\logix.ram_r[746] ),
    .A1(\logix.ram_r[745] ),
    .S(net249),
    .X(_1780_));
 sg13g2_mux2_1 _7987_ (.A0(\logix.ram_r[747] ),
    .A1(\logix.ram_r[746] ),
    .S(net249),
    .X(_1781_));
 sg13g2_mux2_1 _7988_ (.A0(\logix.ram_r[748] ),
    .A1(\logix.ram_r[747] ),
    .S(net249),
    .X(_1782_));
 sg13g2_mux2_1 _7989_ (.A0(\logix.ram_r[749] ),
    .A1(\logix.ram_r[748] ),
    .S(net249),
    .X(_1783_));
 sg13g2_mux2_1 _7990_ (.A0(\logix.ram_r[74] ),
    .A1(\logix.ram_r[73] ),
    .S(_2280_),
    .X(_1784_));
 sg13g2_mux2_1 _7991_ (.A0(\logix.ram_r[750] ),
    .A1(\logix.ram_r[749] ),
    .S(net249),
    .X(_1785_));
 sg13g2_mux2_1 _7992_ (.A0(\logix.ram_r[751] ),
    .A1(\logix.ram_r[750] ),
    .S(_2280_),
    .X(_1786_));
 sg13g2_buf_1 _7993_ (.A(_2274_),
    .X(_2281_));
 sg13g2_mux2_1 _7994_ (.A0(\logix.ram_r[752] ),
    .A1(\logix.ram_r[751] ),
    .S(net248),
    .X(_1787_));
 sg13g2_mux2_1 _7995_ (.A0(\logix.ram_r[753] ),
    .A1(\logix.ram_r[752] ),
    .S(net248),
    .X(_1788_));
 sg13g2_mux2_1 _7996_ (.A0(\logix.ram_r[754] ),
    .A1(\logix.ram_r[753] ),
    .S(net248),
    .X(_1789_));
 sg13g2_mux2_1 _7997_ (.A0(\logix.ram_r[755] ),
    .A1(\logix.ram_r[754] ),
    .S(net248),
    .X(_1790_));
 sg13g2_mux2_1 _7998_ (.A0(\logix.ram_r[756] ),
    .A1(\logix.ram_r[755] ),
    .S(net248),
    .X(_1791_));
 sg13g2_mux2_1 _7999_ (.A0(\logix.ram_r[757] ),
    .A1(\logix.ram_r[756] ),
    .S(net248),
    .X(_1792_));
 sg13g2_mux2_1 _8000_ (.A0(\logix.ram_r[758] ),
    .A1(\logix.ram_r[757] ),
    .S(net248),
    .X(_1793_));
 sg13g2_mux2_1 _8001_ (.A0(\logix.ram_r[759] ),
    .A1(\logix.ram_r[758] ),
    .S(_2281_),
    .X(_1794_));
 sg13g2_mux2_1 _8002_ (.A0(\logix.ram_r[75] ),
    .A1(\logix.ram_r[74] ),
    .S(_2281_),
    .X(_1795_));
 sg13g2_mux2_1 _8003_ (.A0(\logix.ram_r[760] ),
    .A1(\logix.ram_r[759] ),
    .S(net248),
    .X(_1796_));
 sg13g2_buf_1 _8004_ (.A(_2064_),
    .X(_2282_));
 sg13g2_buf_1 _8005_ (.A(_2282_),
    .X(_2283_));
 sg13g2_mux2_1 _8006_ (.A0(\logix.ram_r[761] ),
    .A1(\logix.ram_r[760] ),
    .S(net247),
    .X(_1797_));
 sg13g2_mux2_1 _8007_ (.A0(\logix.ram_r[762] ),
    .A1(\logix.ram_r[761] ),
    .S(net247),
    .X(_1798_));
 sg13g2_mux2_1 _8008_ (.A0(\logix.ram_r[763] ),
    .A1(\logix.ram_r[762] ),
    .S(net247),
    .X(_1799_));
 sg13g2_mux2_1 _8009_ (.A0(\logix.ram_r[764] ),
    .A1(\logix.ram_r[763] ),
    .S(net247),
    .X(_1800_));
 sg13g2_mux2_1 _8010_ (.A0(\logix.ram_r[765] ),
    .A1(\logix.ram_r[764] ),
    .S(net247),
    .X(_1801_));
 sg13g2_mux2_1 _8011_ (.A0(\logix.ram_r[766] ),
    .A1(\logix.ram_r[765] ),
    .S(net247),
    .X(_1802_));
 sg13g2_mux2_1 _8012_ (.A0(\logix.ram_r[767] ),
    .A1(\logix.ram_r[766] ),
    .S(net247),
    .X(_1803_));
 sg13g2_mux2_1 _8013_ (.A0(\logix.ram_r[768] ),
    .A1(\logix.ram_r[767] ),
    .S(_2283_),
    .X(_1804_));
 sg13g2_mux2_1 _8014_ (.A0(\logix.ram_r[769] ),
    .A1(\logix.ram_r[768] ),
    .S(_2283_),
    .X(_1805_));
 sg13g2_mux2_1 _8015_ (.A0(\logix.ram_r[76] ),
    .A1(\logix.ram_r[75] ),
    .S(net247),
    .X(_1806_));
 sg13g2_buf_1 _8016_ (.A(_2282_),
    .X(_2284_));
 sg13g2_mux2_1 _8017_ (.A0(\logix.ram_r[770] ),
    .A1(\logix.ram_r[769] ),
    .S(net246),
    .X(_1807_));
 sg13g2_mux2_1 _8018_ (.A0(\logix.ram_r[771] ),
    .A1(\logix.ram_r[770] ),
    .S(net246),
    .X(_1808_));
 sg13g2_mux2_1 _8019_ (.A0(\logix.ram_r[772] ),
    .A1(\logix.ram_r[771] ),
    .S(net246),
    .X(_1809_));
 sg13g2_mux2_1 _8020_ (.A0(\logix.ram_r[773] ),
    .A1(\logix.ram_r[772] ),
    .S(net246),
    .X(_1810_));
 sg13g2_mux2_1 _8021_ (.A0(\logix.ram_r[774] ),
    .A1(\logix.ram_r[773] ),
    .S(net246),
    .X(_1811_));
 sg13g2_mux2_1 _8022_ (.A0(\logix.ram_r[775] ),
    .A1(\logix.ram_r[774] ),
    .S(net246),
    .X(_1812_));
 sg13g2_mux2_1 _8023_ (.A0(\logix.ram_r[776] ),
    .A1(\logix.ram_r[775] ),
    .S(net246),
    .X(_1813_));
 sg13g2_mux2_1 _8024_ (.A0(\logix.ram_r[777] ),
    .A1(\logix.ram_r[776] ),
    .S(net246),
    .X(_1814_));
 sg13g2_mux2_1 _8025_ (.A0(\logix.ram_r[778] ),
    .A1(\logix.ram_r[777] ),
    .S(_2284_),
    .X(_1815_));
 sg13g2_mux2_1 _8026_ (.A0(\logix.ram_r[779] ),
    .A1(\logix.ram_r[778] ),
    .S(_2284_),
    .X(_1816_));
 sg13g2_buf_1 _8027_ (.A(_2282_),
    .X(_2285_));
 sg13g2_mux2_1 _8028_ (.A0(\logix.ram_r[77] ),
    .A1(\logix.ram_r[76] ),
    .S(_2285_),
    .X(_1817_));
 sg13g2_mux2_1 _8029_ (.A0(\logix.ram_r[780] ),
    .A1(\logix.ram_r[779] ),
    .S(net245),
    .X(_1818_));
 sg13g2_mux2_1 _8030_ (.A0(\logix.ram_r[781] ),
    .A1(\logix.ram_r[780] ),
    .S(net245),
    .X(_1819_));
 sg13g2_mux2_1 _8031_ (.A0(\logix.ram_r[782] ),
    .A1(\logix.ram_r[781] ),
    .S(net245),
    .X(_1820_));
 sg13g2_mux2_1 _8032_ (.A0(\logix.ram_r[783] ),
    .A1(\logix.ram_r[782] ),
    .S(net245),
    .X(_1821_));
 sg13g2_mux2_1 _8033_ (.A0(\logix.ram_r[784] ),
    .A1(\logix.ram_r[783] ),
    .S(net245),
    .X(_1822_));
 sg13g2_mux2_1 _8034_ (.A0(\logix.ram_r[785] ),
    .A1(\logix.ram_r[784] ),
    .S(net245),
    .X(_1823_));
 sg13g2_mux2_1 _8035_ (.A0(\logix.ram_r[786] ),
    .A1(\logix.ram_r[785] ),
    .S(net245),
    .X(_1824_));
 sg13g2_mux2_1 _8036_ (.A0(\logix.ram_r[787] ),
    .A1(\logix.ram_r[786] ),
    .S(_2285_),
    .X(_1825_));
 sg13g2_mux2_1 _8037_ (.A0(\logix.ram_r[788] ),
    .A1(\logix.ram_r[787] ),
    .S(net245),
    .X(_1826_));
 sg13g2_buf_1 _8038_ (.A(_2282_),
    .X(_2286_));
 sg13g2_mux2_1 _8039_ (.A0(\logix.ram_r[789] ),
    .A1(\logix.ram_r[788] ),
    .S(net244),
    .X(_1827_));
 sg13g2_mux2_1 _8040_ (.A0(\logix.ram_r[78] ),
    .A1(\logix.ram_r[77] ),
    .S(_2286_),
    .X(_1828_));
 sg13g2_mux2_1 _8041_ (.A0(\logix.ram_r[790] ),
    .A1(\logix.ram_r[789] ),
    .S(net244),
    .X(_1829_));
 sg13g2_mux2_1 _8042_ (.A0(\logix.ram_r[791] ),
    .A1(\logix.ram_r[790] ),
    .S(net244),
    .X(_1830_));
 sg13g2_mux2_1 _8043_ (.A0(\logix.ram_r[792] ),
    .A1(\logix.ram_r[791] ),
    .S(_2286_),
    .X(_1831_));
 sg13g2_mux2_1 _8044_ (.A0(\logix.ram_r[793] ),
    .A1(\logix.ram_r[792] ),
    .S(net244),
    .X(_1832_));
 sg13g2_mux2_1 _8045_ (.A0(\logix.ram_r[794] ),
    .A1(\logix.ram_r[793] ),
    .S(net244),
    .X(_1833_));
 sg13g2_mux2_1 _8046_ (.A0(\logix.ram_r[795] ),
    .A1(\logix.ram_r[794] ),
    .S(net244),
    .X(_1834_));
 sg13g2_mux2_1 _8047_ (.A0(\logix.ram_r[796] ),
    .A1(\logix.ram_r[795] ),
    .S(net244),
    .X(_1835_));
 sg13g2_mux2_1 _8048_ (.A0(\logix.ram_r[797] ),
    .A1(\logix.ram_r[796] ),
    .S(net244),
    .X(_1836_));
 sg13g2_buf_1 _8049_ (.A(_2282_),
    .X(_2287_));
 sg13g2_mux2_1 _8050_ (.A0(\logix.ram_r[798] ),
    .A1(\logix.ram_r[797] ),
    .S(net243),
    .X(_1837_));
 sg13g2_mux2_1 _8051_ (.A0(\logix.ram_r[799] ),
    .A1(\logix.ram_r[798] ),
    .S(net243),
    .X(_1838_));
 sg13g2_mux2_1 _8052_ (.A0(\logix.ram_r[79] ),
    .A1(\logix.ram_r[78] ),
    .S(net243),
    .X(_1839_));
 sg13g2_mux2_1 _8053_ (.A0(\logix.ram_r[7] ),
    .A1(\logix.ram_r[6] ),
    .S(net243),
    .X(_1840_));
 sg13g2_mux2_1 _8054_ (.A0(\logix.ram_r[800] ),
    .A1(\logix.ram_r[799] ),
    .S(net243),
    .X(_1841_));
 sg13g2_mux2_1 _8055_ (.A0(\logix.ram_r[801] ),
    .A1(\logix.ram_r[800] ),
    .S(net243),
    .X(_1842_));
 sg13g2_mux2_1 _8056_ (.A0(\logix.ram_r[802] ),
    .A1(\logix.ram_r[801] ),
    .S(net243),
    .X(_1843_));
 sg13g2_mux2_1 _8057_ (.A0(\logix.ram_r[803] ),
    .A1(\logix.ram_r[802] ),
    .S(net243),
    .X(_1844_));
 sg13g2_mux2_1 _8058_ (.A0(\logix.ram_r[804] ),
    .A1(\logix.ram_r[803] ),
    .S(_2287_),
    .X(_1845_));
 sg13g2_mux2_1 _8059_ (.A0(\logix.ram_r[805] ),
    .A1(\logix.ram_r[804] ),
    .S(_2287_),
    .X(_1846_));
 sg13g2_buf_1 _8060_ (.A(_2282_),
    .X(_2288_));
 sg13g2_mux2_1 _8061_ (.A0(\logix.ram_r[806] ),
    .A1(\logix.ram_r[805] ),
    .S(_2288_),
    .X(_1847_));
 sg13g2_mux2_1 _8062_ (.A0(\logix.ram_r[807] ),
    .A1(\logix.ram_r[806] ),
    .S(net242),
    .X(_1848_));
 sg13g2_mux2_1 _8063_ (.A0(\logix.ram_r[808] ),
    .A1(\logix.ram_r[807] ),
    .S(net242),
    .X(_1849_));
 sg13g2_mux2_1 _8064_ (.A0(\logix.ram_r[809] ),
    .A1(\logix.ram_r[808] ),
    .S(net242),
    .X(_1850_));
 sg13g2_mux2_1 _8065_ (.A0(\logix.ram_r[80] ),
    .A1(\logix.ram_r[79] ),
    .S(_2288_),
    .X(_1851_));
 sg13g2_mux2_1 _8066_ (.A0(\logix.ram_r[810] ),
    .A1(\logix.ram_r[809] ),
    .S(net242),
    .X(_1852_));
 sg13g2_mux2_1 _8067_ (.A0(\logix.ram_r[811] ),
    .A1(\logix.ram_r[810] ),
    .S(net242),
    .X(_1853_));
 sg13g2_mux2_1 _8068_ (.A0(\logix.ram_r[812] ),
    .A1(\logix.ram_r[811] ),
    .S(net242),
    .X(_1854_));
 sg13g2_mux2_1 _8069_ (.A0(\logix.ram_r[813] ),
    .A1(\logix.ram_r[812] ),
    .S(net242),
    .X(_1855_));
 sg13g2_mux2_1 _8070_ (.A0(\logix.ram_r[814] ),
    .A1(\logix.ram_r[813] ),
    .S(net242),
    .X(_1856_));
 sg13g2_buf_1 _8071_ (.A(_2282_),
    .X(_2289_));
 sg13g2_mux2_1 _8072_ (.A0(\logix.ram_r[815] ),
    .A1(\logix.ram_r[814] ),
    .S(net241),
    .X(_1857_));
 sg13g2_mux2_1 _8073_ (.A0(\logix.ram_r[816] ),
    .A1(\logix.ram_r[815] ),
    .S(net241),
    .X(_1858_));
 sg13g2_mux2_1 _8074_ (.A0(\logix.ram_r[817] ),
    .A1(\logix.ram_r[816] ),
    .S(net241),
    .X(_1859_));
 sg13g2_mux2_1 _8075_ (.A0(\logix.ram_r[818] ),
    .A1(\logix.ram_r[817] ),
    .S(net241),
    .X(_1860_));
 sg13g2_mux2_1 _8076_ (.A0(\logix.ram_r[819] ),
    .A1(\logix.ram_r[818] ),
    .S(_2289_),
    .X(_1861_));
 sg13g2_mux2_1 _8077_ (.A0(\logix.ram_r[81] ),
    .A1(\logix.ram_r[80] ),
    .S(net241),
    .X(_1862_));
 sg13g2_mux2_1 _8078_ (.A0(\logix.ram_r[820] ),
    .A1(\logix.ram_r[819] ),
    .S(net241),
    .X(_1863_));
 sg13g2_mux2_1 _8079_ (.A0(\logix.ram_r[821] ),
    .A1(\logix.ram_r[820] ),
    .S(_2289_),
    .X(_1864_));
 sg13g2_mux2_1 _8080_ (.A0(\logix.ram_r[822] ),
    .A1(\logix.ram_r[821] ),
    .S(net241),
    .X(_1865_));
 sg13g2_mux2_1 _8081_ (.A0(\logix.ram_r[823] ),
    .A1(\logix.ram_r[822] ),
    .S(net241),
    .X(_1866_));
 sg13g2_buf_1 _8082_ (.A(_2064_),
    .X(_2290_));
 sg13g2_buf_1 _8083_ (.A(_2290_),
    .X(_2291_));
 sg13g2_mux2_1 _8084_ (.A0(\logix.ram_r[824] ),
    .A1(\logix.ram_r[823] ),
    .S(net240),
    .X(_1867_));
 sg13g2_mux2_1 _8085_ (.A0(\logix.ram_r[825] ),
    .A1(\logix.ram_r[824] ),
    .S(net240),
    .X(_1868_));
 sg13g2_mux2_1 _8086_ (.A0(\logix.ram_r[826] ),
    .A1(\logix.ram_r[825] ),
    .S(net240),
    .X(_1869_));
 sg13g2_mux2_1 _8087_ (.A0(\logix.ram_r[827] ),
    .A1(\logix.ram_r[826] ),
    .S(net240),
    .X(_1870_));
 sg13g2_mux2_1 _8088_ (.A0(\logix.ram_r[828] ),
    .A1(\logix.ram_r[827] ),
    .S(net240),
    .X(_1871_));
 sg13g2_mux2_1 _8089_ (.A0(\logix.ram_r[829] ),
    .A1(\logix.ram_r[828] ),
    .S(net240),
    .X(_1872_));
 sg13g2_mux2_1 _8090_ (.A0(\logix.ram_r[82] ),
    .A1(\logix.ram_r[81] ),
    .S(_2291_),
    .X(_1873_));
 sg13g2_mux2_1 _8091_ (.A0(\logix.ram_r[830] ),
    .A1(\logix.ram_r[829] ),
    .S(net240),
    .X(_1874_));
 sg13g2_mux2_1 _8092_ (.A0(\logix.ram_r[831] ),
    .A1(\logix.ram_r[830] ),
    .S(net240),
    .X(_1875_));
 sg13g2_mux2_1 _8093_ (.A0(\logix.ram_r[832] ),
    .A1(\logix.ram_r[831] ),
    .S(_2291_),
    .X(_1876_));
 sg13g2_buf_1 _8094_ (.A(_2290_),
    .X(_2292_));
 sg13g2_mux2_1 _8095_ (.A0(\logix.ram_r[833] ),
    .A1(\logix.ram_r[832] ),
    .S(net239),
    .X(_1877_));
 sg13g2_mux2_1 _8096_ (.A0(\logix.ram_r[834] ),
    .A1(\logix.ram_r[833] ),
    .S(net239),
    .X(_1878_));
 sg13g2_mux2_1 _8097_ (.A0(\logix.ram_r[835] ),
    .A1(\logix.ram_r[834] ),
    .S(net239),
    .X(_1879_));
 sg13g2_mux2_1 _8098_ (.A0(\logix.ram_r[836] ),
    .A1(\logix.ram_r[835] ),
    .S(net239),
    .X(_1880_));
 sg13g2_mux2_1 _8099_ (.A0(\logix.ram_r[837] ),
    .A1(\logix.ram_r[836] ),
    .S(net239),
    .X(_1881_));
 sg13g2_mux2_1 _8100_ (.A0(\logix.ram_r[838] ),
    .A1(\logix.ram_r[837] ),
    .S(net239),
    .X(_1882_));
 sg13g2_mux2_1 _8101_ (.A0(\logix.ram_r[839] ),
    .A1(\logix.ram_r[838] ),
    .S(net239),
    .X(_1883_));
 sg13g2_mux2_1 _8102_ (.A0(\logix.ram_r[83] ),
    .A1(\logix.ram_r[82] ),
    .S(_2292_),
    .X(_1884_));
 sg13g2_mux2_1 _8103_ (.A0(\logix.ram_r[840] ),
    .A1(\logix.ram_r[839] ),
    .S(net239),
    .X(_1885_));
 sg13g2_mux2_1 _8104_ (.A0(\logix.ram_r[841] ),
    .A1(\logix.ram_r[840] ),
    .S(_2292_),
    .X(_1886_));
 sg13g2_buf_1 _8105_ (.A(_2290_),
    .X(_2293_));
 sg13g2_mux2_1 _8106_ (.A0(\logix.ram_r[842] ),
    .A1(\logix.ram_r[841] ),
    .S(net238),
    .X(_1887_));
 sg13g2_mux2_1 _8107_ (.A0(\logix.ram_r[843] ),
    .A1(\logix.ram_r[842] ),
    .S(net238),
    .X(_1888_));
 sg13g2_mux2_1 _8108_ (.A0(\logix.ram_r[844] ),
    .A1(\logix.ram_r[843] ),
    .S(_2293_),
    .X(_1889_));
 sg13g2_mux2_1 _8109_ (.A0(\logix.ram_r[845] ),
    .A1(\logix.ram_r[844] ),
    .S(net238),
    .X(_1890_));
 sg13g2_mux2_1 _8110_ (.A0(\logix.ram_r[846] ),
    .A1(\logix.ram_r[845] ),
    .S(net238),
    .X(_1891_));
 sg13g2_mux2_1 _8111_ (.A0(\logix.ram_r[847] ),
    .A1(\logix.ram_r[846] ),
    .S(net238),
    .X(_1892_));
 sg13g2_mux2_1 _8112_ (.A0(\logix.ram_r[848] ),
    .A1(\logix.ram_r[847] ),
    .S(net238),
    .X(_1893_));
 sg13g2_mux2_1 _8113_ (.A0(\logix.ram_r[849] ),
    .A1(\logix.ram_r[848] ),
    .S(_2293_),
    .X(_1894_));
 sg13g2_mux2_1 _8114_ (.A0(\logix.ram_r[84] ),
    .A1(\logix.ram_r[83] ),
    .S(net238),
    .X(_1895_));
 sg13g2_mux2_1 _8115_ (.A0(\logix.ram_r[850] ),
    .A1(\logix.ram_r[849] ),
    .S(net238),
    .X(_1896_));
 sg13g2_buf_1 _8116_ (.A(_2290_),
    .X(_2294_));
 sg13g2_mux2_1 _8117_ (.A0(\logix.ram_r[851] ),
    .A1(\logix.ram_r[850] ),
    .S(net237),
    .X(_1897_));
 sg13g2_mux2_1 _8118_ (.A0(\logix.ram_r[852] ),
    .A1(\logix.ram_r[851] ),
    .S(net237),
    .X(_1898_));
 sg13g2_mux2_1 _8119_ (.A0(\logix.ram_r[853] ),
    .A1(\logix.ram_r[852] ),
    .S(net237),
    .X(_1899_));
 sg13g2_mux2_1 _8120_ (.A0(\logix.ram_r[854] ),
    .A1(\logix.ram_r[853] ),
    .S(net237),
    .X(_1900_));
 sg13g2_mux2_1 _8121_ (.A0(\logix.ram_r[855] ),
    .A1(\logix.ram_r[854] ),
    .S(net237),
    .X(_1901_));
 sg13g2_mux2_1 _8122_ (.A0(\logix.ram_r[856] ),
    .A1(\logix.ram_r[855] ),
    .S(net237),
    .X(_1902_));
 sg13g2_mux2_1 _8123_ (.A0(\logix.ram_r[857] ),
    .A1(\logix.ram_r[856] ),
    .S(_2294_),
    .X(_1903_));
 sg13g2_mux2_1 _8124_ (.A0(\logix.ram_r[858] ),
    .A1(\logix.ram_r[857] ),
    .S(net237),
    .X(_1904_));
 sg13g2_mux2_1 _8125_ (.A0(\logix.ram_r[859] ),
    .A1(\logix.ram_r[858] ),
    .S(net237),
    .X(_1905_));
 sg13g2_mux2_1 _8126_ (.A0(\logix.ram_r[85] ),
    .A1(\logix.ram_r[84] ),
    .S(_2294_),
    .X(_1906_));
 sg13g2_buf_1 _8127_ (.A(_2290_),
    .X(_2295_));
 sg13g2_mux2_1 _8128_ (.A0(\logix.ram_r[860] ),
    .A1(\logix.ram_r[859] ),
    .S(net236),
    .X(_1907_));
 sg13g2_mux2_1 _8129_ (.A0(\logix.ram_r[861] ),
    .A1(\logix.ram_r[860] ),
    .S(net236),
    .X(_1908_));
 sg13g2_mux2_1 _8130_ (.A0(\logix.ram_r[862] ),
    .A1(\logix.ram_r[861] ),
    .S(net236),
    .X(_1909_));
 sg13g2_mux2_1 _8131_ (.A0(\logix.ram_r[863] ),
    .A1(\logix.ram_r[862] ),
    .S(net236),
    .X(_1910_));
 sg13g2_mux2_1 _8132_ (.A0(\logix.ram_r[864] ),
    .A1(\logix.ram_r[863] ),
    .S(_2295_),
    .X(_1911_));
 sg13g2_mux2_1 _8133_ (.A0(\logix.ram_r[865] ),
    .A1(\logix.ram_r[864] ),
    .S(net236),
    .X(_1912_));
 sg13g2_mux2_1 _8134_ (.A0(\logix.ram_r[866] ),
    .A1(\logix.ram_r[865] ),
    .S(_2295_),
    .X(_1913_));
 sg13g2_mux2_1 _8135_ (.A0(\logix.ram_r[867] ),
    .A1(\logix.ram_r[866] ),
    .S(net236),
    .X(_1914_));
 sg13g2_mux2_1 _8136_ (.A0(\logix.ram_r[868] ),
    .A1(\logix.ram_r[867] ),
    .S(net236),
    .X(_1915_));
 sg13g2_mux2_1 _8137_ (.A0(\logix.ram_r[869] ),
    .A1(\logix.ram_r[868] ),
    .S(net236),
    .X(_1916_));
 sg13g2_buf_1 _8138_ (.A(_2290_),
    .X(_2296_));
 sg13g2_mux2_1 _8139_ (.A0(\logix.ram_r[86] ),
    .A1(\logix.ram_r[85] ),
    .S(_2296_),
    .X(_1917_));
 sg13g2_mux2_1 _8140_ (.A0(\logix.ram_r[870] ),
    .A1(\logix.ram_r[869] ),
    .S(net235),
    .X(_1918_));
 sg13g2_mux2_1 _8141_ (.A0(\logix.ram_r[871] ),
    .A1(\logix.ram_r[870] ),
    .S(net235),
    .X(_1919_));
 sg13g2_mux2_1 _8142_ (.A0(\logix.ram_r[872] ),
    .A1(\logix.ram_r[871] ),
    .S(net235),
    .X(_1920_));
 sg13g2_mux2_1 _8143_ (.A0(\logix.ram_r[873] ),
    .A1(\logix.ram_r[872] ),
    .S(net235),
    .X(_1921_));
 sg13g2_mux2_1 _8144_ (.A0(\logix.ram_r[874] ),
    .A1(\logix.ram_r[873] ),
    .S(net235),
    .X(_1922_));
 sg13g2_mux2_1 _8145_ (.A0(\logix.ram_r[875] ),
    .A1(\logix.ram_r[874] ),
    .S(net235),
    .X(_1923_));
 sg13g2_mux2_1 _8146_ (.A0(\logix.ram_r[876] ),
    .A1(\logix.ram_r[875] ),
    .S(net235),
    .X(_1924_));
 sg13g2_mux2_1 _8147_ (.A0(\logix.ram_r[877] ),
    .A1(\logix.ram_r[876] ),
    .S(net235),
    .X(_1925_));
 sg13g2_mux2_1 _8148_ (.A0(\logix.ram_r[878] ),
    .A1(\logix.ram_r[877] ),
    .S(_2296_),
    .X(_1926_));
 sg13g2_buf_1 _8149_ (.A(_2290_),
    .X(_2297_));
 sg13g2_mux2_1 _8150_ (.A0(\logix.ram_r[879] ),
    .A1(\logix.ram_r[878] ),
    .S(net234),
    .X(_1927_));
 sg13g2_mux2_1 _8151_ (.A0(\logix.ram_r[87] ),
    .A1(\logix.ram_r[86] ),
    .S(_2297_),
    .X(_1928_));
 sg13g2_mux2_1 _8152_ (.A0(\logix.ram_r[880] ),
    .A1(\logix.ram_r[879] ),
    .S(net234),
    .X(_1929_));
 sg13g2_mux2_1 _8153_ (.A0(\logix.ram_r[881] ),
    .A1(\logix.ram_r[880] ),
    .S(net234),
    .X(_1930_));
 sg13g2_mux2_1 _8154_ (.A0(\logix.ram_r[882] ),
    .A1(\logix.ram_r[881] ),
    .S(net234),
    .X(_1931_));
 sg13g2_mux2_1 _8155_ (.A0(\logix.ram_r[883] ),
    .A1(\logix.ram_r[882] ),
    .S(net234),
    .X(_1932_));
 sg13g2_mux2_1 _8156_ (.A0(\logix.ram_r[884] ),
    .A1(\logix.ram_r[883] ),
    .S(net234),
    .X(_1933_));
 sg13g2_mux2_1 _8157_ (.A0(\logix.ram_r[885] ),
    .A1(\logix.ram_r[884] ),
    .S(net234),
    .X(_1934_));
 sg13g2_mux2_1 _8158_ (.A0(\logix.ram_r[886] ),
    .A1(\logix.ram_r[885] ),
    .S(net234),
    .X(_1935_));
 sg13g2_mux2_1 _8159_ (.A0(\logix.ram_r[887] ),
    .A1(\logix.ram_r[886] ),
    .S(_2297_),
    .X(_1936_));
 sg13g2_buf_1 _8160_ (.A(_2064_),
    .X(_2298_));
 sg13g2_buf_1 _8161_ (.A(_2298_),
    .X(_2299_));
 sg13g2_mux2_1 _8162_ (.A0(\logix.ram_r[888] ),
    .A1(\logix.ram_r[887] ),
    .S(net233),
    .X(_1937_));
 sg13g2_mux2_1 _8163_ (.A0(\logix.ram_r[889] ),
    .A1(\logix.ram_r[888] ),
    .S(net233),
    .X(_1938_));
 sg13g2_mux2_1 _8164_ (.A0(\logix.ram_r[88] ),
    .A1(\logix.ram_r[87] ),
    .S(_2299_),
    .X(_1939_));
 sg13g2_mux2_1 _8165_ (.A0(\logix.ram_r[890] ),
    .A1(\logix.ram_r[889] ),
    .S(net233),
    .X(_1940_));
 sg13g2_mux2_1 _8166_ (.A0(\logix.ram_r[891] ),
    .A1(\logix.ram_r[890] ),
    .S(net233),
    .X(_1941_));
 sg13g2_mux2_1 _8167_ (.A0(\logix.ram_r[892] ),
    .A1(\logix.ram_r[891] ),
    .S(net233),
    .X(_1942_));
 sg13g2_mux2_1 _8168_ (.A0(\logix.ram_r[893] ),
    .A1(\logix.ram_r[892] ),
    .S(net233),
    .X(_1943_));
 sg13g2_mux2_1 _8169_ (.A0(\logix.ram_r[894] ),
    .A1(\logix.ram_r[893] ),
    .S(net233),
    .X(_1944_));
 sg13g2_mux2_1 _8170_ (.A0(\logix.ram_r[895] ),
    .A1(\logix.ram_r[894] ),
    .S(_2299_),
    .X(_1945_));
 sg13g2_mux2_1 _8171_ (.A0(\logix.ram_r[896] ),
    .A1(\logix.ram_r[895] ),
    .S(net233),
    .X(_1946_));
 sg13g2_buf_1 _8172_ (.A(_2298_),
    .X(_2300_));
 sg13g2_mux2_1 _8173_ (.A0(\logix.ram_r[897] ),
    .A1(\logix.ram_r[896] ),
    .S(_2300_),
    .X(_1947_));
 sg13g2_mux2_1 _8174_ (.A0(\logix.ram_r[898] ),
    .A1(\logix.ram_r[897] ),
    .S(_2300_),
    .X(_1948_));
 sg13g2_mux2_1 _8175_ (.A0(\logix.ram_r[899] ),
    .A1(\logix.ram_r[898] ),
    .S(net232),
    .X(_1949_));
 sg13g2_mux2_1 _8176_ (.A0(\logix.ram_r[89] ),
    .A1(\logix.ram_r[88] ),
    .S(net232),
    .X(_1950_));
 sg13g2_mux2_1 _8177_ (.A0(\logix.ram_r[8] ),
    .A1(\logix.ram_r[7] ),
    .S(net232),
    .X(_1951_));
 sg13g2_mux2_1 _8178_ (.A0(\logix.ram_r[900] ),
    .A1(\logix.ram_r[899] ),
    .S(net232),
    .X(_1952_));
 sg13g2_mux2_1 _8179_ (.A0(\logix.ram_r[901] ),
    .A1(\logix.ram_r[900] ),
    .S(net232),
    .X(_1953_));
 sg13g2_mux2_1 _8180_ (.A0(\logix.ram_r[902] ),
    .A1(\logix.ram_r[901] ),
    .S(net232),
    .X(_1954_));
 sg13g2_mux2_1 _8181_ (.A0(\logix.ram_r[903] ),
    .A1(\logix.ram_r[902] ),
    .S(net232),
    .X(_1955_));
 sg13g2_mux2_1 _8182_ (.A0(\logix.ram_r[904] ),
    .A1(\logix.ram_r[903] ),
    .S(net232),
    .X(_1956_));
 sg13g2_buf_1 _8183_ (.A(_2298_),
    .X(_2301_));
 sg13g2_mux2_1 _8184_ (.A0(\logix.ram_r[905] ),
    .A1(\logix.ram_r[904] ),
    .S(_2301_),
    .X(_1957_));
 sg13g2_mux2_1 _8185_ (.A0(\logix.ram_r[906] ),
    .A1(\logix.ram_r[905] ),
    .S(net231),
    .X(_1958_));
 sg13g2_mux2_1 _8186_ (.A0(\logix.ram_r[907] ),
    .A1(\logix.ram_r[906] ),
    .S(net231),
    .X(_1959_));
 sg13g2_mux2_1 _8187_ (.A0(\logix.ram_r[908] ),
    .A1(\logix.ram_r[907] ),
    .S(net231),
    .X(_1960_));
 sg13g2_mux2_1 _8188_ (.A0(\logix.ram_r[909] ),
    .A1(\logix.ram_r[908] ),
    .S(net231),
    .X(_1961_));
 sg13g2_mux2_1 _8189_ (.A0(\logix.ram_r[90] ),
    .A1(\logix.ram_r[89] ),
    .S(net231),
    .X(_1962_));
 sg13g2_mux2_1 _8190_ (.A0(\logix.ram_r[910] ),
    .A1(\logix.ram_r[909] ),
    .S(net231),
    .X(_1963_));
 sg13g2_mux2_1 _8191_ (.A0(\logix.ram_r[911] ),
    .A1(\logix.ram_r[910] ),
    .S(net231),
    .X(_1964_));
 sg13g2_mux2_1 _8192_ (.A0(\logix.ram_r[912] ),
    .A1(\logix.ram_r[911] ),
    .S(net231),
    .X(_1965_));
 sg13g2_mux2_1 _8193_ (.A0(\logix.ram_r[913] ),
    .A1(\logix.ram_r[912] ),
    .S(_2301_),
    .X(_1966_));
 sg13g2_buf_1 _8194_ (.A(_2298_),
    .X(_2302_));
 sg13g2_mux2_1 _8195_ (.A0(\logix.ram_r[914] ),
    .A1(\logix.ram_r[913] ),
    .S(_2302_),
    .X(_1967_));
 sg13g2_mux2_1 _8196_ (.A0(\logix.ram_r[915] ),
    .A1(\logix.ram_r[914] ),
    .S(net230),
    .X(_1968_));
 sg13g2_mux2_1 _8197_ (.A0(\logix.ram_r[916] ),
    .A1(\logix.ram_r[915] ),
    .S(net230),
    .X(_1969_));
 sg13g2_mux2_1 _8198_ (.A0(\logix.ram_r[917] ),
    .A1(\logix.ram_r[916] ),
    .S(net230),
    .X(_1970_));
 sg13g2_mux2_1 _8199_ (.A0(\logix.ram_r[918] ),
    .A1(\logix.ram_r[917] ),
    .S(net230),
    .X(_1971_));
 sg13g2_mux2_1 _8200_ (.A0(\logix.ram_r[919] ),
    .A1(\logix.ram_r[918] ),
    .S(net230),
    .X(_1972_));
 sg13g2_mux2_1 _8201_ (.A0(\logix.ram_r[91] ),
    .A1(\logix.ram_r[90] ),
    .S(net230),
    .X(_1973_));
 sg13g2_mux2_1 _8202_ (.A0(\logix.ram_r[920] ),
    .A1(\logix.ram_r[919] ),
    .S(_2302_),
    .X(_1974_));
 sg13g2_mux2_1 _8203_ (.A0(\logix.ram_r[921] ),
    .A1(\logix.ram_r[920] ),
    .S(net230),
    .X(_1975_));
 sg13g2_mux2_1 _8204_ (.A0(\logix.ram_r[922] ),
    .A1(\logix.ram_r[921] ),
    .S(net230),
    .X(_1976_));
 sg13g2_buf_1 _8205_ (.A(_2298_),
    .X(_2303_));
 sg13g2_mux2_1 _8206_ (.A0(\logix.ram_r[923] ),
    .A1(\logix.ram_r[922] ),
    .S(_2303_),
    .X(_1977_));
 sg13g2_mux2_1 _8207_ (.A0(\logix.ram_r[924] ),
    .A1(\logix.ram_r[923] ),
    .S(net229),
    .X(_1978_));
 sg13g2_mux2_1 _8208_ (.A0(\logix.ram_r[925] ),
    .A1(\logix.ram_r[924] ),
    .S(net229),
    .X(_1979_));
 sg13g2_mux2_1 _8209_ (.A0(\logix.ram_r[926] ),
    .A1(\logix.ram_r[925] ),
    .S(net229),
    .X(_1980_));
 sg13g2_mux2_1 _8210_ (.A0(\logix.ram_r[927] ),
    .A1(\logix.ram_r[926] ),
    .S(net229),
    .X(_1981_));
 sg13g2_mux2_1 _8211_ (.A0(\logix.ram_r[928] ),
    .A1(\logix.ram_r[927] ),
    .S(net229),
    .X(_1982_));
 sg13g2_mux2_1 _8212_ (.A0(\logix.ram_r[929] ),
    .A1(\logix.ram_r[928] ),
    .S(net229),
    .X(_1983_));
 sg13g2_mux2_1 _8213_ (.A0(\logix.ram_r[92] ),
    .A1(\logix.ram_r[91] ),
    .S(_2303_),
    .X(_1984_));
 sg13g2_mux2_1 _8214_ (.A0(\logix.ram_r[930] ),
    .A1(\logix.ram_r[929] ),
    .S(net229),
    .X(_1985_));
 sg13g2_mux2_1 _8215_ (.A0(\logix.ram_r[931] ),
    .A1(\logix.ram_r[930] ),
    .S(net229),
    .X(_1986_));
 sg13g2_buf_1 _8216_ (.A(_2298_),
    .X(_2304_));
 sg13g2_mux2_1 _8217_ (.A0(\logix.ram_r[932] ),
    .A1(\logix.ram_r[931] ),
    .S(net228),
    .X(_1987_));
 sg13g2_mux2_1 _8218_ (.A0(\logix.ram_r[933] ),
    .A1(\logix.ram_r[932] ),
    .S(net228),
    .X(_1988_));
 sg13g2_mux2_1 _8219_ (.A0(\logix.ram_r[934] ),
    .A1(\logix.ram_r[933] ),
    .S(net228),
    .X(_1989_));
 sg13g2_mux2_1 _8220_ (.A0(\logix.ram_r[935] ),
    .A1(\logix.ram_r[934] ),
    .S(net228),
    .X(_1990_));
 sg13g2_mux2_1 _8221_ (.A0(\logix.ram_r[936] ),
    .A1(\logix.ram_r[935] ),
    .S(net228),
    .X(_1991_));
 sg13g2_mux2_1 _8222_ (.A0(\logix.ram_r[937] ),
    .A1(\logix.ram_r[936] ),
    .S(net228),
    .X(_1992_));
 sg13g2_mux2_1 _8223_ (.A0(\logix.ram_r[938] ),
    .A1(\logix.ram_r[937] ),
    .S(net228),
    .X(_1993_));
 sg13g2_mux2_1 _8224_ (.A0(\logix.ram_r[939] ),
    .A1(\logix.ram_r[938] ),
    .S(net228),
    .X(_1994_));
 sg13g2_mux2_1 _8225_ (.A0(\logix.ram_r[93] ),
    .A1(\logix.ram_r[92] ),
    .S(_2304_),
    .X(_1995_));
 sg13g2_mux2_1 _8226_ (.A0(\logix.ram_r[940] ),
    .A1(\logix.ram_r[939] ),
    .S(_2304_),
    .X(_1996_));
 sg13g2_buf_1 _8227_ (.A(_2298_),
    .X(_2305_));
 sg13g2_mux2_1 _8228_ (.A0(\logix.ram_r[941] ),
    .A1(\logix.ram_r[940] ),
    .S(net227),
    .X(_1997_));
 sg13g2_mux2_1 _8229_ (.A0(\logix.ram_r[942] ),
    .A1(\logix.ram_r[941] ),
    .S(net227),
    .X(_1998_));
 sg13g2_mux2_1 _8230_ (.A0(\logix.ram_r[943] ),
    .A1(\logix.ram_r[942] ),
    .S(net227),
    .X(_1999_));
 sg13g2_mux2_1 _8231_ (.A0(\logix.ram_r[944] ),
    .A1(\logix.ram_r[943] ),
    .S(net227),
    .X(_2000_));
 sg13g2_mux2_1 _8232_ (.A0(\logix.ram_r[945] ),
    .A1(\logix.ram_r[944] ),
    .S(net227),
    .X(_2001_));
 sg13g2_mux2_1 _8233_ (.A0(\logix.ram_r[946] ),
    .A1(\logix.ram_r[945] ),
    .S(net227),
    .X(_2002_));
 sg13g2_mux2_1 _8234_ (.A0(\logix.ram_r[947] ),
    .A1(\logix.ram_r[946] ),
    .S(net227),
    .X(_2003_));
 sg13g2_mux2_1 _8235_ (.A0(\logix.ram_r[948] ),
    .A1(\logix.ram_r[947] ),
    .S(net227),
    .X(_2004_));
 sg13g2_mux2_1 _8236_ (.A0(\logix.ram_r[949] ),
    .A1(\logix.ram_r[948] ),
    .S(_2305_),
    .X(_2005_));
 sg13g2_mux2_1 _8237_ (.A0(\logix.ram_r[94] ),
    .A1(\logix.ram_r[93] ),
    .S(_2305_),
    .X(_2006_));
 sg13g2_buf_1 _8238_ (.A(_2070_),
    .X(_2306_));
 sg13g2_mux2_1 _8239_ (.A0(\logix.ram_r[950] ),
    .A1(\logix.ram_r[949] ),
    .S(_2306_),
    .X(_2007_));
 sg13g2_mux2_1 _8240_ (.A0(\logix.ram_r[951] ),
    .A1(\logix.ram_r[950] ),
    .S(net226),
    .X(_2008_));
 sg13g2_mux2_1 _8241_ (.A0(\logix.ram_r[952] ),
    .A1(\logix.ram_r[951] ),
    .S(_2306_),
    .X(_2009_));
 sg13g2_mux2_1 _8242_ (.A0(\logix.ram_r[953] ),
    .A1(\logix.ram_r[952] ),
    .S(net226),
    .X(_2010_));
 sg13g2_mux2_1 _8243_ (.A0(\logix.ram_r[954] ),
    .A1(\logix.ram_r[953] ),
    .S(net226),
    .X(_2011_));
 sg13g2_mux2_1 _8244_ (.A0(\logix.ram_r[955] ),
    .A1(\logix.ram_r[954] ),
    .S(net226),
    .X(_2012_));
 sg13g2_mux2_1 _8245_ (.A0(\logix.ram_r[956] ),
    .A1(\logix.ram_r[955] ),
    .S(net226),
    .X(_2013_));
 sg13g2_mux2_1 _8246_ (.A0(\logix.ram_r[957] ),
    .A1(\logix.ram_r[956] ),
    .S(net226),
    .X(_2014_));
 sg13g2_mux2_1 _8247_ (.A0(\logix.ram_r[958] ),
    .A1(\logix.ram_r[957] ),
    .S(net226),
    .X(_2015_));
 sg13g2_mux2_1 _8248_ (.A0(\logix.ram_r[959] ),
    .A1(\logix.ram_r[958] ),
    .S(net226),
    .X(_2016_));
 sg13g2_buf_1 _8249_ (.A(_2070_),
    .X(_2307_));
 sg13g2_mux2_1 _8250_ (.A0(\logix.ram_r[95] ),
    .A1(\logix.ram_r[94] ),
    .S(net225),
    .X(_2017_));
 sg13g2_mux2_1 _8251_ (.A0(\logix.ram_r[960] ),
    .A1(\logix.ram_r[959] ),
    .S(net225),
    .X(_2018_));
 sg13g2_mux2_1 _8252_ (.A0(\logix.ram_r[961] ),
    .A1(\logix.ram_r[960] ),
    .S(net225),
    .X(_2019_));
 sg13g2_mux2_1 _8253_ (.A0(\logix.ram_r[962] ),
    .A1(\logix.ram_r[961] ),
    .S(net225),
    .X(_2020_));
 sg13g2_mux2_1 _8254_ (.A0(\logix.ram_r[963] ),
    .A1(\logix.ram_r[962] ),
    .S(net225),
    .X(_2021_));
 sg13g2_mux2_1 _8255_ (.A0(\logix.ram_r[964] ),
    .A1(\logix.ram_r[963] ),
    .S(net225),
    .X(_2022_));
 sg13g2_mux2_1 _8256_ (.A0(\logix.ram_r[965] ),
    .A1(\logix.ram_r[964] ),
    .S(_2307_),
    .X(_2023_));
 sg13g2_mux2_1 _8257_ (.A0(\logix.ram_r[966] ),
    .A1(\logix.ram_r[965] ),
    .S(_2307_),
    .X(_2024_));
 sg13g2_mux2_1 _8258_ (.A0(\logix.ram_r[967] ),
    .A1(\logix.ram_r[966] ),
    .S(net225),
    .X(_2025_));
 sg13g2_mux2_1 _8259_ (.A0(\logix.ram_r[968] ),
    .A1(\logix.ram_r[967] ),
    .S(net225),
    .X(_2026_));
 sg13g2_buf_1 _8260_ (.A(_2070_),
    .X(_2308_));
 sg13g2_mux2_1 _8261_ (.A0(\logix.ram_r[969] ),
    .A1(\logix.ram_r[968] ),
    .S(net224),
    .X(_2027_));
 sg13g2_mux2_1 _8262_ (.A0(\logix.ram_r[96] ),
    .A1(\logix.ram_r[95] ),
    .S(_2308_),
    .X(_2028_));
 sg13g2_mux2_1 _8263_ (.A0(\logix.ram_r[970] ),
    .A1(\logix.ram_r[969] ),
    .S(net224),
    .X(_2029_));
 sg13g2_mux2_1 _8264_ (.A0(\logix.ram_r[971] ),
    .A1(\logix.ram_r[970] ),
    .S(net224),
    .X(_2030_));
 sg13g2_mux2_1 _8265_ (.A0(\logix.ram_r[972] ),
    .A1(\logix.ram_r[971] ),
    .S(net224),
    .X(_2031_));
 sg13g2_mux2_1 _8266_ (.A0(\logix.ram_r[973] ),
    .A1(\logix.ram_r[972] ),
    .S(net224),
    .X(_2032_));
 sg13g2_mux2_1 _8267_ (.A0(\logix.ram_r[974] ),
    .A1(\logix.ram_r[973] ),
    .S(net224),
    .X(_2033_));
 sg13g2_mux2_1 _8268_ (.A0(\logix.ram_r[975] ),
    .A1(\logix.ram_r[974] ),
    .S(net224),
    .X(_2034_));
 sg13g2_mux2_1 _8269_ (.A0(\logix.ram_r[976] ),
    .A1(\logix.ram_r[975] ),
    .S(_2308_),
    .X(_2035_));
 sg13g2_mux2_1 _8270_ (.A0(\logix.ram_r[977] ),
    .A1(\logix.ram_r[976] ),
    .S(net224),
    .X(_2036_));
 sg13g2_buf_1 _8271_ (.A(_2070_),
    .X(_2309_));
 sg13g2_mux2_1 _8272_ (.A0(\logix.ram_r[978] ),
    .A1(\logix.ram_r[977] ),
    .S(_2309_),
    .X(_2037_));
 sg13g2_mux2_1 _8273_ (.A0(\logix.ram_r[979] ),
    .A1(\logix.ram_r[978] ),
    .S(net223),
    .X(_2038_));
 sg13g2_mux2_1 _8274_ (.A0(\logix.ram_r[97] ),
    .A1(\logix.ram_r[96] ),
    .S(_2309_),
    .X(_2039_));
 sg13g2_mux2_1 _8275_ (.A0(\logix.ram_r[980] ),
    .A1(\logix.ram_r[979] ),
    .S(net223),
    .X(_2040_));
 sg13g2_mux2_1 _8276_ (.A0(\logix.ram_r[981] ),
    .A1(\logix.ram_r[980] ),
    .S(net223),
    .X(_2041_));
 sg13g2_mux2_1 _8277_ (.A0(\logix.ram_r[982] ),
    .A1(\logix.ram_r[981] ),
    .S(net223),
    .X(_2042_));
 sg13g2_mux2_1 _8278_ (.A0(\logix.ram_r[983] ),
    .A1(\logix.ram_r[982] ),
    .S(net223),
    .X(_2043_));
 sg13g2_mux2_1 _8279_ (.A0(\logix.ram_r[984] ),
    .A1(\logix.ram_r[983] ),
    .S(net223),
    .X(_2044_));
 sg13g2_mux2_1 _8280_ (.A0(\logix.ram_r[985] ),
    .A1(\logix.ram_r[984] ),
    .S(net223),
    .X(_2045_));
 sg13g2_mux2_1 _8281_ (.A0(\logix.ram_r[986] ),
    .A1(\logix.ram_r[985] ),
    .S(net223),
    .X(_2046_));
 sg13g2_buf_1 _8282_ (.A(_2070_),
    .X(_2310_));
 sg13g2_mux2_1 _8283_ (.A0(\logix.ram_r[987] ),
    .A1(\logix.ram_r[986] ),
    .S(net222),
    .X(_2047_));
 sg13g2_mux2_1 _8284_ (.A0(\logix.ram_r[988] ),
    .A1(\logix.ram_r[987] ),
    .S(net222),
    .X(_2048_));
 sg13g2_mux2_1 _8285_ (.A0(\logix.ram_r[989] ),
    .A1(\logix.ram_r[988] ),
    .S(net222),
    .X(_2049_));
 sg13g2_mux2_1 _8286_ (.A0(\logix.ram_r[98] ),
    .A1(\logix.ram_r[97] ),
    .S(_2310_),
    .X(_2050_));
 sg13g2_mux2_1 _8287_ (.A0(\logix.ram_r[990] ),
    .A1(\logix.ram_r[989] ),
    .S(net222),
    .X(_2051_));
 sg13g2_mux2_1 _8288_ (.A0(\logix.ram_r[991] ),
    .A1(\logix.ram_r[990] ),
    .S(net222),
    .X(_2052_));
 sg13g2_mux2_1 _8289_ (.A0(\logix.ram_r[992] ),
    .A1(\logix.ram_r[991] ),
    .S(net222),
    .X(_2053_));
 sg13g2_mux2_1 _8290_ (.A0(\logix.ram_r[993] ),
    .A1(\logix.ram_r[992] ),
    .S(net222),
    .X(_2054_));
 sg13g2_mux2_1 _8291_ (.A0(\logix.ram_r[994] ),
    .A1(\logix.ram_r[993] ),
    .S(net222),
    .X(_2055_));
 sg13g2_mux2_1 _8292_ (.A0(\logix.ram_r[995] ),
    .A1(\logix.ram_r[994] ),
    .S(_2310_),
    .X(_2056_));
 sg13g2_mux2_1 _8293_ (.A0(\logix.ram_r[996] ),
    .A1(\logix.ram_r[995] ),
    .S(net413),
    .X(_2057_));
 sg13g2_mux2_1 _8294_ (.A0(\logix.ram_r[997] ),
    .A1(\logix.ram_r[996] ),
    .S(net413),
    .X(_2058_));
 sg13g2_mux2_1 _8295_ (.A0(\logix.ram_r[998] ),
    .A1(\logix.ram_r[997] ),
    .S(net413),
    .X(_2059_));
 sg13g2_mux2_1 _8296_ (.A0(\logix.ram_r[999] ),
    .A1(\logix.ram_r[998] ),
    .S(net413),
    .X(_2060_));
 sg13g2_mux2_1 _8297_ (.A0(\logix.ram_r[99] ),
    .A1(\logix.ram_r[98] ),
    .S(net413),
    .X(_2061_));
 sg13g2_mux2_1 _8298_ (.A0(\logix.ram_r[9] ),
    .A1(\logix.ram_r[8] ),
    .S(_2065_),
    .X(_2062_));
 sg13g2_nor4_1 _8299_ (.A(\logix.feedback_r[5] ),
    .B(\logix.feedback_r[4] ),
    .C(\logix.feedback_r[7] ),
    .D(\logix.feedback_r[6] ),
    .Y(_2311_));
 sg13g2_buf_2 _8300_ (.A(\logix.feedback_r[0] ),
    .X(_2312_));
 sg13g2_nor4_1 _8301_ (.A(\logix.feedback_r[1] ),
    .B(_2312_),
    .C(\logix.feedback_r[3] ),
    .D(\logix.feedback_r[2] ),
    .Y(_2313_));
 sg13g2_nand2_1 _8302_ (.Y(net11),
    .A(_2311_),
    .B(_2313_));
 sg13g2_nand4_1 _8303_ (.B(\logix.feedback_r[4] ),
    .C(\logix.feedback_r[7] ),
    .A(\logix.feedback_r[5] ),
    .Y(_2314_),
    .D(\logix.feedback_r[6] ));
 sg13g2_nand4_1 _8304_ (.B(_2312_),
    .C(\logix.feedback_r[3] ),
    .A(\logix.feedback_r[1] ),
    .Y(_2315_),
    .D(\logix.feedback_r[2] ));
 sg13g2_nor2_1 _8305_ (.A(_2314_),
    .B(_2315_),
    .Y(net12));
 sg13g2_xor2_1 _8306_ (.B(\logix.feedback_r[6] ),
    .A(\logix.feedback_r[7] ),
    .X(_2316_));
 sg13g2_xnor2_1 _8307_ (.Y(_2317_),
    .A(\logix.feedback_r[5] ),
    .B(\logix.feedback_r[4] ));
 sg13g2_xnor2_1 _8308_ (.Y(_2318_),
    .A(_2316_),
    .B(_2317_));
 sg13g2_xnor2_1 _8309_ (.Y(_2319_),
    .A(\logix.feedback_r[3] ),
    .B(\logix.feedback_r[2] ));
 sg13g2_xnor2_1 _8310_ (.Y(_2320_),
    .A(\logix.feedback_r[1] ),
    .B(_2312_));
 sg13g2_xnor2_1 _8311_ (.Y(_2321_),
    .A(_2319_),
    .B(_2320_));
 sg13g2_xnor2_1 _8312_ (.Y(net13),
    .A(_2318_),
    .B(_2321_));
 sg13g2_nand2b_1 _8313_ (.Y(_2322_),
    .B(_2206_),
    .A_N(_0001_));
 sg13g2_nand2b_1 _8314_ (.Y(_2323_),
    .B(net3),
    .A_N(_2206_));
 sg13g2_nand2_2 _8315_ (.Y(_2324_),
    .A(_2322_),
    .B(_2323_));
 sg13g2_buf_8 _8316_ (.A(_2324_),
    .X(_2325_));
 sg13g2_buf_1 _8317_ (.A(_2325_),
    .X(_2326_));
 sg13g2_buf_8 _8318_ (.A(net204),
    .X(_2327_));
 sg13g2_mux2_1 _8319_ (.A0(net1),
    .A1(_2312_),
    .S(_2204_),
    .X(_2328_));
 sg13g2_buf_8 _8320_ (.A(_2328_),
    .X(_2329_));
 sg13g2_buf_16 _8321_ (.X(_2330_),
    .A(_2329_));
 sg13g2_buf_16 _8322_ (.X(_2331_),
    .A(_2330_));
 sg13g2_buf_8 _8323_ (.A(_2331_),
    .X(_2332_));
 sg13g2_nor2_1 _8324_ (.A(net2),
    .B(_2205_),
    .Y(_2333_));
 sg13g2_and2_1 _8325_ (.A(_0000_),
    .B(_2205_),
    .X(_2334_));
 sg13g2_nor2_2 _8326_ (.A(_2333_),
    .B(_2334_),
    .Y(_2335_));
 sg13g2_buf_8 _8327_ (.A(_2335_),
    .X(_2336_));
 sg13g2_buf_8 _8328_ (.A(_2336_),
    .X(_2337_));
 sg13g2_buf_8 _8329_ (.A(_2337_),
    .X(_2338_));
 sg13g2_mux4_1 _8330_ (.S0(net178),
    .A0(\logix.ram_r[384] ),
    .A1(\logix.ram_r[392] ),
    .A2(\logix.ram_r[400] ),
    .A3(\logix.ram_r[408] ),
    .S1(net177),
    .X(_2339_));
 sg13g2_nor2_1 _8331_ (.A(net179),
    .B(_2339_),
    .Y(_2340_));
 sg13g2_nor2b_1 _8332_ (.A(_2204_),
    .B_N(net1),
    .Y(_2341_));
 sg13g2_a21oi_2 _8333_ (.B1(_2341_),
    .Y(_2342_),
    .A2(_2204_),
    .A1(_2312_));
 sg13g2_nand2_1 _8334_ (.Y(_2343_),
    .A(_2325_),
    .B(_2342_));
 sg13g2_buf_2 _8335_ (.A(_2343_),
    .X(_2344_));
 sg13g2_buf_8 _8336_ (.A(_2344_),
    .X(_2345_));
 sg13g2_buf_16 _8337_ (.X(_2346_),
    .A(_2336_));
 sg13g2_buf_8 _8338_ (.A(_2346_),
    .X(_2347_));
 sg13g2_mux2_1 _8339_ (.A0(\logix.ram_r[416] ),
    .A1(\logix.ram_r[432] ),
    .S(net176),
    .X(_2348_));
 sg13g2_nor2_1 _8340_ (.A(net83),
    .B(_2348_),
    .Y(_2349_));
 sg13g2_buf_16 _8341_ (.X(_2350_),
    .A(_2329_));
 sg13g2_nand2_1 _8342_ (.Y(_2351_),
    .A(_2324_),
    .B(_2350_));
 sg13g2_buf_2 _8343_ (.A(_2351_),
    .X(_2352_));
 sg13g2_buf_1 _8344_ (.A(_2352_),
    .X(_2353_));
 sg13g2_buf_16 _8345_ (.X(_2354_),
    .A(_2336_));
 sg13g2_buf_8 _8346_ (.A(_2354_),
    .X(_2355_));
 sg13g2_mux2_1 _8347_ (.A0(\logix.ram_r[424] ),
    .A1(\logix.ram_r[440] ),
    .S(net175),
    .X(_2356_));
 sg13g2_or2_1 _8348_ (.X(_2357_),
    .B(_2207_),
    .A(net4));
 sg13g2_buf_8 _8349_ (.A(_2357_),
    .X(_2358_));
 sg13g2_nand2_1 _8350_ (.Y(_2359_),
    .A(_0002_),
    .B(_2207_));
 sg13g2_buf_2 _8351_ (.A(_2359_),
    .X(_2360_));
 sg13g2_nand2_1 _8352_ (.Y(_2361_),
    .A(_2358_),
    .B(_2360_));
 sg13g2_buf_2 _8353_ (.A(_2361_),
    .X(_2362_));
 sg13g2_buf_2 _8354_ (.A(_2362_),
    .X(_2363_));
 sg13g2_o21ai_1 _8355_ (.B1(net174),
    .Y(_2364_),
    .A1(net82),
    .A2(_2356_));
 sg13g2_nor3_1 _8356_ (.A(_2340_),
    .B(_2349_),
    .C(_2364_),
    .Y(_2365_));
 sg13g2_or2_1 _8357_ (.X(_2366_),
    .B(_2206_),
    .A(net3));
 sg13g2_buf_1 _8358_ (.A(_2366_),
    .X(_2367_));
 sg13g2_nand2_1 _8359_ (.Y(_2368_),
    .A(_0001_),
    .B(_2206_));
 sg13g2_nand4_1 _8360_ (.B(_2368_),
    .C(_2358_),
    .A(_2367_),
    .Y(_2369_),
    .D(_2360_));
 sg13g2_buf_1 _8361_ (.A(_2369_),
    .X(_2370_));
 sg13g2_nor2_1 _8362_ (.A(_2336_),
    .B(_2370_),
    .Y(_2371_));
 sg13g2_buf_1 _8363_ (.A(_2371_),
    .X(_2372_));
 sg13g2_buf_1 _8364_ (.A(_2372_),
    .X(_2373_));
 sg13g2_buf_8 _8365_ (.A(_2350_),
    .X(_2374_));
 sg13g2_buf_8 _8366_ (.A(net203),
    .X(_2375_));
 sg13g2_mux2_1 _8367_ (.A0(\logix.ram_r[480] ),
    .A1(\logix.ram_r[488] ),
    .S(net173),
    .X(_2376_));
 sg13g2_or2_1 _8368_ (.X(_2377_),
    .B(_2334_),
    .A(_2333_));
 sg13g2_buf_2 _8369_ (.A(_2377_),
    .X(_2378_));
 sg13g2_nand4_1 _8370_ (.B(_2323_),
    .C(_2358_),
    .A(_2322_),
    .Y(_2379_),
    .D(_2360_));
 sg13g2_buf_1 _8371_ (.A(_2379_),
    .X(_2380_));
 sg13g2_nor2_1 _8372_ (.A(net207),
    .B(net202),
    .Y(_2381_));
 sg13g2_buf_2 _8373_ (.A(_2381_),
    .X(_2382_));
 sg13g2_buf_8 _8374_ (.A(_2382_),
    .X(_2383_));
 sg13g2_buf_8 _8375_ (.A(_2350_),
    .X(_2384_));
 sg13g2_buf_8 _8376_ (.A(net201),
    .X(_2385_));
 sg13g2_mux2_1 _8377_ (.A0(\logix.ram_r[464] ),
    .A1(\logix.ram_r[472] ),
    .S(net172),
    .X(_2386_));
 sg13g2_a22oi_1 _8378_ (.Y(_2387_),
    .B1(net47),
    .B2(_2386_),
    .A2(_2376_),
    .A1(_2373_));
 sg13g2_nor2_1 _8379_ (.A(_2336_),
    .B(net202),
    .Y(_2388_));
 sg13g2_buf_8 _8380_ (.A(_2388_),
    .X(_2389_));
 sg13g2_buf_8 _8381_ (.A(_2389_),
    .X(_2390_));
 sg13g2_buf_8 _8382_ (.A(_2330_),
    .X(_2391_));
 sg13g2_buf_8 _8383_ (.A(_2391_),
    .X(_2392_));
 sg13g2_mux2_1 _8384_ (.A0(\logix.ram_r[448] ),
    .A1(\logix.ram_r[456] ),
    .S(net171),
    .X(_2393_));
 sg13g2_nor2_1 _8385_ (.A(net207),
    .B(_2370_),
    .Y(_2394_));
 sg13g2_buf_1 _8386_ (.A(_2394_),
    .X(_2395_));
 sg13g2_buf_1 _8387_ (.A(_2395_),
    .X(_2396_));
 sg13g2_mux2_1 _8388_ (.A0(\logix.ram_r[496] ),
    .A1(\logix.ram_r[504] ),
    .S(net172),
    .X(_2397_));
 sg13g2_a22oi_1 _8389_ (.Y(_2398_),
    .B1(net45),
    .B2(_2397_),
    .A2(_2393_),
    .A1(net46));
 sg13g2_nand2_1 _8390_ (.Y(_2399_),
    .A(_2387_),
    .B(_2398_));
 sg13g2_nor2_1 _8391_ (.A(net6),
    .B(_2209_),
    .Y(_2400_));
 sg13g2_a21o_1 _8392_ (.A2(_2209_),
    .A1(_0004_),
    .B1(_2400_),
    .X(_2401_));
 sg13g2_buf_1 _8393_ (.A(_2401_),
    .X(_2402_));
 sg13g2_nor2_1 _8394_ (.A(net5),
    .B(_2208_),
    .Y(_2403_));
 sg13g2_a21o_1 _8395_ (.A2(_2208_),
    .A1(_0003_),
    .B1(_2403_),
    .X(_2404_));
 sg13g2_buf_1 _8396_ (.A(_2404_),
    .X(_2405_));
 sg13g2_nor2_1 _8397_ (.A(_2402_),
    .B(_2405_),
    .Y(_2406_));
 sg13g2_buf_1 _8398_ (.A(_2406_),
    .X(_2407_));
 sg13g2_buf_1 _8399_ (.A(_2407_),
    .X(_2408_));
 sg13g2_o21ai_1 _8400_ (.B1(net81),
    .Y(_2409_),
    .A1(_2365_),
    .A2(_2399_));
 sg13g2_and2_1 _8401_ (.A(_2358_),
    .B(_2360_),
    .X(_2410_));
 sg13g2_buf_2 _8402_ (.A(_2410_),
    .X(_2411_));
 sg13g2_buf_1 _8403_ (.A(_2411_),
    .X(_2412_));
 sg13g2_buf_8 _8404_ (.A(_2337_),
    .X(_2413_));
 sg13g2_buf_2 _8405_ (.A(_2325_),
    .X(_2414_));
 sg13g2_mux4_1 _8406_ (.S0(net168),
    .A0(\logix.ram_r[256] ),
    .A1(\logix.ram_r[272] ),
    .A2(\logix.ram_r[288] ),
    .A3(\logix.ram_r[304] ),
    .S1(net199),
    .X(_2415_));
 sg13g2_buf_8 _8407_ (.A(_2336_),
    .X(_2416_));
 sg13g2_buf_8 _8408_ (.A(_2416_),
    .X(_2417_));
 sg13g2_mux4_1 _8409_ (.S0(net167),
    .A0(\logix.ram_r[264] ),
    .A1(\logix.ram_r[280] ),
    .A2(\logix.ram_r[296] ),
    .A3(\logix.ram_r[312] ),
    .S1(net199),
    .X(_2418_));
 sg13g2_buf_8 _8410_ (.A(_2331_),
    .X(_2419_));
 sg13g2_buf_8 _8411_ (.A(net166),
    .X(_2420_));
 sg13g2_buf_8 _8412_ (.A(_2420_),
    .X(_2421_));
 sg13g2_mux2_1 _8413_ (.A0(_2415_),
    .A1(_2418_),
    .S(_2421_),
    .X(_2422_));
 sg13g2_buf_1 _8414_ (.A(net202),
    .X(_2423_));
 sg13g2_buf_8 _8415_ (.A(_2330_),
    .X(_2424_));
 sg13g2_buf_8 _8416_ (.A(net198),
    .X(_2425_));
 sg13g2_buf_8 _8417_ (.A(_2336_),
    .X(_2426_));
 sg13g2_buf_8 _8418_ (.A(_2426_),
    .X(_2427_));
 sg13g2_mux4_1 _8419_ (.S0(net164),
    .A0(\logix.ram_r[320] ),
    .A1(\logix.ram_r[328] ),
    .A2(\logix.ram_r[336] ),
    .A3(\logix.ram_r[344] ),
    .S1(_2427_),
    .X(_2428_));
 sg13g2_nor2_1 _8420_ (.A(_2423_),
    .B(_2428_),
    .Y(_2429_));
 sg13g2_and4_1 _8421_ (.A(_2367_),
    .B(_2368_),
    .C(_2358_),
    .D(_2360_),
    .X(_2430_));
 sg13g2_buf_8 _8422_ (.A(_2430_),
    .X(_2431_));
 sg13g2_nand2_1 _8423_ (.Y(_2432_),
    .A(net198),
    .B(_2431_));
 sg13g2_buf_2 _8424_ (.A(_2432_),
    .X(_2433_));
 sg13g2_buf_8 _8425_ (.A(_2433_),
    .X(_2434_));
 sg13g2_buf_8 _8426_ (.A(_2426_),
    .X(_2435_));
 sg13g2_mux2_1 _8427_ (.A0(\logix.ram_r[360] ),
    .A1(\logix.ram_r[376] ),
    .S(net162),
    .X(_2436_));
 sg13g2_nor2_1 _8428_ (.A(net43),
    .B(_2436_),
    .Y(_2437_));
 sg13g2_nand2_1 _8429_ (.Y(_2438_),
    .A(_2342_),
    .B(_2431_));
 sg13g2_buf_2 _8430_ (.A(_2438_),
    .X(_2439_));
 sg13g2_buf_8 _8431_ (.A(_2439_),
    .X(_2440_));
 sg13g2_mux2_1 _8432_ (.A0(\logix.ram_r[352] ),
    .A1(\logix.ram_r[368] ),
    .S(net176),
    .X(_2441_));
 sg13g2_a21oi_2 _8433_ (.B1(_2403_),
    .Y(_2442_),
    .A2(_2208_),
    .A1(_0003_));
 sg13g2_nor2_1 _8434_ (.A(_2402_),
    .B(_2442_),
    .Y(_2443_));
 sg13g2_buf_2 _8435_ (.A(_2443_),
    .X(_2444_));
 sg13g2_buf_8 _8436_ (.A(_2444_),
    .X(_2445_));
 sg13g2_o21ai_1 _8437_ (.B1(net79),
    .Y(_2446_),
    .A1(_2440_),
    .A2(_2441_));
 sg13g2_nor3_1 _8438_ (.A(_2429_),
    .B(_2437_),
    .C(_2446_),
    .Y(_2447_));
 sg13g2_o21ai_1 _8439_ (.B1(_2447_),
    .Y(_2448_),
    .A1(net169),
    .A2(_2422_));
 sg13g2_nor2_1 _8440_ (.A(net8),
    .B(_2212_),
    .Y(_2449_));
 sg13g2_a21o_1 _8441_ (.A2(_2212_),
    .A1(_0006_),
    .B1(_2449_),
    .X(_2450_));
 sg13g2_buf_1 _8442_ (.A(_2450_),
    .X(_2451_));
 sg13g2_nand2_1 _8443_ (.Y(_2452_),
    .A(_0005_),
    .B(_2211_));
 sg13g2_o21ai_1 _8444_ (.B1(_2452_),
    .Y(_2453_),
    .A1(net7),
    .A2(_2211_));
 sg13g2_buf_2 _8445_ (.A(_2453_),
    .X(_2454_));
 sg13g2_nand2_2 _8446_ (.Y(_2455_),
    .A(_2451_),
    .B(_2454_));
 sg13g2_inv_4 _8447_ (.A(_2455_),
    .Y(_2456_));
 sg13g2_nand2_1 _8448_ (.Y(_2457_),
    .A(_2367_),
    .B(_2368_));
 sg13g2_buf_2 _8449_ (.A(_2457_),
    .X(_2458_));
 sg13g2_nor2_1 _8450_ (.A(_2458_),
    .B(_2411_),
    .Y(_2459_));
 sg13g2_buf_8 _8451_ (.A(_2459_),
    .X(_2460_));
 sg13g2_buf_8 _8452_ (.A(net78),
    .X(_2461_));
 sg13g2_buf_16 _8453_ (.X(_2462_),
    .A(_2330_));
 sg13g2_buf_8 _8454_ (.A(_2462_),
    .X(_2463_));
 sg13g2_mux4_1 _8455_ (.S0(net161),
    .A0(\logix.ram_r[32] ),
    .A1(\logix.ram_r[40] ),
    .A2(\logix.ram_r[48] ),
    .A3(\logix.ram_r[56] ),
    .S1(net168),
    .X(_2464_));
 sg13g2_nor2_1 _8456_ (.A(_2324_),
    .B(_2411_),
    .Y(_2465_));
 sg13g2_buf_8 _8457_ (.A(_2465_),
    .X(_2466_));
 sg13g2_buf_8 _8458_ (.A(net77),
    .X(_2467_));
 sg13g2_buf_8 _8459_ (.A(net198),
    .X(_2468_));
 sg13g2_buf_8 _8460_ (.A(_2426_),
    .X(_2469_));
 sg13g2_mux4_1 _8461_ (.S0(net160),
    .A0(\logix.ram_r[0] ),
    .A1(\logix.ram_r[8] ),
    .A2(\logix.ram_r[16] ),
    .A3(\logix.ram_r[24] ),
    .S1(net159),
    .X(_2470_));
 sg13g2_a22oi_1 _8462_ (.Y(_2471_),
    .B1(net40),
    .B2(_2470_),
    .A2(_2464_),
    .A1(net41));
 sg13g2_buf_8 _8463_ (.A(_2431_),
    .X(_2472_));
 sg13g2_buf_2 _8464_ (.A(net158),
    .X(_2473_));
 sg13g2_buf_8 _8465_ (.A(_2462_),
    .X(_2474_));
 sg13g2_buf_8 _8466_ (.A(_2416_),
    .X(_2475_));
 sg13g2_mux4_1 _8467_ (.S0(net157),
    .A0(\logix.ram_r[96] ),
    .A1(\logix.ram_r[104] ),
    .A2(\logix.ram_r[112] ),
    .A3(\logix.ram_r[120] ),
    .S1(net156),
    .X(_2476_));
 sg13g2_buf_8 _8468_ (.A(_2331_),
    .X(_2477_));
 sg13g2_mux4_1 _8469_ (.S0(net155),
    .A0(\logix.ram_r[64] ),
    .A1(\logix.ram_r[72] ),
    .A2(\logix.ram_r[80] ),
    .A3(\logix.ram_r[88] ),
    .S1(_2435_),
    .X(_2478_));
 sg13g2_and4_1 _8470_ (.A(_2322_),
    .B(_2323_),
    .C(_2358_),
    .D(_2360_),
    .X(_2479_));
 sg13g2_buf_2 _8471_ (.A(_2479_),
    .X(_2480_));
 sg13g2_buf_8 _8472_ (.A(_2480_),
    .X(_2481_));
 sg13g2_buf_1 _8473_ (.A(net154),
    .X(_2482_));
 sg13g2_a22oi_1 _8474_ (.Y(_2483_),
    .B1(_2478_),
    .B2(net75),
    .A2(_2476_),
    .A1(net76));
 sg13g2_nand2_1 _8475_ (.Y(_2484_),
    .A(_2402_),
    .B(_2405_));
 sg13g2_buf_1 _8476_ (.A(_2484_),
    .X(_2485_));
 sg13g2_buf_2 _8477_ (.A(_2485_),
    .X(_2486_));
 sg13g2_a21oi_1 _8478_ (.A1(_2471_),
    .A2(_2483_),
    .Y(_2487_),
    .B1(_2486_));
 sg13g2_buf_8 _8479_ (.A(net78),
    .X(_2488_));
 sg13g2_buf_8 _8480_ (.A(_2337_),
    .X(_2489_));
 sg13g2_mux4_1 _8481_ (.S0(net178),
    .A0(\logix.ram_r[160] ),
    .A1(\logix.ram_r[168] ),
    .A2(\logix.ram_r[176] ),
    .A3(\logix.ram_r[184] ),
    .S1(net153),
    .X(_2490_));
 sg13g2_mux4_1 _8482_ (.S0(net160),
    .A0(\logix.ram_r[128] ),
    .A1(\logix.ram_r[136] ),
    .A2(\logix.ram_r[144] ),
    .A3(\logix.ram_r[152] ),
    .S1(net163),
    .X(_2491_));
 sg13g2_buf_8 _8483_ (.A(net77),
    .X(_2492_));
 sg13g2_a22oi_1 _8484_ (.Y(_2493_),
    .B1(_2491_),
    .B2(net38),
    .A2(_2490_),
    .A1(net39));
 sg13g2_buf_1 _8485_ (.A(net158),
    .X(_2494_));
 sg13g2_mux4_1 _8486_ (.S0(net161),
    .A0(\logix.ram_r[224] ),
    .A1(\logix.ram_r[232] ),
    .A2(\logix.ram_r[240] ),
    .A3(\logix.ram_r[248] ),
    .S1(net168),
    .X(_2495_));
 sg13g2_buf_8 _8487_ (.A(_2424_),
    .X(_2496_));
 sg13g2_buf_8 _8488_ (.A(_2426_),
    .X(_2497_));
 sg13g2_mux4_1 _8489_ (.S0(net152),
    .A0(\logix.ram_r[192] ),
    .A1(\logix.ram_r[200] ),
    .A2(\logix.ram_r[208] ),
    .A3(\logix.ram_r[216] ),
    .S1(net151),
    .X(_2498_));
 sg13g2_buf_2 _8490_ (.A(net154),
    .X(_2499_));
 sg13g2_a22oi_1 _8491_ (.Y(_2500_),
    .B1(_2498_),
    .B2(net72),
    .A2(_2495_),
    .A1(net73));
 sg13g2_nand2_1 _8492_ (.Y(_2501_),
    .A(_2402_),
    .B(_2442_));
 sg13g2_buf_2 _8493_ (.A(_2501_),
    .X(_2502_));
 sg13g2_buf_2 _8494_ (.A(_2502_),
    .X(_2503_));
 sg13g2_a21oi_1 _8495_ (.A1(_2493_),
    .A2(_2500_),
    .Y(_2504_),
    .B1(net71));
 sg13g2_nor2_1 _8496_ (.A(_2487_),
    .B(_2504_),
    .Y(_2505_));
 sg13g2_nand4_1 _8497_ (.B(_2448_),
    .C(_2456_),
    .A(_2409_),
    .Y(_2506_),
    .D(_2505_));
 sg13g2_buf_8 _8498_ (.A(net204),
    .X(_2507_));
 sg13g2_buf_8 _8499_ (.A(_2462_),
    .X(_2508_));
 sg13g2_buf_8 _8500_ (.A(_2416_),
    .X(_2509_));
 sg13g2_mux4_1 _8501_ (.S0(net149),
    .A0(\logix.ram_r[896] ),
    .A1(\logix.ram_r[904] ),
    .A2(\logix.ram_r[912] ),
    .A3(\logix.ram_r[920] ),
    .S1(net148),
    .X(_2510_));
 sg13g2_nor2_1 _8502_ (.A(_2507_),
    .B(_2510_),
    .Y(_2511_));
 sg13g2_buf_8 _8503_ (.A(_2346_),
    .X(_2512_));
 sg13g2_mux2_1 _8504_ (.A0(\logix.ram_r[928] ),
    .A1(\logix.ram_r[944] ),
    .S(net147),
    .X(_2513_));
 sg13g2_nor2_1 _8505_ (.A(net83),
    .B(_2513_),
    .Y(_2514_));
 sg13g2_buf_8 _8506_ (.A(_2335_),
    .X(_2515_));
 sg13g2_buf_2 _8507_ (.A(_2515_),
    .X(_2516_));
 sg13g2_mux2_1 _8508_ (.A0(\logix.ram_r[936] ),
    .A1(\logix.ram_r[952] ),
    .S(net197),
    .X(_2517_));
 sg13g2_o21ai_1 _8509_ (.B1(net174),
    .Y(_2518_),
    .A1(net82),
    .A2(_2517_));
 sg13g2_nor3_1 _8510_ (.A(_2511_),
    .B(_2514_),
    .C(_2518_),
    .Y(_2519_));
 sg13g2_buf_1 _8511_ (.A(_2372_),
    .X(_2520_));
 sg13g2_buf_8 _8512_ (.A(net200),
    .X(_2521_));
 sg13g2_mux2_1 _8513_ (.A0(\logix.ram_r[992] ),
    .A1(\logix.ram_r[1000] ),
    .S(net146),
    .X(_2522_));
 sg13g2_buf_8 _8514_ (.A(_2350_),
    .X(_2523_));
 sg13g2_buf_8 _8515_ (.A(_2523_),
    .X(_2524_));
 sg13g2_mux2_1 _8516_ (.A0(\logix.ram_r[976] ),
    .A1(\logix.ram_r[984] ),
    .S(net145),
    .X(_2525_));
 sg13g2_a22oi_1 _8517_ (.Y(_2526_),
    .B1(_2525_),
    .B2(_2383_),
    .A2(_2522_),
    .A1(net37));
 sg13g2_buf_8 _8518_ (.A(_2330_),
    .X(_2527_));
 sg13g2_buf_8 _8519_ (.A(net195),
    .X(_2528_));
 sg13g2_mux2_1 _8520_ (.A0(\logix.ram_r[960] ),
    .A1(\logix.ram_r[968] ),
    .S(_2528_),
    .X(_2529_));
 sg13g2_mux2_1 _8521_ (.A0(\logix.ram_r[1008] ),
    .A1(\logix.ram_r[1016] ),
    .S(net173),
    .X(_2530_));
 sg13g2_a22oi_1 _8522_ (.Y(_2531_),
    .B1(_2530_),
    .B2(net45),
    .A2(_2529_),
    .A1(net46));
 sg13g2_nand2_1 _8523_ (.Y(_2532_),
    .A(_2526_),
    .B(_2531_));
 sg13g2_o21ai_1 _8524_ (.B1(net81),
    .Y(_2533_),
    .A1(_2519_),
    .A2(_2532_));
 sg13g2_buf_8 _8525_ (.A(_2416_),
    .X(_2534_));
 sg13g2_buf_2 _8526_ (.A(_2325_),
    .X(_2535_));
 sg13g2_mux4_1 _8527_ (.S0(net143),
    .A0(\logix.ram_r[768] ),
    .A1(\logix.ram_r[784] ),
    .A2(\logix.ram_r[800] ),
    .A3(\logix.ram_r[816] ),
    .S1(net194),
    .X(_2536_));
 sg13g2_buf_8 _8528_ (.A(_2416_),
    .X(_2537_));
 sg13g2_mux4_1 _8529_ (.S0(_2537_),
    .A0(\logix.ram_r[776] ),
    .A1(\logix.ram_r[792] ),
    .A2(\logix.ram_r[808] ),
    .A3(\logix.ram_r[824] ),
    .S1(net194),
    .X(_2538_));
 sg13g2_mux2_1 _8530_ (.A0(_2536_),
    .A1(_2538_),
    .S(net44),
    .X(_2539_));
 sg13g2_buf_8 _8531_ (.A(net198),
    .X(_2540_));
 sg13g2_mux4_1 _8532_ (.S0(net141),
    .A0(\logix.ram_r[832] ),
    .A1(\logix.ram_r[840] ),
    .A2(\logix.ram_r[848] ),
    .A3(\logix.ram_r[856] ),
    .S1(net151),
    .X(_2541_));
 sg13g2_nor2_1 _8533_ (.A(net165),
    .B(_2541_),
    .Y(_2542_));
 sg13g2_buf_8 _8534_ (.A(_2337_),
    .X(_2543_));
 sg13g2_mux2_1 _8535_ (.A0(\logix.ram_r[872] ),
    .A1(\logix.ram_r[888] ),
    .S(net140),
    .X(_2544_));
 sg13g2_nor2_1 _8536_ (.A(net43),
    .B(_2544_),
    .Y(_2545_));
 sg13g2_mux2_1 _8537_ (.A0(\logix.ram_r[864] ),
    .A1(\logix.ram_r[880] ),
    .S(net147),
    .X(_2546_));
 sg13g2_buf_8 _8538_ (.A(_2444_),
    .X(_2547_));
 sg13g2_o21ai_1 _8539_ (.B1(net70),
    .Y(_2548_),
    .A1(net42),
    .A2(_2546_));
 sg13g2_nor3_1 _8540_ (.A(_2542_),
    .B(_2545_),
    .C(_2548_),
    .Y(_2549_));
 sg13g2_o21ai_1 _8541_ (.B1(_2549_),
    .Y(_2550_),
    .A1(net169),
    .A2(_2539_));
 sg13g2_a21oi_2 _8542_ (.B1(_2449_),
    .Y(_2551_),
    .A2(_2212_),
    .A1(_0006_));
 sg13g2_nor2_1 _8543_ (.A(_2551_),
    .B(_2454_),
    .Y(_2552_));
 sg13g2_buf_2 _8544_ (.A(_2552_),
    .X(_2553_));
 sg13g2_buf_8 _8545_ (.A(_2460_),
    .X(_2554_));
 sg13g2_buf_8 _8546_ (.A(_2462_),
    .X(_2555_));
 sg13g2_buf_8 _8547_ (.A(_2416_),
    .X(_2556_));
 sg13g2_mux4_1 _8548_ (.S0(net139),
    .A0(\logix.ram_r[672] ),
    .A1(\logix.ram_r[680] ),
    .A2(\logix.ram_r[688] ),
    .A3(\logix.ram_r[696] ),
    .S1(net138),
    .X(_2557_));
 sg13g2_buf_2 _8549_ (.A(_2426_),
    .X(_2558_));
 sg13g2_mux4_1 _8550_ (.S0(net166),
    .A0(\logix.ram_r[640] ),
    .A1(\logix.ram_r[648] ),
    .A2(\logix.ram_r[656] ),
    .A3(\logix.ram_r[664] ),
    .S1(net137),
    .X(_2559_));
 sg13g2_a22oi_1 _8551_ (.Y(_2560_),
    .B1(_2559_),
    .B2(net40),
    .A2(_2557_),
    .A1(net36));
 sg13g2_buf_1 _8552_ (.A(net158),
    .X(_2561_));
 sg13g2_buf_16 _8553_ (.X(_2562_),
    .A(_2330_));
 sg13g2_buf_8 _8554_ (.A(_2562_),
    .X(_2563_));
 sg13g2_buf_8 _8555_ (.A(_2346_),
    .X(_2564_));
 sg13g2_mux4_1 _8556_ (.S0(net136),
    .A0(\logix.ram_r[736] ),
    .A1(\logix.ram_r[744] ),
    .A2(\logix.ram_r[752] ),
    .A3(\logix.ram_r[760] ),
    .S1(net135),
    .X(_2565_));
 sg13g2_buf_8 _8557_ (.A(_2331_),
    .X(_2566_));
 sg13g2_mux4_1 _8558_ (.S0(_2566_),
    .A0(\logix.ram_r[704] ),
    .A1(\logix.ram_r[712] ),
    .A2(\logix.ram_r[720] ),
    .A3(\logix.ram_r[728] ),
    .S1(net140),
    .X(_2567_));
 sg13g2_buf_2 _8559_ (.A(net154),
    .X(_2568_));
 sg13g2_a22oi_1 _8560_ (.Y(_2569_),
    .B1(_2567_),
    .B2(net68),
    .A2(_2565_),
    .A1(net69));
 sg13g2_buf_1 _8561_ (.A(_2502_),
    .X(_2570_));
 sg13g2_a21oi_1 _8562_ (.A1(_2560_),
    .A2(_2569_),
    .Y(_2571_),
    .B1(net67));
 sg13g2_mux4_1 _8563_ (.S0(net149),
    .A0(\logix.ram_r[544] ),
    .A1(\logix.ram_r[552] ),
    .A2(\logix.ram_r[560] ),
    .A3(\logix.ram_r[568] ),
    .S1(net148),
    .X(_2572_));
 sg13g2_buf_8 _8564_ (.A(_2331_),
    .X(_2573_));
 sg13g2_buf_8 _8565_ (.A(_2426_),
    .X(_2574_));
 sg13g2_mux4_1 _8566_ (.S0(net133),
    .A0(\logix.ram_r[512] ),
    .A1(\logix.ram_r[520] ),
    .A2(\logix.ram_r[528] ),
    .A3(\logix.ram_r[536] ),
    .S1(net132),
    .X(_2575_));
 sg13g2_a22oi_1 _8567_ (.Y(_2576_),
    .B1(_2575_),
    .B2(net40),
    .A2(_2572_),
    .A1(net36));
 sg13g2_buf_8 _8568_ (.A(_2462_),
    .X(_2577_));
 sg13g2_mux4_1 _8569_ (.S0(net131),
    .A0(\logix.ram_r[608] ),
    .A1(\logix.ram_r[616] ),
    .A2(\logix.ram_r[624] ),
    .A3(\logix.ram_r[632] ),
    .S1(net138),
    .X(_2578_));
 sg13g2_buf_8 _8570_ (.A(_2337_),
    .X(_2579_));
 sg13g2_mux4_1 _8571_ (.S0(net166),
    .A0(\logix.ram_r[576] ),
    .A1(\logix.ram_r[584] ),
    .A2(\logix.ram_r[592] ),
    .A3(\logix.ram_r[600] ),
    .S1(net130),
    .X(_2580_));
 sg13g2_a22oi_1 _8572_ (.Y(_2581_),
    .B1(_2580_),
    .B2(net68),
    .A2(_2578_),
    .A1(net76));
 sg13g2_buf_1 _8573_ (.A(_2485_),
    .X(_2582_));
 sg13g2_a21oi_1 _8574_ (.A1(_2576_),
    .A2(_2581_),
    .Y(_2583_),
    .B1(net66));
 sg13g2_nor2_1 _8575_ (.A(_2571_),
    .B(_2583_),
    .Y(_2584_));
 sg13g2_nand4_1 _8576_ (.B(_2550_),
    .C(_2553_),
    .A(_2533_),
    .Y(_2585_),
    .D(_2584_));
 sg13g2_buf_8 _8577_ (.A(net203),
    .X(_2586_));
 sg13g2_buf_8 _8578_ (.A(_2515_),
    .X(_2587_));
 sg13g2_buf_8 _8579_ (.A(net193),
    .X(_2588_));
 sg13g2_mux4_1 _8580_ (.S0(net129),
    .A0(\logix.ram_r[1952] ),
    .A1(\logix.ram_r[1960] ),
    .A2(\logix.ram_r[1968] ),
    .A3(\logix.ram_r[1976] ),
    .S1(net128),
    .X(_2589_));
 sg13g2_buf_8 _8581_ (.A(_2516_),
    .X(_2590_));
 sg13g2_mux4_1 _8582_ (.S0(net172),
    .A0(\logix.ram_r[1920] ),
    .A1(\logix.ram_r[1928] ),
    .A2(\logix.ram_r[1936] ),
    .A3(\logix.ram_r[1944] ),
    .S1(net127),
    .X(_2591_));
 sg13g2_a22oi_1 _8583_ (.Y(_2592_),
    .B1(_2591_),
    .B2(net38),
    .A2(_2589_),
    .A1(net39));
 sg13g2_buf_2 _8584_ (.A(_2431_),
    .X(_2593_));
 sg13g2_buf_1 _8585_ (.A(net126),
    .X(_2594_));
 sg13g2_buf_8 _8586_ (.A(_2527_),
    .X(_2595_));
 sg13g2_buf_8 _8587_ (.A(_2515_),
    .X(_2596_));
 sg13g2_buf_2 _8588_ (.A(net192),
    .X(_2597_));
 sg13g2_mux4_1 _8589_ (.S0(net125),
    .A0(\logix.ram_r[2016] ),
    .A1(\logix.ram_r[2024] ),
    .A2(\logix.ram_r[2032] ),
    .A3(\logix.ram_r[2040] ),
    .S1(net124),
    .X(_2598_));
 sg13g2_mux4_1 _8590_ (.S0(net145),
    .A0(\logix.ram_r[1984] ),
    .A1(\logix.ram_r[1992] ),
    .A2(\logix.ram_r[2000] ),
    .A3(\logix.ram_r[2008] ),
    .S1(net127),
    .X(_2599_));
 sg13g2_a22oi_1 _8591_ (.Y(_2600_),
    .B1(_2599_),
    .B2(net72),
    .A2(_2598_),
    .A1(net65));
 sg13g2_a21oi_1 _8592_ (.A1(_0004_),
    .A2(_2209_),
    .Y(_2601_),
    .B1(_2400_));
 sg13g2_nand2_1 _8593_ (.Y(_2602_),
    .A(_2601_),
    .B(_2442_));
 sg13g2_buf_2 _8594_ (.A(_2602_),
    .X(_2603_));
 sg13g2_a21o_1 _8595_ (.A2(_2600_),
    .A1(_2592_),
    .B1(_2603_),
    .X(_2604_));
 sg13g2_buf_1 _8596_ (.A(_2458_),
    .X(_2605_));
 sg13g2_mux4_1 _8597_ (.S0(net157),
    .A0(\logix.ram_r[1536] ),
    .A1(\logix.ram_r[1544] ),
    .A2(\logix.ram_r[1552] ),
    .A3(\logix.ram_r[1560] ),
    .S1(net156),
    .X(_2606_));
 sg13g2_nand2_1 _8598_ (.Y(_2607_),
    .A(net123),
    .B(_2606_));
 sg13g2_buf_8 _8599_ (.A(_2562_),
    .X(_2608_));
 sg13g2_buf_8 _8600_ (.A(_2346_),
    .X(_2609_));
 sg13g2_mux4_1 _8601_ (.S0(_2608_),
    .A0(\logix.ram_r[1568] ),
    .A1(\logix.ram_r[1576] ),
    .A2(\logix.ram_r[1584] ),
    .A3(\logix.ram_r[1592] ),
    .S1(net121),
    .X(_2610_));
 sg13g2_nand2_1 _8602_ (.Y(_2611_),
    .A(_2507_),
    .B(_2610_));
 sg13g2_buf_1 _8603_ (.A(_2411_),
    .X(_2612_));
 sg13g2_a21oi_1 _8604_ (.A1(_2607_),
    .A2(_2611_),
    .Y(_2613_),
    .B1(net120));
 sg13g2_buf_8 _8605_ (.A(_2389_),
    .X(_2614_));
 sg13g2_buf_8 _8606_ (.A(_2330_),
    .X(_2615_));
 sg13g2_buf_8 _8607_ (.A(net191),
    .X(_2616_));
 sg13g2_mux2_1 _8608_ (.A0(\logix.ram_r[1600] ),
    .A1(\logix.ram_r[1608] ),
    .S(net119),
    .X(_2617_));
 sg13g2_mux2_1 _8609_ (.A0(\logix.ram_r[1648] ),
    .A1(\logix.ram_r[1656] ),
    .S(net129),
    .X(_2618_));
 sg13g2_buf_1 _8610_ (.A(_2395_),
    .X(_2619_));
 sg13g2_a22oi_1 _8611_ (.Y(_2620_),
    .B1(_2618_),
    .B2(net34),
    .A2(_2617_),
    .A1(net35));
 sg13g2_buf_1 _8612_ (.A(_2372_),
    .X(_2621_));
 sg13g2_mux2_1 _8613_ (.A0(\logix.ram_r[1632] ),
    .A1(\logix.ram_r[1640] ),
    .S(net119),
    .X(_2622_));
 sg13g2_mux2_1 _8614_ (.A0(\logix.ram_r[1616] ),
    .A1(\logix.ram_r[1624] ),
    .S(net144),
    .X(_2623_));
 sg13g2_buf_8 _8615_ (.A(_2382_),
    .X(_2624_));
 sg13g2_a22oi_1 _8616_ (.Y(_2625_),
    .B1(_2623_),
    .B2(_2624_),
    .A2(_2622_),
    .A1(_2621_));
 sg13g2_nand2_1 _8617_ (.Y(_2626_),
    .A(_2620_),
    .B(_2625_));
 sg13g2_nor2_1 _8618_ (.A(_2601_),
    .B(_2442_),
    .Y(_2627_));
 sg13g2_o21ai_1 _8619_ (.B1(_2627_),
    .Y(_2628_),
    .A1(_2613_),
    .A2(_2626_));
 sg13g2_buf_8 _8620_ (.A(_2362_),
    .X(_2629_));
 sg13g2_buf_8 _8621_ (.A(_2462_),
    .X(_2630_));
 sg13g2_buf_8 _8622_ (.A(_2337_),
    .X(_2631_));
 sg13g2_mux4_1 _8623_ (.S0(net117),
    .A0(\logix.ram_r[1792] ),
    .A1(\logix.ram_r[1800] ),
    .A2(\logix.ram_r[1808] ),
    .A3(\logix.ram_r[1816] ),
    .S1(net116),
    .X(_2632_));
 sg13g2_nand2_1 _8624_ (.Y(_2633_),
    .A(net123),
    .B(_2632_));
 sg13g2_buf_8 _8625_ (.A(_2462_),
    .X(_2634_));
 sg13g2_mux4_1 _8626_ (.S0(net115),
    .A0(\logix.ram_r[1824] ),
    .A1(\logix.ram_r[1832] ),
    .A2(\logix.ram_r[1840] ),
    .A3(\logix.ram_r[1848] ),
    .S1(net167),
    .X(_2635_));
 sg13g2_nand2_1 _8627_ (.Y(_2636_),
    .A(net179),
    .B(_2635_));
 sg13g2_nand3_1 _8628_ (.B(_2633_),
    .C(_2636_),
    .A(net118),
    .Y(_2637_));
 sg13g2_nor2_1 _8629_ (.A(net191),
    .B(_2380_),
    .Y(_2638_));
 sg13g2_buf_4 _8630_ (.X(_2639_),
    .A(_2638_));
 sg13g2_buf_8 _8631_ (.A(_2346_),
    .X(_2640_));
 sg13g2_buf_8 _8632_ (.A(net114),
    .X(_2641_));
 sg13g2_buf_8 _8633_ (.A(_2336_),
    .X(_2642_));
 sg13g2_buf_8 _8634_ (.A(net190),
    .X(_2643_));
 sg13g2_nand2b_1 _8635_ (.Y(_2644_),
    .B(net113),
    .A_N(\logix.ram_r[1872] ));
 sg13g2_o21ai_1 _8636_ (.B1(_2644_),
    .Y(_2645_),
    .A1(\logix.ram_r[1856] ),
    .A2(net64));
 sg13g2_nor2_1 _8637_ (.A(_2342_),
    .B(net202),
    .Y(_2646_));
 sg13g2_buf_8 _8638_ (.A(_2646_),
    .X(_2647_));
 sg13g2_buf_8 _8639_ (.A(_2337_),
    .X(_2648_));
 sg13g2_buf_8 _8640_ (.A(net112),
    .X(_2649_));
 sg13g2_buf_8 _8641_ (.A(net190),
    .X(_2650_));
 sg13g2_nand2b_1 _8642_ (.Y(_2651_),
    .B(net111),
    .A_N(\logix.ram_r[1880] ));
 sg13g2_o21ai_1 _8643_ (.B1(_2651_),
    .Y(_2652_),
    .A1(\logix.ram_r[1864] ),
    .A2(net63));
 sg13g2_a22oi_1 _8644_ (.Y(_2653_),
    .B1(_2647_),
    .B2(_2652_),
    .A2(_2645_),
    .A1(_2639_));
 sg13g2_buf_2 _8645_ (.A(net193),
    .X(_2654_));
 sg13g2_mux4_1 _8646_ (.S0(net171),
    .A0(\logix.ram_r[1888] ),
    .A1(\logix.ram_r[1896] ),
    .A2(\logix.ram_r[1904] ),
    .A3(\logix.ram_r[1912] ),
    .S1(net110),
    .X(_2655_));
 sg13g2_nand2b_1 _8647_ (.Y(_2656_),
    .B(net65),
    .A_N(_2655_));
 sg13g2_nand4_1 _8648_ (.B(_2637_),
    .C(_2653_),
    .A(net79),
    .Y(_2657_),
    .D(_2656_));
 sg13g2_buf_8 _8649_ (.A(net78),
    .X(_2658_));
 sg13g2_mux4_1 _8650_ (.S0(net122),
    .A0(\logix.ram_r[1696] ),
    .A1(\logix.ram_r[1704] ),
    .A2(\logix.ram_r[1712] ),
    .A3(\logix.ram_r[1720] ),
    .S1(net121),
    .X(_2659_));
 sg13g2_mux4_1 _8651_ (.S0(net134),
    .A0(\logix.ram_r[1664] ),
    .A1(\logix.ram_r[1672] ),
    .A2(\logix.ram_r[1680] ),
    .A3(\logix.ram_r[1688] ),
    .S1(net177),
    .X(_2660_));
 sg13g2_buf_8 _8652_ (.A(net77),
    .X(_2661_));
 sg13g2_a22oi_1 _8653_ (.Y(_2662_),
    .B1(_2660_),
    .B2(net30),
    .A2(_2659_),
    .A1(net31));
 sg13g2_buf_1 _8654_ (.A(net158),
    .X(_2663_));
 sg13g2_buf_8 _8655_ (.A(_2562_),
    .X(_2664_));
 sg13g2_mux4_1 _8656_ (.S0(net109),
    .A0(\logix.ram_r[1760] ),
    .A1(\logix.ram_r[1768] ),
    .A2(\logix.ram_r[1776] ),
    .A3(\logix.ram_r[1784] ),
    .S1(net147),
    .X(_2665_));
 sg13g2_mux4_1 _8657_ (.S0(net149),
    .A0(\logix.ram_r[1728] ),
    .A1(\logix.ram_r[1736] ),
    .A2(\logix.ram_r[1744] ),
    .A3(\logix.ram_r[1752] ),
    .S1(net167),
    .X(_2666_));
 sg13g2_buf_2 _8658_ (.A(net154),
    .X(_2667_));
 sg13g2_a22oi_1 _8659_ (.Y(_2668_),
    .B1(_2666_),
    .B2(net61),
    .A2(_2665_),
    .A1(net62));
 sg13g2_a21oi_1 _8660_ (.A1(_2662_),
    .A2(_2668_),
    .Y(_2669_),
    .B1(net67));
 sg13g2_or2_1 _8661_ (.X(_2670_),
    .B(_2454_),
    .A(_2451_));
 sg13g2_nor2_1 _8662_ (.A(_2669_),
    .B(_2670_),
    .Y(_2671_));
 sg13g2_nand4_1 _8663_ (.B(_2628_),
    .C(_2657_),
    .A(_2604_),
    .Y(_2672_),
    .D(_2671_));
 sg13g2_mux4_1 _8664_ (.S0(net160),
    .A0(\logix.ram_r[1408] ),
    .A1(\logix.ram_r[1416] ),
    .A2(\logix.ram_r[1424] ),
    .A3(\logix.ram_r[1432] ),
    .S1(net163),
    .X(_2673_));
 sg13g2_nand2_1 _8665_ (.Y(_2674_),
    .A(net123),
    .B(_2673_));
 sg13g2_mux4_1 _8666_ (.S0(net141),
    .A0(\logix.ram_r[1440] ),
    .A1(\logix.ram_r[1448] ),
    .A2(\logix.ram_r[1456] ),
    .A3(\logix.ram_r[1464] ),
    .S1(net151),
    .X(_2675_));
 sg13g2_nand2_1 _8667_ (.Y(_2676_),
    .A(net179),
    .B(_2675_));
 sg13g2_nand3_1 _8668_ (.B(_2674_),
    .C(_2676_),
    .A(_2629_),
    .Y(_2677_));
 sg13g2_buf_8 _8669_ (.A(_2639_),
    .X(_2678_));
 sg13g2_nand2b_1 _8670_ (.Y(_2679_),
    .B(net124),
    .A_N(\logix.ram_r[1488] ));
 sg13g2_o21ai_1 _8671_ (.B1(_2679_),
    .Y(_2680_),
    .A1(\logix.ram_r[1472] ),
    .A2(net63));
 sg13g2_buf_8 _8672_ (.A(net151),
    .X(_2681_));
 sg13g2_nand2b_1 _8673_ (.Y(_2682_),
    .B(net110),
    .A_N(\logix.ram_r[1496] ));
 sg13g2_o21ai_1 _8674_ (.B1(_2682_),
    .Y(_2683_),
    .A1(\logix.ram_r[1480] ),
    .A2(net60));
 sg13g2_buf_1 _8675_ (.A(_2647_),
    .X(_2684_));
 sg13g2_a22oi_1 _8676_ (.Y(_2685_),
    .B1(_2683_),
    .B2(net28),
    .A2(_2680_),
    .A1(net29));
 sg13g2_buf_8 _8677_ (.A(_2354_),
    .X(_2686_));
 sg13g2_buf_8 _8678_ (.A(net108),
    .X(_2687_));
 sg13g2_mux4_1 _8679_ (.S0(_2385_),
    .A0(\logix.ram_r[1504] ),
    .A1(\logix.ram_r[1512] ),
    .A2(\logix.ram_r[1520] ),
    .A3(\logix.ram_r[1528] ),
    .S1(_2687_),
    .X(_2688_));
 sg13g2_nand2b_1 _8680_ (.Y(_2689_),
    .B(net65),
    .A_N(_2688_));
 sg13g2_nand4_1 _8681_ (.B(_2677_),
    .C(_2685_),
    .A(_2408_),
    .Y(_2690_),
    .D(_2689_));
 sg13g2_mux4_1 _8682_ (.S0(net178),
    .A0(\logix.ram_r[1280] ),
    .A1(\logix.ram_r[1288] ),
    .A2(\logix.ram_r[1296] ),
    .A3(\logix.ram_r[1304] ),
    .S1(net177),
    .X(_2691_));
 sg13g2_nand2_1 _8683_ (.Y(_2692_),
    .A(net123),
    .B(_2691_));
 sg13g2_mux4_1 _8684_ (.S0(net117),
    .A0(\logix.ram_r[1312] ),
    .A1(\logix.ram_r[1320] ),
    .A2(\logix.ram_r[1328] ),
    .A3(\logix.ram_r[1336] ),
    .S1(net116),
    .X(_2693_));
 sg13g2_nand2_1 _8685_ (.Y(_2694_),
    .A(net179),
    .B(_2693_));
 sg13g2_a21oi_1 _8686_ (.A1(_2692_),
    .A2(_2694_),
    .Y(_2695_),
    .B1(net120));
 sg13g2_buf_8 _8687_ (.A(_2389_),
    .X(_2696_));
 sg13g2_mux2_1 _8688_ (.A0(\logix.ram_r[1344] ),
    .A1(\logix.ram_r[1352] ),
    .S(net119),
    .X(_2697_));
 sg13g2_mux2_1 _8689_ (.A0(\logix.ram_r[1376] ),
    .A1(\logix.ram_r[1384] ),
    .S(net125),
    .X(_2698_));
 sg13g2_a22oi_1 _8690_ (.Y(_2699_),
    .B1(_2698_),
    .B2(net48),
    .A2(_2697_),
    .A1(net27));
 sg13g2_buf_8 _8691_ (.A(_2395_),
    .X(_2700_));
 sg13g2_mux2_1 _8692_ (.A0(\logix.ram_r[1392] ),
    .A1(\logix.ram_r[1400] ),
    .S(net164),
    .X(_2701_));
 sg13g2_buf_8 _8693_ (.A(_2615_),
    .X(_2702_));
 sg13g2_mux2_1 _8694_ (.A0(\logix.ram_r[1360] ),
    .A1(\logix.ram_r[1368] ),
    .S(net107),
    .X(_2703_));
 sg13g2_a22oi_1 _8695_ (.Y(_2704_),
    .B1(_2703_),
    .B2(net32),
    .A2(_2701_),
    .A1(net26));
 sg13g2_nand2_2 _8696_ (.Y(_2705_),
    .A(_2551_),
    .B(_2454_));
 sg13g2_inv_4 _8697_ (.A(_2705_),
    .Y(_2706_));
 sg13g2_nand3_1 _8698_ (.B(_2704_),
    .C(_2706_),
    .A(_2699_),
    .Y(_2707_));
 sg13g2_nand2_1 _8699_ (.Y(_2708_),
    .A(_2601_),
    .B(_2405_));
 sg13g2_buf_1 _8700_ (.A(_2708_),
    .X(_2709_));
 sg13g2_nand2_2 _8701_ (.Y(_2710_),
    .A(_2709_),
    .B(_2706_));
 sg13g2_o21ai_1 _8702_ (.B1(_2710_),
    .Y(_2711_),
    .A1(_2695_),
    .A2(_2707_));
 sg13g2_buf_8 _8703_ (.A(_2331_),
    .X(_2712_));
 sg13g2_mux4_1 _8704_ (.S0(_2712_),
    .A0(\logix.ram_r[1184] ),
    .A1(\logix.ram_r[1192] ),
    .A2(\logix.ram_r[1200] ),
    .A3(\logix.ram_r[1208] ),
    .S1(net140),
    .X(_2713_));
 sg13g2_mux4_1 _8705_ (.S0(net141),
    .A0(\logix.ram_r[1152] ),
    .A1(\logix.ram_r[1160] ),
    .A2(\logix.ram_r[1168] ),
    .A3(\logix.ram_r[1176] ),
    .S1(net151),
    .X(_2714_));
 sg13g2_buf_8 _8706_ (.A(net77),
    .X(_2715_));
 sg13g2_a22oi_1 _8707_ (.Y(_2716_),
    .B1(_2714_),
    .B2(net25),
    .A2(_2713_),
    .A1(net41));
 sg13g2_mux4_1 _8708_ (.S0(net149),
    .A0(\logix.ram_r[1248] ),
    .A1(\logix.ram_r[1256] ),
    .A2(\logix.ram_r[1264] ),
    .A3(\logix.ram_r[1272] ),
    .S1(net167),
    .X(_2717_));
 sg13g2_mux4_1 _8709_ (.S0(net155),
    .A0(\logix.ram_r[1216] ),
    .A1(\logix.ram_r[1224] ),
    .A2(\logix.ram_r[1232] ),
    .A3(\logix.ram_r[1240] ),
    .S1(net162),
    .X(_2718_));
 sg13g2_a22oi_1 _8710_ (.Y(_2719_),
    .B1(_2718_),
    .B2(net75),
    .A2(_2717_),
    .A1(net76));
 sg13g2_a21oi_1 _8711_ (.A1(_2716_),
    .A2(_2719_),
    .Y(_2720_),
    .B1(net71));
 sg13g2_buf_8 _8712_ (.A(_2331_),
    .X(_2721_));
 sg13g2_mux4_1 _8713_ (.S0(net105),
    .A0(\logix.ram_r[1056] ),
    .A1(\logix.ram_r[1064] ),
    .A2(\logix.ram_r[1072] ),
    .A3(\logix.ram_r[1080] ),
    .S1(net130),
    .X(_2722_));
 sg13g2_mux4_1 _8714_ (.S0(_2425_),
    .A0(\logix.ram_r[1024] ),
    .A1(\logix.ram_r[1032] ),
    .A2(\logix.ram_r[1040] ),
    .A3(\logix.ram_r[1048] ),
    .S1(_2427_),
    .X(_2723_));
 sg13g2_a22oi_1 _8715_ (.Y(_2724_),
    .B1(_2723_),
    .B2(net38),
    .A2(_2722_),
    .A1(net39));
 sg13g2_mux4_1 _8716_ (.S0(net106),
    .A0(\logix.ram_r[1120] ),
    .A1(\logix.ram_r[1128] ),
    .A2(\logix.ram_r[1136] ),
    .A3(\logix.ram_r[1144] ),
    .S1(_2648_),
    .X(_2725_));
 sg13g2_mux4_1 _8717_ (.S0(net141),
    .A0(\logix.ram_r[1088] ),
    .A1(\logix.ram_r[1096] ),
    .A2(\logix.ram_r[1104] ),
    .A3(\logix.ram_r[1112] ),
    .S1(net151),
    .X(_2726_));
 sg13g2_a22oi_1 _8718_ (.Y(_2727_),
    .B1(_2726_),
    .B2(net72),
    .A2(_2725_),
    .A1(net73));
 sg13g2_a21oi_1 _8719_ (.A1(_2724_),
    .A2(_2727_),
    .Y(_2728_),
    .B1(net74));
 sg13g2_nor2_1 _8720_ (.A(_2720_),
    .B(_2728_),
    .Y(_2729_));
 sg13g2_nand3_1 _8721_ (.B(_2711_),
    .C(_2729_),
    .A(_2690_),
    .Y(_2730_));
 sg13g2_and4_1 _8722_ (.A(_2506_),
    .B(_2585_),
    .C(_2672_),
    .D(_2730_),
    .X(net14));
 sg13g2_mux4_1 _8723_ (.S0(net115),
    .A0(\logix.ram_r[897] ),
    .A1(\logix.ram_r[905] ),
    .A2(\logix.ram_r[913] ),
    .A3(\logix.ram_r[921] ),
    .S1(net167),
    .X(_2731_));
 sg13g2_nor2_1 _8724_ (.A(net150),
    .B(_2731_),
    .Y(_2732_));
 sg13g2_buf_8 _8725_ (.A(_2354_),
    .X(_2733_));
 sg13g2_mux2_1 _8726_ (.A0(\logix.ram_r[929] ),
    .A1(\logix.ram_r[945] ),
    .S(net104),
    .X(_2734_));
 sg13g2_nor2_1 _8727_ (.A(net83),
    .B(_2734_),
    .Y(_2735_));
 sg13g2_buf_2 _8728_ (.A(_2515_),
    .X(_2736_));
 sg13g2_mux2_1 _8729_ (.A0(\logix.ram_r[937] ),
    .A1(\logix.ram_r[953] ),
    .S(net189),
    .X(_2737_));
 sg13g2_o21ai_1 _8730_ (.B1(net174),
    .Y(_2738_),
    .A1(net82),
    .A2(_2737_));
 sg13g2_nor3_1 _8731_ (.A(_2732_),
    .B(_2735_),
    .C(_2738_),
    .Y(_2739_));
 sg13g2_mux2_1 _8732_ (.A0(\logix.ram_r[993] ),
    .A1(\logix.ram_r[1001] ),
    .S(_2595_),
    .X(_2740_));
 sg13g2_mux2_1 _8733_ (.A0(\logix.ram_r[977] ),
    .A1(\logix.ram_r[985] ),
    .S(net145),
    .X(_2741_));
 sg13g2_buf_8 _8734_ (.A(_2382_),
    .X(_2742_));
 sg13g2_a22oi_1 _8735_ (.Y(_2743_),
    .B1(_2741_),
    .B2(net24),
    .A2(_2740_),
    .A1(net37));
 sg13g2_buf_8 _8736_ (.A(net195),
    .X(_2744_));
 sg13g2_mux2_1 _8737_ (.A0(\logix.ram_r[961] ),
    .A1(\logix.ram_r[969] ),
    .S(net103),
    .X(_2745_));
 sg13g2_mux2_1 _8738_ (.A0(\logix.ram_r[1009] ),
    .A1(\logix.ram_r[1017] ),
    .S(net173),
    .X(_2746_));
 sg13g2_a22oi_1 _8739_ (.Y(_2747_),
    .B1(_2746_),
    .B2(net34),
    .A2(_2745_),
    .A1(net35));
 sg13g2_nand2_1 _8740_ (.Y(_2748_),
    .A(_2743_),
    .B(_2747_));
 sg13g2_o21ai_1 _8741_ (.B1(net81),
    .Y(_2749_),
    .A1(_2739_),
    .A2(_2748_));
 sg13g2_buf_8 _8742_ (.A(_2416_),
    .X(_2750_));
 sg13g2_mux4_1 _8743_ (.S0(_2750_),
    .A0(\logix.ram_r[769] ),
    .A1(\logix.ram_r[785] ),
    .A2(\logix.ram_r[801] ),
    .A3(\logix.ram_r[817] ),
    .S1(net199),
    .X(_2751_));
 sg13g2_mux4_1 _8744_ (.S0(_2534_),
    .A0(\logix.ram_r[777] ),
    .A1(\logix.ram_r[793] ),
    .A2(\logix.ram_r[809] ),
    .A3(\logix.ram_r[825] ),
    .S1(net194),
    .X(_2752_));
 sg13g2_mux2_1 _8745_ (.A0(_2751_),
    .A1(_2752_),
    .S(net44),
    .X(_2753_));
 sg13g2_mux4_1 _8746_ (.S0(net141),
    .A0(\logix.ram_r[833] ),
    .A1(\logix.ram_r[841] ),
    .A2(\logix.ram_r[849] ),
    .A3(\logix.ram_r[857] ),
    .S1(_2469_),
    .X(_2754_));
 sg13g2_nor2_1 _8747_ (.A(net165),
    .B(_2754_),
    .Y(_2755_));
 sg13g2_mux2_1 _8748_ (.A0(\logix.ram_r[873] ),
    .A1(\logix.ram_r[889] ),
    .S(net177),
    .X(_2756_));
 sg13g2_nor2_1 _8749_ (.A(net43),
    .B(_2756_),
    .Y(_2757_));
 sg13g2_buf_8 _8750_ (.A(_2346_),
    .X(_2758_));
 sg13g2_mux2_1 _8751_ (.A0(\logix.ram_r[865] ),
    .A1(\logix.ram_r[881] ),
    .S(net101),
    .X(_2759_));
 sg13g2_o21ai_1 _8752_ (.B1(net70),
    .Y(_2760_),
    .A1(net42),
    .A2(_2759_));
 sg13g2_nor3_1 _8753_ (.A(_2755_),
    .B(_2757_),
    .C(_2760_),
    .Y(_2761_));
 sg13g2_o21ai_1 _8754_ (.B1(_2761_),
    .Y(_2762_),
    .A1(net169),
    .A2(_2753_));
 sg13g2_mux4_1 _8755_ (.S0(net161),
    .A0(\logix.ram_r[673] ),
    .A1(\logix.ram_r[681] ),
    .A2(\logix.ram_r[689] ),
    .A3(\logix.ram_r[697] ),
    .S1(net168),
    .X(_2763_));
 sg13g2_mux4_1 _8756_ (.S0(net152),
    .A0(\logix.ram_r[641] ),
    .A1(\logix.ram_r[649] ),
    .A2(\logix.ram_r[657] ),
    .A3(\logix.ram_r[665] ),
    .S1(_2497_),
    .X(_2764_));
 sg13g2_a22oi_1 _8757_ (.Y(_2765_),
    .B1(_2764_),
    .B2(_2715_),
    .A2(_2763_),
    .A1(net41));
 sg13g2_mux4_1 _8758_ (.S0(_2555_),
    .A0(\logix.ram_r[737] ),
    .A1(\logix.ram_r[745] ),
    .A2(\logix.ram_r[753] ),
    .A3(\logix.ram_r[761] ),
    .S1(net156),
    .X(_2766_));
 sg13g2_mux4_1 _8759_ (.S0(net155),
    .A0(\logix.ram_r[705] ),
    .A1(\logix.ram_r[713] ),
    .A2(\logix.ram_r[721] ),
    .A3(\logix.ram_r[729] ),
    .S1(net162),
    .X(_2767_));
 sg13g2_a22oi_1 _8760_ (.Y(_2768_),
    .B1(_2767_),
    .B2(net75),
    .A2(_2766_),
    .A1(net76));
 sg13g2_a21oi_1 _8761_ (.A1(_2765_),
    .A2(_2768_),
    .Y(_2769_),
    .B1(_2503_));
 sg13g2_mux4_1 _8762_ (.S0(net178),
    .A0(\logix.ram_r[545] ),
    .A1(\logix.ram_r[553] ),
    .A2(\logix.ram_r[561] ),
    .A3(\logix.ram_r[569] ),
    .S1(net153),
    .X(_2770_));
 sg13g2_mux4_1 _8763_ (.S0(net160),
    .A0(\logix.ram_r[513] ),
    .A1(\logix.ram_r[521] ),
    .A2(\logix.ram_r[529] ),
    .A3(\logix.ram_r[537] ),
    .S1(net163),
    .X(_2771_));
 sg13g2_a22oi_1 _8764_ (.Y(_2772_),
    .B1(_2771_),
    .B2(net25),
    .A2(_2770_),
    .A1(net41));
 sg13g2_mux4_1 _8765_ (.S0(net117),
    .A0(\logix.ram_r[609] ),
    .A1(\logix.ram_r[617] ),
    .A2(\logix.ram_r[625] ),
    .A3(\logix.ram_r[633] ),
    .S1(net168),
    .X(_2773_));
 sg13g2_mux4_1 _8766_ (.S0(net152),
    .A0(\logix.ram_r[577] ),
    .A1(\logix.ram_r[585] ),
    .A2(\logix.ram_r[593] ),
    .A3(\logix.ram_r[601] ),
    .S1(net132),
    .X(_2774_));
 sg13g2_a22oi_1 _8767_ (.Y(_2775_),
    .B1(_2774_),
    .B2(net75),
    .A2(_2773_),
    .A1(net73));
 sg13g2_a21oi_1 _8768_ (.A1(_2772_),
    .A2(_2775_),
    .Y(_2776_),
    .B1(net74));
 sg13g2_nor2_1 _8769_ (.A(_2769_),
    .B(_2776_),
    .Y(_2777_));
 sg13g2_nand4_1 _8770_ (.B(_2749_),
    .C(_2762_),
    .A(_2553_),
    .Y(_2778_),
    .D(_2777_));
 sg13g2_nor2_1 _8771_ (.A(_2451_),
    .B(_2454_),
    .Y(_2779_));
 sg13g2_buf_2 _8772_ (.A(_2779_),
    .X(_2780_));
 sg13g2_buf_1 _8773_ (.A(_2325_),
    .X(_2781_));
 sg13g2_buf_8 _8774_ (.A(_2562_),
    .X(_2782_));
 sg13g2_mux4_1 _8775_ (.S0(net100),
    .A0(\logix.ram_r[1921] ),
    .A1(\logix.ram_r[1929] ),
    .A2(\logix.ram_r[1937] ),
    .A3(\logix.ram_r[1945] ),
    .S1(net176),
    .X(_2783_));
 sg13g2_nor2_1 _8776_ (.A(net188),
    .B(_2783_),
    .Y(_2784_));
 sg13g2_buf_8 _8777_ (.A(_2354_),
    .X(_2785_));
 sg13g2_mux2_1 _8778_ (.A0(\logix.ram_r[1953] ),
    .A1(\logix.ram_r[1969] ),
    .S(net99),
    .X(_2786_));
 sg13g2_nor2_1 _8779_ (.A(net83),
    .B(_2786_),
    .Y(_2787_));
 sg13g2_mux2_1 _8780_ (.A0(\logix.ram_r[1961] ),
    .A1(\logix.ram_r[1977] ),
    .S(net193),
    .X(_2788_));
 sg13g2_buf_1 _8781_ (.A(_2362_),
    .X(_2789_));
 sg13g2_o21ai_1 _8782_ (.B1(net98),
    .Y(_2790_),
    .A1(net82),
    .A2(_2788_));
 sg13g2_nor3_1 _8783_ (.A(_2784_),
    .B(_2787_),
    .C(_2790_),
    .Y(_2791_));
 sg13g2_mux2_1 _8784_ (.A0(\logix.ram_r[2017] ),
    .A1(\logix.ram_r[2025] ),
    .S(net103),
    .X(_2792_));
 sg13g2_mux2_1 _8785_ (.A0(\logix.ram_r[2001] ),
    .A1(\logix.ram_r[2009] ),
    .S(net171),
    .X(_2793_));
 sg13g2_a22oi_1 _8786_ (.Y(_2794_),
    .B1(_2793_),
    .B2(net24),
    .A2(_2792_),
    .A1(net37));
 sg13g2_mux2_1 _8787_ (.A0(\logix.ram_r[1985] ),
    .A1(\logix.ram_r[1993] ),
    .S(net107),
    .X(_2795_));
 sg13g2_mux2_1 _8788_ (.A0(\logix.ram_r[2033] ),
    .A1(\logix.ram_r[2041] ),
    .S(net129),
    .X(_2796_));
 sg13g2_a22oi_1 _8789_ (.Y(_2797_),
    .B1(_2796_),
    .B2(net34),
    .A2(_2795_),
    .A1(net35));
 sg13g2_nand2_1 _8790_ (.Y(_2798_),
    .A(_2794_),
    .B(_2797_));
 sg13g2_o21ai_1 _8791_ (.B1(net81),
    .Y(_2799_),
    .A1(_2791_),
    .A2(_2798_));
 sg13g2_buf_1 _8792_ (.A(_2325_),
    .X(_2800_));
 sg13g2_mux4_1 _8793_ (.S0(net121),
    .A0(\logix.ram_r[1793] ),
    .A1(\logix.ram_r[1809] ),
    .A2(\logix.ram_r[1825] ),
    .A3(\logix.ram_r[1841] ),
    .S1(net187),
    .X(_2801_));
 sg13g2_mux4_1 _8794_ (.S0(net135),
    .A0(\logix.ram_r[1801] ),
    .A1(\logix.ram_r[1817] ),
    .A2(\logix.ram_r[1833] ),
    .A3(\logix.ram_r[1849] ),
    .S1(net187),
    .X(_2802_));
 sg13g2_mux2_1 _8795_ (.A0(_2801_),
    .A1(_2802_),
    .S(net44),
    .X(_2803_));
 sg13g2_mux4_1 _8796_ (.S0(net133),
    .A0(\logix.ram_r[1857] ),
    .A1(\logix.ram_r[1865] ),
    .A2(\logix.ram_r[1873] ),
    .A3(\logix.ram_r[1881] ),
    .S1(net162),
    .X(_2804_));
 sg13g2_nor2_1 _8797_ (.A(net165),
    .B(_2804_),
    .Y(_2805_));
 sg13g2_mux2_1 _8798_ (.A0(\logix.ram_r[1897] ),
    .A1(\logix.ram_r[1913] ),
    .S(net148),
    .X(_2806_));
 sg13g2_nor2_1 _8799_ (.A(net43),
    .B(_2806_),
    .Y(_2807_));
 sg13g2_buf_8 _8800_ (.A(_2354_),
    .X(_2808_));
 sg13g2_mux2_1 _8801_ (.A0(\logix.ram_r[1889] ),
    .A1(\logix.ram_r[1905] ),
    .S(net97),
    .X(_2809_));
 sg13g2_o21ai_1 _8802_ (.B1(net70),
    .Y(_2810_),
    .A1(net42),
    .A2(_2809_));
 sg13g2_nor3_1 _8803_ (.A(_2805_),
    .B(_2807_),
    .C(_2810_),
    .Y(_2811_));
 sg13g2_o21ai_1 _8804_ (.B1(_2811_),
    .Y(_2812_),
    .A1(net169),
    .A2(_2803_));
 sg13g2_mux4_1 _8805_ (.S0(net131),
    .A0(\logix.ram_r[1697] ),
    .A1(\logix.ram_r[1705] ),
    .A2(\logix.ram_r[1713] ),
    .A3(\logix.ram_r[1721] ),
    .S1(net138),
    .X(_2813_));
 sg13g2_mux4_1 _8806_ (.S0(net166),
    .A0(\logix.ram_r[1665] ),
    .A1(\logix.ram_r[1673] ),
    .A2(\logix.ram_r[1681] ),
    .A3(\logix.ram_r[1689] ),
    .S1(net137),
    .X(_2814_));
 sg13g2_a22oi_1 _8807_ (.Y(_2815_),
    .B1(_2814_),
    .B2(net30),
    .A2(_2813_),
    .A1(net31));
 sg13g2_mux4_1 _8808_ (.S0(net136),
    .A0(\logix.ram_r[1761] ),
    .A1(\logix.ram_r[1769] ),
    .A2(\logix.ram_r[1777] ),
    .A3(\logix.ram_r[1785] ),
    .S1(net135),
    .X(_2816_));
 sg13g2_mux4_1 _8809_ (.S0(net134),
    .A0(\logix.ram_r[1729] ),
    .A1(\logix.ram_r[1737] ),
    .A2(\logix.ram_r[1745] ),
    .A3(\logix.ram_r[1753] ),
    .S1(net140),
    .X(_2817_));
 sg13g2_a22oi_1 _8810_ (.Y(_2818_),
    .B1(_2817_),
    .B2(net61),
    .A2(_2816_),
    .A1(net69));
 sg13g2_a21oi_1 _8811_ (.A1(_2815_),
    .A2(_2818_),
    .Y(_2819_),
    .B1(net67));
 sg13g2_mux4_1 _8812_ (.S0(net149),
    .A0(\logix.ram_r[1569] ),
    .A1(\logix.ram_r[1577] ),
    .A2(\logix.ram_r[1585] ),
    .A3(\logix.ram_r[1593] ),
    .S1(net148),
    .X(_2820_));
 sg13g2_mux4_1 _8813_ (.S0(net133),
    .A0(\logix.ram_r[1537] ),
    .A1(\logix.ram_r[1545] ),
    .A2(\logix.ram_r[1553] ),
    .A3(\logix.ram_r[1561] ),
    .S1(net132),
    .X(_2821_));
 sg13g2_a22oi_1 _8814_ (.Y(_2822_),
    .B1(_2821_),
    .B2(net40),
    .A2(_2820_),
    .A1(net36));
 sg13g2_mux4_1 _8815_ (.S0(net131),
    .A0(\logix.ram_r[1633] ),
    .A1(\logix.ram_r[1641] ),
    .A2(\logix.ram_r[1649] ),
    .A3(\logix.ram_r[1657] ),
    .S1(net138),
    .X(_2823_));
 sg13g2_mux4_1 _8816_ (.S0(net105),
    .A0(\logix.ram_r[1601] ),
    .A1(\logix.ram_r[1609] ),
    .A2(\logix.ram_r[1617] ),
    .A3(\logix.ram_r[1625] ),
    .S1(net130),
    .X(_2824_));
 sg13g2_a22oi_1 _8817_ (.Y(_2825_),
    .B1(_2824_),
    .B2(net68),
    .A2(_2823_),
    .A1(net76));
 sg13g2_a21oi_1 _8818_ (.A1(_2822_),
    .A2(_2825_),
    .Y(_2826_),
    .B1(net66));
 sg13g2_nor2_1 _8819_ (.A(_2819_),
    .B(_2826_),
    .Y(_2827_));
 sg13g2_nand4_1 _8820_ (.B(_2799_),
    .C(_2812_),
    .A(_2780_),
    .Y(_2828_),
    .D(_2827_));
 sg13g2_mux4_1 _8821_ (.S0(net160),
    .A0(\logix.ram_r[1409] ),
    .A1(\logix.ram_r[1417] ),
    .A2(\logix.ram_r[1425] ),
    .A3(\logix.ram_r[1433] ),
    .S1(net163),
    .X(_2829_));
 sg13g2_nand2_1 _8822_ (.Y(_2830_),
    .A(net123),
    .B(_2829_));
 sg13g2_mux4_1 _8823_ (.S0(net160),
    .A0(\logix.ram_r[1441] ),
    .A1(\logix.ram_r[1449] ),
    .A2(\logix.ram_r[1457] ),
    .A3(\logix.ram_r[1465] ),
    .S1(net163),
    .X(_2831_));
 sg13g2_nand2_1 _8824_ (.Y(_2832_),
    .A(net179),
    .B(_2831_));
 sg13g2_nand3_1 _8825_ (.B(_2830_),
    .C(_2832_),
    .A(_2629_),
    .Y(_2833_));
 sg13g2_nand2b_1 _8826_ (.Y(_2834_),
    .B(net124),
    .A_N(\logix.ram_r[1489] ));
 sg13g2_o21ai_1 _8827_ (.B1(_2834_),
    .Y(_2835_),
    .A1(\logix.ram_r[1473] ),
    .A2(net63));
 sg13g2_nand2b_1 _8828_ (.Y(_2836_),
    .B(net110),
    .A_N(\logix.ram_r[1497] ));
 sg13g2_o21ai_1 _8829_ (.B1(_2836_),
    .Y(_2837_),
    .A1(\logix.ram_r[1481] ),
    .A2(net60));
 sg13g2_a22oi_1 _8830_ (.Y(_2838_),
    .B1(_2837_),
    .B2(net28),
    .A2(_2835_),
    .A1(net29));
 sg13g2_mux4_1 _8831_ (.S0(_2385_),
    .A0(\logix.ram_r[1505] ),
    .A1(\logix.ram_r[1513] ),
    .A2(\logix.ram_r[1521] ),
    .A3(\logix.ram_r[1529] ),
    .S1(net59),
    .X(_2839_));
 sg13g2_nand2b_1 _8832_ (.Y(_2840_),
    .B(net65),
    .A_N(_2839_));
 sg13g2_nand4_1 _8833_ (.B(_2833_),
    .C(_2838_),
    .A(net81),
    .Y(_2841_),
    .D(_2840_));
 sg13g2_mux4_1 _8834_ (.S0(net105),
    .A0(\logix.ram_r[1281] ),
    .A1(\logix.ram_r[1289] ),
    .A2(\logix.ram_r[1297] ),
    .A3(\logix.ram_r[1305] ),
    .S1(net130),
    .X(_2842_));
 sg13g2_nand2_1 _8835_ (.Y(_2843_),
    .A(net123),
    .B(_2842_));
 sg13g2_mux4_1 _8836_ (.S0(net106),
    .A0(\logix.ram_r[1313] ),
    .A1(\logix.ram_r[1321] ),
    .A2(\logix.ram_r[1329] ),
    .A3(\logix.ram_r[1337] ),
    .S1(net112),
    .X(_2844_));
 sg13g2_nand2_1 _8837_ (.Y(_2845_),
    .A(net179),
    .B(_2844_));
 sg13g2_a21oi_1 _8838_ (.A1(_2843_),
    .A2(_2845_),
    .Y(_2846_),
    .B1(net120));
 sg13g2_buf_8 _8839_ (.A(net191),
    .X(_2847_));
 sg13g2_mux2_1 _8840_ (.A0(\logix.ram_r[1345] ),
    .A1(\logix.ram_r[1353] ),
    .S(net96),
    .X(_2848_));
 sg13g2_mux2_1 _8841_ (.A0(\logix.ram_r[1377] ),
    .A1(\logix.ram_r[1385] ),
    .S(net103),
    .X(_2849_));
 sg13g2_a22oi_1 _8842_ (.Y(_2850_),
    .B1(_2849_),
    .B2(net37),
    .A2(_2848_),
    .A1(net27));
 sg13g2_mux2_1 _8843_ (.A0(\logix.ram_r[1393] ),
    .A1(\logix.ram_r[1401] ),
    .S(net164),
    .X(_2851_));
 sg13g2_mux2_1 _8844_ (.A0(\logix.ram_r[1361] ),
    .A1(\logix.ram_r[1369] ),
    .S(net107),
    .X(_2852_));
 sg13g2_a22oi_1 _8845_ (.Y(_2853_),
    .B1(_2852_),
    .B2(net32),
    .A2(_2851_),
    .A1(net26));
 sg13g2_nand3_1 _8846_ (.B(_2850_),
    .C(_2853_),
    .A(_2706_),
    .Y(_2854_));
 sg13g2_o21ai_1 _8847_ (.B1(_2710_),
    .Y(_2855_),
    .A1(_2846_),
    .A2(_2854_));
 sg13g2_mux4_1 _8848_ (.S0(net134),
    .A0(\logix.ram_r[1185] ),
    .A1(\logix.ram_r[1193] ),
    .A2(\logix.ram_r[1201] ),
    .A3(\logix.ram_r[1209] ),
    .S1(net177),
    .X(_2856_));
 sg13g2_mux4_1 _8849_ (.S0(_2540_),
    .A0(\logix.ram_r[1153] ),
    .A1(\logix.ram_r[1161] ),
    .A2(\logix.ram_r[1169] ),
    .A3(\logix.ram_r[1177] ),
    .S1(net159),
    .X(_2857_));
 sg13g2_a22oi_1 _8850_ (.Y(_2858_),
    .B1(_2857_),
    .B2(net25),
    .A2(_2856_),
    .A1(net41));
 sg13g2_mux4_1 _8851_ (.S0(net117),
    .A0(\logix.ram_r[1249] ),
    .A1(\logix.ram_r[1257] ),
    .A2(\logix.ram_r[1265] ),
    .A3(\logix.ram_r[1273] ),
    .S1(net116),
    .X(_2859_));
 sg13g2_mux4_1 _8852_ (.S0(net152),
    .A0(\logix.ram_r[1217] ),
    .A1(\logix.ram_r[1225] ),
    .A2(\logix.ram_r[1233] ),
    .A3(\logix.ram_r[1241] ),
    .S1(net132),
    .X(_2860_));
 sg13g2_a22oi_1 _8853_ (.Y(_2861_),
    .B1(_2860_),
    .B2(net75),
    .A2(_2859_),
    .A1(net76));
 sg13g2_a21oi_1 _8854_ (.A1(_2858_),
    .A2(_2861_),
    .Y(_2862_),
    .B1(net71));
 sg13g2_mux4_1 _8855_ (.S0(_2477_),
    .A0(\logix.ram_r[1057] ),
    .A1(\logix.ram_r[1065] ),
    .A2(\logix.ram_r[1073] ),
    .A3(\logix.ram_r[1081] ),
    .S1(net162),
    .X(_2863_));
 sg13g2_mux4_1 _8856_ (.S0(net164),
    .A0(\logix.ram_r[1025] ),
    .A1(\logix.ram_r[1033] ),
    .A2(\logix.ram_r[1041] ),
    .A3(\logix.ram_r[1049] ),
    .S1(net163),
    .X(_2864_));
 sg13g2_a22oi_1 _8857_ (.Y(_2865_),
    .B1(_2864_),
    .B2(net38),
    .A2(_2863_),
    .A1(net39));
 sg13g2_mux4_1 _8858_ (.S0(net134),
    .A0(\logix.ram_r[1121] ),
    .A1(\logix.ram_r[1129] ),
    .A2(\logix.ram_r[1137] ),
    .A3(\logix.ram_r[1145] ),
    .S1(net177),
    .X(_2866_));
 sg13g2_mux4_1 _8859_ (.S0(_2540_),
    .A0(\logix.ram_r[1089] ),
    .A1(\logix.ram_r[1097] ),
    .A2(\logix.ram_r[1105] ),
    .A3(\logix.ram_r[1113] ),
    .S1(_2469_),
    .X(_2867_));
 sg13g2_a22oi_1 _8860_ (.Y(_2868_),
    .B1(_2867_),
    .B2(net72),
    .A2(_2866_),
    .A1(net73));
 sg13g2_a21oi_1 _8861_ (.A1(_2865_),
    .A2(_2868_),
    .Y(_2869_),
    .B1(net74));
 sg13g2_nor2_1 _8862_ (.A(_2862_),
    .B(_2869_),
    .Y(_2870_));
 sg13g2_nand3_1 _8863_ (.B(_2855_),
    .C(_2870_),
    .A(_2841_),
    .Y(_2871_));
 sg13g2_mux4_1 _8864_ (.S0(_2595_),
    .A0(\logix.ram_r[33] ),
    .A1(\logix.ram_r[41] ),
    .A2(\logix.ram_r[49] ),
    .A3(\logix.ram_r[57] ),
    .S1(net124),
    .X(_2872_));
 sg13g2_mux4_1 _8865_ (.S0(net145),
    .A0(\logix.ram_r[1] ),
    .A1(\logix.ram_r[9] ),
    .A2(\logix.ram_r[17] ),
    .A3(\logix.ram_r[25] ),
    .S1(net127),
    .X(_2873_));
 sg13g2_a22oi_1 _8866_ (.Y(_2874_),
    .B1(_2873_),
    .B2(net38),
    .A2(_2872_),
    .A1(net39));
 sg13g2_mux4_1 _8867_ (.S0(net144),
    .A0(\logix.ram_r[97] ),
    .A1(\logix.ram_r[105] ),
    .A2(\logix.ram_r[113] ),
    .A3(\logix.ram_r[121] ),
    .S1(net124),
    .X(_2875_));
 sg13g2_mux4_1 _8868_ (.S0(_2375_),
    .A0(\logix.ram_r[65] ),
    .A1(\logix.ram_r[73] ),
    .A2(\logix.ram_r[81] ),
    .A3(\logix.ram_r[89] ),
    .S1(net110),
    .X(_2876_));
 sg13g2_a22oi_1 _8869_ (.Y(_2877_),
    .B1(_2876_),
    .B2(net72),
    .A2(_2875_),
    .A1(net73));
 sg13g2_a21o_1 _8870_ (.A2(_2877_),
    .A1(_2874_),
    .B1(net74),
    .X(_2878_));
 sg13g2_buf_1 _8871_ (.A(_2458_),
    .X(_2879_));
 sg13g2_mux4_1 _8872_ (.S0(net131),
    .A0(\logix.ram_r[385] ),
    .A1(\logix.ram_r[393] ),
    .A2(\logix.ram_r[401] ),
    .A3(\logix.ram_r[409] ),
    .S1(net142),
    .X(_2880_));
 sg13g2_nand2_1 _8873_ (.Y(_2881_),
    .A(net95),
    .B(_2880_));
 sg13g2_mux4_1 _8874_ (.S0(net136),
    .A0(\logix.ram_r[417] ),
    .A1(\logix.ram_r[425] ),
    .A2(\logix.ram_r[433] ),
    .A3(\logix.ram_r[441] ),
    .S1(net135),
    .X(_2882_));
 sg13g2_nand2_1 _8875_ (.Y(_2883_),
    .A(net150),
    .B(_2882_));
 sg13g2_a21oi_1 _8876_ (.A1(_2881_),
    .A2(_2883_),
    .Y(_2884_),
    .B1(_2411_));
 sg13g2_mux2_1 _8877_ (.A0(\logix.ram_r[449] ),
    .A1(\logix.ram_r[457] ),
    .S(net119),
    .X(_2885_));
 sg13g2_mux2_1 _8878_ (.A0(\logix.ram_r[497] ),
    .A1(\logix.ram_r[505] ),
    .S(net146),
    .X(_2886_));
 sg13g2_a22oi_1 _8879_ (.Y(_2887_),
    .B1(_2886_),
    .B2(net26),
    .A2(_2885_),
    .A1(net27));
 sg13g2_mux2_1 _8880_ (.A0(\logix.ram_r[481] ),
    .A1(\logix.ram_r[489] ),
    .S(net96),
    .X(_2888_));
 sg13g2_mux2_1 _8881_ (.A0(\logix.ram_r[465] ),
    .A1(\logix.ram_r[473] ),
    .S(net144),
    .X(_2889_));
 sg13g2_a22oi_1 _8882_ (.Y(_2890_),
    .B1(_2889_),
    .B2(net32),
    .A2(_2888_),
    .A1(net33));
 sg13g2_nand2_1 _8883_ (.Y(_2891_),
    .A(_2887_),
    .B(_2890_));
 sg13g2_o21ai_1 _8884_ (.B1(net170),
    .Y(_2892_),
    .A1(_2884_),
    .A2(_2891_));
 sg13g2_mux4_1 _8885_ (.S0(net115),
    .A0(\logix.ram_r[257] ),
    .A1(\logix.ram_r[265] ),
    .A2(\logix.ram_r[273] ),
    .A3(\logix.ram_r[281] ),
    .S1(net167),
    .X(_2893_));
 sg13g2_nand2_1 _8886_ (.Y(_2894_),
    .A(net123),
    .B(_2893_));
 sg13g2_mux4_1 _8887_ (.S0(_2474_),
    .A0(\logix.ram_r[289] ),
    .A1(\logix.ram_r[297] ),
    .A2(\logix.ram_r[305] ),
    .A3(\logix.ram_r[313] ),
    .S1(_2475_),
    .X(_2895_));
 sg13g2_nand2_1 _8888_ (.Y(_2896_),
    .A(net179),
    .B(_2895_));
 sg13g2_nand3_1 _8889_ (.B(_2894_),
    .C(_2896_),
    .A(net174),
    .Y(_2897_));
 sg13g2_nand2b_1 _8890_ (.Y(_2898_),
    .B(net163),
    .A_N(\logix.ram_r[337] ));
 sg13g2_o21ai_1 _8891_ (.B1(_2898_),
    .Y(_2899_),
    .A1(\logix.ram_r[321] ),
    .A2(net59));
 sg13g2_buf_8 _8892_ (.A(_2475_),
    .X(_2900_));
 sg13g2_nand2b_1 _8893_ (.Y(_2901_),
    .B(_2650_),
    .A_N(\logix.ram_r[345] ));
 sg13g2_o21ai_1 _8894_ (.B1(_2901_),
    .Y(_2902_),
    .A1(\logix.ram_r[329] ),
    .A2(net58));
 sg13g2_a22oi_1 _8895_ (.Y(_2903_),
    .B1(_2902_),
    .B2(_2647_),
    .A2(_2899_),
    .A1(_2639_));
 sg13g2_mux4_1 _8896_ (.S0(net146),
    .A0(\logix.ram_r[353] ),
    .A1(\logix.ram_r[361] ),
    .A2(\logix.ram_r[369] ),
    .A3(\logix.ram_r[377] ),
    .S1(net128),
    .X(_2904_));
 sg13g2_nand2b_1 _8897_ (.Y(_2905_),
    .B(net65),
    .A_N(_2904_));
 sg13g2_nand4_1 _8898_ (.B(_2897_),
    .C(_2903_),
    .A(net79),
    .Y(_2906_),
    .D(_2905_));
 sg13g2_mux4_1 _8899_ (.S0(net100),
    .A0(\logix.ram_r[161] ),
    .A1(\logix.ram_r[169] ),
    .A2(\logix.ram_r[177] ),
    .A3(\logix.ram_r[185] ),
    .S1(net142),
    .X(_2907_));
 sg13g2_mux4_1 _8900_ (.S0(net105),
    .A0(\logix.ram_r[129] ),
    .A1(\logix.ram_r[137] ),
    .A2(\logix.ram_r[145] ),
    .A3(\logix.ram_r[153] ),
    .S1(net130),
    .X(_2908_));
 sg13g2_a22oi_1 _8901_ (.Y(_2909_),
    .B1(_2908_),
    .B2(net30),
    .A2(_2907_),
    .A1(net31));
 sg13g2_buf_8 _8902_ (.A(_2562_),
    .X(_2910_));
 sg13g2_mux4_1 _8903_ (.S0(net94),
    .A0(\logix.ram_r[225] ),
    .A1(\logix.ram_r[233] ),
    .A2(\logix.ram_r[241] ),
    .A3(\logix.ram_r[249] ),
    .S1(net114),
    .X(_2911_));
 sg13g2_mux4_1 _8904_ (.S0(net106),
    .A0(\logix.ram_r[193] ),
    .A1(\logix.ram_r[201] ),
    .A2(\logix.ram_r[209] ),
    .A3(\logix.ram_r[217] ),
    .S1(net112),
    .X(_2912_));
 sg13g2_a22oi_1 _8905_ (.Y(_2913_),
    .B1(_2912_),
    .B2(net61),
    .A2(_2911_),
    .A1(net62));
 sg13g2_a21oi_1 _8906_ (.A1(_2909_),
    .A2(_2913_),
    .Y(_2914_),
    .B1(net67));
 sg13g2_nor2_1 _8907_ (.A(_2455_),
    .B(_2914_),
    .Y(_2915_));
 sg13g2_nand4_1 _8908_ (.B(_2892_),
    .C(_2906_),
    .A(_2878_),
    .Y(_2916_),
    .D(_2915_));
 sg13g2_and4_1 _8909_ (.A(_2778_),
    .B(_2828_),
    .C(_2871_),
    .D(_2916_),
    .X(net15));
 sg13g2_buf_2 _8910_ (.A(_2515_),
    .X(_2917_));
 sg13g2_mux4_1 _8911_ (.S0(net195),
    .A0(\logix.ram_r[898] ),
    .A1(\logix.ram_r[906] ),
    .A2(\logix.ram_r[914] ),
    .A3(\logix.ram_r[922] ),
    .S1(net186),
    .X(_2918_));
 sg13g2_nor2_1 _8912_ (.A(net188),
    .B(_2918_),
    .Y(_2919_));
 sg13g2_mux2_1 _8913_ (.A0(\logix.ram_r[930] ),
    .A1(\logix.ram_r[946] ),
    .S(net190),
    .X(_2920_));
 sg13g2_nor2_1 _8914_ (.A(_2344_),
    .B(_2920_),
    .Y(_2921_));
 sg13g2_mux2_1 _8915_ (.A0(\logix.ram_r[938] ),
    .A1(\logix.ram_r[954] ),
    .S(net190),
    .X(_2922_));
 sg13g2_o21ai_1 _8916_ (.B1(_2362_),
    .Y(_2923_),
    .A1(_2352_),
    .A2(_2922_));
 sg13g2_nor3_1 _8917_ (.A(_2919_),
    .B(_2921_),
    .C(_2923_),
    .Y(_2924_));
 sg13g2_mux2_1 _8918_ (.A0(\logix.ram_r[994] ),
    .A1(\logix.ram_r[1002] ),
    .S(net133),
    .X(_2925_));
 sg13g2_mux2_1 _8919_ (.A0(\logix.ram_r[978] ),
    .A1(\logix.ram_r[986] ),
    .S(_2425_),
    .X(_2926_));
 sg13g2_a22oi_1 _8920_ (.Y(_2927_),
    .B1(_2926_),
    .B2(_2624_),
    .A2(_2925_),
    .A1(_2621_));
 sg13g2_mux2_1 _8921_ (.A0(\logix.ram_r[962] ),
    .A1(\logix.ram_r[970] ),
    .S(net166),
    .X(_2928_));
 sg13g2_mux2_1 _8922_ (.A0(\logix.ram_r[1010] ),
    .A1(\logix.ram_r[1018] ),
    .S(net164),
    .X(_2929_));
 sg13g2_a22oi_1 _8923_ (.Y(_2930_),
    .B1(_2929_),
    .B2(net26),
    .A2(_2928_),
    .A1(net27));
 sg13g2_nand2_1 _8924_ (.Y(_2931_),
    .A(_2927_),
    .B(_2930_));
 sg13g2_o21ai_1 _8925_ (.B1(net170),
    .Y(_2932_),
    .A1(_2924_),
    .A2(_2931_));
 sg13g2_mux4_1 _8926_ (.S0(net192),
    .A0(\logix.ram_r[770] ),
    .A1(\logix.ram_r[786] ),
    .A2(\logix.ram_r[802] ),
    .A3(\logix.ram_r[818] ),
    .S1(net204),
    .X(_2933_));
 sg13g2_mux4_1 _8927_ (.S0(net192),
    .A0(\logix.ram_r[778] ),
    .A1(\logix.ram_r[794] ),
    .A2(\logix.ram_r[810] ),
    .A3(\logix.ram_r[826] ),
    .S1(_2325_),
    .X(_2934_));
 sg13g2_buf_8 _8928_ (.A(_2468_),
    .X(_2935_));
 sg13g2_mux2_1 _8929_ (.A0(_2933_),
    .A1(_2934_),
    .S(net57),
    .X(_2936_));
 sg13g2_buf_8 _8930_ (.A(_2350_),
    .X(_2937_));
 sg13g2_buf_8 _8931_ (.A(_2354_),
    .X(_2938_));
 sg13g2_mux4_1 _8932_ (.S0(net185),
    .A0(\logix.ram_r[834] ),
    .A1(\logix.ram_r[842] ),
    .A2(\logix.ram_r[850] ),
    .A3(\logix.ram_r[858] ),
    .S1(net93),
    .X(_2939_));
 sg13g2_nor2_1 _8933_ (.A(net202),
    .B(_2939_),
    .Y(_2940_));
 sg13g2_buf_8 _8934_ (.A(_2515_),
    .X(_2941_));
 sg13g2_mux2_1 _8935_ (.A0(\logix.ram_r[874] ),
    .A1(\logix.ram_r[890] ),
    .S(net184),
    .X(_2942_));
 sg13g2_nor2_1 _8936_ (.A(_2433_),
    .B(_2942_),
    .Y(_2943_));
 sg13g2_mux2_1 _8937_ (.A0(\logix.ram_r[866] ),
    .A1(\logix.ram_r[882] ),
    .S(net190),
    .X(_2944_));
 sg13g2_o21ai_1 _8938_ (.B1(_2444_),
    .Y(_2945_),
    .A1(_2439_),
    .A2(_2944_));
 sg13g2_nor3_1 _8939_ (.A(_2940_),
    .B(_2943_),
    .C(_2945_),
    .Y(_2946_));
 sg13g2_o21ai_1 _8940_ (.B1(_2946_),
    .Y(_2947_),
    .A1(net120),
    .A2(_2936_));
 sg13g2_mux4_1 _8941_ (.S0(net200),
    .A0(\logix.ram_r[674] ),
    .A1(\logix.ram_r[682] ),
    .A2(\logix.ram_r[690] ),
    .A3(\logix.ram_r[698] ),
    .S1(net186),
    .X(_2948_));
 sg13g2_mux4_1 _8942_ (.S0(net201),
    .A0(\logix.ram_r[642] ),
    .A1(\logix.ram_r[650] ),
    .A2(\logix.ram_r[658] ),
    .A3(\logix.ram_r[666] ),
    .S1(net197),
    .X(_2949_));
 sg13g2_a22oi_1 _8943_ (.Y(_2950_),
    .B1(_2949_),
    .B2(_2466_),
    .A2(_2948_),
    .A1(net78));
 sg13g2_mux4_1 _8944_ (.S0(_2527_),
    .A0(\logix.ram_r[738] ),
    .A1(\logix.ram_r[746] ),
    .A2(\logix.ram_r[754] ),
    .A3(\logix.ram_r[762] ),
    .S1(net192),
    .X(_2951_));
 sg13g2_mux4_1 _8945_ (.S0(_2523_),
    .A0(\logix.ram_r[706] ),
    .A1(\logix.ram_r[714] ),
    .A2(\logix.ram_r[722] ),
    .A3(\logix.ram_r[730] ),
    .S1(_2736_),
    .X(_2952_));
 sg13g2_a22oi_1 _8946_ (.Y(_2953_),
    .B1(_2952_),
    .B2(net154),
    .A2(_2951_),
    .A1(net126));
 sg13g2_a21oi_1 _8947_ (.A1(_2950_),
    .A2(_2953_),
    .Y(_2954_),
    .B1(_2502_));
 sg13g2_buf_2 _8948_ (.A(_2459_),
    .X(_2955_));
 sg13g2_mux4_1 _8949_ (.S0(net203),
    .A0(\logix.ram_r[546] ),
    .A1(\logix.ram_r[554] ),
    .A2(\logix.ram_r[562] ),
    .A3(\logix.ram_r[570] ),
    .S1(net184),
    .X(_2956_));
 sg13g2_buf_8 _8950_ (.A(_2350_),
    .X(_2957_));
 sg13g2_mux4_1 _8951_ (.S0(net183),
    .A0(\logix.ram_r[514] ),
    .A1(\logix.ram_r[522] ),
    .A2(\logix.ram_r[530] ),
    .A3(\logix.ram_r[538] ),
    .S1(net175),
    .X(_2958_));
 sg13g2_buf_2 _8952_ (.A(_2465_),
    .X(_2959_));
 sg13g2_a22oi_1 _8953_ (.Y(_2960_),
    .B1(_2958_),
    .B2(net55),
    .A2(_2956_),
    .A1(net56));
 sg13g2_mux4_1 _8954_ (.S0(net200),
    .A0(\logix.ram_r[610] ),
    .A1(\logix.ram_r[618] ),
    .A2(\logix.ram_r[626] ),
    .A3(\logix.ram_r[634] ),
    .S1(net193),
    .X(_2961_));
 sg13g2_buf_8 _8955_ (.A(_2350_),
    .X(_2962_));
 sg13g2_buf_8 _8956_ (.A(_2354_),
    .X(_2963_));
 sg13g2_mux4_1 _8957_ (.S0(net182),
    .A0(\logix.ram_r[578] ),
    .A1(\logix.ram_r[586] ),
    .A2(\logix.ram_r[594] ),
    .A3(\logix.ram_r[602] ),
    .S1(_2963_),
    .X(_2964_));
 sg13g2_buf_2 _8958_ (.A(_2480_),
    .X(_2965_));
 sg13g2_a22oi_1 _8959_ (.Y(_2966_),
    .B1(_2964_),
    .B2(net91),
    .A2(_2961_),
    .A1(net126));
 sg13g2_buf_2 _8960_ (.A(_2485_),
    .X(_2967_));
 sg13g2_a21oi_1 _8961_ (.A1(_2960_),
    .A2(_2966_),
    .Y(_2968_),
    .B1(net54));
 sg13g2_nor2_1 _8962_ (.A(_2954_),
    .B(_2968_),
    .Y(_2969_));
 sg13g2_and4_1 _8963_ (.A(_2553_),
    .B(_2932_),
    .C(_2947_),
    .D(_2969_),
    .X(_2970_));
 sg13g2_nand2b_1 _8964_ (.Y(_2971_),
    .B(net59),
    .A_N(\logix.ram_r[1490] ));
 sg13g2_o21ai_1 _8965_ (.B1(_2971_),
    .Y(_2972_),
    .A1(\logix.ram_r[1474] ),
    .A2(net60));
 sg13g2_buf_8 _8966_ (.A(net111),
    .X(_2973_));
 sg13g2_nand2b_1 _8967_ (.Y(_2974_),
    .B(net58),
    .A_N(\logix.ram_r[1498] ));
 sg13g2_o21ai_1 _8968_ (.B1(_2974_),
    .Y(_2975_),
    .A1(\logix.ram_r[1482] ),
    .A2(net53));
 sg13g2_a221oi_1 _8969_ (.B2(net28),
    .C1(_2603_),
    .B1(_2975_),
    .A1(net29),
    .Y(_2976_),
    .A2(_2972_));
 sg13g2_buf_1 _8970_ (.A(_2358_),
    .X(_2977_));
 sg13g2_buf_2 _8971_ (.A(_2360_),
    .X(_2978_));
 sg13g2_mux4_1 _8972_ (.S0(net96),
    .A0(\logix.ram_r[1442] ),
    .A1(\logix.ram_r[1450] ),
    .A2(\logix.ram_r[1458] ),
    .A3(\logix.ram_r[1466] ),
    .S1(net113),
    .X(_2979_));
 sg13g2_buf_8 _8973_ (.A(_2535_),
    .X(_2980_));
 sg13g2_mux4_1 _8974_ (.S0(net200),
    .A0(\logix.ram_r[1410] ),
    .A1(\logix.ram_r[1418] ),
    .A2(\logix.ram_r[1426] ),
    .A3(\logix.ram_r[1434] ),
    .S1(net186),
    .X(_2981_));
 sg13g2_and2_1 _8975_ (.A(_2458_),
    .B(_2981_),
    .X(_2982_));
 sg13g2_a221oi_1 _8976_ (.B2(_2980_),
    .C1(_2982_),
    .B1(_2979_),
    .A1(_2977_),
    .Y(_2983_),
    .A2(_2978_));
 sg13g2_buf_1 _8977_ (.A(_2370_),
    .X(_2984_));
 sg13g2_buf_8 _8978_ (.A(_2562_),
    .X(_2985_));
 sg13g2_buf_8 _8979_ (.A(net88),
    .X(_2986_));
 sg13g2_mux4_1 _8980_ (.S0(_2986_),
    .A0(\logix.ram_r[1506] ),
    .A1(\logix.ram_r[1514] ),
    .A2(\logix.ram_r[1522] ),
    .A3(\logix.ram_r[1530] ),
    .S1(_2641_),
    .X(_2987_));
 sg13g2_nor2_1 _8981_ (.A(_2984_),
    .B(_2987_),
    .Y(_2988_));
 sg13g2_nor2_1 _8982_ (.A(_2983_),
    .B(_2988_),
    .Y(_2989_));
 sg13g2_buf_2 _8983_ (.A(_2515_),
    .X(_2990_));
 sg13g2_mux4_1 _8984_ (.S0(net196),
    .A0(\logix.ram_r[1282] ),
    .A1(\logix.ram_r[1290] ),
    .A2(\logix.ram_r[1298] ),
    .A3(\logix.ram_r[1306] ),
    .S1(net181),
    .X(_2991_));
 sg13g2_buf_8 _8985_ (.A(_2350_),
    .X(_2992_));
 sg13g2_mux4_1 _8986_ (.S0(net180),
    .A0(\logix.ram_r[1314] ),
    .A1(\logix.ram_r[1322] ),
    .A2(\logix.ram_r[1330] ),
    .A3(\logix.ram_r[1338] ),
    .S1(net181),
    .X(_2993_));
 sg13g2_mux2_1 _8987_ (.A0(_2991_),
    .A1(_2993_),
    .S(net194),
    .X(_2994_));
 sg13g2_nand2_1 _8988_ (.Y(_2995_),
    .A(net118),
    .B(_2994_));
 sg13g2_mux2_1 _8989_ (.A0(\logix.ram_r[1346] ),
    .A1(\logix.ram_r[1354] ),
    .S(net52),
    .X(_2996_));
 sg13g2_buf_8 _8990_ (.A(_2463_),
    .X(_2997_));
 sg13g2_mux2_1 _8991_ (.A0(\logix.ram_r[1394] ),
    .A1(\logix.ram_r[1402] ),
    .S(net51),
    .X(_2998_));
 sg13g2_a22oi_1 _8992_ (.Y(_2999_),
    .B1(_2998_),
    .B2(net45),
    .A2(_2996_),
    .A1(net46));
 sg13g2_mux2_1 _8993_ (.A0(\logix.ram_r[1378] ),
    .A1(\logix.ram_r[1386] ),
    .S(net52),
    .X(_3000_));
 sg13g2_mux2_1 _8994_ (.A0(\logix.ram_r[1362] ),
    .A1(\logix.ram_r[1370] ),
    .S(net51),
    .X(_3001_));
 sg13g2_a22oi_1 _8995_ (.Y(_3002_),
    .B1(_3001_),
    .B2(net47),
    .A2(_3000_),
    .A1(net48));
 sg13g2_nand4_1 _8996_ (.B(_2995_),
    .C(_2999_),
    .A(_2706_),
    .Y(_3003_),
    .D(_3002_));
 sg13g2_mux4_1 _8997_ (.S0(net196),
    .A0(\logix.ram_r[1186] ),
    .A1(\logix.ram_r[1194] ),
    .A2(\logix.ram_r[1202] ),
    .A3(\logix.ram_r[1210] ),
    .S1(net189),
    .X(_3004_));
 sg13g2_mux4_1 _8998_ (.S0(net88),
    .A0(\logix.ram_r[1154] ),
    .A1(\logix.ram_r[1162] ),
    .A2(\logix.ram_r[1170] ),
    .A3(\logix.ram_r[1178] ),
    .S1(net108),
    .X(_3005_));
 sg13g2_a22oi_1 _8999_ (.Y(_3006_),
    .B1(_3005_),
    .B2(net55),
    .A2(_3004_),
    .A1(net56));
 sg13g2_mux4_1 _9000_ (.S0(net203),
    .A0(\logix.ram_r[1250] ),
    .A1(\logix.ram_r[1258] ),
    .A2(\logix.ram_r[1266] ),
    .A3(\logix.ram_r[1274] ),
    .S1(net184),
    .X(_3007_));
 sg13g2_mux4_1 _9001_ (.S0(net183),
    .A0(\logix.ram_r[1218] ),
    .A1(\logix.ram_r[1226] ),
    .A2(\logix.ram_r[1234] ),
    .A3(\logix.ram_r[1242] ),
    .S1(net175),
    .X(_3008_));
 sg13g2_a22oi_1 _9002_ (.Y(_3009_),
    .B1(_3008_),
    .B2(net91),
    .A2(_3007_),
    .A1(net126));
 sg13g2_buf_2 _9003_ (.A(_2502_),
    .X(_3010_));
 sg13g2_a21oi_1 _9004_ (.A1(_3006_),
    .A2(_3009_),
    .Y(_3011_),
    .B1(_3010_));
 sg13g2_mux4_1 _9005_ (.S0(net201),
    .A0(\logix.ram_r[1058] ),
    .A1(\logix.ram_r[1066] ),
    .A2(\logix.ram_r[1074] ),
    .A3(\logix.ram_r[1082] ),
    .S1(net197),
    .X(_3012_));
 sg13g2_buf_8 _9006_ (.A(_2562_),
    .X(_3013_));
 sg13g2_buf_8 _9007_ (.A(_2346_),
    .X(_3014_));
 sg13g2_mux4_1 _9008_ (.S0(net87),
    .A0(\logix.ram_r[1026] ),
    .A1(\logix.ram_r[1034] ),
    .A2(\logix.ram_r[1042] ),
    .A3(\logix.ram_r[1050] ),
    .S1(net86),
    .X(_3015_));
 sg13g2_a22oi_1 _9009_ (.Y(_3016_),
    .B1(_3015_),
    .B2(net55),
    .A2(_3012_),
    .A1(net56));
 sg13g2_mux4_1 _9010_ (.S0(net180),
    .A0(\logix.ram_r[1122] ),
    .A1(\logix.ram_r[1130] ),
    .A2(\logix.ram_r[1138] ),
    .A3(\logix.ram_r[1146] ),
    .S1(_2990_),
    .X(_3017_));
 sg13g2_mux4_1 _9011_ (.S0(net183),
    .A0(\logix.ram_r[1090] ),
    .A1(\logix.ram_r[1098] ),
    .A2(\logix.ram_r[1106] ),
    .A3(\logix.ram_r[1114] ),
    .S1(net108),
    .X(_3018_));
 sg13g2_a22oi_1 _9012_ (.Y(_3019_),
    .B1(_3018_),
    .B2(net91),
    .A2(_3017_),
    .A1(_2593_));
 sg13g2_a21oi_1 _9013_ (.A1(_3016_),
    .A2(_3019_),
    .Y(_3020_),
    .B1(net54));
 sg13g2_or2_1 _9014_ (.X(_3021_),
    .B(_3020_),
    .A(_3011_));
 sg13g2_a221oi_1 _9015_ (.B2(_2710_),
    .C1(_3021_),
    .B1(_3003_),
    .A1(_2976_),
    .Y(_3022_),
    .A2(_2989_));
 sg13g2_nand2b_1 _9016_ (.Y(_3023_),
    .B(net64),
    .A_N(\logix.ram_r[1874] ));
 sg13g2_o21ai_1 _9017_ (.B1(_3023_),
    .Y(_3024_),
    .A1(\logix.ram_r[1858] ),
    .A2(net60));
 sg13g2_nand2b_1 _9018_ (.Y(_3025_),
    .B(net63),
    .A_N(\logix.ram_r[1882] ));
 sg13g2_o21ai_1 _9019_ (.B1(_3025_),
    .Y(_3026_),
    .A1(\logix.ram_r[1866] ),
    .A2(net53));
 sg13g2_a221oi_1 _9020_ (.B2(net28),
    .C1(_2709_),
    .B1(_3026_),
    .A1(net29),
    .Y(_3027_),
    .A2(_3024_));
 sg13g2_mux4_1 _9021_ (.S0(net107),
    .A0(\logix.ram_r[1826] ),
    .A1(\logix.ram_r[1834] ),
    .A2(\logix.ram_r[1842] ),
    .A3(\logix.ram_r[1850] ),
    .S1(net111),
    .X(_3028_));
 sg13g2_mux4_1 _9022_ (.S0(net180),
    .A0(\logix.ram_r[1794] ),
    .A1(\logix.ram_r[1802] ),
    .A2(\logix.ram_r[1810] ),
    .A3(\logix.ram_r[1818] ),
    .S1(net181),
    .X(_3029_));
 sg13g2_and2_1 _9023_ (.A(net95),
    .B(_3029_),
    .X(_3030_));
 sg13g2_a221oi_1 _9024_ (.B2(net90),
    .C1(_3030_),
    .B1(_3028_),
    .A1(net206),
    .Y(_3031_),
    .A2(net205));
 sg13g2_buf_8 _9025_ (.A(net122),
    .X(_3032_));
 sg13g2_mux4_1 _9026_ (.S0(net49),
    .A0(\logix.ram_r[1890] ),
    .A1(\logix.ram_r[1898] ),
    .A2(\logix.ram_r[1906] ),
    .A3(\logix.ram_r[1914] ),
    .S1(net58),
    .X(_3033_));
 sg13g2_nor2_1 _9027_ (.A(net89),
    .B(_3033_),
    .Y(_3034_));
 sg13g2_nor2_1 _9028_ (.A(_3031_),
    .B(_3034_),
    .Y(_3035_));
 sg13g2_mux4_1 _9029_ (.S0(net185),
    .A0(\logix.ram_r[1922] ),
    .A1(\logix.ram_r[1930] ),
    .A2(\logix.ram_r[1938] ),
    .A3(\logix.ram_r[1946] ),
    .S1(net93),
    .X(_3036_));
 sg13g2_mux4_1 _9030_ (.S0(net182),
    .A0(\logix.ram_r[1954] ),
    .A1(\logix.ram_r[1962] ),
    .A2(\logix.ram_r[1970] ),
    .A3(\logix.ram_r[1978] ),
    .S1(net92),
    .X(_3037_));
 sg13g2_mux2_1 _9031_ (.A0(_3036_),
    .A1(_3037_),
    .S(net199),
    .X(_3038_));
 sg13g2_nand2_1 _9032_ (.Y(_3039_),
    .A(net118),
    .B(_3038_));
 sg13g2_mux2_1 _9033_ (.A0(\logix.ram_r[1986] ),
    .A1(\logix.ram_r[1994] ),
    .S(net51),
    .X(_3040_));
 sg13g2_mux2_1 _9034_ (.A0(\logix.ram_r[2034] ),
    .A1(\logix.ram_r[2042] ),
    .S(net80),
    .X(_3041_));
 sg13g2_a22oi_1 _9035_ (.Y(_3042_),
    .B1(_3041_),
    .B2(net45),
    .A2(_3040_),
    .A1(net46));
 sg13g2_mux2_1 _9036_ (.A0(\logix.ram_r[2018] ),
    .A1(\logix.ram_r[2026] ),
    .S(net49),
    .X(_3043_));
 sg13g2_mux2_1 _9037_ (.A0(\logix.ram_r[2002] ),
    .A1(\logix.ram_r[2010] ),
    .S(net80),
    .X(_3044_));
 sg13g2_a22oi_1 _9038_ (.Y(_3045_),
    .B1(_3044_),
    .B2(net47),
    .A2(_3043_),
    .A1(net48));
 sg13g2_nand4_1 _9039_ (.B(_3039_),
    .C(_3042_),
    .A(_2780_),
    .Y(_3046_),
    .D(_3045_));
 sg13g2_nand2_1 _9040_ (.Y(_3047_),
    .A(_2603_),
    .B(_2780_));
 sg13g2_buf_8 _9041_ (.A(net78),
    .X(_3048_));
 sg13g2_mux4_1 _9042_ (.S0(net185),
    .A0(\logix.ram_r[1570] ),
    .A1(\logix.ram_r[1578] ),
    .A2(\logix.ram_r[1586] ),
    .A3(\logix.ram_r[1594] ),
    .S1(net175),
    .X(_3049_));
 sg13g2_mux4_1 _9043_ (.S0(net136),
    .A0(\logix.ram_r[1538] ),
    .A1(\logix.ram_r[1546] ),
    .A2(\logix.ram_r[1554] ),
    .A3(\logix.ram_r[1562] ),
    .S1(net101),
    .X(_3050_));
 sg13g2_buf_8 _9044_ (.A(net77),
    .X(_3051_));
 sg13g2_a22oi_1 _9045_ (.Y(_3052_),
    .B1(_3050_),
    .B2(net22),
    .A2(_3049_),
    .A1(net23));
 sg13g2_buf_2 _9046_ (.A(_2431_),
    .X(_3053_));
 sg13g2_mux4_1 _9047_ (.S0(net201),
    .A0(\logix.ram_r[1634] ),
    .A1(\logix.ram_r[1642] ),
    .A2(\logix.ram_r[1650] ),
    .A3(\logix.ram_r[1658] ),
    .S1(net197),
    .X(_3054_));
 sg13g2_mux4_1 _9048_ (.S0(net87),
    .A0(\logix.ram_r[1602] ),
    .A1(\logix.ram_r[1610] ),
    .A2(\logix.ram_r[1618] ),
    .A3(\logix.ram_r[1626] ),
    .S1(net86),
    .X(_3055_));
 sg13g2_buf_2 _9049_ (.A(_2480_),
    .X(_3056_));
 sg13g2_a22oi_1 _9050_ (.Y(_3057_),
    .B1(_3055_),
    .B2(net84),
    .A2(_3054_),
    .A1(net85));
 sg13g2_a21oi_1 _9051_ (.A1(_3052_),
    .A2(_3057_),
    .Y(_3058_),
    .B1(net54));
 sg13g2_mux4_1 _9052_ (.S0(net183),
    .A0(\logix.ram_r[1698] ),
    .A1(\logix.ram_r[1706] ),
    .A2(\logix.ram_r[1714] ),
    .A3(\logix.ram_r[1722] ),
    .S1(net99),
    .X(_3059_));
 sg13g2_mux4_1 _9053_ (.S0(net100),
    .A0(\logix.ram_r[1666] ),
    .A1(\logix.ram_r[1674] ),
    .A2(\logix.ram_r[1682] ),
    .A3(\logix.ram_r[1690] ),
    .S1(net176),
    .X(_3060_));
 sg13g2_a22oi_1 _9054_ (.Y(_3061_),
    .B1(_3060_),
    .B2(net22),
    .A2(_3059_),
    .A1(net23));
 sg13g2_mux4_1 _9055_ (.S0(net182),
    .A0(\logix.ram_r[1762] ),
    .A1(\logix.ram_r[1770] ),
    .A2(\logix.ram_r[1778] ),
    .A3(\logix.ram_r[1786] ),
    .S1(net93),
    .X(_3062_));
 sg13g2_mux4_1 _9056_ (.S0(net94),
    .A0(\logix.ram_r[1730] ),
    .A1(\logix.ram_r[1738] ),
    .A2(\logix.ram_r[1746] ),
    .A3(\logix.ram_r[1754] ),
    .S1(net147),
    .X(_3063_));
 sg13g2_a22oi_1 _9057_ (.Y(_3064_),
    .B1(_3063_),
    .B2(net84),
    .A2(_3062_),
    .A1(net85));
 sg13g2_a21oi_1 _9058_ (.A1(_3061_),
    .A2(_3064_),
    .Y(_3065_),
    .B1(net50));
 sg13g2_or2_1 _9059_ (.X(_3066_),
    .B(_3065_),
    .A(_3058_));
 sg13g2_a221oi_1 _9060_ (.B2(_3047_),
    .C1(_3066_),
    .B1(_3046_),
    .A1(_3027_),
    .Y(_3067_),
    .A2(_3035_));
 sg13g2_nand2b_1 _9061_ (.Y(_3068_),
    .B(net58),
    .A_N(\logix.ram_r[338] ));
 sg13g2_o21ai_1 _9062_ (.B1(_3068_),
    .Y(_3069_),
    .A1(\logix.ram_r[322] ),
    .A2(net53));
 sg13g2_nand2b_1 _9063_ (.Y(_3070_),
    .B(_2681_),
    .A_N(\logix.ram_r[346] ));
 sg13g2_o21ai_1 _9064_ (.B1(_3070_),
    .Y(_3071_),
    .A1(\logix.ram_r[330] ),
    .A2(net53));
 sg13g2_a221oi_1 _9065_ (.B2(_2684_),
    .C1(_2709_),
    .B1(_3071_),
    .A1(net29),
    .Y(_3072_),
    .A2(_3069_));
 sg13g2_mux4_1 _9066_ (.S0(net146),
    .A0(\logix.ram_r[290] ),
    .A1(\logix.ram_r[298] ),
    .A2(\logix.ram_r[306] ),
    .A3(\logix.ram_r[314] ),
    .S1(net128),
    .X(_3073_));
 sg13g2_mux4_1 _9067_ (.S0(net185),
    .A0(\logix.ram_r[258] ),
    .A1(\logix.ram_r[266] ),
    .A2(\logix.ram_r[274] ),
    .A3(\logix.ram_r[282] ),
    .S1(net93),
    .X(_3074_));
 sg13g2_and2_1 _9068_ (.A(net95),
    .B(_3074_),
    .X(_3075_));
 sg13g2_a221oi_1 _9069_ (.B2(net90),
    .C1(_3075_),
    .B1(_3073_),
    .A1(net206),
    .Y(_3076_),
    .A2(net205));
 sg13g2_mux4_1 _9070_ (.S0(_2997_),
    .A0(\logix.ram_r[354] ),
    .A1(\logix.ram_r[362] ),
    .A2(\logix.ram_r[370] ),
    .A3(\logix.ram_r[378] ),
    .S1(net63),
    .X(_3077_));
 sg13g2_nor2_1 _9071_ (.A(net89),
    .B(_3077_),
    .Y(_3078_));
 sg13g2_nor2_1 _9072_ (.A(_3076_),
    .B(_3078_),
    .Y(_3079_));
 sg13g2_mux4_1 _9073_ (.S0(net109),
    .A0(\logix.ram_r[386] ),
    .A1(\logix.ram_r[394] ),
    .A2(\logix.ram_r[402] ),
    .A3(\logix.ram_r[410] ),
    .S1(net104),
    .X(_3080_));
 sg13g2_mux4_1 _9074_ (.S0(net88),
    .A0(\logix.ram_r[418] ),
    .A1(\logix.ram_r[426] ),
    .A2(\logix.ram_r[434] ),
    .A3(\logix.ram_r[442] ),
    .S1(net97),
    .X(_3081_));
 sg13g2_mux2_1 _9075_ (.A0(_3080_),
    .A1(_3081_),
    .S(net188),
    .X(_3082_));
 sg13g2_nand2_1 _9076_ (.Y(_3083_),
    .A(net118),
    .B(_3082_));
 sg13g2_mux2_1 _9077_ (.A0(\logix.ram_r[450] ),
    .A1(\logix.ram_r[458] ),
    .S(_2420_),
    .X(_3084_));
 sg13g2_mux2_1 _9078_ (.A0(\logix.ram_r[498] ),
    .A1(\logix.ram_r[506] ),
    .S(net57),
    .X(_3085_));
 sg13g2_a22oi_1 _9079_ (.Y(_3086_),
    .B1(_3085_),
    .B2(_2396_),
    .A2(_3084_),
    .A1(_2390_));
 sg13g2_mux2_1 _9080_ (.A0(\logix.ram_r[482] ),
    .A1(\logix.ram_r[490] ),
    .S(net80),
    .X(_3087_));
 sg13g2_mux2_1 _9081_ (.A0(\logix.ram_r[466] ),
    .A1(\logix.ram_r[474] ),
    .S(net57),
    .X(_3088_));
 sg13g2_a22oi_1 _9082_ (.Y(_3089_),
    .B1(_3088_),
    .B2(_2383_),
    .A2(_3087_),
    .A1(net48));
 sg13g2_nand4_1 _9083_ (.B(_3083_),
    .C(_3086_),
    .A(_2456_),
    .Y(_3090_),
    .D(_3089_));
 sg13g2_nand2_1 _9084_ (.Y(_3091_),
    .A(_2603_),
    .B(_2456_));
 sg13g2_mux4_1 _9085_ (.S0(net109),
    .A0(\logix.ram_r[34] ),
    .A1(\logix.ram_r[42] ),
    .A2(\logix.ram_r[50] ),
    .A3(\logix.ram_r[58] ),
    .S1(net147),
    .X(_3092_));
 sg13g2_mux4_1 _9086_ (.S0(net149),
    .A0(\logix.ram_r[2] ),
    .A1(\logix.ram_r[10] ),
    .A2(\logix.ram_r[18] ),
    .A3(\logix.ram_r[26] ),
    .S1(net116),
    .X(_3093_));
 sg13g2_a22oi_1 _9087_ (.Y(_3094_),
    .B1(_3093_),
    .B2(net22),
    .A2(_3092_),
    .A1(net23));
 sg13g2_mux4_1 _9088_ (.S0(net88),
    .A0(\logix.ram_r[98] ),
    .A1(\logix.ram_r[106] ),
    .A2(\logix.ram_r[114] ),
    .A3(\logix.ram_r[122] ),
    .S1(net108),
    .X(_3095_));
 sg13g2_mux4_1 _9089_ (.S0(net139),
    .A0(\logix.ram_r[66] ),
    .A1(\logix.ram_r[74] ),
    .A2(\logix.ram_r[82] ),
    .A3(\logix.ram_r[90] ),
    .S1(net138),
    .X(_3096_));
 sg13g2_a22oi_1 _9090_ (.Y(_3097_),
    .B1(_3096_),
    .B2(net84),
    .A2(_3095_),
    .A1(net85));
 sg13g2_a21oi_1 _9091_ (.A1(_3094_),
    .A2(_3097_),
    .Y(_3098_),
    .B1(net66));
 sg13g2_mux4_1 _9092_ (.S0(net136),
    .A0(\logix.ram_r[162] ),
    .A1(\logix.ram_r[170] ),
    .A2(\logix.ram_r[178] ),
    .A3(\logix.ram_r[186] ),
    .S1(net101),
    .X(_3099_));
 sg13g2_mux4_1 _9093_ (.S0(net106),
    .A0(\logix.ram_r[130] ),
    .A1(\logix.ram_r[138] ),
    .A2(\logix.ram_r[146] ),
    .A3(\logix.ram_r[154] ),
    .S1(net112),
    .X(_3100_));
 sg13g2_a22oi_1 _9094_ (.Y(_3101_),
    .B1(_3100_),
    .B2(net30),
    .A2(_3099_),
    .A1(net31));
 sg13g2_mux4_1 _9095_ (.S0(net87),
    .A0(\logix.ram_r[226] ),
    .A1(\logix.ram_r[234] ),
    .A2(\logix.ram_r[242] ),
    .A3(\logix.ram_r[250] ),
    .S1(net86),
    .X(_3102_));
 sg13g2_mux4_1 _9096_ (.S0(net115),
    .A0(\logix.ram_r[194] ),
    .A1(\logix.ram_r[202] ),
    .A2(\logix.ram_r[210] ),
    .A3(\logix.ram_r[218] ),
    .S1(net102),
    .X(_3103_));
 sg13g2_a22oi_1 _9097_ (.Y(_3104_),
    .B1(_3103_),
    .B2(net61),
    .A2(_3102_),
    .A1(net62));
 sg13g2_a21oi_1 _9098_ (.A1(_3101_),
    .A2(_3104_),
    .Y(_3105_),
    .B1(net67));
 sg13g2_or2_1 _9099_ (.X(_3106_),
    .B(_3105_),
    .A(_3098_));
 sg13g2_a221oi_1 _9100_ (.B2(_3091_),
    .C1(_3106_),
    .B1(_3090_),
    .A1(_3072_),
    .Y(_3107_),
    .A2(_3079_));
 sg13g2_nor4_2 _9101_ (.A(_2970_),
    .B(_3022_),
    .C(_3067_),
    .Y(net16),
    .D(_3107_));
 sg13g2_nand2b_1 _9102_ (.Y(_3108_),
    .B(net127),
    .A_N(\logix.ram_r[1875] ));
 sg13g2_o21ai_1 _9103_ (.B1(_3108_),
    .Y(_3109_),
    .A1(\logix.ram_r[1859] ),
    .A2(net60));
 sg13g2_nand2b_1 _9104_ (.Y(_3110_),
    .B(net64),
    .A_N(\logix.ram_r[1883] ));
 sg13g2_o21ai_1 _9105_ (.B1(_3110_),
    .Y(_3111_),
    .A1(\logix.ram_r[1867] ),
    .A2(net53));
 sg13g2_a221oi_1 _9106_ (.B2(net28),
    .C1(_2709_),
    .B1(_3111_),
    .A1(net29),
    .Y(_3112_),
    .A2(_3109_));
 sg13g2_mux4_1 _9107_ (.S0(net164),
    .A0(\logix.ram_r[1827] ),
    .A1(\logix.ram_r[1835] ),
    .A2(\logix.ram_r[1843] ),
    .A3(\logix.ram_r[1851] ),
    .S1(net113),
    .X(_3113_));
 sg13g2_mux4_1 _9108_ (.S0(net195),
    .A0(\logix.ram_r[1795] ),
    .A1(\logix.ram_r[1803] ),
    .A2(\logix.ram_r[1811] ),
    .A3(\logix.ram_r[1819] ),
    .S1(net192),
    .X(_3114_));
 sg13g2_and2_1 _9109_ (.A(_2458_),
    .B(_3114_),
    .X(_3115_));
 sg13g2_a221oi_1 _9110_ (.B2(net90),
    .C1(_3115_),
    .B1(_3113_),
    .A1(net206),
    .Y(_3116_),
    .A2(net205));
 sg13g2_mux4_1 _9111_ (.S0(net52),
    .A0(\logix.ram_r[1891] ),
    .A1(\logix.ram_r[1899] ),
    .A2(\logix.ram_r[1907] ),
    .A3(\logix.ram_r[1915] ),
    .S1(net59),
    .X(_3117_));
 sg13g2_nor2_1 _9112_ (.A(net89),
    .B(_3117_),
    .Y(_3118_));
 sg13g2_nor2_1 _9113_ (.A(_3116_),
    .B(_3118_),
    .Y(_3119_));
 sg13g2_mux4_1 _9114_ (.S0(net180),
    .A0(\logix.ram_r[1923] ),
    .A1(\logix.ram_r[1931] ),
    .A2(\logix.ram_r[1939] ),
    .A3(\logix.ram_r[1947] ),
    .S1(net181),
    .X(_3120_));
 sg13g2_mux4_1 _9115_ (.S0(net203),
    .A0(\logix.ram_r[1955] ),
    .A1(\logix.ram_r[1963] ),
    .A2(\logix.ram_r[1971] ),
    .A3(\logix.ram_r[1979] ),
    .S1(net193),
    .X(_3121_));
 sg13g2_mux2_1 _9116_ (.A0(_3120_),
    .A1(_3121_),
    .S(net194),
    .X(_3122_));
 sg13g2_nand2_1 _9117_ (.Y(_3123_),
    .A(net174),
    .B(_3122_));
 sg13g2_mux2_1 _9118_ (.A0(\logix.ram_r[1987] ),
    .A1(\logix.ram_r[1995] ),
    .S(net52),
    .X(_3124_));
 sg13g2_mux2_1 _9119_ (.A0(\logix.ram_r[2035] ),
    .A1(\logix.ram_r[2043] ),
    .S(net51),
    .X(_3125_));
 sg13g2_a22oi_1 _9120_ (.Y(_3126_),
    .B1(_3125_),
    .B2(net45),
    .A2(_3124_),
    .A1(net46));
 sg13g2_mux2_1 _9121_ (.A0(\logix.ram_r[2019] ),
    .A1(\logix.ram_r[2027] ),
    .S(net52),
    .X(_3127_));
 sg13g2_mux2_1 _9122_ (.A0(\logix.ram_r[2003] ),
    .A1(\logix.ram_r[2011] ),
    .S(net51),
    .X(_3128_));
 sg13g2_a22oi_1 _9123_ (.Y(_3129_),
    .B1(_3128_),
    .B2(net47),
    .A2(_3127_),
    .A1(net48));
 sg13g2_nand4_1 _9124_ (.B(_3123_),
    .C(_3126_),
    .A(_2780_),
    .Y(_3130_),
    .D(_3129_));
 sg13g2_mux4_1 _9125_ (.S0(net196),
    .A0(\logix.ram_r[1571] ),
    .A1(\logix.ram_r[1579] ),
    .A2(\logix.ram_r[1587] ),
    .A3(\logix.ram_r[1595] ),
    .S1(net181),
    .X(_3131_));
 sg13g2_mux4_1 _9126_ (.S0(net183),
    .A0(\logix.ram_r[1539] ),
    .A1(\logix.ram_r[1547] ),
    .A2(\logix.ram_r[1555] ),
    .A3(\logix.ram_r[1563] ),
    .S1(net108),
    .X(_3132_));
 sg13g2_a22oi_1 _9127_ (.Y(_3133_),
    .B1(_3132_),
    .B2(net55),
    .A2(_3131_),
    .A1(net56));
 sg13g2_mux4_1 _9128_ (.S0(net203),
    .A0(\logix.ram_r[1635] ),
    .A1(\logix.ram_r[1643] ),
    .A2(\logix.ram_r[1651] ),
    .A3(\logix.ram_r[1659] ),
    .S1(net193),
    .X(_3134_));
 sg13g2_mux4_1 _9129_ (.S0(net185),
    .A0(\logix.ram_r[1603] ),
    .A1(\logix.ram_r[1611] ),
    .A2(\logix.ram_r[1619] ),
    .A3(\logix.ram_r[1627] ),
    .S1(net93),
    .X(_3135_));
 sg13g2_a22oi_1 _9130_ (.Y(_3136_),
    .B1(_3135_),
    .B2(net91),
    .A2(_3134_),
    .A1(net126));
 sg13g2_a21oi_1 _9131_ (.A1(_3133_),
    .A2(_3136_),
    .Y(_3137_),
    .B1(net54));
 sg13g2_mux4_1 _9132_ (.S0(net201),
    .A0(\logix.ram_r[1699] ),
    .A1(\logix.ram_r[1707] ),
    .A2(\logix.ram_r[1715] ),
    .A3(\logix.ram_r[1723] ),
    .S1(net197),
    .X(_3138_));
 sg13g2_mux4_1 _9133_ (.S0(net88),
    .A0(\logix.ram_r[1667] ),
    .A1(\logix.ram_r[1675] ),
    .A2(\logix.ram_r[1683] ),
    .A3(\logix.ram_r[1691] ),
    .S1(net108),
    .X(_3139_));
 sg13g2_a22oi_1 _9134_ (.Y(_3140_),
    .B1(_3139_),
    .B2(net55),
    .A2(_3138_),
    .A1(net56));
 sg13g2_mux4_1 _9135_ (.S0(net180),
    .A0(\logix.ram_r[1763] ),
    .A1(\logix.ram_r[1771] ),
    .A2(\logix.ram_r[1779] ),
    .A3(\logix.ram_r[1787] ),
    .S1(net184),
    .X(_3141_));
 sg13g2_mux4_1 _9136_ (.S0(net183),
    .A0(\logix.ram_r[1731] ),
    .A1(\logix.ram_r[1739] ),
    .A2(\logix.ram_r[1747] ),
    .A3(\logix.ram_r[1755] ),
    .S1(net99),
    .X(_3142_));
 sg13g2_a22oi_1 _9137_ (.Y(_3143_),
    .B1(_3142_),
    .B2(net91),
    .A2(_3141_),
    .A1(net126));
 sg13g2_a21oi_1 _9138_ (.A1(_3140_),
    .A2(_3143_),
    .Y(_3144_),
    .B1(net50));
 sg13g2_or2_1 _9139_ (.X(_3145_),
    .B(_3144_),
    .A(_3137_));
 sg13g2_a221oi_1 _9140_ (.B2(_3047_),
    .C1(_3145_),
    .B1(_3130_),
    .A1(_3112_),
    .Y(_3146_),
    .A2(_3119_));
 sg13g2_nand2b_1 _9141_ (.Y(_3147_),
    .B(_2451_),
    .A_N(_2454_));
 sg13g2_mux4_1 _9142_ (.S0(net191),
    .A0(\logix.ram_r[899] ),
    .A1(\logix.ram_r[907] ),
    .A2(\logix.ram_r[915] ),
    .A3(\logix.ram_r[923] ),
    .S1(net190),
    .X(_3148_));
 sg13g2_mux4_1 _9143_ (.S0(net191),
    .A0(\logix.ram_r[931] ),
    .A1(\logix.ram_r[939] ),
    .A2(\logix.ram_r[947] ),
    .A3(\logix.ram_r[955] ),
    .S1(net190),
    .X(_3149_));
 sg13g2_mux2_1 _9144_ (.A0(_3148_),
    .A1(_3149_),
    .S(net204),
    .X(_3150_));
 sg13g2_mux2_1 _9145_ (.A0(\logix.ram_r[963] ),
    .A1(\logix.ram_r[971] ),
    .S(net198),
    .X(_3151_));
 sg13g2_nand3_1 _9146_ (.B(_2480_),
    .C(_3151_),
    .A(net207),
    .Y(_3152_));
 sg13g2_mux2_1 _9147_ (.A0(\logix.ram_r[1011] ),
    .A1(\logix.ram_r[1019] ),
    .S(net198),
    .X(_3153_));
 sg13g2_nand3_1 _9148_ (.B(net158),
    .C(_3153_),
    .A(net162),
    .Y(_3154_));
 sg13g2_mux2_1 _9149_ (.A0(\logix.ram_r[995] ),
    .A1(\logix.ram_r[1003] ),
    .S(net198),
    .X(_3155_));
 sg13g2_nand3_1 _9150_ (.B(net158),
    .C(_3155_),
    .A(net207),
    .Y(_3156_));
 sg13g2_mux2_1 _9151_ (.A0(\logix.ram_r[979] ),
    .A1(\logix.ram_r[987] ),
    .S(net198),
    .X(_3157_));
 sg13g2_nand3_1 _9152_ (.B(_2480_),
    .C(_3157_),
    .A(net153),
    .Y(_3158_));
 sg13g2_nand4_1 _9153_ (.B(_3154_),
    .C(_3156_),
    .A(_3152_),
    .Y(_3159_),
    .D(_3158_));
 sg13g2_a21oi_1 _9154_ (.A1(net174),
    .A2(_3150_),
    .Y(_3160_),
    .B1(_3159_));
 sg13g2_mux4_1 _9155_ (.S0(net195),
    .A0(\logix.ram_r[547] ),
    .A1(\logix.ram_r[555] ),
    .A2(\logix.ram_r[563] ),
    .A3(\logix.ram_r[571] ),
    .S1(net192),
    .X(_3161_));
 sg13g2_mux4_1 _9156_ (.S0(net196),
    .A0(\logix.ram_r[515] ),
    .A1(\logix.ram_r[523] ),
    .A2(\logix.ram_r[531] ),
    .A3(\logix.ram_r[539] ),
    .S1(net189),
    .X(_3162_));
 sg13g2_a22oi_1 _9157_ (.Y(_3163_),
    .B1(_3162_),
    .B2(net77),
    .A2(_3161_),
    .A1(net78));
 sg13g2_mux4_1 _9158_ (.S0(net191),
    .A0(\logix.ram_r[611] ),
    .A1(\logix.ram_r[619] ),
    .A2(\logix.ram_r[627] ),
    .A3(\logix.ram_r[635] ),
    .S1(_2642_),
    .X(_3164_));
 sg13g2_mux4_1 _9159_ (.S0(net203),
    .A0(\logix.ram_r[579] ),
    .A1(\logix.ram_r[587] ),
    .A2(\logix.ram_r[595] ),
    .A3(\logix.ram_r[603] ),
    .S1(net184),
    .X(_3165_));
 sg13g2_a22oi_1 _9160_ (.Y(_3166_),
    .B1(_3165_),
    .B2(net154),
    .A2(_3164_),
    .A1(_2472_));
 sg13g2_a21o_1 _9161_ (.A2(_3166_),
    .A1(_3163_),
    .B1(_2485_),
    .X(_3167_));
 sg13g2_o21ai_1 _9162_ (.B1(_3167_),
    .Y(_3168_),
    .A1(_2603_),
    .A2(_3160_));
 sg13g2_mux4_1 _9163_ (.S0(net171),
    .A0(\logix.ram_r[675] ),
    .A1(\logix.ram_r[683] ),
    .A2(\logix.ram_r[691] ),
    .A3(\logix.ram_r[699] ),
    .S1(net110),
    .X(_3169_));
 sg13g2_mux4_1 _9164_ (.S0(net172),
    .A0(\logix.ram_r[643] ),
    .A1(\logix.ram_r[651] ),
    .A2(\logix.ram_r[659] ),
    .A3(\logix.ram_r[667] ),
    .S1(net127),
    .X(_3170_));
 sg13g2_a22oi_1 _9165_ (.Y(_3171_),
    .B1(_3170_),
    .B2(net38),
    .A2(_3169_),
    .A1(net39));
 sg13g2_mux4_1 _9166_ (.S0(net125),
    .A0(\logix.ram_r[739] ),
    .A1(\logix.ram_r[747] ),
    .A2(\logix.ram_r[755] ),
    .A3(\logix.ram_r[763] ),
    .S1(_2597_),
    .X(_3172_));
 sg13g2_mux4_1 _9167_ (.S0(_2524_),
    .A0(\logix.ram_r[707] ),
    .A1(\logix.ram_r[715] ),
    .A2(\logix.ram_r[723] ),
    .A3(\logix.ram_r[731] ),
    .S1(_2590_),
    .X(_3173_));
 sg13g2_a22oi_1 _9168_ (.Y(_3174_),
    .B1(_3173_),
    .B2(net72),
    .A2(_3172_),
    .A1(_2594_));
 sg13g2_a21oi_1 _9169_ (.A1(_3171_),
    .A2(_3174_),
    .Y(_3175_),
    .B1(net71));
 sg13g2_mux4_1 _9170_ (.S0(_2702_),
    .A0(\logix.ram_r[803] ),
    .A1(\logix.ram_r[811] ),
    .A2(\logix.ram_r[819] ),
    .A3(\logix.ram_r[827] ),
    .S1(_2650_),
    .X(_3176_));
 sg13g2_mux4_1 _9171_ (.S0(_2992_),
    .A0(\logix.ram_r[771] ),
    .A1(\logix.ram_r[779] ),
    .A2(\logix.ram_r[787] ),
    .A3(\logix.ram_r[795] ),
    .S1(net184),
    .X(_3177_));
 sg13g2_and2_1 _9172_ (.A(_2458_),
    .B(_3177_),
    .X(_3178_));
 sg13g2_a221oi_1 _9173_ (.B2(net90),
    .C1(_3178_),
    .B1(_3176_),
    .A1(net206),
    .Y(_3179_),
    .A2(net205));
 sg13g2_nand2_1 _9174_ (.Y(_3180_),
    .A(\logix.ram_r[835] ),
    .B(net207));
 sg13g2_nand2_1 _9175_ (.Y(_3181_),
    .A(\logix.ram_r[851] ),
    .B(_2643_));
 sg13g2_nand3_1 _9176_ (.B(_3180_),
    .C(_3181_),
    .A(_2639_),
    .Y(_3182_));
 sg13g2_nand2_1 _9177_ (.Y(_3183_),
    .A(\logix.ram_r[843] ),
    .B(net207));
 sg13g2_nand2_1 _9178_ (.Y(_3184_),
    .A(\logix.ram_r[859] ),
    .B(_2643_));
 sg13g2_nand3_1 _9179_ (.B(_3183_),
    .C(_3184_),
    .A(_2647_),
    .Y(_3185_));
 sg13g2_nand3_1 _9180_ (.B(_3182_),
    .C(_3185_),
    .A(net79),
    .Y(_3186_));
 sg13g2_mux4_1 _9181_ (.S0(_3032_),
    .A0(\logix.ram_r[867] ),
    .A1(\logix.ram_r[875] ),
    .A2(\logix.ram_r[883] ),
    .A3(\logix.ram_r[891] ),
    .S1(net63),
    .X(_3187_));
 sg13g2_nor2_1 _9182_ (.A(net89),
    .B(_3187_),
    .Y(_3188_));
 sg13g2_nor3_1 _9183_ (.A(_3179_),
    .B(_3186_),
    .C(_3188_),
    .Y(_3189_));
 sg13g2_nor4_1 _9184_ (.A(_3147_),
    .B(_3168_),
    .C(_3175_),
    .D(_3189_),
    .Y(_3190_));
 sg13g2_nand2b_1 _9185_ (.Y(_3191_),
    .B(net64),
    .A_N(\logix.ram_r[1491] ));
 sg13g2_o21ai_1 _9186_ (.B1(_3191_),
    .Y(_3192_),
    .A1(\logix.ram_r[1475] ),
    .A2(net60));
 sg13g2_nand2b_1 _9187_ (.Y(_3193_),
    .B(net63),
    .A_N(\logix.ram_r[1499] ));
 sg13g2_o21ai_1 _9188_ (.B1(_3193_),
    .Y(_3194_),
    .A1(\logix.ram_r[1483] ),
    .A2(net53));
 sg13g2_a221oi_1 _9189_ (.B2(net28),
    .C1(_2603_),
    .B1(_3194_),
    .A1(_2678_),
    .Y(_3195_),
    .A2(_3192_));
 sg13g2_mux4_1 _9190_ (.S0(net107),
    .A0(\logix.ram_r[1443] ),
    .A1(\logix.ram_r[1451] ),
    .A2(\logix.ram_r[1459] ),
    .A3(\logix.ram_r[1467] ),
    .S1(net111),
    .X(_3196_));
 sg13g2_mux4_1 _9191_ (.S0(net180),
    .A0(\logix.ram_r[1411] ),
    .A1(\logix.ram_r[1419] ),
    .A2(\logix.ram_r[1427] ),
    .A3(\logix.ram_r[1435] ),
    .S1(_2990_),
    .X(_3197_));
 sg13g2_and2_1 _9192_ (.A(net95),
    .B(_3197_),
    .X(_3198_));
 sg13g2_a221oi_1 _9193_ (.B2(net90),
    .C1(_3198_),
    .B1(_3196_),
    .A1(net206),
    .Y(_3199_),
    .A2(net205));
 sg13g2_mux4_1 _9194_ (.S0(net49),
    .A0(\logix.ram_r[1507] ),
    .A1(\logix.ram_r[1515] ),
    .A2(\logix.ram_r[1523] ),
    .A3(\logix.ram_r[1531] ),
    .S1(_2900_),
    .X(_3200_));
 sg13g2_nor2_1 _9195_ (.A(net89),
    .B(_3200_),
    .Y(_3201_));
 sg13g2_nor2_1 _9196_ (.A(_3199_),
    .B(_3201_),
    .Y(_3202_));
 sg13g2_mux4_1 _9197_ (.S0(net182),
    .A0(\logix.ram_r[1283] ),
    .A1(\logix.ram_r[1291] ),
    .A2(\logix.ram_r[1299] ),
    .A3(\logix.ram_r[1307] ),
    .S1(net93),
    .X(_3203_));
 sg13g2_mux4_1 _9198_ (.S0(net182),
    .A0(\logix.ram_r[1315] ),
    .A1(\logix.ram_r[1323] ),
    .A2(\logix.ram_r[1331] ),
    .A3(\logix.ram_r[1339] ),
    .S1(net92),
    .X(_3204_));
 sg13g2_mux2_1 _9199_ (.A0(_3203_),
    .A1(_3204_),
    .S(net199),
    .X(_3205_));
 sg13g2_nand2_1 _9200_ (.Y(_3206_),
    .A(net118),
    .B(_3205_));
 sg13g2_mux2_1 _9201_ (.A0(\logix.ram_r[1347] ),
    .A1(\logix.ram_r[1355] ),
    .S(net49),
    .X(_3207_));
 sg13g2_mux2_1 _9202_ (.A0(\logix.ram_r[1395] ),
    .A1(\logix.ram_r[1403] ),
    .S(net80),
    .X(_3208_));
 sg13g2_a22oi_1 _9203_ (.Y(_3209_),
    .B1(_3208_),
    .B2(net45),
    .A2(_3207_),
    .A1(net46));
 sg13g2_mux2_1 _9204_ (.A0(\logix.ram_r[1379] ),
    .A1(\logix.ram_r[1387] ),
    .S(net49),
    .X(_3210_));
 sg13g2_mux2_1 _9205_ (.A0(\logix.ram_r[1363] ),
    .A1(\logix.ram_r[1371] ),
    .S(net80),
    .X(_3211_));
 sg13g2_a22oi_1 _9206_ (.Y(_3212_),
    .B1(_3211_),
    .B2(net47),
    .A2(_3210_),
    .A1(net48));
 sg13g2_nand4_1 _9207_ (.B(_3206_),
    .C(_3209_),
    .A(_2706_),
    .Y(_3213_),
    .D(_3212_));
 sg13g2_mux4_1 _9208_ (.S0(net185),
    .A0(\logix.ram_r[1187] ),
    .A1(\logix.ram_r[1195] ),
    .A2(\logix.ram_r[1203] ),
    .A3(\logix.ram_r[1211] ),
    .S1(net175),
    .X(_3214_));
 sg13g2_mux4_1 _9209_ (.S0(net136),
    .A0(\logix.ram_r[1155] ),
    .A1(\logix.ram_r[1163] ),
    .A2(\logix.ram_r[1171] ),
    .A3(\logix.ram_r[1179] ),
    .S1(net101),
    .X(_3215_));
 sg13g2_a22oi_1 _9210_ (.Y(_3216_),
    .B1(_3215_),
    .B2(net55),
    .A2(_3214_),
    .A1(net56));
 sg13g2_mux4_1 _9211_ (.S0(net201),
    .A0(\logix.ram_r[1251] ),
    .A1(\logix.ram_r[1259] ),
    .A2(\logix.ram_r[1267] ),
    .A3(\logix.ram_r[1275] ),
    .S1(_2516_),
    .X(_3217_));
 sg13g2_mux4_1 _9212_ (.S0(_3013_),
    .A0(\logix.ram_r[1219] ),
    .A1(\logix.ram_r[1227] ),
    .A2(\logix.ram_r[1235] ),
    .A3(\logix.ram_r[1243] ),
    .S1(_3014_),
    .X(_3218_));
 sg13g2_a22oi_1 _9213_ (.Y(_3219_),
    .B1(_3218_),
    .B2(net91),
    .A2(_3217_),
    .A1(net85));
 sg13g2_a21oi_1 _9214_ (.A1(_3216_),
    .A2(_3219_),
    .Y(_3220_),
    .B1(_3010_));
 sg13g2_mux4_1 _9215_ (.S0(_2957_),
    .A0(\logix.ram_r[1059] ),
    .A1(\logix.ram_r[1067] ),
    .A2(\logix.ram_r[1075] ),
    .A3(\logix.ram_r[1083] ),
    .S1(_2785_),
    .X(_3221_));
 sg13g2_mux4_1 _9216_ (.S0(net100),
    .A0(\logix.ram_r[1027] ),
    .A1(\logix.ram_r[1035] ),
    .A2(\logix.ram_r[1043] ),
    .A3(\logix.ram_r[1051] ),
    .S1(net176),
    .X(_3222_));
 sg13g2_a22oi_1 _9217_ (.Y(_3223_),
    .B1(_3222_),
    .B2(net22),
    .A2(_3221_),
    .A1(net23));
 sg13g2_mux4_1 _9218_ (.S0(_2962_),
    .A0(\logix.ram_r[1123] ),
    .A1(\logix.ram_r[1131] ),
    .A2(\logix.ram_r[1139] ),
    .A3(\logix.ram_r[1147] ),
    .S1(net93),
    .X(_3224_));
 sg13g2_mux4_1 _9219_ (.S0(_2910_),
    .A0(\logix.ram_r[1091] ),
    .A1(\logix.ram_r[1099] ),
    .A2(\logix.ram_r[1107] ),
    .A3(\logix.ram_r[1115] ),
    .S1(net147),
    .X(_3225_));
 sg13g2_a22oi_1 _9220_ (.Y(_3226_),
    .B1(_3225_),
    .B2(_3056_),
    .A2(_3224_),
    .A1(net85));
 sg13g2_a21oi_1 _9221_ (.A1(_3223_),
    .A2(_3226_),
    .Y(_3227_),
    .B1(net54));
 sg13g2_or2_1 _9222_ (.X(_3228_),
    .B(_3227_),
    .A(_3220_));
 sg13g2_a221oi_1 _9223_ (.B2(_2710_),
    .C1(_3228_),
    .B1(_3213_),
    .A1(_3195_),
    .Y(_3229_),
    .A2(_3202_));
 sg13g2_nand2b_1 _9224_ (.Y(_3230_),
    .B(net58),
    .A_N(\logix.ram_r[339] ));
 sg13g2_o21ai_1 _9225_ (.B1(_3230_),
    .Y(_3231_),
    .A1(\logix.ram_r[323] ),
    .A2(_2973_));
 sg13g2_nand2b_1 _9226_ (.Y(_3232_),
    .B(_2649_),
    .A_N(\logix.ram_r[347] ));
 sg13g2_o21ai_1 _9227_ (.B1(_3232_),
    .Y(_3233_),
    .A1(\logix.ram_r[331] ),
    .A2(_2973_));
 sg13g2_a221oi_1 _9228_ (.B2(_2684_),
    .C1(_2709_),
    .B1(_3233_),
    .A1(_2678_),
    .Y(_3234_),
    .A2(_3231_));
 sg13g2_mux4_1 _9229_ (.S0(_2521_),
    .A0(\logix.ram_r[291] ),
    .A1(\logix.ram_r[299] ),
    .A2(\logix.ram_r[307] ),
    .A3(\logix.ram_r[315] ),
    .S1(net124),
    .X(_3235_));
 sg13g2_mux4_1 _9230_ (.S0(net185),
    .A0(\logix.ram_r[259] ),
    .A1(\logix.ram_r[267] ),
    .A2(\logix.ram_r[275] ),
    .A3(\logix.ram_r[283] ),
    .S1(_2938_),
    .X(_3236_));
 sg13g2_and2_1 _9231_ (.A(_2879_),
    .B(_3236_),
    .X(_3237_));
 sg13g2_a221oi_1 _9232_ (.B2(_2980_),
    .C1(_3237_),
    .B1(_3235_),
    .A1(_2977_),
    .Y(_3238_),
    .A2(_2978_));
 sg13g2_mux4_1 _9233_ (.S0(_2997_),
    .A0(\logix.ram_r[355] ),
    .A1(\logix.ram_r[363] ),
    .A2(\logix.ram_r[371] ),
    .A3(\logix.ram_r[379] ),
    .S1(_2649_),
    .X(_3239_));
 sg13g2_nor2_1 _9234_ (.A(_2984_),
    .B(_3239_),
    .Y(_3240_));
 sg13g2_nor2_1 _9235_ (.A(_3238_),
    .B(_3240_),
    .Y(_3241_));
 sg13g2_mux4_1 _9236_ (.S0(net109),
    .A0(\logix.ram_r[387] ),
    .A1(\logix.ram_r[395] ),
    .A2(\logix.ram_r[403] ),
    .A3(\logix.ram_r[411] ),
    .S1(net104),
    .X(_3242_));
 sg13g2_mux4_1 _9237_ (.S0(net88),
    .A0(\logix.ram_r[419] ),
    .A1(\logix.ram_r[427] ),
    .A2(\logix.ram_r[435] ),
    .A3(\logix.ram_r[443] ),
    .S1(net97),
    .X(_3243_));
 sg13g2_mux2_1 _9238_ (.A0(_3242_),
    .A1(_3243_),
    .S(net188),
    .X(_3244_));
 sg13g2_nand2_1 _9239_ (.Y(_3245_),
    .A(net118),
    .B(_3244_));
 sg13g2_mux2_1 _9240_ (.A0(\logix.ram_r[451] ),
    .A1(\logix.ram_r[459] ),
    .S(net80),
    .X(_3246_));
 sg13g2_mux2_1 _9241_ (.A0(\logix.ram_r[499] ),
    .A1(\logix.ram_r[507] ),
    .S(net57),
    .X(_3247_));
 sg13g2_a22oi_1 _9242_ (.Y(_3248_),
    .B1(_3247_),
    .B2(_2396_),
    .A2(_3246_),
    .A1(_2390_));
 sg13g2_mux2_1 _9243_ (.A0(\logix.ram_r[483] ),
    .A1(\logix.ram_r[491] ),
    .S(net51),
    .X(_3249_));
 sg13g2_mux2_1 _9244_ (.A0(\logix.ram_r[467] ),
    .A1(\logix.ram_r[475] ),
    .S(net57),
    .X(_3250_));
 sg13g2_a22oi_1 _9245_ (.Y(_3251_),
    .B1(_3250_),
    .B2(net47),
    .A2(_3249_),
    .A1(_2373_));
 sg13g2_nand4_1 _9246_ (.B(_3245_),
    .C(_3248_),
    .A(_2456_),
    .Y(_3252_),
    .D(_3251_));
 sg13g2_mux4_1 _9247_ (.S0(net109),
    .A0(\logix.ram_r[35] ),
    .A1(\logix.ram_r[43] ),
    .A2(\logix.ram_r[51] ),
    .A3(\logix.ram_r[59] ),
    .S1(_2512_),
    .X(_3253_));
 sg13g2_mux4_1 _9248_ (.S0(net149),
    .A0(\logix.ram_r[3] ),
    .A1(\logix.ram_r[11] ),
    .A2(\logix.ram_r[19] ),
    .A3(\logix.ram_r[27] ),
    .S1(net148),
    .X(_3254_));
 sg13g2_a22oi_1 _9249_ (.Y(_3255_),
    .B1(_3254_),
    .B2(_3051_),
    .A2(_3253_),
    .A1(_3048_));
 sg13g2_mux4_1 _9250_ (.S0(net88),
    .A0(\logix.ram_r[99] ),
    .A1(\logix.ram_r[107] ),
    .A2(\logix.ram_r[115] ),
    .A3(\logix.ram_r[123] ),
    .S1(net108),
    .X(_3256_));
 sg13g2_mux4_1 _9251_ (.S0(net139),
    .A0(\logix.ram_r[67] ),
    .A1(\logix.ram_r[75] ),
    .A2(\logix.ram_r[83] ),
    .A3(\logix.ram_r[91] ),
    .S1(net138),
    .X(_3257_));
 sg13g2_a22oi_1 _9252_ (.Y(_3258_),
    .B1(_3257_),
    .B2(_3056_),
    .A2(_3256_),
    .A1(_3053_));
 sg13g2_a21oi_1 _9253_ (.A1(_3255_),
    .A2(_3258_),
    .Y(_3259_),
    .B1(net54));
 sg13g2_mux4_1 _9254_ (.S0(net136),
    .A0(\logix.ram_r[163] ),
    .A1(\logix.ram_r[171] ),
    .A2(\logix.ram_r[179] ),
    .A3(\logix.ram_r[187] ),
    .S1(net101),
    .X(_3260_));
 sg13g2_mux4_1 _9255_ (.S0(net106),
    .A0(\logix.ram_r[131] ),
    .A1(\logix.ram_r[139] ),
    .A2(\logix.ram_r[147] ),
    .A3(\logix.ram_r[155] ),
    .S1(net112),
    .X(_3261_));
 sg13g2_a22oi_1 _9256_ (.Y(_3262_),
    .B1(_3261_),
    .B2(net22),
    .A2(_3260_),
    .A1(net23));
 sg13g2_mux4_1 _9257_ (.S0(net87),
    .A0(\logix.ram_r[227] ),
    .A1(\logix.ram_r[235] ),
    .A2(\logix.ram_r[243] ),
    .A3(\logix.ram_r[251] ),
    .S1(net86),
    .X(_3263_));
 sg13g2_mux4_1 _9258_ (.S0(net157),
    .A0(\logix.ram_r[195] ),
    .A1(\logix.ram_r[203] ),
    .A2(\logix.ram_r[211] ),
    .A3(\logix.ram_r[219] ),
    .S1(net102),
    .X(_3264_));
 sg13g2_a22oi_1 _9259_ (.Y(_3265_),
    .B1(_3264_),
    .B2(net84),
    .A2(_3263_),
    .A1(net62));
 sg13g2_a21oi_1 _9260_ (.A1(_3262_),
    .A2(_3265_),
    .Y(_3266_),
    .B1(net50));
 sg13g2_or2_1 _9261_ (.X(_3267_),
    .B(_3266_),
    .A(_3259_));
 sg13g2_a221oi_1 _9262_ (.B2(_3091_),
    .C1(_3267_),
    .B1(_3252_),
    .A1(_3234_),
    .Y(_3268_),
    .A2(_3241_));
 sg13g2_nor4_2 _9263_ (.A(_3146_),
    .B(_3190_),
    .C(_3229_),
    .Y(net17),
    .D(_3268_));
 sg13g2_mux4_1 _9264_ (.S0(net195),
    .A0(\logix.ram_r[388] ),
    .A1(\logix.ram_r[396] ),
    .A2(\logix.ram_r[404] ),
    .A3(\logix.ram_r[412] ),
    .S1(net192),
    .X(_3269_));
 sg13g2_nor2_1 _9265_ (.A(net199),
    .B(_3269_),
    .Y(_3270_));
 sg13g2_mux2_1 _9266_ (.A0(\logix.ram_r[420] ),
    .A1(\logix.ram_r[436] ),
    .S(net190),
    .X(_3271_));
 sg13g2_nor2_1 _9267_ (.A(_2344_),
    .B(_3271_),
    .Y(_3272_));
 sg13g2_mux2_1 _9268_ (.A0(\logix.ram_r[428] ),
    .A1(\logix.ram_r[444] ),
    .S(_2426_),
    .X(_3273_));
 sg13g2_o21ai_1 _9269_ (.B1(_2362_),
    .Y(_3274_),
    .A1(_2352_),
    .A2(_3273_));
 sg13g2_nor3_1 _9270_ (.A(_3270_),
    .B(_3272_),
    .C(_3274_),
    .Y(_3275_));
 sg13g2_mux2_1 _9271_ (.A0(\logix.ram_r[484] ),
    .A1(\logix.ram_r[492] ),
    .S(net133),
    .X(_3276_));
 sg13g2_mux2_1 _9272_ (.A0(\logix.ram_r[468] ),
    .A1(\logix.ram_r[476] ),
    .S(net164),
    .X(_3277_));
 sg13g2_a22oi_1 _9273_ (.Y(_3278_),
    .B1(_3277_),
    .B2(net32),
    .A2(_3276_),
    .A1(net33));
 sg13g2_mux2_1 _9274_ (.A0(\logix.ram_r[452] ),
    .A1(\logix.ram_r[460] ),
    .S(net166),
    .X(_3279_));
 sg13g2_mux2_1 _9275_ (.A0(\logix.ram_r[500] ),
    .A1(\logix.ram_r[508] ),
    .S(net164),
    .X(_3280_));
 sg13g2_a22oi_1 _9276_ (.Y(_3281_),
    .B1(_3280_),
    .B2(_2700_),
    .A2(_3279_),
    .A1(_2696_));
 sg13g2_nand2_1 _9277_ (.Y(_3282_),
    .A(_3278_),
    .B(_3281_));
 sg13g2_o21ai_1 _9278_ (.B1(net170),
    .Y(_3283_),
    .A1(_3275_),
    .A2(_3282_));
 sg13g2_mux4_1 _9279_ (.S0(_2596_),
    .A0(\logix.ram_r[260] ),
    .A1(\logix.ram_r[276] ),
    .A2(\logix.ram_r[292] ),
    .A3(\logix.ram_r[308] ),
    .S1(net204),
    .X(_3284_));
 sg13g2_mux4_1 _9280_ (.S0(_2596_),
    .A0(\logix.ram_r[268] ),
    .A1(\logix.ram_r[284] ),
    .A2(\logix.ram_r[300] ),
    .A3(\logix.ram_r[316] ),
    .S1(_2325_),
    .X(_3285_));
 sg13g2_mux2_1 _9281_ (.A0(_3284_),
    .A1(_3285_),
    .S(net57),
    .X(_3286_));
 sg13g2_mux4_1 _9282_ (.S0(_2937_),
    .A0(\logix.ram_r[324] ),
    .A1(\logix.ram_r[332] ),
    .A2(\logix.ram_r[340] ),
    .A3(\logix.ram_r[348] ),
    .S1(_2938_),
    .X(_3287_));
 sg13g2_nor2_1 _9283_ (.A(net202),
    .B(_3287_),
    .Y(_3288_));
 sg13g2_mux2_1 _9284_ (.A0(\logix.ram_r[364] ),
    .A1(\logix.ram_r[380] ),
    .S(net184),
    .X(_3289_));
 sg13g2_nor2_1 _9285_ (.A(_2433_),
    .B(_3289_),
    .Y(_3290_));
 sg13g2_mux2_1 _9286_ (.A0(\logix.ram_r[356] ),
    .A1(\logix.ram_r[372] ),
    .S(_2642_),
    .X(_3291_));
 sg13g2_o21ai_1 _9287_ (.B1(_2444_),
    .Y(_3292_),
    .A1(_2439_),
    .A2(_3291_));
 sg13g2_nor3_1 _9288_ (.A(_3288_),
    .B(_3290_),
    .C(_3292_),
    .Y(_3293_));
 sg13g2_o21ai_1 _9289_ (.B1(_3293_),
    .Y(_3294_),
    .A1(_2612_),
    .A2(_3286_));
 sg13g2_mux4_1 _9290_ (.S0(net200),
    .A0(\logix.ram_r[164] ),
    .A1(\logix.ram_r[172] ),
    .A2(\logix.ram_r[180] ),
    .A3(\logix.ram_r[188] ),
    .S1(net186),
    .X(_3295_));
 sg13g2_mux4_1 _9291_ (.S0(net201),
    .A0(\logix.ram_r[132] ),
    .A1(\logix.ram_r[140] ),
    .A2(\logix.ram_r[148] ),
    .A3(\logix.ram_r[156] ),
    .S1(net197),
    .X(_3296_));
 sg13g2_a22oi_1 _9292_ (.Y(_3297_),
    .B1(_3296_),
    .B2(net77),
    .A2(_3295_),
    .A1(net78));
 sg13g2_mux4_1 _9293_ (.S0(net195),
    .A0(\logix.ram_r[228] ),
    .A1(\logix.ram_r[236] ),
    .A2(\logix.ram_r[244] ),
    .A3(\logix.ram_r[252] ),
    .S1(net192),
    .X(_3298_));
 sg13g2_mux4_1 _9294_ (.S0(net196),
    .A0(\logix.ram_r[196] ),
    .A1(\logix.ram_r[204] ),
    .A2(\logix.ram_r[212] ),
    .A3(\logix.ram_r[220] ),
    .S1(net189),
    .X(_3299_));
 sg13g2_a22oi_1 _9295_ (.Y(_3300_),
    .B1(_3299_),
    .B2(net154),
    .A2(_3298_),
    .A1(net158));
 sg13g2_a21oi_1 _9296_ (.A1(_3297_),
    .A2(_3300_),
    .Y(_3301_),
    .B1(_2502_));
 sg13g2_mux4_1 _9297_ (.S0(net203),
    .A0(\logix.ram_r[36] ),
    .A1(\logix.ram_r[44] ),
    .A2(\logix.ram_r[52] ),
    .A3(\logix.ram_r[60] ),
    .S1(_2941_),
    .X(_3302_));
 sg13g2_mux4_1 _9298_ (.S0(_2937_),
    .A0(\logix.ram_r[4] ),
    .A1(\logix.ram_r[12] ),
    .A2(\logix.ram_r[20] ),
    .A3(\logix.ram_r[28] ),
    .S1(net175),
    .X(_3303_));
 sg13g2_a22oi_1 _9299_ (.Y(_3304_),
    .B1(_3303_),
    .B2(net77),
    .A2(_3302_),
    .A1(net78));
 sg13g2_mux4_1 _9300_ (.S0(net200),
    .A0(\logix.ram_r[100] ),
    .A1(\logix.ram_r[108] ),
    .A2(\logix.ram_r[116] ),
    .A3(\logix.ram_r[124] ),
    .S1(net186),
    .X(_3305_));
 sg13g2_mux4_1 _9301_ (.S0(_2384_),
    .A0(\logix.ram_r[68] ),
    .A1(\logix.ram_r[76] ),
    .A2(\logix.ram_r[84] ),
    .A3(\logix.ram_r[92] ),
    .S1(net92),
    .X(_3306_));
 sg13g2_a22oi_1 _9302_ (.Y(_3307_),
    .B1(_3306_),
    .B2(net154),
    .A2(_3305_),
    .A1(net126));
 sg13g2_a21oi_1 _9303_ (.A1(_3304_),
    .A2(_3307_),
    .Y(_3308_),
    .B1(net54));
 sg13g2_nor2_1 _9304_ (.A(_3301_),
    .B(_3308_),
    .Y(_3309_));
 sg13g2_and4_1 _9305_ (.A(_2456_),
    .B(_3283_),
    .C(_3294_),
    .D(_3309_),
    .X(_3310_));
 sg13g2_nand2b_1 _9306_ (.Y(_3311_),
    .B(net59),
    .A_N(\logix.ram_r[1492] ));
 sg13g2_o21ai_1 _9307_ (.B1(_3311_),
    .Y(_3312_),
    .A1(\logix.ram_r[1476] ),
    .A2(net60));
 sg13g2_nand2b_1 _9308_ (.Y(_3313_),
    .B(net64),
    .A_N(\logix.ram_r[1500] ));
 sg13g2_o21ai_1 _9309_ (.B1(_3313_),
    .Y(_3314_),
    .A1(\logix.ram_r[1484] ),
    .A2(net53));
 sg13g2_a221oi_1 _9310_ (.B2(net28),
    .C1(_2603_),
    .B1(_3314_),
    .A1(net29),
    .Y(_3315_),
    .A2(_3312_));
 sg13g2_mux4_1 _9311_ (.S0(_2847_),
    .A0(\logix.ram_r[1444] ),
    .A1(\logix.ram_r[1452] ),
    .A2(\logix.ram_r[1460] ),
    .A3(\logix.ram_r[1468] ),
    .S1(net113),
    .X(_3316_));
 sg13g2_mux4_1 _9312_ (.S0(net200),
    .A0(\logix.ram_r[1412] ),
    .A1(\logix.ram_r[1420] ),
    .A2(\logix.ram_r[1428] ),
    .A3(\logix.ram_r[1436] ),
    .S1(_2917_),
    .X(_3317_));
 sg13g2_and2_1 _9313_ (.A(_2458_),
    .B(_3317_),
    .X(_3318_));
 sg13g2_a221oi_1 _9314_ (.B2(net90),
    .C1(_3318_),
    .B1(_3316_),
    .A1(net206),
    .Y(_3319_),
    .A2(net205));
 sg13g2_mux4_1 _9315_ (.S0(_2986_),
    .A0(\logix.ram_r[1508] ),
    .A1(\logix.ram_r[1516] ),
    .A2(\logix.ram_r[1524] ),
    .A3(\logix.ram_r[1532] ),
    .S1(net64),
    .X(_3320_));
 sg13g2_nor2_1 _9316_ (.A(net89),
    .B(_3320_),
    .Y(_3321_));
 sg13g2_nor2_1 _9317_ (.A(_3319_),
    .B(_3321_),
    .Y(_3322_));
 sg13g2_mux4_1 _9318_ (.S0(net196),
    .A0(\logix.ram_r[1284] ),
    .A1(\logix.ram_r[1292] ),
    .A2(\logix.ram_r[1300] ),
    .A3(\logix.ram_r[1308] ),
    .S1(net181),
    .X(_3323_));
 sg13g2_mux4_1 _9319_ (.S0(net180),
    .A0(\logix.ram_r[1316] ),
    .A1(\logix.ram_r[1324] ),
    .A2(\logix.ram_r[1332] ),
    .A3(\logix.ram_r[1340] ),
    .S1(net184),
    .X(_3324_));
 sg13g2_mux2_1 _9320_ (.A0(_3323_),
    .A1(_3324_),
    .S(net194),
    .X(_3325_));
 sg13g2_nand2_1 _9321_ (.Y(_3326_),
    .A(net118),
    .B(_3325_));
 sg13g2_mux2_1 _9322_ (.A0(\logix.ram_r[1348] ),
    .A1(\logix.ram_r[1356] ),
    .S(net52),
    .X(_3327_));
 sg13g2_mux2_1 _9323_ (.A0(\logix.ram_r[1396] ),
    .A1(\logix.ram_r[1404] ),
    .S(net51),
    .X(_3328_));
 sg13g2_a22oi_1 _9324_ (.Y(_3329_),
    .B1(_3328_),
    .B2(net45),
    .A2(_3327_),
    .A1(net46));
 sg13g2_mux2_1 _9325_ (.A0(\logix.ram_r[1380] ),
    .A1(\logix.ram_r[1388] ),
    .S(net52),
    .X(_3330_));
 sg13g2_mux2_1 _9326_ (.A0(\logix.ram_r[1364] ),
    .A1(\logix.ram_r[1372] ),
    .S(net51),
    .X(_3331_));
 sg13g2_a22oi_1 _9327_ (.Y(_3332_),
    .B1(_3331_),
    .B2(net47),
    .A2(_3330_),
    .A1(net48));
 sg13g2_nand4_1 _9328_ (.B(_3326_),
    .C(_3329_),
    .A(_2706_),
    .Y(_3333_),
    .D(_3332_));
 sg13g2_mux4_1 _9329_ (.S0(net196),
    .A0(\logix.ram_r[1188] ),
    .A1(\logix.ram_r[1196] ),
    .A2(\logix.ram_r[1204] ),
    .A3(\logix.ram_r[1212] ),
    .S1(_2736_),
    .X(_3334_));
 sg13g2_mux4_1 _9330_ (.S0(net88),
    .A0(\logix.ram_r[1156] ),
    .A1(\logix.ram_r[1164] ),
    .A2(\logix.ram_r[1172] ),
    .A3(\logix.ram_r[1180] ),
    .S1(net108),
    .X(_3335_));
 sg13g2_a22oi_1 _9331_ (.Y(_3336_),
    .B1(_3335_),
    .B2(net55),
    .A2(_3334_),
    .A1(net56));
 sg13g2_mux4_1 _9332_ (.S0(_2374_),
    .A0(\logix.ram_r[1252] ),
    .A1(\logix.ram_r[1260] ),
    .A2(\logix.ram_r[1268] ),
    .A3(\logix.ram_r[1276] ),
    .S1(_2941_),
    .X(_3337_));
 sg13g2_mux4_1 _9333_ (.S0(_2957_),
    .A0(\logix.ram_r[1220] ),
    .A1(\logix.ram_r[1228] ),
    .A2(\logix.ram_r[1236] ),
    .A3(\logix.ram_r[1244] ),
    .S1(_2355_),
    .X(_3338_));
 sg13g2_a22oi_1 _9334_ (.Y(_3339_),
    .B1(_3338_),
    .B2(_2965_),
    .A2(_3337_),
    .A1(_2593_));
 sg13g2_a21oi_1 _9335_ (.A1(_3336_),
    .A2(_3339_),
    .Y(_3340_),
    .B1(net50));
 sg13g2_mux4_1 _9336_ (.S0(_2384_),
    .A0(\logix.ram_r[1060] ),
    .A1(\logix.ram_r[1068] ),
    .A2(\logix.ram_r[1076] ),
    .A3(\logix.ram_r[1084] ),
    .S1(net197),
    .X(_3341_));
 sg13g2_mux4_1 _9337_ (.S0(net87),
    .A0(\logix.ram_r[1028] ),
    .A1(\logix.ram_r[1036] ),
    .A2(\logix.ram_r[1044] ),
    .A3(\logix.ram_r[1052] ),
    .S1(net86),
    .X(_3342_));
 sg13g2_a22oi_1 _9338_ (.Y(_3343_),
    .B1(_3342_),
    .B2(_2959_),
    .A2(_3341_),
    .A1(_2955_));
 sg13g2_mux4_1 _9339_ (.S0(_2992_),
    .A0(\logix.ram_r[1124] ),
    .A1(\logix.ram_r[1132] ),
    .A2(\logix.ram_r[1140] ),
    .A3(\logix.ram_r[1148] ),
    .S1(net181),
    .X(_3344_));
 sg13g2_mux4_1 _9340_ (.S0(net183),
    .A0(\logix.ram_r[1092] ),
    .A1(\logix.ram_r[1100] ),
    .A2(\logix.ram_r[1108] ),
    .A3(\logix.ram_r[1116] ),
    .S1(_2785_),
    .X(_3345_));
 sg13g2_a22oi_1 _9341_ (.Y(_3346_),
    .B1(_3345_),
    .B2(net91),
    .A2(_3344_),
    .A1(net126));
 sg13g2_a21oi_1 _9342_ (.A1(_3343_),
    .A2(_3346_),
    .Y(_3347_),
    .B1(_2967_));
 sg13g2_or2_1 _9343_ (.X(_3348_),
    .B(_3347_),
    .A(_3340_));
 sg13g2_a221oi_1 _9344_ (.B2(_2710_),
    .C1(_3348_),
    .B1(_3333_),
    .A1(_3315_),
    .Y(_3349_),
    .A2(_3322_));
 sg13g2_nand2b_1 _9345_ (.Y(_3350_),
    .B(net64),
    .A_N(\logix.ram_r[1876] ));
 sg13g2_o21ai_1 _9346_ (.B1(_3350_),
    .Y(_3351_),
    .A1(\logix.ram_r[1860] ),
    .A2(net60));
 sg13g2_nand2b_1 _9347_ (.Y(_3352_),
    .B(net63),
    .A_N(\logix.ram_r[1884] ));
 sg13g2_o21ai_1 _9348_ (.B1(_3352_),
    .Y(_3353_),
    .A1(\logix.ram_r[1868] ),
    .A2(net53));
 sg13g2_a221oi_1 _9349_ (.B2(net28),
    .C1(_2709_),
    .B1(_3353_),
    .A1(net29),
    .Y(_3354_),
    .A2(_3351_));
 sg13g2_mux4_1 _9350_ (.S0(net107),
    .A0(\logix.ram_r[1828] ),
    .A1(\logix.ram_r[1836] ),
    .A2(\logix.ram_r[1844] ),
    .A3(\logix.ram_r[1852] ),
    .S1(net111),
    .X(_3355_));
 sg13g2_mux4_1 _9351_ (.S0(net180),
    .A0(\logix.ram_r[1796] ),
    .A1(\logix.ram_r[1804] ),
    .A2(\logix.ram_r[1812] ),
    .A3(\logix.ram_r[1820] ),
    .S1(net181),
    .X(_3356_));
 sg13g2_and2_1 _9352_ (.A(net95),
    .B(_3356_),
    .X(_3357_));
 sg13g2_a221oi_1 _9353_ (.B2(net90),
    .C1(_3357_),
    .B1(_3355_),
    .A1(net206),
    .Y(_3358_),
    .A2(net205));
 sg13g2_mux4_1 _9354_ (.S0(net49),
    .A0(\logix.ram_r[1892] ),
    .A1(\logix.ram_r[1900] ),
    .A2(\logix.ram_r[1908] ),
    .A3(\logix.ram_r[1916] ),
    .S1(net58),
    .X(_3359_));
 sg13g2_nor2_1 _9355_ (.A(net89),
    .B(_3359_),
    .Y(_3360_));
 sg13g2_nor2_1 _9356_ (.A(_3358_),
    .B(_3360_),
    .Y(_3361_));
 sg13g2_mux4_1 _9357_ (.S0(net182),
    .A0(\logix.ram_r[1924] ),
    .A1(\logix.ram_r[1932] ),
    .A2(\logix.ram_r[1940] ),
    .A3(\logix.ram_r[1948] ),
    .S1(net93),
    .X(_3362_));
 sg13g2_mux4_1 _9358_ (.S0(net182),
    .A0(\logix.ram_r[1956] ),
    .A1(\logix.ram_r[1964] ),
    .A2(\logix.ram_r[1972] ),
    .A3(\logix.ram_r[1980] ),
    .S1(net92),
    .X(_3363_));
 sg13g2_mux2_1 _9359_ (.A0(_3362_),
    .A1(_3363_),
    .S(net199),
    .X(_3364_));
 sg13g2_nand2_1 _9360_ (.Y(_3365_),
    .A(net118),
    .B(_3364_));
 sg13g2_mux2_1 _9361_ (.A0(\logix.ram_r[1988] ),
    .A1(\logix.ram_r[1996] ),
    .S(net49),
    .X(_3366_));
 sg13g2_mux2_1 _9362_ (.A0(\logix.ram_r[2036] ),
    .A1(\logix.ram_r[2044] ),
    .S(net80),
    .X(_3367_));
 sg13g2_a22oi_1 _9363_ (.Y(_3368_),
    .B1(_3367_),
    .B2(net45),
    .A2(_3366_),
    .A1(net46));
 sg13g2_mux2_1 _9364_ (.A0(\logix.ram_r[2020] ),
    .A1(\logix.ram_r[2028] ),
    .S(net49),
    .X(_3369_));
 sg13g2_mux2_1 _9365_ (.A0(\logix.ram_r[2004] ),
    .A1(\logix.ram_r[2012] ),
    .S(net80),
    .X(_3370_));
 sg13g2_a22oi_1 _9366_ (.Y(_3371_),
    .B1(_3370_),
    .B2(net47),
    .A2(_3369_),
    .A1(net48));
 sg13g2_nand4_1 _9367_ (.B(_3365_),
    .C(_3368_),
    .A(_2780_),
    .Y(_3372_),
    .D(_3371_));
 sg13g2_mux4_1 _9368_ (.S0(net185),
    .A0(\logix.ram_r[1572] ),
    .A1(\logix.ram_r[1580] ),
    .A2(\logix.ram_r[1588] ),
    .A3(\logix.ram_r[1596] ),
    .S1(net175),
    .X(_3373_));
 sg13g2_mux4_1 _9369_ (.S0(net94),
    .A0(\logix.ram_r[1540] ),
    .A1(\logix.ram_r[1548] ),
    .A2(\logix.ram_r[1556] ),
    .A3(\logix.ram_r[1564] ),
    .S1(net101),
    .X(_3374_));
 sg13g2_a22oi_1 _9370_ (.Y(_3375_),
    .B1(_3374_),
    .B2(net55),
    .A2(_3373_),
    .A1(net56));
 sg13g2_mux4_1 _9371_ (.S0(net201),
    .A0(\logix.ram_r[1636] ),
    .A1(\logix.ram_r[1644] ),
    .A2(\logix.ram_r[1652] ),
    .A3(\logix.ram_r[1660] ),
    .S1(net197),
    .X(_3376_));
 sg13g2_mux4_1 _9372_ (.S0(net87),
    .A0(\logix.ram_r[1604] ),
    .A1(\logix.ram_r[1612] ),
    .A2(\logix.ram_r[1620] ),
    .A3(\logix.ram_r[1628] ),
    .S1(net86),
    .X(_3377_));
 sg13g2_a22oi_1 _9373_ (.Y(_3378_),
    .B1(_3377_),
    .B2(net91),
    .A2(_3376_),
    .A1(net85));
 sg13g2_a21oi_1 _9374_ (.A1(_3375_),
    .A2(_3378_),
    .Y(_3379_),
    .B1(net54));
 sg13g2_mux4_1 _9375_ (.S0(net183),
    .A0(\logix.ram_r[1700] ),
    .A1(\logix.ram_r[1708] ),
    .A2(\logix.ram_r[1716] ),
    .A3(\logix.ram_r[1724] ),
    .S1(net99),
    .X(_3380_));
 sg13g2_mux4_1 _9376_ (.S0(net122),
    .A0(\logix.ram_r[1668] ),
    .A1(\logix.ram_r[1676] ),
    .A2(\logix.ram_r[1684] ),
    .A3(\logix.ram_r[1692] ),
    .S1(net176),
    .X(_3381_));
 sg13g2_a22oi_1 _9377_ (.Y(_3382_),
    .B1(_3381_),
    .B2(net22),
    .A2(_3380_),
    .A1(net23));
 sg13g2_mux4_1 _9378_ (.S0(net182),
    .A0(\logix.ram_r[1764] ),
    .A1(\logix.ram_r[1772] ),
    .A2(\logix.ram_r[1780] ),
    .A3(\logix.ram_r[1788] ),
    .S1(net92),
    .X(_3383_));
 sg13g2_mux4_1 _9379_ (.S0(net109),
    .A0(\logix.ram_r[1732] ),
    .A1(\logix.ram_r[1740] ),
    .A2(\logix.ram_r[1748] ),
    .A3(\logix.ram_r[1756] ),
    .S1(net147),
    .X(_3384_));
 sg13g2_a22oi_1 _9380_ (.Y(_3385_),
    .B1(_3384_),
    .B2(net84),
    .A2(_3383_),
    .A1(net85));
 sg13g2_a21oi_1 _9381_ (.A1(_3382_),
    .A2(_3385_),
    .Y(_3386_),
    .B1(net50));
 sg13g2_or2_1 _9382_ (.X(_3387_),
    .B(_3386_),
    .A(_3379_));
 sg13g2_a221oi_1 _9383_ (.B2(_3047_),
    .C1(_3387_),
    .B1(_3372_),
    .A1(_3354_),
    .Y(_3388_),
    .A2(_3361_));
 sg13g2_mux4_1 _9384_ (.S0(_2391_),
    .A0(\logix.ram_r[900] ),
    .A1(\logix.ram_r[908] ),
    .A2(\logix.ram_r[916] ),
    .A3(\logix.ram_r[924] ),
    .S1(net193),
    .X(_3389_));
 sg13g2_mux4_1 _9385_ (.S0(net200),
    .A0(\logix.ram_r[932] ),
    .A1(\logix.ram_r[940] ),
    .A2(\logix.ram_r[948] ),
    .A3(\logix.ram_r[956] ),
    .S1(_2917_),
    .X(_3390_));
 sg13g2_mux2_1 _9386_ (.A0(_3389_),
    .A1(_3390_),
    .S(net187),
    .X(_3391_));
 sg13g2_mux2_1 _9387_ (.A0(\logix.ram_r[964] ),
    .A1(\logix.ram_r[972] ),
    .S(net195),
    .X(_3392_));
 sg13g2_nand3_1 _9388_ (.B(_2481_),
    .C(_3392_),
    .A(net207),
    .Y(_3393_));
 sg13g2_mux2_1 _9389_ (.A0(\logix.ram_r[1012] ),
    .A1(\logix.ram_r[1020] ),
    .S(_2615_),
    .X(_3394_));
 sg13g2_nand3_1 _9390_ (.B(_2472_),
    .C(_3394_),
    .A(net113),
    .Y(_3395_));
 sg13g2_mux2_1 _9391_ (.A0(\logix.ram_r[996] ),
    .A1(\logix.ram_r[1004] ),
    .S(net191),
    .X(_3396_));
 sg13g2_nand3_1 _9392_ (.B(net158),
    .C(_3396_),
    .A(net207),
    .Y(_3397_));
 sg13g2_mux2_1 _9393_ (.A0(\logix.ram_r[980] ),
    .A1(\logix.ram_r[988] ),
    .S(net191),
    .X(_3398_));
 sg13g2_nand3_1 _9394_ (.B(_2481_),
    .C(_3398_),
    .A(net163),
    .Y(_3399_));
 sg13g2_nand4_1 _9395_ (.B(_3395_),
    .C(_3397_),
    .A(_3393_),
    .Y(_3400_),
    .D(_3399_));
 sg13g2_a21oi_1 _9396_ (.A1(net174),
    .A2(_3391_),
    .Y(_3401_),
    .B1(_3400_));
 sg13g2_mux4_1 _9397_ (.S0(_2962_),
    .A0(\logix.ram_r[548] ),
    .A1(\logix.ram_r[556] ),
    .A2(\logix.ram_r[564] ),
    .A3(\logix.ram_r[572] ),
    .S1(_2963_),
    .X(_3402_));
 sg13g2_mux4_1 _9398_ (.S0(_2664_),
    .A0(\logix.ram_r[516] ),
    .A1(\logix.ram_r[524] ),
    .A2(\logix.ram_r[532] ),
    .A3(\logix.ram_r[540] ),
    .S1(_2512_),
    .X(_3403_));
 sg13g2_a22oi_1 _9399_ (.Y(_3404_),
    .B1(_3403_),
    .B2(_2959_),
    .A2(_3402_),
    .A1(_2955_));
 sg13g2_mux4_1 _9400_ (.S0(net196),
    .A0(\logix.ram_r[612] ),
    .A1(\logix.ram_r[620] ),
    .A2(\logix.ram_r[628] ),
    .A3(\logix.ram_r[636] ),
    .S1(net189),
    .X(_3405_));
 sg13g2_mux4_1 _9401_ (.S0(_2985_),
    .A0(\logix.ram_r[580] ),
    .A1(\logix.ram_r[588] ),
    .A2(\logix.ram_r[596] ),
    .A3(\logix.ram_r[604] ),
    .S1(_2686_),
    .X(_3406_));
 sg13g2_a22oi_1 _9402_ (.Y(_3407_),
    .B1(_3406_),
    .B2(_2965_),
    .A2(_3405_),
    .A1(_3053_));
 sg13g2_a21o_1 _9403_ (.A2(_3407_),
    .A1(_3404_),
    .B1(_2967_),
    .X(_3408_));
 sg13g2_o21ai_1 _9404_ (.B1(_3408_),
    .Y(_3409_),
    .A1(_2603_),
    .A2(_3401_));
 sg13g2_mux4_1 _9405_ (.S0(net172),
    .A0(\logix.ram_r[676] ),
    .A1(\logix.ram_r[684] ),
    .A2(\logix.ram_r[692] ),
    .A3(\logix.ram_r[700] ),
    .S1(net59),
    .X(_3410_));
 sg13g2_mux4_1 _9406_ (.S0(_3032_),
    .A0(\logix.ram_r[644] ),
    .A1(\logix.ram_r[652] ),
    .A2(\logix.ram_r[660] ),
    .A3(\logix.ram_r[668] ),
    .S1(net64),
    .X(_3411_));
 sg13g2_a22oi_1 _9407_ (.Y(_3412_),
    .B1(_3411_),
    .B2(_2492_),
    .A2(_3410_),
    .A1(_2488_));
 sg13g2_mux4_1 _9408_ (.S0(net172),
    .A0(\logix.ram_r[740] ),
    .A1(\logix.ram_r[748] ),
    .A2(\logix.ram_r[756] ),
    .A3(\logix.ram_r[764] ),
    .S1(_2590_),
    .X(_3413_));
 sg13g2_mux4_1 _9409_ (.S0(net52),
    .A0(\logix.ram_r[708] ),
    .A1(\logix.ram_r[716] ),
    .A2(\logix.ram_r[724] ),
    .A3(\logix.ram_r[732] ),
    .S1(_2641_),
    .X(_3414_));
 sg13g2_a22oi_1 _9410_ (.Y(_3415_),
    .B1(_3414_),
    .B2(net72),
    .A2(_3413_),
    .A1(_2594_));
 sg13g2_a21oi_1 _9411_ (.A1(_3412_),
    .A2(_3415_),
    .Y(_3416_),
    .B1(net71));
 sg13g2_mux4_1 _9412_ (.S0(net173),
    .A0(\logix.ram_r[804] ),
    .A1(\logix.ram_r[812] ),
    .A2(\logix.ram_r[820] ),
    .A3(\logix.ram_r[828] ),
    .S1(net110),
    .X(_3417_));
 sg13g2_mux4_1 _9413_ (.S0(_2985_),
    .A0(\logix.ram_r[772] ),
    .A1(\logix.ram_r[780] ),
    .A2(\logix.ram_r[788] ),
    .A3(\logix.ram_r[796] ),
    .S1(_2686_),
    .X(_3418_));
 sg13g2_and2_1 _9414_ (.A(_2879_),
    .B(_3418_),
    .X(_3419_));
 sg13g2_a221oi_1 _9415_ (.B2(net90),
    .C1(_3419_),
    .B1(_3417_),
    .A1(net206),
    .Y(_3420_),
    .A2(net205));
 sg13g2_nand2_1 _9416_ (.Y(_3421_),
    .A(\logix.ram_r[836] ),
    .B(_2378_));
 sg13g2_nand2_1 _9417_ (.Y(_3422_),
    .A(\logix.ram_r[852] ),
    .B(net128));
 sg13g2_nand3_1 _9418_ (.B(_3421_),
    .C(_3422_),
    .A(_2639_),
    .Y(_3423_));
 sg13g2_nand2_1 _9419_ (.Y(_3424_),
    .A(\logix.ram_r[844] ),
    .B(_2378_));
 sg13g2_nand2_1 _9420_ (.Y(_3425_),
    .A(\logix.ram_r[860] ),
    .B(_2588_));
 sg13g2_nand3_1 _9421_ (.B(_3424_),
    .C(_3425_),
    .A(_2647_),
    .Y(_3426_));
 sg13g2_nand3_1 _9422_ (.B(_3423_),
    .C(_3426_),
    .A(_2445_),
    .Y(_3427_));
 sg13g2_mux4_1 _9423_ (.S0(_2935_),
    .A0(\logix.ram_r[868] ),
    .A1(\logix.ram_r[876] ),
    .A2(\logix.ram_r[884] ),
    .A3(\logix.ram_r[892] ),
    .S1(_2681_),
    .X(_3428_));
 sg13g2_nor2_1 _9424_ (.A(net89),
    .B(_3428_),
    .Y(_3429_));
 sg13g2_nor3_1 _9425_ (.A(_3420_),
    .B(_3427_),
    .C(_3429_),
    .Y(_3430_));
 sg13g2_nor4_1 _9426_ (.A(_3147_),
    .B(_3409_),
    .C(_3416_),
    .D(_3430_),
    .Y(_3431_));
 sg13g2_nor4_2 _9427_ (.A(_3310_),
    .B(_3349_),
    .C(_3388_),
    .Y(net18),
    .D(_3431_));
 sg13g2_mux4_1 _9428_ (.S0(net115),
    .A0(\logix.ram_r[1285] ),
    .A1(\logix.ram_r[1293] ),
    .A2(\logix.ram_r[1301] ),
    .A3(\logix.ram_r[1309] ),
    .S1(net102),
    .X(_3432_));
 sg13g2_nor2_1 _9429_ (.A(net150),
    .B(_3432_),
    .Y(_3433_));
 sg13g2_mux2_1 _9430_ (.A0(\logix.ram_r[1317] ),
    .A1(\logix.ram_r[1333] ),
    .S(net104),
    .X(_3434_));
 sg13g2_nor2_1 _9431_ (.A(net83),
    .B(_3434_),
    .Y(_3435_));
 sg13g2_mux2_1 _9432_ (.A0(\logix.ram_r[1325] ),
    .A1(\logix.ram_r[1341] ),
    .S(net189),
    .X(_3436_));
 sg13g2_o21ai_1 _9433_ (.B1(net98),
    .Y(_3437_),
    .A1(net82),
    .A2(_3436_));
 sg13g2_nor3_1 _9434_ (.A(_3433_),
    .B(_3435_),
    .C(_3437_),
    .Y(_3438_));
 sg13g2_mux2_1 _9435_ (.A0(\logix.ram_r[1381] ),
    .A1(\logix.ram_r[1389] ),
    .S(net125),
    .X(_3439_));
 sg13g2_mux2_1 _9436_ (.A0(\logix.ram_r[1365] ),
    .A1(\logix.ram_r[1373] ),
    .S(net145),
    .X(_3440_));
 sg13g2_a22oi_1 _9437_ (.Y(_3441_),
    .B1(_3440_),
    .B2(net24),
    .A2(_3439_),
    .A1(net37));
 sg13g2_mux2_1 _9438_ (.A0(\logix.ram_r[1349] ),
    .A1(\logix.ram_r[1357] ),
    .S(net103),
    .X(_3442_));
 sg13g2_mux2_1 _9439_ (.A0(\logix.ram_r[1397] ),
    .A1(\logix.ram_r[1405] ),
    .S(net173),
    .X(_3443_));
 sg13g2_a22oi_1 _9440_ (.Y(_3444_),
    .B1(_3443_),
    .B2(net34),
    .A2(_3442_),
    .A1(net35));
 sg13g2_nand2_1 _9441_ (.Y(_3445_),
    .A(_3441_),
    .B(_3444_));
 sg13g2_o21ai_1 _9442_ (.B1(net79),
    .Y(_3446_),
    .A1(_3438_),
    .A2(_3445_));
 sg13g2_mux4_1 _9443_ (.S0(net102),
    .A0(\logix.ram_r[1413] ),
    .A1(\logix.ram_r[1429] ),
    .A2(\logix.ram_r[1445] ),
    .A3(\logix.ram_r[1461] ),
    .S1(net199),
    .X(_3447_));
 sg13g2_mux4_1 _9444_ (.S0(net143),
    .A0(\logix.ram_r[1421] ),
    .A1(\logix.ram_r[1437] ),
    .A2(\logix.ram_r[1453] ),
    .A3(\logix.ram_r[1469] ),
    .S1(_2535_),
    .X(_3448_));
 sg13g2_mux2_1 _9445_ (.A0(_3447_),
    .A1(_3448_),
    .S(net44),
    .X(_3449_));
 sg13g2_mux4_1 _9446_ (.S0(net141),
    .A0(\logix.ram_r[1477] ),
    .A1(\logix.ram_r[1485] ),
    .A2(\logix.ram_r[1493] ),
    .A3(\logix.ram_r[1501] ),
    .S1(net159),
    .X(_3450_));
 sg13g2_nor2_1 _9447_ (.A(net165),
    .B(_3450_),
    .Y(_3451_));
 sg13g2_mux2_1 _9448_ (.A0(\logix.ram_r[1517] ),
    .A1(\logix.ram_r[1533] ),
    .S(net177),
    .X(_3452_));
 sg13g2_nor2_1 _9449_ (.A(net43),
    .B(_3452_),
    .Y(_3453_));
 sg13g2_mux2_1 _9450_ (.A0(\logix.ram_r[1509] ),
    .A1(\logix.ram_r[1525] ),
    .S(net101),
    .X(_3454_));
 sg13g2_o21ai_1 _9451_ (.B1(_2406_),
    .Y(_3455_),
    .A1(net42),
    .A2(_3454_));
 sg13g2_nor3_1 _9452_ (.A(_3451_),
    .B(_3453_),
    .C(_3455_),
    .Y(_3456_));
 sg13g2_o21ai_1 _9453_ (.B1(_3456_),
    .Y(_3457_),
    .A1(net169),
    .A2(_3449_));
 sg13g2_mux4_1 _9454_ (.S0(net161),
    .A0(\logix.ram_r[1061] ),
    .A1(\logix.ram_r[1069] ),
    .A2(\logix.ram_r[1077] ),
    .A3(\logix.ram_r[1085] ),
    .S1(net168),
    .X(_3458_));
 sg13g2_mux4_1 _9455_ (.S0(net152),
    .A0(\logix.ram_r[1029] ),
    .A1(\logix.ram_r[1037] ),
    .A2(\logix.ram_r[1045] ),
    .A3(\logix.ram_r[1053] ),
    .S1(_2497_),
    .X(_3459_));
 sg13g2_a22oi_1 _9456_ (.Y(_3460_),
    .B1(_3459_),
    .B2(net25),
    .A2(_3458_),
    .A1(_2461_));
 sg13g2_mux4_1 _9457_ (.S0(net139),
    .A0(\logix.ram_r[1125] ),
    .A1(\logix.ram_r[1133] ),
    .A2(\logix.ram_r[1141] ),
    .A3(\logix.ram_r[1149] ),
    .S1(net143),
    .X(_3461_));
 sg13g2_mux4_1 _9458_ (.S0(net155),
    .A0(\logix.ram_r[1093] ),
    .A1(\logix.ram_r[1101] ),
    .A2(\logix.ram_r[1109] ),
    .A3(\logix.ram_r[1117] ),
    .S1(net137),
    .X(_3462_));
 sg13g2_a22oi_1 _9459_ (.Y(_3463_),
    .B1(_3462_),
    .B2(_2482_),
    .A2(_3461_),
    .A1(net76));
 sg13g2_a21oi_1 _9460_ (.A1(_3460_),
    .A2(_3463_),
    .Y(_3464_),
    .B1(net74));
 sg13g2_mux4_1 _9461_ (.S0(net178),
    .A0(\logix.ram_r[1189] ),
    .A1(\logix.ram_r[1197] ),
    .A2(\logix.ram_r[1205] ),
    .A3(\logix.ram_r[1213] ),
    .S1(net153),
    .X(_3465_));
 sg13g2_mux4_1 _9462_ (.S0(_2468_),
    .A0(\logix.ram_r[1157] ),
    .A1(\logix.ram_r[1165] ),
    .A2(\logix.ram_r[1173] ),
    .A3(\logix.ram_r[1181] ),
    .S1(net159),
    .X(_3466_));
 sg13g2_a22oi_1 _9463_ (.Y(_3467_),
    .B1(_3466_),
    .B2(net25),
    .A2(_3465_),
    .A1(net41));
 sg13g2_mux4_1 _9464_ (.S0(net117),
    .A0(\logix.ram_r[1253] ),
    .A1(\logix.ram_r[1261] ),
    .A2(\logix.ram_r[1269] ),
    .A3(\logix.ram_r[1277] ),
    .S1(net116),
    .X(_3468_));
 sg13g2_mux4_1 _9465_ (.S0(net152),
    .A0(\logix.ram_r[1221] ),
    .A1(\logix.ram_r[1229] ),
    .A2(\logix.ram_r[1237] ),
    .A3(\logix.ram_r[1245] ),
    .S1(net132),
    .X(_3469_));
 sg13g2_a22oi_1 _9466_ (.Y(_3470_),
    .B1(_3469_),
    .B2(net75),
    .A2(_3468_),
    .A1(net73));
 sg13g2_a21oi_1 _9467_ (.A1(_3467_),
    .A2(_3470_),
    .Y(_3471_),
    .B1(net71));
 sg13g2_nor2_1 _9468_ (.A(_3464_),
    .B(_3471_),
    .Y(_3472_));
 sg13g2_nand4_1 _9469_ (.B(_3446_),
    .C(_3457_),
    .A(_2706_),
    .Y(_3473_),
    .D(_3472_));
 sg13g2_mux4_1 _9470_ (.S0(net100),
    .A0(\logix.ram_r[901] ),
    .A1(\logix.ram_r[909] ),
    .A2(\logix.ram_r[917] ),
    .A3(\logix.ram_r[925] ),
    .S1(_2347_),
    .X(_3474_));
 sg13g2_nor2_1 _9471_ (.A(net188),
    .B(_3474_),
    .Y(_3475_));
 sg13g2_mux2_1 _9472_ (.A0(\logix.ram_r[933] ),
    .A1(\logix.ram_r[949] ),
    .S(net99),
    .X(_3476_));
 sg13g2_nor2_1 _9473_ (.A(_2345_),
    .B(_3476_),
    .Y(_3477_));
 sg13g2_mux2_1 _9474_ (.A0(\logix.ram_r[941] ),
    .A1(\logix.ram_r[957] ),
    .S(_2587_),
    .X(_3478_));
 sg13g2_o21ai_1 _9475_ (.B1(net98),
    .Y(_3479_),
    .A1(_2353_),
    .A2(_3478_));
 sg13g2_nor3_1 _9476_ (.A(_3475_),
    .B(_3477_),
    .C(_3479_),
    .Y(_3480_));
 sg13g2_mux2_1 _9477_ (.A0(\logix.ram_r[997] ),
    .A1(\logix.ram_r[1005] ),
    .S(net103),
    .X(_3481_));
 sg13g2_mux2_1 _9478_ (.A0(\logix.ram_r[981] ),
    .A1(\logix.ram_r[989] ),
    .S(net171),
    .X(_3482_));
 sg13g2_a22oi_1 _9479_ (.Y(_3483_),
    .B1(_3482_),
    .B2(net24),
    .A2(_3481_),
    .A1(_2520_));
 sg13g2_mux2_1 _9480_ (.A0(\logix.ram_r[965] ),
    .A1(\logix.ram_r[973] ),
    .S(_2702_),
    .X(_3484_));
 sg13g2_mux2_1 _9481_ (.A0(\logix.ram_r[1013] ),
    .A1(\logix.ram_r[1021] ),
    .S(net129),
    .X(_3485_));
 sg13g2_a22oi_1 _9482_ (.Y(_3486_),
    .B1(_3485_),
    .B2(net34),
    .A2(_3484_),
    .A1(net35));
 sg13g2_nand2_1 _9483_ (.Y(_3487_),
    .A(_3483_),
    .B(_3486_));
 sg13g2_o21ai_1 _9484_ (.B1(net81),
    .Y(_3488_),
    .A1(_3480_),
    .A2(_3487_));
 sg13g2_mux4_1 _9485_ (.S0(net121),
    .A0(\logix.ram_r[773] ),
    .A1(\logix.ram_r[789] ),
    .A2(\logix.ram_r[805] ),
    .A3(\logix.ram_r[821] ),
    .S1(net187),
    .X(_3489_));
 sg13g2_mux4_1 _9486_ (.S0(net101),
    .A0(\logix.ram_r[781] ),
    .A1(\logix.ram_r[797] ),
    .A2(\logix.ram_r[813] ),
    .A3(\logix.ram_r[829] ),
    .S1(net187),
    .X(_3490_));
 sg13g2_mux2_1 _9487_ (.A0(_3489_),
    .A1(_3490_),
    .S(net44),
    .X(_3491_));
 sg13g2_mux4_1 _9488_ (.S0(net133),
    .A0(\logix.ram_r[837] ),
    .A1(\logix.ram_r[845] ),
    .A2(\logix.ram_r[853] ),
    .A3(\logix.ram_r[861] ),
    .S1(net162),
    .X(_3492_));
 sg13g2_nor2_1 _9489_ (.A(net165),
    .B(_3492_),
    .Y(_3493_));
 sg13g2_mux2_1 _9490_ (.A0(\logix.ram_r[877] ),
    .A1(\logix.ram_r[893] ),
    .S(_2509_),
    .X(_3494_));
 sg13g2_nor2_1 _9491_ (.A(net43),
    .B(_3494_),
    .Y(_3495_));
 sg13g2_mux2_1 _9492_ (.A0(\logix.ram_r[869] ),
    .A1(\logix.ram_r[885] ),
    .S(net97),
    .X(_3496_));
 sg13g2_o21ai_1 _9493_ (.B1(net70),
    .Y(_3497_),
    .A1(net42),
    .A2(_3496_));
 sg13g2_nor3_1 _9494_ (.A(_3493_),
    .B(_3495_),
    .C(_3497_),
    .Y(_3498_));
 sg13g2_o21ai_1 _9495_ (.B1(_3498_),
    .Y(_3499_),
    .A1(net169),
    .A2(_3491_));
 sg13g2_mux4_1 _9496_ (.S0(net131),
    .A0(\logix.ram_r[677] ),
    .A1(\logix.ram_r[685] ),
    .A2(\logix.ram_r[693] ),
    .A3(\logix.ram_r[701] ),
    .S1(_2556_),
    .X(_3500_));
 sg13g2_mux4_1 _9497_ (.S0(net166),
    .A0(\logix.ram_r[645] ),
    .A1(\logix.ram_r[653] ),
    .A2(\logix.ram_r[661] ),
    .A3(\logix.ram_r[669] ),
    .S1(net137),
    .X(_3501_));
 sg13g2_a22oi_1 _9498_ (.Y(_3502_),
    .B1(_3501_),
    .B2(net30),
    .A2(_3500_),
    .A1(net31));
 sg13g2_mux4_1 _9499_ (.S0(_2563_),
    .A0(\logix.ram_r[741] ),
    .A1(\logix.ram_r[749] ),
    .A2(\logix.ram_r[757] ),
    .A3(\logix.ram_r[765] ),
    .S1(net135),
    .X(_3503_));
 sg13g2_mux4_1 _9500_ (.S0(_2566_),
    .A0(\logix.ram_r[709] ),
    .A1(\logix.ram_r[717] ),
    .A2(\logix.ram_r[725] ),
    .A3(\logix.ram_r[733] ),
    .S1(_2543_),
    .X(_3504_));
 sg13g2_a22oi_1 _9501_ (.Y(_3505_),
    .B1(_3504_),
    .B2(_2667_),
    .A2(_3503_),
    .A1(_2561_));
 sg13g2_a21oi_1 _9502_ (.A1(_3502_),
    .A2(_3505_),
    .Y(_3506_),
    .B1(_2570_));
 sg13g2_mux4_1 _9503_ (.S0(net149),
    .A0(\logix.ram_r[549] ),
    .A1(\logix.ram_r[557] ),
    .A2(\logix.ram_r[565] ),
    .A3(\logix.ram_r[573] ),
    .S1(net148),
    .X(_3507_));
 sg13g2_mux4_1 _9504_ (.S0(net133),
    .A0(\logix.ram_r[517] ),
    .A1(\logix.ram_r[525] ),
    .A2(\logix.ram_r[533] ),
    .A3(\logix.ram_r[541] ),
    .S1(net132),
    .X(_3508_));
 sg13g2_a22oi_1 _9505_ (.Y(_3509_),
    .B1(_3508_),
    .B2(net40),
    .A2(_3507_),
    .A1(net36));
 sg13g2_mux4_1 _9506_ (.S0(net131),
    .A0(\logix.ram_r[613] ),
    .A1(\logix.ram_r[621] ),
    .A2(\logix.ram_r[629] ),
    .A3(\logix.ram_r[637] ),
    .S1(net142),
    .X(_3510_));
 sg13g2_mux4_1 _9507_ (.S0(net105),
    .A0(\logix.ram_r[581] ),
    .A1(\logix.ram_r[589] ),
    .A2(\logix.ram_r[597] ),
    .A3(\logix.ram_r[605] ),
    .S1(net130),
    .X(_3511_));
 sg13g2_a22oi_1 _9508_ (.Y(_3512_),
    .B1(_3511_),
    .B2(net68),
    .A2(_3510_),
    .A1(net69));
 sg13g2_a21oi_1 _9509_ (.A1(_3509_),
    .A2(_3512_),
    .Y(_3513_),
    .B1(net66));
 sg13g2_nor2_1 _9510_ (.A(_3506_),
    .B(_3513_),
    .Y(_3514_));
 sg13g2_nand4_1 _9511_ (.B(_3488_),
    .C(_3499_),
    .A(_2553_),
    .Y(_3515_),
    .D(_3514_));
 sg13g2_mux4_1 _9512_ (.S0(net129),
    .A0(\logix.ram_r[37] ),
    .A1(\logix.ram_r[45] ),
    .A2(\logix.ram_r[53] ),
    .A3(\logix.ram_r[61] ),
    .S1(net128),
    .X(_3516_));
 sg13g2_mux4_1 _9513_ (.S0(net172),
    .A0(\logix.ram_r[5] ),
    .A1(\logix.ram_r[13] ),
    .A2(\logix.ram_r[21] ),
    .A3(\logix.ram_r[29] ),
    .S1(net127),
    .X(_3517_));
 sg13g2_a22oi_1 _9514_ (.Y(_3518_),
    .B1(_3517_),
    .B2(net38),
    .A2(_3516_),
    .A1(net39));
 sg13g2_mux4_1 _9515_ (.S0(net125),
    .A0(\logix.ram_r[101] ),
    .A1(\logix.ram_r[109] ),
    .A2(\logix.ram_r[117] ),
    .A3(\logix.ram_r[125] ),
    .S1(_2597_),
    .X(_3519_));
 sg13g2_mux4_1 _9516_ (.S0(_2524_),
    .A0(\logix.ram_r[69] ),
    .A1(\logix.ram_r[77] ),
    .A2(\logix.ram_r[85] ),
    .A3(\logix.ram_r[93] ),
    .S1(net110),
    .X(_3520_));
 sg13g2_a22oi_1 _9517_ (.Y(_3521_),
    .B1(_3520_),
    .B2(_2499_),
    .A2(_3519_),
    .A1(net73));
 sg13g2_a21o_1 _9518_ (.A2(_3521_),
    .A1(_3518_),
    .B1(net74),
    .X(_3522_));
 sg13g2_mux4_1 _9519_ (.S0(net157),
    .A0(\logix.ram_r[389] ),
    .A1(\logix.ram_r[397] ),
    .A2(\logix.ram_r[405] ),
    .A3(\logix.ram_r[413] ),
    .S1(net156),
    .X(_3523_));
 sg13g2_nand2_1 _9520_ (.Y(_3524_),
    .A(net95),
    .B(_3523_));
 sg13g2_mux4_1 _9521_ (.S0(net122),
    .A0(\logix.ram_r[421] ),
    .A1(\logix.ram_r[429] ),
    .A2(\logix.ram_r[437] ),
    .A3(\logix.ram_r[445] ),
    .S1(net121),
    .X(_3525_));
 sg13g2_nand2_1 _9522_ (.Y(_3526_),
    .A(net150),
    .B(_3525_));
 sg13g2_a21oi_1 _9523_ (.A1(_3524_),
    .A2(_3526_),
    .Y(_3527_),
    .B1(net120));
 sg13g2_mux2_1 _9524_ (.A0(\logix.ram_r[453] ),
    .A1(\logix.ram_r[461] ),
    .S(_2616_),
    .X(_3528_));
 sg13g2_mux2_1 _9525_ (.A0(\logix.ram_r[501] ),
    .A1(\logix.ram_r[509] ),
    .S(net129),
    .X(_3529_));
 sg13g2_a22oi_1 _9526_ (.Y(_3530_),
    .B1(_3529_),
    .B2(net34),
    .A2(_3528_),
    .A1(net35));
 sg13g2_mux2_1 _9527_ (.A0(\logix.ram_r[485] ),
    .A1(\logix.ram_r[493] ),
    .S(net96),
    .X(_3531_));
 sg13g2_mux2_1 _9528_ (.A0(\logix.ram_r[469] ),
    .A1(\logix.ram_r[477] ),
    .S(net144),
    .X(_3532_));
 sg13g2_a22oi_1 _9529_ (.Y(_3533_),
    .B1(_3532_),
    .B2(net32),
    .A2(_3531_),
    .A1(net33));
 sg13g2_nand2_1 _9530_ (.Y(_3534_),
    .A(_3530_),
    .B(_3533_));
 sg13g2_o21ai_1 _9531_ (.B1(net170),
    .Y(_3535_),
    .A1(_3527_),
    .A2(_3534_));
 sg13g2_mux4_1 _9532_ (.S0(net117),
    .A0(\logix.ram_r[261] ),
    .A1(\logix.ram_r[269] ),
    .A2(\logix.ram_r[277] ),
    .A3(\logix.ram_r[285] ),
    .S1(net116),
    .X(_3536_));
 sg13g2_nand2_1 _9533_ (.Y(_3537_),
    .A(_2605_),
    .B(_3536_));
 sg13g2_mux4_1 _9534_ (.S0(_2634_),
    .A0(\logix.ram_r[293] ),
    .A1(\logix.ram_r[301] ),
    .A2(\logix.ram_r[309] ),
    .A3(\logix.ram_r[317] ),
    .S1(_2417_),
    .X(_3538_));
 sg13g2_nand2_1 _9535_ (.Y(_3539_),
    .A(_2327_),
    .B(_3538_));
 sg13g2_nand3_1 _9536_ (.B(_3537_),
    .C(_3539_),
    .A(_2363_),
    .Y(_3540_));
 sg13g2_nand2b_1 _9537_ (.Y(_3541_),
    .B(net113),
    .A_N(\logix.ram_r[341] ));
 sg13g2_o21ai_1 _9538_ (.B1(_3541_),
    .Y(_3542_),
    .A1(\logix.ram_r[325] ),
    .A2(net59));
 sg13g2_nand2b_1 _9539_ (.Y(_3543_),
    .B(net111),
    .A_N(\logix.ram_r[349] ));
 sg13g2_o21ai_1 _9540_ (.B1(_3543_),
    .Y(_3544_),
    .A1(\logix.ram_r[333] ),
    .A2(_2900_));
 sg13g2_a22oi_1 _9541_ (.Y(_3545_),
    .B1(_3544_),
    .B2(_2647_),
    .A2(_3542_),
    .A1(_2639_));
 sg13g2_mux4_1 _9542_ (.S0(_2392_),
    .A0(\logix.ram_r[357] ),
    .A1(\logix.ram_r[365] ),
    .A2(\logix.ram_r[373] ),
    .A3(\logix.ram_r[381] ),
    .S1(_2654_),
    .X(_3546_));
 sg13g2_nand2b_1 _9543_ (.Y(_3547_),
    .B(net65),
    .A_N(_3546_));
 sg13g2_nand4_1 _9544_ (.B(_3540_),
    .C(_3545_),
    .A(_2445_),
    .Y(_3548_),
    .D(_3547_));
 sg13g2_mux4_1 _9545_ (.S0(net139),
    .A0(\logix.ram_r[165] ),
    .A1(\logix.ram_r[173] ),
    .A2(\logix.ram_r[181] ),
    .A3(\logix.ram_r[189] ),
    .S1(net143),
    .X(_3549_));
 sg13g2_mux4_1 _9546_ (.S0(net155),
    .A0(\logix.ram_r[133] ),
    .A1(\logix.ram_r[141] ),
    .A2(\logix.ram_r[149] ),
    .A3(\logix.ram_r[157] ),
    .S1(net137),
    .X(_3550_));
 sg13g2_a22oi_1 _9547_ (.Y(_3551_),
    .B1(_3550_),
    .B2(net40),
    .A2(_3549_),
    .A1(net36));
 sg13g2_mux4_1 _9548_ (.S0(net122),
    .A0(\logix.ram_r[229] ),
    .A1(\logix.ram_r[237] ),
    .A2(\logix.ram_r[245] ),
    .A3(\logix.ram_r[253] ),
    .S1(net135),
    .X(_3552_));
 sg13g2_mux4_1 _9549_ (.S0(net134),
    .A0(\logix.ram_r[197] ),
    .A1(\logix.ram_r[205] ),
    .A2(\logix.ram_r[213] ),
    .A3(\logix.ram_r[221] ),
    .S1(net140),
    .X(_3553_));
 sg13g2_a22oi_1 _9550_ (.Y(_3554_),
    .B1(_3553_),
    .B2(net68),
    .A2(_3552_),
    .A1(net69));
 sg13g2_a21oi_1 _9551_ (.A1(_3551_),
    .A2(_3554_),
    .Y(_3555_),
    .B1(net67));
 sg13g2_nor2_1 _9552_ (.A(_2455_),
    .B(_3555_),
    .Y(_3556_));
 sg13g2_nand4_1 _9553_ (.B(_3535_),
    .C(_3548_),
    .A(_3522_),
    .Y(_3557_),
    .D(_3556_));
 sg13g2_mux4_1 _9554_ (.S0(net109),
    .A0(\logix.ram_r[1925] ),
    .A1(\logix.ram_r[1933] ),
    .A2(\logix.ram_r[1941] ),
    .A3(\logix.ram_r[1949] ),
    .S1(net147),
    .X(_3558_));
 sg13g2_nor2_1 _9555_ (.A(net188),
    .B(_3558_),
    .Y(_3559_));
 sg13g2_mux2_1 _9556_ (.A0(\logix.ram_r[1957] ),
    .A1(\logix.ram_r[1973] ),
    .S(net92),
    .X(_3560_));
 sg13g2_nor2_1 _9557_ (.A(_2344_),
    .B(_3560_),
    .Y(_3561_));
 sg13g2_mux2_1 _9558_ (.A0(\logix.ram_r[1965] ),
    .A1(\logix.ram_r[1981] ),
    .S(net186),
    .X(_3562_));
 sg13g2_o21ai_1 _9559_ (.B1(net98),
    .Y(_3563_),
    .A1(_2352_),
    .A2(_3562_));
 sg13g2_nor3_1 _9560_ (.A(_3559_),
    .B(_3561_),
    .C(_3563_),
    .Y(_3564_));
 sg13g2_mux2_1 _9561_ (.A0(\logix.ram_r[2021] ),
    .A1(\logix.ram_r[2029] ),
    .S(net119),
    .X(_3565_));
 sg13g2_mux2_1 _9562_ (.A0(\logix.ram_r[2005] ),
    .A1(\logix.ram_r[2013] ),
    .S(net146),
    .X(_3566_));
 sg13g2_a22oi_1 _9563_ (.Y(_3567_),
    .B1(_3566_),
    .B2(net24),
    .A2(_3565_),
    .A1(net33));
 sg13g2_mux2_1 _9564_ (.A0(\logix.ram_r[1989] ),
    .A1(\logix.ram_r[1997] ),
    .S(net96),
    .X(_3568_));
 sg13g2_mux2_1 _9565_ (.A0(\logix.ram_r[2037] ),
    .A1(\logix.ram_r[2045] ),
    .S(net144),
    .X(_3569_));
 sg13g2_a22oi_1 _9566_ (.Y(_3570_),
    .B1(_3569_),
    .B2(net26),
    .A2(_3568_),
    .A1(net27));
 sg13g2_nand2_1 _9567_ (.Y(_3571_),
    .A(_3567_),
    .B(_3570_));
 sg13g2_o21ai_1 _9568_ (.B1(net170),
    .Y(_3572_),
    .A1(_3564_),
    .A2(_3571_));
 sg13g2_mux4_1 _9569_ (.S0(net104),
    .A0(\logix.ram_r[1797] ),
    .A1(\logix.ram_r[1813] ),
    .A2(\logix.ram_r[1829] ),
    .A3(\logix.ram_r[1845] ),
    .S1(net187),
    .X(_3573_));
 sg13g2_mux4_1 _9570_ (.S0(net97),
    .A0(\logix.ram_r[1805] ),
    .A1(\logix.ram_r[1821] ),
    .A2(\logix.ram_r[1837] ),
    .A3(\logix.ram_r[1853] ),
    .S1(net204),
    .X(_3574_));
 sg13g2_mux2_1 _9571_ (.A0(_3573_),
    .A1(_3574_),
    .S(net57),
    .X(_3575_));
 sg13g2_mux4_1 _9572_ (.S0(net178),
    .A0(\logix.ram_r[1861] ),
    .A1(\logix.ram_r[1869] ),
    .A2(\logix.ram_r[1877] ),
    .A3(\logix.ram_r[1885] ),
    .S1(net153),
    .X(_3576_));
 sg13g2_nor2_1 _9573_ (.A(net202),
    .B(_3576_),
    .Y(_3577_));
 sg13g2_mux2_1 _9574_ (.A0(\logix.ram_r[1901] ),
    .A1(\logix.ram_r[1917] ),
    .S(net142),
    .X(_3578_));
 sg13g2_nor2_1 _9575_ (.A(_2433_),
    .B(_3578_),
    .Y(_3579_));
 sg13g2_mux2_1 _9576_ (.A0(\logix.ram_r[1893] ),
    .A1(\logix.ram_r[1909] ),
    .S(net99),
    .X(_3580_));
 sg13g2_o21ai_1 _9577_ (.B1(net70),
    .Y(_3581_),
    .A1(_2439_),
    .A2(_3580_));
 sg13g2_nor3_1 _9578_ (.A(_3577_),
    .B(_3579_),
    .C(_3581_),
    .Y(_3582_));
 sg13g2_o21ai_1 _9579_ (.B1(_3582_),
    .Y(_3583_),
    .A1(net120),
    .A2(_3575_));
 sg13g2_mux4_1 _9580_ (.S0(net94),
    .A0(\logix.ram_r[1701] ),
    .A1(\logix.ram_r[1709] ),
    .A2(\logix.ram_r[1717] ),
    .A3(\logix.ram_r[1725] ),
    .S1(net114),
    .X(_3584_));
 sg13g2_mux4_1 _9581_ (.S0(net106),
    .A0(\logix.ram_r[1669] ),
    .A1(\logix.ram_r[1677] ),
    .A2(\logix.ram_r[1685] ),
    .A3(\logix.ram_r[1693] ),
    .S1(net112),
    .X(_3585_));
 sg13g2_a22oi_1 _9582_ (.Y(_3586_),
    .B1(_3585_),
    .B2(net22),
    .A2(_3584_),
    .A1(net23));
 sg13g2_mux4_1 _9583_ (.S0(net87),
    .A0(\logix.ram_r[1765] ),
    .A1(\logix.ram_r[1773] ),
    .A2(\logix.ram_r[1781] ),
    .A3(\logix.ram_r[1789] ),
    .S1(net86),
    .X(_3587_));
 sg13g2_mux4_1 _9584_ (.S0(net157),
    .A0(\logix.ram_r[1733] ),
    .A1(\logix.ram_r[1741] ),
    .A2(\logix.ram_r[1749] ),
    .A3(\logix.ram_r[1757] ),
    .S1(net102),
    .X(_3588_));
 sg13g2_a22oi_1 _9585_ (.Y(_3589_),
    .B1(_3588_),
    .B2(net84),
    .A2(_3587_),
    .A1(net62));
 sg13g2_a21oi_1 _9586_ (.A1(_3586_),
    .A2(_3589_),
    .Y(_3590_),
    .B1(net50));
 sg13g2_mux4_1 _9587_ (.S0(net100),
    .A0(\logix.ram_r[1573] ),
    .A1(\logix.ram_r[1581] ),
    .A2(\logix.ram_r[1589] ),
    .A3(\logix.ram_r[1597] ),
    .S1(net142),
    .X(_3591_));
 sg13g2_mux4_1 _9588_ (.S0(net105),
    .A0(\logix.ram_r[1541] ),
    .A1(\logix.ram_r[1549] ),
    .A2(\logix.ram_r[1557] ),
    .A3(\logix.ram_r[1565] ),
    .S1(net130),
    .X(_3592_));
 sg13g2_a22oi_1 _9589_ (.Y(_3593_),
    .B1(_3592_),
    .B2(net30),
    .A2(_3591_),
    .A1(net31));
 sg13g2_mux4_1 _9590_ (.S0(net94),
    .A0(\logix.ram_r[1637] ),
    .A1(\logix.ram_r[1645] ),
    .A2(\logix.ram_r[1653] ),
    .A3(\logix.ram_r[1661] ),
    .S1(net114),
    .X(_3594_));
 sg13g2_mux4_1 _9591_ (.S0(net161),
    .A0(\logix.ram_r[1605] ),
    .A1(\logix.ram_r[1613] ),
    .A2(\logix.ram_r[1621] ),
    .A3(\logix.ram_r[1629] ),
    .S1(net112),
    .X(_3595_));
 sg13g2_a22oi_1 _9592_ (.Y(_3596_),
    .B1(_3595_),
    .B2(net61),
    .A2(_3594_),
    .A1(net62));
 sg13g2_a21oi_1 _9593_ (.A1(_3593_),
    .A2(_3596_),
    .Y(_3597_),
    .B1(net66));
 sg13g2_nor2_1 _9594_ (.A(_3590_),
    .B(_3597_),
    .Y(_3598_));
 sg13g2_nand4_1 _9595_ (.B(_3572_),
    .C(_3583_),
    .A(_2780_),
    .Y(_3599_),
    .D(_3598_));
 sg13g2_and4_1 _9596_ (.A(_3473_),
    .B(_3515_),
    .C(_3557_),
    .D(_3599_),
    .X(net19));
 sg13g2_mux4_1 _9597_ (.S0(net115),
    .A0(\logix.ram_r[1286] ),
    .A1(\logix.ram_r[1294] ),
    .A2(\logix.ram_r[1302] ),
    .A3(\logix.ram_r[1310] ),
    .S1(net102),
    .X(_3600_));
 sg13g2_nor2_1 _9598_ (.A(net150),
    .B(_3600_),
    .Y(_3601_));
 sg13g2_mux2_1 _9599_ (.A0(\logix.ram_r[1318] ),
    .A1(\logix.ram_r[1334] ),
    .S(net104),
    .X(_3602_));
 sg13g2_nor2_1 _9600_ (.A(net83),
    .B(_3602_),
    .Y(_3603_));
 sg13g2_mux2_1 _9601_ (.A0(\logix.ram_r[1326] ),
    .A1(\logix.ram_r[1342] ),
    .S(net189),
    .X(_3604_));
 sg13g2_o21ai_1 _9602_ (.B1(net98),
    .Y(_3605_),
    .A1(net82),
    .A2(_3604_));
 sg13g2_nor3_1 _9603_ (.A(_3601_),
    .B(_3603_),
    .C(_3605_),
    .Y(_3606_));
 sg13g2_mux2_1 _9604_ (.A0(\logix.ram_r[1382] ),
    .A1(\logix.ram_r[1390] ),
    .S(net125),
    .X(_3607_));
 sg13g2_mux2_1 _9605_ (.A0(\logix.ram_r[1366] ),
    .A1(\logix.ram_r[1374] ),
    .S(net145),
    .X(_3608_));
 sg13g2_a22oi_1 _9606_ (.Y(_3609_),
    .B1(_3608_),
    .B2(net24),
    .A2(_3607_),
    .A1(net37));
 sg13g2_mux2_1 _9607_ (.A0(\logix.ram_r[1350] ),
    .A1(\logix.ram_r[1358] ),
    .S(net103),
    .X(_3610_));
 sg13g2_mux2_1 _9608_ (.A0(\logix.ram_r[1398] ),
    .A1(\logix.ram_r[1406] ),
    .S(net173),
    .X(_3611_));
 sg13g2_a22oi_1 _9609_ (.Y(_3612_),
    .B1(_3611_),
    .B2(net34),
    .A2(_3610_),
    .A1(net35));
 sg13g2_nand2_1 _9610_ (.Y(_3613_),
    .A(_3609_),
    .B(_3612_));
 sg13g2_o21ai_1 _9611_ (.B1(net79),
    .Y(_3614_),
    .A1(_3606_),
    .A2(_3613_));
 sg13g2_mux4_1 _9612_ (.S0(_2750_),
    .A0(\logix.ram_r[1414] ),
    .A1(\logix.ram_r[1430] ),
    .A2(\logix.ram_r[1446] ),
    .A3(\logix.ram_r[1462] ),
    .S1(_2414_),
    .X(_3615_));
 sg13g2_mux4_1 _9613_ (.S0(net143),
    .A0(\logix.ram_r[1422] ),
    .A1(\logix.ram_r[1438] ),
    .A2(\logix.ram_r[1454] ),
    .A3(\logix.ram_r[1470] ),
    .S1(net194),
    .X(_3616_));
 sg13g2_mux2_1 _9614_ (.A0(_3615_),
    .A1(_3616_),
    .S(net44),
    .X(_3617_));
 sg13g2_mux4_1 _9615_ (.S0(net141),
    .A0(\logix.ram_r[1478] ),
    .A1(\logix.ram_r[1486] ),
    .A2(\logix.ram_r[1494] ),
    .A3(\logix.ram_r[1502] ),
    .S1(net159),
    .X(_3618_));
 sg13g2_nor2_1 _9616_ (.A(net165),
    .B(_3618_),
    .Y(_3619_));
 sg13g2_mux2_1 _9617_ (.A0(\logix.ram_r[1518] ),
    .A1(\logix.ram_r[1534] ),
    .S(net177),
    .X(_3620_));
 sg13g2_nor2_1 _9618_ (.A(net43),
    .B(_3620_),
    .Y(_3621_));
 sg13g2_mux2_1 _9619_ (.A0(\logix.ram_r[1510] ),
    .A1(\logix.ram_r[1526] ),
    .S(net114),
    .X(_3622_));
 sg13g2_o21ai_1 _9620_ (.B1(_2406_),
    .Y(_3623_),
    .A1(net42),
    .A2(_3622_));
 sg13g2_nor3_1 _9621_ (.A(_3619_),
    .B(_3621_),
    .C(_3623_),
    .Y(_3624_));
 sg13g2_o21ai_1 _9622_ (.B1(_3624_),
    .Y(_3625_),
    .A1(net169),
    .A2(_3617_));
 sg13g2_mux4_1 _9623_ (.S0(_2463_),
    .A0(\logix.ram_r[1062] ),
    .A1(\logix.ram_r[1070] ),
    .A2(\logix.ram_r[1078] ),
    .A3(\logix.ram_r[1086] ),
    .S1(_2413_),
    .X(_3626_));
 sg13g2_mux4_1 _9624_ (.S0(net152),
    .A0(\logix.ram_r[1030] ),
    .A1(\logix.ram_r[1038] ),
    .A2(\logix.ram_r[1046] ),
    .A3(\logix.ram_r[1054] ),
    .S1(net151),
    .X(_3627_));
 sg13g2_a22oi_1 _9625_ (.Y(_3628_),
    .B1(_3627_),
    .B2(_2715_),
    .A2(_3626_),
    .A1(_2461_));
 sg13g2_mux4_1 _9626_ (.S0(_2555_),
    .A0(\logix.ram_r[1126] ),
    .A1(\logix.ram_r[1134] ),
    .A2(\logix.ram_r[1142] ),
    .A3(\logix.ram_r[1150] ),
    .S1(net143),
    .X(_3629_));
 sg13g2_mux4_1 _9627_ (.S0(net155),
    .A0(\logix.ram_r[1094] ),
    .A1(\logix.ram_r[1102] ),
    .A2(\logix.ram_r[1110] ),
    .A3(\logix.ram_r[1118] ),
    .S1(_2558_),
    .X(_3630_));
 sg13g2_a22oi_1 _9628_ (.Y(_3631_),
    .B1(_3630_),
    .B2(_2482_),
    .A2(_3629_),
    .A1(_2473_));
 sg13g2_a21oi_1 _9629_ (.A1(_3628_),
    .A2(_3631_),
    .Y(_3632_),
    .B1(_2486_));
 sg13g2_mux4_1 _9630_ (.S0(_2332_),
    .A0(\logix.ram_r[1190] ),
    .A1(\logix.ram_r[1198] ),
    .A2(\logix.ram_r[1206] ),
    .A3(\logix.ram_r[1214] ),
    .S1(net153),
    .X(_3633_));
 sg13g2_mux4_1 _9631_ (.S0(net160),
    .A0(\logix.ram_r[1158] ),
    .A1(\logix.ram_r[1166] ),
    .A2(\logix.ram_r[1174] ),
    .A3(\logix.ram_r[1182] ),
    .S1(net159),
    .X(_3634_));
 sg13g2_a22oi_1 _9632_ (.Y(_3635_),
    .B1(_3634_),
    .B2(net25),
    .A2(_3633_),
    .A1(net41));
 sg13g2_mux4_1 _9633_ (.S0(_2630_),
    .A0(\logix.ram_r[1254] ),
    .A1(\logix.ram_r[1262] ),
    .A2(\logix.ram_r[1270] ),
    .A3(\logix.ram_r[1278] ),
    .S1(_2631_),
    .X(_3636_));
 sg13g2_mux4_1 _9634_ (.S0(_2496_),
    .A0(\logix.ram_r[1222] ),
    .A1(\logix.ram_r[1230] ),
    .A2(\logix.ram_r[1238] ),
    .A3(\logix.ram_r[1246] ),
    .S1(_2574_),
    .X(_3637_));
 sg13g2_a22oi_1 _9635_ (.Y(_3638_),
    .B1(_3637_),
    .B2(net75),
    .A2(_3636_),
    .A1(_2494_));
 sg13g2_a21oi_1 _9636_ (.A1(_3635_),
    .A2(_3638_),
    .Y(_3639_),
    .B1(net71));
 sg13g2_nor2_1 _9637_ (.A(_3632_),
    .B(_3639_),
    .Y(_3640_));
 sg13g2_nand4_1 _9638_ (.B(_3614_),
    .C(_3625_),
    .A(_2706_),
    .Y(_3641_),
    .D(_3640_));
 sg13g2_mux4_1 _9639_ (.S0(net100),
    .A0(\logix.ram_r[390] ),
    .A1(\logix.ram_r[398] ),
    .A2(\logix.ram_r[406] ),
    .A3(\logix.ram_r[414] ),
    .S1(net176),
    .X(_3642_));
 sg13g2_nor2_1 _9640_ (.A(net188),
    .B(_3642_),
    .Y(_3643_));
 sg13g2_mux2_1 _9641_ (.A0(\logix.ram_r[422] ),
    .A1(\logix.ram_r[438] ),
    .S(net99),
    .X(_3644_));
 sg13g2_nor2_1 _9642_ (.A(net83),
    .B(_3644_),
    .Y(_3645_));
 sg13g2_mux2_1 _9643_ (.A0(\logix.ram_r[430] ),
    .A1(\logix.ram_r[446] ),
    .S(net193),
    .X(_3646_));
 sg13g2_o21ai_1 _9644_ (.B1(net98),
    .Y(_3647_),
    .A1(net82),
    .A2(_3646_));
 sg13g2_nor3_1 _9645_ (.A(_3643_),
    .B(_3645_),
    .C(_3647_),
    .Y(_3648_));
 sg13g2_mux2_1 _9646_ (.A0(\logix.ram_r[486] ),
    .A1(\logix.ram_r[494] ),
    .S(net103),
    .X(_3649_));
 sg13g2_mux2_1 _9647_ (.A0(\logix.ram_r[470] ),
    .A1(\logix.ram_r[478] ),
    .S(net171),
    .X(_3650_));
 sg13g2_a22oi_1 _9648_ (.Y(_3651_),
    .B1(_3650_),
    .B2(net24),
    .A2(_3649_),
    .A1(net37));
 sg13g2_mux2_1 _9649_ (.A0(\logix.ram_r[454] ),
    .A1(\logix.ram_r[462] ),
    .S(net107),
    .X(_3652_));
 sg13g2_mux2_1 _9650_ (.A0(\logix.ram_r[502] ),
    .A1(\logix.ram_r[510] ),
    .S(_2586_),
    .X(_3653_));
 sg13g2_a22oi_1 _9651_ (.Y(_3654_),
    .B1(_3653_),
    .B2(_2619_),
    .A2(_3652_),
    .A1(_2614_));
 sg13g2_nand2_1 _9652_ (.Y(_3655_),
    .A(_3651_),
    .B(_3654_));
 sg13g2_o21ai_1 _9653_ (.B1(net81),
    .Y(_3656_),
    .A1(_3648_),
    .A2(_3655_));
 sg13g2_mux4_1 _9654_ (.S0(net121),
    .A0(\logix.ram_r[262] ),
    .A1(\logix.ram_r[278] ),
    .A2(\logix.ram_r[294] ),
    .A3(\logix.ram_r[310] ),
    .S1(net187),
    .X(_3657_));
 sg13g2_mux4_1 _9655_ (.S0(_2758_),
    .A0(\logix.ram_r[270] ),
    .A1(\logix.ram_r[286] ),
    .A2(\logix.ram_r[302] ),
    .A3(\logix.ram_r[318] ),
    .S1(net187),
    .X(_3658_));
 sg13g2_mux2_1 _9656_ (.A0(_3657_),
    .A1(_3658_),
    .S(net44),
    .X(_3659_));
 sg13g2_mux4_1 _9657_ (.S0(_2573_),
    .A0(\logix.ram_r[326] ),
    .A1(\logix.ram_r[334] ),
    .A2(\logix.ram_r[342] ),
    .A3(\logix.ram_r[350] ),
    .S1(_2435_),
    .X(_3660_));
 sg13g2_nor2_1 _9658_ (.A(net165),
    .B(_3660_),
    .Y(_3661_));
 sg13g2_mux2_1 _9659_ (.A0(\logix.ram_r[366] ),
    .A1(\logix.ram_r[382] ),
    .S(_2509_),
    .X(_3662_));
 sg13g2_nor2_1 _9660_ (.A(_2434_),
    .B(_3662_),
    .Y(_3663_));
 sg13g2_mux2_1 _9661_ (.A0(\logix.ram_r[358] ),
    .A1(\logix.ram_r[374] ),
    .S(net97),
    .X(_3664_));
 sg13g2_o21ai_1 _9662_ (.B1(net70),
    .Y(_3665_),
    .A1(net42),
    .A2(_3664_));
 sg13g2_nor3_1 _9663_ (.A(_3661_),
    .B(_3663_),
    .C(_3665_),
    .Y(_3666_));
 sg13g2_o21ai_1 _9664_ (.B1(_3666_),
    .Y(_3667_),
    .A1(net169),
    .A2(_3659_));
 sg13g2_mux4_1 _9665_ (.S0(net131),
    .A0(\logix.ram_r[166] ),
    .A1(\logix.ram_r[174] ),
    .A2(\logix.ram_r[182] ),
    .A3(\logix.ram_r[190] ),
    .S1(net138),
    .X(_3668_));
 sg13g2_mux4_1 _9666_ (.S0(net166),
    .A0(\logix.ram_r[134] ),
    .A1(\logix.ram_r[142] ),
    .A2(\logix.ram_r[150] ),
    .A3(\logix.ram_r[158] ),
    .S1(net137),
    .X(_3669_));
 sg13g2_a22oi_1 _9667_ (.Y(_3670_),
    .B1(_3669_),
    .B2(net30),
    .A2(_3668_),
    .A1(net31));
 sg13g2_mux4_1 _9668_ (.S0(net136),
    .A0(\logix.ram_r[230] ),
    .A1(\logix.ram_r[238] ),
    .A2(\logix.ram_r[246] ),
    .A3(\logix.ram_r[254] ),
    .S1(net135),
    .X(_3671_));
 sg13g2_mux4_1 _9669_ (.S0(net134),
    .A0(\logix.ram_r[198] ),
    .A1(\logix.ram_r[206] ),
    .A2(\logix.ram_r[214] ),
    .A3(\logix.ram_r[222] ),
    .S1(net140),
    .X(_3672_));
 sg13g2_a22oi_1 _9670_ (.Y(_3673_),
    .B1(_3672_),
    .B2(net61),
    .A2(_3671_),
    .A1(net69));
 sg13g2_a21oi_1 _9671_ (.A1(_3670_),
    .A2(_3673_),
    .Y(_3674_),
    .B1(net67));
 sg13g2_mux4_1 _9672_ (.S0(_2508_),
    .A0(\logix.ram_r[38] ),
    .A1(\logix.ram_r[46] ),
    .A2(\logix.ram_r[54] ),
    .A3(\logix.ram_r[62] ),
    .S1(net148),
    .X(_3675_));
 sg13g2_mux4_1 _9673_ (.S0(net133),
    .A0(\logix.ram_r[6] ),
    .A1(\logix.ram_r[14] ),
    .A2(\logix.ram_r[22] ),
    .A3(\logix.ram_r[30] ),
    .S1(net132),
    .X(_3676_));
 sg13g2_a22oi_1 _9674_ (.Y(_3677_),
    .B1(_3676_),
    .B2(net40),
    .A2(_3675_),
    .A1(net36));
 sg13g2_mux4_1 _9675_ (.S0(_2577_),
    .A0(\logix.ram_r[102] ),
    .A1(\logix.ram_r[110] ),
    .A2(\logix.ram_r[118] ),
    .A3(\logix.ram_r[126] ),
    .S1(net142),
    .X(_3678_));
 sg13g2_mux4_1 _9676_ (.S0(net105),
    .A0(\logix.ram_r[70] ),
    .A1(\logix.ram_r[78] ),
    .A2(\logix.ram_r[86] ),
    .A3(\logix.ram_r[94] ),
    .S1(net130),
    .X(_3679_));
 sg13g2_a22oi_1 _9677_ (.Y(_3680_),
    .B1(_3679_),
    .B2(net68),
    .A2(_3678_),
    .A1(net69));
 sg13g2_a21oi_1 _9678_ (.A1(_3677_),
    .A2(_3680_),
    .Y(_3681_),
    .B1(net66));
 sg13g2_nor2_1 _9679_ (.A(_3674_),
    .B(_3681_),
    .Y(_3682_));
 sg13g2_nand4_1 _9680_ (.B(_3656_),
    .C(_3667_),
    .A(_2456_),
    .Y(_3683_),
    .D(_3682_));
 sg13g2_mux4_1 _9681_ (.S0(net146),
    .A0(\logix.ram_r[1574] ),
    .A1(\logix.ram_r[1582] ),
    .A2(\logix.ram_r[1590] ),
    .A3(\logix.ram_r[1598] ),
    .S1(net128),
    .X(_3684_));
 sg13g2_mux4_1 _9682_ (.S0(net172),
    .A0(\logix.ram_r[1542] ),
    .A1(\logix.ram_r[1550] ),
    .A2(\logix.ram_r[1558] ),
    .A3(\logix.ram_r[1566] ),
    .S1(net127),
    .X(_3685_));
 sg13g2_a22oi_1 _9683_ (.Y(_3686_),
    .B1(_3685_),
    .B2(net38),
    .A2(_3684_),
    .A1(net39));
 sg13g2_mux4_1 _9684_ (.S0(net125),
    .A0(\logix.ram_r[1638] ),
    .A1(\logix.ram_r[1646] ),
    .A2(\logix.ram_r[1654] ),
    .A3(\logix.ram_r[1662] ),
    .S1(net124),
    .X(_3687_));
 sg13g2_mux4_1 _9685_ (.S0(net173),
    .A0(\logix.ram_r[1606] ),
    .A1(\logix.ram_r[1614] ),
    .A2(\logix.ram_r[1622] ),
    .A3(\logix.ram_r[1630] ),
    .S1(net110),
    .X(_3688_));
 sg13g2_a22oi_1 _9686_ (.Y(_3689_),
    .B1(_3688_),
    .B2(net72),
    .A2(_3687_),
    .A1(net73));
 sg13g2_a21o_1 _9687_ (.A2(_3689_),
    .A1(_3686_),
    .B1(net74),
    .X(_3690_));
 sg13g2_mux4_1 _9688_ (.S0(net157),
    .A0(\logix.ram_r[1926] ),
    .A1(\logix.ram_r[1934] ),
    .A2(\logix.ram_r[1942] ),
    .A3(\logix.ram_r[1950] ),
    .S1(net156),
    .X(_3691_));
 sg13g2_nand2_1 _9689_ (.Y(_3692_),
    .A(net95),
    .B(_3691_));
 sg13g2_mux4_1 _9690_ (.S0(net122),
    .A0(\logix.ram_r[1958] ),
    .A1(\logix.ram_r[1966] ),
    .A2(\logix.ram_r[1974] ),
    .A3(\logix.ram_r[1982] ),
    .S1(net121),
    .X(_3693_));
 sg13g2_nand2_1 _9691_ (.Y(_3694_),
    .A(net150),
    .B(_3693_));
 sg13g2_a21oi_1 _9692_ (.A1(_3692_),
    .A2(_3694_),
    .Y(_3695_),
    .B1(net120));
 sg13g2_mux2_1 _9693_ (.A0(\logix.ram_r[1990] ),
    .A1(\logix.ram_r[1998] ),
    .S(net119),
    .X(_3696_));
 sg13g2_mux2_1 _9694_ (.A0(\logix.ram_r[2038] ),
    .A1(\logix.ram_r[2046] ),
    .S(net129),
    .X(_3697_));
 sg13g2_a22oi_1 _9695_ (.Y(_3698_),
    .B1(_3697_),
    .B2(net26),
    .A2(_3696_),
    .A1(net27));
 sg13g2_mux2_1 _9696_ (.A0(\logix.ram_r[2022] ),
    .A1(\logix.ram_r[2030] ),
    .S(net96),
    .X(_3699_));
 sg13g2_mux2_1 _9697_ (.A0(\logix.ram_r[2006] ),
    .A1(\logix.ram_r[2014] ),
    .S(net144),
    .X(_3700_));
 sg13g2_a22oi_1 _9698_ (.Y(_3701_),
    .B1(_3700_),
    .B2(net32),
    .A2(_3699_),
    .A1(net33));
 sg13g2_nand2_1 _9699_ (.Y(_3702_),
    .A(_3698_),
    .B(_3701_));
 sg13g2_o21ai_1 _9700_ (.B1(net170),
    .Y(_3703_),
    .A1(_3695_),
    .A2(_3702_));
 sg13g2_mux4_1 _9701_ (.S0(net117),
    .A0(\logix.ram_r[1798] ),
    .A1(\logix.ram_r[1806] ),
    .A2(\logix.ram_r[1814] ),
    .A3(\logix.ram_r[1822] ),
    .S1(net116),
    .X(_3704_));
 sg13g2_nand2_1 _9702_ (.Y(_3705_),
    .A(net123),
    .B(_3704_));
 sg13g2_mux4_1 _9703_ (.S0(net115),
    .A0(\logix.ram_r[1830] ),
    .A1(\logix.ram_r[1838] ),
    .A2(\logix.ram_r[1846] ),
    .A3(\logix.ram_r[1854] ),
    .S1(net167),
    .X(_3706_));
 sg13g2_nand2_1 _9704_ (.Y(_3707_),
    .A(net179),
    .B(_3706_));
 sg13g2_nand3_1 _9705_ (.B(_3705_),
    .C(_3707_),
    .A(net174),
    .Y(_3708_));
 sg13g2_nand2b_1 _9706_ (.Y(_3709_),
    .B(net113),
    .A_N(\logix.ram_r[1878] ));
 sg13g2_o21ai_1 _9707_ (.B1(_3709_),
    .Y(_3710_),
    .A1(\logix.ram_r[1862] ),
    .A2(net59));
 sg13g2_nand2b_1 _9708_ (.Y(_3711_),
    .B(net111),
    .A_N(\logix.ram_r[1886] ));
 sg13g2_o21ai_1 _9709_ (.B1(_3711_),
    .Y(_3712_),
    .A1(\logix.ram_r[1870] ),
    .A2(net58));
 sg13g2_a22oi_1 _9710_ (.Y(_3713_),
    .B1(_3712_),
    .B2(_2647_),
    .A2(_3710_),
    .A1(_2639_));
 sg13g2_mux4_1 _9711_ (.S0(net171),
    .A0(\logix.ram_r[1894] ),
    .A1(\logix.ram_r[1902] ),
    .A2(\logix.ram_r[1910] ),
    .A3(\logix.ram_r[1918] ),
    .S1(net128),
    .X(_3714_));
 sg13g2_nand2b_1 _9712_ (.Y(_3715_),
    .B(net65),
    .A_N(_3714_));
 sg13g2_nand4_1 _9713_ (.B(_3708_),
    .C(_3713_),
    .A(net79),
    .Y(_3716_),
    .D(_3715_));
 sg13g2_mux4_1 _9714_ (.S0(net139),
    .A0(\logix.ram_r[1702] ),
    .A1(\logix.ram_r[1710] ),
    .A2(\logix.ram_r[1718] ),
    .A3(\logix.ram_r[1726] ),
    .S1(net143),
    .X(_3717_));
 sg13g2_mux4_1 _9715_ (.S0(net155),
    .A0(\logix.ram_r[1670] ),
    .A1(\logix.ram_r[1678] ),
    .A2(\logix.ram_r[1686] ),
    .A3(\logix.ram_r[1694] ),
    .S1(net137),
    .X(_3718_));
 sg13g2_a22oi_1 _9716_ (.Y(_3719_),
    .B1(_3718_),
    .B2(net40),
    .A2(_3717_),
    .A1(net36));
 sg13g2_mux4_1 _9717_ (.S0(net122),
    .A0(\logix.ram_r[1766] ),
    .A1(\logix.ram_r[1774] ),
    .A2(\logix.ram_r[1782] ),
    .A3(\logix.ram_r[1790] ),
    .S1(net135),
    .X(_3720_));
 sg13g2_mux4_1 _9718_ (.S0(net134),
    .A0(\logix.ram_r[1734] ),
    .A1(\logix.ram_r[1742] ),
    .A2(\logix.ram_r[1750] ),
    .A3(\logix.ram_r[1758] ),
    .S1(net140),
    .X(_3721_));
 sg13g2_a22oi_1 _9719_ (.Y(_3722_),
    .B1(_3721_),
    .B2(net68),
    .A2(_3720_),
    .A1(net69));
 sg13g2_a21oi_1 _9720_ (.A1(_3719_),
    .A2(_3722_),
    .Y(_3723_),
    .B1(net67));
 sg13g2_nor2_1 _9721_ (.A(_2670_),
    .B(_3723_),
    .Y(_3724_));
 sg13g2_nand4_1 _9722_ (.B(_3703_),
    .C(_3716_),
    .A(_3690_),
    .Y(_3725_),
    .D(_3724_));
 sg13g2_mux4_1 _9723_ (.S0(_2664_),
    .A0(\logix.ram_r[902] ),
    .A1(\logix.ram_r[910] ),
    .A2(\logix.ram_r[918] ),
    .A3(\logix.ram_r[926] ),
    .S1(_2733_),
    .X(_3726_));
 sg13g2_nor2_1 _9724_ (.A(_2781_),
    .B(_3726_),
    .Y(_3727_));
 sg13g2_mux2_1 _9725_ (.A0(\logix.ram_r[934] ),
    .A1(\logix.ram_r[950] ),
    .S(net92),
    .X(_3728_));
 sg13g2_nor2_1 _9726_ (.A(_2344_),
    .B(_3728_),
    .Y(_3729_));
 sg13g2_mux2_1 _9727_ (.A0(\logix.ram_r[942] ),
    .A1(\logix.ram_r[958] ),
    .S(net186),
    .X(_3730_));
 sg13g2_o21ai_1 _9728_ (.B1(_2789_),
    .Y(_3731_),
    .A1(_2352_),
    .A2(_3730_));
 sg13g2_nor3_1 _9729_ (.A(_3727_),
    .B(_3729_),
    .C(_3731_),
    .Y(_3732_));
 sg13g2_mux2_1 _9730_ (.A0(\logix.ram_r[998] ),
    .A1(\logix.ram_r[1006] ),
    .S(_2616_),
    .X(_3733_));
 sg13g2_mux2_1 _9731_ (.A0(\logix.ram_r[982] ),
    .A1(\logix.ram_r[990] ),
    .S(net146),
    .X(_3734_));
 sg13g2_a22oi_1 _9732_ (.Y(_3735_),
    .B1(_3734_),
    .B2(_2742_),
    .A2(_3733_),
    .A1(net33));
 sg13g2_mux2_1 _9733_ (.A0(\logix.ram_r[966] ),
    .A1(\logix.ram_r[974] ),
    .S(_2847_),
    .X(_3736_));
 sg13g2_mux2_1 _9734_ (.A0(\logix.ram_r[1014] ),
    .A1(\logix.ram_r[1022] ),
    .S(net144),
    .X(_3737_));
 sg13g2_a22oi_1 _9735_ (.Y(_3738_),
    .B1(_3737_),
    .B2(_2700_),
    .A2(_3736_),
    .A1(_2696_));
 sg13g2_nand2_1 _9736_ (.Y(_3739_),
    .A(_3735_),
    .B(_3738_));
 sg13g2_o21ai_1 _9737_ (.B1(_2407_),
    .Y(_3740_),
    .A1(_3732_),
    .A2(_3739_));
 sg13g2_mux4_1 _9738_ (.S0(_2733_),
    .A0(\logix.ram_r[774] ),
    .A1(\logix.ram_r[790] ),
    .A2(\logix.ram_r[806] ),
    .A3(\logix.ram_r[822] ),
    .S1(_2326_),
    .X(_3741_));
 sg13g2_mux4_1 _9739_ (.S0(_2808_),
    .A0(\logix.ram_r[782] ),
    .A1(\logix.ram_r[798] ),
    .A2(\logix.ram_r[814] ),
    .A3(\logix.ram_r[830] ),
    .S1(_2326_),
    .X(_3742_));
 sg13g2_mux2_1 _9740_ (.A0(_3741_),
    .A1(_3742_),
    .S(_2935_),
    .X(_3743_));
 sg13g2_mux4_1 _9741_ (.S0(_2332_),
    .A0(\logix.ram_r[838] ),
    .A1(\logix.ram_r[846] ),
    .A2(\logix.ram_r[854] ),
    .A3(\logix.ram_r[862] ),
    .S1(_2489_),
    .X(_3744_));
 sg13g2_nor2_1 _9742_ (.A(_2380_),
    .B(_3744_),
    .Y(_3745_));
 sg13g2_mux2_1 _9743_ (.A0(\logix.ram_r[878] ),
    .A1(\logix.ram_r[894] ),
    .S(_2347_),
    .X(_3746_));
 sg13g2_nor2_1 _9744_ (.A(_2433_),
    .B(_3746_),
    .Y(_3747_));
 sg13g2_mux2_1 _9745_ (.A0(\logix.ram_r[870] ),
    .A1(\logix.ram_r[886] ),
    .S(_2355_),
    .X(_3748_));
 sg13g2_o21ai_1 _9746_ (.B1(net70),
    .Y(_3749_),
    .A1(_2439_),
    .A2(_3748_));
 sg13g2_nor3_1 _9747_ (.A(_3745_),
    .B(_3747_),
    .C(_3749_),
    .Y(_3750_));
 sg13g2_o21ai_1 _9748_ (.B1(_3750_),
    .Y(_3751_),
    .A1(_2612_),
    .A2(_3743_));
 sg13g2_mux4_1 _9749_ (.S0(_2910_),
    .A0(\logix.ram_r[678] ),
    .A1(\logix.ram_r[686] ),
    .A2(\logix.ram_r[694] ),
    .A3(\logix.ram_r[702] ),
    .S1(net114),
    .X(_3752_));
 sg13g2_mux4_1 _9750_ (.S0(net106),
    .A0(\logix.ram_r[646] ),
    .A1(\logix.ram_r[654] ),
    .A2(\logix.ram_r[662] ),
    .A3(\logix.ram_r[670] ),
    .S1(_2648_),
    .X(_3753_));
 sg13g2_a22oi_1 _9751_ (.Y(_3754_),
    .B1(_3753_),
    .B2(_3051_),
    .A2(_3752_),
    .A1(_3048_));
 sg13g2_mux4_1 _9752_ (.S0(_3013_),
    .A0(\logix.ram_r[742] ),
    .A1(\logix.ram_r[750] ),
    .A2(\logix.ram_r[758] ),
    .A3(\logix.ram_r[766] ),
    .S1(_3014_),
    .X(_3755_));
 sg13g2_mux4_1 _9753_ (.S0(_2474_),
    .A0(\logix.ram_r[710] ),
    .A1(\logix.ram_r[718] ),
    .A2(\logix.ram_r[726] ),
    .A3(\logix.ram_r[734] ),
    .S1(net156),
    .X(_3756_));
 sg13g2_a22oi_1 _9754_ (.Y(_3757_),
    .B1(_3756_),
    .B2(net84),
    .A2(_3755_),
    .A1(net62));
 sg13g2_a21oi_1 _9755_ (.A1(_3754_),
    .A2(_3757_),
    .Y(_3758_),
    .B1(net50));
 sg13g2_mux4_1 _9756_ (.S0(_2782_),
    .A0(\logix.ram_r[550] ),
    .A1(\logix.ram_r[558] ),
    .A2(\logix.ram_r[566] ),
    .A3(\logix.ram_r[574] ),
    .S1(net142),
    .X(_3759_));
 sg13g2_mux4_1 _9757_ (.S0(_2721_),
    .A0(\logix.ram_r[518] ),
    .A1(\logix.ram_r[526] ),
    .A2(\logix.ram_r[534] ),
    .A3(\logix.ram_r[542] ),
    .S1(_2489_),
    .X(_3760_));
 sg13g2_a22oi_1 _9758_ (.Y(_3761_),
    .B1(_3760_),
    .B2(_2661_),
    .A2(_3759_),
    .A1(_2658_));
 sg13g2_mux4_1 _9759_ (.S0(net94),
    .A0(\logix.ram_r[614] ),
    .A1(\logix.ram_r[622] ),
    .A2(\logix.ram_r[630] ),
    .A3(\logix.ram_r[638] ),
    .S1(_2640_),
    .X(_3762_));
 sg13g2_mux4_1 _9760_ (.S0(net161),
    .A0(\logix.ram_r[582] ),
    .A1(\logix.ram_r[590] ),
    .A2(\logix.ram_r[598] ),
    .A3(\logix.ram_r[606] ),
    .S1(_2413_),
    .X(_3763_));
 sg13g2_a22oi_1 _9761_ (.Y(_3764_),
    .B1(_3763_),
    .B2(_2667_),
    .A2(_3762_),
    .A1(_2663_));
 sg13g2_a21oi_1 _9762_ (.A1(_3761_),
    .A2(_3764_),
    .Y(_3765_),
    .B1(_2582_));
 sg13g2_nor2_1 _9763_ (.A(_3758_),
    .B(_3765_),
    .Y(_3766_));
 sg13g2_nand4_1 _9764_ (.B(_3740_),
    .C(_3751_),
    .A(_2553_),
    .Y(_3767_),
    .D(_3766_));
 sg13g2_and4_1 _9765_ (.A(_3641_),
    .B(_3683_),
    .C(_3725_),
    .D(_3767_),
    .X(net20));
 sg13g2_mux4_1 _9766_ (.S0(net115),
    .A0(\logix.ram_r[391] ),
    .A1(\logix.ram_r[399] ),
    .A2(\logix.ram_r[407] ),
    .A3(\logix.ram_r[415] ),
    .S1(net102),
    .X(_3768_));
 sg13g2_nor2_1 _9767_ (.A(net150),
    .B(_3768_),
    .Y(_3769_));
 sg13g2_mux2_1 _9768_ (.A0(\logix.ram_r[423] ),
    .A1(\logix.ram_r[439] ),
    .S(net86),
    .X(_3770_));
 sg13g2_nor2_1 _9769_ (.A(net83),
    .B(_3770_),
    .Y(_3771_));
 sg13g2_mux2_1 _9770_ (.A0(\logix.ram_r[431] ),
    .A1(\logix.ram_r[447] ),
    .S(net189),
    .X(_3772_));
 sg13g2_o21ai_1 _9771_ (.B1(net98),
    .Y(_3773_),
    .A1(net82),
    .A2(_3772_));
 sg13g2_nor3_1 _9772_ (.A(_3769_),
    .B(_3771_),
    .C(_3773_),
    .Y(_3774_));
 sg13g2_mux2_1 _9773_ (.A0(\logix.ram_r[487] ),
    .A1(\logix.ram_r[495] ),
    .S(net125),
    .X(_3775_));
 sg13g2_mux2_1 _9774_ (.A0(\logix.ram_r[471] ),
    .A1(\logix.ram_r[479] ),
    .S(net145),
    .X(_3776_));
 sg13g2_a22oi_1 _9775_ (.Y(_3777_),
    .B1(_3776_),
    .B2(net24),
    .A2(_3775_),
    .A1(net37));
 sg13g2_mux2_1 _9776_ (.A0(\logix.ram_r[455] ),
    .A1(\logix.ram_r[463] ),
    .S(_2744_),
    .X(_3778_));
 sg13g2_mux2_1 _9777_ (.A0(\logix.ram_r[503] ),
    .A1(\logix.ram_r[511] ),
    .S(net173),
    .X(_3779_));
 sg13g2_a22oi_1 _9778_ (.Y(_3780_),
    .B1(_3779_),
    .B2(net34),
    .A2(_3778_),
    .A1(net35));
 sg13g2_nand2_1 _9779_ (.Y(_3781_),
    .A(_3777_),
    .B(_3780_));
 sg13g2_o21ai_1 _9780_ (.B1(net81),
    .Y(_3782_),
    .A1(_3774_),
    .A2(_3781_));
 sg13g2_mux4_1 _9781_ (.S0(net102),
    .A0(\logix.ram_r[263] ),
    .A1(\logix.ram_r[279] ),
    .A2(\logix.ram_r[295] ),
    .A3(\logix.ram_r[311] ),
    .S1(_2414_),
    .X(_3783_));
 sg13g2_mux4_1 _9782_ (.S0(_2534_),
    .A0(\logix.ram_r[271] ),
    .A1(\logix.ram_r[287] ),
    .A2(\logix.ram_r[303] ),
    .A3(\logix.ram_r[319] ),
    .S1(net194),
    .X(_3784_));
 sg13g2_mux2_1 _9783_ (.A0(_3783_),
    .A1(_3784_),
    .S(_2421_),
    .X(_3785_));
 sg13g2_mux4_1 _9784_ (.S0(net141),
    .A0(\logix.ram_r[327] ),
    .A1(\logix.ram_r[335] ),
    .A2(\logix.ram_r[343] ),
    .A3(\logix.ram_r[351] ),
    .S1(net159),
    .X(_3786_));
 sg13g2_nor2_1 _9785_ (.A(_2423_),
    .B(_3786_),
    .Y(_3787_));
 sg13g2_mux2_1 _9786_ (.A0(\logix.ram_r[367] ),
    .A1(\logix.ram_r[383] ),
    .S(_2338_),
    .X(_3788_));
 sg13g2_nor2_1 _9787_ (.A(_2434_),
    .B(_3788_),
    .Y(_3789_));
 sg13g2_mux2_1 _9788_ (.A0(\logix.ram_r[359] ),
    .A1(\logix.ram_r[375] ),
    .S(_2640_),
    .X(_3790_));
 sg13g2_o21ai_1 _9789_ (.B1(_2547_),
    .Y(_3791_),
    .A1(_2440_),
    .A2(_3790_));
 sg13g2_nor3_1 _9790_ (.A(_3787_),
    .B(_3789_),
    .C(_3791_),
    .Y(_3792_));
 sg13g2_o21ai_1 _9791_ (.B1(_3792_),
    .Y(_3793_),
    .A1(_2412_),
    .A2(_3785_));
 sg13g2_mux4_1 _9792_ (.S0(net161),
    .A0(\logix.ram_r[167] ),
    .A1(\logix.ram_r[175] ),
    .A2(\logix.ram_r[183] ),
    .A3(\logix.ram_r[191] ),
    .S1(net168),
    .X(_3794_));
 sg13g2_mux4_1 _9793_ (.S0(net152),
    .A0(\logix.ram_r[135] ),
    .A1(\logix.ram_r[143] ),
    .A2(\logix.ram_r[151] ),
    .A3(\logix.ram_r[159] ),
    .S1(net151),
    .X(_3795_));
 sg13g2_a22oi_1 _9794_ (.Y(_3796_),
    .B1(_3795_),
    .B2(net25),
    .A2(_3794_),
    .A1(net36));
 sg13g2_mux4_1 _9795_ (.S0(net139),
    .A0(\logix.ram_r[231] ),
    .A1(\logix.ram_r[239] ),
    .A2(\logix.ram_r[247] ),
    .A3(\logix.ram_r[255] ),
    .S1(net143),
    .X(_3797_));
 sg13g2_mux4_1 _9796_ (.S0(net155),
    .A0(\logix.ram_r[199] ),
    .A1(\logix.ram_r[207] ),
    .A2(\logix.ram_r[215] ),
    .A3(\logix.ram_r[223] ),
    .S1(net137),
    .X(_3798_));
 sg13g2_a22oi_1 _9797_ (.Y(_3799_),
    .B1(_3798_),
    .B2(net68),
    .A2(_3797_),
    .A1(net76));
 sg13g2_a21oi_1 _9798_ (.A1(_3796_),
    .A2(_3799_),
    .Y(_3800_),
    .B1(net71));
 sg13g2_mux4_1 _9799_ (.S0(net178),
    .A0(\logix.ram_r[39] ),
    .A1(\logix.ram_r[47] ),
    .A2(\logix.ram_r[55] ),
    .A3(\logix.ram_r[63] ),
    .S1(_2338_),
    .X(_3801_));
 sg13g2_mux4_1 _9800_ (.S0(net160),
    .A0(\logix.ram_r[7] ),
    .A1(\logix.ram_r[15] ),
    .A2(\logix.ram_r[23] ),
    .A3(\logix.ram_r[31] ),
    .S1(net159),
    .X(_3802_));
 sg13g2_a22oi_1 _9801_ (.Y(_3803_),
    .B1(_3802_),
    .B2(net25),
    .A2(_3801_),
    .A1(net41));
 sg13g2_mux4_1 _9802_ (.S0(_2630_),
    .A0(\logix.ram_r[103] ),
    .A1(\logix.ram_r[111] ),
    .A2(\logix.ram_r[119] ),
    .A3(\logix.ram_r[127] ),
    .S1(_2631_),
    .X(_3804_));
 sg13g2_mux4_1 _9803_ (.S0(_2496_),
    .A0(\logix.ram_r[71] ),
    .A1(\logix.ram_r[79] ),
    .A2(\logix.ram_r[87] ),
    .A3(\logix.ram_r[95] ),
    .S1(net132),
    .X(_3805_));
 sg13g2_a22oi_1 _9804_ (.Y(_3806_),
    .B1(_3805_),
    .B2(net75),
    .A2(_3804_),
    .A1(_2473_));
 sg13g2_a21oi_1 _9805_ (.A1(_3803_),
    .A2(_3806_),
    .Y(_3807_),
    .B1(net74));
 sg13g2_nor2_1 _9806_ (.A(_3800_),
    .B(_3807_),
    .Y(_3808_));
 sg13g2_nand4_1 _9807_ (.B(_3782_),
    .C(_3793_),
    .A(_2456_),
    .Y(_3809_),
    .D(_3808_));
 sg13g2_mux4_1 _9808_ (.S0(_2782_),
    .A0(\logix.ram_r[903] ),
    .A1(\logix.ram_r[911] ),
    .A2(\logix.ram_r[919] ),
    .A3(\logix.ram_r[927] ),
    .S1(_2609_),
    .X(_3810_));
 sg13g2_nor2_1 _9809_ (.A(_2781_),
    .B(_3810_),
    .Y(_3811_));
 sg13g2_mux2_1 _9810_ (.A0(\logix.ram_r[935] ),
    .A1(\logix.ram_r[951] ),
    .S(net99),
    .X(_3812_));
 sg13g2_nor2_1 _9811_ (.A(_2345_),
    .B(_3812_),
    .Y(_3813_));
 sg13g2_mux2_1 _9812_ (.A0(\logix.ram_r[943] ),
    .A1(\logix.ram_r[959] ),
    .S(_2587_),
    .X(_3814_));
 sg13g2_o21ai_1 _9813_ (.B1(_2789_),
    .Y(_3815_),
    .A1(_2353_),
    .A2(_3814_));
 sg13g2_nor3_1 _9814_ (.A(_3811_),
    .B(_3813_),
    .C(_3815_),
    .Y(_3816_));
 sg13g2_mux2_1 _9815_ (.A0(\logix.ram_r[999] ),
    .A1(\logix.ram_r[1007] ),
    .S(_2744_),
    .X(_3817_));
 sg13g2_mux2_1 _9816_ (.A0(\logix.ram_r[983] ),
    .A1(\logix.ram_r[991] ),
    .S(net171),
    .X(_3818_));
 sg13g2_a22oi_1 _9817_ (.Y(_3819_),
    .B1(_3818_),
    .B2(_2742_),
    .A2(_3817_),
    .A1(_2520_));
 sg13g2_mux2_1 _9818_ (.A0(\logix.ram_r[967] ),
    .A1(\logix.ram_r[975] ),
    .S(net107),
    .X(_3820_));
 sg13g2_mux2_1 _9819_ (.A0(\logix.ram_r[1015] ),
    .A1(\logix.ram_r[1023] ),
    .S(_2586_),
    .X(_3821_));
 sg13g2_a22oi_1 _9820_ (.Y(_3822_),
    .B1(_3821_),
    .B2(_2619_),
    .A2(_3820_),
    .A1(_2614_));
 sg13g2_nand2_1 _9821_ (.Y(_3823_),
    .A(_3819_),
    .B(_3822_));
 sg13g2_o21ai_1 _9822_ (.B1(_2408_),
    .Y(_3824_),
    .A1(_3816_),
    .A2(_3823_));
 sg13g2_mux4_1 _9823_ (.S0(_2609_),
    .A0(\logix.ram_r[775] ),
    .A1(\logix.ram_r[791] ),
    .A2(\logix.ram_r[807] ),
    .A3(\logix.ram_r[823] ),
    .S1(_2800_),
    .X(_3825_));
 sg13g2_mux4_1 _9824_ (.S0(_2758_),
    .A0(\logix.ram_r[783] ),
    .A1(\logix.ram_r[799] ),
    .A2(\logix.ram_r[815] ),
    .A3(\logix.ram_r[831] ),
    .S1(_2800_),
    .X(_3826_));
 sg13g2_mux2_1 _9825_ (.A0(_3825_),
    .A1(_3826_),
    .S(net44),
    .X(_3827_));
 sg13g2_mux4_1 _9826_ (.S0(_2477_),
    .A0(\logix.ram_r[839] ),
    .A1(\logix.ram_r[847] ),
    .A2(\logix.ram_r[855] ),
    .A3(\logix.ram_r[863] ),
    .S1(net162),
    .X(_3828_));
 sg13g2_nor2_1 _9827_ (.A(net165),
    .B(_3828_),
    .Y(_3829_));
 sg13g2_mux2_1 _9828_ (.A0(\logix.ram_r[879] ),
    .A1(\logix.ram_r[895] ),
    .S(_2417_),
    .X(_3830_));
 sg13g2_nor2_1 _9829_ (.A(net43),
    .B(_3830_),
    .Y(_3831_));
 sg13g2_mux2_1 _9830_ (.A0(\logix.ram_r[871] ),
    .A1(\logix.ram_r[887] ),
    .S(_2808_),
    .X(_3832_));
 sg13g2_o21ai_1 _9831_ (.B1(_2547_),
    .Y(_3833_),
    .A1(net42),
    .A2(_3832_));
 sg13g2_nor3_1 _9832_ (.A(_3829_),
    .B(_3831_),
    .C(_3833_),
    .Y(_3834_));
 sg13g2_o21ai_1 _9833_ (.B1(_3834_),
    .Y(_3835_),
    .A1(_2412_),
    .A2(_3827_));
 sg13g2_mux4_1 _9834_ (.S0(net131),
    .A0(\logix.ram_r[679] ),
    .A1(\logix.ram_r[687] ),
    .A2(\logix.ram_r[695] ),
    .A3(\logix.ram_r[703] ),
    .S1(net138),
    .X(_3836_));
 sg13g2_mux4_1 _9835_ (.S0(_2419_),
    .A0(\logix.ram_r[647] ),
    .A1(\logix.ram_r[655] ),
    .A2(\logix.ram_r[663] ),
    .A3(\logix.ram_r[671] ),
    .S1(_2579_),
    .X(_3837_));
 sg13g2_a22oi_1 _9836_ (.Y(_3838_),
    .B1(_3837_),
    .B2(_2661_),
    .A2(_3836_),
    .A1(_2658_));
 sg13g2_mux4_1 _9837_ (.S0(_2563_),
    .A0(\logix.ram_r[743] ),
    .A1(\logix.ram_r[751] ),
    .A2(\logix.ram_r[759] ),
    .A3(\logix.ram_r[767] ),
    .S1(_2564_),
    .X(_3839_));
 sg13g2_mux4_1 _9838_ (.S0(_2712_),
    .A0(\logix.ram_r[711] ),
    .A1(\logix.ram_r[719] ),
    .A2(\logix.ram_r[727] ),
    .A3(\logix.ram_r[735] ),
    .S1(_2543_),
    .X(_3840_));
 sg13g2_a22oi_1 _9839_ (.Y(_3841_),
    .B1(_3840_),
    .B2(net61),
    .A2(_3839_),
    .A1(_2663_));
 sg13g2_a21oi_1 _9840_ (.A1(_3838_),
    .A2(_3841_),
    .Y(_3842_),
    .B1(_2570_));
 sg13g2_mux4_1 _9841_ (.S0(_2508_),
    .A0(\logix.ram_r[551] ),
    .A1(\logix.ram_r[559] ),
    .A2(\logix.ram_r[567] ),
    .A3(\logix.ram_r[575] ),
    .S1(net148),
    .X(_3843_));
 sg13g2_mux4_1 _9842_ (.S0(_2573_),
    .A0(\logix.ram_r[519] ),
    .A1(\logix.ram_r[527] ),
    .A2(\logix.ram_r[535] ),
    .A3(\logix.ram_r[543] ),
    .S1(_2574_),
    .X(_3844_));
 sg13g2_a22oi_1 _9843_ (.Y(_3845_),
    .B1(_3844_),
    .B2(_2467_),
    .A2(_3843_),
    .A1(_2554_));
 sg13g2_mux4_1 _9844_ (.S0(_2577_),
    .A0(\logix.ram_r[615] ),
    .A1(\logix.ram_r[623] ),
    .A2(\logix.ram_r[631] ),
    .A3(\logix.ram_r[639] ),
    .S1(_2537_),
    .X(_3846_));
 sg13g2_mux4_1 _9845_ (.S0(_2721_),
    .A0(\logix.ram_r[583] ),
    .A1(\logix.ram_r[591] ),
    .A2(\logix.ram_r[599] ),
    .A3(\logix.ram_r[607] ),
    .S1(_2579_),
    .X(_3847_));
 sg13g2_a22oi_1 _9846_ (.Y(_3848_),
    .B1(_3847_),
    .B2(_2568_),
    .A2(_3846_),
    .A1(_2561_));
 sg13g2_a21oi_1 _9847_ (.A1(_3845_),
    .A2(_3848_),
    .Y(_3849_),
    .B1(_2582_));
 sg13g2_nor2_1 _9848_ (.A(_3842_),
    .B(_3849_),
    .Y(_3850_));
 sg13g2_nand4_1 _9849_ (.B(_3824_),
    .C(_3835_),
    .A(_2553_),
    .Y(_3851_),
    .D(_3850_));
 sg13g2_mux4_1 _9850_ (.S0(_2521_),
    .A0(\logix.ram_r[1191] ),
    .A1(\logix.ram_r[1199] ),
    .A2(\logix.ram_r[1207] ),
    .A3(\logix.ram_r[1215] ),
    .S1(_2588_),
    .X(_3852_));
 sg13g2_mux4_1 _9851_ (.S0(net145),
    .A0(\logix.ram_r[1159] ),
    .A1(\logix.ram_r[1167] ),
    .A2(\logix.ram_r[1175] ),
    .A3(\logix.ram_r[1183] ),
    .S1(net127),
    .X(_3853_));
 sg13g2_a22oi_1 _9852_ (.Y(_3854_),
    .B1(_3853_),
    .B2(_2492_),
    .A2(_3852_),
    .A1(_2488_));
 sg13g2_mux4_1 _9853_ (.S0(_2528_),
    .A0(\logix.ram_r[1255] ),
    .A1(\logix.ram_r[1263] ),
    .A2(\logix.ram_r[1271] ),
    .A3(\logix.ram_r[1279] ),
    .S1(net124),
    .X(_3855_));
 sg13g2_mux4_1 _9854_ (.S0(_2375_),
    .A0(\logix.ram_r[1223] ),
    .A1(\logix.ram_r[1231] ),
    .A2(\logix.ram_r[1239] ),
    .A3(\logix.ram_r[1247] ),
    .S1(_2654_),
    .X(_3856_));
 sg13g2_a22oi_1 _9855_ (.Y(_3857_),
    .B1(_3856_),
    .B2(_2499_),
    .A2(_3855_),
    .A1(_2494_));
 sg13g2_a21o_1 _9856_ (.A2(_3857_),
    .A1(_3854_),
    .B1(_2503_),
    .X(_3858_));
 sg13g2_mux4_1 _9857_ (.S0(net157),
    .A0(\logix.ram_r[1287] ),
    .A1(\logix.ram_r[1295] ),
    .A2(\logix.ram_r[1303] ),
    .A3(\logix.ram_r[1311] ),
    .S1(net156),
    .X(_3859_));
 sg13g2_nand2_1 _9858_ (.Y(_3860_),
    .A(net95),
    .B(_3859_));
 sg13g2_mux4_1 _9859_ (.S0(net122),
    .A0(\logix.ram_r[1319] ),
    .A1(\logix.ram_r[1327] ),
    .A2(\logix.ram_r[1335] ),
    .A3(\logix.ram_r[1343] ),
    .S1(net121),
    .X(_3861_));
 sg13g2_nand2_1 _9860_ (.Y(_3862_),
    .A(net150),
    .B(_3861_));
 sg13g2_a21oi_1 _9861_ (.A1(_3860_),
    .A2(_3862_),
    .Y(_3863_),
    .B1(_2411_));
 sg13g2_mux2_1 _9862_ (.A0(\logix.ram_r[1351] ),
    .A1(\logix.ram_r[1359] ),
    .S(net119),
    .X(_3864_));
 sg13g2_mux2_1 _9863_ (.A0(\logix.ram_r[1399] ),
    .A1(\logix.ram_r[1407] ),
    .S(net129),
    .X(_3865_));
 sg13g2_a22oi_1 _9864_ (.Y(_3866_),
    .B1(_3865_),
    .B2(net26),
    .A2(_3864_),
    .A1(net27));
 sg13g2_mux2_1 _9865_ (.A0(\logix.ram_r[1383] ),
    .A1(\logix.ram_r[1391] ),
    .S(net96),
    .X(_3867_));
 sg13g2_mux2_1 _9866_ (.A0(\logix.ram_r[1367] ),
    .A1(\logix.ram_r[1375] ),
    .S(net144),
    .X(_3868_));
 sg13g2_a22oi_1 _9867_ (.Y(_3869_),
    .B1(_3868_),
    .B2(net32),
    .A2(_3867_),
    .A1(net33));
 sg13g2_nand2_1 _9868_ (.Y(_3870_),
    .A(_3866_),
    .B(_3869_));
 sg13g2_o21ai_1 _9869_ (.B1(net79),
    .Y(_3871_),
    .A1(_3863_),
    .A2(_3870_));
 sg13g2_mux4_1 _9870_ (.S0(net117),
    .A0(\logix.ram_r[1415] ),
    .A1(\logix.ram_r[1423] ),
    .A2(\logix.ram_r[1431] ),
    .A3(\logix.ram_r[1439] ),
    .S1(net116),
    .X(_3872_));
 sg13g2_nand2_1 _9871_ (.Y(_3873_),
    .A(_2605_),
    .B(_3872_));
 sg13g2_mux4_1 _9872_ (.S0(_2634_),
    .A0(\logix.ram_r[1447] ),
    .A1(\logix.ram_r[1455] ),
    .A2(\logix.ram_r[1463] ),
    .A3(\logix.ram_r[1471] ),
    .S1(net167),
    .X(_3874_));
 sg13g2_nand2_1 _9873_ (.Y(_3875_),
    .A(_2327_),
    .B(_3874_));
 sg13g2_nand3_1 _9874_ (.B(_3873_),
    .C(_3875_),
    .A(_2363_),
    .Y(_3876_));
 sg13g2_nand2b_1 _9875_ (.Y(_3877_),
    .B(net113),
    .A_N(\logix.ram_r[1495] ));
 sg13g2_o21ai_1 _9876_ (.B1(_3877_),
    .Y(_3878_),
    .A1(\logix.ram_r[1479] ),
    .A2(_2687_));
 sg13g2_nand2b_1 _9877_ (.Y(_3879_),
    .B(net111),
    .A_N(\logix.ram_r[1503] ));
 sg13g2_o21ai_1 _9878_ (.B1(_3879_),
    .Y(_3880_),
    .A1(\logix.ram_r[1487] ),
    .A2(net58));
 sg13g2_a22oi_1 _9879_ (.Y(_3881_),
    .B1(_3880_),
    .B2(_2647_),
    .A2(_3878_),
    .A1(_2639_));
 sg13g2_mux4_1 _9880_ (.S0(_2392_),
    .A0(\logix.ram_r[1511] ),
    .A1(\logix.ram_r[1519] ),
    .A2(\logix.ram_r[1527] ),
    .A3(\logix.ram_r[1535] ),
    .S1(net128),
    .X(_3882_));
 sg13g2_nand2b_1 _9881_ (.Y(_3883_),
    .B(net65),
    .A_N(_3882_));
 sg13g2_nand4_1 _9882_ (.B(_3876_),
    .C(_3881_),
    .A(net170),
    .Y(_3884_),
    .D(_3883_));
 sg13g2_mux4_1 _9883_ (.S0(net139),
    .A0(\logix.ram_r[1063] ),
    .A1(\logix.ram_r[1071] ),
    .A2(\logix.ram_r[1079] ),
    .A3(\logix.ram_r[1087] ),
    .S1(_2556_),
    .X(_3885_));
 sg13g2_mux4_1 _9884_ (.S0(_2419_),
    .A0(\logix.ram_r[1031] ),
    .A1(\logix.ram_r[1039] ),
    .A2(\logix.ram_r[1047] ),
    .A3(\logix.ram_r[1055] ),
    .S1(_2558_),
    .X(_3886_));
 sg13g2_a22oi_1 _9885_ (.Y(_3887_),
    .B1(_3886_),
    .B2(_2467_),
    .A2(_3885_),
    .A1(_2554_));
 sg13g2_mux4_1 _9886_ (.S0(_2608_),
    .A0(\logix.ram_r[1127] ),
    .A1(\logix.ram_r[1135] ),
    .A2(\logix.ram_r[1143] ),
    .A3(\logix.ram_r[1151] ),
    .S1(_2564_),
    .X(_3888_));
 sg13g2_mux4_1 _9887_ (.S0(net134),
    .A0(\logix.ram_r[1095] ),
    .A1(\logix.ram_r[1103] ),
    .A2(\logix.ram_r[1111] ),
    .A3(\logix.ram_r[1119] ),
    .S1(net140),
    .X(_3889_));
 sg13g2_a22oi_1 _9888_ (.Y(_3890_),
    .B1(_3889_),
    .B2(_2568_),
    .A2(_3888_),
    .A1(net69));
 sg13g2_a21oi_1 _9889_ (.A1(_3887_),
    .A2(_3890_),
    .Y(_3891_),
    .B1(net66));
 sg13g2_nor2_1 _9890_ (.A(_2705_),
    .B(_3891_),
    .Y(_3892_));
 sg13g2_nand4_1 _9891_ (.B(_3871_),
    .C(_3884_),
    .A(_3858_),
    .Y(_3893_),
    .D(_3892_));
 sg13g2_mux4_1 _9892_ (.S0(net109),
    .A0(\logix.ram_r[1927] ),
    .A1(\logix.ram_r[1935] ),
    .A2(\logix.ram_r[1943] ),
    .A3(\logix.ram_r[1951] ),
    .S1(net104),
    .X(_3894_));
 sg13g2_nor2_1 _9893_ (.A(net188),
    .B(_3894_),
    .Y(_3895_));
 sg13g2_mux2_1 _9894_ (.A0(\logix.ram_r[1959] ),
    .A1(\logix.ram_r[1975] ),
    .S(net92),
    .X(_3896_));
 sg13g2_nor2_1 _9895_ (.A(_2344_),
    .B(_3896_),
    .Y(_3897_));
 sg13g2_mux2_1 _9896_ (.A0(\logix.ram_r[1967] ),
    .A1(\logix.ram_r[1983] ),
    .S(net186),
    .X(_3898_));
 sg13g2_o21ai_1 _9897_ (.B1(net98),
    .Y(_3899_),
    .A1(_2352_),
    .A2(_3898_));
 sg13g2_nor3_1 _9898_ (.A(_3895_),
    .B(_3897_),
    .C(_3899_),
    .Y(_3900_));
 sg13g2_mux2_1 _9899_ (.A0(\logix.ram_r[2023] ),
    .A1(\logix.ram_r[2031] ),
    .S(net119),
    .X(_3901_));
 sg13g2_mux2_1 _9900_ (.A0(\logix.ram_r[2007] ),
    .A1(\logix.ram_r[2015] ),
    .S(net146),
    .X(_3902_));
 sg13g2_a22oi_1 _9901_ (.Y(_3903_),
    .B1(_3902_),
    .B2(net32),
    .A2(_3901_),
    .A1(net33));
 sg13g2_mux2_1 _9902_ (.A0(\logix.ram_r[1991] ),
    .A1(\logix.ram_r[1999] ),
    .S(net96),
    .X(_3904_));
 sg13g2_mux2_1 _9903_ (.A0(\logix.ram_r[2039] ),
    .A1(\logix.ram_r[2047] ),
    .S(net103),
    .X(_3905_));
 sg13g2_a22oi_1 _9904_ (.Y(_3906_),
    .B1(_3905_),
    .B2(net26),
    .A2(_3904_),
    .A1(net27));
 sg13g2_nand2_1 _9905_ (.Y(_3907_),
    .A(_3903_),
    .B(_3906_));
 sg13g2_o21ai_1 _9906_ (.B1(net170),
    .Y(_3908_),
    .A1(_3900_),
    .A2(_3907_));
 sg13g2_mux4_1 _9907_ (.S0(net104),
    .A0(\logix.ram_r[1799] ),
    .A1(\logix.ram_r[1815] ),
    .A2(\logix.ram_r[1831] ),
    .A3(\logix.ram_r[1847] ),
    .S1(net204),
    .X(_3909_));
 sg13g2_mux4_1 _9908_ (.S0(net97),
    .A0(\logix.ram_r[1807] ),
    .A1(\logix.ram_r[1823] ),
    .A2(\logix.ram_r[1839] ),
    .A3(\logix.ram_r[1855] ),
    .S1(net204),
    .X(_3910_));
 sg13g2_mux2_1 _9909_ (.A0(_3909_),
    .A1(_3910_),
    .S(net57),
    .X(_3911_));
 sg13g2_mux4_1 _9910_ (.S0(net178),
    .A0(\logix.ram_r[1863] ),
    .A1(\logix.ram_r[1871] ),
    .A2(\logix.ram_r[1879] ),
    .A3(\logix.ram_r[1887] ),
    .S1(net153),
    .X(_3912_));
 sg13g2_nor2_1 _9911_ (.A(net202),
    .B(_3912_),
    .Y(_3913_));
 sg13g2_mux2_1 _9912_ (.A0(\logix.ram_r[1903] ),
    .A1(\logix.ram_r[1919] ),
    .S(net176),
    .X(_3914_));
 sg13g2_nor2_1 _9913_ (.A(_2433_),
    .B(_3914_),
    .Y(_3915_));
 sg13g2_mux2_1 _9914_ (.A0(\logix.ram_r[1895] ),
    .A1(\logix.ram_r[1911] ),
    .S(net175),
    .X(_3916_));
 sg13g2_o21ai_1 _9915_ (.B1(net70),
    .Y(_3917_),
    .A1(_2439_),
    .A2(_3916_));
 sg13g2_nor3_1 _9916_ (.A(_3913_),
    .B(_3915_),
    .C(_3917_),
    .Y(_3918_));
 sg13g2_o21ai_1 _9917_ (.B1(_3918_),
    .Y(_3919_),
    .A1(net120),
    .A2(_3911_));
 sg13g2_mux4_1 _9918_ (.S0(net94),
    .A0(\logix.ram_r[1703] ),
    .A1(\logix.ram_r[1711] ),
    .A2(\logix.ram_r[1719] ),
    .A3(\logix.ram_r[1727] ),
    .S1(net114),
    .X(_3920_));
 sg13g2_mux4_1 _9919_ (.S0(net106),
    .A0(\logix.ram_r[1671] ),
    .A1(\logix.ram_r[1679] ),
    .A2(\logix.ram_r[1687] ),
    .A3(\logix.ram_r[1695] ),
    .S1(net112),
    .X(_3921_));
 sg13g2_a22oi_1 _9920_ (.Y(_3922_),
    .B1(_3921_),
    .B2(net22),
    .A2(_3920_),
    .A1(net23));
 sg13g2_mux4_1 _9921_ (.S0(net87),
    .A0(\logix.ram_r[1767] ),
    .A1(\logix.ram_r[1775] ),
    .A2(\logix.ram_r[1783] ),
    .A3(\logix.ram_r[1791] ),
    .S1(net97),
    .X(_3923_));
 sg13g2_mux4_1 _9922_ (.S0(net157),
    .A0(\logix.ram_r[1735] ),
    .A1(\logix.ram_r[1743] ),
    .A2(\logix.ram_r[1751] ),
    .A3(\logix.ram_r[1759] ),
    .S1(net156),
    .X(_3924_));
 sg13g2_a22oi_1 _9923_ (.Y(_3925_),
    .B1(_3924_),
    .B2(net84),
    .A2(_3923_),
    .A1(net85));
 sg13g2_a21oi_1 _9924_ (.A1(_3922_),
    .A2(_3925_),
    .Y(_3926_),
    .B1(net50));
 sg13g2_mux4_1 _9925_ (.S0(net100),
    .A0(\logix.ram_r[1575] ),
    .A1(\logix.ram_r[1583] ),
    .A2(\logix.ram_r[1591] ),
    .A3(\logix.ram_r[1599] ),
    .S1(net142),
    .X(_3927_));
 sg13g2_mux4_1 _9926_ (.S0(net105),
    .A0(\logix.ram_r[1543] ),
    .A1(\logix.ram_r[1551] ),
    .A2(\logix.ram_r[1559] ),
    .A3(\logix.ram_r[1567] ),
    .S1(net153),
    .X(_3928_));
 sg13g2_a22oi_1 _9927_ (.Y(_3929_),
    .B1(_3928_),
    .B2(net30),
    .A2(_3927_),
    .A1(net31));
 sg13g2_mux4_1 _9928_ (.S0(net94),
    .A0(\logix.ram_r[1639] ),
    .A1(\logix.ram_r[1647] ),
    .A2(\logix.ram_r[1655] ),
    .A3(\logix.ram_r[1663] ),
    .S1(net114),
    .X(_3930_));
 sg13g2_mux4_1 _9929_ (.S0(net161),
    .A0(\logix.ram_r[1607] ),
    .A1(\logix.ram_r[1615] ),
    .A2(\logix.ram_r[1623] ),
    .A3(\logix.ram_r[1631] ),
    .S1(net168),
    .X(_3931_));
 sg13g2_a22oi_1 _9930_ (.Y(_3932_),
    .B1(_3931_),
    .B2(net61),
    .A2(_3930_),
    .A1(net62));
 sg13g2_a21oi_1 _9931_ (.A1(_3929_),
    .A2(_3932_),
    .Y(_3933_),
    .B1(net66));
 sg13g2_nor2_1 _9932_ (.A(_3926_),
    .B(_3933_),
    .Y(_3934_));
 sg13g2_nand4_1 _9933_ (.B(_3908_),
    .C(_3919_),
    .A(_2780_),
    .Y(_3935_),
    .D(_3934_));
 sg13g2_and4_1 _9934_ (.A(_3809_),
    .B(_3851_),
    .C(_3893_),
    .D(_3935_),
    .X(net21));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_tiehi _9942__787 (.L_HI(net787));
 sg13g2_buf_1 _9937_ (.A(net777),
    .X(uio_oe[0]));
 sg13g2_buf_1 _9938_ (.A(net778),
    .X(uio_oe[1]));
 sg13g2_buf_1 _9939_ (.A(net779),
    .X(uio_oe[2]));
 sg13g2_buf_1 _9940_ (.A(net780),
    .X(uio_oe[3]));
 sg13g2_buf_1 _9941_ (.A(net781),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9942_ (.A(net787),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9943_ (.A(net788),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9944_ (.A(net789),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9945_ (.A(net782),
    .X(uio_out[0]));
 sg13g2_buf_1 _9946_ (.A(net783),
    .X(uio_out[1]));
 sg13g2_buf_1 _9947_ (.A(net784),
    .X(uio_out[2]));
 sg13g2_buf_1 _9948_ (.A(net785),
    .X(uio_out[3]));
 sg13g2_buf_1 _9949_ (.A(net786),
    .X(uio_out[4]));
 sg13g2_dfrbp_1 \logix.feedback_r[0]$_DFF_P_  (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net790),
    .D(net14),
    .Q_N(_5992_),
    .Q(\logix.feedback_r[0] ));
 sg13g2_dfrbp_1 \logix.feedback_r[1]$_DFF_P_  (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net791),
    .D(net15),
    .Q_N(_0000_),
    .Q(\logix.feedback_r[1] ));
 sg13g2_dfrbp_1 \logix.feedback_r[2]$_DFF_P_  (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net792),
    .D(net16),
    .Q_N(_0001_),
    .Q(\logix.feedback_r[2] ));
 sg13g2_dfrbp_1 \logix.feedback_r[3]$_DFF_P_  (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net793),
    .D(net17),
    .Q_N(_0002_),
    .Q(\logix.feedback_r[3] ));
 sg13g2_dfrbp_1 \logix.feedback_r[4]$_DFF_P_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net794),
    .D(net18),
    .Q_N(_0003_),
    .Q(\logix.feedback_r[4] ));
 sg13g2_dfrbp_1 \logix.feedback_r[5]$_DFF_P_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net795),
    .D(net19),
    .Q_N(_0004_),
    .Q(\logix.feedback_r[5] ));
 sg13g2_dfrbp_1 \logix.feedback_r[6]$_DFF_P_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net796),
    .D(net20),
    .Q_N(_0005_),
    .Q(\logix.feedback_r[6] ));
 sg13g2_dfrbp_1 \logix.feedback_r[7]$_DFF_P_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net797),
    .D(net21),
    .Q_N(_0006_),
    .Q(\logix.feedback_r[7] ));
 sg13g2_dfrbp_1 \logix.ram_r[0]$_DFFE_PP_  (.CLK(net576),
    .RESET_B(net798),
    .D(_0007_),
    .Q_N(_5991_),
    .Q(\logix.ram_r[0] ));
 sg13g2_dfrbp_1 \logix.ram_r[1000]$_DFFE_PP_  (.CLK(net576),
    .RESET_B(net799),
    .D(_0008_),
    .Q_N(_5990_),
    .Q(\logix.ram_r[1000] ));
 sg13g2_dfrbp_1 \logix.ram_r[1001]$_DFFE_PP_  (.CLK(net576),
    .RESET_B(net800),
    .D(_0009_),
    .Q_N(_5989_),
    .Q(\logix.ram_r[1001] ));
 sg13g2_dfrbp_1 \logix.ram_r[1002]$_DFFE_PP_  (.CLK(net575),
    .RESET_B(net801),
    .D(_0010_),
    .Q_N(_5988_),
    .Q(\logix.ram_r[1002] ));
 sg13g2_dfrbp_1 \logix.ram_r[1003]$_DFFE_PP_  (.CLK(net575),
    .RESET_B(net802),
    .D(_0011_),
    .Q_N(_5987_),
    .Q(\logix.ram_r[1003] ));
 sg13g2_dfrbp_1 \logix.ram_r[1004]$_DFFE_PP_  (.CLK(net634),
    .RESET_B(net803),
    .D(_0012_),
    .Q_N(_5986_),
    .Q(\logix.ram_r[1004] ));
 sg13g2_dfrbp_1 \logix.ram_r[1005]$_DFFE_PP_  (.CLK(net576),
    .RESET_B(net804),
    .D(_0013_),
    .Q_N(_5985_),
    .Q(\logix.ram_r[1005] ));
 sg13g2_dfrbp_1 \logix.ram_r[1006]$_DFFE_PP_  (.CLK(net576),
    .RESET_B(net805),
    .D(_0014_),
    .Q_N(_5984_),
    .Q(\logix.ram_r[1006] ));
 sg13g2_dfrbp_1 \logix.ram_r[1007]$_DFFE_PP_  (.CLK(net576),
    .RESET_B(net806),
    .D(_0015_),
    .Q_N(_5983_),
    .Q(\logix.ram_r[1007] ));
 sg13g2_dfrbp_1 \logix.ram_r[1008]$_DFFE_PP_  (.CLK(net636),
    .RESET_B(net807),
    .D(_0016_),
    .Q_N(_5982_),
    .Q(\logix.ram_r[1008] ));
 sg13g2_dfrbp_1 \logix.ram_r[1009]$_DFFE_PP_  (.CLK(net641),
    .RESET_B(net808),
    .D(_0017_),
    .Q_N(_5981_),
    .Q(\logix.ram_r[1009] ));
 sg13g2_dfrbp_1 \logix.ram_r[100]$_DFFE_PP_  (.CLK(net694),
    .RESET_B(net809),
    .D(_0018_),
    .Q_N(_5980_),
    .Q(\logix.ram_r[100] ));
 sg13g2_dfrbp_1 \logix.ram_r[1010]$_DFFE_PP_  (.CLK(net641),
    .RESET_B(net810),
    .D(_0019_),
    .Q_N(_5979_),
    .Q(\logix.ram_r[1010] ));
 sg13g2_dfrbp_1 \logix.ram_r[1011]$_DFFE_PP_  (.CLK(net639),
    .RESET_B(net811),
    .D(_0020_),
    .Q_N(_5978_),
    .Q(\logix.ram_r[1011] ));
 sg13g2_dfrbp_1 \logix.ram_r[1012]$_DFFE_PP_  (.CLK(net639),
    .RESET_B(net812),
    .D(_0021_),
    .Q_N(_5977_),
    .Q(\logix.ram_r[1012] ));
 sg13g2_dfrbp_1 \logix.ram_r[1013]$_DFFE_PP_  (.CLK(net642),
    .RESET_B(net813),
    .D(_0022_),
    .Q_N(_5976_),
    .Q(\logix.ram_r[1013] ));
 sg13g2_dfrbp_1 \logix.ram_r[1014]$_DFFE_PP_  (.CLK(net659),
    .RESET_B(net814),
    .D(_0023_),
    .Q_N(_5975_),
    .Q(\logix.ram_r[1014] ));
 sg13g2_dfrbp_1 \logix.ram_r[1015]$_DFFE_PP_  (.CLK(net642),
    .RESET_B(net815),
    .D(_0024_),
    .Q_N(_5974_),
    .Q(\logix.ram_r[1015] ));
 sg13g2_dfrbp_1 \logix.ram_r[1016]$_DFFE_PP_  (.CLK(net642),
    .RESET_B(net816),
    .D(_0025_),
    .Q_N(_5973_),
    .Q(\logix.ram_r[1016] ));
 sg13g2_dfrbp_1 \logix.ram_r[1017]$_DFFE_PP_  (.CLK(net641),
    .RESET_B(net817),
    .D(_0026_),
    .Q_N(_5972_),
    .Q(\logix.ram_r[1017] ));
 sg13g2_dfrbp_1 \logix.ram_r[1018]$_DFFE_PP_  (.CLK(net641),
    .RESET_B(net818),
    .D(_0027_),
    .Q_N(_5971_),
    .Q(\logix.ram_r[1018] ));
 sg13g2_dfrbp_1 \logix.ram_r[1019]$_DFFE_PP_  (.CLK(net639),
    .RESET_B(net819),
    .D(_0028_),
    .Q_N(_5970_),
    .Q(\logix.ram_r[1019] ));
 sg13g2_dfrbp_1 \logix.ram_r[101]$_DFFE_PP_  (.CLK(net695),
    .RESET_B(net820),
    .D(_0029_),
    .Q_N(_5969_),
    .Q(\logix.ram_r[101] ));
 sg13g2_dfrbp_1 \logix.ram_r[1020]$_DFFE_PP_  (.CLK(net640),
    .RESET_B(net821),
    .D(_0030_),
    .Q_N(_5968_),
    .Q(\logix.ram_r[1020] ));
 sg13g2_dfrbp_1 \logix.ram_r[1021]$_DFFE_PP_  (.CLK(net642),
    .RESET_B(net822),
    .D(_0031_),
    .Q_N(_5967_),
    .Q(\logix.ram_r[1021] ));
 sg13g2_dfrbp_1 \logix.ram_r[1022]$_DFFE_PP_  (.CLK(net659),
    .RESET_B(net823),
    .D(_0032_),
    .Q_N(_5966_),
    .Q(\logix.ram_r[1022] ));
 sg13g2_dfrbp_1 \logix.ram_r[1023]$_DFFE_PP_  (.CLK(net660),
    .RESET_B(net824),
    .D(_0033_),
    .Q_N(_5965_),
    .Q(\logix.ram_r[1023] ));
 sg13g2_dfrbp_1 \logix.ram_r[1024]$_DFFE_PP_  (.CLK(net693),
    .RESET_B(net825),
    .D(_0034_),
    .Q_N(_5964_),
    .Q(\logix.ram_r[1024] ));
 sg13g2_dfrbp_1 \logix.ram_r[1025]$_DFFE_PP_  (.CLK(net693),
    .RESET_B(net826),
    .D(_0035_),
    .Q_N(_5963_),
    .Q(\logix.ram_r[1025] ));
 sg13g2_dfrbp_1 \logix.ram_r[1026]$_DFFE_PP_  (.CLK(net693),
    .RESET_B(net827),
    .D(_0036_),
    .Q_N(_5962_),
    .Q(\logix.ram_r[1026] ));
 sg13g2_dfrbp_1 \logix.ram_r[1027]$_DFFE_PP_  (.CLK(net684),
    .RESET_B(net828),
    .D(_0037_),
    .Q_N(_5961_),
    .Q(\logix.ram_r[1027] ));
 sg13g2_dfrbp_1 \logix.ram_r[1028]$_DFFE_PP_  (.CLK(net684),
    .RESET_B(net829),
    .D(_0038_),
    .Q_N(_5960_),
    .Q(\logix.ram_r[1028] ));
 sg13g2_dfrbp_1 \logix.ram_r[1029]$_DFFE_PP_  (.CLK(net690),
    .RESET_B(net830),
    .D(_0039_),
    .Q_N(_5959_),
    .Q(\logix.ram_r[1029] ));
 sg13g2_dfrbp_1 \logix.ram_r[102]$_DFFE_PP_  (.CLK(net693),
    .RESET_B(net831),
    .D(_0040_),
    .Q_N(_5958_),
    .Q(\logix.ram_r[102] ));
 sg13g2_dfrbp_1 \logix.ram_r[1030]$_DFFE_PP_  (.CLK(net690),
    .RESET_B(net832),
    .D(_0041_),
    .Q_N(_5957_),
    .Q(\logix.ram_r[1030] ));
 sg13g2_dfrbp_1 \logix.ram_r[1031]$_DFFE_PP_  (.CLK(net689),
    .RESET_B(net833),
    .D(_0042_),
    .Q_N(_5956_),
    .Q(\logix.ram_r[1031] ));
 sg13g2_dfrbp_1 \logix.ram_r[1032]$_DFFE_PP_  (.CLK(net684),
    .RESET_B(net834),
    .D(_0043_),
    .Q_N(_5955_),
    .Q(\logix.ram_r[1032] ));
 sg13g2_dfrbp_1 \logix.ram_r[1033]$_DFFE_PP_  (.CLK(net684),
    .RESET_B(net835),
    .D(_0044_),
    .Q_N(_5954_),
    .Q(\logix.ram_r[1033] ));
 sg13g2_dfrbp_1 \logix.ram_r[1034]$_DFFE_PP_  (.CLK(net684),
    .RESET_B(net836),
    .D(_0045_),
    .Q_N(_5953_),
    .Q(\logix.ram_r[1034] ));
 sg13g2_dfrbp_1 \logix.ram_r[1035]$_DFFE_PP_  (.CLK(net684),
    .RESET_B(net837),
    .D(_0046_),
    .Q_N(_5952_),
    .Q(\logix.ram_r[1035] ));
 sg13g2_dfrbp_1 \logix.ram_r[1036]$_DFFE_PP_  (.CLK(net689),
    .RESET_B(net838),
    .D(_0047_),
    .Q_N(_5951_),
    .Q(\logix.ram_r[1036] ));
 sg13g2_dfrbp_1 \logix.ram_r[1037]$_DFFE_PP_  (.CLK(net690),
    .RESET_B(net839),
    .D(_0048_),
    .Q_N(_5950_),
    .Q(\logix.ram_r[1037] ));
 sg13g2_dfrbp_1 \logix.ram_r[1038]$_DFFE_PP_  (.CLK(net690),
    .RESET_B(net840),
    .D(_0049_),
    .Q_N(_5949_),
    .Q(\logix.ram_r[1038] ));
 sg13g2_dfrbp_1 \logix.ram_r[1039]$_DFFE_PP_  (.CLK(net689),
    .RESET_B(net841),
    .D(_0050_),
    .Q_N(_5948_),
    .Q(\logix.ram_r[1039] ));
 sg13g2_dfrbp_1 \logix.ram_r[103]$_DFFE_PP_  (.CLK(net697),
    .RESET_B(net842),
    .D(_0051_),
    .Q_N(_5947_),
    .Q(\logix.ram_r[103] ));
 sg13g2_dfrbp_1 \logix.ram_r[1040]$_DFFE_PP_  (.CLK(net689),
    .RESET_B(net843),
    .D(_0052_),
    .Q_N(_5946_),
    .Q(\logix.ram_r[1040] ));
 sg13g2_dfrbp_1 \logix.ram_r[1041]$_DFFE_PP_  (.CLK(net685),
    .RESET_B(net844),
    .D(_0053_),
    .Q_N(_5945_),
    .Q(\logix.ram_r[1041] ));
 sg13g2_dfrbp_1 \logix.ram_r[1042]$_DFFE_PP_  (.CLK(net685),
    .RESET_B(net845),
    .D(_0054_),
    .Q_N(_5944_),
    .Q(\logix.ram_r[1042] ));
 sg13g2_dfrbp_1 \logix.ram_r[1043]$_DFFE_PP_  (.CLK(net689),
    .RESET_B(net846),
    .D(_0055_),
    .Q_N(_5943_),
    .Q(\logix.ram_r[1043] ));
 sg13g2_dfrbp_1 \logix.ram_r[1044]$_DFFE_PP_  (.CLK(net690),
    .RESET_B(net847),
    .D(_0056_),
    .Q_N(_5942_),
    .Q(\logix.ram_r[1044] ));
 sg13g2_dfrbp_1 \logix.ram_r[1045]$_DFFE_PP_  (.CLK(net706),
    .RESET_B(net848),
    .D(_0057_),
    .Q_N(_5941_),
    .Q(\logix.ram_r[1045] ));
 sg13g2_dfrbp_1 \logix.ram_r[1046]$_DFFE_PP_  (.CLK(net690),
    .RESET_B(net849),
    .D(_0058_),
    .Q_N(_5940_),
    .Q(\logix.ram_r[1046] ));
 sg13g2_dfrbp_1 \logix.ram_r[1047]$_DFFE_PP_  (.CLK(net691),
    .RESET_B(net850),
    .D(_0059_),
    .Q_N(_5939_),
    .Q(\logix.ram_r[1047] ));
 sg13g2_dfrbp_1 \logix.ram_r[1048]$_DFFE_PP_  (.CLK(net689),
    .RESET_B(net851),
    .D(_0060_),
    .Q_N(_5938_),
    .Q(\logix.ram_r[1048] ));
 sg13g2_dfrbp_1 \logix.ram_r[1049]$_DFFE_PP_  (.CLK(net690),
    .RESET_B(net852),
    .D(_0061_),
    .Q_N(_5937_),
    .Q(\logix.ram_r[1049] ));
 sg13g2_dfrbp_1 \logix.ram_r[104]$_DFFE_PP_  (.CLK(net697),
    .RESET_B(net853),
    .D(_0062_),
    .Q_N(_5936_),
    .Q(\logix.ram_r[104] ));
 sg13g2_dfrbp_1 \logix.ram_r[1050]$_DFFE_PP_  (.CLK(net689),
    .RESET_B(net854),
    .D(_0063_),
    .Q_N(_5935_),
    .Q(\logix.ram_r[1050] ));
 sg13g2_dfrbp_1 \logix.ram_r[1051]$_DFFE_PP_  (.CLK(net689),
    .RESET_B(net855),
    .D(_0064_),
    .Q_N(_5934_),
    .Q(\logix.ram_r[1051] ));
 sg13g2_dfrbp_1 \logix.ram_r[1052]$_DFFE_PP_  (.CLK(net691),
    .RESET_B(net856),
    .D(_0065_),
    .Q_N(_5933_),
    .Q(\logix.ram_r[1052] ));
 sg13g2_dfrbp_1 \logix.ram_r[1053]$_DFFE_PP_  (.CLK(net706),
    .RESET_B(net857),
    .D(_0066_),
    .Q_N(_5932_),
    .Q(\logix.ram_r[1053] ));
 sg13g2_dfrbp_1 \logix.ram_r[1054]$_DFFE_PP_  (.CLK(net706),
    .RESET_B(net858),
    .D(_0067_),
    .Q_N(_5931_),
    .Q(\logix.ram_r[1054] ));
 sg13g2_dfrbp_1 \logix.ram_r[1055]$_DFFE_PP_  (.CLK(net706),
    .RESET_B(net859),
    .D(_0068_),
    .Q_N(_5930_),
    .Q(\logix.ram_r[1055] ));
 sg13g2_dfrbp_1 \logix.ram_r[1056]$_DFFE_PP_  (.CLK(net706),
    .RESET_B(net860),
    .D(_0069_),
    .Q_N(_5929_),
    .Q(\logix.ram_r[1056] ));
 sg13g2_dfrbp_1 \logix.ram_r[1057]$_DFFE_PP_  (.CLK(net715),
    .RESET_B(net861),
    .D(_0070_),
    .Q_N(_5928_),
    .Q(\logix.ram_r[1057] ));
 sg13g2_dfrbp_1 \logix.ram_r[1058]$_DFFE_PP_  (.CLK(net710),
    .RESET_B(net862),
    .D(_0071_),
    .Q_N(_5927_),
    .Q(\logix.ram_r[1058] ));
 sg13g2_dfrbp_1 \logix.ram_r[1059]$_DFFE_PP_  (.CLK(net710),
    .RESET_B(net863),
    .D(_0072_),
    .Q_N(_5926_),
    .Q(\logix.ram_r[1059] ));
 sg13g2_dfrbp_1 \logix.ram_r[105]$_DFFE_PP_  (.CLK(net716),
    .RESET_B(net864),
    .D(_0073_),
    .Q_N(_5925_),
    .Q(\logix.ram_r[105] ));
 sg13g2_dfrbp_1 \logix.ram_r[1060]$_DFFE_PP_  (.CLK(net710),
    .RESET_B(net865),
    .D(_0074_),
    .Q_N(_5924_),
    .Q(\logix.ram_r[1060] ));
 sg13g2_dfrbp_1 \logix.ram_r[1061]$_DFFE_PP_  (.CLK(net710),
    .RESET_B(net866),
    .D(_0075_),
    .Q_N(_5923_),
    .Q(\logix.ram_r[1061] ));
 sg13g2_dfrbp_1 \logix.ram_r[1062]$_DFFE_PP_  (.CLK(net706),
    .RESET_B(net867),
    .D(_0076_),
    .Q_N(_5922_),
    .Q(\logix.ram_r[1062] ));
 sg13g2_dfrbp_1 \logix.ram_r[1063]$_DFFE_PP_  (.CLK(net706),
    .RESET_B(net868),
    .D(_0077_),
    .Q_N(_5921_),
    .Q(\logix.ram_r[1063] ));
 sg13g2_dfrbp_1 \logix.ram_r[1064]$_DFFE_PP_  (.CLK(net715),
    .RESET_B(net869),
    .D(_0078_),
    .Q_N(_5920_),
    .Q(\logix.ram_r[1064] ));
 sg13g2_dfrbp_1 \logix.ram_r[1065]$_DFFE_PP_  (.CLK(net719),
    .RESET_B(net870),
    .D(_0079_),
    .Q_N(_5919_),
    .Q(\logix.ram_r[1065] ));
 sg13g2_dfrbp_1 \logix.ram_r[1066]$_DFFE_PP_  (.CLK(net720),
    .RESET_B(net871),
    .D(_0080_),
    .Q_N(_5918_),
    .Q(\logix.ram_r[1066] ));
 sg13g2_dfrbp_1 \logix.ram_r[1067]$_DFFE_PP_  (.CLK(net711),
    .RESET_B(net872),
    .D(_0081_),
    .Q_N(_5917_),
    .Q(\logix.ram_r[1067] ));
 sg13g2_dfrbp_1 \logix.ram_r[1068]$_DFFE_PP_  (.CLK(net711),
    .RESET_B(net873),
    .D(_0082_),
    .Q_N(_5916_),
    .Q(\logix.ram_r[1068] ));
 sg13g2_dfrbp_1 \logix.ram_r[1069]$_DFFE_PP_  (.CLK(net711),
    .RESET_B(net874),
    .D(_0083_),
    .Q_N(_5915_),
    .Q(\logix.ram_r[1069] ));
 sg13g2_dfrbp_1 \logix.ram_r[106]$_DFFE_PP_  (.CLK(net715),
    .RESET_B(net875),
    .D(_0084_),
    .Q_N(_5914_),
    .Q(\logix.ram_r[106] ));
 sg13g2_dfrbp_1 \logix.ram_r[1070]$_DFFE_PP_  (.CLK(net706),
    .RESET_B(net876),
    .D(_0085_),
    .Q_N(_5913_),
    .Q(\logix.ram_r[1070] ));
 sg13g2_dfrbp_1 \logix.ram_r[1071]$_DFFE_PP_  (.CLK(net707),
    .RESET_B(net877),
    .D(_0086_),
    .Q_N(_5912_),
    .Q(\logix.ram_r[1071] ));
 sg13g2_dfrbp_1 \logix.ram_r[1072]$_DFFE_PP_  (.CLK(net712),
    .RESET_B(net878),
    .D(_0087_),
    .Q_N(_5911_),
    .Q(\logix.ram_r[1072] ));
 sg13g2_dfrbp_1 \logix.ram_r[1073]$_DFFE_PP_  (.CLK(net719),
    .RESET_B(net879),
    .D(_0088_),
    .Q_N(_5910_),
    .Q(\logix.ram_r[1073] ));
 sg13g2_dfrbp_1 \logix.ram_r[1074]$_DFFE_PP_  (.CLK(net720),
    .RESET_B(net880),
    .D(_0089_),
    .Q_N(_5909_),
    .Q(\logix.ram_r[1074] ));
 sg13g2_dfrbp_1 \logix.ram_r[1075]$_DFFE_PP_  (.CLK(net720),
    .RESET_B(net881),
    .D(_0090_),
    .Q_N(_5908_),
    .Q(\logix.ram_r[1075] ));
 sg13g2_dfrbp_1 \logix.ram_r[1076]$_DFFE_PP_  (.CLK(net711),
    .RESET_B(net882),
    .D(_0091_),
    .Q_N(_5907_),
    .Q(\logix.ram_r[1076] ));
 sg13g2_dfrbp_1 \logix.ram_r[1077]$_DFFE_PP_  (.CLK(net712),
    .RESET_B(net883),
    .D(_0092_),
    .Q_N(_5906_),
    .Q(\logix.ram_r[1077] ));
 sg13g2_dfrbp_1 \logix.ram_r[1078]$_DFFE_PP_  (.CLK(net707),
    .RESET_B(net884),
    .D(_0093_),
    .Q_N(_5905_),
    .Q(\logix.ram_r[1078] ));
 sg13g2_dfrbp_1 \logix.ram_r[1079]$_DFFE_PP_  (.CLK(net707),
    .RESET_B(net885),
    .D(_0094_),
    .Q_N(_5904_),
    .Q(\logix.ram_r[1079] ));
 sg13g2_dfrbp_1 \logix.ram_r[107]$_DFFE_PP_  (.CLK(net715),
    .RESET_B(net886),
    .D(_0095_),
    .Q_N(_5903_),
    .Q(\logix.ram_r[107] ));
 sg13g2_dfrbp_1 \logix.ram_r[1080]$_DFFE_PP_  (.CLK(net712),
    .RESET_B(net887),
    .D(_0096_),
    .Q_N(_5902_),
    .Q(\logix.ram_r[1080] ));
 sg13g2_dfrbp_1 \logix.ram_r[1081]$_DFFE_PP_  (.CLK(net719),
    .RESET_B(net888),
    .D(_0097_),
    .Q_N(_5901_),
    .Q(\logix.ram_r[1081] ));
 sg13g2_dfrbp_1 \logix.ram_r[1082]$_DFFE_PP_  (.CLK(net720),
    .RESET_B(net889),
    .D(_0098_),
    .Q_N(_5900_),
    .Q(\logix.ram_r[1082] ));
 sg13g2_dfrbp_1 \logix.ram_r[1083]$_DFFE_PP_  (.CLK(net712),
    .RESET_B(net890),
    .D(_0099_),
    .Q_N(_5899_),
    .Q(\logix.ram_r[1083] ));
 sg13g2_dfrbp_1 \logix.ram_r[1084]$_DFFE_PP_  (.CLK(net711),
    .RESET_B(net891),
    .D(_0100_),
    .Q_N(_5898_),
    .Q(\logix.ram_r[1084] ));
 sg13g2_dfrbp_1 \logix.ram_r[1085]$_DFFE_PP_  (.CLK(net711),
    .RESET_B(net892),
    .D(_0101_),
    .Q_N(_5897_),
    .Q(\logix.ram_r[1085] ));
 sg13g2_dfrbp_1 \logix.ram_r[1086]$_DFFE_PP_  (.CLK(net707),
    .RESET_B(net893),
    .D(_0102_),
    .Q_N(_5896_),
    .Q(\logix.ram_r[1086] ));
 sg13g2_dfrbp_1 \logix.ram_r[1087]$_DFFE_PP_  (.CLK(net707),
    .RESET_B(net894),
    .D(_0103_),
    .Q_N(_5895_),
    .Q(\logix.ram_r[1087] ));
 sg13g2_dfrbp_1 \logix.ram_r[1088]$_DFFE_PP_  (.CLK(net710),
    .RESET_B(net895),
    .D(_0104_),
    .Q_N(_5894_),
    .Q(\logix.ram_r[1088] ));
 sg13g2_dfrbp_1 \logix.ram_r[1089]$_DFFE_PP_  (.CLK(net710),
    .RESET_B(net896),
    .D(_0105_),
    .Q_N(_5893_),
    .Q(\logix.ram_r[1089] ));
 sg13g2_dfrbp_1 \logix.ram_r[108]$_DFFE_PP_  (.CLK(net715),
    .RESET_B(net897),
    .D(_0106_),
    .Q_N(_5892_),
    .Q(\logix.ram_r[108] ));
 sg13g2_dfrbp_1 \logix.ram_r[1090]$_DFFE_PP_  (.CLK(net711),
    .RESET_B(net898),
    .D(_0107_),
    .Q_N(_5891_),
    .Q(\logix.ram_r[1090] ));
 sg13g2_dfrbp_1 \logix.ram_r[1091]$_DFFE_PP_  (.CLK(net709),
    .RESET_B(net899),
    .D(_0108_),
    .Q_N(_5890_),
    .Q(\logix.ram_r[1091] ));
 sg13g2_dfrbp_1 \logix.ram_r[1092]$_DFFE_PP_  (.CLK(net708),
    .RESET_B(net900),
    .D(_0109_),
    .Q_N(_5889_),
    .Q(\logix.ram_r[1092] ));
 sg13g2_dfrbp_1 \logix.ram_r[1093]$_DFFE_PP_  (.CLK(net708),
    .RESET_B(net901),
    .D(_0110_),
    .Q_N(_5888_),
    .Q(\logix.ram_r[1093] ));
 sg13g2_dfrbp_1 \logix.ram_r[1094]$_DFFE_PP_  (.CLK(net704),
    .RESET_B(net902),
    .D(_0111_),
    .Q_N(_5887_),
    .Q(\logix.ram_r[1094] ));
 sg13g2_dfrbp_1 \logix.ram_r[1095]$_DFFE_PP_  (.CLK(net704),
    .RESET_B(net903),
    .D(_0112_),
    .Q_N(_5886_),
    .Q(\logix.ram_r[1095] ));
 sg13g2_dfrbp_1 \logix.ram_r[1096]$_DFFE_PP_  (.CLK(net708),
    .RESET_B(net904),
    .D(_0113_),
    .Q_N(_5885_),
    .Q(\logix.ram_r[1096] ));
 sg13g2_dfrbp_1 \logix.ram_r[1097]$_DFFE_PP_  (.CLK(net710),
    .RESET_B(net905),
    .D(_0114_),
    .Q_N(_5884_),
    .Q(\logix.ram_r[1097] ));
 sg13g2_dfrbp_1 \logix.ram_r[1098]$_DFFE_PP_  (.CLK(net709),
    .RESET_B(net906),
    .D(_0115_),
    .Q_N(_5883_),
    .Q(\logix.ram_r[1098] ));
 sg13g2_dfrbp_1 \logix.ram_r[1099]$_DFFE_PP_  (.CLK(net709),
    .RESET_B(net907),
    .D(_0116_),
    .Q_N(_5882_),
    .Q(\logix.ram_r[1099] ));
 sg13g2_dfrbp_1 \logix.ram_r[109]$_DFFE_PP_  (.CLK(net697),
    .RESET_B(net908),
    .D(_0117_),
    .Q_N(_5881_),
    .Q(\logix.ram_r[109] ));
 sg13g2_dfrbp_1 \logix.ram_r[10]$_DFFE_PP_  (.CLK(net658),
    .RESET_B(net909),
    .D(_0118_),
    .Q_N(_5880_),
    .Q(\logix.ram_r[10] ));
 sg13g2_dfrbp_1 \logix.ram_r[1100]$_DFFE_PP_  (.CLK(net708),
    .RESET_B(net910),
    .D(_0119_),
    .Q_N(_5879_),
    .Q(\logix.ram_r[1100] ));
 sg13g2_dfrbp_1 \logix.ram_r[1101]$_DFFE_PP_  (.CLK(net708),
    .RESET_B(net911),
    .D(_0120_),
    .Q_N(_5878_),
    .Q(\logix.ram_r[1101] ));
 sg13g2_dfrbp_1 \logix.ram_r[1102]$_DFFE_PP_  (.CLK(net704),
    .RESET_B(net912),
    .D(_0121_),
    .Q_N(_5877_),
    .Q(\logix.ram_r[1102] ));
 sg13g2_dfrbp_1 \logix.ram_r[1103]$_DFFE_PP_  (.CLK(net704),
    .RESET_B(net913),
    .D(_0122_),
    .Q_N(_5876_),
    .Q(\logix.ram_r[1103] ));
 sg13g2_dfrbp_1 \logix.ram_r[1104]$_DFFE_PP_  (.CLK(net705),
    .RESET_B(net914),
    .D(_0123_),
    .Q_N(_5875_),
    .Q(\logix.ram_r[1104] ));
 sg13g2_dfrbp_1 \logix.ram_r[1105]$_DFFE_PP_  (.CLK(net710),
    .RESET_B(net915),
    .D(_0124_),
    .Q_N(_5874_),
    .Q(\logix.ram_r[1105] ));
 sg13g2_dfrbp_1 \logix.ram_r[1106]$_DFFE_PP_  (.CLK(net708),
    .RESET_B(net916),
    .D(_0125_),
    .Q_N(_5873_),
    .Q(\logix.ram_r[1106] ));
 sg13g2_dfrbp_1 \logix.ram_r[1107]$_DFFE_PP_  (.CLK(net708),
    .RESET_B(net917),
    .D(_0126_),
    .Q_N(_5872_),
    .Q(\logix.ram_r[1107] ));
 sg13g2_dfrbp_1 \logix.ram_r[1108]$_DFFE_PP_  (.CLK(net709),
    .RESET_B(net918),
    .D(_0127_),
    .Q_N(_5871_),
    .Q(\logix.ram_r[1108] ));
 sg13g2_dfrbp_1 \logix.ram_r[1109]$_DFFE_PP_  (.CLK(net709),
    .RESET_B(net919),
    .D(_0128_),
    .Q_N(_5870_),
    .Q(\logix.ram_r[1109] ));
 sg13g2_dfrbp_1 \logix.ram_r[110]$_DFFE_PP_  (.CLK(net697),
    .RESET_B(net920),
    .D(_0129_),
    .Q_N(_5869_),
    .Q(\logix.ram_r[110] ));
 sg13g2_dfrbp_1 \logix.ram_r[1110]$_DFFE_PP_  (.CLK(net704),
    .RESET_B(net921),
    .D(_0130_),
    .Q_N(_5868_),
    .Q(\logix.ram_r[1110] ));
 sg13g2_dfrbp_1 \logix.ram_r[1111]$_DFFE_PP_  (.CLK(net708),
    .RESET_B(net922),
    .D(_0131_),
    .Q_N(_5867_),
    .Q(\logix.ram_r[1111] ));
 sg13g2_dfrbp_1 \logix.ram_r[1112]$_DFFE_PP_  (.CLK(net709),
    .RESET_B(net923),
    .D(_0132_),
    .Q_N(_5866_),
    .Q(\logix.ram_r[1112] ));
 sg13g2_dfrbp_1 \logix.ram_r[1113]$_DFFE_PP_  (.CLK(net711),
    .RESET_B(net924),
    .D(_0133_),
    .Q_N(_5865_),
    .Q(\logix.ram_r[1113] ));
 sg13g2_dfrbp_1 \logix.ram_r[1114]$_DFFE_PP_  (.CLK(net709),
    .RESET_B(net925),
    .D(_0134_),
    .Q_N(_5864_),
    .Q(\logix.ram_r[1114] ));
 sg13g2_dfrbp_1 \logix.ram_r[1115]$_DFFE_PP_  (.CLK(net713),
    .RESET_B(net926),
    .D(_0135_),
    .Q_N(_5863_),
    .Q(\logix.ram_r[1115] ));
 sg13g2_dfrbp_1 \logix.ram_r[1116]$_DFFE_PP_  (.CLK(net713),
    .RESET_B(net927),
    .D(_0136_),
    .Q_N(_5862_),
    .Q(\logix.ram_r[1116] ));
 sg13g2_dfrbp_1 \logix.ram_r[1117]$_DFFE_PP_  (.CLK(net704),
    .RESET_B(net928),
    .D(_0137_),
    .Q_N(_5861_),
    .Q(\logix.ram_r[1117] ));
 sg13g2_dfrbp_1 \logix.ram_r[1118]$_DFFE_PP_  (.CLK(net704),
    .RESET_B(net929),
    .D(_0138_),
    .Q_N(_5860_),
    .Q(\logix.ram_r[1118] ));
 sg13g2_dfrbp_1 \logix.ram_r[1119]$_DFFE_PP_  (.CLK(net704),
    .RESET_B(net930),
    .D(_0139_),
    .Q_N(_5859_),
    .Q(\logix.ram_r[1119] ));
 sg13g2_dfrbp_1 \logix.ram_r[111]$_DFFE_PP_  (.CLK(net716),
    .RESET_B(net931),
    .D(_0140_),
    .Q_N(_5858_),
    .Q(\logix.ram_r[111] ));
 sg13g2_dfrbp_1 \logix.ram_r[1120]$_DFFE_PP_  (.CLK(net703),
    .RESET_B(net932),
    .D(_0141_),
    .Q_N(_5857_),
    .Q(\logix.ram_r[1120] ));
 sg13g2_dfrbp_1 \logix.ram_r[1121]$_DFFE_PP_  (.CLK(net703),
    .RESET_B(net933),
    .D(_0142_),
    .Q_N(_5856_),
    .Q(\logix.ram_r[1121] ));
 sg13g2_dfrbp_1 \logix.ram_r[1122]$_DFFE_PP_  (.CLK(net703),
    .RESET_B(net934),
    .D(_0143_),
    .Q_N(_5855_),
    .Q(\logix.ram_r[1122] ));
 sg13g2_dfrbp_1 \logix.ram_r[1123]$_DFFE_PP_  (.CLK(net703),
    .RESET_B(net935),
    .D(_0144_),
    .Q_N(_5854_),
    .Q(\logix.ram_r[1123] ));
 sg13g2_dfrbp_1 \logix.ram_r[1124]$_DFFE_PP_  (.CLK(net703),
    .RESET_B(net936),
    .D(_0145_),
    .Q_N(_5853_),
    .Q(\logix.ram_r[1124] ));
 sg13g2_dfrbp_1 \logix.ram_r[1125]$_DFFE_PP_  (.CLK(net703),
    .RESET_B(net937),
    .D(_0146_),
    .Q_N(_5852_),
    .Q(\logix.ram_r[1125] ));
 sg13g2_dfrbp_1 \logix.ram_r[1126]$_DFFE_PP_  (.CLK(net686),
    .RESET_B(net938),
    .D(_0147_),
    .Q_N(_5851_),
    .Q(\logix.ram_r[1126] ));
 sg13g2_dfrbp_1 \logix.ram_r[1127]$_DFFE_PP_  (.CLK(net681),
    .RESET_B(net939),
    .D(_0148_),
    .Q_N(_5850_),
    .Q(\logix.ram_r[1127] ));
 sg13g2_dfrbp_1 \logix.ram_r[1128]$_DFFE_PP_  (.CLK(net686),
    .RESET_B(net940),
    .D(_0149_),
    .Q_N(_5849_),
    .Q(\logix.ram_r[1128] ));
 sg13g2_dfrbp_1 \logix.ram_r[1129]$_DFFE_PP_  (.CLK(net686),
    .RESET_B(net941),
    .D(_0150_),
    .Q_N(_5848_),
    .Q(\logix.ram_r[1129] ));
 sg13g2_dfrbp_1 \logix.ram_r[112]$_DFFE_PP_  (.CLK(net697),
    .RESET_B(net942),
    .D(_0151_),
    .Q_N(_5847_),
    .Q(\logix.ram_r[112] ));
 sg13g2_dfrbp_1 \logix.ram_r[1130]$_DFFE_PP_  (.CLK(net687),
    .RESET_B(net943),
    .D(_0152_),
    .Q_N(_5846_),
    .Q(\logix.ram_r[1130] ));
 sg13g2_dfrbp_1 \logix.ram_r[1131]$_DFFE_PP_  (.CLK(net687),
    .RESET_B(net944),
    .D(_0153_),
    .Q_N(_5845_),
    .Q(\logix.ram_r[1131] ));
 sg13g2_dfrbp_1 \logix.ram_r[1132]$_DFFE_PP_  (.CLK(net687),
    .RESET_B(net945),
    .D(_0154_),
    .Q_N(_5844_),
    .Q(\logix.ram_r[1132] ));
 sg13g2_dfrbp_1 \logix.ram_r[1133]$_DFFE_PP_  (.CLK(net687),
    .RESET_B(net946),
    .D(_0155_),
    .Q_N(_5843_),
    .Q(\logix.ram_r[1133] ));
 sg13g2_dfrbp_1 \logix.ram_r[1134]$_DFFE_PP_  (.CLK(net686),
    .RESET_B(net947),
    .D(_0156_),
    .Q_N(_5842_),
    .Q(\logix.ram_r[1134] ));
 sg13g2_dfrbp_1 \logix.ram_r[1135]$_DFFE_PP_  (.CLK(net681),
    .RESET_B(net948),
    .D(_0157_),
    .Q_N(_5841_),
    .Q(\logix.ram_r[1135] ));
 sg13g2_dfrbp_1 \logix.ram_r[1136]$_DFFE_PP_  (.CLK(net686),
    .RESET_B(net949),
    .D(_0158_),
    .Q_N(_5840_),
    .Q(\logix.ram_r[1136] ));
 sg13g2_dfrbp_1 \logix.ram_r[1137]$_DFFE_PP_  (.CLK(net686),
    .RESET_B(net950),
    .D(_0159_),
    .Q_N(_5839_),
    .Q(\logix.ram_r[1137] ));
 sg13g2_dfrbp_1 \logix.ram_r[1138]$_DFFE_PP_  (.CLK(net687),
    .RESET_B(net951),
    .D(_0160_),
    .Q_N(_5838_),
    .Q(\logix.ram_r[1138] ));
 sg13g2_dfrbp_1 \logix.ram_r[1139]$_DFFE_PP_  (.CLK(net687),
    .RESET_B(net952),
    .D(_0161_),
    .Q_N(_5837_),
    .Q(\logix.ram_r[1139] ));
 sg13g2_dfrbp_1 \logix.ram_r[113]$_DFFE_PP_  (.CLK(net697),
    .RESET_B(net953),
    .D(_0162_),
    .Q_N(_5836_),
    .Q(\logix.ram_r[113] ));
 sg13g2_dfrbp_1 \logix.ram_r[1140]$_DFFE_PP_  (.CLK(net705),
    .RESET_B(net954),
    .D(_0163_),
    .Q_N(_5835_),
    .Q(\logix.ram_r[1140] ));
 sg13g2_dfrbp_1 \logix.ram_r[1141]$_DFFE_PP_  (.CLK(net688),
    .RESET_B(net955),
    .D(_0164_),
    .Q_N(_5834_),
    .Q(\logix.ram_r[1141] ));
 sg13g2_dfrbp_1 \logix.ram_r[1142]$_DFFE_PP_  (.CLK(net688),
    .RESET_B(net956),
    .D(_0165_),
    .Q_N(_5833_),
    .Q(\logix.ram_r[1142] ));
 sg13g2_dfrbp_1 \logix.ram_r[1143]$_DFFE_PP_  (.CLK(net686),
    .RESET_B(net957),
    .D(_0166_),
    .Q_N(_5832_),
    .Q(\logix.ram_r[1143] ));
 sg13g2_dfrbp_1 \logix.ram_r[1144]$_DFFE_PP_  (.CLK(net686),
    .RESET_B(net958),
    .D(_0167_),
    .Q_N(_5831_),
    .Q(\logix.ram_r[1144] ));
 sg13g2_dfrbp_1 \logix.ram_r[1145]$_DFFE_PP_  (.CLK(net687),
    .RESET_B(net959),
    .D(_0168_),
    .Q_N(_5830_),
    .Q(\logix.ram_r[1145] ));
 sg13g2_dfrbp_1 \logix.ram_r[1146]$_DFFE_PP_  (.CLK(net687),
    .RESET_B(net960),
    .D(_0169_),
    .Q_N(_5829_),
    .Q(\logix.ram_r[1146] ));
 sg13g2_dfrbp_1 \logix.ram_r[1147]$_DFFE_PP_  (.CLK(net703),
    .RESET_B(net961),
    .D(_0170_),
    .Q_N(_5828_),
    .Q(\logix.ram_r[1147] ));
 sg13g2_dfrbp_1 \logix.ram_r[1148]$_DFFE_PP_  (.CLK(net703),
    .RESET_B(net962),
    .D(_0171_),
    .Q_N(_5827_),
    .Q(\logix.ram_r[1148] ));
 sg13g2_dfrbp_1 \logix.ram_r[1149]$_DFFE_PP_  (.CLK(net705),
    .RESET_B(net963),
    .D(_0172_),
    .Q_N(_5826_),
    .Q(\logix.ram_r[1149] ));
 sg13g2_dfrbp_1 \logix.ram_r[114]$_DFFE_PP_  (.CLK(net698),
    .RESET_B(net964),
    .D(_0173_),
    .Q_N(_5825_),
    .Q(\logix.ram_r[114] ));
 sg13g2_dfrbp_1 \logix.ram_r[1150]$_DFFE_PP_  (.CLK(net688),
    .RESET_B(net965),
    .D(_0174_),
    .Q_N(_5824_),
    .Q(\logix.ram_r[1150] ));
 sg13g2_dfrbp_1 \logix.ram_r[1151]$_DFFE_PP_  (.CLK(net688),
    .RESET_B(net966),
    .D(_0175_),
    .Q_N(_5823_),
    .Q(\logix.ram_r[1151] ));
 sg13g2_dfrbp_1 \logix.ram_r[1152]$_DFFE_PP_  (.CLK(net688),
    .RESET_B(net967),
    .D(_0176_),
    .Q_N(_5822_),
    .Q(\logix.ram_r[1152] ));
 sg13g2_dfrbp_1 \logix.ram_r[1153]$_DFFE_PP_  (.CLK(net752),
    .RESET_B(net968),
    .D(_0177_),
    .Q_N(_5821_),
    .Q(\logix.ram_r[1153] ));
 sg13g2_dfrbp_1 \logix.ram_r[1154]$_DFFE_PP_  (.CLK(net752),
    .RESET_B(net969),
    .D(_0178_),
    .Q_N(_5820_),
    .Q(\logix.ram_r[1154] ));
 sg13g2_dfrbp_1 \logix.ram_r[1155]$_DFFE_PP_  (.CLK(net752),
    .RESET_B(net970),
    .D(_0179_),
    .Q_N(_5819_),
    .Q(\logix.ram_r[1155] ));
 sg13g2_dfrbp_1 \logix.ram_r[1156]$_DFFE_PP_  (.CLK(net752),
    .RESET_B(net971),
    .D(_0180_),
    .Q_N(_5818_),
    .Q(\logix.ram_r[1156] ));
 sg13g2_dfrbp_1 \logix.ram_r[1157]$_DFFE_PP_  (.CLK(net752),
    .RESET_B(net972),
    .D(_0181_),
    .Q_N(_5817_),
    .Q(\logix.ram_r[1157] ));
 sg13g2_dfrbp_1 \logix.ram_r[1158]$_DFFE_PP_  (.CLK(net755),
    .RESET_B(net973),
    .D(_0182_),
    .Q_N(_5816_),
    .Q(\logix.ram_r[1158] ));
 sg13g2_dfrbp_1 \logix.ram_r[1159]$_DFFE_PP_  (.CLK(net755),
    .RESET_B(net974),
    .D(_0183_),
    .Q_N(_5815_),
    .Q(\logix.ram_r[1159] ));
 sg13g2_dfrbp_1 \logix.ram_r[115]$_DFFE_PP_  (.CLK(net716),
    .RESET_B(net975),
    .D(_0184_),
    .Q_N(_5814_),
    .Q(\logix.ram_r[115] ));
 sg13g2_dfrbp_1 \logix.ram_r[1160]$_DFFE_PP_  (.CLK(net752),
    .RESET_B(net976),
    .D(_0185_),
    .Q_N(_5813_),
    .Q(\logix.ram_r[1160] ));
 sg13g2_dfrbp_1 \logix.ram_r[1161]$_DFFE_PP_  (.CLK(net753),
    .RESET_B(net977),
    .D(_0186_),
    .Q_N(_5812_),
    .Q(\logix.ram_r[1161] ));
 sg13g2_dfrbp_1 \logix.ram_r[1162]$_DFFE_PP_  (.CLK(net753),
    .RESET_B(net978),
    .D(_0187_),
    .Q_N(_5811_),
    .Q(\logix.ram_r[1162] ));
 sg13g2_dfrbp_1 \logix.ram_r[1163]$_DFFE_PP_  (.CLK(net753),
    .RESET_B(net979),
    .D(_0188_),
    .Q_N(_5810_),
    .Q(\logix.ram_r[1163] ));
 sg13g2_dfrbp_1 \logix.ram_r[1164]$_DFFE_PP_  (.CLK(net754),
    .RESET_B(net980),
    .D(_0189_),
    .Q_N(_5809_),
    .Q(\logix.ram_r[1164] ));
 sg13g2_dfrbp_1 \logix.ram_r[1165]$_DFFE_PP_  (.CLK(net756),
    .RESET_B(net981),
    .D(_0190_),
    .Q_N(_5808_),
    .Q(\logix.ram_r[1165] ));
 sg13g2_dfrbp_1 \logix.ram_r[1166]$_DFFE_PP_  (.CLK(net758),
    .RESET_B(net982),
    .D(_0191_),
    .Q_N(_5807_),
    .Q(\logix.ram_r[1166] ));
 sg13g2_dfrbp_1 \logix.ram_r[1167]$_DFFE_PP_  (.CLK(net755),
    .RESET_B(net983),
    .D(_0192_),
    .Q_N(_5806_),
    .Q(\logix.ram_r[1167] ));
 sg13g2_dfrbp_1 \logix.ram_r[1168]$_DFFE_PP_  (.CLK(net752),
    .RESET_B(net984),
    .D(_0193_),
    .Q_N(_5805_),
    .Q(\logix.ram_r[1168] ));
 sg13g2_dfrbp_1 \logix.ram_r[1169]$_DFFE_PP_  (.CLK(net753),
    .RESET_B(net985),
    .D(_0194_),
    .Q_N(_5804_),
    .Q(\logix.ram_r[1169] ));
 sg13g2_dfrbp_1 \logix.ram_r[116]$_DFFE_PP_  (.CLK(net699),
    .RESET_B(net986),
    .D(_0195_),
    .Q_N(_5803_),
    .Q(\logix.ram_r[116] ));
 sg13g2_dfrbp_1 \logix.ram_r[1170]$_DFFE_PP_  (.CLK(net753),
    .RESET_B(net987),
    .D(_0196_),
    .Q_N(_5802_),
    .Q(\logix.ram_r[1170] ));
 sg13g2_dfrbp_1 \logix.ram_r[1171]$_DFFE_PP_  (.CLK(net754),
    .RESET_B(net988),
    .D(_0197_),
    .Q_N(_5801_),
    .Q(\logix.ram_r[1171] ));
 sg13g2_dfrbp_1 \logix.ram_r[1172]$_DFFE_PP_  (.CLK(net754),
    .RESET_B(net989),
    .D(_0198_),
    .Q_N(_5800_),
    .Q(\logix.ram_r[1172] ));
 sg13g2_dfrbp_1 \logix.ram_r[1173]$_DFFE_PP_  (.CLK(net756),
    .RESET_B(net990),
    .D(_0199_),
    .Q_N(_5799_),
    .Q(\logix.ram_r[1173] ));
 sg13g2_dfrbp_1 \logix.ram_r[1174]$_DFFE_PP_  (.CLK(net756),
    .RESET_B(net991),
    .D(_0200_),
    .Q_N(_5798_),
    .Q(\logix.ram_r[1174] ));
 sg13g2_dfrbp_1 \logix.ram_r[1175]$_DFFE_PP_  (.CLK(net758),
    .RESET_B(net992),
    .D(_0201_),
    .Q_N(_5797_),
    .Q(\logix.ram_r[1175] ));
 sg13g2_dfrbp_1 \logix.ram_r[1176]$_DFFE_PP_  (.CLK(net752),
    .RESET_B(net993),
    .D(_0202_),
    .Q_N(_5796_),
    .Q(\logix.ram_r[1176] ));
 sg13g2_dfrbp_1 \logix.ram_r[1177]$_DFFE_PP_  (.CLK(net753),
    .RESET_B(net994),
    .D(_0203_),
    .Q_N(_5795_),
    .Q(\logix.ram_r[1177] ));
 sg13g2_dfrbp_1 \logix.ram_r[1178]$_DFFE_PP_  (.CLK(net753),
    .RESET_B(net995),
    .D(_0204_),
    .Q_N(_5794_),
    .Q(\logix.ram_r[1178] ));
 sg13g2_dfrbp_1 \logix.ram_r[1179]$_DFFE_PP_  (.CLK(net753),
    .RESET_B(net996),
    .D(_0205_),
    .Q_N(_5793_),
    .Q(\logix.ram_r[1179] ));
 sg13g2_dfrbp_1 \logix.ram_r[117]$_DFFE_PP_  (.CLK(net695),
    .RESET_B(net997),
    .D(_0206_),
    .Q_N(_5792_),
    .Q(\logix.ram_r[117] ));
 sg13g2_dfrbp_1 \logix.ram_r[1180]$_DFFE_PP_  (.CLK(net754),
    .RESET_B(net998),
    .D(_0207_),
    .Q_N(_5791_),
    .Q(\logix.ram_r[1180] ));
 sg13g2_dfrbp_1 \logix.ram_r[1181]$_DFFE_PP_  (.CLK(net756),
    .RESET_B(net999),
    .D(_0208_),
    .Q_N(_5790_),
    .Q(\logix.ram_r[1181] ));
 sg13g2_dfrbp_1 \logix.ram_r[1182]$_DFFE_PP_  (.CLK(net756),
    .RESET_B(net1000),
    .D(_0209_),
    .Q_N(_5789_),
    .Q(\logix.ram_r[1182] ));
 sg13g2_dfrbp_1 \logix.ram_r[1183]$_DFFE_PP_  (.CLK(net758),
    .RESET_B(net1001),
    .D(_0210_),
    .Q_N(_5788_),
    .Q(\logix.ram_r[1183] ));
 sg13g2_dfrbp_1 \logix.ram_r[1184]$_DFFE_PP_  (.CLK(net748),
    .RESET_B(net1002),
    .D(_0211_),
    .Q_N(_5787_),
    .Q(\logix.ram_r[1184] ));
 sg13g2_dfrbp_1 \logix.ram_r[1185]$_DFFE_PP_  (.CLK(net748),
    .RESET_B(net1003),
    .D(_0212_),
    .Q_N(_5786_),
    .Q(\logix.ram_r[1185] ));
 sg13g2_dfrbp_1 \logix.ram_r[1186]$_DFFE_PP_  (.CLK(net749),
    .RESET_B(net1004),
    .D(_0213_),
    .Q_N(_5785_),
    .Q(\logix.ram_r[1186] ));
 sg13g2_dfrbp_1 \logix.ram_r[1187]$_DFFE_PP_  (.CLK(net749),
    .RESET_B(net1005),
    .D(_0214_),
    .Q_N(_5784_),
    .Q(\logix.ram_r[1187] ));
 sg13g2_dfrbp_1 \logix.ram_r[1188]$_DFFE_PP_  (.CLK(net749),
    .RESET_B(net1006),
    .D(_0215_),
    .Q_N(_5783_),
    .Q(\logix.ram_r[1188] ));
 sg13g2_dfrbp_1 \logix.ram_r[1189]$_DFFE_PP_  (.CLK(net750),
    .RESET_B(net1007),
    .D(_0216_),
    .Q_N(_5782_),
    .Q(\logix.ram_r[1189] ));
 sg13g2_dfrbp_1 \logix.ram_r[118]$_DFFE_PP_  (.CLK(net699),
    .RESET_B(net1008),
    .D(_0217_),
    .Q_N(_5781_),
    .Q(\logix.ram_r[118] ));
 sg13g2_dfrbp_1 \logix.ram_r[1190]$_DFFE_PP_  (.CLK(net733),
    .RESET_B(net1009),
    .D(_0218_),
    .Q_N(_5780_),
    .Q(\logix.ram_r[1190] ));
 sg13g2_dfrbp_1 \logix.ram_r[1191]$_DFFE_PP_  (.CLK(net734),
    .RESET_B(net1010),
    .D(_0219_),
    .Q_N(_5779_),
    .Q(\logix.ram_r[1191] ));
 sg13g2_dfrbp_1 \logix.ram_r[1192]$_DFFE_PP_  (.CLK(net732),
    .RESET_B(net1011),
    .D(_0220_),
    .Q_N(_5778_),
    .Q(\logix.ram_r[1192] ));
 sg13g2_dfrbp_1 \logix.ram_r[1193]$_DFFE_PP_  (.CLK(net732),
    .RESET_B(net1012),
    .D(_0221_),
    .Q_N(_5777_),
    .Q(\logix.ram_r[1193] ));
 sg13g2_dfrbp_1 \logix.ram_r[1194]$_DFFE_PP_  (.CLK(net748),
    .RESET_B(net1013),
    .D(_0222_),
    .Q_N(_5776_),
    .Q(\logix.ram_r[1194] ));
 sg13g2_dfrbp_1 \logix.ram_r[1195]$_DFFE_PP_  (.CLK(net748),
    .RESET_B(net1014),
    .D(_0223_),
    .Q_N(_5775_),
    .Q(\logix.ram_r[1195] ));
 sg13g2_dfrbp_1 \logix.ram_r[1196]$_DFFE_PP_  (.CLK(net748),
    .RESET_B(net1015),
    .D(_0224_),
    .Q_N(_5774_),
    .Q(\logix.ram_r[1196] ));
 sg13g2_dfrbp_1 \logix.ram_r[1197]$_DFFE_PP_  (.CLK(net751),
    .RESET_B(net1016),
    .D(_0225_),
    .Q_N(_5773_),
    .Q(\logix.ram_r[1197] ));
 sg13g2_dfrbp_1 \logix.ram_r[1198]$_DFFE_PP_  (.CLK(net733),
    .RESET_B(net1017),
    .D(_0226_),
    .Q_N(_5772_),
    .Q(\logix.ram_r[1198] ));
 sg13g2_dfrbp_1 \logix.ram_r[1199]$_DFFE_PP_  (.CLK(net733),
    .RESET_B(net1018),
    .D(_0227_),
    .Q_N(_5771_),
    .Q(\logix.ram_r[1199] ));
 sg13g2_dfrbp_1 \logix.ram_r[119]$_DFFE_PP_  (.CLK(net699),
    .RESET_B(net1019),
    .D(_0228_),
    .Q_N(_5770_),
    .Q(\logix.ram_r[119] ));
 sg13g2_dfrbp_1 \logix.ram_r[11]$_DFFE_PP_  (.CLK(net658),
    .RESET_B(net1020),
    .D(_0229_),
    .Q_N(_5769_),
    .Q(\logix.ram_r[11] ));
 sg13g2_dfrbp_1 \logix.ram_r[1200]$_DFFE_PP_  (.CLK(net732),
    .RESET_B(net1021),
    .D(_0230_),
    .Q_N(_5768_),
    .Q(\logix.ram_r[1200] ));
 sg13g2_dfrbp_1 \logix.ram_r[1201]$_DFFE_PP_  (.CLK(net732),
    .RESET_B(net1022),
    .D(_0231_),
    .Q_N(_5767_),
    .Q(\logix.ram_r[1201] ));
 sg13g2_dfrbp_1 \logix.ram_r[1202]$_DFFE_PP_  (.CLK(net748),
    .RESET_B(net1023),
    .D(_0232_),
    .Q_N(_5766_),
    .Q(\logix.ram_r[1202] ));
 sg13g2_dfrbp_1 \logix.ram_r[1203]$_DFFE_PP_  (.CLK(net748),
    .RESET_B(net1024),
    .D(_0233_),
    .Q_N(_5765_),
    .Q(\logix.ram_r[1203] ));
 sg13g2_dfrbp_1 \logix.ram_r[1204]$_DFFE_PP_  (.CLK(net748),
    .RESET_B(net1025),
    .D(_0234_),
    .Q_N(_5764_),
    .Q(\logix.ram_r[1204] ));
 sg13g2_dfrbp_1 \logix.ram_r[1205]$_DFFE_PP_  (.CLK(net751),
    .RESET_B(net1026),
    .D(_0235_),
    .Q_N(_5763_),
    .Q(\logix.ram_r[1205] ));
 sg13g2_dfrbp_1 \logix.ram_r[1206]$_DFFE_PP_  (.CLK(net733),
    .RESET_B(net1027),
    .D(_0236_),
    .Q_N(_5762_),
    .Q(\logix.ram_r[1206] ));
 sg13g2_dfrbp_1 \logix.ram_r[1207]$_DFFE_PP_  (.CLK(net733),
    .RESET_B(net1028),
    .D(_0237_),
    .Q_N(_5761_),
    .Q(\logix.ram_r[1207] ));
 sg13g2_dfrbp_1 \logix.ram_r[1208]$_DFFE_PP_  (.CLK(net732),
    .RESET_B(net1029),
    .D(_0238_),
    .Q_N(_5760_),
    .Q(\logix.ram_r[1208] ));
 sg13g2_dfrbp_1 \logix.ram_r[1209]$_DFFE_PP_  (.CLK(net735),
    .RESET_B(net1030),
    .D(_0239_),
    .Q_N(_5759_),
    .Q(\logix.ram_r[1209] ));
 sg13g2_dfrbp_1 \logix.ram_r[120]$_DFFE_PP_  (.CLK(net699),
    .RESET_B(net1031),
    .D(_0240_),
    .Q_N(_5758_),
    .Q(\logix.ram_r[120] ));
 sg13g2_dfrbp_1 \logix.ram_r[1210]$_DFFE_PP_  (.CLK(net749),
    .RESET_B(net1032),
    .D(_0241_),
    .Q_N(_5757_),
    .Q(\logix.ram_r[1210] ));
 sg13g2_dfrbp_1 \logix.ram_r[1211]$_DFFE_PP_  (.CLK(net749),
    .RESET_B(net1033),
    .D(_0242_),
    .Q_N(_5756_),
    .Q(\logix.ram_r[1211] ));
 sg13g2_dfrbp_1 \logix.ram_r[1212]$_DFFE_PP_  (.CLK(net749),
    .RESET_B(net1034),
    .D(_0243_),
    .Q_N(_5755_),
    .Q(\logix.ram_r[1212] ));
 sg13g2_dfrbp_1 \logix.ram_r[1213]$_DFFE_PP_  (.CLK(net750),
    .RESET_B(net1035),
    .D(_0244_),
    .Q_N(_5754_),
    .Q(\logix.ram_r[1213] ));
 sg13g2_dfrbp_1 \logix.ram_r[1214]$_DFFE_PP_  (.CLK(net750),
    .RESET_B(net1036),
    .D(_0245_),
    .Q_N(_5753_),
    .Q(\logix.ram_r[1214] ));
 sg13g2_dfrbp_1 \logix.ram_r[1215]$_DFFE_PP_  (.CLK(net750),
    .RESET_B(net1037),
    .D(_0246_),
    .Q_N(_5752_),
    .Q(\logix.ram_r[1215] ));
 sg13g2_dfrbp_1 \logix.ram_r[1216]$_DFFE_PP_  (.CLK(net724),
    .RESET_B(net1038),
    .D(_0247_),
    .Q_N(_5751_),
    .Q(\logix.ram_r[1216] ));
 sg13g2_dfrbp_1 \logix.ram_r[1217]$_DFFE_PP_  (.CLK(net719),
    .RESET_B(net1039),
    .D(_0248_),
    .Q_N(_5750_),
    .Q(\logix.ram_r[1217] ));
 sg13g2_dfrbp_1 \logix.ram_r[1218]$_DFFE_PP_  (.CLK(net719),
    .RESET_B(net1040),
    .D(_0249_),
    .Q_N(_5749_),
    .Q(\logix.ram_r[1218] ));
 sg13g2_dfrbp_1 \logix.ram_r[1219]$_DFFE_PP_  (.CLK(net719),
    .RESET_B(net1041),
    .D(_0250_),
    .Q_N(_5748_),
    .Q(\logix.ram_r[1219] ));
 sg13g2_dfrbp_1 \logix.ram_r[121]$_DFFE_PP_  (.CLK(net698),
    .RESET_B(net1042),
    .D(_0251_),
    .Q_N(_5747_),
    .Q(\logix.ram_r[121] ));
 sg13g2_dfrbp_1 \logix.ram_r[1220]$_DFFE_PP_  (.CLK(net720),
    .RESET_B(net1043),
    .D(_0252_),
    .Q_N(_5746_),
    .Q(\logix.ram_r[1220] ));
 sg13g2_dfrbp_1 \logix.ram_r[1221]$_DFFE_PP_  (.CLK(net724),
    .RESET_B(net1044),
    .D(_0253_),
    .Q_N(_5745_),
    .Q(\logix.ram_r[1221] ));
 sg13g2_dfrbp_1 \logix.ram_r[1222]$_DFFE_PP_  (.CLK(net724),
    .RESET_B(net1045),
    .D(_0254_),
    .Q_N(_5744_),
    .Q(\logix.ram_r[1222] ));
 sg13g2_dfrbp_1 \logix.ram_r[1223]$_DFFE_PP_  (.CLK(net724),
    .RESET_B(net1046),
    .D(_0255_),
    .Q_N(_5743_),
    .Q(\logix.ram_r[1223] ));
 sg13g2_dfrbp_1 \logix.ram_r[1224]$_DFFE_PP_  (.CLK(net724),
    .RESET_B(net1047),
    .D(_0256_),
    .Q_N(_5742_),
    .Q(\logix.ram_r[1224] ));
 sg13g2_dfrbp_1 \logix.ram_r[1225]$_DFFE_PP_  (.CLK(net722),
    .RESET_B(net1048),
    .D(_0257_),
    .Q_N(_5741_),
    .Q(\logix.ram_r[1225] ));
 sg13g2_dfrbp_1 \logix.ram_r[1226]$_DFFE_PP_  (.CLK(net719),
    .RESET_B(net1049),
    .D(_0258_),
    .Q_N(_5740_),
    .Q(\logix.ram_r[1226] ));
 sg13g2_dfrbp_1 \logix.ram_r[1227]$_DFFE_PP_  (.CLK(net719),
    .RESET_B(net1050),
    .D(_0259_),
    .Q_N(_5739_),
    .Q(\logix.ram_r[1227] ));
 sg13g2_dfrbp_1 \logix.ram_r[1228]$_DFFE_PP_  (.CLK(net721),
    .RESET_B(net1051),
    .D(_0260_),
    .Q_N(_5738_),
    .Q(\logix.ram_r[1228] ));
 sg13g2_dfrbp_1 \logix.ram_r[1229]$_DFFE_PP_  (.CLK(net723),
    .RESET_B(net1052),
    .D(_0261_),
    .Q_N(_5737_),
    .Q(\logix.ram_r[1229] ));
 sg13g2_dfrbp_1 \logix.ram_r[122]$_DFFE_PP_  (.CLK(net698),
    .RESET_B(net1053),
    .D(_0262_),
    .Q_N(_5736_),
    .Q(\logix.ram_r[122] ));
 sg13g2_dfrbp_1 \logix.ram_r[1230]$_DFFE_PP_  (.CLK(net723),
    .RESET_B(net1054),
    .D(_0263_),
    .Q_N(_5735_),
    .Q(\logix.ram_r[1230] ));
 sg13g2_dfrbp_1 \logix.ram_r[1231]$_DFFE_PP_  (.CLK(net723),
    .RESET_B(net1055),
    .D(_0264_),
    .Q_N(_5734_),
    .Q(\logix.ram_r[1231] ));
 sg13g2_dfrbp_1 \logix.ram_r[1232]$_DFFE_PP_  (.CLK(net724),
    .RESET_B(net1056),
    .D(_0265_),
    .Q_N(_5733_),
    .Q(\logix.ram_r[1232] ));
 sg13g2_dfrbp_1 \logix.ram_r[1233]$_DFFE_PP_  (.CLK(net722),
    .RESET_B(net1057),
    .D(_0266_),
    .Q_N(_5732_),
    .Q(\logix.ram_r[1233] ));
 sg13g2_dfrbp_1 \logix.ram_r[1234]$_DFFE_PP_  (.CLK(net722),
    .RESET_B(net1058),
    .D(_0267_),
    .Q_N(_5731_),
    .Q(\logix.ram_r[1234] ));
 sg13g2_dfrbp_1 \logix.ram_r[1235]$_DFFE_PP_  (.CLK(net720),
    .RESET_B(net1059),
    .D(_0268_),
    .Q_N(_5730_),
    .Q(\logix.ram_r[1235] ));
 sg13g2_dfrbp_1 \logix.ram_r[1236]$_DFFE_PP_  (.CLK(net721),
    .RESET_B(net1060),
    .D(_0269_),
    .Q_N(_5729_),
    .Q(\logix.ram_r[1236] ));
 sg13g2_dfrbp_1 \logix.ram_r[1237]$_DFFE_PP_  (.CLK(net723),
    .RESET_B(net1061),
    .D(_0270_),
    .Q_N(_5728_),
    .Q(\logix.ram_r[1237] ));
 sg13g2_dfrbp_1 \logix.ram_r[1238]$_DFFE_PP_  (.CLK(net723),
    .RESET_B(net1062),
    .D(_0271_),
    .Q_N(_5727_),
    .Q(\logix.ram_r[1238] ));
 sg13g2_dfrbp_1 \logix.ram_r[1239]$_DFFE_PP_  (.CLK(net725),
    .RESET_B(net1063),
    .D(_0272_),
    .Q_N(_5726_),
    .Q(\logix.ram_r[1239] ));
 sg13g2_dfrbp_1 \logix.ram_r[123]$_DFFE_PP_  (.CLK(net698),
    .RESET_B(net1064),
    .D(_0273_),
    .Q_N(_5725_),
    .Q(\logix.ram_r[123] ));
 sg13g2_dfrbp_1 \logix.ram_r[1240]$_DFFE_PP_  (.CLK(net724),
    .RESET_B(net1065),
    .D(_0274_),
    .Q_N(_5724_),
    .Q(\logix.ram_r[1240] ));
 sg13g2_dfrbp_1 \logix.ram_r[1241]$_DFFE_PP_  (.CLK(net721),
    .RESET_B(net1066),
    .D(_0275_),
    .Q_N(_5723_),
    .Q(\logix.ram_r[1241] ));
 sg13g2_dfrbp_1 \logix.ram_r[1242]$_DFFE_PP_  (.CLK(net720),
    .RESET_B(net1067),
    .D(_0276_),
    .Q_N(_5722_),
    .Q(\logix.ram_r[1242] ));
 sg13g2_dfrbp_1 \logix.ram_r[1243]$_DFFE_PP_  (.CLK(net720),
    .RESET_B(net1068),
    .D(_0277_),
    .Q_N(_5721_),
    .Q(\logix.ram_r[1243] ));
 sg13g2_dfrbp_1 \logix.ram_r[1244]$_DFFE_PP_  (.CLK(net721),
    .RESET_B(net1069),
    .D(_0278_),
    .Q_N(_5720_),
    .Q(\logix.ram_r[1244] ));
 sg13g2_dfrbp_1 \logix.ram_r[1245]$_DFFE_PP_  (.CLK(net721),
    .RESET_B(net1070),
    .D(_0279_),
    .Q_N(_5719_),
    .Q(\logix.ram_r[1245] ));
 sg13g2_dfrbp_1 \logix.ram_r[1246]$_DFFE_PP_  (.CLK(net723),
    .RESET_B(net1071),
    .D(_0280_),
    .Q_N(_5718_),
    .Q(\logix.ram_r[1246] ));
 sg13g2_dfrbp_1 \logix.ram_r[1247]$_DFFE_PP_  (.CLK(net723),
    .RESET_B(net1072),
    .D(_0281_),
    .Q_N(_5717_),
    .Q(\logix.ram_r[1247] ));
 sg13g2_dfrbp_1 \logix.ram_r[1248]$_DFFE_PP_  (.CLK(net723),
    .RESET_B(net1073),
    .D(_0282_),
    .Q_N(_5716_),
    .Q(\logix.ram_r[1248] ));
 sg13g2_dfrbp_1 \logix.ram_r[1249]$_DFFE_PP_  (.CLK(net716),
    .RESET_B(net1074),
    .D(_0283_),
    .Q_N(_5715_),
    .Q(\logix.ram_r[1249] ));
 sg13g2_dfrbp_1 \logix.ram_r[124]$_DFFE_PP_  (.CLK(net698),
    .RESET_B(net1075),
    .D(_0284_),
    .Q_N(_5714_),
    .Q(\logix.ram_r[124] ));
 sg13g2_dfrbp_1 \logix.ram_r[1250]$_DFFE_PP_  (.CLK(net716),
    .RESET_B(net1076),
    .D(_0285_),
    .Q_N(_5713_),
    .Q(\logix.ram_r[1250] ));
 sg13g2_dfrbp_1 \logix.ram_r[1251]$_DFFE_PP_  (.CLK(net715),
    .RESET_B(net1077),
    .D(_0286_),
    .Q_N(_5712_),
    .Q(\logix.ram_r[1251] ));
 sg13g2_dfrbp_1 \logix.ram_r[1252]$_DFFE_PP_  (.CLK(net718),
    .RESET_B(net1078),
    .D(_0287_),
    .Q_N(_5711_),
    .Q(\logix.ram_r[1252] ));
 sg13g2_dfrbp_1 \logix.ram_r[1253]$_DFFE_PP_  (.CLK(net718),
    .RESET_B(net1079),
    .D(_0288_),
    .Q_N(_5710_),
    .Q(\logix.ram_r[1253] ));
 sg13g2_dfrbp_1 \logix.ram_r[1254]$_DFFE_PP_  (.CLK(net718),
    .RESET_B(net1080),
    .D(_0289_),
    .Q_N(_5709_),
    .Q(\logix.ram_r[1254] ));
 sg13g2_dfrbp_1 \logix.ram_r[1255]$_DFFE_PP_  (.CLK(net699),
    .RESET_B(net1081),
    .D(_0290_),
    .Q_N(_5708_),
    .Q(\logix.ram_r[1255] ));
 sg13g2_dfrbp_1 \logix.ram_r[1256]$_DFFE_PP_  (.CLK(net700),
    .RESET_B(net1082),
    .D(_0291_),
    .Q_N(_5707_),
    .Q(\logix.ram_r[1256] ));
 sg13g2_dfrbp_1 \logix.ram_r[1257]$_DFFE_PP_  (.CLK(net700),
    .RESET_B(net1083),
    .D(_0292_),
    .Q_N(_5706_),
    .Q(\logix.ram_r[1257] ));
 sg13g2_dfrbp_1 \logix.ram_r[1258]$_DFFE_PP_  (.CLK(net716),
    .RESET_B(net1084),
    .D(_0293_),
    .Q_N(_5705_),
    .Q(\logix.ram_r[1258] ));
 sg13g2_dfrbp_1 \logix.ram_r[1259]$_DFFE_PP_  (.CLK(net717),
    .RESET_B(net1085),
    .D(_0294_),
    .Q_N(_5704_),
    .Q(\logix.ram_r[1259] ));
 sg13g2_dfrbp_1 \logix.ram_r[125]$_DFFE_PP_  (.CLK(net699),
    .RESET_B(net1086),
    .D(_0295_),
    .Q_N(_5703_),
    .Q(\logix.ram_r[125] ));
 sg13g2_dfrbp_1 \logix.ram_r[1260]$_DFFE_PP_  (.CLK(net717),
    .RESET_B(net1087),
    .D(_0296_),
    .Q_N(_5702_),
    .Q(\logix.ram_r[1260] ));
 sg13g2_dfrbp_1 \logix.ram_r[1261]$_DFFE_PP_  (.CLK(net717),
    .RESET_B(net1088),
    .D(_0297_),
    .Q_N(_5701_),
    .Q(\logix.ram_r[1261] ));
 sg13g2_dfrbp_1 \logix.ram_r[1262]$_DFFE_PP_  (.CLK(net717),
    .RESET_B(net1089),
    .D(_0298_),
    .Q_N(_5700_),
    .Q(\logix.ram_r[1262] ));
 sg13g2_dfrbp_1 \logix.ram_r[1263]$_DFFE_PP_  (.CLK(net700),
    .RESET_B(net1090),
    .D(_0299_),
    .Q_N(_5699_),
    .Q(\logix.ram_r[1263] ));
 sg13g2_dfrbp_1 \logix.ram_r[1264]$_DFFE_PP_  (.CLK(net700),
    .RESET_B(net1091),
    .D(_0300_),
    .Q_N(_5698_),
    .Q(\logix.ram_r[1264] ));
 sg13g2_dfrbp_1 \logix.ram_r[1265]$_DFFE_PP_  (.CLK(net700),
    .RESET_B(net1092),
    .D(_0301_),
    .Q_N(_5697_),
    .Q(\logix.ram_r[1265] ));
 sg13g2_dfrbp_1 \logix.ram_r[1266]$_DFFE_PP_  (.CLK(net716),
    .RESET_B(net1093),
    .D(_0302_),
    .Q_N(_5696_),
    .Q(\logix.ram_r[1266] ));
 sg13g2_dfrbp_1 \logix.ram_r[1267]$_DFFE_PP_  (.CLK(net715),
    .RESET_B(net1094),
    .D(_0303_),
    .Q_N(_5695_),
    .Q(\logix.ram_r[1267] ));
 sg13g2_dfrbp_1 \logix.ram_r[1268]$_DFFE_PP_  (.CLK(net717),
    .RESET_B(net1095),
    .D(_0304_),
    .Q_N(_5694_),
    .Q(\logix.ram_r[1268] ));
 sg13g2_dfrbp_1 \logix.ram_r[1269]$_DFFE_PP_  (.CLK(net717),
    .RESET_B(net1096),
    .D(_0305_),
    .Q_N(_5693_),
    .Q(\logix.ram_r[1269] ));
 sg13g2_dfrbp_1 \logix.ram_r[126]$_DFFE_PP_  (.CLK(net697),
    .RESET_B(net1097),
    .D(_0306_),
    .Q_N(_5692_),
    .Q(\logix.ram_r[126] ));
 sg13g2_dfrbp_1 \logix.ram_r[1270]$_DFFE_PP_  (.CLK(net718),
    .RESET_B(net1098),
    .D(_0307_),
    .Q_N(_5691_),
    .Q(\logix.ram_r[1270] ));
 sg13g2_dfrbp_1 \logix.ram_r[1271]$_DFFE_PP_  (.CLK(net700),
    .RESET_B(net1099),
    .D(_0308_),
    .Q_N(_5690_),
    .Q(\logix.ram_r[1271] ));
 sg13g2_dfrbp_1 \logix.ram_r[1272]$_DFFE_PP_  (.CLK(net700),
    .RESET_B(net1100),
    .D(_0309_),
    .Q_N(_5689_),
    .Q(\logix.ram_r[1272] ));
 sg13g2_dfrbp_1 \logix.ram_r[1273]$_DFFE_PP_  (.CLK(net718),
    .RESET_B(net1101),
    .D(_0310_),
    .Q_N(_5688_),
    .Q(\logix.ram_r[1273] ));
 sg13g2_dfrbp_1 \logix.ram_r[1274]$_DFFE_PP_  (.CLK(net715),
    .RESET_B(net1102),
    .D(_0311_),
    .Q_N(_5687_),
    .Q(\logix.ram_r[1274] ));
 sg13g2_dfrbp_1 \logix.ram_r[1275]$_DFFE_PP_  (.CLK(net725),
    .RESET_B(net1103),
    .D(_0312_),
    .Q_N(_5686_),
    .Q(\logix.ram_r[1275] ));
 sg13g2_dfrbp_1 \logix.ram_r[1276]$_DFFE_PP_  (.CLK(net717),
    .RESET_B(net1104),
    .D(_0313_),
    .Q_N(_5685_),
    .Q(\logix.ram_r[1276] ));
 sg13g2_dfrbp_1 \logix.ram_r[1277]$_DFFE_PP_  (.CLK(net717),
    .RESET_B(net1105),
    .D(_0314_),
    .Q_N(_5684_),
    .Q(\logix.ram_r[1277] ));
 sg13g2_dfrbp_1 \logix.ram_r[1278]$_DFFE_PP_  (.CLK(net718),
    .RESET_B(net1106),
    .D(_0315_),
    .Q_N(_5683_),
    .Q(\logix.ram_r[1278] ));
 sg13g2_dfrbp_1 \logix.ram_r[1279]$_DFFE_PP_  (.CLK(net718),
    .RESET_B(net1107),
    .D(_0316_),
    .Q_N(_5682_),
    .Q(\logix.ram_r[1279] ));
 sg13g2_dfrbp_1 \logix.ram_r[127]$_DFFE_PP_  (.CLK(net697),
    .RESET_B(net1108),
    .D(_0317_),
    .Q_N(_5681_),
    .Q(\logix.ram_r[127] ));
 sg13g2_dfrbp_1 \logix.ram_r[1280]$_DFFE_PP_  (.CLK(net615),
    .RESET_B(net1109),
    .D(_0318_),
    .Q_N(_5680_),
    .Q(\logix.ram_r[1280] ));
 sg13g2_dfrbp_1 \logix.ram_r[1281]$_DFFE_PP_  (.CLK(net443),
    .RESET_B(net1110),
    .D(_0319_),
    .Q_N(_5679_),
    .Q(\logix.ram_r[1281] ));
 sg13g2_dfrbp_1 \logix.ram_r[1282]$_DFFE_PP_  (.CLK(net418),
    .RESET_B(net1111),
    .D(_0320_),
    .Q_N(_5678_),
    .Q(\logix.ram_r[1282] ));
 sg13g2_dfrbp_1 \logix.ram_r[1283]$_DFFE_PP_  (.CLK(net418),
    .RESET_B(net1112),
    .D(_0321_),
    .Q_N(_5677_),
    .Q(\logix.ram_r[1283] ));
 sg13g2_dfrbp_1 \logix.ram_r[1284]$_DFFE_PP_  (.CLK(net419),
    .RESET_B(net1113),
    .D(_0322_),
    .Q_N(_5676_),
    .Q(\logix.ram_r[1284] ));
 sg13g2_dfrbp_1 \logix.ram_r[1285]$_DFFE_PP_  (.CLK(net419),
    .RESET_B(net1114),
    .D(_0323_),
    .Q_N(_5675_),
    .Q(\logix.ram_r[1285] ));
 sg13g2_dfrbp_1 \logix.ram_r[1286]$_DFFE_PP_  (.CLK(net423),
    .RESET_B(net1115),
    .D(_0324_),
    .Q_N(_5674_),
    .Q(\logix.ram_r[1286] ));
 sg13g2_dfrbp_1 \logix.ram_r[1287]$_DFFE_PP_  (.CLK(net424),
    .RESET_B(net1116),
    .D(_0325_),
    .Q_N(_5673_),
    .Q(\logix.ram_r[1287] ));
 sg13g2_dfrbp_1 \logix.ram_r[1288]$_DFFE_PP_  (.CLK(net443),
    .RESET_B(net1117),
    .D(_0326_),
    .Q_N(_5672_),
    .Q(\logix.ram_r[1288] ));
 sg13g2_dfrbp_1 \logix.ram_r[1289]$_DFFE_PP_  (.CLK(net443),
    .RESET_B(net1118),
    .D(_0327_),
    .Q_N(_5671_),
    .Q(\logix.ram_r[1289] ));
 sg13g2_dfrbp_1 \logix.ram_r[128]$_DFFE_PP_  (.CLK(net543),
    .RESET_B(net1119),
    .D(_0328_),
    .Q_N(_5670_),
    .Q(\logix.ram_r[128] ));
 sg13g2_dfrbp_1 \logix.ram_r[1290]$_DFFE_PP_  (.CLK(net418),
    .RESET_B(net1120),
    .D(_0329_),
    .Q_N(_5669_),
    .Q(\logix.ram_r[1290] ));
 sg13g2_dfrbp_1 \logix.ram_r[1291]$_DFFE_PP_  (.CLK(net418),
    .RESET_B(net1121),
    .D(_0330_),
    .Q_N(_5668_),
    .Q(\logix.ram_r[1291] ));
 sg13g2_dfrbp_1 \logix.ram_r[1292]$_DFFE_PP_  (.CLK(net419),
    .RESET_B(net1122),
    .D(_0331_),
    .Q_N(_5667_),
    .Q(\logix.ram_r[1292] ));
 sg13g2_dfrbp_1 \logix.ram_r[1293]$_DFFE_PP_  (.CLK(net423),
    .RESET_B(net1123),
    .D(_0332_),
    .Q_N(_5666_),
    .Q(\logix.ram_r[1293] ));
 sg13g2_dfrbp_1 \logix.ram_r[1294]$_DFFE_PP_  (.CLK(net423),
    .RESET_B(net1124),
    .D(_0333_),
    .Q_N(_5665_),
    .Q(\logix.ram_r[1294] ));
 sg13g2_dfrbp_1 \logix.ram_r[1295]$_DFFE_PP_  (.CLK(net424),
    .RESET_B(net1125),
    .D(_0334_),
    .Q_N(_5664_),
    .Q(\logix.ram_r[1295] ));
 sg13g2_dfrbp_1 \logix.ram_r[1296]$_DFFE_PP_  (.CLK(net443),
    .RESET_B(net1126),
    .D(_0335_),
    .Q_N(_5663_),
    .Q(\logix.ram_r[1296] ));
 sg13g2_dfrbp_1 \logix.ram_r[1297]$_DFFE_PP_  (.CLK(net443),
    .RESET_B(net1127),
    .D(_0336_),
    .Q_N(_5662_),
    .Q(\logix.ram_r[1297] ));
 sg13g2_dfrbp_1 \logix.ram_r[1298]$_DFFE_PP_  (.CLK(net418),
    .RESET_B(net1128),
    .D(_0337_),
    .Q_N(_5661_),
    .Q(\logix.ram_r[1298] ));
 sg13g2_dfrbp_1 \logix.ram_r[1299]$_DFFE_PP_  (.CLK(net418),
    .RESET_B(net1129),
    .D(_0338_),
    .Q_N(_5660_),
    .Q(\logix.ram_r[1299] ));
 sg13g2_dfrbp_1 \logix.ram_r[129]$_DFFE_PP_  (.CLK(net539),
    .RESET_B(net1130),
    .D(_0339_),
    .Q_N(_5659_),
    .Q(\logix.ram_r[129] ));
 sg13g2_dfrbp_1 \logix.ram_r[12]$_DFFE_PP_  (.CLK(net634),
    .RESET_B(net1131),
    .D(_0340_),
    .Q_N(_5658_),
    .Q(\logix.ram_r[12] ));
 sg13g2_dfrbp_1 \logix.ram_r[1300]$_DFFE_PP_  (.CLK(net419),
    .RESET_B(net1132),
    .D(_0341_),
    .Q_N(_5657_),
    .Q(\logix.ram_r[1300] ));
 sg13g2_dfrbp_1 \logix.ram_r[1301]$_DFFE_PP_  (.CLK(net423),
    .RESET_B(net1133),
    .D(_0342_),
    .Q_N(_5656_),
    .Q(\logix.ram_r[1301] ));
 sg13g2_dfrbp_1 \logix.ram_r[1302]$_DFFE_PP_  (.CLK(net423),
    .RESET_B(net1134),
    .D(_0343_),
    .Q_N(_5655_),
    .Q(\logix.ram_r[1302] ));
 sg13g2_dfrbp_1 \logix.ram_r[1303]$_DFFE_PP_  (.CLK(net424),
    .RESET_B(net1135),
    .D(_0344_),
    .Q_N(_5654_),
    .Q(\logix.ram_r[1303] ));
 sg13g2_dfrbp_1 \logix.ram_r[1304]$_DFFE_PP_  (.CLK(net443),
    .RESET_B(net1136),
    .D(_0345_),
    .Q_N(_5653_),
    .Q(\logix.ram_r[1304] ));
 sg13g2_dfrbp_1 \logix.ram_r[1305]$_DFFE_PP_  (.CLK(net443),
    .RESET_B(net1137),
    .D(_0346_),
    .Q_N(_5652_),
    .Q(\logix.ram_r[1305] ));
 sg13g2_dfrbp_1 \logix.ram_r[1306]$_DFFE_PP_  (.CLK(net419),
    .RESET_B(net1138),
    .D(_0347_),
    .Q_N(_5651_),
    .Q(\logix.ram_r[1306] ));
 sg13g2_dfrbp_1 \logix.ram_r[1307]$_DFFE_PP_  (.CLK(net419),
    .RESET_B(net1139),
    .D(_0348_),
    .Q_N(_5650_),
    .Q(\logix.ram_r[1307] ));
 sg13g2_dfrbp_1 \logix.ram_r[1308]$_DFFE_PP_  (.CLK(net419),
    .RESET_B(net1140),
    .D(_0349_),
    .Q_N(_5649_),
    .Q(\logix.ram_r[1308] ));
 sg13g2_dfrbp_1 \logix.ram_r[1309]$_DFFE_PP_  (.CLK(net423),
    .RESET_B(net1141),
    .D(_0350_),
    .Q_N(_5648_),
    .Q(\logix.ram_r[1309] ));
 sg13g2_dfrbp_1 \logix.ram_r[130]$_DFFE_PP_  (.CLK(net518),
    .RESET_B(net1142),
    .D(_0351_),
    .Q_N(_5647_),
    .Q(\logix.ram_r[130] ));
 sg13g2_dfrbp_1 \logix.ram_r[1310]$_DFFE_PP_  (.CLK(net424),
    .RESET_B(net1143),
    .D(_0352_),
    .Q_N(_5646_),
    .Q(\logix.ram_r[1310] ));
 sg13g2_dfrbp_1 \logix.ram_r[1311]$_DFFE_PP_  (.CLK(net424),
    .RESET_B(net1144),
    .D(_0353_),
    .Q_N(_5645_),
    .Q(\logix.ram_r[1311] ));
 sg13g2_dfrbp_1 \logix.ram_r[1312]$_DFFE_PP_  (.CLK(net451),
    .RESET_B(net1145),
    .D(_0354_),
    .Q_N(_5644_),
    .Q(\logix.ram_r[1312] ));
 sg13g2_dfrbp_1 \logix.ram_r[1313]$_DFFE_PP_  (.CLK(net451),
    .RESET_B(net1146),
    .D(_0355_),
    .Q_N(_5643_),
    .Q(\logix.ram_r[1313] ));
 sg13g2_dfrbp_1 \logix.ram_r[1314]$_DFFE_PP_  (.CLK(net426),
    .RESET_B(net1147),
    .D(_0356_),
    .Q_N(_5642_),
    .Q(\logix.ram_r[1314] ));
 sg13g2_dfrbp_1 \logix.ram_r[1315]$_DFFE_PP_  (.CLK(net426),
    .RESET_B(net1148),
    .D(_0357_),
    .Q_N(_5641_),
    .Q(\logix.ram_r[1315] ));
 sg13g2_dfrbp_1 \logix.ram_r[1316]$_DFFE_PP_  (.CLK(net426),
    .RESET_B(net1149),
    .D(_0358_),
    .Q_N(_5640_),
    .Q(\logix.ram_r[1316] ));
 sg13g2_dfrbp_1 \logix.ram_r[1317]$_DFFE_PP_  (.CLK(net433),
    .RESET_B(net1150),
    .D(_0359_),
    .Q_N(_5639_),
    .Q(\logix.ram_r[1317] ));
 sg13g2_dfrbp_1 \logix.ram_r[1318]$_DFFE_PP_  (.CLK(net434),
    .RESET_B(net1151),
    .D(_0360_),
    .Q_N(_5638_),
    .Q(\logix.ram_r[1318] ));
 sg13g2_dfrbp_1 \logix.ram_r[1319]$_DFFE_PP_  (.CLK(net434),
    .RESET_B(net1152),
    .D(_0361_),
    .Q_N(_5637_),
    .Q(\logix.ram_r[1319] ));
 sg13g2_dfrbp_1 \logix.ram_r[131]$_DFFE_PP_  (.CLK(net519),
    .RESET_B(net1153),
    .D(_0362_),
    .Q_N(_5636_),
    .Q(\logix.ram_r[131] ));
 sg13g2_dfrbp_1 \logix.ram_r[1320]$_DFFE_PP_  (.CLK(net451),
    .RESET_B(net1154),
    .D(_0363_),
    .Q_N(_5635_),
    .Q(\logix.ram_r[1320] ));
 sg13g2_dfrbp_1 \logix.ram_r[1321]$_DFFE_PP_  (.CLK(net451),
    .RESET_B(net1155),
    .D(_0364_),
    .Q_N(_5634_),
    .Q(\logix.ram_r[1321] ));
 sg13g2_dfrbp_1 \logix.ram_r[1322]$_DFFE_PP_  (.CLK(net426),
    .RESET_B(net1156),
    .D(_0365_),
    .Q_N(_5633_),
    .Q(\logix.ram_r[1322] ));
 sg13g2_dfrbp_1 \logix.ram_r[1323]$_DFFE_PP_  (.CLK(net426),
    .RESET_B(net1157),
    .D(_0366_),
    .Q_N(_5632_),
    .Q(\logix.ram_r[1323] ));
 sg13g2_dfrbp_1 \logix.ram_r[1324]$_DFFE_PP_  (.CLK(net428),
    .RESET_B(net1158),
    .D(_0367_),
    .Q_N(_5631_),
    .Q(\logix.ram_r[1324] ));
 sg13g2_dfrbp_1 \logix.ram_r[1325]$_DFFE_PP_  (.CLK(net433),
    .RESET_B(net1159),
    .D(_0368_),
    .Q_N(_5630_),
    .Q(\logix.ram_r[1325] ));
 sg13g2_dfrbp_1 \logix.ram_r[1326]$_DFFE_PP_  (.CLK(net434),
    .RESET_B(net1160),
    .D(_0369_),
    .Q_N(_5629_),
    .Q(\logix.ram_r[1326] ));
 sg13g2_dfrbp_1 \logix.ram_r[1327]$_DFFE_PP_  (.CLK(net451),
    .RESET_B(net1161),
    .D(_0370_),
    .Q_N(_5628_),
    .Q(\logix.ram_r[1327] ));
 sg13g2_dfrbp_1 \logix.ram_r[1328]$_DFFE_PP_  (.CLK(net452),
    .RESET_B(net1162),
    .D(_0371_),
    .Q_N(_5627_),
    .Q(\logix.ram_r[1328] ));
 sg13g2_dfrbp_1 \logix.ram_r[1329]$_DFFE_PP_  (.CLK(net451),
    .RESET_B(net1163),
    .D(_0372_),
    .Q_N(_5626_),
    .Q(\logix.ram_r[1329] ));
 sg13g2_dfrbp_1 \logix.ram_r[132]$_DFFE_PP_  (.CLK(net519),
    .RESET_B(net1164),
    .D(_0373_),
    .Q_N(_5625_),
    .Q(\logix.ram_r[132] ));
 sg13g2_dfrbp_1 \logix.ram_r[1330]$_DFFE_PP_  (.CLK(net426),
    .RESET_B(net1165),
    .D(_0374_),
    .Q_N(_5624_),
    .Q(\logix.ram_r[1330] ));
 sg13g2_dfrbp_1 \logix.ram_r[1331]$_DFFE_PP_  (.CLK(net426),
    .RESET_B(net1166),
    .D(_0375_),
    .Q_N(_5623_),
    .Q(\logix.ram_r[1331] ));
 sg13g2_dfrbp_1 \logix.ram_r[1332]$_DFFE_PP_  (.CLK(net428),
    .RESET_B(net1167),
    .D(_0376_),
    .Q_N(_5622_),
    .Q(\logix.ram_r[1332] ));
 sg13g2_dfrbp_1 \logix.ram_r[1333]$_DFFE_PP_  (.CLK(net433),
    .RESET_B(net1168),
    .D(_0377_),
    .Q_N(_5621_),
    .Q(\logix.ram_r[1333] ));
 sg13g2_dfrbp_1 \logix.ram_r[1334]$_DFFE_PP_  (.CLK(net434),
    .RESET_B(net1169),
    .D(_0378_),
    .Q_N(_5620_),
    .Q(\logix.ram_r[1334] ));
 sg13g2_dfrbp_1 \logix.ram_r[1335]$_DFFE_PP_  (.CLK(net434),
    .RESET_B(net1170),
    .D(_0379_),
    .Q_N(_5619_),
    .Q(\logix.ram_r[1335] ));
 sg13g2_dfrbp_1 \logix.ram_r[1336]$_DFFE_PP_  (.CLK(net451),
    .RESET_B(net1171),
    .D(_0380_),
    .Q_N(_5618_),
    .Q(\logix.ram_r[1336] ));
 sg13g2_dfrbp_1 \logix.ram_r[1337]$_DFFE_PP_  (.CLK(net451),
    .RESET_B(net1172),
    .D(_0381_),
    .Q_N(_5617_),
    .Q(\logix.ram_r[1337] ));
 sg13g2_dfrbp_1 \logix.ram_r[1338]$_DFFE_PP_  (.CLK(net433),
    .RESET_B(net1173),
    .D(_0382_),
    .Q_N(_5616_),
    .Q(\logix.ram_r[1338] ));
 sg13g2_dfrbp_1 \logix.ram_r[1339]$_DFFE_PP_  (.CLK(net428),
    .RESET_B(net1174),
    .D(_0383_),
    .Q_N(_5615_),
    .Q(\logix.ram_r[1339] ));
 sg13g2_dfrbp_1 \logix.ram_r[133]$_DFFE_PP_  (.CLK(net518),
    .RESET_B(net1175),
    .D(_0384_),
    .Q_N(_5614_),
    .Q(\logix.ram_r[133] ));
 sg13g2_dfrbp_1 \logix.ram_r[1340]$_DFFE_PP_  (.CLK(net428),
    .RESET_B(net1176),
    .D(_0385_),
    .Q_N(_5613_),
    .Q(\logix.ram_r[1340] ));
 sg13g2_dfrbp_1 \logix.ram_r[1341]$_DFFE_PP_  (.CLK(net433),
    .RESET_B(net1177),
    .D(_0386_),
    .Q_N(_5612_),
    .Q(\logix.ram_r[1341] ));
 sg13g2_dfrbp_1 \logix.ram_r[1342]$_DFFE_PP_  (.CLK(net437),
    .RESET_B(net1178),
    .D(_0387_),
    .Q_N(_5611_),
    .Q(\logix.ram_r[1342] ));
 sg13g2_dfrbp_1 \logix.ram_r[1343]$_DFFE_PP_  (.CLK(net437),
    .RESET_B(net1179),
    .D(_0388_),
    .Q_N(_5610_),
    .Q(\logix.ram_r[1343] ));
 sg13g2_dfrbp_1 \logix.ram_r[1344]$_DFFE_PP_  (.CLK(net467),
    .RESET_B(net1180),
    .D(_0389_),
    .Q_N(_5609_),
    .Q(\logix.ram_r[1344] ));
 sg13g2_dfrbp_1 \logix.ram_r[1345]$_DFFE_PP_  (.CLK(net483),
    .RESET_B(net1181),
    .D(_0390_),
    .Q_N(_5608_),
    .Q(\logix.ram_r[1345] ));
 sg13g2_dfrbp_1 \logix.ram_r[1346]$_DFFE_PP_  (.CLK(net483),
    .RESET_B(net1182),
    .D(_0391_),
    .Q_N(_5607_),
    .Q(\logix.ram_r[1346] ));
 sg13g2_dfrbp_1 \logix.ram_r[1347]$_DFFE_PP_  (.CLK(net478),
    .RESET_B(net1183),
    .D(_0392_),
    .Q_N(_5606_),
    .Q(\logix.ram_r[1347] ));
 sg13g2_dfrbp_1 \logix.ram_r[1348]$_DFFE_PP_  (.CLK(net480),
    .RESET_B(net1184),
    .D(_0393_),
    .Q_N(_5605_),
    .Q(\logix.ram_r[1348] ));
 sg13g2_dfrbp_1 \logix.ram_r[1349]$_DFFE_PP_  (.CLK(net480),
    .RESET_B(net1185),
    .D(_0394_),
    .Q_N(_5604_),
    .Q(\logix.ram_r[1349] ));
 sg13g2_dfrbp_1 \logix.ram_r[134]$_DFFE_PP_  (.CLK(net521),
    .RESET_B(net1186),
    .D(_0395_),
    .Q_N(_5603_),
    .Q(\logix.ram_r[134] ));
 sg13g2_dfrbp_1 \logix.ram_r[1350]$_DFFE_PP_  (.CLK(net480),
    .RESET_B(net1187),
    .D(_0396_),
    .Q_N(_5602_),
    .Q(\logix.ram_r[1350] ));
 sg13g2_dfrbp_1 \logix.ram_r[1351]$_DFFE_PP_  (.CLK(net495),
    .RESET_B(net1188),
    .D(_0397_),
    .Q_N(_5601_),
    .Q(\logix.ram_r[1351] ));
 sg13g2_dfrbp_1 \logix.ram_r[1352]$_DFFE_PP_  (.CLK(net495),
    .RESET_B(net1189),
    .D(_0398_),
    .Q_N(_5600_),
    .Q(\logix.ram_r[1352] ));
 sg13g2_dfrbp_1 \logix.ram_r[1353]$_DFFE_PP_  (.CLK(net480),
    .RESET_B(net1190),
    .D(_0399_),
    .Q_N(_5599_),
    .Q(\logix.ram_r[1353] ));
 sg13g2_dfrbp_1 \logix.ram_r[1354]$_DFFE_PP_  (.CLK(net481),
    .RESET_B(net1191),
    .D(_0400_),
    .Q_N(_5598_),
    .Q(\logix.ram_r[1354] ));
 sg13g2_dfrbp_1 \logix.ram_r[1355]$_DFFE_PP_  (.CLK(net475),
    .RESET_B(net1192),
    .D(_0401_),
    .Q_N(_5597_),
    .Q(\logix.ram_r[1355] ));
 sg13g2_dfrbp_1 \logix.ram_r[1356]$_DFFE_PP_  (.CLK(net475),
    .RESET_B(net1193),
    .D(_0402_),
    .Q_N(_5596_),
    .Q(\logix.ram_r[1356] ));
 sg13g2_dfrbp_1 \logix.ram_r[1357]$_DFFE_PP_  (.CLK(net480),
    .RESET_B(net1194),
    .D(_0403_),
    .Q_N(_5595_),
    .Q(\logix.ram_r[1357] ));
 sg13g2_dfrbp_1 \logix.ram_r[1358]$_DFFE_PP_  (.CLK(net480),
    .RESET_B(net1195),
    .D(_0404_),
    .Q_N(_5594_),
    .Q(\logix.ram_r[1358] ));
 sg13g2_dfrbp_1 \logix.ram_r[1359]$_DFFE_PP_  (.CLK(net481),
    .RESET_B(net1196),
    .D(_0405_),
    .Q_N(_5593_),
    .Q(\logix.ram_r[1359] ));
 sg13g2_dfrbp_1 \logix.ram_r[135]$_DFFE_PP_  (.CLK(net458),
    .RESET_B(net1197),
    .D(_0406_),
    .Q_N(_5592_),
    .Q(\logix.ram_r[135] ));
 sg13g2_dfrbp_1 \logix.ram_r[1360]$_DFFE_PP_  (.CLK(net483),
    .RESET_B(net1198),
    .D(_0407_),
    .Q_N(_5591_),
    .Q(\logix.ram_r[1360] ));
 sg13g2_dfrbp_1 \logix.ram_r[1361]$_DFFE_PP_  (.CLK(net483),
    .RESET_B(net1199),
    .D(_0408_),
    .Q_N(_5590_),
    .Q(\logix.ram_r[1361] ));
 sg13g2_dfrbp_1 \logix.ram_r[1362]$_DFFE_PP_  (.CLK(net482),
    .RESET_B(net1200),
    .D(_0409_),
    .Q_N(_5589_),
    .Q(\logix.ram_r[1362] ));
 sg13g2_dfrbp_1 \logix.ram_r[1363]$_DFFE_PP_  (.CLK(net478),
    .RESET_B(net1201),
    .D(_0410_),
    .Q_N(_5588_),
    .Q(\logix.ram_r[1363] ));
 sg13g2_dfrbp_1 \logix.ram_r[1364]$_DFFE_PP_  (.CLK(net478),
    .RESET_B(net1202),
    .D(_0411_),
    .Q_N(_5587_),
    .Q(\logix.ram_r[1364] ));
 sg13g2_dfrbp_1 \logix.ram_r[1365]$_DFFE_PP_  (.CLK(net477),
    .RESET_B(net1203),
    .D(_0412_),
    .Q_N(_5586_),
    .Q(\logix.ram_r[1365] ));
 sg13g2_dfrbp_1 \logix.ram_r[1366]$_DFFE_PP_  (.CLK(net482),
    .RESET_B(net1204),
    .D(_0413_),
    .Q_N(_5585_),
    .Q(\logix.ram_r[1366] ));
 sg13g2_dfrbp_1 \logix.ram_r[1367]$_DFFE_PP_  (.CLK(net482),
    .RESET_B(net1205),
    .D(_0414_),
    .Q_N(_5584_),
    .Q(\logix.ram_r[1367] ));
 sg13g2_dfrbp_1 \logix.ram_r[1368]$_DFFE_PP_  (.CLK(net483),
    .RESET_B(net1206),
    .D(_0415_),
    .Q_N(_5583_),
    .Q(\logix.ram_r[1368] ));
 sg13g2_dfrbp_1 \logix.ram_r[1369]$_DFFE_PP_  (.CLK(net483),
    .RESET_B(net1207),
    .D(_0416_),
    .Q_N(_5582_),
    .Q(\logix.ram_r[1369] ));
 sg13g2_dfrbp_1 \logix.ram_r[136]$_DFFE_PP_  (.CLK(net491),
    .RESET_B(net1208),
    .D(_0417_),
    .Q_N(_5581_),
    .Q(\logix.ram_r[136] ));
 sg13g2_dfrbp_1 \logix.ram_r[1370]$_DFFE_PP_  (.CLK(net484),
    .RESET_B(net1209),
    .D(_0418_),
    .Q_N(_5580_),
    .Q(\logix.ram_r[1370] ));
 sg13g2_dfrbp_1 \logix.ram_r[1371]$_DFFE_PP_  (.CLK(net477),
    .RESET_B(net1210),
    .D(_0419_),
    .Q_N(_5579_),
    .Q(\logix.ram_r[1371] ));
 sg13g2_dfrbp_1 \logix.ram_r[1372]$_DFFE_PP_  (.CLK(net477),
    .RESET_B(net1211),
    .D(_0420_),
    .Q_N(_5578_),
    .Q(\logix.ram_r[1372] ));
 sg13g2_dfrbp_1 \logix.ram_r[1373]$_DFFE_PP_  (.CLK(net477),
    .RESET_B(net1212),
    .D(_0421_),
    .Q_N(_5577_),
    .Q(\logix.ram_r[1373] ));
 sg13g2_dfrbp_1 \logix.ram_r[1374]$_DFFE_PP_  (.CLK(net478),
    .RESET_B(net1213),
    .D(_0422_),
    .Q_N(_5576_),
    .Q(\logix.ram_r[1374] ));
 sg13g2_dfrbp_1 \logix.ram_r[1375]$_DFFE_PP_  (.CLK(net478),
    .RESET_B(net1214),
    .D(_0423_),
    .Q_N(_5575_),
    .Q(\logix.ram_r[1375] ));
 sg13g2_dfrbp_1 \logix.ram_r[1376]$_DFFE_PP_  (.CLK(net477),
    .RESET_B(net1215),
    .D(_0424_),
    .Q_N(_5574_),
    .Q(\logix.ram_r[1376] ));
 sg13g2_dfrbp_1 \logix.ram_r[1377]$_DFFE_PP_  (.CLK(net476),
    .RESET_B(net1216),
    .D(_0425_),
    .Q_N(_5573_),
    .Q(\logix.ram_r[1377] ));
 sg13g2_dfrbp_1 \logix.ram_r[1378]$_DFFE_PP_  (.CLK(net476),
    .RESET_B(net1217),
    .D(_0426_),
    .Q_N(_5572_),
    .Q(\logix.ram_r[1378] ));
 sg13g2_dfrbp_1 \logix.ram_r[1379]$_DFFE_PP_  (.CLK(net473),
    .RESET_B(net1218),
    .D(_0427_),
    .Q_N(_5571_),
    .Q(\logix.ram_r[1379] ));
 sg13g2_dfrbp_1 \logix.ram_r[137]$_DFFE_PP_  (.CLK(net494),
    .RESET_B(net1219),
    .D(_0428_),
    .Q_N(_5570_),
    .Q(\logix.ram_r[137] ));
 sg13g2_dfrbp_1 \logix.ram_r[1380]$_DFFE_PP_  (.CLK(net473),
    .RESET_B(net1220),
    .D(_0429_),
    .Q_N(_5569_),
    .Q(\logix.ram_r[1380] ));
 sg13g2_dfrbp_1 \logix.ram_r[1381]$_DFFE_PP_  (.CLK(net476),
    .RESET_B(net1221),
    .D(_0430_),
    .Q_N(_5568_),
    .Q(\logix.ram_r[1381] ));
 sg13g2_dfrbp_1 \logix.ram_r[1382]$_DFFE_PP_  (.CLK(net476),
    .RESET_B(net1222),
    .D(_0431_),
    .Q_N(_5567_),
    .Q(\logix.ram_r[1382] ));
 sg13g2_dfrbp_1 \logix.ram_r[1383]$_DFFE_PP_  (.CLK(net476),
    .RESET_B(net1223),
    .D(_0432_),
    .Q_N(_5566_),
    .Q(\logix.ram_r[1383] ));
 sg13g2_dfrbp_1 \logix.ram_r[1384]$_DFFE_PP_  (.CLK(net474),
    .RESET_B(net1224),
    .D(_0433_),
    .Q_N(_5565_),
    .Q(\logix.ram_r[1384] ));
 sg13g2_dfrbp_1 \logix.ram_r[1385]$_DFFE_PP_  (.CLK(net474),
    .RESET_B(net1225),
    .D(_0434_),
    .Q_N(_5564_),
    .Q(\logix.ram_r[1385] ));
 sg13g2_dfrbp_1 \logix.ram_r[1386]$_DFFE_PP_  (.CLK(net474),
    .RESET_B(net1226),
    .D(_0435_),
    .Q_N(_5563_),
    .Q(\logix.ram_r[1386] ));
 sg13g2_dfrbp_1 \logix.ram_r[1387]$_DFFE_PP_  (.CLK(net475),
    .RESET_B(net1227),
    .D(_0436_),
    .Q_N(_5562_),
    .Q(\logix.ram_r[1387] ));
 sg13g2_dfrbp_1 \logix.ram_r[1388]$_DFFE_PP_  (.CLK(net474),
    .RESET_B(net1228),
    .D(_0437_),
    .Q_N(_5561_),
    .Q(\logix.ram_r[1388] ));
 sg13g2_dfrbp_1 \logix.ram_r[1389]$_DFFE_PP_  (.CLK(net476),
    .RESET_B(net1229),
    .D(_0438_),
    .Q_N(_5560_),
    .Q(\logix.ram_r[1389] ));
 sg13g2_dfrbp_1 \logix.ram_r[138]$_DFFE_PP_  (.CLK(net494),
    .RESET_B(net1230),
    .D(_0439_),
    .Q_N(_5559_),
    .Q(\logix.ram_r[138] ));
 sg13g2_dfrbp_1 \logix.ram_r[1390]$_DFFE_PP_  (.CLK(net476),
    .RESET_B(net1231),
    .D(_0440_),
    .Q_N(_5558_),
    .Q(\logix.ram_r[1390] ));
 sg13g2_dfrbp_1 \logix.ram_r[1391]$_DFFE_PP_  (.CLK(net476),
    .RESET_B(net1232),
    .D(_0441_),
    .Q_N(_5557_),
    .Q(\logix.ram_r[1391] ));
 sg13g2_dfrbp_1 \logix.ram_r[1392]$_DFFE_PP_  (.CLK(net483),
    .RESET_B(net1233),
    .D(_0442_),
    .Q_N(_5556_),
    .Q(\logix.ram_r[1392] ));
 sg13g2_dfrbp_1 \logix.ram_r[1393]$_DFFE_PP_  (.CLK(net482),
    .RESET_B(net1234),
    .D(_0443_),
    .Q_N(_5555_),
    .Q(\logix.ram_r[1393] ));
 sg13g2_dfrbp_1 \logix.ram_r[1394]$_DFFE_PP_  (.CLK(net478),
    .RESET_B(net1235),
    .D(_0444_),
    .Q_N(_5554_),
    .Q(\logix.ram_r[1394] ));
 sg13g2_dfrbp_1 \logix.ram_r[1395]$_DFFE_PP_  (.CLK(net479),
    .RESET_B(net1236),
    .D(_0445_),
    .Q_N(_5553_),
    .Q(\logix.ram_r[1395] ));
 sg13g2_dfrbp_1 \logix.ram_r[1396]$_DFFE_PP_  (.CLK(net482),
    .RESET_B(net1237),
    .D(_0446_),
    .Q_N(_5552_),
    .Q(\logix.ram_r[1396] ));
 sg13g2_dfrbp_1 \logix.ram_r[1397]$_DFFE_PP_  (.CLK(net482),
    .RESET_B(net1238),
    .D(_0447_),
    .Q_N(_5551_),
    .Q(\logix.ram_r[1397] ));
 sg13g2_dfrbp_1 \logix.ram_r[1398]$_DFFE_PP_  (.CLK(net497),
    .RESET_B(net1239),
    .D(_0448_),
    .Q_N(_5550_),
    .Q(\logix.ram_r[1398] ));
 sg13g2_dfrbp_1 \logix.ram_r[1399]$_DFFE_PP_  (.CLK(net497),
    .RESET_B(net1240),
    .D(_0449_),
    .Q_N(_5549_),
    .Q(\logix.ram_r[1399] ));
 sg13g2_dfrbp_1 \logix.ram_r[139]$_DFFE_PP_  (.CLK(net570),
    .RESET_B(net1241),
    .D(_0450_),
    .Q_N(_5548_),
    .Q(\logix.ram_r[139] ));
 sg13g2_dfrbp_1 \logix.ram_r[13]$_DFFE_PP_  (.CLK(net634),
    .RESET_B(net1242),
    .D(_0451_),
    .Q_N(_5547_),
    .Q(\logix.ram_r[13] ));
 sg13g2_dfrbp_1 \logix.ram_r[1400]$_DFFE_PP_  (.CLK(net483),
    .RESET_B(net1243),
    .D(_0452_),
    .Q_N(_5546_),
    .Q(\logix.ram_r[1400] ));
 sg13g2_dfrbp_1 \logix.ram_r[1401]$_DFFE_PP_  (.CLK(net484),
    .RESET_B(net1244),
    .D(_0453_),
    .Q_N(_5545_),
    .Q(\logix.ram_r[1401] ));
 sg13g2_dfrbp_1 \logix.ram_r[1402]$_DFFE_PP_  (.CLK(net479),
    .RESET_B(net1245),
    .D(_0454_),
    .Q_N(_5544_),
    .Q(\logix.ram_r[1402] ));
 sg13g2_dfrbp_1 \logix.ram_r[1403]$_DFFE_PP_  (.CLK(net482),
    .RESET_B(net1246),
    .D(_0455_),
    .Q_N(_5543_),
    .Q(\logix.ram_r[1403] ));
 sg13g2_dfrbp_1 \logix.ram_r[1404]$_DFFE_PP_  (.CLK(net482),
    .RESET_B(net1247),
    .D(_0456_),
    .Q_N(_5542_),
    .Q(\logix.ram_r[1404] ));
 sg13g2_dfrbp_1 \logix.ram_r[1405]$_DFFE_PP_  (.CLK(net497),
    .RESET_B(net1248),
    .D(_0457_),
    .Q_N(_5541_),
    .Q(\logix.ram_r[1405] ));
 sg13g2_dfrbp_1 \logix.ram_r[1406]$_DFFE_PP_  (.CLK(net497),
    .RESET_B(net1249),
    .D(_0458_),
    .Q_N(_5540_),
    .Q(\logix.ram_r[1406] ));
 sg13g2_dfrbp_1 \logix.ram_r[1407]$_DFFE_PP_  (.CLK(net497),
    .RESET_B(net1250),
    .D(_0459_),
    .Q_N(_5539_),
    .Q(\logix.ram_r[1407] ));
 sg13g2_dfrbp_1 \logix.ram_r[1408]$_DFFE_PP_  (.CLK(net495),
    .RESET_B(net1251),
    .D(_0460_),
    .Q_N(_5538_),
    .Q(\logix.ram_r[1408] ));
 sg13g2_dfrbp_1 \logix.ram_r[1409]$_DFFE_PP_  (.CLK(net651),
    .RESET_B(net1252),
    .D(_0461_),
    .Q_N(_5537_),
    .Q(\logix.ram_r[1409] ));
 sg13g2_dfrbp_1 \logix.ram_r[140]$_DFFE_PP_  (.CLK(net570),
    .RESET_B(net1253),
    .D(_0462_),
    .Q_N(_5536_),
    .Q(\logix.ram_r[140] ));
 sg13g2_dfrbp_1 \logix.ram_r[1410]$_DFFE_PP_  (.CLK(net651),
    .RESET_B(net1254),
    .D(_0463_),
    .Q_N(_5535_),
    .Q(\logix.ram_r[1410] ));
 sg13g2_dfrbp_1 \logix.ram_r[1411]$_DFFE_PP_  (.CLK(net642),
    .RESET_B(net1255),
    .D(_0464_),
    .Q_N(_5534_),
    .Q(\logix.ram_r[1411] ));
 sg13g2_dfrbp_1 \logix.ram_r[1412]$_DFFE_PP_  (.CLK(net642),
    .RESET_B(net1256),
    .D(_0465_),
    .Q_N(_5533_),
    .Q(\logix.ram_r[1412] ));
 sg13g2_dfrbp_1 \logix.ram_r[1413]$_DFFE_PP_  (.CLK(net641),
    .RESET_B(net1257),
    .D(_0466_),
    .Q_N(_5532_),
    .Q(\logix.ram_r[1413] ));
 sg13g2_dfrbp_1 \logix.ram_r[1414]$_DFFE_PP_  (.CLK(net636),
    .RESET_B(net1258),
    .D(_0467_),
    .Q_N(_5531_),
    .Q(\logix.ram_r[1414] ));
 sg13g2_dfrbp_1 \logix.ram_r[1415]$_DFFE_PP_  (.CLK(net652),
    .RESET_B(net1259),
    .D(_0468_),
    .Q_N(_5530_),
    .Q(\logix.ram_r[1415] ));
 sg13g2_dfrbp_1 \logix.ram_r[1416]$_DFFE_PP_  (.CLK(net651),
    .RESET_B(net1260),
    .D(_0469_),
    .Q_N(_5529_),
    .Q(\logix.ram_r[1416] ));
 sg13g2_dfrbp_1 \logix.ram_r[1417]$_DFFE_PP_  (.CLK(net651),
    .RESET_B(net1261),
    .D(_0470_),
    .Q_N(_5528_),
    .Q(\logix.ram_r[1417] ));
 sg13g2_dfrbp_1 \logix.ram_r[1418]$_DFFE_PP_  (.CLK(net668),
    .RESET_B(net1262),
    .D(_0471_),
    .Q_N(_5527_),
    .Q(\logix.ram_r[1418] ));
 sg13g2_dfrbp_1 \logix.ram_r[1419]$_DFFE_PP_  (.CLK(net659),
    .RESET_B(net1263),
    .D(_0472_),
    .Q_N(_5526_),
    .Q(\logix.ram_r[1419] ));
 sg13g2_dfrbp_1 \logix.ram_r[141]$_DFFE_PP_  (.CLK(net571),
    .RESET_B(net1264),
    .D(_0473_),
    .Q_N(_5525_),
    .Q(\logix.ram_r[141] ));
 sg13g2_dfrbp_1 \logix.ram_r[1420]$_DFFE_PP_  (.CLK(net659),
    .RESET_B(net1265),
    .D(_0474_),
    .Q_N(_5524_),
    .Q(\logix.ram_r[1420] ));
 sg13g2_dfrbp_1 \logix.ram_r[1421]$_DFFE_PP_  (.CLK(net642),
    .RESET_B(net1266),
    .D(_0475_),
    .Q_N(_5523_),
    .Q(\logix.ram_r[1421] ));
 sg13g2_dfrbp_1 \logix.ram_r[1422]$_DFFE_PP_  (.CLK(net652),
    .RESET_B(net1267),
    .D(_0476_),
    .Q_N(_5522_),
    .Q(\logix.ram_r[1422] ));
 sg13g2_dfrbp_1 \logix.ram_r[1423]$_DFFE_PP_  (.CLK(net652),
    .RESET_B(net1268),
    .D(_0477_),
    .Q_N(_5521_),
    .Q(\logix.ram_r[1423] ));
 sg13g2_dfrbp_1 \logix.ram_r[1424]$_DFFE_PP_  (.CLK(net651),
    .RESET_B(net1269),
    .D(_0478_),
    .Q_N(_5520_),
    .Q(\logix.ram_r[1424] ));
 sg13g2_dfrbp_1 \logix.ram_r[1425]$_DFFE_PP_  (.CLK(net651),
    .RESET_B(net1270),
    .D(_0479_),
    .Q_N(_5519_),
    .Q(\logix.ram_r[1425] ));
 sg13g2_dfrbp_1 \logix.ram_r[1426]$_DFFE_PP_  (.CLK(net668),
    .RESET_B(net1271),
    .D(_0480_),
    .Q_N(_5518_),
    .Q(\logix.ram_r[1426] ));
 sg13g2_dfrbp_1 \logix.ram_r[1427]$_DFFE_PP_  (.CLK(net642),
    .RESET_B(net1272),
    .D(_0481_),
    .Q_N(_5517_),
    .Q(\logix.ram_r[1427] ));
 sg13g2_dfrbp_1 \logix.ram_r[1428]$_DFFE_PP_  (.CLK(net643),
    .RESET_B(net1273),
    .D(_0482_),
    .Q_N(_5516_),
    .Q(\logix.ram_r[1428] ));
 sg13g2_dfrbp_1 \logix.ram_r[1429]$_DFFE_PP_  (.CLK(net643),
    .RESET_B(net1274),
    .D(_0483_),
    .Q_N(_5515_),
    .Q(\logix.ram_r[1429] ));
 sg13g2_dfrbp_1 \logix.ram_r[142]$_DFFE_PP_  (.CLK(net545),
    .RESET_B(net1275),
    .D(_0484_),
    .Q_N(_5514_),
    .Q(\logix.ram_r[142] ));
 sg13g2_dfrbp_1 \logix.ram_r[1430]$_DFFE_PP_  (.CLK(net637),
    .RESET_B(net1276),
    .D(_0485_),
    .Q_N(_5513_),
    .Q(\logix.ram_r[1430] ));
 sg13g2_dfrbp_1 \logix.ram_r[1431]$_DFFE_PP_  (.CLK(net652),
    .RESET_B(net1277),
    .D(_0486_),
    .Q_N(_5512_),
    .Q(\logix.ram_r[1431] ));
 sg13g2_dfrbp_1 \logix.ram_r[1432]$_DFFE_PP_  (.CLK(net652),
    .RESET_B(net1278),
    .D(_0487_),
    .Q_N(_5511_),
    .Q(\logix.ram_r[1432] ));
 sg13g2_dfrbp_1 \logix.ram_r[1433]$_DFFE_PP_  (.CLK(net651),
    .RESET_B(net1279),
    .D(_0488_),
    .Q_N(_5510_),
    .Q(\logix.ram_r[1433] ));
 sg13g2_dfrbp_1 \logix.ram_r[1434]$_DFFE_PP_  (.CLK(net668),
    .RESET_B(net1280),
    .D(_0489_),
    .Q_N(_5509_),
    .Q(\logix.ram_r[1434] ));
 sg13g2_dfrbp_1 \logix.ram_r[1435]$_DFFE_PP_  (.CLK(net659),
    .RESET_B(net1281),
    .D(_0490_),
    .Q_N(_5508_),
    .Q(\logix.ram_r[1435] ));
 sg13g2_dfrbp_1 \logix.ram_r[1436]$_DFFE_PP_  (.CLK(net659),
    .RESET_B(net1282),
    .D(_0491_),
    .Q_N(_5507_),
    .Q(\logix.ram_r[1436] ));
 sg13g2_dfrbp_1 \logix.ram_r[1437]$_DFFE_PP_  (.CLK(net651),
    .RESET_B(net1283),
    .D(_0492_),
    .Q_N(_5506_),
    .Q(\logix.ram_r[1437] ));
 sg13g2_dfrbp_1 \logix.ram_r[1438]$_DFFE_PP_  (.CLK(net645),
    .RESET_B(net1284),
    .D(_0493_),
    .Q_N(_5505_),
    .Q(\logix.ram_r[1438] ));
 sg13g2_dfrbp_1 \logix.ram_r[1439]$_DFFE_PP_  (.CLK(net652),
    .RESET_B(net1285),
    .D(_0494_),
    .Q_N(_5504_),
    .Q(\logix.ram_r[1439] ));
 sg13g2_dfrbp_1 \logix.ram_r[143]$_DFFE_PP_  (.CLK(net574),
    .RESET_B(net1286),
    .D(_0495_),
    .Q_N(_5503_),
    .Q(\logix.ram_r[143] ));
 sg13g2_dfrbp_1 \logix.ram_r[1440]$_DFFE_PP_  (.CLK(net646),
    .RESET_B(net1287),
    .D(_0496_),
    .Q_N(_5502_),
    .Q(\logix.ram_r[1440] ));
 sg13g2_dfrbp_1 \logix.ram_r[1441]$_DFFE_PP_  (.CLK(net584),
    .RESET_B(net1288),
    .D(_0497_),
    .Q_N(_5501_),
    .Q(\logix.ram_r[1441] ));
 sg13g2_dfrbp_1 \logix.ram_r[1442]$_DFFE_PP_  (.CLK(net584),
    .RESET_B(net1289),
    .D(_0498_),
    .Q_N(_5500_),
    .Q(\logix.ram_r[1442] ));
 sg13g2_dfrbp_1 \logix.ram_r[1443]$_DFFE_PP_  (.CLK(net584),
    .RESET_B(net1290),
    .D(_0499_),
    .Q_N(_5499_),
    .Q(\logix.ram_r[1443] ));
 sg13g2_dfrbp_1 \logix.ram_r[1444]$_DFFE_PP_  (.CLK(net577),
    .RESET_B(net1291),
    .D(_0500_),
    .Q_N(_5498_),
    .Q(\logix.ram_r[1444] ));
 sg13g2_dfrbp_1 \logix.ram_r[1445]$_DFFE_PP_  (.CLK(net636),
    .RESET_B(net1292),
    .D(_0501_),
    .Q_N(_5497_),
    .Q(\logix.ram_r[1445] ));
 sg13g2_dfrbp_1 \logix.ram_r[1446]$_DFFE_PP_  (.CLK(net637),
    .RESET_B(net1293),
    .D(_0502_),
    .Q_N(_5496_),
    .Q(\logix.ram_r[1446] ));
 sg13g2_dfrbp_1 \logix.ram_r[1447]$_DFFE_PP_  (.CLK(net645),
    .RESET_B(net1294),
    .D(_0503_),
    .Q_N(_5495_),
    .Q(\logix.ram_r[1447] ));
 sg13g2_dfrbp_1 \logix.ram_r[1448]$_DFFE_PP_  (.CLK(net645),
    .RESET_B(net1295),
    .D(_0504_),
    .Q_N(_5494_),
    .Q(\logix.ram_r[1448] ));
 sg13g2_dfrbp_1 \logix.ram_r[1449]$_DFFE_PP_  (.CLK(net584),
    .RESET_B(net1296),
    .D(_0505_),
    .Q_N(_5493_),
    .Q(\logix.ram_r[1449] ));
 sg13g2_dfrbp_1 \logix.ram_r[144]$_DFFE_PP_  (.CLK(net574),
    .RESET_B(net1297),
    .D(_0506_),
    .Q_N(_5492_),
    .Q(\logix.ram_r[144] ));
 sg13g2_dfrbp_1 \logix.ram_r[1450]$_DFFE_PP_  (.CLK(net585),
    .RESET_B(net1298),
    .D(_0507_),
    .Q_N(_5491_),
    .Q(\logix.ram_r[1450] ));
 sg13g2_dfrbp_1 \logix.ram_r[1451]$_DFFE_PP_  (.CLK(net585),
    .RESET_B(net1299),
    .D(_0508_),
    .Q_N(_5490_),
    .Q(\logix.ram_r[1451] ));
 sg13g2_dfrbp_1 \logix.ram_r[1452]$_DFFE_PP_  (.CLK(net585),
    .RESET_B(net1300),
    .D(_0509_),
    .Q_N(_5489_),
    .Q(\logix.ram_r[1452] ));
 sg13g2_dfrbp_1 \logix.ram_r[1453]$_DFFE_PP_  (.CLK(net645),
    .RESET_B(net1301),
    .D(_0510_),
    .Q_N(_5488_),
    .Q(\logix.ram_r[1453] ));
 sg13g2_dfrbp_1 \logix.ram_r[1454]$_DFFE_PP_  (.CLK(net645),
    .RESET_B(net1302),
    .D(_0511_),
    .Q_N(_5487_),
    .Q(\logix.ram_r[1454] ));
 sg13g2_dfrbp_1 \logix.ram_r[1455]$_DFFE_PP_  (.CLK(net645),
    .RESET_B(net1303),
    .D(_0512_),
    .Q_N(_5486_),
    .Q(\logix.ram_r[1455] ));
 sg13g2_dfrbp_1 \logix.ram_r[1456]$_DFFE_PP_  (.CLK(net645),
    .RESET_B(net1304),
    .D(_0513_),
    .Q_N(_5485_),
    .Q(\logix.ram_r[1456] ));
 sg13g2_dfrbp_1 \logix.ram_r[1457]$_DFFE_PP_  (.CLK(net584),
    .RESET_B(net1305),
    .D(_0514_),
    .Q_N(_5484_),
    .Q(\logix.ram_r[1457] ));
 sg13g2_dfrbp_1 \logix.ram_r[1458]$_DFFE_PP_  (.CLK(net585),
    .RESET_B(net1306),
    .D(_0515_),
    .Q_N(_5483_),
    .Q(\logix.ram_r[1458] ));
 sg13g2_dfrbp_1 \logix.ram_r[1459]$_DFFE_PP_  (.CLK(net585),
    .RESET_B(net1307),
    .D(_0516_),
    .Q_N(_5482_),
    .Q(\logix.ram_r[1459] ));
 sg13g2_dfrbp_1 \logix.ram_r[145]$_DFFE_PP_  (.CLK(net574),
    .RESET_B(net1308),
    .D(_0517_),
    .Q_N(_5481_),
    .Q(\logix.ram_r[145] ));
 sg13g2_dfrbp_1 \logix.ram_r[1460]$_DFFE_PP_  (.CLK(net577),
    .RESET_B(net1309),
    .D(_0518_),
    .Q_N(_5480_),
    .Q(\logix.ram_r[1460] ));
 sg13g2_dfrbp_1 \logix.ram_r[1461]$_DFFE_PP_  (.CLK(net636),
    .RESET_B(net1310),
    .D(_0519_),
    .Q_N(_5479_),
    .Q(\logix.ram_r[1461] ));
 sg13g2_dfrbp_1 \logix.ram_r[1462]$_DFFE_PP_  (.CLK(net646),
    .RESET_B(net1311),
    .D(_0520_),
    .Q_N(_5478_),
    .Q(\logix.ram_r[1462] ));
 sg13g2_dfrbp_1 \logix.ram_r[1463]$_DFFE_PP_  (.CLK(net646),
    .RESET_B(net1312),
    .D(_0521_),
    .Q_N(_5477_),
    .Q(\logix.ram_r[1463] ));
 sg13g2_dfrbp_1 \logix.ram_r[1464]$_DFFE_PP_  (.CLK(net646),
    .RESET_B(net1313),
    .D(_0522_),
    .Q_N(_5476_),
    .Q(\logix.ram_r[1464] ));
 sg13g2_dfrbp_1 \logix.ram_r[1465]$_DFFE_PP_  (.CLK(net646),
    .RESET_B(net1314),
    .D(_0523_),
    .Q_N(_5475_),
    .Q(\logix.ram_r[1465] ));
 sg13g2_dfrbp_1 \logix.ram_r[1466]$_DFFE_PP_  (.CLK(net584),
    .RESET_B(net1315),
    .D(_0524_),
    .Q_N(_5474_),
    .Q(\logix.ram_r[1466] ));
 sg13g2_dfrbp_1 \logix.ram_r[1467]$_DFFE_PP_  (.CLK(net584),
    .RESET_B(net1316),
    .D(_0525_),
    .Q_N(_5473_),
    .Q(\logix.ram_r[1467] ));
 sg13g2_dfrbp_1 \logix.ram_r[1468]$_DFFE_PP_  (.CLK(net584),
    .RESET_B(net1317),
    .D(_0526_),
    .Q_N(_5472_),
    .Q(\logix.ram_r[1468] ));
 sg13g2_dfrbp_1 \logix.ram_r[1469]$_DFFE_PP_  (.CLK(net580),
    .RESET_B(net1318),
    .D(_0527_),
    .Q_N(_5471_),
    .Q(\logix.ram_r[1469] ));
 sg13g2_dfrbp_1 \logix.ram_r[146]$_DFFE_PP_  (.CLK(net540),
    .RESET_B(net1319),
    .D(_0528_),
    .Q_N(_5470_),
    .Q(\logix.ram_r[146] ));
 sg13g2_dfrbp_1 \logix.ram_r[1470]$_DFFE_PP_  (.CLK(net580),
    .RESET_B(net1320),
    .D(_0529_),
    .Q_N(_5469_),
    .Q(\logix.ram_r[1470] ));
 sg13g2_dfrbp_1 \logix.ram_r[1471]$_DFFE_PP_  (.CLK(net581),
    .RESET_B(net1321),
    .D(_0530_),
    .Q_N(_5468_),
    .Q(\logix.ram_r[1471] ));
 sg13g2_dfrbp_1 \logix.ram_r[1472]$_DFFE_PP_  (.CLK(net581),
    .RESET_B(net1322),
    .D(_0531_),
    .Q_N(_5467_),
    .Q(\logix.ram_r[1472] ));
 sg13g2_dfrbp_1 \logix.ram_r[1473]$_DFFE_PP_  (.CLK(net581),
    .RESET_B(net1323),
    .D(_0532_),
    .Q_N(_5466_),
    .Q(\logix.ram_r[1473] ));
 sg13g2_dfrbp_1 \logix.ram_r[1474]$_DFFE_PP_  (.CLK(net581),
    .RESET_B(net1324),
    .D(_0533_),
    .Q_N(_5465_),
    .Q(\logix.ram_r[1474] ));
 sg13g2_dfrbp_1 \logix.ram_r[1475]$_DFFE_PP_  (.CLK(net582),
    .RESET_B(net1325),
    .D(_0534_),
    .Q_N(_5464_),
    .Q(\logix.ram_r[1475] ));
 sg13g2_dfrbp_1 \logix.ram_r[1476]$_DFFE_PP_  (.CLK(net586),
    .RESET_B(net1326),
    .D(_0535_),
    .Q_N(_5463_),
    .Q(\logix.ram_r[1476] ));
 sg13g2_dfrbp_1 \logix.ram_r[1477]$_DFFE_PP_  (.CLK(net586),
    .RESET_B(net1327),
    .D(_0536_),
    .Q_N(_5462_),
    .Q(\logix.ram_r[1477] ));
 sg13g2_dfrbp_1 \logix.ram_r[1478]$_DFFE_PP_  (.CLK(net586),
    .RESET_B(net1328),
    .D(_0537_),
    .Q_N(_5461_),
    .Q(\logix.ram_r[1478] ));
 sg13g2_dfrbp_1 \logix.ram_r[1479]$_DFFE_PP_  (.CLK(net587),
    .RESET_B(net1329),
    .D(_0538_),
    .Q_N(_5460_),
    .Q(\logix.ram_r[1479] ));
 sg13g2_dfrbp_1 \logix.ram_r[147]$_DFFE_PP_  (.CLK(net540),
    .RESET_B(net1330),
    .D(_0539_),
    .Q_N(_5459_),
    .Q(\logix.ram_r[147] ));
 sg13g2_dfrbp_1 \logix.ram_r[1480]$_DFFE_PP_  (.CLK(net586),
    .RESET_B(net1331),
    .D(_0540_),
    .Q_N(_5458_),
    .Q(\logix.ram_r[1480] ));
 sg13g2_dfrbp_1 \logix.ram_r[1481]$_DFFE_PP_  (.CLK(net583),
    .RESET_B(net1332),
    .D(_0541_),
    .Q_N(_5457_),
    .Q(\logix.ram_r[1481] ));
 sg13g2_dfrbp_1 \logix.ram_r[1482]$_DFFE_PP_  (.CLK(net583),
    .RESET_B(net1333),
    .D(_0542_),
    .Q_N(_5456_),
    .Q(\logix.ram_r[1482] ));
 sg13g2_dfrbp_1 \logix.ram_r[1483]$_DFFE_PP_  (.CLK(net582),
    .RESET_B(net1334),
    .D(_0543_),
    .Q_N(_5455_),
    .Q(\logix.ram_r[1483] ));
 sg13g2_dfrbp_1 \logix.ram_r[1484]$_DFFE_PP_  (.CLK(net582),
    .RESET_B(net1335),
    .D(_0544_),
    .Q_N(_5454_),
    .Q(\logix.ram_r[1484] ));
 sg13g2_dfrbp_1 \logix.ram_r[1485]$_DFFE_PP_  (.CLK(net586),
    .RESET_B(net1336),
    .D(_0545_),
    .Q_N(_5453_),
    .Q(\logix.ram_r[1485] ));
 sg13g2_dfrbp_1 \logix.ram_r[1486]$_DFFE_PP_  (.CLK(net587),
    .RESET_B(net1337),
    .D(_0546_),
    .Q_N(_5452_),
    .Q(\logix.ram_r[1486] ));
 sg13g2_dfrbp_1 \logix.ram_r[1487]$_DFFE_PP_  (.CLK(net587),
    .RESET_B(net1338),
    .D(_0547_),
    .Q_N(_5451_),
    .Q(\logix.ram_r[1487] ));
 sg13g2_dfrbp_1 \logix.ram_r[1488]$_DFFE_PP_  (.CLK(net587),
    .RESET_B(net1339),
    .D(_0548_),
    .Q_N(_5450_),
    .Q(\logix.ram_r[1488] ));
 sg13g2_dfrbp_1 \logix.ram_r[1489]$_DFFE_PP_  (.CLK(net581),
    .RESET_B(net1340),
    .D(_0549_),
    .Q_N(_5449_),
    .Q(\logix.ram_r[1489] ));
 sg13g2_dfrbp_1 \logix.ram_r[148]$_DFFE_PP_  (.CLK(net540),
    .RESET_B(net1341),
    .D(_0550_),
    .Q_N(_5448_),
    .Q(\logix.ram_r[148] ));
 sg13g2_dfrbp_1 \logix.ram_r[1490]$_DFFE_PP_  (.CLK(net582),
    .RESET_B(net1342),
    .D(_0551_),
    .Q_N(_5447_),
    .Q(\logix.ram_r[1490] ));
 sg13g2_dfrbp_1 \logix.ram_r[1491]$_DFFE_PP_  (.CLK(net582),
    .RESET_B(net1343),
    .D(_0552_),
    .Q_N(_5446_),
    .Q(\logix.ram_r[1491] ));
 sg13g2_dfrbp_1 \logix.ram_r[1492]$_DFFE_PP_  (.CLK(net586),
    .RESET_B(net1344),
    .D(_0553_),
    .Q_N(_5445_),
    .Q(\logix.ram_r[1492] ));
 sg13g2_dfrbp_1 \logix.ram_r[1493]$_DFFE_PP_  (.CLK(net586),
    .RESET_B(net1345),
    .D(_0554_),
    .Q_N(_5444_),
    .Q(\logix.ram_r[1493] ));
 sg13g2_dfrbp_1 \logix.ram_r[1494]$_DFFE_PP_  (.CLK(net587),
    .RESET_B(net1346),
    .D(_0555_),
    .Q_N(_5443_),
    .Q(\logix.ram_r[1494] ));
 sg13g2_dfrbp_1 \logix.ram_r[1495]$_DFFE_PP_  (.CLK(net587),
    .RESET_B(net1347),
    .D(_0556_),
    .Q_N(_5442_),
    .Q(\logix.ram_r[1495] ));
 sg13g2_dfrbp_1 \logix.ram_r[1496]$_DFFE_PP_  (.CLK(net586),
    .RESET_B(net1348),
    .D(_0557_),
    .Q_N(_5441_),
    .Q(\logix.ram_r[1496] ));
 sg13g2_dfrbp_1 \logix.ram_r[1497]$_DFFE_PP_  (.CLK(net582),
    .RESET_B(net1349),
    .D(_0558_),
    .Q_N(_5440_),
    .Q(\logix.ram_r[1497] ));
 sg13g2_dfrbp_1 \logix.ram_r[1498]$_DFFE_PP_  (.CLK(net582),
    .RESET_B(net1350),
    .D(_0559_),
    .Q_N(_5439_),
    .Q(\logix.ram_r[1498] ));
 sg13g2_dfrbp_1 \logix.ram_r[1499]$_DFFE_PP_  (.CLK(net582),
    .RESET_B(net1351),
    .D(_0560_),
    .Q_N(_5438_),
    .Q(\logix.ram_r[1499] ));
 sg13g2_dfrbp_1 \logix.ram_r[149]$_DFFE_PP_  (.CLK(net541),
    .RESET_B(net1352),
    .D(_0561_),
    .Q_N(_5437_),
    .Q(\logix.ram_r[149] ));
 sg13g2_dfrbp_1 \logix.ram_r[14]$_DFFE_PP_  (.CLK(net604),
    .RESET_B(net1353),
    .D(_0562_),
    .Q_N(_5436_),
    .Q(\logix.ram_r[14] ));
 sg13g2_dfrbp_1 \logix.ram_r[1500]$_DFFE_PP_  (.CLK(net583),
    .RESET_B(net1354),
    .D(_0563_),
    .Q_N(_5435_),
    .Q(\logix.ram_r[1500] ));
 sg13g2_dfrbp_1 \logix.ram_r[1501]$_DFFE_PP_  (.CLK(net587),
    .RESET_B(net1355),
    .D(_0564_),
    .Q_N(_5434_),
    .Q(\logix.ram_r[1501] ));
 sg13g2_dfrbp_1 \logix.ram_r[1502]$_DFFE_PP_  (.CLK(net588),
    .RESET_B(net1356),
    .D(_0565_),
    .Q_N(_5433_),
    .Q(\logix.ram_r[1502] ));
 sg13g2_dfrbp_1 \logix.ram_r[1503]$_DFFE_PP_  (.CLK(net588),
    .RESET_B(net1357),
    .D(_0566_),
    .Q_N(_5432_),
    .Q(\logix.ram_r[1503] ));
 sg13g2_dfrbp_1 \logix.ram_r[1504]$_DFFE_PP_  (.CLK(net647),
    .RESET_B(net1358),
    .D(_0567_),
    .Q_N(_5431_),
    .Q(\logix.ram_r[1504] ));
 sg13g2_dfrbp_1 \logix.ram_r[1505]$_DFFE_PP_  (.CLK(net648),
    .RESET_B(net1359),
    .D(_0568_),
    .Q_N(_5430_),
    .Q(\logix.ram_r[1505] ));
 sg13g2_dfrbp_1 \logix.ram_r[1506]$_DFFE_PP_  (.CLK(net648),
    .RESET_B(net1360),
    .D(_0569_),
    .Q_N(_5429_),
    .Q(\logix.ram_r[1506] ));
 sg13g2_dfrbp_1 \logix.ram_r[1507]$_DFFE_PP_  (.CLK(net648),
    .RESET_B(net1361),
    .D(_0570_),
    .Q_N(_5428_),
    .Q(\logix.ram_r[1507] ));
 sg13g2_dfrbp_1 \logix.ram_r[1508]$_DFFE_PP_  (.CLK(net647),
    .RESET_B(net1362),
    .D(_0571_),
    .Q_N(_5427_),
    .Q(\logix.ram_r[1508] ));
 sg13g2_dfrbp_1 \logix.ram_r[1509]$_DFFE_PP_  (.CLK(net647),
    .RESET_B(net1363),
    .D(_0572_),
    .Q_N(_5426_),
    .Q(\logix.ram_r[1509] ));
 sg13g2_dfrbp_1 \logix.ram_r[150]$_DFFE_PP_  (.CLK(net541),
    .RESET_B(net1364),
    .D(_0573_),
    .Q_N(_5425_),
    .Q(\logix.ram_r[150] ));
 sg13g2_dfrbp_1 \logix.ram_r[1510]$_DFFE_PP_  (.CLK(net647),
    .RESET_B(net1365),
    .D(_0574_),
    .Q_N(_5424_),
    .Q(\logix.ram_r[1510] ));
 sg13g2_dfrbp_1 \logix.ram_r[1511]$_DFFE_PP_  (.CLK(net648),
    .RESET_B(net1366),
    .D(_0575_),
    .Q_N(_5423_),
    .Q(\logix.ram_r[1511] ));
 sg13g2_dfrbp_1 \logix.ram_r[1512]$_DFFE_PP_  (.CLK(net649),
    .RESET_B(net1367),
    .D(_0576_),
    .Q_N(_5422_),
    .Q(\logix.ram_r[1512] ));
 sg13g2_dfrbp_1 \logix.ram_r[1513]$_DFFE_PP_  (.CLK(net653),
    .RESET_B(net1368),
    .D(_0577_),
    .Q_N(_5421_),
    .Q(\logix.ram_r[1513] ));
 sg13g2_dfrbp_1 \logix.ram_r[1514]$_DFFE_PP_  (.CLK(net653),
    .RESET_B(net1369),
    .D(_0578_),
    .Q_N(_5420_),
    .Q(\logix.ram_r[1514] ));
 sg13g2_dfrbp_1 \logix.ram_r[1515]$_DFFE_PP_  (.CLK(net653),
    .RESET_B(net1370),
    .D(_0579_),
    .Q_N(_5419_),
    .Q(\logix.ram_r[1515] ));
 sg13g2_dfrbp_1 \logix.ram_r[1516]$_DFFE_PP_  (.CLK(net653),
    .RESET_B(net1371),
    .D(_0580_),
    .Q_N(_5418_),
    .Q(\logix.ram_r[1516] ));
 sg13g2_dfrbp_1 \logix.ram_r[1517]$_DFFE_PP_  (.CLK(net648),
    .RESET_B(net1372),
    .D(_0581_),
    .Q_N(_5417_),
    .Q(\logix.ram_r[1517] ));
 sg13g2_dfrbp_1 \logix.ram_r[1518]$_DFFE_PP_  (.CLK(net647),
    .RESET_B(net1373),
    .D(_0582_),
    .Q_N(_5416_),
    .Q(\logix.ram_r[1518] ));
 sg13g2_dfrbp_1 \logix.ram_r[1519]$_DFFE_PP_  (.CLK(net646),
    .RESET_B(net1374),
    .D(_0583_),
    .Q_N(_5415_),
    .Q(\logix.ram_r[1519] ));
 sg13g2_dfrbp_1 \logix.ram_r[151]$_DFFE_PP_  (.CLK(net545),
    .RESET_B(net1375),
    .D(_0584_),
    .Q_N(_5414_),
    .Q(\logix.ram_r[151] ));
 sg13g2_dfrbp_1 \logix.ram_r[1520]$_DFFE_PP_  (.CLK(net652),
    .RESET_B(net1376),
    .D(_0585_),
    .Q_N(_5413_),
    .Q(\logix.ram_r[1520] ));
 sg13g2_dfrbp_1 \logix.ram_r[1521]$_DFFE_PP_  (.CLK(net653),
    .RESET_B(net1377),
    .D(_0586_),
    .Q_N(_5412_),
    .Q(\logix.ram_r[1521] ));
 sg13g2_dfrbp_1 \logix.ram_r[1522]$_DFFE_PP_  (.CLK(net653),
    .RESET_B(net1378),
    .D(_0587_),
    .Q_N(_5411_),
    .Q(\logix.ram_r[1522] ));
 sg13g2_dfrbp_1 \logix.ram_r[1523]$_DFFE_PP_  (.CLK(net655),
    .RESET_B(net1379),
    .D(_0588_),
    .Q_N(_5410_),
    .Q(\logix.ram_r[1523] ));
 sg13g2_dfrbp_1 \logix.ram_r[1524]$_DFFE_PP_  (.CLK(net649),
    .RESET_B(net1380),
    .D(_0589_),
    .Q_N(_5409_),
    .Q(\logix.ram_r[1524] ));
 sg13g2_dfrbp_1 \logix.ram_r[1525]$_DFFE_PP_  (.CLK(net648),
    .RESET_B(net1381),
    .D(_0590_),
    .Q_N(_5408_),
    .Q(\logix.ram_r[1525] ));
 sg13g2_dfrbp_1 \logix.ram_r[1526]$_DFFE_PP_  (.CLK(net647),
    .RESET_B(net1382),
    .D(_0591_),
    .Q_N(_5407_),
    .Q(\logix.ram_r[1526] ));
 sg13g2_dfrbp_1 \logix.ram_r[1527]$_DFFE_PP_  (.CLK(net649),
    .RESET_B(net1383),
    .D(_0592_),
    .Q_N(_5406_),
    .Q(\logix.ram_r[1527] ));
 sg13g2_dfrbp_1 \logix.ram_r[1528]$_DFFE_PP_  (.CLK(net652),
    .RESET_B(net1384),
    .D(_0593_),
    .Q_N(_5405_),
    .Q(\logix.ram_r[1528] ));
 sg13g2_dfrbp_1 \logix.ram_r[1529]$_DFFE_PP_  (.CLK(net653),
    .RESET_B(net1385),
    .D(_0594_),
    .Q_N(_5404_),
    .Q(\logix.ram_r[1529] ));
 sg13g2_dfrbp_1 \logix.ram_r[152]$_DFFE_PP_  (.CLK(net545),
    .RESET_B(net1386),
    .D(_0595_),
    .Q_N(_5403_),
    .Q(\logix.ram_r[152] ));
 sg13g2_dfrbp_1 \logix.ram_r[1530]$_DFFE_PP_  (.CLK(net653),
    .RESET_B(net1387),
    .D(_0596_),
    .Q_N(_5402_),
    .Q(\logix.ram_r[1530] ));
 sg13g2_dfrbp_1 \logix.ram_r[1531]$_DFFE_PP_  (.CLK(net649),
    .RESET_B(net1388),
    .D(_0597_),
    .Q_N(_5401_),
    .Q(\logix.ram_r[1531] ));
 sg13g2_dfrbp_1 \logix.ram_r[1532]$_DFFE_PP_  (.CLK(net648),
    .RESET_B(net1389),
    .D(_0598_),
    .Q_N(_5400_),
    .Q(\logix.ram_r[1532] ));
 sg13g2_dfrbp_1 \logix.ram_r[1533]$_DFFE_PP_  (.CLK(net647),
    .RESET_B(net1390),
    .D(_0599_),
    .Q_N(_5399_),
    .Q(\logix.ram_r[1533] ));
 sg13g2_dfrbp_1 \logix.ram_r[1534]$_DFFE_PP_  (.CLK(net647),
    .RESET_B(net1391),
    .D(_0600_),
    .Q_N(_5398_),
    .Q(\logix.ram_r[1534] ));
 sg13g2_dfrbp_1 \logix.ram_r[1535]$_DFFE_PP_  (.CLK(net645),
    .RESET_B(net1392),
    .D(_0601_),
    .Q_N(_5397_),
    .Q(\logix.ram_r[1535] ));
 sg13g2_dfrbp_1 \logix.ram_r[1536]$_DFFE_PP_  (.CLK(net534),
    .RESET_B(net1393),
    .D(_0602_),
    .Q_N(_5396_),
    .Q(\logix.ram_r[1536] ));
 sg13g2_dfrbp_1 \logix.ram_r[1537]$_DFFE_PP_  (.CLK(net534),
    .RESET_B(net1394),
    .D(_0603_),
    .Q_N(_5395_),
    .Q(\logix.ram_r[1537] ));
 sg13g2_dfrbp_1 \logix.ram_r[1538]$_DFFE_PP_  (.CLK(net593),
    .RESET_B(net1395),
    .D(_0604_),
    .Q_N(_5394_),
    .Q(\logix.ram_r[1538] ));
 sg13g2_dfrbp_1 \logix.ram_r[1539]$_DFFE_PP_  (.CLK(net593),
    .RESET_B(net1396),
    .D(_0605_),
    .Q_N(_5393_),
    .Q(\logix.ram_r[1539] ));
 sg13g2_dfrbp_1 \logix.ram_r[153]$_DFFE_PP_  (.CLK(net545),
    .RESET_B(net1397),
    .D(_0606_),
    .Q_N(_5392_),
    .Q(\logix.ram_r[153] ));
 sg13g2_dfrbp_1 \logix.ram_r[1540]$_DFFE_PP_  (.CLK(net529),
    .RESET_B(net1398),
    .D(_0607_),
    .Q_N(_5391_),
    .Q(\logix.ram_r[1540] ));
 sg13g2_dfrbp_1 \logix.ram_r[1541]$_DFFE_PP_  (.CLK(net529),
    .RESET_B(net1399),
    .D(_0608_),
    .Q_N(_5390_),
    .Q(\logix.ram_r[1541] ));
 sg13g2_dfrbp_1 \logix.ram_r[1542]$_DFFE_PP_  (.CLK(net529),
    .RESET_B(net1400),
    .D(_0609_),
    .Q_N(_5389_),
    .Q(\logix.ram_r[1542] ));
 sg13g2_dfrbp_1 \logix.ram_r[1543]$_DFFE_PP_  (.CLK(net529),
    .RESET_B(net1401),
    .D(_0610_),
    .Q_N(_5388_),
    .Q(\logix.ram_r[1543] ));
 sg13g2_dfrbp_1 \logix.ram_r[1544]$_DFFE_PP_  (.CLK(net533),
    .RESET_B(net1402),
    .D(_0611_),
    .Q_N(_5387_),
    .Q(\logix.ram_r[1544] ));
 sg13g2_dfrbp_1 \logix.ram_r[1545]$_DFFE_PP_  (.CLK(net535),
    .RESET_B(net1403),
    .D(_0612_),
    .Q_N(_5386_),
    .Q(\logix.ram_r[1545] ));
 sg13g2_dfrbp_1 \logix.ram_r[1546]$_DFFE_PP_  (.CLK(net534),
    .RESET_B(net1404),
    .D(_0613_),
    .Q_N(_5385_),
    .Q(\logix.ram_r[1546] ));
 sg13g2_dfrbp_1 \logix.ram_r[1547]$_DFFE_PP_  (.CLK(net534),
    .RESET_B(net1405),
    .D(_0614_),
    .Q_N(_5384_),
    .Q(\logix.ram_r[1547] ));
 sg13g2_dfrbp_1 \logix.ram_r[1548]$_DFFE_PP_  (.CLK(net534),
    .RESET_B(net1406),
    .D(_0615_),
    .Q_N(_5383_),
    .Q(\logix.ram_r[1548] ));
 sg13g2_dfrbp_1 \logix.ram_r[1549]$_DFFE_PP_  (.CLK(net529),
    .RESET_B(net1407),
    .D(_0616_),
    .Q_N(_5382_),
    .Q(\logix.ram_r[1549] ));
 sg13g2_dfrbp_1 \logix.ram_r[154]$_DFFE_PP_  (.CLK(net541),
    .RESET_B(net1408),
    .D(_0617_),
    .Q_N(_5381_),
    .Q(\logix.ram_r[154] ));
 sg13g2_dfrbp_1 \logix.ram_r[1550]$_DFFE_PP_  (.CLK(net532),
    .RESET_B(net1409),
    .D(_0618_),
    .Q_N(_5380_),
    .Q(\logix.ram_r[1550] ));
 sg13g2_dfrbp_1 \logix.ram_r[1551]$_DFFE_PP_  (.CLK(net533),
    .RESET_B(net1410),
    .D(_0619_),
    .Q_N(_5379_),
    .Q(\logix.ram_r[1551] ));
 sg13g2_dfrbp_1 \logix.ram_r[1552]$_DFFE_PP_  (.CLK(net533),
    .RESET_B(net1411),
    .D(_0620_),
    .Q_N(_5378_),
    .Q(\logix.ram_r[1552] ));
 sg13g2_dfrbp_1 \logix.ram_r[1553]$_DFFE_PP_  (.CLK(net535),
    .RESET_B(net1412),
    .D(_0621_),
    .Q_N(_5377_),
    .Q(\logix.ram_r[1553] ));
 sg13g2_dfrbp_1 \logix.ram_r[1554]$_DFFE_PP_  (.CLK(net534),
    .RESET_B(net1413),
    .D(_0622_),
    .Q_N(_5376_),
    .Q(\logix.ram_r[1554] ));
 sg13g2_dfrbp_1 \logix.ram_r[1555]$_DFFE_PP_  (.CLK(net534),
    .RESET_B(net1414),
    .D(_0623_),
    .Q_N(_5375_),
    .Q(\logix.ram_r[1555] ));
 sg13g2_dfrbp_1 \logix.ram_r[1556]$_DFFE_PP_  (.CLK(net533),
    .RESET_B(net1415),
    .D(_0624_),
    .Q_N(_5374_),
    .Q(\logix.ram_r[1556] ));
 sg13g2_dfrbp_1 \logix.ram_r[1557]$_DFFE_PP_  (.CLK(net532),
    .RESET_B(net1416),
    .D(_0625_),
    .Q_N(_5373_),
    .Q(\logix.ram_r[1557] ));
 sg13g2_dfrbp_1 \logix.ram_r[1558]$_DFFE_PP_  (.CLK(net533),
    .RESET_B(net1417),
    .D(_0626_),
    .Q_N(_5372_),
    .Q(\logix.ram_r[1558] ));
 sg13g2_dfrbp_1 \logix.ram_r[1559]$_DFFE_PP_  (.CLK(net533),
    .RESET_B(net1418),
    .D(_0627_),
    .Q_N(_5371_),
    .Q(\logix.ram_r[1559] ));
 sg13g2_dfrbp_1 \logix.ram_r[155]$_DFFE_PP_  (.CLK(net539),
    .RESET_B(net1419),
    .D(_0628_),
    .Q_N(_5370_),
    .Q(\logix.ram_r[155] ));
 sg13g2_dfrbp_1 \logix.ram_r[1560]$_DFFE_PP_  (.CLK(net535),
    .RESET_B(net1420),
    .D(_0629_),
    .Q_N(_5369_),
    .Q(\logix.ram_r[1560] ));
 sg13g2_dfrbp_1 \logix.ram_r[1561]$_DFFE_PP_  (.CLK(net534),
    .RESET_B(net1421),
    .D(_0630_),
    .Q_N(_5368_),
    .Q(\logix.ram_r[1561] ));
 sg13g2_dfrbp_1 \logix.ram_r[1562]$_DFFE_PP_  (.CLK(net593),
    .RESET_B(net1422),
    .D(_0631_),
    .Q_N(_5367_),
    .Q(\logix.ram_r[1562] ));
 sg13g2_dfrbp_1 \logix.ram_r[1563]$_DFFE_PP_  (.CLK(net593),
    .RESET_B(net1423),
    .D(_0632_),
    .Q_N(_5366_),
    .Q(\logix.ram_r[1563] ));
 sg13g2_dfrbp_1 \logix.ram_r[1564]$_DFFE_PP_  (.CLK(net593),
    .RESET_B(net1424),
    .D(_0633_),
    .Q_N(_5365_),
    .Q(\logix.ram_r[1564] ));
 sg13g2_dfrbp_1 \logix.ram_r[1565]$_DFFE_PP_  (.CLK(net532),
    .RESET_B(net1425),
    .D(_0634_),
    .Q_N(_5364_),
    .Q(\logix.ram_r[1565] ));
 sg13g2_dfrbp_1 \logix.ram_r[1566]$_DFFE_PP_  (.CLK(net533),
    .RESET_B(net1426),
    .D(_0635_),
    .Q_N(_5363_),
    .Q(\logix.ram_r[1566] ));
 sg13g2_dfrbp_1 \logix.ram_r[1567]$_DFFE_PP_  (.CLK(net533),
    .RESET_B(net1427),
    .D(_0636_),
    .Q_N(_5362_),
    .Q(\logix.ram_r[1567] ));
 sg13g2_dfrbp_1 \logix.ram_r[1568]$_DFFE_PP_  (.CLK(net535),
    .RESET_B(net1428),
    .D(_0637_),
    .Q_N(_5361_),
    .Q(\logix.ram_r[1568] ));
 sg13g2_dfrbp_1 \logix.ram_r[1569]$_DFFE_PP_  (.CLK(net536),
    .RESET_B(net1429),
    .D(_0638_),
    .Q_N(_5360_),
    .Q(\logix.ram_r[1569] ));
 sg13g2_dfrbp_1 \logix.ram_r[156]$_DFFE_PP_  (.CLK(net539),
    .RESET_B(net1430),
    .D(_0639_),
    .Q_N(_5359_),
    .Q(\logix.ram_r[156] ));
 sg13g2_dfrbp_1 \logix.ram_r[1570]$_DFFE_PP_  (.CLK(net536),
    .RESET_B(net1431),
    .D(_0640_),
    .Q_N(_5358_),
    .Q(\logix.ram_r[1570] ));
 sg13g2_dfrbp_1 \logix.ram_r[1571]$_DFFE_PP_  (.CLK(net530),
    .RESET_B(net1432),
    .D(_0641_),
    .Q_N(_5357_),
    .Q(\logix.ram_r[1571] ));
 sg13g2_dfrbp_1 \logix.ram_r[1572]$_DFFE_PP_  (.CLK(net530),
    .RESET_B(net1433),
    .D(_0642_),
    .Q_N(_5356_),
    .Q(\logix.ram_r[1572] ));
 sg13g2_dfrbp_1 \logix.ram_r[1573]$_DFFE_PP_  (.CLK(net530),
    .RESET_B(net1434),
    .D(_0643_),
    .Q_N(_5355_),
    .Q(\logix.ram_r[1573] ));
 sg13g2_dfrbp_1 \logix.ram_r[1574]$_DFFE_PP_  (.CLK(net538),
    .RESET_B(net1435),
    .D(_0644_),
    .Q_N(_5354_),
    .Q(\logix.ram_r[1574] ));
 sg13g2_dfrbp_1 \logix.ram_r[1575]$_DFFE_PP_  (.CLK(net539),
    .RESET_B(net1436),
    .D(_0645_),
    .Q_N(_5353_),
    .Q(\logix.ram_r[1575] ));
 sg13g2_dfrbp_1 \logix.ram_r[1576]$_DFFE_PP_  (.CLK(net536),
    .RESET_B(net1437),
    .D(_0646_),
    .Q_N(_5352_),
    .Q(\logix.ram_r[1576] ));
 sg13g2_dfrbp_1 \logix.ram_r[1577]$_DFFE_PP_  (.CLK(net536),
    .RESET_B(net1438),
    .D(_0647_),
    .Q_N(_5351_),
    .Q(\logix.ram_r[1577] ));
 sg13g2_dfrbp_1 \logix.ram_r[1578]$_DFFE_PP_  (.CLK(net536),
    .RESET_B(net1439),
    .D(_0648_),
    .Q_N(_5350_),
    .Q(\logix.ram_r[1578] ));
 sg13g2_dfrbp_1 \logix.ram_r[1579]$_DFFE_PP_  (.CLK(net530),
    .RESET_B(net1440),
    .D(_0649_),
    .Q_N(_5349_),
    .Q(\logix.ram_r[1579] ));
 sg13g2_dfrbp_1 \logix.ram_r[157]$_DFFE_PP_  (.CLK(net539),
    .RESET_B(net1441),
    .D(_0650_),
    .Q_N(_5348_),
    .Q(\logix.ram_r[157] ));
 sg13g2_dfrbp_1 \logix.ram_r[1580]$_DFFE_PP_  (.CLK(net530),
    .RESET_B(net1442),
    .D(_0651_),
    .Q_N(_5347_),
    .Q(\logix.ram_r[1580] ));
 sg13g2_dfrbp_1 \logix.ram_r[1581]$_DFFE_PP_  (.CLK(net530),
    .RESET_B(net1443),
    .D(_0652_),
    .Q_N(_5346_),
    .Q(\logix.ram_r[1581] ));
 sg13g2_dfrbp_1 \logix.ram_r[1582]$_DFFE_PP_  (.CLK(net538),
    .RESET_B(net1444),
    .D(_0653_),
    .Q_N(_5345_),
    .Q(\logix.ram_r[1582] ));
 sg13g2_dfrbp_1 \logix.ram_r[1583]$_DFFE_PP_  (.CLK(net542),
    .RESET_B(net1445),
    .D(_0654_),
    .Q_N(_5344_),
    .Q(\logix.ram_r[1583] ));
 sg13g2_dfrbp_1 \logix.ram_r[1584]$_DFFE_PP_  (.CLK(net536),
    .RESET_B(net1446),
    .D(_0655_),
    .Q_N(_5343_),
    .Q(\logix.ram_r[1584] ));
 sg13g2_dfrbp_1 \logix.ram_r[1585]$_DFFE_PP_  (.CLK(net536),
    .RESET_B(net1447),
    .D(_0656_),
    .Q_N(_5342_),
    .Q(\logix.ram_r[1585] ));
 sg13g2_dfrbp_1 \logix.ram_r[1586]$_DFFE_PP_  (.CLK(net536),
    .RESET_B(net1448),
    .D(_0657_),
    .Q_N(_5341_),
    .Q(\logix.ram_r[1586] ));
 sg13g2_dfrbp_1 \logix.ram_r[1587]$_DFFE_PP_  (.CLK(net531),
    .RESET_B(net1449),
    .D(_0658_),
    .Q_N(_5340_),
    .Q(\logix.ram_r[1587] ));
 sg13g2_dfrbp_1 \logix.ram_r[1588]$_DFFE_PP_  (.CLK(net531),
    .RESET_B(net1450),
    .D(_0659_),
    .Q_N(_5339_),
    .Q(\logix.ram_r[1588] ));
 sg13g2_dfrbp_1 \logix.ram_r[1589]$_DFFE_PP_  (.CLK(net531),
    .RESET_B(net1451),
    .D(_0660_),
    .Q_N(_5338_),
    .Q(\logix.ram_r[1589] ));
 sg13g2_dfrbp_1 \logix.ram_r[158]$_DFFE_PP_  (.CLK(net542),
    .RESET_B(net1452),
    .D(_0661_),
    .Q_N(_5337_),
    .Q(\logix.ram_r[158] ));
 sg13g2_dfrbp_1 \logix.ram_r[1590]$_DFFE_PP_  (.CLK(net531),
    .RESET_B(net1453),
    .D(_0662_),
    .Q_N(_5336_),
    .Q(\logix.ram_r[1590] ));
 sg13g2_dfrbp_1 \logix.ram_r[1591]$_DFFE_PP_  (.CLK(net537),
    .RESET_B(net1454),
    .D(_0663_),
    .Q_N(_5335_),
    .Q(\logix.ram_r[1591] ));
 sg13g2_dfrbp_1 \logix.ram_r[1592]$_DFFE_PP_  (.CLK(net537),
    .RESET_B(net1455),
    .D(_0664_),
    .Q_N(_5334_),
    .Q(\logix.ram_r[1592] ));
 sg13g2_dfrbp_1 \logix.ram_r[1593]$_DFFE_PP_  (.CLK(net537),
    .RESET_B(net1456),
    .D(_0665_),
    .Q_N(_5333_),
    .Q(\logix.ram_r[1593] ));
 sg13g2_dfrbp_1 \logix.ram_r[1594]$_DFFE_PP_  (.CLK(net537),
    .RESET_B(net1457),
    .D(_0666_),
    .Q_N(_5332_),
    .Q(\logix.ram_r[1594] ));
 sg13g2_dfrbp_1 \logix.ram_r[1595]$_DFFE_PP_  (.CLK(net531),
    .RESET_B(net1458),
    .D(_0667_),
    .Q_N(_5331_),
    .Q(\logix.ram_r[1595] ));
 sg13g2_dfrbp_1 \logix.ram_r[1596]$_DFFE_PP_  (.CLK(net530),
    .RESET_B(net1459),
    .D(_0668_),
    .Q_N(_5330_),
    .Q(\logix.ram_r[1596] ));
 sg13g2_dfrbp_1 \logix.ram_r[1597]$_DFFE_PP_  (.CLK(net530),
    .RESET_B(net1460),
    .D(_0669_),
    .Q_N(_5329_),
    .Q(\logix.ram_r[1597] ));
 sg13g2_dfrbp_1 \logix.ram_r[1598]$_DFFE_PP_  (.CLK(net538),
    .RESET_B(net1461),
    .D(_0670_),
    .Q_N(_5328_),
    .Q(\logix.ram_r[1598] ));
 sg13g2_dfrbp_1 \logix.ram_r[1599]$_DFFE_PP_  (.CLK(net538),
    .RESET_B(net1462),
    .D(_0671_),
    .Q_N(_5327_),
    .Q(\logix.ram_r[1599] ));
 sg13g2_dfrbp_1 \logix.ram_r[159]$_DFFE_PP_  (.CLK(net543),
    .RESET_B(net1463),
    .D(_0672_),
    .Q_N(_5326_),
    .Q(\logix.ram_r[159] ));
 sg13g2_dfrbp_1 \logix.ram_r[15]$_DFFE_PP_  (.CLK(net604),
    .RESET_B(net1464),
    .D(_0673_),
    .Q_N(_5325_),
    .Q(\logix.ram_r[15] ));
 sg13g2_dfrbp_1 \logix.ram_r[1600]$_DFFE_PP_  (.CLK(net538),
    .RESET_B(net1465),
    .D(_0674_),
    .Q_N(_5324_),
    .Q(\logix.ram_r[1600] ));
 sg13g2_dfrbp_1 \logix.ram_r[1601]$_DFFE_PP_  (.CLK(net523),
    .RESET_B(net1466),
    .D(_0675_),
    .Q_N(_5323_),
    .Q(\logix.ram_r[1601] ));
 sg13g2_dfrbp_1 \logix.ram_r[1602]$_DFFE_PP_  (.CLK(net515),
    .RESET_B(net1467),
    .D(_0676_),
    .Q_N(_5322_),
    .Q(\logix.ram_r[1602] ));
 sg13g2_dfrbp_1 \logix.ram_r[1603]$_DFFE_PP_  (.CLK(net516),
    .RESET_B(net1468),
    .D(_0677_),
    .Q_N(_5321_),
    .Q(\logix.ram_r[1603] ));
 sg13g2_dfrbp_1 \logix.ram_r[1604]$_DFFE_PP_  (.CLK(net515),
    .RESET_B(net1469),
    .D(_0678_),
    .Q_N(_5320_),
    .Q(\logix.ram_r[1604] ));
 sg13g2_dfrbp_1 \logix.ram_r[1605]$_DFFE_PP_  (.CLK(net509),
    .RESET_B(net1470),
    .D(_0679_),
    .Q_N(_5319_),
    .Q(\logix.ram_r[1605] ));
 sg13g2_dfrbp_1 \logix.ram_r[1606]$_DFFE_PP_  (.CLK(net509),
    .RESET_B(net1471),
    .D(_0680_),
    .Q_N(_5318_),
    .Q(\logix.ram_r[1606] ));
 sg13g2_dfrbp_1 \logix.ram_r[1607]$_DFFE_PP_  (.CLK(net519),
    .RESET_B(net1472),
    .D(_0681_),
    .Q_N(_5317_),
    .Q(\logix.ram_r[1607] ));
 sg13g2_dfrbp_1 \logix.ram_r[1608]$_DFFE_PP_  (.CLK(net523),
    .RESET_B(net1473),
    .D(_0682_),
    .Q_N(_5316_),
    .Q(\logix.ram_r[1608] ));
 sg13g2_dfrbp_1 \logix.ram_r[1609]$_DFFE_PP_  (.CLK(net523),
    .RESET_B(net1474),
    .D(_0683_),
    .Q_N(_5315_),
    .Q(\logix.ram_r[1609] ));
 sg13g2_dfrbp_1 \logix.ram_r[160]$_DFFE_PP_  (.CLK(net519),
    .RESET_B(net1475),
    .D(_0684_),
    .Q_N(_5314_),
    .Q(\logix.ram_r[160] ));
 sg13g2_dfrbp_1 \logix.ram_r[1610]$_DFFE_PP_  (.CLK(net515),
    .RESET_B(net1476),
    .D(_0685_),
    .Q_N(_5313_),
    .Q(\logix.ram_r[1610] ));
 sg13g2_dfrbp_1 \logix.ram_r[1611]$_DFFE_PP_  (.CLK(net516),
    .RESET_B(net1477),
    .D(_0686_),
    .Q_N(_5312_),
    .Q(\logix.ram_r[1611] ));
 sg13g2_dfrbp_1 \logix.ram_r[1612]$_DFFE_PP_  (.CLK(net515),
    .RESET_B(net1478),
    .D(_0687_),
    .Q_N(_5311_),
    .Q(\logix.ram_r[1612] ));
 sg13g2_dfrbp_1 \logix.ram_r[1613]$_DFFE_PP_  (.CLK(net509),
    .RESET_B(net1479),
    .D(_0688_),
    .Q_N(_5310_),
    .Q(\logix.ram_r[1613] ));
 sg13g2_dfrbp_1 \logix.ram_r[1614]$_DFFE_PP_  (.CLK(net509),
    .RESET_B(net1480),
    .D(_0689_),
    .Q_N(_5309_),
    .Q(\logix.ram_r[1614] ));
 sg13g2_dfrbp_1 \logix.ram_r[1615]$_DFFE_PP_  (.CLK(net511),
    .RESET_B(net1481),
    .D(_0690_),
    .Q_N(_5308_),
    .Q(\logix.ram_r[1615] ));
 sg13g2_dfrbp_1 \logix.ram_r[1616]$_DFFE_PP_  (.CLK(net523),
    .RESET_B(net1482),
    .D(_0691_),
    .Q_N(_5307_),
    .Q(\logix.ram_r[1616] ));
 sg13g2_dfrbp_1 \logix.ram_r[1617]$_DFFE_PP_  (.CLK(net523),
    .RESET_B(net1483),
    .D(_0692_),
    .Q_N(_5306_),
    .Q(\logix.ram_r[1617] ));
 sg13g2_dfrbp_1 \logix.ram_r[1618]$_DFFE_PP_  (.CLK(net515),
    .RESET_B(net1484),
    .D(_0693_),
    .Q_N(_5305_),
    .Q(\logix.ram_r[1618] ));
 sg13g2_dfrbp_1 \logix.ram_r[1619]$_DFFE_PP_  (.CLK(net515),
    .RESET_B(net1485),
    .D(_0694_),
    .Q_N(_5304_),
    .Q(\logix.ram_r[1619] ));
 sg13g2_dfrbp_1 \logix.ram_r[161]$_DFFE_PP_  (.CLK(net519),
    .RESET_B(net1486),
    .D(_0695_),
    .Q_N(_5303_),
    .Q(\logix.ram_r[161] ));
 sg13g2_dfrbp_1 \logix.ram_r[1620]$_DFFE_PP_  (.CLK(net515),
    .RESET_B(net1487),
    .D(_0696_),
    .Q_N(_5302_),
    .Q(\logix.ram_r[1620] ));
 sg13g2_dfrbp_1 \logix.ram_r[1621]$_DFFE_PP_  (.CLK(net509),
    .RESET_B(net1488),
    .D(_0697_),
    .Q_N(_5301_),
    .Q(\logix.ram_r[1621] ));
 sg13g2_dfrbp_1 \logix.ram_r[1622]$_DFFE_PP_  (.CLK(net511),
    .RESET_B(net1489),
    .D(_0698_),
    .Q_N(_5300_),
    .Q(\logix.ram_r[1622] ));
 sg13g2_dfrbp_1 \logix.ram_r[1623]$_DFFE_PP_  (.CLK(net515),
    .RESET_B(net1490),
    .D(_0699_),
    .Q_N(_5299_),
    .Q(\logix.ram_r[1623] ));
 sg13g2_dfrbp_1 \logix.ram_r[1624]$_DFFE_PP_  (.CLK(net523),
    .RESET_B(net1491),
    .D(_0700_),
    .Q_N(_5298_),
    .Q(\logix.ram_r[1624] ));
 sg13g2_dfrbp_1 \logix.ram_r[1625]$_DFFE_PP_  (.CLK(net524),
    .RESET_B(net1492),
    .D(_0701_),
    .Q_N(_5297_),
    .Q(\logix.ram_r[1625] ));
 sg13g2_dfrbp_1 \logix.ram_r[1626]$_DFFE_PP_  (.CLK(net516),
    .RESET_B(net1493),
    .D(_0702_),
    .Q_N(_5296_),
    .Q(\logix.ram_r[1626] ));
 sg13g2_dfrbp_1 \logix.ram_r[1627]$_DFFE_PP_  (.CLK(net516),
    .RESET_B(net1494),
    .D(_0703_),
    .Q_N(_5295_),
    .Q(\logix.ram_r[1627] ));
 sg13g2_dfrbp_1 \logix.ram_r[1628]$_DFFE_PP_  (.CLK(net516),
    .RESET_B(net1495),
    .D(_0704_),
    .Q_N(_5294_),
    .Q(\logix.ram_r[1628] ));
 sg13g2_dfrbp_1 \logix.ram_r[1629]$_DFFE_PP_  (.CLK(net509),
    .RESET_B(net1496),
    .D(_0705_),
    .Q_N(_5293_),
    .Q(\logix.ram_r[1629] ));
 sg13g2_dfrbp_1 \logix.ram_r[162]$_DFFE_PP_  (.CLK(net518),
    .RESET_B(net1497),
    .D(_0706_),
    .Q_N(_5292_),
    .Q(\logix.ram_r[162] ));
 sg13g2_dfrbp_1 \logix.ram_r[1630]$_DFFE_PP_  (.CLK(net510),
    .RESET_B(net1498),
    .D(_0707_),
    .Q_N(_5291_),
    .Q(\logix.ram_r[1630] ));
 sg13g2_dfrbp_1 \logix.ram_r[1631]$_DFFE_PP_  (.CLK(net510),
    .RESET_B(net1499),
    .D(_0708_),
    .Q_N(_5290_),
    .Q(\logix.ram_r[1631] ));
 sg13g2_dfrbp_1 \logix.ram_r[1632]$_DFFE_PP_  (.CLK(net510),
    .RESET_B(net1500),
    .D(_0709_),
    .Q_N(_5289_),
    .Q(\logix.ram_r[1632] ));
 sg13g2_dfrbp_1 \logix.ram_r[1633]$_DFFE_PP_  (.CLK(net449),
    .RESET_B(net1501),
    .D(_0710_),
    .Q_N(_5288_),
    .Q(\logix.ram_r[1633] ));
 sg13g2_dfrbp_1 \logix.ram_r[1634]$_DFFE_PP_  (.CLK(net449),
    .RESET_B(net1502),
    .D(_0711_),
    .Q_N(_5287_),
    .Q(\logix.ram_r[1634] ));
 sg13g2_dfrbp_1 \logix.ram_r[1635]$_DFFE_PP_  (.CLK(net442),
    .RESET_B(net1503),
    .D(_0712_),
    .Q_N(_5286_),
    .Q(\logix.ram_r[1635] ));
 sg13g2_dfrbp_1 \logix.ram_r[1636]$_DFFE_PP_  (.CLK(net442),
    .RESET_B(net1504),
    .D(_0713_),
    .Q_N(_5285_),
    .Q(\logix.ram_r[1636] ));
 sg13g2_dfrbp_1 \logix.ram_r[1637]$_DFFE_PP_  (.CLK(net442),
    .RESET_B(net1505),
    .D(_0714_),
    .Q_N(_5284_),
    .Q(\logix.ram_r[1637] ));
 sg13g2_dfrbp_1 \logix.ram_r[1638]$_DFFE_PP_  (.CLK(net442),
    .RESET_B(net1506),
    .D(_0715_),
    .Q_N(_5283_),
    .Q(\logix.ram_r[1638] ));
 sg13g2_dfrbp_1 \logix.ram_r[1639]$_DFFE_PP_  (.CLK(net442),
    .RESET_B(net1507),
    .D(_0716_),
    .Q_N(_5282_),
    .Q(\logix.ram_r[1639] ));
 sg13g2_dfrbp_1 \logix.ram_r[163]$_DFFE_PP_  (.CLK(net518),
    .RESET_B(net1508),
    .D(_0717_),
    .Q_N(_5281_),
    .Q(\logix.ram_r[163] ));
 sg13g2_dfrbp_1 \logix.ram_r[1640]$_DFFE_PP_  (.CLK(net456),
    .RESET_B(net1509),
    .D(_0718_),
    .Q_N(_5280_),
    .Q(\logix.ram_r[1640] ));
 sg13g2_dfrbp_1 \logix.ram_r[1641]$_DFFE_PP_  (.CLK(net457),
    .RESET_B(net1510),
    .D(_0719_),
    .Q_N(_5279_),
    .Q(\logix.ram_r[1641] ));
 sg13g2_dfrbp_1 \logix.ram_r[1642]$_DFFE_PP_  (.CLK(net449),
    .RESET_B(net1511),
    .D(_0720_),
    .Q_N(_5278_),
    .Q(\logix.ram_r[1642] ));
 sg13g2_dfrbp_1 \logix.ram_r[1643]$_DFFE_PP_  (.CLK(net448),
    .RESET_B(net1512),
    .D(_0721_),
    .Q_N(_5277_),
    .Q(\logix.ram_r[1643] ));
 sg13g2_dfrbp_1 \logix.ram_r[1644]$_DFFE_PP_  (.CLK(net448),
    .RESET_B(net1513),
    .D(_0722_),
    .Q_N(_5276_),
    .Q(\logix.ram_r[1644] ));
 sg13g2_dfrbp_1 \logix.ram_r[1645]$_DFFE_PP_  (.CLK(net444),
    .RESET_B(net1514),
    .D(_0723_),
    .Q_N(_5275_),
    .Q(\logix.ram_r[1645] ));
 sg13g2_dfrbp_1 \logix.ram_r[1646]$_DFFE_PP_  (.CLK(net444),
    .RESET_B(net1515),
    .D(_0724_),
    .Q_N(_5274_),
    .Q(\logix.ram_r[1646] ));
 sg13g2_dfrbp_1 \logix.ram_r[1647]$_DFFE_PP_  (.CLK(net456),
    .RESET_B(net1516),
    .D(_0725_),
    .Q_N(_5273_),
    .Q(\logix.ram_r[1647] ));
 sg13g2_dfrbp_1 \logix.ram_r[1648]$_DFFE_PP_  (.CLK(net457),
    .RESET_B(net1517),
    .D(_0726_),
    .Q_N(_5272_),
    .Q(\logix.ram_r[1648] ));
 sg13g2_dfrbp_1 \logix.ram_r[1649]$_DFFE_PP_  (.CLK(net457),
    .RESET_B(net1518),
    .D(_0727_),
    .Q_N(_5271_),
    .Q(\logix.ram_r[1649] ));
 sg13g2_dfrbp_1 \logix.ram_r[164]$_DFFE_PP_  (.CLK(net518),
    .RESET_B(net1519),
    .D(_0728_),
    .Q_N(_5270_),
    .Q(\logix.ram_r[164] ));
 sg13g2_dfrbp_1 \logix.ram_r[1650]$_DFFE_PP_  (.CLK(net449),
    .RESET_B(net1520),
    .D(_0729_),
    .Q_N(_5269_),
    .Q(\logix.ram_r[1650] ));
 sg13g2_dfrbp_1 \logix.ram_r[1651]$_DFFE_PP_  (.CLK(net448),
    .RESET_B(net1521),
    .D(_0730_),
    .Q_N(_5268_),
    .Q(\logix.ram_r[1651] ));
 sg13g2_dfrbp_1 \logix.ram_r[1652]$_DFFE_PP_  (.CLK(net448),
    .RESET_B(net1522),
    .D(_0731_),
    .Q_N(_5267_),
    .Q(\logix.ram_r[1652] ));
 sg13g2_dfrbp_1 \logix.ram_r[1653]$_DFFE_PP_  (.CLK(net442),
    .RESET_B(net1523),
    .D(_0732_),
    .Q_N(_5266_),
    .Q(\logix.ram_r[1653] ));
 sg13g2_dfrbp_1 \logix.ram_r[1654]$_DFFE_PP_  (.CLK(net444),
    .RESET_B(net1524),
    .D(_0733_),
    .Q_N(_5265_),
    .Q(\logix.ram_r[1654] ));
 sg13g2_dfrbp_1 \logix.ram_r[1655]$_DFFE_PP_  (.CLK(net448),
    .RESET_B(net1525),
    .D(_0734_),
    .Q_N(_5264_),
    .Q(\logix.ram_r[1655] ));
 sg13g2_dfrbp_1 \logix.ram_r[1656]$_DFFE_PP_  (.CLK(net456),
    .RESET_B(net1526),
    .D(_0735_),
    .Q_N(_5263_),
    .Q(\logix.ram_r[1656] ));
 sg13g2_dfrbp_1 \logix.ram_r[1657]$_DFFE_PP_  (.CLK(net449),
    .RESET_B(net1527),
    .D(_0736_),
    .Q_N(_5262_),
    .Q(\logix.ram_r[1657] ));
 sg13g2_dfrbp_1 \logix.ram_r[1658]$_DFFE_PP_  (.CLK(net449),
    .RESET_B(net1528),
    .D(_0737_),
    .Q_N(_5261_),
    .Q(\logix.ram_r[1658] ));
 sg13g2_dfrbp_1 \logix.ram_r[1659]$_DFFE_PP_  (.CLK(net449),
    .RESET_B(net1529),
    .D(_0738_),
    .Q_N(_5260_),
    .Q(\logix.ram_r[1659] ));
 sg13g2_dfrbp_1 \logix.ram_r[165]$_DFFE_PP_  (.CLK(net510),
    .RESET_B(net1530),
    .D(_0739_),
    .Q_N(_5259_),
    .Q(\logix.ram_r[165] ));
 sg13g2_dfrbp_1 \logix.ram_r[1660]$_DFFE_PP_  (.CLK(net448),
    .RESET_B(net1531),
    .D(_0740_),
    .Q_N(_5258_),
    .Q(\logix.ram_r[1660] ));
 sg13g2_dfrbp_1 \logix.ram_r[1661]$_DFFE_PP_  (.CLK(net448),
    .RESET_B(net1532),
    .D(_0741_),
    .Q_N(_5257_),
    .Q(\logix.ram_r[1661] ));
 sg13g2_dfrbp_1 \logix.ram_r[1662]$_DFFE_PP_  (.CLK(net448),
    .RESET_B(net1533),
    .D(_0742_),
    .Q_N(_5256_),
    .Q(\logix.ram_r[1662] ));
 sg13g2_dfrbp_1 \logix.ram_r[1663]$_DFFE_PP_  (.CLK(net445),
    .RESET_B(net1534),
    .D(_0743_),
    .Q_N(_5255_),
    .Q(\logix.ram_r[1663] ));
 sg13g2_dfrbp_1 \logix.ram_r[1664]$_DFFE_PP_  (.CLK(net508),
    .RESET_B(net1535),
    .D(_0744_),
    .Q_N(_5254_),
    .Q(\logix.ram_r[1664] ));
 sg13g2_dfrbp_1 \logix.ram_r[1665]$_DFFE_PP_  (.CLK(net512),
    .RESET_B(net1536),
    .D(_0745_),
    .Q_N(_5253_),
    .Q(\logix.ram_r[1665] ));
 sg13g2_dfrbp_1 \logix.ram_r[1666]$_DFFE_PP_  (.CLK(net512),
    .RESET_B(net1537),
    .D(_0746_),
    .Q_N(_5252_),
    .Q(\logix.ram_r[1666] ));
 sg13g2_dfrbp_1 \logix.ram_r[1667]$_DFFE_PP_  (.CLK(net513),
    .RESET_B(net1538),
    .D(_0747_),
    .Q_N(_5251_),
    .Q(\logix.ram_r[1667] ));
 sg13g2_dfrbp_1 \logix.ram_r[1668]$_DFFE_PP_  (.CLK(net513),
    .RESET_B(net1539),
    .D(_0748_),
    .Q_N(_5250_),
    .Q(\logix.ram_r[1668] ));
 sg13g2_dfrbp_1 \logix.ram_r[1669]$_DFFE_PP_  (.CLK(net513),
    .RESET_B(net1540),
    .D(_0749_),
    .Q_N(_5249_),
    .Q(\logix.ram_r[1669] ));
 sg13g2_dfrbp_1 \logix.ram_r[166]$_DFFE_PP_  (.CLK(net510),
    .RESET_B(net1541),
    .D(_0750_),
    .Q_N(_5248_),
    .Q(\logix.ram_r[166] ));
 sg13g2_dfrbp_1 \logix.ram_r[1670]$_DFFE_PP_  (.CLK(net513),
    .RESET_B(net1542),
    .D(_0751_),
    .Q_N(_5247_),
    .Q(\logix.ram_r[1670] ));
 sg13g2_dfrbp_1 \logix.ram_r[1671]$_DFFE_PP_  (.CLK(net513),
    .RESET_B(net1543),
    .D(_0752_),
    .Q_N(_5246_),
    .Q(\logix.ram_r[1671] ));
 sg13g2_dfrbp_1 \logix.ram_r[1672]$_DFFE_PP_  (.CLK(net508),
    .RESET_B(net1544),
    .D(_0753_),
    .Q_N(_5245_),
    .Q(\logix.ram_r[1672] ));
 sg13g2_dfrbp_1 \logix.ram_r[1673]$_DFFE_PP_  (.CLK(net512),
    .RESET_B(net1545),
    .D(_0754_),
    .Q_N(_5244_),
    .Q(\logix.ram_r[1673] ));
 sg13g2_dfrbp_1 \logix.ram_r[1674]$_DFFE_PP_  (.CLK(net514),
    .RESET_B(net1546),
    .D(_0755_),
    .Q_N(_5243_),
    .Q(\logix.ram_r[1674] ));
 sg13g2_dfrbp_1 \logix.ram_r[1675]$_DFFE_PP_  (.CLK(net513),
    .RESET_B(net1547),
    .D(_0756_),
    .Q_N(_5242_),
    .Q(\logix.ram_r[1675] ));
 sg13g2_dfrbp_1 \logix.ram_r[1676]$_DFFE_PP_  (.CLK(net528),
    .RESET_B(net1548),
    .D(_0757_),
    .Q_N(_5241_),
    .Q(\logix.ram_r[1676] ));
 sg13g2_dfrbp_1 \logix.ram_r[1677]$_DFFE_PP_  (.CLK(net528),
    .RESET_B(net1549),
    .D(_0758_),
    .Q_N(_5240_),
    .Q(\logix.ram_r[1677] ));
 sg13g2_dfrbp_1 \logix.ram_r[1678]$_DFFE_PP_  (.CLK(net528),
    .RESET_B(net1550),
    .D(_0759_),
    .Q_N(_5239_),
    .Q(\logix.ram_r[1678] ));
 sg13g2_dfrbp_1 \logix.ram_r[1679]$_DFFE_PP_  (.CLK(net513),
    .RESET_B(net1551),
    .D(_0760_),
    .Q_N(_5238_),
    .Q(\logix.ram_r[1679] ));
 sg13g2_dfrbp_1 \logix.ram_r[167]$_DFFE_PP_  (.CLK(net510),
    .RESET_B(net1552),
    .D(_0761_),
    .Q_N(_5237_),
    .Q(\logix.ram_r[167] ));
 sg13g2_dfrbp_1 \logix.ram_r[1680]$_DFFE_PP_  (.CLK(net508),
    .RESET_B(net1553),
    .D(_0762_),
    .Q_N(_5236_),
    .Q(\logix.ram_r[1680] ));
 sg13g2_dfrbp_1 \logix.ram_r[1681]$_DFFE_PP_  (.CLK(net512),
    .RESET_B(net1554),
    .D(_0763_),
    .Q_N(_5235_),
    .Q(\logix.ram_r[1681] ));
 sg13g2_dfrbp_1 \logix.ram_r[1682]$_DFFE_PP_  (.CLK(net514),
    .RESET_B(net1555),
    .D(_0764_),
    .Q_N(_5234_),
    .Q(\logix.ram_r[1682] ));
 sg13g2_dfrbp_1 \logix.ram_r[1683]$_DFFE_PP_  (.CLK(net514),
    .RESET_B(net1556),
    .D(_0765_),
    .Q_N(_5233_),
    .Q(\logix.ram_r[1683] ));
 sg13g2_dfrbp_1 \logix.ram_r[1684]$_DFFE_PP_  (.CLK(net528),
    .RESET_B(net1557),
    .D(_0766_),
    .Q_N(_5232_),
    .Q(\logix.ram_r[1684] ));
 sg13g2_dfrbp_1 \logix.ram_r[1685]$_DFFE_PP_  (.CLK(net528),
    .RESET_B(net1558),
    .D(_0767_),
    .Q_N(_5231_),
    .Q(\logix.ram_r[1685] ));
 sg13g2_dfrbp_1 \logix.ram_r[1686]$_DFFE_PP_  (.CLK(net528),
    .RESET_B(net1559),
    .D(_0768_),
    .Q_N(_5230_),
    .Q(\logix.ram_r[1686] ));
 sg13g2_dfrbp_1 \logix.ram_r[1687]$_DFFE_PP_  (.CLK(net512),
    .RESET_B(net1560),
    .D(_0769_),
    .Q_N(_5229_),
    .Q(\logix.ram_r[1687] ));
 sg13g2_dfrbp_1 \logix.ram_r[1688]$_DFFE_PP_  (.CLK(net512),
    .RESET_B(net1561),
    .D(_0770_),
    .Q_N(_5228_),
    .Q(\logix.ram_r[1688] ));
 sg13g2_dfrbp_1 \logix.ram_r[1689]$_DFFE_PP_  (.CLK(net512),
    .RESET_B(net1562),
    .D(_0771_),
    .Q_N(_5227_),
    .Q(\logix.ram_r[1689] ));
 sg13g2_dfrbp_1 \logix.ram_r[168]$_DFFE_PP_  (.CLK(net509),
    .RESET_B(net1563),
    .D(_0772_),
    .Q_N(_5226_),
    .Q(\logix.ram_r[168] ));
 sg13g2_dfrbp_1 \logix.ram_r[1690]$_DFFE_PP_  (.CLK(net513),
    .RESET_B(net1564),
    .D(_0773_),
    .Q_N(_5225_),
    .Q(\logix.ram_r[1690] ));
 sg13g2_dfrbp_1 \logix.ram_r[1691]$_DFFE_PP_  (.CLK(net529),
    .RESET_B(net1565),
    .D(_0774_),
    .Q_N(_5224_),
    .Q(\logix.ram_r[1691] ));
 sg13g2_dfrbp_1 \logix.ram_r[1692]$_DFFE_PP_  (.CLK(net529),
    .RESET_B(net1566),
    .D(_0775_),
    .Q_N(_5223_),
    .Q(\logix.ram_r[1692] ));
 sg13g2_dfrbp_1 \logix.ram_r[1693]$_DFFE_PP_  (.CLK(net528),
    .RESET_B(net1567),
    .D(_0776_),
    .Q_N(_5222_),
    .Q(\logix.ram_r[1693] ));
 sg13g2_dfrbp_1 \logix.ram_r[1694]$_DFFE_PP_  (.CLK(net528),
    .RESET_B(net1568),
    .D(_0777_),
    .Q_N(_5221_),
    .Q(\logix.ram_r[1694] ));
 sg13g2_dfrbp_1 \logix.ram_r[1695]$_DFFE_PP_  (.CLK(net512),
    .RESET_B(net1569),
    .D(_0778_),
    .Q_N(_5220_),
    .Q(\logix.ram_r[1695] ));
 sg13g2_dfrbp_1 \logix.ram_r[1696]$_DFFE_PP_  (.CLK(net508),
    .RESET_B(net1570),
    .D(_0779_),
    .Q_N(_5219_),
    .Q(\logix.ram_r[1696] ));
 sg13g2_dfrbp_1 \logix.ram_r[1697]$_DFFE_PP_  (.CLK(net508),
    .RESET_B(net1571),
    .D(_0780_),
    .Q_N(_5218_),
    .Q(\logix.ram_r[1697] ));
 sg13g2_dfrbp_1 \logix.ram_r[1698]$_DFFE_PP_  (.CLK(net508),
    .RESET_B(net1572),
    .D(_0781_),
    .Q_N(_5217_),
    .Q(\logix.ram_r[1698] ));
 sg13g2_dfrbp_1 \logix.ram_r[1699]$_DFFE_PP_  (.CLK(net445),
    .RESET_B(net1573),
    .D(_0782_),
    .Q_N(_5216_),
    .Q(\logix.ram_r[1699] ));
 sg13g2_dfrbp_1 \logix.ram_r[169]$_DFFE_PP_  (.CLK(net509),
    .RESET_B(net1574),
    .D(_0783_),
    .Q_N(_5215_),
    .Q(\logix.ram_r[169] ));
 sg13g2_dfrbp_1 \logix.ram_r[16]$_DFFE_PP_  (.CLK(net604),
    .RESET_B(net1575),
    .D(_0784_),
    .Q_N(_5214_),
    .Q(\logix.ram_r[16] ));
 sg13g2_dfrbp_1 \logix.ram_r[1700]$_DFFE_PP_  (.CLK(net445),
    .RESET_B(net1576),
    .D(_0785_),
    .Q_N(_5213_),
    .Q(\logix.ram_r[1700] ));
 sg13g2_dfrbp_1 \logix.ram_r[1701]$_DFFE_PP_  (.CLK(net445),
    .RESET_B(net1577),
    .D(_0786_),
    .Q_N(_5212_),
    .Q(\logix.ram_r[1701] ));
 sg13g2_dfrbp_1 \logix.ram_r[1702]$_DFFE_PP_  (.CLK(net446),
    .RESET_B(net1578),
    .D(_0787_),
    .Q_N(_5211_),
    .Q(\logix.ram_r[1702] ));
 sg13g2_dfrbp_1 \logix.ram_r[1703]$_DFFE_PP_  (.CLK(net507),
    .RESET_B(net1579),
    .D(_0788_),
    .Q_N(_5210_),
    .Q(\logix.ram_r[1703] ));
 sg13g2_dfrbp_1 \logix.ram_r[1704]$_DFFE_PP_  (.CLK(net507),
    .RESET_B(net1580),
    .D(_0789_),
    .Q_N(_5209_),
    .Q(\logix.ram_r[1704] ));
 sg13g2_dfrbp_1 \logix.ram_r[1705]$_DFFE_PP_  (.CLK(net507),
    .RESET_B(net1581),
    .D(_0790_),
    .Q_N(_5208_),
    .Q(\logix.ram_r[1705] ));
 sg13g2_dfrbp_1 \logix.ram_r[1706]$_DFFE_PP_  (.CLK(net446),
    .RESET_B(net1582),
    .D(_0791_),
    .Q_N(_5207_),
    .Q(\logix.ram_r[1706] ));
 sg13g2_dfrbp_1 \logix.ram_r[1707]$_DFFE_PP_  (.CLK(net446),
    .RESET_B(net1583),
    .D(_0792_),
    .Q_N(_5206_),
    .Q(\logix.ram_r[1707] ));
 sg13g2_dfrbp_1 \logix.ram_r[1708]$_DFFE_PP_  (.CLK(net445),
    .RESET_B(net1584),
    .D(_0793_),
    .Q_N(_5205_),
    .Q(\logix.ram_r[1708] ));
 sg13g2_dfrbp_1 \logix.ram_r[1709]$_DFFE_PP_  (.CLK(net446),
    .RESET_B(net1585),
    .D(_0794_),
    .Q_N(_5204_),
    .Q(\logix.ram_r[1709] ));
 sg13g2_dfrbp_1 \logix.ram_r[170]$_DFFE_PP_  (.CLK(net510),
    .RESET_B(net1586),
    .D(_0795_),
    .Q_N(_5203_),
    .Q(\logix.ram_r[170] ));
 sg13g2_dfrbp_1 \logix.ram_r[1710]$_DFFE_PP_  (.CLK(net446),
    .RESET_B(net1587),
    .D(_0796_),
    .Q_N(_5202_),
    .Q(\logix.ram_r[1710] ));
 sg13g2_dfrbp_1 \logix.ram_r[1711]$_DFFE_PP_  (.CLK(net507),
    .RESET_B(net1588),
    .D(_0797_),
    .Q_N(_5201_),
    .Q(\logix.ram_r[1711] ));
 sg13g2_dfrbp_1 \logix.ram_r[1712]$_DFFE_PP_  (.CLK(net507),
    .RESET_B(net1589),
    .D(_0798_),
    .Q_N(_5200_),
    .Q(\logix.ram_r[1712] ));
 sg13g2_dfrbp_1 \logix.ram_r[1713]$_DFFE_PP_  (.CLK(net507),
    .RESET_B(net1590),
    .D(_0799_),
    .Q_N(_5199_),
    .Q(\logix.ram_r[1713] ));
 sg13g2_dfrbp_1 \logix.ram_r[1714]$_DFFE_PP_  (.CLK(net507),
    .RESET_B(net1591),
    .D(_0800_),
    .Q_N(_5198_),
    .Q(\logix.ram_r[1714] ));
 sg13g2_dfrbp_1 \logix.ram_r[1715]$_DFFE_PP_  (.CLK(net447),
    .RESET_B(net1592),
    .D(_0801_),
    .Q_N(_5197_),
    .Q(\logix.ram_r[1715] ));
 sg13g2_dfrbp_1 \logix.ram_r[1716]$_DFFE_PP_  (.CLK(net446),
    .RESET_B(net1593),
    .D(_0802_),
    .Q_N(_5196_),
    .Q(\logix.ram_r[1716] ));
 sg13g2_dfrbp_1 \logix.ram_r[1717]$_DFFE_PP_  (.CLK(net446),
    .RESET_B(net1594),
    .D(_0803_),
    .Q_N(_5195_),
    .Q(\logix.ram_r[1717] ));
 sg13g2_dfrbp_1 \logix.ram_r[1718]$_DFFE_PP_  (.CLK(net446),
    .RESET_B(net1595),
    .D(_0804_),
    .Q_N(_5194_),
    .Q(\logix.ram_r[1718] ));
 sg13g2_dfrbp_1 \logix.ram_r[1719]$_DFFE_PP_  (.CLK(net507),
    .RESET_B(net1596),
    .D(_0805_),
    .Q_N(_5193_),
    .Q(\logix.ram_r[1719] ));
 sg13g2_dfrbp_1 \logix.ram_r[171]$_DFFE_PP_  (.CLK(net510),
    .RESET_B(net1597),
    .D(_0806_),
    .Q_N(_5192_),
    .Q(\logix.ram_r[171] ));
 sg13g2_dfrbp_1 \logix.ram_r[1720]$_DFFE_PP_  (.CLK(net511),
    .RESET_B(net1598),
    .D(_0807_),
    .Q_N(_5191_),
    .Q(\logix.ram_r[1720] ));
 sg13g2_dfrbp_1 \logix.ram_r[1721]$_DFFE_PP_  (.CLK(net511),
    .RESET_B(net1599),
    .D(_0808_),
    .Q_N(_5190_),
    .Q(\logix.ram_r[1721] ));
 sg13g2_dfrbp_1 \logix.ram_r[1722]$_DFFE_PP_  (.CLK(net508),
    .RESET_B(net1600),
    .D(_0809_),
    .Q_N(_5189_),
    .Q(\logix.ram_r[1722] ));
 sg13g2_dfrbp_1 \logix.ram_r[1723]$_DFFE_PP_  (.CLK(net447),
    .RESET_B(net1601),
    .D(_0810_),
    .Q_N(_5188_),
    .Q(\logix.ram_r[1723] ));
 sg13g2_dfrbp_1 \logix.ram_r[1724]$_DFFE_PP_  (.CLK(net447),
    .RESET_B(net1602),
    .D(_0811_),
    .Q_N(_5187_),
    .Q(\logix.ram_r[1724] ));
 sg13g2_dfrbp_1 \logix.ram_r[1725]$_DFFE_PP_  (.CLK(net445),
    .RESET_B(net1603),
    .D(_0812_),
    .Q_N(_5186_),
    .Q(\logix.ram_r[1725] ));
 sg13g2_dfrbp_1 \logix.ram_r[1726]$_DFFE_PP_  (.CLK(net445),
    .RESET_B(net1604),
    .D(_0813_),
    .Q_N(_5185_),
    .Q(\logix.ram_r[1726] ));
 sg13g2_dfrbp_1 \logix.ram_r[1727]$_DFFE_PP_  (.CLK(net445),
    .RESET_B(net1605),
    .D(_0814_),
    .Q_N(_5184_),
    .Q(\logix.ram_r[1727] ));
 sg13g2_dfrbp_1 \logix.ram_r[1728]$_DFFE_PP_  (.CLK(net440),
    .RESET_B(net1606),
    .D(_0815_),
    .Q_N(_5183_),
    .Q(\logix.ram_r[1728] ));
 sg13g2_dfrbp_1 \logix.ram_r[1729]$_DFFE_PP_  (.CLK(net440),
    .RESET_B(net1607),
    .D(_0816_),
    .Q_N(_5182_),
    .Q(\logix.ram_r[1729] ));
 sg13g2_dfrbp_1 \logix.ram_r[172]$_DFFE_PP_  (.CLK(net442),
    .RESET_B(net1608),
    .D(_0817_),
    .Q_N(_5181_),
    .Q(\logix.ram_r[172] ));
 sg13g2_dfrbp_1 \logix.ram_r[1730]$_DFFE_PP_  (.CLK(net440),
    .RESET_B(net1609),
    .D(_0818_),
    .Q_N(_5180_),
    .Q(\logix.ram_r[1730] ));
 sg13g2_dfrbp_1 \logix.ram_r[1731]$_DFFE_PP_  (.CLK(net439),
    .RESET_B(net1610),
    .D(_0819_),
    .Q_N(_5179_),
    .Q(\logix.ram_r[1731] ));
 sg13g2_dfrbp_1 \logix.ram_r[1732]$_DFFE_PP_  (.CLK(net421),
    .RESET_B(net1611),
    .D(_0820_),
    .Q_N(_5178_),
    .Q(\logix.ram_r[1732] ));
 sg13g2_dfrbp_1 \logix.ram_r[1733]$_DFFE_PP_  (.CLK(net421),
    .RESET_B(net1612),
    .D(_0821_),
    .Q_N(_5177_),
    .Q(\logix.ram_r[1733] ));
 sg13g2_dfrbp_1 \logix.ram_r[1734]$_DFFE_PP_  (.CLK(net422),
    .RESET_B(net1613),
    .D(_0822_),
    .Q_N(_5176_),
    .Q(\logix.ram_r[1734] ));
 sg13g2_dfrbp_1 \logix.ram_r[1735]$_DFFE_PP_  (.CLK(net439),
    .RESET_B(net1614),
    .D(_0823_),
    .Q_N(_5175_),
    .Q(\logix.ram_r[1735] ));
 sg13g2_dfrbp_1 \logix.ram_r[1736]$_DFFE_PP_  (.CLK(net440),
    .RESET_B(net1615),
    .D(_0824_),
    .Q_N(_5174_),
    .Q(\logix.ram_r[1736] ));
 sg13g2_dfrbp_1 \logix.ram_r[1737]$_DFFE_PP_  (.CLK(net440),
    .RESET_B(net1616),
    .D(_0825_),
    .Q_N(_5173_),
    .Q(\logix.ram_r[1737] ));
 sg13g2_dfrbp_1 \logix.ram_r[1738]$_DFFE_PP_  (.CLK(net440),
    .RESET_B(net1617),
    .D(_0826_),
    .Q_N(_5172_),
    .Q(\logix.ram_r[1738] ));
 sg13g2_dfrbp_1 \logix.ram_r[1739]$_DFFE_PP_  (.CLK(net439),
    .RESET_B(net1618),
    .D(_0827_),
    .Q_N(_5171_),
    .Q(\logix.ram_r[1739] ));
 sg13g2_dfrbp_1 \logix.ram_r[173]$_DFFE_PP_  (.CLK(net443),
    .RESET_B(net1619),
    .D(_0828_),
    .Q_N(_5170_),
    .Q(\logix.ram_r[173] ));
 sg13g2_dfrbp_1 \logix.ram_r[1740]$_DFFE_PP_  (.CLK(net422),
    .RESET_B(net1620),
    .D(_0829_),
    .Q_N(_5169_),
    .Q(\logix.ram_r[1740] ));
 sg13g2_dfrbp_1 \logix.ram_r[1741]$_DFFE_PP_  (.CLK(net422),
    .RESET_B(net1621),
    .D(_0830_),
    .Q_N(_5168_),
    .Q(\logix.ram_r[1741] ));
 sg13g2_dfrbp_1 \logix.ram_r[1742]$_DFFE_PP_  (.CLK(net422),
    .RESET_B(net1622),
    .D(_0831_),
    .Q_N(_5167_),
    .Q(\logix.ram_r[1742] ));
 sg13g2_dfrbp_1 \logix.ram_r[1743]$_DFFE_PP_  (.CLK(net439),
    .RESET_B(net1623),
    .D(_0832_),
    .Q_N(_5166_),
    .Q(\logix.ram_r[1743] ));
 sg13g2_dfrbp_1 \logix.ram_r[1744]$_DFFE_PP_  (.CLK(net439),
    .RESET_B(net1624),
    .D(_0833_),
    .Q_N(_5165_),
    .Q(\logix.ram_r[1744] ));
 sg13g2_dfrbp_1 \logix.ram_r[1745]$_DFFE_PP_  (.CLK(net441),
    .RESET_B(net1625),
    .D(_0834_),
    .Q_N(_5164_),
    .Q(\logix.ram_r[1745] ));
 sg13g2_dfrbp_1 \logix.ram_r[1746]$_DFFE_PP_  (.CLK(net439),
    .RESET_B(net1626),
    .D(_0835_),
    .Q_N(_5163_),
    .Q(\logix.ram_r[1746] ));
 sg13g2_dfrbp_1 \logix.ram_r[1747]$_DFFE_PP_  (.CLK(net439),
    .RESET_B(net1627),
    .D(_0836_),
    .Q_N(_5162_),
    .Q(\logix.ram_r[1747] ));
 sg13g2_dfrbp_1 \logix.ram_r[1748]$_DFFE_PP_  (.CLK(net422),
    .RESET_B(net1628),
    .D(_0837_),
    .Q_N(_5161_),
    .Q(\logix.ram_r[1748] ));
 sg13g2_dfrbp_1 \logix.ram_r[1749]$_DFFE_PP_  (.CLK(net422),
    .RESET_B(net1629),
    .D(_0838_),
    .Q_N(_5160_),
    .Q(\logix.ram_r[1749] ));
 sg13g2_dfrbp_1 \logix.ram_r[174]$_DFFE_PP_  (.CLK(net442),
    .RESET_B(net1630),
    .D(_0839_),
    .Q_N(_5159_),
    .Q(\logix.ram_r[174] ));
 sg13g2_dfrbp_1 \logix.ram_r[1750]$_DFFE_PP_  (.CLK(net422),
    .RESET_B(net1631),
    .D(_0840_),
    .Q_N(_5158_),
    .Q(\logix.ram_r[1750] ));
 sg13g2_dfrbp_1 \logix.ram_r[1751]$_DFFE_PP_  (.CLK(net441),
    .RESET_B(net1632),
    .D(_0841_),
    .Q_N(_5157_),
    .Q(\logix.ram_r[1751] ));
 sg13g2_dfrbp_1 \logix.ram_r[1752]$_DFFE_PP_  (.CLK(net441),
    .RESET_B(net1633),
    .D(_0842_),
    .Q_N(_5156_),
    .Q(\logix.ram_r[1752] ));
 sg13g2_dfrbp_1 \logix.ram_r[1753]$_DFFE_PP_  (.CLK(net440),
    .RESET_B(net1634),
    .D(_0843_),
    .Q_N(_5155_),
    .Q(\logix.ram_r[1753] ));
 sg13g2_dfrbp_1 \logix.ram_r[1754]$_DFFE_PP_  (.CLK(net440),
    .RESET_B(net1635),
    .D(_0844_),
    .Q_N(_5154_),
    .Q(\logix.ram_r[1754] ));
 sg13g2_dfrbp_1 \logix.ram_r[1755]$_DFFE_PP_  (.CLK(net439),
    .RESET_B(net1636),
    .D(_0845_),
    .Q_N(_5153_),
    .Q(\logix.ram_r[1755] ));
 sg13g2_dfrbp_1 \logix.ram_r[1756]$_DFFE_PP_  (.CLK(net422),
    .RESET_B(net1637),
    .D(_0846_),
    .Q_N(_5152_),
    .Q(\logix.ram_r[1756] ));
 sg13g2_dfrbp_1 \logix.ram_r[1757]$_DFFE_PP_  (.CLK(net421),
    .RESET_B(net1638),
    .D(_0847_),
    .Q_N(_5151_),
    .Q(\logix.ram_r[1757] ));
 sg13g2_dfrbp_1 \logix.ram_r[1758]$_DFFE_PP_  (.CLK(net421),
    .RESET_B(net1639),
    .D(_0848_),
    .Q_N(_5150_),
    .Q(\logix.ram_r[1758] ));
 sg13g2_dfrbp_1 \logix.ram_r[1759]$_DFFE_PP_  (.CLK(net421),
    .RESET_B(net1640),
    .D(_0849_),
    .Q_N(_5149_),
    .Q(\logix.ram_r[1759] ));
 sg13g2_dfrbp_1 \logix.ram_r[175]$_DFFE_PP_  (.CLK(net424),
    .RESET_B(net1641),
    .D(_0850_),
    .Q_N(_5148_),
    .Q(\logix.ram_r[175] ));
 sg13g2_dfrbp_1 \logix.ram_r[1760]$_DFFE_PP_  (.CLK(net421),
    .RESET_B(net1642),
    .D(_0851_),
    .Q_N(_5147_),
    .Q(\logix.ram_r[1760] ));
 sg13g2_dfrbp_1 \logix.ram_r[1761]$_DFFE_PP_  (.CLK(net416),
    .RESET_B(net1643),
    .D(_0852_),
    .Q_N(_5146_),
    .Q(\logix.ram_r[1761] ));
 sg13g2_dfrbp_1 \logix.ram_r[1762]$_DFFE_PP_  (.CLK(net414),
    .RESET_B(net1644),
    .D(_0853_),
    .Q_N(_5145_),
    .Q(\logix.ram_r[1762] ));
 sg13g2_dfrbp_1 \logix.ram_r[1763]$_DFFE_PP_  (.CLK(net414),
    .RESET_B(net1645),
    .D(_0854_),
    .Q_N(_5144_),
    .Q(\logix.ram_r[1763] ));
 sg13g2_dfrbp_1 \logix.ram_r[1764]$_DFFE_PP_  (.CLK(net415),
    .RESET_B(net1646),
    .D(_0855_),
    .Q_N(_5143_),
    .Q(\logix.ram_r[1764] ));
 sg13g2_dfrbp_1 \logix.ram_r[1765]$_DFFE_PP_  (.CLK(net415),
    .RESET_B(net1647),
    .D(_0856_),
    .Q_N(_5142_),
    .Q(\logix.ram_r[1765] ));
 sg13g2_dfrbp_1 \logix.ram_r[1766]$_DFFE_PP_  (.CLK(net415),
    .RESET_B(net1648),
    .D(_0857_),
    .Q_N(_5141_),
    .Q(\logix.ram_r[1766] ));
 sg13g2_dfrbp_1 \logix.ram_r[1767]$_DFFE_PP_  (.CLK(net416),
    .RESET_B(net1649),
    .D(_0858_),
    .Q_N(_5140_),
    .Q(\logix.ram_r[1767] ));
 sg13g2_dfrbp_1 \logix.ram_r[1768]$_DFFE_PP_  (.CLK(net416),
    .RESET_B(net1650),
    .D(_0859_),
    .Q_N(_5139_),
    .Q(\logix.ram_r[1768] ));
 sg13g2_dfrbp_1 \logix.ram_r[1769]$_DFFE_PP_  (.CLK(net416),
    .RESET_B(net1651),
    .D(_0860_),
    .Q_N(_5138_),
    .Q(\logix.ram_r[1769] ));
 sg13g2_dfrbp_1 \logix.ram_r[176]$_DFFE_PP_  (.CLK(net424),
    .RESET_B(net1652),
    .D(_0861_),
    .Q_N(_5137_),
    .Q(\logix.ram_r[176] ));
 sg13g2_dfrbp_1 \logix.ram_r[1770]$_DFFE_PP_  (.CLK(net414),
    .RESET_B(net1653),
    .D(_0862_),
    .Q_N(_5136_),
    .Q(\logix.ram_r[1770] ));
 sg13g2_dfrbp_1 \logix.ram_r[1771]$_DFFE_PP_  (.CLK(net414),
    .RESET_B(net1654),
    .D(_0863_),
    .Q_N(_5135_),
    .Q(\logix.ram_r[1771] ));
 sg13g2_dfrbp_1 \logix.ram_r[1772]$_DFFE_PP_  (.CLK(net415),
    .RESET_B(net1655),
    .D(_0864_),
    .Q_N(_5134_),
    .Q(\logix.ram_r[1772] ));
 sg13g2_dfrbp_1 \logix.ram_r[1773]$_DFFE_PP_  (.CLK(net418),
    .RESET_B(net1656),
    .D(_0865_),
    .Q_N(_5133_),
    .Q(\logix.ram_r[1773] ));
 sg13g2_dfrbp_1 \logix.ram_r[1774]$_DFFE_PP_  (.CLK(net420),
    .RESET_B(net1657),
    .D(_0866_),
    .Q_N(_5132_),
    .Q(\logix.ram_r[1774] ));
 sg13g2_dfrbp_1 \logix.ram_r[1775]$_DFFE_PP_  (.CLK(net421),
    .RESET_B(net1658),
    .D(_0867_),
    .Q_N(_5131_),
    .Q(\logix.ram_r[1775] ));
 sg13g2_dfrbp_1 \logix.ram_r[1776]$_DFFE_PP_  (.CLK(net416),
    .RESET_B(net1659),
    .D(_0868_),
    .Q_N(_5130_),
    .Q(\logix.ram_r[1776] ));
 sg13g2_dfrbp_1 \logix.ram_r[1777]$_DFFE_PP_  (.CLK(net416),
    .RESET_B(net1660),
    .D(_0869_),
    .Q_N(_5129_),
    .Q(\logix.ram_r[1777] ));
 sg13g2_dfrbp_1 \logix.ram_r[1778]$_DFFE_PP_  (.CLK(net414),
    .RESET_B(net1661),
    .D(_0870_),
    .Q_N(_5128_),
    .Q(\logix.ram_r[1778] ));
 sg13g2_dfrbp_1 \logix.ram_r[1779]$_DFFE_PP_  (.CLK(net414),
    .RESET_B(net1662),
    .D(_0871_),
    .Q_N(_5127_),
    .Q(\logix.ram_r[1779] ));
 sg13g2_dfrbp_1 \logix.ram_r[177]$_DFFE_PP_  (.CLK(net425),
    .RESET_B(net1663),
    .D(_0872_),
    .Q_N(_5126_),
    .Q(\logix.ram_r[177] ));
 sg13g2_dfrbp_1 \logix.ram_r[1780]$_DFFE_PP_  (.CLK(net415),
    .RESET_B(net1664),
    .D(_0873_),
    .Q_N(_5125_),
    .Q(\logix.ram_r[1780] ));
 sg13g2_dfrbp_1 \logix.ram_r[1781]$_DFFE_PP_  (.CLK(net417),
    .RESET_B(net1665),
    .D(_0874_),
    .Q_N(_5124_),
    .Q(\logix.ram_r[1781] ));
 sg13g2_dfrbp_1 \logix.ram_r[1782]$_DFFE_PP_  (.CLK(net417),
    .RESET_B(net1666),
    .D(_0875_),
    .Q_N(_5123_),
    .Q(\logix.ram_r[1782] ));
 sg13g2_dfrbp_1 \logix.ram_r[1783]$_DFFE_PP_  (.CLK(net421),
    .RESET_B(net1667),
    .D(_0876_),
    .Q_N(_5122_),
    .Q(\logix.ram_r[1783] ));
 sg13g2_dfrbp_1 \logix.ram_r[1784]$_DFFE_PP_  (.CLK(net416),
    .RESET_B(net1668),
    .D(_0877_),
    .Q_N(_5121_),
    .Q(\logix.ram_r[1784] ));
 sg13g2_dfrbp_1 \logix.ram_r[1785]$_DFFE_PP_  (.CLK(net416),
    .RESET_B(net1669),
    .D(_0878_),
    .Q_N(_5120_),
    .Q(\logix.ram_r[1785] ));
 sg13g2_dfrbp_1 \logix.ram_r[1786]$_DFFE_PP_  (.CLK(net414),
    .RESET_B(net1670),
    .D(_0879_),
    .Q_N(_5119_),
    .Q(\logix.ram_r[1786] ));
 sg13g2_dfrbp_1 \logix.ram_r[1787]$_DFFE_PP_  (.CLK(net414),
    .RESET_B(net1671),
    .D(_0880_),
    .Q_N(_5118_),
    .Q(\logix.ram_r[1787] ));
 sg13g2_dfrbp_1 \logix.ram_r[1788]$_DFFE_PP_  (.CLK(net415),
    .RESET_B(net1672),
    .D(_0881_),
    .Q_N(_5117_),
    .Q(\logix.ram_r[1788] ));
 sg13g2_dfrbp_1 \logix.ram_r[1789]$_DFFE_PP_  (.CLK(net418),
    .RESET_B(net1673),
    .D(_0882_),
    .Q_N(_5116_),
    .Q(\logix.ram_r[1789] ));
 sg13g2_dfrbp_1 \logix.ram_r[178]$_DFFE_PP_  (.CLK(net425),
    .RESET_B(net1674),
    .D(_0883_),
    .Q_N(_5115_),
    .Q(\logix.ram_r[178] ));
 sg13g2_dfrbp_1 \logix.ram_r[1790]$_DFFE_PP_  (.CLK(net420),
    .RESET_B(net1675),
    .D(_0884_),
    .Q_N(_5114_),
    .Q(\logix.ram_r[1790] ));
 sg13g2_dfrbp_1 \logix.ram_r[1791]$_DFFE_PP_  (.CLK(net423),
    .RESET_B(net1676),
    .D(_0885_),
    .Q_N(_5113_),
    .Q(\logix.ram_r[1791] ));
 sg13g2_dfrbp_1 \logix.ram_r[1792]$_DFFE_PP_  (.CLK(net423),
    .RESET_B(net1677),
    .D(_0886_),
    .Q_N(_5112_),
    .Q(\logix.ram_r[1792] ));
 sg13g2_dfrbp_1 \logix.ram_r[1793]$_DFFE_PP_  (.CLK(net489),
    .RESET_B(net1678),
    .D(_0887_),
    .Q_N(_5111_),
    .Q(\logix.ram_r[1793] ));
 sg13g2_dfrbp_1 \logix.ram_r[1794]$_DFFE_PP_  (.CLK(net486),
    .RESET_B(net1679),
    .D(_0888_),
    .Q_N(_5110_),
    .Q(\logix.ram_r[1794] ));
 sg13g2_dfrbp_1 \logix.ram_r[1795]$_DFFE_PP_  (.CLK(net487),
    .RESET_B(net1680),
    .D(_0889_),
    .Q_N(_5109_),
    .Q(\logix.ram_r[1795] ));
 sg13g2_dfrbp_1 \logix.ram_r[1796]$_DFFE_PP_  (.CLK(net491),
    .RESET_B(net1681),
    .D(_0890_),
    .Q_N(_5108_),
    .Q(\logix.ram_r[1796] ));
 sg13g2_dfrbp_1 \logix.ram_r[1797]$_DFFE_PP_  (.CLK(net492),
    .RESET_B(net1682),
    .D(_0891_),
    .Q_N(_5107_),
    .Q(\logix.ram_r[1797] ));
 sg13g2_dfrbp_1 \logix.ram_r[1798]$_DFFE_PP_  (.CLK(net489),
    .RESET_B(net1683),
    .D(_0892_),
    .Q_N(_5106_),
    .Q(\logix.ram_r[1798] ));
 sg13g2_dfrbp_1 \logix.ram_r[1799]$_DFFE_PP_  (.CLK(net489),
    .RESET_B(net1684),
    .D(_0893_),
    .Q_N(_5105_),
    .Q(\logix.ram_r[1799] ));
 sg13g2_dfrbp_1 \logix.ram_r[179]$_DFFE_PP_  (.CLK(net550),
    .RESET_B(net1685),
    .D(_0894_),
    .Q_N(_5104_),
    .Q(\logix.ram_r[179] ));
 sg13g2_dfrbp_1 \logix.ram_r[17]$_DFFE_PP_  (.CLK(net640),
    .RESET_B(net1686),
    .D(_0895_),
    .Q_N(_5103_),
    .Q(\logix.ram_r[17] ));
 sg13g2_dfrbp_1 \logix.ram_r[1800]$_DFFE_PP_  (.CLK(net489),
    .RESET_B(net1687),
    .D(_0896_),
    .Q_N(_5102_),
    .Q(\logix.ram_r[1800] ));
 sg13g2_dfrbp_1 \logix.ram_r[1801]$_DFFE_PP_  (.CLK(net489),
    .RESET_B(net1688),
    .D(_0897_),
    .Q_N(_5101_),
    .Q(\logix.ram_r[1801] ));
 sg13g2_dfrbp_1 \logix.ram_r[1802]$_DFFE_PP_  (.CLK(net486),
    .RESET_B(net1689),
    .D(_0898_),
    .Q_N(_5100_),
    .Q(\logix.ram_r[1802] ));
 sg13g2_dfrbp_1 \logix.ram_r[1803]$_DFFE_PP_  (.CLK(net486),
    .RESET_B(net1690),
    .D(_0899_),
    .Q_N(_5099_),
    .Q(\logix.ram_r[1803] ));
 sg13g2_dfrbp_1 \logix.ram_r[1804]$_DFFE_PP_  (.CLK(net491),
    .RESET_B(net1691),
    .D(_0900_),
    .Q_N(_5098_),
    .Q(\logix.ram_r[1804] ));
 sg13g2_dfrbp_1 \logix.ram_r[1805]$_DFFE_PP_  (.CLK(net491),
    .RESET_B(net1692),
    .D(_0901_),
    .Q_N(_5097_),
    .Q(\logix.ram_r[1805] ));
 sg13g2_dfrbp_1 \logix.ram_r[1806]$_DFFE_PP_  (.CLK(net495),
    .RESET_B(net1693),
    .D(_0902_),
    .Q_N(_5096_),
    .Q(\logix.ram_r[1806] ));
 sg13g2_dfrbp_1 \logix.ram_r[1807]$_DFFE_PP_  (.CLK(net496),
    .RESET_B(net1694),
    .D(_0903_),
    .Q_N(_5095_),
    .Q(\logix.ram_r[1807] ));
 sg13g2_dfrbp_1 \logix.ram_r[1808]$_DFFE_PP_  (.CLK(net495),
    .RESET_B(net1695),
    .D(_0904_),
    .Q_N(_5094_),
    .Q(\logix.ram_r[1808] ));
 sg13g2_dfrbp_1 \logix.ram_r[1809]$_DFFE_PP_  (.CLK(net488),
    .RESET_B(net1696),
    .D(_0905_),
    .Q_N(_5093_),
    .Q(\logix.ram_r[1809] ));
 sg13g2_dfrbp_1 \logix.ram_r[180]$_DFFE_PP_  (.CLK(net550),
    .RESET_B(net1697),
    .D(_0906_),
    .Q_N(_5092_),
    .Q(\logix.ram_r[180] ));
 sg13g2_dfrbp_1 \logix.ram_r[1810]$_DFFE_PP_  (.CLK(net488),
    .RESET_B(net1698),
    .D(_0907_),
    .Q_N(_5091_),
    .Q(\logix.ram_r[1810] ));
 sg13g2_dfrbp_1 \logix.ram_r[1811]$_DFFE_PP_  (.CLK(net487),
    .RESET_B(net1699),
    .D(_0908_),
    .Q_N(_5090_),
    .Q(\logix.ram_r[1811] ));
 sg13g2_dfrbp_1 \logix.ram_r[1812]$_DFFE_PP_  (.CLK(net487),
    .RESET_B(net1700),
    .D(_0909_),
    .Q_N(_5089_),
    .Q(\logix.ram_r[1812] ));
 sg13g2_dfrbp_1 \logix.ram_r[1813]$_DFFE_PP_  (.CLK(net488),
    .RESET_B(net1701),
    .D(_0910_),
    .Q_N(_5088_),
    .Q(\logix.ram_r[1813] ));
 sg13g2_dfrbp_1 \logix.ram_r[1814]$_DFFE_PP_  (.CLK(net488),
    .RESET_B(net1702),
    .D(_0911_),
    .Q_N(_5087_),
    .Q(\logix.ram_r[1814] ));
 sg13g2_dfrbp_1 \logix.ram_r[1815]$_DFFE_PP_  (.CLK(net488),
    .RESET_B(net1703),
    .D(_0912_),
    .Q_N(_5086_),
    .Q(\logix.ram_r[1815] ));
 sg13g2_dfrbp_1 \logix.ram_r[1816]$_DFFE_PP_  (.CLK(net488),
    .RESET_B(net1704),
    .D(_0913_),
    .Q_N(_5085_),
    .Q(\logix.ram_r[1816] ));
 sg13g2_dfrbp_1 \logix.ram_r[1817]$_DFFE_PP_  (.CLK(net488),
    .RESET_B(net1705),
    .D(_0914_),
    .Q_N(_5084_),
    .Q(\logix.ram_r[1817] ));
 sg13g2_dfrbp_1 \logix.ram_r[1818]$_DFFE_PP_  (.CLK(net487),
    .RESET_B(net1706),
    .D(_0915_),
    .Q_N(_5083_),
    .Q(\logix.ram_r[1818] ));
 sg13g2_dfrbp_1 \logix.ram_r[1819]$_DFFE_PP_  (.CLK(net487),
    .RESET_B(net1707),
    .D(_0916_),
    .Q_N(_5082_),
    .Q(\logix.ram_r[1819] ));
 sg13g2_dfrbp_1 \logix.ram_r[181]$_DFFE_PP_  (.CLK(net550),
    .RESET_B(net1708),
    .D(_0917_),
    .Q_N(_5081_),
    .Q(\logix.ram_r[181] ));
 sg13g2_dfrbp_1 \logix.ram_r[1820]$_DFFE_PP_  (.CLK(net491),
    .RESET_B(net1709),
    .D(_0918_),
    .Q_N(_5080_),
    .Q(\logix.ram_r[1820] ));
 sg13g2_dfrbp_1 \logix.ram_r[1821]$_DFFE_PP_  (.CLK(net491),
    .RESET_B(net1710),
    .D(_0919_),
    .Q_N(_5079_),
    .Q(\logix.ram_r[1821] ));
 sg13g2_dfrbp_1 \logix.ram_r[1822]$_DFFE_PP_  (.CLK(net488),
    .RESET_B(net1711),
    .D(_0920_),
    .Q_N(_5078_),
    .Q(\logix.ram_r[1822] ));
 sg13g2_dfrbp_1 \logix.ram_r[1823]$_DFFE_PP_  (.CLK(net490),
    .RESET_B(net1712),
    .D(_0921_),
    .Q_N(_5077_),
    .Q(\logix.ram_r[1823] ));
 sg13g2_dfrbp_1 \logix.ram_r[1824]$_DFFE_PP_  (.CLK(net492),
    .RESET_B(net1713),
    .D(_0922_),
    .Q_N(_5076_),
    .Q(\logix.ram_r[1824] ));
 sg13g2_dfrbp_1 \logix.ram_r[1825]$_DFFE_PP_  (.CLK(net492),
    .RESET_B(net1714),
    .D(_0923_),
    .Q_N(_5075_),
    .Q(\logix.ram_r[1825] ));
 sg13g2_dfrbp_1 \logix.ram_r[1826]$_DFFE_PP_  (.CLK(net553),
    .RESET_B(net1715),
    .D(_0924_),
    .Q_N(_5074_),
    .Q(\logix.ram_r[1826] ));
 sg13g2_dfrbp_1 \logix.ram_r[1827]$_DFFE_PP_  (.CLK(net553),
    .RESET_B(net1716),
    .D(_0925_),
    .Q_N(_5073_),
    .Q(\logix.ram_r[1827] ));
 sg13g2_dfrbp_1 \logix.ram_r[1828]$_DFFE_PP_  (.CLK(net553),
    .RESET_B(net1717),
    .D(_0926_),
    .Q_N(_5072_),
    .Q(\logix.ram_r[1828] ));
 sg13g2_dfrbp_1 \logix.ram_r[1829]$_DFFE_PP_  (.CLK(net492),
    .RESET_B(net1718),
    .D(_0927_),
    .Q_N(_5071_),
    .Q(\logix.ram_r[1829] ));
 sg13g2_dfrbp_1 \logix.ram_r[182]$_DFFE_PP_  (.CLK(net550),
    .RESET_B(net1719),
    .D(_0928_),
    .Q_N(_5070_),
    .Q(\logix.ram_r[182] ));
 sg13g2_dfrbp_1 \logix.ram_r[1830]$_DFFE_PP_  (.CLK(net492),
    .RESET_B(net1720),
    .D(_0929_),
    .Q_N(_5069_),
    .Q(\logix.ram_r[1830] ));
 sg13g2_dfrbp_1 \logix.ram_r[1831]$_DFFE_PP_  (.CLK(net492),
    .RESET_B(net1721),
    .D(_0930_),
    .Q_N(_5068_),
    .Q(\logix.ram_r[1831] ));
 sg13g2_dfrbp_1 \logix.ram_r[1832]$_DFFE_PP_  (.CLK(net493),
    .RESET_B(net1722),
    .D(_0931_),
    .Q_N(_5067_),
    .Q(\logix.ram_r[1832] ));
 sg13g2_dfrbp_1 \logix.ram_r[1833]$_DFFE_PP_  (.CLK(net493),
    .RESET_B(net1723),
    .D(_0932_),
    .Q_N(_5066_),
    .Q(\logix.ram_r[1833] ));
 sg13g2_dfrbp_1 \logix.ram_r[1834]$_DFFE_PP_  (.CLK(net553),
    .RESET_B(net1724),
    .D(_0933_),
    .Q_N(_5065_),
    .Q(\logix.ram_r[1834] ));
 sg13g2_dfrbp_1 \logix.ram_r[1835]$_DFFE_PP_  (.CLK(net553),
    .RESET_B(net1725),
    .D(_0934_),
    .Q_N(_5064_),
    .Q(\logix.ram_r[1835] ));
 sg13g2_dfrbp_1 \logix.ram_r[1836]$_DFFE_PP_  (.CLK(net553),
    .RESET_B(net1726),
    .D(_0935_),
    .Q_N(_5063_),
    .Q(\logix.ram_r[1836] ));
 sg13g2_dfrbp_1 \logix.ram_r[1837]$_DFFE_PP_  (.CLK(net501),
    .RESET_B(net1727),
    .D(_0936_),
    .Q_N(_5062_),
    .Q(\logix.ram_r[1837] ));
 sg13g2_dfrbp_1 \logix.ram_r[1838]$_DFFE_PP_  (.CLK(net500),
    .RESET_B(net1728),
    .D(_0937_),
    .Q_N(_5061_),
    .Q(\logix.ram_r[1838] ));
 sg13g2_dfrbp_1 \logix.ram_r[1839]$_DFFE_PP_  (.CLK(net500),
    .RESET_B(net1729),
    .D(_0938_),
    .Q_N(_5060_),
    .Q(\logix.ram_r[1839] ));
 sg13g2_dfrbp_1 \logix.ram_r[183]$_DFFE_PP_  (.CLK(net550),
    .RESET_B(net1730),
    .D(_0939_),
    .Q_N(_5059_),
    .Q(\logix.ram_r[183] ));
 sg13g2_dfrbp_1 \logix.ram_r[1840]$_DFFE_PP_  (.CLK(net492),
    .RESET_B(net1731),
    .D(_0940_),
    .Q_N(_5058_),
    .Q(\logix.ram_r[1840] ));
 sg13g2_dfrbp_1 \logix.ram_r[1841]$_DFFE_PP_  (.CLK(net493),
    .RESET_B(net1732),
    .D(_0941_),
    .Q_N(_5057_),
    .Q(\logix.ram_r[1841] ));
 sg13g2_dfrbp_1 \logix.ram_r[1842]$_DFFE_PP_  (.CLK(net553),
    .RESET_B(net1733),
    .D(_0942_),
    .Q_N(_5056_),
    .Q(\logix.ram_r[1842] ));
 sg13g2_dfrbp_1 \logix.ram_r[1843]$_DFFE_PP_  (.CLK(net559),
    .RESET_B(net1734),
    .D(_0943_),
    .Q_N(_5055_),
    .Q(\logix.ram_r[1843] ));
 sg13g2_dfrbp_1 \logix.ram_r[1844]$_DFFE_PP_  (.CLK(net559),
    .RESET_B(net1735),
    .D(_0944_),
    .Q_N(_5054_),
    .Q(\logix.ram_r[1844] ));
 sg13g2_dfrbp_1 \logix.ram_r[1845]$_DFFE_PP_  (.CLK(net501),
    .RESET_B(net1736),
    .D(_0945_),
    .Q_N(_5053_),
    .Q(\logix.ram_r[1845] ));
 sg13g2_dfrbp_1 \logix.ram_r[1846]$_DFFE_PP_  (.CLK(net500),
    .RESET_B(net1737),
    .D(_0946_),
    .Q_N(_5052_),
    .Q(\logix.ram_r[1846] ));
 sg13g2_dfrbp_1 \logix.ram_r[1847]$_DFFE_PP_  (.CLK(net492),
    .RESET_B(net1738),
    .D(_0947_),
    .Q_N(_5051_),
    .Q(\logix.ram_r[1847] ));
 sg13g2_dfrbp_1 \logix.ram_r[1848]$_DFFE_PP_  (.CLK(net493),
    .RESET_B(net1739),
    .D(_0948_),
    .Q_N(_5050_),
    .Q(\logix.ram_r[1848] ));
 sg13g2_dfrbp_1 \logix.ram_r[1849]$_DFFE_PP_  (.CLK(net493),
    .RESET_B(net1740),
    .D(_0949_),
    .Q_N(_5049_),
    .Q(\logix.ram_r[1849] ));
 sg13g2_dfrbp_1 \logix.ram_r[184]$_DFFE_PP_  (.CLK(net551),
    .RESET_B(net1741),
    .D(_0950_),
    .Q_N(_5048_),
    .Q(\logix.ram_r[184] ));
 sg13g2_dfrbp_1 \logix.ram_r[1850]$_DFFE_PP_  (.CLK(net553),
    .RESET_B(net1742),
    .D(_0951_),
    .Q_N(_5047_),
    .Q(\logix.ram_r[1850] ));
 sg13g2_dfrbp_1 \logix.ram_r[1851]$_DFFE_PP_  (.CLK(net552),
    .RESET_B(net1743),
    .D(_0952_),
    .Q_N(_5046_),
    .Q(\logix.ram_r[1851] ));
 sg13g2_dfrbp_1 \logix.ram_r[1852]$_DFFE_PP_  (.CLK(net552),
    .RESET_B(net1744),
    .D(_0953_),
    .Q_N(_5045_),
    .Q(\logix.ram_r[1852] ));
 sg13g2_dfrbp_1 \logix.ram_r[1853]$_DFFE_PP_  (.CLK(net501),
    .RESET_B(net1745),
    .D(_0954_),
    .Q_N(_5044_),
    .Q(\logix.ram_r[1853] ));
 sg13g2_dfrbp_1 \logix.ram_r[1854]$_DFFE_PP_  (.CLK(net500),
    .RESET_B(net1746),
    .D(_0955_),
    .Q_N(_5043_),
    .Q(\logix.ram_r[1854] ));
 sg13g2_dfrbp_1 \logix.ram_r[1855]$_DFFE_PP_  (.CLK(net501),
    .RESET_B(net1747),
    .D(_0956_),
    .Q_N(_5042_),
    .Q(\logix.ram_r[1855] ));
 sg13g2_dfrbp_1 \logix.ram_r[1856]$_DFFE_PP_  (.CLK(net564),
    .RESET_B(net1748),
    .D(_0957_),
    .Q_N(_5041_),
    .Q(\logix.ram_r[1856] ));
 sg13g2_dfrbp_1 \logix.ram_r[1857]$_DFFE_PP_  (.CLK(net567),
    .RESET_B(net1749),
    .D(_0958_),
    .Q_N(_5040_),
    .Q(\logix.ram_r[1857] ));
 sg13g2_dfrbp_1 \logix.ram_r[1858]$_DFFE_PP_  (.CLK(net566),
    .RESET_B(net1750),
    .D(_0959_),
    .Q_N(_5039_),
    .Q(\logix.ram_r[1858] ));
 sg13g2_dfrbp_1 \logix.ram_r[1859]$_DFFE_PP_  (.CLK(net566),
    .RESET_B(net1751),
    .D(_0960_),
    .Q_N(_5038_),
    .Q(\logix.ram_r[1859] ));
 sg13g2_dfrbp_1 \logix.ram_r[185]$_DFFE_PP_  (.CLK(net552),
    .RESET_B(net1752),
    .D(_0961_),
    .Q_N(_5037_),
    .Q(\logix.ram_r[185] ));
 sg13g2_dfrbp_1 \logix.ram_r[1860]$_DFFE_PP_  (.CLK(net566),
    .RESET_B(net1753),
    .D(_0962_),
    .Q_N(_5036_),
    .Q(\logix.ram_r[1860] ));
 sg13g2_dfrbp_1 \logix.ram_r[1861]$_DFFE_PP_  (.CLK(net560),
    .RESET_B(net1754),
    .D(_0963_),
    .Q_N(_5035_),
    .Q(\logix.ram_r[1861] ));
 sg13g2_dfrbp_1 \logix.ram_r[1862]$_DFFE_PP_  (.CLK(net560),
    .RESET_B(net1755),
    .D(_0964_),
    .Q_N(_5034_),
    .Q(\logix.ram_r[1862] ));
 sg13g2_dfrbp_1 \logix.ram_r[1863]$_DFFE_PP_  (.CLK(net567),
    .RESET_B(net1756),
    .D(_0965_),
    .Q_N(_5033_),
    .Q(\logix.ram_r[1863] ));
 sg13g2_dfrbp_1 \logix.ram_r[1864]$_DFFE_PP_  (.CLK(net567),
    .RESET_B(net1757),
    .D(_0966_),
    .Q_N(_5032_),
    .Q(\logix.ram_r[1864] ));
 sg13g2_dfrbp_1 \logix.ram_r[1865]$_DFFE_PP_  (.CLK(net567),
    .RESET_B(net1758),
    .D(_0967_),
    .Q_N(_5031_),
    .Q(\logix.ram_r[1865] ));
 sg13g2_dfrbp_1 \logix.ram_r[1866]$_DFFE_PP_  (.CLK(net566),
    .RESET_B(net1759),
    .D(_0968_),
    .Q_N(_5030_),
    .Q(\logix.ram_r[1866] ));
 sg13g2_dfrbp_1 \logix.ram_r[1867]$_DFFE_PP_  (.CLK(net583),
    .RESET_B(net1760),
    .D(_0969_),
    .Q_N(_5029_),
    .Q(\logix.ram_r[1867] ));
 sg13g2_dfrbp_1 \logix.ram_r[1868]$_DFFE_PP_  (.CLK(net583),
    .RESET_B(net1761),
    .D(_0970_),
    .Q_N(_5028_),
    .Q(\logix.ram_r[1868] ));
 sg13g2_dfrbp_1 \logix.ram_r[1869]$_DFFE_PP_  (.CLK(net560),
    .RESET_B(net1762),
    .D(_0971_),
    .Q_N(_5027_),
    .Q(\logix.ram_r[1869] ));
 sg13g2_dfrbp_1 \logix.ram_r[186]$_DFFE_PP_  (.CLK(net552),
    .RESET_B(net1763),
    .D(_0972_),
    .Q_N(_5026_),
    .Q(\logix.ram_r[186] ));
 sg13g2_dfrbp_1 \logix.ram_r[1870]$_DFFE_PP_  (.CLK(net560),
    .RESET_B(net1764),
    .D(_0973_),
    .Q_N(_5025_),
    .Q(\logix.ram_r[1870] ));
 sg13g2_dfrbp_1 \logix.ram_r[1871]$_DFFE_PP_  (.CLK(net561),
    .RESET_B(net1765),
    .D(_0974_),
    .Q_N(_5024_),
    .Q(\logix.ram_r[1871] ));
 sg13g2_dfrbp_1 \logix.ram_r[1872]$_DFFE_PP_  (.CLK(net567),
    .RESET_B(net1766),
    .D(_0975_),
    .Q_N(_5023_),
    .Q(\logix.ram_r[1872] ));
 sg13g2_dfrbp_1 \logix.ram_r[1873]$_DFFE_PP_  (.CLK(net566),
    .RESET_B(net1767),
    .D(_0976_),
    .Q_N(_5022_),
    .Q(\logix.ram_r[1873] ));
 sg13g2_dfrbp_1 \logix.ram_r[1874]$_DFFE_PP_  (.CLK(net566),
    .RESET_B(net1768),
    .D(_0977_),
    .Q_N(_5021_),
    .Q(\logix.ram_r[1874] ));
 sg13g2_dfrbp_1 \logix.ram_r[1875]$_DFFE_PP_  (.CLK(net566),
    .RESET_B(net1769),
    .D(_0978_),
    .Q_N(_5020_),
    .Q(\logix.ram_r[1875] ));
 sg13g2_dfrbp_1 \logix.ram_r[1876]$_DFFE_PP_  (.CLK(net566),
    .RESET_B(net1770),
    .D(_0979_),
    .Q_N(_5019_),
    .Q(\logix.ram_r[1876] ));
 sg13g2_dfrbp_1 \logix.ram_r[1877]$_DFFE_PP_  (.CLK(net561),
    .RESET_B(net1771),
    .D(_0980_),
    .Q_N(_5018_),
    .Q(\logix.ram_r[1877] ));
 sg13g2_dfrbp_1 \logix.ram_r[1878]$_DFFE_PP_  (.CLK(net561),
    .RESET_B(net1772),
    .D(_0981_),
    .Q_N(_5017_),
    .Q(\logix.ram_r[1878] ));
 sg13g2_dfrbp_1 \logix.ram_r[1879]$_DFFE_PP_  (.CLK(net561),
    .RESET_B(net1773),
    .D(_0982_),
    .Q_N(_5016_),
    .Q(\logix.ram_r[1879] ));
 sg13g2_dfrbp_1 \logix.ram_r[187]$_DFFE_PP_  (.CLK(net552),
    .RESET_B(net1774),
    .D(_0983_),
    .Q_N(_5015_),
    .Q(\logix.ram_r[187] ));
 sg13g2_dfrbp_1 \logix.ram_r[1880]$_DFFE_PP_  (.CLK(net567),
    .RESET_B(net1775),
    .D(_0984_),
    .Q_N(_5014_),
    .Q(\logix.ram_r[1880] ));
 sg13g2_dfrbp_1 \logix.ram_r[1881]$_DFFE_PP_  (.CLK(net568),
    .RESET_B(net1776),
    .D(_0985_),
    .Q_N(_5013_),
    .Q(\logix.ram_r[1881] ));
 sg13g2_dfrbp_1 \logix.ram_r[1882]$_DFFE_PP_  (.CLK(net568),
    .RESET_B(net1777),
    .D(_0986_),
    .Q_N(_5012_),
    .Q(\logix.ram_r[1882] ));
 sg13g2_dfrbp_1 \logix.ram_r[1883]$_DFFE_PP_  (.CLK(net583),
    .RESET_B(net1778),
    .D(_0987_),
    .Q_N(_5011_),
    .Q(\logix.ram_r[1883] ));
 sg13g2_dfrbp_1 \logix.ram_r[1884]$_DFFE_PP_  (.CLK(net583),
    .RESET_B(net1779),
    .D(_0988_),
    .Q_N(_5010_),
    .Q(\logix.ram_r[1884] ));
 sg13g2_dfrbp_1 \logix.ram_r[1885]$_DFFE_PP_  (.CLK(net562),
    .RESET_B(net1780),
    .D(_0989_),
    .Q_N(_5009_),
    .Q(\logix.ram_r[1885] ));
 sg13g2_dfrbp_1 \logix.ram_r[1886]$_DFFE_PP_  (.CLK(net562),
    .RESET_B(net1781),
    .D(_0990_),
    .Q_N(_5008_),
    .Q(\logix.ram_r[1886] ));
 sg13g2_dfrbp_1 \logix.ram_r[1887]$_DFFE_PP_  (.CLK(net562),
    .RESET_B(net1782),
    .D(_0991_),
    .Q_N(_5007_),
    .Q(\logix.ram_r[1887] ));
 sg13g2_dfrbp_1 \logix.ram_r[1888]$_DFFE_PP_  (.CLK(net562),
    .RESET_B(net1783),
    .D(_0992_),
    .Q_N(_5006_),
    .Q(\logix.ram_r[1888] ));
 sg13g2_dfrbp_1 \logix.ram_r[1889]$_DFFE_PP_  (.CLK(net562),
    .RESET_B(net1784),
    .D(_0993_),
    .Q_N(_5005_),
    .Q(\logix.ram_r[1889] ));
 sg13g2_dfrbp_1 \logix.ram_r[188]$_DFFE_PP_  (.CLK(net552),
    .RESET_B(net1785),
    .D(_0994_),
    .Q_N(_5004_),
    .Q(\logix.ram_r[188] ));
 sg13g2_dfrbp_1 \logix.ram_r[1890]$_DFFE_PP_  (.CLK(net562),
    .RESET_B(net1786),
    .D(_0995_),
    .Q_N(_5003_),
    .Q(\logix.ram_r[1890] ));
 sg13g2_dfrbp_1 \logix.ram_r[1891]$_DFFE_PP_  (.CLK(net560),
    .RESET_B(net1787),
    .D(_0996_),
    .Q_N(_5002_),
    .Q(\logix.ram_r[1891] ));
 sg13g2_dfrbp_1 \logix.ram_r[1892]$_DFFE_PP_  (.CLK(net559),
    .RESET_B(net1788),
    .D(_0997_),
    .Q_N(_5001_),
    .Q(\logix.ram_r[1892] ));
 sg13g2_dfrbp_1 \logix.ram_r[1893]$_DFFE_PP_  (.CLK(net564),
    .RESET_B(net1789),
    .D(_0998_),
    .Q_N(_5000_),
    .Q(\logix.ram_r[1893] ));
 sg13g2_dfrbp_1 \logix.ram_r[1894]$_DFFE_PP_  (.CLK(net564),
    .RESET_B(net1790),
    .D(_0999_),
    .Q_N(_4999_),
    .Q(\logix.ram_r[1894] ));
 sg13g2_dfrbp_1 \logix.ram_r[1895]$_DFFE_PP_  (.CLK(net565),
    .RESET_B(net1791),
    .D(_1000_),
    .Q_N(_4998_),
    .Q(\logix.ram_r[1895] ));
 sg13g2_dfrbp_1 \logix.ram_r[1896]$_DFFE_PP_  (.CLK(net580),
    .RESET_B(net1792),
    .D(_1001_),
    .Q_N(_4997_),
    .Q(\logix.ram_r[1896] ));
 sg13g2_dfrbp_1 \logix.ram_r[1897]$_DFFE_PP_  (.CLK(net580),
    .RESET_B(net1793),
    .D(_1002_),
    .Q_N(_4996_),
    .Q(\logix.ram_r[1897] ));
 sg13g2_dfrbp_1 \logix.ram_r[1898]$_DFFE_PP_  (.CLK(net559),
    .RESET_B(net1794),
    .D(_1003_),
    .Q_N(_4995_),
    .Q(\logix.ram_r[1898] ));
 sg13g2_dfrbp_1 \logix.ram_r[1899]$_DFFE_PP_  (.CLK(net559),
    .RESET_B(net1795),
    .D(_1004_),
    .Q_N(_4994_),
    .Q(\logix.ram_r[1899] ));
 sg13g2_dfrbp_1 \logix.ram_r[189]$_DFFE_PP_  (.CLK(net521),
    .RESET_B(net1796),
    .D(_1005_),
    .Q_N(_4993_),
    .Q(\logix.ram_r[189] ));
 sg13g2_dfrbp_1 \logix.ram_r[18]$_DFFE_PP_  (.CLK(net657),
    .RESET_B(net1797),
    .D(_1006_),
    .Q_N(_4992_),
    .Q(\logix.ram_r[18] ));
 sg13g2_dfrbp_1 \logix.ram_r[1900]$_DFFE_PP_  (.CLK(net559),
    .RESET_B(net1798),
    .D(_1007_),
    .Q_N(_4991_),
    .Q(\logix.ram_r[1900] ));
 sg13g2_dfrbp_1 \logix.ram_r[1901]$_DFFE_PP_  (.CLK(net559),
    .RESET_B(net1799),
    .D(_1008_),
    .Q_N(_4990_),
    .Q(\logix.ram_r[1901] ));
 sg13g2_dfrbp_1 \logix.ram_r[1902]$_DFFE_PP_  (.CLK(net564),
    .RESET_B(net1800),
    .D(_1009_),
    .Q_N(_4989_),
    .Q(\logix.ram_r[1902] ));
 sg13g2_dfrbp_1 \logix.ram_r[1903]$_DFFE_PP_  (.CLK(net564),
    .RESET_B(net1801),
    .D(_1010_),
    .Q_N(_4988_),
    .Q(\logix.ram_r[1903] ));
 sg13g2_dfrbp_1 \logix.ram_r[1904]$_DFFE_PP_  (.CLK(net567),
    .RESET_B(net1802),
    .D(_1011_),
    .Q_N(_4987_),
    .Q(\logix.ram_r[1904] ));
 sg13g2_dfrbp_1 \logix.ram_r[1905]$_DFFE_PP_  (.CLK(net562),
    .RESET_B(net1803),
    .D(_1012_),
    .Q_N(_4986_),
    .Q(\logix.ram_r[1905] ));
 sg13g2_dfrbp_1 \logix.ram_r[1906]$_DFFE_PP_  (.CLK(net560),
    .RESET_B(net1804),
    .D(_1013_),
    .Q_N(_4985_),
    .Q(\logix.ram_r[1906] ));
 sg13g2_dfrbp_1 \logix.ram_r[1907]$_DFFE_PP_  (.CLK(net560),
    .RESET_B(net1805),
    .D(_1014_),
    .Q_N(_4984_),
    .Q(\logix.ram_r[1907] ));
 sg13g2_dfrbp_1 \logix.ram_r[1908]$_DFFE_PP_  (.CLK(net559),
    .RESET_B(net1806),
    .D(_1015_),
    .Q_N(_4983_),
    .Q(\logix.ram_r[1908] ));
 sg13g2_dfrbp_1 \logix.ram_r[1909]$_DFFE_PP_  (.CLK(net564),
    .RESET_B(net1807),
    .D(_1016_),
    .Q_N(_4982_),
    .Q(\logix.ram_r[1909] ));
 sg13g2_dfrbp_1 \logix.ram_r[190]$_DFFE_PP_  (.CLK(net520),
    .RESET_B(net1808),
    .D(_1017_),
    .Q_N(_4981_),
    .Q(\logix.ram_r[190] ));
 sg13g2_dfrbp_1 \logix.ram_r[1910]$_DFFE_PP_  (.CLK(net564),
    .RESET_B(net1809),
    .D(_1018_),
    .Q_N(_4980_),
    .Q(\logix.ram_r[1910] ));
 sg13g2_dfrbp_1 \logix.ram_r[1911]$_DFFE_PP_  (.CLK(net565),
    .RESET_B(net1810),
    .D(_1019_),
    .Q_N(_4979_),
    .Q(\logix.ram_r[1911] ));
 sg13g2_dfrbp_1 \logix.ram_r[1912]$_DFFE_PP_  (.CLK(net564),
    .RESET_B(net1811),
    .D(_1020_),
    .Q_N(_4978_),
    .Q(\logix.ram_r[1912] ));
 sg13g2_dfrbp_1 \logix.ram_r[1913]$_DFFE_PP_  (.CLK(net565),
    .RESET_B(net1812),
    .D(_1021_),
    .Q_N(_4977_),
    .Q(\logix.ram_r[1913] ));
 sg13g2_dfrbp_1 \logix.ram_r[1914]$_DFFE_PP_  (.CLK(net567),
    .RESET_B(net1813),
    .D(_1022_),
    .Q_N(_4976_),
    .Q(\logix.ram_r[1914] ));
 sg13g2_dfrbp_1 \logix.ram_r[1915]$_DFFE_PP_  (.CLK(net560),
    .RESET_B(net1814),
    .D(_1023_),
    .Q_N(_4975_),
    .Q(\logix.ram_r[1915] ));
 sg13g2_dfrbp_1 \logix.ram_r[1916]$_DFFE_PP_  (.CLK(net563),
    .RESET_B(net1815),
    .D(_1024_),
    .Q_N(_4974_),
    .Q(\logix.ram_r[1916] ));
 sg13g2_dfrbp_1 \logix.ram_r[1917]$_DFFE_PP_  (.CLK(net552),
    .RESET_B(net1816),
    .D(_1025_),
    .Q_N(_4973_),
    .Q(\logix.ram_r[1917] ));
 sg13g2_dfrbp_1 \logix.ram_r[1918]$_DFFE_PP_  (.CLK(net557),
    .RESET_B(net1817),
    .D(_1026_),
    .Q_N(_4972_),
    .Q(\logix.ram_r[1918] ));
 sg13g2_dfrbp_1 \logix.ram_r[1919]$_DFFE_PP_  (.CLK(net552),
    .RESET_B(net1818),
    .D(_1027_),
    .Q_N(_4971_),
    .Q(\logix.ram_r[1919] ));
 sg13g2_dfrbp_1 \logix.ram_r[191]$_DFFE_PP_  (.CLK(net520),
    .RESET_B(net1819),
    .D(_1028_),
    .Q_N(_4970_),
    .Q(\logix.ram_r[191] ));
 sg13g2_dfrbp_1 \logix.ram_r[1920]$_DFFE_PP_  (.CLK(net487),
    .RESET_B(net1820),
    .D(_1029_),
    .Q_N(_4969_),
    .Q(\logix.ram_r[1920] ));
 sg13g2_dfrbp_1 \logix.ram_r[1921]$_DFFE_PP_  (.CLK(net453),
    .RESET_B(net1821),
    .D(_1030_),
    .Q_N(_4968_),
    .Q(\logix.ram_r[1921] ));
 sg13g2_dfrbp_1 \logix.ram_r[1922]$_DFFE_PP_  (.CLK(net429),
    .RESET_B(net1822),
    .D(_1031_),
    .Q_N(_4967_),
    .Q(\logix.ram_r[1922] ));
 sg13g2_dfrbp_1 \logix.ram_r[1923]$_DFFE_PP_  (.CLK(net429),
    .RESET_B(net1823),
    .D(_1032_),
    .Q_N(_4966_),
    .Q(\logix.ram_r[1923] ));
 sg13g2_dfrbp_1 \logix.ram_r[1924]$_DFFE_PP_  (.CLK(net426),
    .RESET_B(net1824),
    .D(_1033_),
    .Q_N(_4965_),
    .Q(\logix.ram_r[1924] ));
 sg13g2_dfrbp_1 \logix.ram_r[1925]$_DFFE_PP_  (.CLK(net427),
    .RESET_B(net1825),
    .D(_1034_),
    .Q_N(_4964_),
    .Q(\logix.ram_r[1925] ));
 sg13g2_dfrbp_1 \logix.ram_r[1926]$_DFFE_PP_  (.CLK(net433),
    .RESET_B(net1826),
    .D(_1035_),
    .Q_N(_4963_),
    .Q(\logix.ram_r[1926] ));
 sg13g2_dfrbp_1 \logix.ram_r[1927]$_DFFE_PP_  (.CLK(net433),
    .RESET_B(net1827),
    .D(_1036_),
    .Q_N(_4962_),
    .Q(\logix.ram_r[1927] ));
 sg13g2_dfrbp_1 \logix.ram_r[1928]$_DFFE_PP_  (.CLK(net436),
    .RESET_B(net1828),
    .D(_1037_),
    .Q_N(_4961_),
    .Q(\logix.ram_r[1928] ));
 sg13g2_dfrbp_1 \logix.ram_r[1929]$_DFFE_PP_  (.CLK(net453),
    .RESET_B(net1829),
    .D(_1038_),
    .Q_N(_4960_),
    .Q(\logix.ram_r[1929] ));
 sg13g2_dfrbp_1 \logix.ram_r[192]$_DFFE_PP_  (.CLK(net454),
    .RESET_B(net1830),
    .D(_1039_),
    .Q_N(_4959_),
    .Q(\logix.ram_r[192] ));
 sg13g2_dfrbp_1 \logix.ram_r[1930]$_DFFE_PP_  (.CLK(net429),
    .RESET_B(net1831),
    .D(_1040_),
    .Q_N(_4958_),
    .Q(\logix.ram_r[1930] ));
 sg13g2_dfrbp_1 \logix.ram_r[1931]$_DFFE_PP_  (.CLK(net429),
    .RESET_B(net1832),
    .D(_1041_),
    .Q_N(_4957_),
    .Q(\logix.ram_r[1931] ));
 sg13g2_dfrbp_1 \logix.ram_r[1932]$_DFFE_PP_  (.CLK(net427),
    .RESET_B(net1833),
    .D(_1042_),
    .Q_N(_4956_),
    .Q(\logix.ram_r[1932] ));
 sg13g2_dfrbp_1 \logix.ram_r[1933]$_DFFE_PP_  (.CLK(net427),
    .RESET_B(net1834),
    .D(_1043_),
    .Q_N(_4955_),
    .Q(\logix.ram_r[1933] ));
 sg13g2_dfrbp_1 \logix.ram_r[1934]$_DFFE_PP_  (.CLK(net433),
    .RESET_B(net1835),
    .D(_1044_),
    .Q_N(_4954_),
    .Q(\logix.ram_r[1934] ));
 sg13g2_dfrbp_1 \logix.ram_r[1935]$_DFFE_PP_  (.CLK(net434),
    .RESET_B(net1836),
    .D(_1045_),
    .Q_N(_4953_),
    .Q(\logix.ram_r[1935] ));
 sg13g2_dfrbp_1 \logix.ram_r[1936]$_DFFE_PP_  (.CLK(net436),
    .RESET_B(net1837),
    .D(_1046_),
    .Q_N(_4952_),
    .Q(\logix.ram_r[1936] ));
 sg13g2_dfrbp_1 \logix.ram_r[1937]$_DFFE_PP_  (.CLK(net453),
    .RESET_B(net1838),
    .D(_1047_),
    .Q_N(_4951_),
    .Q(\logix.ram_r[1937] ));
 sg13g2_dfrbp_1 \logix.ram_r[1938]$_DFFE_PP_  (.CLK(net431),
    .RESET_B(net1839),
    .D(_1048_),
    .Q_N(_4950_),
    .Q(\logix.ram_r[1938] ));
 sg13g2_dfrbp_1 \logix.ram_r[1939]$_DFFE_PP_  (.CLK(net431),
    .RESET_B(net1840),
    .D(_1049_),
    .Q_N(_4949_),
    .Q(\logix.ram_r[1939] ));
 sg13g2_dfrbp_1 \logix.ram_r[193]$_DFFE_PP_  (.CLK(net453),
    .RESET_B(net1841),
    .D(_1050_),
    .Q_N(_4948_),
    .Q(\logix.ram_r[193] ));
 sg13g2_dfrbp_1 \logix.ram_r[1940]$_DFFE_PP_  (.CLK(net428),
    .RESET_B(net1842),
    .D(_1051_),
    .Q_N(_4947_),
    .Q(\logix.ram_r[1940] ));
 sg13g2_dfrbp_1 \logix.ram_r[1941]$_DFFE_PP_  (.CLK(net428),
    .RESET_B(net1843),
    .D(_1052_),
    .Q_N(_4946_),
    .Q(\logix.ram_r[1941] ));
 sg13g2_dfrbp_1 \logix.ram_r[1942]$_DFFE_PP_  (.CLK(net434),
    .RESET_B(net1844),
    .D(_1053_),
    .Q_N(_4945_),
    .Q(\logix.ram_r[1942] ));
 sg13g2_dfrbp_1 \logix.ram_r[1943]$_DFFE_PP_  (.CLK(net435),
    .RESET_B(net1845),
    .D(_1054_),
    .Q_N(_4944_),
    .Q(\logix.ram_r[1943] ));
 sg13g2_dfrbp_1 \logix.ram_r[1944]$_DFFE_PP_  (.CLK(net435),
    .RESET_B(net1846),
    .D(_1055_),
    .Q_N(_4943_),
    .Q(\logix.ram_r[1944] ));
 sg13g2_dfrbp_1 \logix.ram_r[1945]$_DFFE_PP_  (.CLK(net453),
    .RESET_B(net1847),
    .D(_1056_),
    .Q_N(_4942_),
    .Q(\logix.ram_r[1945] ));
 sg13g2_dfrbp_1 \logix.ram_r[1946]$_DFFE_PP_  (.CLK(net429),
    .RESET_B(net1848),
    .D(_1057_),
    .Q_N(_4941_),
    .Q(\logix.ram_r[1946] ));
 sg13g2_dfrbp_1 \logix.ram_r[1947]$_DFFE_PP_  (.CLK(net429),
    .RESET_B(net1849),
    .D(_1058_),
    .Q_N(_4940_),
    .Q(\logix.ram_r[1947] ));
 sg13g2_dfrbp_1 \logix.ram_r[1948]$_DFFE_PP_  (.CLK(net427),
    .RESET_B(net1850),
    .D(_1059_),
    .Q_N(_4939_),
    .Q(\logix.ram_r[1948] ));
 sg13g2_dfrbp_1 \logix.ram_r[1949]$_DFFE_PP_  (.CLK(net432),
    .RESET_B(net1851),
    .D(_1060_),
    .Q_N(_4938_),
    .Q(\logix.ram_r[1949] ));
 sg13g2_dfrbp_1 \logix.ram_r[194]$_DFFE_PP_  (.CLK(net436),
    .RESET_B(net1852),
    .D(_1061_),
    .Q_N(_4937_),
    .Q(\logix.ram_r[194] ));
 sg13g2_dfrbp_1 \logix.ram_r[1950]$_DFFE_PP_  (.CLK(net435),
    .RESET_B(net1853),
    .D(_1062_),
    .Q_N(_4936_),
    .Q(\logix.ram_r[1950] ));
 sg13g2_dfrbp_1 \logix.ram_r[1951]$_DFFE_PP_  (.CLK(net435),
    .RESET_B(net1854),
    .D(_1063_),
    .Q_N(_4935_),
    .Q(\logix.ram_r[1951] ));
 sg13g2_dfrbp_1 \logix.ram_r[1952]$_DFFE_PP_  (.CLK(net435),
    .RESET_B(net1855),
    .D(_1064_),
    .Q_N(_4934_),
    .Q(\logix.ram_r[1952] ));
 sg13g2_dfrbp_1 \logix.ram_r[1953]$_DFFE_PP_  (.CLK(net435),
    .RESET_B(net1856),
    .D(_1065_),
    .Q_N(_4933_),
    .Q(\logix.ram_r[1953] ));
 sg13g2_dfrbp_1 \logix.ram_r[1954]$_DFFE_PP_  (.CLK(net429),
    .RESET_B(net1857),
    .D(_1066_),
    .Q_N(_4932_),
    .Q(\logix.ram_r[1954] ));
 sg13g2_dfrbp_1 \logix.ram_r[1955]$_DFFE_PP_  (.CLK(net429),
    .RESET_B(net1858),
    .D(_1067_),
    .Q_N(_4931_),
    .Q(\logix.ram_r[1955] ));
 sg13g2_dfrbp_1 \logix.ram_r[1956]$_DFFE_PP_  (.CLK(net462),
    .RESET_B(net1859),
    .D(_1068_),
    .Q_N(_4930_),
    .Q(\logix.ram_r[1956] ));
 sg13g2_dfrbp_1 \logix.ram_r[1957]$_DFFE_PP_  (.CLK(net463),
    .RESET_B(net1860),
    .D(_1069_),
    .Q_N(_4929_),
    .Q(\logix.ram_r[1957] ));
 sg13g2_dfrbp_1 \logix.ram_r[1958]$_DFFE_PP_  (.CLK(net463),
    .RESET_B(net1861),
    .D(_1070_),
    .Q_N(_4928_),
    .Q(\logix.ram_r[1958] ));
 sg13g2_dfrbp_1 \logix.ram_r[1959]$_DFFE_PP_  (.CLK(net431),
    .RESET_B(net1862),
    .D(_1071_),
    .Q_N(_4927_),
    .Q(\logix.ram_r[1959] ));
 sg13g2_dfrbp_1 \logix.ram_r[195]$_DFFE_PP_  (.CLK(net436),
    .RESET_B(net1863),
    .D(_1072_),
    .Q_N(_4926_),
    .Q(\logix.ram_r[195] ));
 sg13g2_dfrbp_1 \logix.ram_r[1960]$_DFFE_PP_  (.CLK(net431),
    .RESET_B(net1864),
    .D(_1073_),
    .Q_N(_4925_),
    .Q(\logix.ram_r[1960] ));
 sg13g2_dfrbp_1 \logix.ram_r[1961]$_DFFE_PP_  (.CLK(net431),
    .RESET_B(net1865),
    .D(_1074_),
    .Q_N(_4924_),
    .Q(\logix.ram_r[1961] ));
 sg13g2_dfrbp_1 \logix.ram_r[1962]$_DFFE_PP_  (.CLK(net430),
    .RESET_B(net1866),
    .D(_1075_),
    .Q_N(_4923_),
    .Q(\logix.ram_r[1962] ));
 sg13g2_dfrbp_1 \logix.ram_r[1963]$_DFFE_PP_  (.CLK(net430),
    .RESET_B(net1867),
    .D(_1076_),
    .Q_N(_4922_),
    .Q(\logix.ram_r[1963] ));
 sg13g2_dfrbp_1 \logix.ram_r[1964]$_DFFE_PP_  (.CLK(net462),
    .RESET_B(net1868),
    .D(_1077_),
    .Q_N(_4921_),
    .Q(\logix.ram_r[1964] ));
 sg13g2_dfrbp_1 \logix.ram_r[1965]$_DFFE_PP_  (.CLK(net462),
    .RESET_B(net1869),
    .D(_1078_),
    .Q_N(_4920_),
    .Q(\logix.ram_r[1965] ));
 sg13g2_dfrbp_1 \logix.ram_r[1966]$_DFFE_PP_  (.CLK(net467),
    .RESET_B(net1870),
    .D(_1079_),
    .Q_N(_4919_),
    .Q(\logix.ram_r[1966] ));
 sg13g2_dfrbp_1 \logix.ram_r[1967]$_DFFE_PP_  (.CLK(net467),
    .RESET_B(net1871),
    .D(_1080_),
    .Q_N(_4918_),
    .Q(\logix.ram_r[1967] ));
 sg13g2_dfrbp_1 \logix.ram_r[1968]$_DFFE_PP_  (.CLK(net435),
    .RESET_B(net1872),
    .D(_1081_),
    .Q_N(_4917_),
    .Q(\logix.ram_r[1968] ));
 sg13g2_dfrbp_1 \logix.ram_r[1969]$_DFFE_PP_  (.CLK(net435),
    .RESET_B(net1873),
    .D(_1082_),
    .Q_N(_4916_),
    .Q(\logix.ram_r[1969] ));
 sg13g2_dfrbp_1 \logix.ram_r[196]$_DFFE_PP_  (.CLK(net436),
    .RESET_B(net1874),
    .D(_1083_),
    .Q_N(_4915_),
    .Q(\logix.ram_r[196] ));
 sg13g2_dfrbp_1 \logix.ram_r[1970]$_DFFE_PP_  (.CLK(net430),
    .RESET_B(net1875),
    .D(_1084_),
    .Q_N(_4914_),
    .Q(\logix.ram_r[1970] ));
 sg13g2_dfrbp_1 \logix.ram_r[1971]$_DFFE_PP_  (.CLK(net462),
    .RESET_B(net1876),
    .D(_1085_),
    .Q_N(_4913_),
    .Q(\logix.ram_r[1971] ));
 sg13g2_dfrbp_1 \logix.ram_r[1972]$_DFFE_PP_  (.CLK(net462),
    .RESET_B(net1877),
    .D(_1086_),
    .Q_N(_4912_),
    .Q(\logix.ram_r[1972] ));
 sg13g2_dfrbp_1 \logix.ram_r[1973]$_DFFE_PP_  (.CLK(net463),
    .RESET_B(net1878),
    .D(_1087_),
    .Q_N(_4911_),
    .Q(\logix.ram_r[1973] ));
 sg13g2_dfrbp_1 \logix.ram_r[1974]$_DFFE_PP_  (.CLK(net463),
    .RESET_B(net1879),
    .D(_1088_),
    .Q_N(_4910_),
    .Q(\logix.ram_r[1974] ));
 sg13g2_dfrbp_1 \logix.ram_r[1975]$_DFFE_PP_  (.CLK(net431),
    .RESET_B(net1880),
    .D(_1089_),
    .Q_N(_4909_),
    .Q(\logix.ram_r[1975] ));
 sg13g2_dfrbp_1 \logix.ram_r[1976]$_DFFE_PP_  (.CLK(net436),
    .RESET_B(net1881),
    .D(_1090_),
    .Q_N(_4908_),
    .Q(\logix.ram_r[1976] ));
 sg13g2_dfrbp_1 \logix.ram_r[1977]$_DFFE_PP_  (.CLK(net432),
    .RESET_B(net1882),
    .D(_1091_),
    .Q_N(_4907_),
    .Q(\logix.ram_r[1977] ));
 sg13g2_dfrbp_1 \logix.ram_r[1978]$_DFFE_PP_  (.CLK(net430),
    .RESET_B(net1883),
    .D(_1092_),
    .Q_N(_4906_),
    .Q(\logix.ram_r[1978] ));
 sg13g2_dfrbp_1 \logix.ram_r[1979]$_DFFE_PP_  (.CLK(net462),
    .RESET_B(net1884),
    .D(_1093_),
    .Q_N(_4905_),
    .Q(\logix.ram_r[1979] ));
 sg13g2_dfrbp_1 \logix.ram_r[197]$_DFFE_PP_  (.CLK(net468),
    .RESET_B(net1885),
    .D(_1094_),
    .Q_N(_4904_),
    .Q(\logix.ram_r[197] ));
 sg13g2_dfrbp_1 \logix.ram_r[1980]$_DFFE_PP_  (.CLK(net463),
    .RESET_B(net1886),
    .D(_1095_),
    .Q_N(_4903_),
    .Q(\logix.ram_r[1980] ));
 sg13g2_dfrbp_1 \logix.ram_r[1981]$_DFFE_PP_  (.CLK(net463),
    .RESET_B(net1887),
    .D(_1096_),
    .Q_N(_4902_),
    .Q(\logix.ram_r[1981] ));
 sg13g2_dfrbp_1 \logix.ram_r[1982]$_DFFE_PP_  (.CLK(net467),
    .RESET_B(net1888),
    .D(_1097_),
    .Q_N(_4901_),
    .Q(\logix.ram_r[1982] ));
 sg13g2_dfrbp_1 \logix.ram_r[1983]$_DFFE_PP_  (.CLK(net467),
    .RESET_B(net1889),
    .D(_1098_),
    .Q_N(_4900_),
    .Q(\logix.ram_r[1983] ));
 sg13g2_dfrbp_1 \logix.ram_r[1984]$_DFFE_PP_  (.CLK(net468),
    .RESET_B(net1890),
    .D(_1099_),
    .Q_N(_4899_),
    .Q(\logix.ram_r[1984] ));
 sg13g2_dfrbp_1 \logix.ram_r[1985]$_DFFE_PP_  (.CLK(net468),
    .RESET_B(net1891),
    .D(_1100_),
    .Q_N(_4898_),
    .Q(\logix.ram_r[1985] ));
 sg13g2_dfrbp_1 \logix.ram_r[1986]$_DFFE_PP_  (.CLK(net463),
    .RESET_B(net1892),
    .D(_1101_),
    .Q_N(_4897_),
    .Q(\logix.ram_r[1986] ));
 sg13g2_dfrbp_1 \logix.ram_r[1987]$_DFFE_PP_  (.CLK(net467),
    .RESET_B(net1893),
    .D(_1102_),
    .Q_N(_4896_),
    .Q(\logix.ram_r[1987] ));
 sg13g2_dfrbp_1 \logix.ram_r[1988]$_DFFE_PP_  (.CLK(net467),
    .RESET_B(net1894),
    .D(_1103_),
    .Q_N(_4895_),
    .Q(\logix.ram_r[1988] ));
 sg13g2_dfrbp_1 \logix.ram_r[1989]$_DFFE_PP_  (.CLK(net467),
    .RESET_B(net1895),
    .D(_1104_),
    .Q_N(_4894_),
    .Q(\logix.ram_r[1989] ));
 sg13g2_dfrbp_1 \logix.ram_r[198]$_DFFE_PP_  (.CLK(net468),
    .RESET_B(net1896),
    .D(_1105_),
    .Q_N(_4893_),
    .Q(\logix.ram_r[198] ));
 sg13g2_dfrbp_1 \logix.ram_r[1990]$_DFFE_PP_  (.CLK(net469),
    .RESET_B(net1897),
    .D(_1106_),
    .Q_N(_4892_),
    .Q(\logix.ram_r[1990] ));
 sg13g2_dfrbp_1 \logix.ram_r[1991]$_DFFE_PP_  (.CLK(net470),
    .RESET_B(net1898),
    .D(_1107_),
    .Q_N(_4891_),
    .Q(\logix.ram_r[1991] ));
 sg13g2_dfrbp_1 \logix.ram_r[1992]$_DFFE_PP_  (.CLK(net470),
    .RESET_B(net1899),
    .D(_1108_),
    .Q_N(_4890_),
    .Q(\logix.ram_r[1992] ));
 sg13g2_dfrbp_1 \logix.ram_r[1993]$_DFFE_PP_  (.CLK(net470),
    .RESET_B(net1900),
    .D(_1109_),
    .Q_N(_4889_),
    .Q(\logix.ram_r[1993] ));
 sg13g2_dfrbp_1 \logix.ram_r[1994]$_DFFE_PP_  (.CLK(net469),
    .RESET_B(net1901),
    .D(_1110_),
    .Q_N(_4888_),
    .Q(\logix.ram_r[1994] ));
 sg13g2_dfrbp_1 \logix.ram_r[1995]$_DFFE_PP_  (.CLK(net469),
    .RESET_B(net1902),
    .D(_1111_),
    .Q_N(_4887_),
    .Q(\logix.ram_r[1995] ));
 sg13g2_dfrbp_1 \logix.ram_r[1996]$_DFFE_PP_  (.CLK(net469),
    .RESET_B(net1903),
    .D(_1112_),
    .Q_N(_4886_),
    .Q(\logix.ram_r[1996] ));
 sg13g2_dfrbp_1 \logix.ram_r[1997]$_DFFE_PP_  (.CLK(net469),
    .RESET_B(net1904),
    .D(_1113_),
    .Q_N(_4885_),
    .Q(\logix.ram_r[1997] ));
 sg13g2_dfrbp_1 \logix.ram_r[1998]$_DFFE_PP_  (.CLK(net470),
    .RESET_B(net1905),
    .D(_1114_),
    .Q_N(_4884_),
    .Q(\logix.ram_r[1998] ));
 sg13g2_dfrbp_1 \logix.ram_r[1999]$_DFFE_PP_  (.CLK(net470),
    .RESET_B(net1906),
    .D(_1115_),
    .Q_N(_4883_),
    .Q(\logix.ram_r[1999] ));
 sg13g2_dfrbp_1 \logix.ram_r[199]$_DFFE_PP_  (.CLK(net486),
    .RESET_B(net1907),
    .D(_1116_),
    .Q_N(_4882_),
    .Q(\logix.ram_r[199] ));
 sg13g2_dfrbp_1 \logix.ram_r[19]$_DFFE_PP_  (.CLK(net640),
    .RESET_B(net1908),
    .D(_1117_),
    .Q_N(_4881_),
    .Q(\logix.ram_r[19] ));
 sg13g2_dfrbp_1 \logix.ram_r[1]$_DFFE_PP_  (.CLK(net657),
    .RESET_B(net1909),
    .D(_1118_),
    .Q_N(_4880_),
    .Q(\logix.ram_r[1] ));
 sg13g2_dfrbp_1 \logix.ram_r[2000]$_DFFE_PP_  (.CLK(net489),
    .RESET_B(net1910),
    .D(_1119_),
    .Q_N(_4879_),
    .Q(\logix.ram_r[2000] ));
 sg13g2_dfrbp_1 \logix.ram_r[2001]$_DFFE_PP_  (.CLK(net489),
    .RESET_B(net1911),
    .D(_1120_),
    .Q_N(_4878_),
    .Q(\logix.ram_r[2001] ));
 sg13g2_dfrbp_1 \logix.ram_r[2002]$_DFFE_PP_  (.CLK(net466),
    .RESET_B(net1912),
    .D(_1121_),
    .Q_N(_4877_),
    .Q(\logix.ram_r[2002] ));
 sg13g2_dfrbp_1 \logix.ram_r[2003]$_DFFE_PP_  (.CLK(net469),
    .RESET_B(net1913),
    .D(_1122_),
    .Q_N(_4876_),
    .Q(\logix.ram_r[2003] ));
 sg13g2_dfrbp_1 \logix.ram_r[2004]$_DFFE_PP_  (.CLK(net469),
    .RESET_B(net1914),
    .D(_1123_),
    .Q_N(_4875_),
    .Q(\logix.ram_r[2004] ));
 sg13g2_dfrbp_1 \logix.ram_r[2005]$_DFFE_PP_  (.CLK(net481),
    .RESET_B(net1915),
    .D(_1124_),
    .Q_N(_4874_),
    .Q(\logix.ram_r[2005] ));
 sg13g2_dfrbp_1 \logix.ram_r[2006]$_DFFE_PP_  (.CLK(net481),
    .RESET_B(net1916),
    .D(_1125_),
    .Q_N(_4873_),
    .Q(\logix.ram_r[2006] ));
 sg13g2_dfrbp_1 \logix.ram_r[2007]$_DFFE_PP_  (.CLK(net495),
    .RESET_B(net1917),
    .D(_1126_),
    .Q_N(_4872_),
    .Q(\logix.ram_r[2007] ));
 sg13g2_dfrbp_1 \logix.ram_r[2008]$_DFFE_PP_  (.CLK(net495),
    .RESET_B(net1918),
    .D(_1127_),
    .Q_N(_4871_),
    .Q(\logix.ram_r[2008] ));
 sg13g2_dfrbp_1 \logix.ram_r[2009]$_DFFE_PP_  (.CLK(net495),
    .RESET_B(net1919),
    .D(_1128_),
    .Q_N(_4870_),
    .Q(\logix.ram_r[2009] ));
 sg13g2_dfrbp_1 \logix.ram_r[200]$_DFFE_PP_  (.CLK(net486),
    .RESET_B(net1920),
    .D(_1129_),
    .Q_N(_4869_),
    .Q(\logix.ram_r[200] ));
 sg13g2_dfrbp_1 \logix.ram_r[2010]$_DFFE_PP_  (.CLK(net466),
    .RESET_B(net1921),
    .D(_1130_),
    .Q_N(_4868_),
    .Q(\logix.ram_r[2010] ));
 sg13g2_dfrbp_1 \logix.ram_r[2011]$_DFFE_PP_  (.CLK(net466),
    .RESET_B(net1922),
    .D(_1131_),
    .Q_N(_4867_),
    .Q(\logix.ram_r[2011] ));
 sg13g2_dfrbp_1 \logix.ram_r[2012]$_DFFE_PP_  (.CLK(net469),
    .RESET_B(net1923),
    .D(_1132_),
    .Q_N(_4866_),
    .Q(\logix.ram_r[2012] ));
 sg13g2_dfrbp_1 \logix.ram_r[2013]$_DFFE_PP_  (.CLK(net470),
    .RESET_B(net1924),
    .D(_1133_),
    .Q_N(_4865_),
    .Q(\logix.ram_r[2013] ));
 sg13g2_dfrbp_1 \logix.ram_r[2014]$_DFFE_PP_  (.CLK(net470),
    .RESET_B(net1925),
    .D(_1134_),
    .Q_N(_4864_),
    .Q(\logix.ram_r[2014] ));
 sg13g2_dfrbp_1 \logix.ram_r[2015]$_DFFE_PP_  (.CLK(net471),
    .RESET_B(net1926),
    .D(_1135_),
    .Q_N(_4863_),
    .Q(\logix.ram_r[2015] ));
 sg13g2_dfrbp_1 \logix.ram_r[2016]$_DFFE_PP_  (.CLK(net465),
    .RESET_B(net1927),
    .D(_1136_),
    .Q_N(_4862_),
    .Q(\logix.ram_r[2016] ));
 sg13g2_dfrbp_1 \logix.ram_r[2017]$_DFFE_PP_  (.CLK(net473),
    .RESET_B(net1928),
    .D(_1137_),
    .Q_N(_4861_),
    .Q(\logix.ram_r[2017] ));
 sg13g2_dfrbp_1 \logix.ram_r[2018]$_DFFE_PP_  (.CLK(net475),
    .RESET_B(net1929),
    .D(_1138_),
    .Q_N(_4860_),
    .Q(\logix.ram_r[2018] ));
 sg13g2_dfrbp_1 \logix.ram_r[2019]$_DFFE_PP_  (.CLK(net475),
    .RESET_B(net1930),
    .D(_1139_),
    .Q_N(_4859_),
    .Q(\logix.ram_r[2019] ));
 sg13g2_dfrbp_1 \logix.ram_r[201]$_DFFE_PP_  (.CLK(net468),
    .RESET_B(net1931),
    .D(_1140_),
    .Q_N(_4858_),
    .Q(\logix.ram_r[201] ));
 sg13g2_dfrbp_1 \logix.ram_r[2020]$_DFFE_PP_  (.CLK(net480),
    .RESET_B(net1932),
    .D(_1141_),
    .Q_N(_4857_),
    .Q(\logix.ram_r[2020] ));
 sg13g2_dfrbp_1 \logix.ram_r[2021]$_DFFE_PP_  (.CLK(net480),
    .RESET_B(net1933),
    .D(_1142_),
    .Q_N(_4856_),
    .Q(\logix.ram_r[2021] ));
 sg13g2_dfrbp_1 \logix.ram_r[2022]$_DFFE_PP_  (.CLK(net481),
    .RESET_B(net1934),
    .D(_1143_),
    .Q_N(_4855_),
    .Q(\logix.ram_r[2022] ));
 sg13g2_dfrbp_1 \logix.ram_r[2023]$_DFFE_PP_  (.CLK(net481),
    .RESET_B(net1935),
    .D(_1144_),
    .Q_N(_4854_),
    .Q(\logix.ram_r[2023] ));
 sg13g2_dfrbp_1 \logix.ram_r[2024]$_DFFE_PP_  (.CLK(net473),
    .RESET_B(net1936),
    .D(_1145_),
    .Q_N(_4853_),
    .Q(\logix.ram_r[2024] ));
 sg13g2_dfrbp_1 \logix.ram_r[2025]$_DFFE_PP_  (.CLK(net473),
    .RESET_B(net1937),
    .D(_1146_),
    .Q_N(_4852_),
    .Q(\logix.ram_r[2025] ));
 sg13g2_dfrbp_1 \logix.ram_r[2026]$_DFFE_PP_  (.CLK(net473),
    .RESET_B(net1938),
    .D(_1147_),
    .Q_N(_4851_),
    .Q(\logix.ram_r[2026] ));
 sg13g2_dfrbp_1 \logix.ram_r[2027]$_DFFE_PP_  (.CLK(net473),
    .RESET_B(net1939),
    .D(_1148_),
    .Q_N(_4850_),
    .Q(\logix.ram_r[2027] ));
 sg13g2_dfrbp_1 \logix.ram_r[2028]$_DFFE_PP_  (.CLK(net473),
    .RESET_B(net1940),
    .D(_1149_),
    .Q_N(_4849_),
    .Q(\logix.ram_r[2028] ));
 sg13g2_dfrbp_1 \logix.ram_r[2029]$_DFFE_PP_  (.CLK(net465),
    .RESET_B(net1941),
    .D(_1150_),
    .Q_N(_4848_),
    .Q(\logix.ram_r[2029] ));
 sg13g2_dfrbp_1 \logix.ram_r[202]$_DFFE_PP_  (.CLK(net468),
    .RESET_B(net1942),
    .D(_1151_),
    .Q_N(_4847_),
    .Q(\logix.ram_r[202] ));
 sg13g2_dfrbp_1 \logix.ram_r[2030]$_DFFE_PP_  (.CLK(net466),
    .RESET_B(net1943),
    .D(_1152_),
    .Q_N(_4846_),
    .Q(\logix.ram_r[2030] ));
 sg13g2_dfrbp_1 \logix.ram_r[2031]$_DFFE_PP_  (.CLK(net466),
    .RESET_B(net1944),
    .D(_1153_),
    .Q_N(_4845_),
    .Q(\logix.ram_r[2031] ));
 sg13g2_dfrbp_1 \logix.ram_r[2032]$_DFFE_PP_  (.CLK(net466),
    .RESET_B(net1945),
    .D(_1154_),
    .Q_N(_4844_),
    .Q(\logix.ram_r[2032] ));
 sg13g2_dfrbp_1 \logix.ram_r[2033]$_DFFE_PP_  (.CLK(net465),
    .RESET_B(net1946),
    .D(_1155_),
    .Q_N(_4843_),
    .Q(\logix.ram_r[2033] ));
 sg13g2_dfrbp_1 \logix.ram_r[2034]$_DFFE_PP_  (.CLK(net465),
    .RESET_B(net1947),
    .D(_1156_),
    .Q_N(_4842_),
    .Q(\logix.ram_r[2034] ));
 sg13g2_dfrbp_1 \logix.ram_r[2035]$_DFFE_PP_  (.CLK(net465),
    .RESET_B(net1948),
    .D(_1157_),
    .Q_N(_4841_),
    .Q(\logix.ram_r[2035] ));
 sg13g2_dfrbp_1 \logix.ram_r[2036]$_DFFE_PP_  (.CLK(net462),
    .RESET_B(net1949),
    .D(_1158_),
    .Q_N(_4840_),
    .Q(\logix.ram_r[2036] ));
 sg13g2_dfrbp_1 \logix.ram_r[2037]$_DFFE_PP_  (.CLK(net463),
    .RESET_B(net1950),
    .D(_1159_),
    .Q_N(_4839_),
    .Q(\logix.ram_r[2037] ));
 sg13g2_dfrbp_1 \logix.ram_r[2038]$_DFFE_PP_  (.CLK(net464),
    .RESET_B(net1951),
    .D(_1160_),
    .Q_N(_4838_),
    .Q(\logix.ram_r[2038] ));
 sg13g2_dfrbp_1 \logix.ram_r[2039]$_DFFE_PP_  (.CLK(net464),
    .RESET_B(net1952),
    .D(_1161_),
    .Q_N(_4837_),
    .Q(\logix.ram_r[2039] ));
 sg13g2_dfrbp_1 \logix.ram_r[203]$_DFFE_PP_  (.CLK(net468),
    .RESET_B(net1953),
    .D(_1162_),
    .Q_N(_4836_),
    .Q(\logix.ram_r[203] ));
 sg13g2_dfrbp_1 \logix.ram_r[2040]$_DFFE_PP_  (.CLK(net466),
    .RESET_B(net1954),
    .D(_1163_),
    .Q_N(_4835_),
    .Q(\logix.ram_r[2040] ));
 sg13g2_dfrbp_1 \logix.ram_r[2041]$_DFFE_PP_  (.CLK(net472),
    .RESET_B(net1955),
    .D(_1164_),
    .Q_N(_4834_),
    .Q(\logix.ram_r[2041] ));
 sg13g2_dfrbp_1 \logix.ram_r[2042]$_DFFE_PP_  (.CLK(net465),
    .RESET_B(net1956),
    .D(_1165_),
    .Q_N(_4833_),
    .Q(\logix.ram_r[2042] ));
 sg13g2_dfrbp_1 \logix.ram_r[2043]$_DFFE_PP_  (.CLK(net465),
    .RESET_B(net1957),
    .D(_1166_),
    .Q_N(_4832_),
    .Q(\logix.ram_r[2043] ));
 sg13g2_dfrbp_1 \logix.ram_r[2044]$_DFFE_PP_  (.CLK(net465),
    .RESET_B(net1958),
    .D(_1167_),
    .Q_N(_4831_),
    .Q(\logix.ram_r[2044] ));
 sg13g2_dfrbp_1 \logix.ram_r[2045]$_DFFE_PP_  (.CLK(net462),
    .RESET_B(net1959),
    .D(_1168_),
    .Q_N(_4830_),
    .Q(\logix.ram_r[2045] ));
 sg13g2_dfrbp_1 \logix.ram_r[2046]$_DFFE_PP_  (.CLK(net464),
    .RESET_B(net1960),
    .D(_1169_),
    .Q_N(_4829_),
    .Q(\logix.ram_r[2046] ));
 sg13g2_dfrbp_1 \logix.ram_r[2047]$_DFFE_PP_  (.CLK(net464),
    .RESET_B(net1961),
    .D(_1170_),
    .Q_N(_4828_),
    .Q(\logix.ram_r[2047] ));
 sg13g2_dfrbp_1 \logix.ram_r[2048]$_DFFE_PP_  (.CLK(net477),
    .RESET_B(net1962),
    .D(_1171_),
    .Q_N(_4827_),
    .Q(\logix.input_sel_cfg_w[0] ));
 sg13g2_dfrbp_1 \logix.ram_r[2049]$_DFFE_PP_  (.CLK(net484),
    .RESET_B(net1963),
    .D(_1172_),
    .Q_N(_4826_),
    .Q(\logix.input_sel_cfg_w[1] ));
 sg13g2_dfrbp_1 \logix.ram_r[204]$_DFFE_PP_  (.CLK(net486),
    .RESET_B(net1964),
    .D(_1173_),
    .Q_N(_4825_),
    .Q(\logix.ram_r[204] ));
 sg13g2_dfrbp_1 \logix.ram_r[2050]$_DFFE_PP_  (.CLK(net503),
    .RESET_B(net1965),
    .D(_1174_),
    .Q_N(_4824_),
    .Q(\logix.input_sel_cfg_w[2] ));
 sg13g2_dfrbp_1 \logix.ram_r[2051]$_DFFE_PP_  (.CLK(net503),
    .RESET_B(net1966),
    .D(_1175_),
    .Q_N(_4823_),
    .Q(\logix.input_sel_cfg_w[3] ));
 sg13g2_dfrbp_1 \logix.ram_r[2052]$_DFFE_PP_  (.CLK(net504),
    .RESET_B(net1967),
    .D(_1176_),
    .Q_N(_4822_),
    .Q(\logix.input_sel_cfg_w[4] ));
 sg13g2_dfrbp_1 \logix.ram_r[2053]$_DFFE_PP_  (.CLK(net504),
    .RESET_B(net1968),
    .D(_1177_),
    .Q_N(_4821_),
    .Q(\logix.input_sel_cfg_w[5] ));
 sg13g2_dfrbp_1 \logix.ram_r[2054]$_DFFE_PP_  (.CLK(net504),
    .RESET_B(net1969),
    .D(_1178_),
    .Q_N(_4820_),
    .Q(\logix.input_sel_cfg_w[6] ));
 sg13g2_dfrbp_1 \logix.ram_r[2055]$_DFFE_PP_  (.CLK(net497),
    .RESET_B(net1970),
    .D(_1179_),
    .Q_N(_4819_),
    .Q(\logix.input_sel_cfg_w[7] ));
 sg13g2_dfrbp_1 \logix.ram_r[205]$_DFFE_PP_  (.CLK(net486),
    .RESET_B(net1971),
    .D(_1180_),
    .Q_N(_4818_),
    .Q(\logix.ram_r[205] ));
 sg13g2_dfrbp_1 \logix.ram_r[206]$_DFFE_PP_  (.CLK(net487),
    .RESET_B(net1972),
    .D(_1181_),
    .Q_N(_4817_),
    .Q(\logix.ram_r[206] ));
 sg13g2_dfrbp_1 \logix.ram_r[207]$_DFFE_PP_  (.CLK(net491),
    .RESET_B(net1973),
    .D(_1182_),
    .Q_N(_4816_),
    .Q(\logix.ram_r[207] ));
 sg13g2_dfrbp_1 \logix.ram_r[208]$_DFFE_PP_  (.CLK(net458),
    .RESET_B(net1974),
    .D(_1183_),
    .Q_N(_4815_),
    .Q(\logix.ram_r[208] ));
 sg13g2_dfrbp_1 \logix.ram_r[209]$_DFFE_PP_  (.CLK(net454),
    .RESET_B(net1975),
    .D(_1184_),
    .Q_N(_4814_),
    .Q(\logix.ram_r[209] ));
 sg13g2_dfrbp_1 \logix.ram_r[20]$_DFFE_PP_  (.CLK(net639),
    .RESET_B(net1976),
    .D(_1185_),
    .Q_N(_4813_),
    .Q(\logix.ram_r[20] ));
 sg13g2_dfrbp_1 \logix.ram_r[210]$_DFFE_PP_  (.CLK(net454),
    .RESET_B(net1977),
    .D(_1186_),
    .Q_N(_4812_),
    .Q(\logix.ram_r[210] ));
 sg13g2_dfrbp_1 \logix.ram_r[211]$_DFFE_PP_  (.CLK(net436),
    .RESET_B(net1978),
    .D(_1187_),
    .Q_N(_4811_),
    .Q(\logix.ram_r[211] ));
 sg13g2_dfrbp_1 \logix.ram_r[212]$_DFFE_PP_  (.CLK(net453),
    .RESET_B(net1979),
    .D(_1188_),
    .Q_N(_4810_),
    .Q(\logix.ram_r[212] ));
 sg13g2_dfrbp_1 \logix.ram_r[213]$_DFFE_PP_  (.CLK(net486),
    .RESET_B(net1980),
    .D(_1189_),
    .Q_N(_4809_),
    .Q(\logix.ram_r[213] ));
 sg13g2_dfrbp_1 \logix.ram_r[214]$_DFFE_PP_  (.CLK(net490),
    .RESET_B(net1981),
    .D(_1190_),
    .Q_N(_4808_),
    .Q(\logix.ram_r[214] ));
 sg13g2_dfrbp_1 \logix.ram_r[215]$_DFFE_PP_  (.CLK(net491),
    .RESET_B(net1982),
    .D(_1191_),
    .Q_N(_4807_),
    .Q(\logix.ram_r[215] ));
 sg13g2_dfrbp_1 \logix.ram_r[216]$_DFFE_PP_  (.CLK(net458),
    .RESET_B(net1983),
    .D(_1192_),
    .Q_N(_4806_),
    .Q(\logix.ram_r[216] ));
 sg13g2_dfrbp_1 \logix.ram_r[217]$_DFFE_PP_  (.CLK(net454),
    .RESET_B(net1984),
    .D(_1193_),
    .Q_N(_4805_),
    .Q(\logix.ram_r[217] ));
 sg13g2_dfrbp_1 \logix.ram_r[218]$_DFFE_PP_  (.CLK(net453),
    .RESET_B(net1985),
    .D(_1194_),
    .Q_N(_4804_),
    .Q(\logix.ram_r[218] ));
 sg13g2_dfrbp_1 \logix.ram_r[219]$_DFFE_PP_  (.CLK(net453),
    .RESET_B(net1986),
    .D(_1195_),
    .Q_N(_4803_),
    .Q(\logix.ram_r[219] ));
 sg13g2_dfrbp_1 \logix.ram_r[21]$_DFFE_PP_  (.CLK(net639),
    .RESET_B(net1987),
    .D(_1196_),
    .Q_N(_4802_),
    .Q(\logix.ram_r[21] ));
 sg13g2_dfrbp_1 \logix.ram_r[220]$_DFFE_PP_  (.CLK(net454),
    .RESET_B(net1988),
    .D(_1197_),
    .Q_N(_4801_),
    .Q(\logix.ram_r[220] ));
 sg13g2_dfrbp_1 \logix.ram_r[221]$_DFFE_PP_  (.CLK(net454),
    .RESET_B(net1989),
    .D(_1198_),
    .Q_N(_4800_),
    .Q(\logix.ram_r[221] ));
 sg13g2_dfrbp_1 \logix.ram_r[222]$_DFFE_PP_  (.CLK(net454),
    .RESET_B(net1990),
    .D(_1199_),
    .Q_N(_4799_),
    .Q(\logix.ram_r[222] ));
 sg13g2_dfrbp_1 \logix.ram_r[223]$_DFFE_PP_  (.CLK(net458),
    .RESET_B(net1991),
    .D(_1200_),
    .Q_N(_4798_),
    .Q(\logix.ram_r[223] ));
 sg13g2_dfrbp_1 \logix.ram_r[224]$_DFFE_PP_  (.CLK(net455),
    .RESET_B(net1992),
    .D(_1201_),
    .Q_N(_4797_),
    .Q(\logix.ram_r[224] ));
 sg13g2_dfrbp_1 \logix.ram_r[225]$_DFFE_PP_  (.CLK(net452),
    .RESET_B(net1993),
    .D(_1202_),
    .Q_N(_4796_),
    .Q(\logix.ram_r[225] ));
 sg13g2_dfrbp_1 \logix.ram_r[226]$_DFFE_PP_  (.CLK(net452),
    .RESET_B(net1994),
    .D(_1203_),
    .Q_N(_4795_),
    .Q(\logix.ram_r[226] ));
 sg13g2_dfrbp_1 \logix.ram_r[227]$_DFFE_PP_  (.CLK(net452),
    .RESET_B(net1995),
    .D(_1204_),
    .Q_N(_4794_),
    .Q(\logix.ram_r[227] ));
 sg13g2_dfrbp_1 \logix.ram_r[228]$_DFFE_PP_  (.CLK(net455),
    .RESET_B(net1996),
    .D(_1205_),
    .Q_N(_4793_),
    .Q(\logix.ram_r[228] ));
 sg13g2_dfrbp_1 \logix.ram_r[229]$_DFFE_PP_  (.CLK(net458),
    .RESET_B(net1997),
    .D(_1206_),
    .Q_N(_4792_),
    .Q(\logix.ram_r[229] ));
 sg13g2_dfrbp_1 \logix.ram_r[22]$_DFFE_PP_  (.CLK(net609),
    .RESET_B(net1998),
    .D(_1207_),
    .Q_N(_4791_),
    .Q(\logix.ram_r[22] ));
 sg13g2_dfrbp_1 \logix.ram_r[230]$_DFFE_PP_  (.CLK(net459),
    .RESET_B(net1999),
    .D(_1208_),
    .Q_N(_4790_),
    .Q(\logix.ram_r[230] ));
 sg13g2_dfrbp_1 \logix.ram_r[231]$_DFFE_PP_  (.CLK(net521),
    .RESET_B(net2000),
    .D(_1209_),
    .Q_N(_4789_),
    .Q(\logix.ram_r[231] ));
 sg13g2_dfrbp_1 \logix.ram_r[232]$_DFFE_PP_  (.CLK(net518),
    .RESET_B(net2001),
    .D(_1210_),
    .Q_N(_4788_),
    .Q(\logix.ram_r[232] ));
 sg13g2_dfrbp_1 \logix.ram_r[233]$_DFFE_PP_  (.CLK(net457),
    .RESET_B(net2002),
    .D(_1211_),
    .Q_N(_4787_),
    .Q(\logix.ram_r[233] ));
 sg13g2_dfrbp_1 \logix.ram_r[234]$_DFFE_PP_  (.CLK(net456),
    .RESET_B(net2003),
    .D(_1212_),
    .Q_N(_4786_),
    .Q(\logix.ram_r[234] ));
 sg13g2_dfrbp_1 \logix.ram_r[235]$_DFFE_PP_  (.CLK(net456),
    .RESET_B(net2004),
    .D(_1213_),
    .Q_N(_4785_),
    .Q(\logix.ram_r[235] ));
 sg13g2_dfrbp_1 \logix.ram_r[236]$_DFFE_PP_  (.CLK(net458),
    .RESET_B(net2005),
    .D(_1214_),
    .Q_N(_4784_),
    .Q(\logix.ram_r[236] ));
 sg13g2_dfrbp_1 \logix.ram_r[237]$_DFFE_PP_  (.CLK(net458),
    .RESET_B(net2006),
    .D(_1215_),
    .Q_N(_4783_),
    .Q(\logix.ram_r[237] ));
 sg13g2_dfrbp_1 \logix.ram_r[238]$_DFFE_PP_  (.CLK(net459),
    .RESET_B(net2007),
    .D(_1216_),
    .Q_N(_4782_),
    .Q(\logix.ram_r[238] ));
 sg13g2_dfrbp_1 \logix.ram_r[239]$_DFFE_PP_  (.CLK(net521),
    .RESET_B(net2008),
    .D(_1217_),
    .Q_N(_4781_),
    .Q(\logix.ram_r[239] ));
 sg13g2_dfrbp_1 \logix.ram_r[23]$_DFFE_PP_  (.CLK(net604),
    .RESET_B(net2009),
    .D(_1218_),
    .Q_N(_4780_),
    .Q(\logix.ram_r[23] ));
 sg13g2_dfrbp_1 \logix.ram_r[240]$_DFFE_PP_  (.CLK(net518),
    .RESET_B(net2010),
    .D(_1219_),
    .Q_N(_4779_),
    .Q(\logix.ram_r[240] ));
 sg13g2_dfrbp_1 \logix.ram_r[241]$_DFFE_PP_  (.CLK(net457),
    .RESET_B(net2011),
    .D(_1220_),
    .Q_N(_4778_),
    .Q(\logix.ram_r[241] ));
 sg13g2_dfrbp_1 \logix.ram_r[242]$_DFFE_PP_  (.CLK(net456),
    .RESET_B(net2012),
    .D(_1221_),
    .Q_N(_4777_),
    .Q(\logix.ram_r[242] ));
 sg13g2_dfrbp_1 \logix.ram_r[243]$_DFFE_PP_  (.CLK(net456),
    .RESET_B(net2013),
    .D(_1222_),
    .Q_N(_4776_),
    .Q(\logix.ram_r[243] ));
 sg13g2_dfrbp_1 \logix.ram_r[244]$_DFFE_PP_  (.CLK(net458),
    .RESET_B(net2014),
    .D(_1223_),
    .Q_N(_4775_),
    .Q(\logix.ram_r[244] ));
 sg13g2_dfrbp_1 \logix.ram_r[245]$_DFFE_PP_  (.CLK(net459),
    .RESET_B(net2015),
    .D(_1224_),
    .Q_N(_4774_),
    .Q(\logix.ram_r[245] ));
 sg13g2_dfrbp_1 \logix.ram_r[246]$_DFFE_PP_  (.CLK(net459),
    .RESET_B(net2016),
    .D(_1225_),
    .Q_N(_4773_),
    .Q(\logix.ram_r[246] ));
 sg13g2_dfrbp_1 \logix.ram_r[247]$_DFFE_PP_  (.CLK(net521),
    .RESET_B(net2017),
    .D(_1226_),
    .Q_N(_4772_),
    .Q(\logix.ram_r[247] ));
 sg13g2_dfrbp_1 \logix.ram_r[248]$_DFFE_PP_  (.CLK(net518),
    .RESET_B(net2018),
    .D(_1227_),
    .Q_N(_4771_),
    .Q(\logix.ram_r[248] ));
 sg13g2_dfrbp_1 \logix.ram_r[249]$_DFFE_PP_  (.CLK(net457),
    .RESET_B(net2019),
    .D(_1228_),
    .Q_N(_4770_),
    .Q(\logix.ram_r[249] ));
 sg13g2_dfrbp_1 \logix.ram_r[24]$_DFFE_PP_  (.CLK(net605),
    .RESET_B(net2020),
    .D(_1229_),
    .Q_N(_4769_),
    .Q(\logix.ram_r[24] ));
 sg13g2_dfrbp_1 \logix.ram_r[250]$_DFFE_PP_  (.CLK(net456),
    .RESET_B(net2021),
    .D(_1230_),
    .Q_N(_4768_),
    .Q(\logix.ram_r[250] ));
 sg13g2_dfrbp_1 \logix.ram_r[251]$_DFFE_PP_  (.CLK(net457),
    .RESET_B(net2022),
    .D(_1231_),
    .Q_N(_4767_),
    .Q(\logix.ram_r[251] ));
 sg13g2_dfrbp_1 \logix.ram_r[252]$_DFFE_PP_  (.CLK(net459),
    .RESET_B(net2023),
    .D(_1232_),
    .Q_N(_4766_),
    .Q(\logix.ram_r[252] ));
 sg13g2_dfrbp_1 \logix.ram_r[253]$_DFFE_PP_  (.CLK(net459),
    .RESET_B(net2024),
    .D(_1233_),
    .Q_N(_4765_),
    .Q(\logix.ram_r[253] ));
 sg13g2_dfrbp_1 \logix.ram_r[254]$_DFFE_PP_  (.CLK(net521),
    .RESET_B(net2025),
    .D(_1234_),
    .Q_N(_4764_),
    .Q(\logix.ram_r[254] ));
 sg13g2_dfrbp_1 \logix.ram_r[255]$_DFFE_PP_  (.CLK(net521),
    .RESET_B(net2026),
    .D(_1235_),
    .Q_N(_4763_),
    .Q(\logix.ram_r[255] ));
 sg13g2_dfrbp_1 \logix.ram_r[256]$_DFFE_PP_  (.CLK(net545),
    .RESET_B(net2027),
    .D(_1236_),
    .Q_N(_4762_),
    .Q(\logix.ram_r[256] ));
 sg13g2_dfrbp_1 \logix.ram_r[257]$_DFFE_PP_  (.CLK(net664),
    .RESET_B(net2028),
    .D(_1237_),
    .Q_N(_4761_),
    .Q(\logix.ram_r[257] ));
 sg13g2_dfrbp_1 \logix.ram_r[258]$_DFFE_PP_  (.CLK(net665),
    .RESET_B(net2029),
    .D(_1238_),
    .Q_N(_4760_),
    .Q(\logix.ram_r[258] ));
 sg13g2_dfrbp_1 \logix.ram_r[259]$_DFFE_PP_  (.CLK(net729),
    .RESET_B(net2030),
    .D(_1239_),
    .Q_N(_4759_),
    .Q(\logix.ram_r[259] ));
 sg13g2_dfrbp_1 \logix.ram_r[25]$_DFFE_PP_  (.CLK(net659),
    .RESET_B(net2031),
    .D(_1240_),
    .Q_N(_4758_),
    .Q(\logix.ram_r[25] ));
 sg13g2_dfrbp_1 \logix.ram_r[260]$_DFFE_PP_  (.CLK(net737),
    .RESET_B(net2032),
    .D(_1241_),
    .Q_N(_4757_),
    .Q(\logix.ram_r[260] ));
 sg13g2_dfrbp_1 \logix.ram_r[261]$_DFFE_PP_  (.CLK(net737),
    .RESET_B(net2033),
    .D(_1242_),
    .Q_N(_4756_),
    .Q(\logix.ram_r[261] ));
 sg13g2_dfrbp_1 \logix.ram_r[262]$_DFFE_PP_  (.CLK(net673),
    .RESET_B(net2034),
    .D(_1243_),
    .Q_N(_4755_),
    .Q(\logix.ram_r[262] ));
 sg13g2_dfrbp_1 \logix.ram_r[263]$_DFFE_PP_  (.CLK(net664),
    .RESET_B(net2035),
    .D(_1244_),
    .Q_N(_4754_),
    .Q(\logix.ram_r[263] ));
 sg13g2_dfrbp_1 \logix.ram_r[264]$_DFFE_PP_  (.CLK(net664),
    .RESET_B(net2036),
    .D(_1245_),
    .Q_N(_4753_),
    .Q(\logix.ram_r[264] ));
 sg13g2_dfrbp_1 \logix.ram_r[265]$_DFFE_PP_  (.CLK(net665),
    .RESET_B(net2037),
    .D(_1246_),
    .Q_N(_4752_),
    .Q(\logix.ram_r[265] ));
 sg13g2_dfrbp_1 \logix.ram_r[266]$_DFFE_PP_  (.CLK(net729),
    .RESET_B(net2038),
    .D(_1247_),
    .Q_N(_4751_),
    .Q(\logix.ram_r[266] ));
 sg13g2_dfrbp_1 \logix.ram_r[267]$_DFFE_PP_  (.CLK(net729),
    .RESET_B(net2039),
    .D(_1248_),
    .Q_N(_4750_),
    .Q(\logix.ram_r[267] ));
 sg13g2_dfrbp_1 \logix.ram_r[268]$_DFFE_PP_  (.CLK(net728),
    .RESET_B(net2040),
    .D(_1249_),
    .Q_N(_4749_),
    .Q(\logix.ram_r[268] ));
 sg13g2_dfrbp_1 \logix.ram_r[269]$_DFFE_PP_  (.CLK(net666),
    .RESET_B(net2041),
    .D(_1250_),
    .Q_N(_4748_),
    .Q(\logix.ram_r[269] ));
 sg13g2_dfrbp_1 \logix.ram_r[26]$_DFFE_PP_  (.CLK(net660),
    .RESET_B(net2042),
    .D(_1251_),
    .Q_N(_4747_),
    .Q(\logix.ram_r[26] ));
 sg13g2_dfrbp_1 \logix.ram_r[270]$_DFFE_PP_  (.CLK(net660),
    .RESET_B(net2043),
    .D(_1252_),
    .Q_N(_4746_),
    .Q(\logix.ram_r[270] ));
 sg13g2_dfrbp_1 \logix.ram_r[271]$_DFFE_PP_  (.CLK(net660),
    .RESET_B(net2044),
    .D(_1253_),
    .Q_N(_4745_),
    .Q(\logix.ram_r[271] ));
 sg13g2_dfrbp_1 \logix.ram_r[272]$_DFFE_PP_  (.CLK(net660),
    .RESET_B(net2045),
    .D(_1254_),
    .Q_N(_4744_),
    .Q(\logix.ram_r[272] ));
 sg13g2_dfrbp_1 \logix.ram_r[273]$_DFFE_PP_  (.CLK(net664),
    .RESET_B(net2046),
    .D(_1255_),
    .Q_N(_4743_),
    .Q(\logix.ram_r[273] ));
 sg13g2_dfrbp_1 \logix.ram_r[274]$_DFFE_PP_  (.CLK(net665),
    .RESET_B(net2047),
    .D(_1256_),
    .Q_N(_4742_),
    .Q(\logix.ram_r[274] ));
 sg13g2_dfrbp_1 \logix.ram_r[275]$_DFFE_PP_  (.CLK(net729),
    .RESET_B(net2048),
    .D(_1257_),
    .Q_N(_4741_),
    .Q(\logix.ram_r[275] ));
 sg13g2_dfrbp_1 \logix.ram_r[276]$_DFFE_PP_  (.CLK(net737),
    .RESET_B(net2049),
    .D(_1258_),
    .Q_N(_4740_),
    .Q(\logix.ram_r[276] ));
 sg13g2_dfrbp_1 \logix.ram_r[277]$_DFFE_PP_  (.CLK(net737),
    .RESET_B(net2050),
    .D(_1259_),
    .Q_N(_4739_),
    .Q(\logix.ram_r[277] ));
 sg13g2_dfrbp_1 \logix.ram_r[278]$_DFFE_PP_  (.CLK(net673),
    .RESET_B(net2051),
    .D(_1260_),
    .Q_N(_4738_),
    .Q(\logix.ram_r[278] ));
 sg13g2_dfrbp_1 \logix.ram_r[279]$_DFFE_PP_  (.CLK(net665),
    .RESET_B(net2052),
    .D(_1261_),
    .Q_N(_4737_),
    .Q(\logix.ram_r[279] ));
 sg13g2_dfrbp_1 \logix.ram_r[27]$_DFFE_PP_  (.CLK(net660),
    .RESET_B(net2053),
    .D(_1262_),
    .Q_N(_4736_),
    .Q(\logix.ram_r[27] ));
 sg13g2_dfrbp_1 \logix.ram_r[280]$_DFFE_PP_  (.CLK(net665),
    .RESET_B(net2054),
    .D(_1263_),
    .Q_N(_4735_),
    .Q(\logix.ram_r[280] ));
 sg13g2_dfrbp_1 \logix.ram_r[281]$_DFFE_PP_  (.CLK(net666),
    .RESET_B(net2055),
    .D(_1264_),
    .Q_N(_4734_),
    .Q(\logix.ram_r[281] ));
 sg13g2_dfrbp_1 \logix.ram_r[282]$_DFFE_PP_  (.CLK(net729),
    .RESET_B(net2056),
    .D(_1265_),
    .Q_N(_4733_),
    .Q(\logix.ram_r[282] ));
 sg13g2_dfrbp_1 \logix.ram_r[283]$_DFFE_PP_  (.CLK(net728),
    .RESET_B(net2057),
    .D(_1266_),
    .Q_N(_4732_),
    .Q(\logix.ram_r[283] ));
 sg13g2_dfrbp_1 \logix.ram_r[284]$_DFFE_PP_  (.CLK(net728),
    .RESET_B(net2058),
    .D(_1267_),
    .Q_N(_4731_),
    .Q(\logix.ram_r[284] ));
 sg13g2_dfrbp_1 \logix.ram_r[285]$_DFFE_PP_  (.CLK(net736),
    .RESET_B(net2059),
    .D(_1268_),
    .Q_N(_4730_),
    .Q(\logix.ram_r[285] ));
 sg13g2_dfrbp_1 \logix.ram_r[286]$_DFFE_PP_  (.CLK(net668),
    .RESET_B(net2060),
    .D(_1269_),
    .Q_N(_4729_),
    .Q(\logix.ram_r[286] ));
 sg13g2_dfrbp_1 \logix.ram_r[287]$_DFFE_PP_  (.CLK(net668),
    .RESET_B(net2061),
    .D(_1270_),
    .Q_N(_4728_),
    .Q(\logix.ram_r[287] ));
 sg13g2_dfrbp_1 \logix.ram_r[288]$_DFFE_PP_  (.CLK(net669),
    .RESET_B(net2062),
    .D(_1271_),
    .Q_N(_4727_),
    .Q(\logix.ram_r[288] ));
 sg13g2_dfrbp_1 \logix.ram_r[289]$_DFFE_PP_  (.CLK(net673),
    .RESET_B(net2063),
    .D(_1272_),
    .Q_N(_4726_),
    .Q(\logix.ram_r[289] ));
 sg13g2_dfrbp_1 \logix.ram_r[28]$_DFFE_PP_  (.CLK(net660),
    .RESET_B(net2064),
    .D(_1273_),
    .Q_N(_4725_),
    .Q(\logix.ram_r[28] ));
 sg13g2_dfrbp_1 \logix.ram_r[290]$_DFFE_PP_  (.CLK(net674),
    .RESET_B(net2065),
    .D(_1274_),
    .Q_N(_4724_),
    .Q(\logix.ram_r[290] ));
 sg13g2_dfrbp_1 \logix.ram_r[291]$_DFFE_PP_  (.CLK(net737),
    .RESET_B(net2066),
    .D(_1275_),
    .Q_N(_4723_),
    .Q(\logix.ram_r[291] ));
 sg13g2_dfrbp_1 \logix.ram_r[292]$_DFFE_PP_  (.CLK(net736),
    .RESET_B(net2067),
    .D(_1276_),
    .Q_N(_4722_),
    .Q(\logix.ram_r[292] ));
 sg13g2_dfrbp_1 \logix.ram_r[293]$_DFFE_PP_  (.CLK(net736),
    .RESET_B(net2068),
    .D(_1277_),
    .Q_N(_4721_),
    .Q(\logix.ram_r[293] ));
 sg13g2_dfrbp_1 \logix.ram_r[294]$_DFFE_PP_  (.CLK(net736),
    .RESET_B(net2069),
    .D(_1278_),
    .Q_N(_4720_),
    .Q(\logix.ram_r[294] ));
 sg13g2_dfrbp_1 \logix.ram_r[295]$_DFFE_PP_  (.CLK(net674),
    .RESET_B(net2070),
    .D(_1279_),
    .Q_N(_4719_),
    .Q(\logix.ram_r[295] ));
 sg13g2_dfrbp_1 \logix.ram_r[296]$_DFFE_PP_  (.CLK(net673),
    .RESET_B(net2071),
    .D(_1280_),
    .Q_N(_4718_),
    .Q(\logix.ram_r[296] ));
 sg13g2_dfrbp_1 \logix.ram_r[297]$_DFFE_PP_  (.CLK(net674),
    .RESET_B(net2072),
    .D(_1281_),
    .Q_N(_4717_),
    .Q(\logix.ram_r[297] ));
 sg13g2_dfrbp_1 \logix.ram_r[298]$_DFFE_PP_  (.CLK(net674),
    .RESET_B(net2073),
    .D(_1282_),
    .Q_N(_4716_),
    .Q(\logix.ram_r[298] ));
 sg13g2_dfrbp_1 \logix.ram_r[299]$_DFFE_PP_  (.CLK(net737),
    .RESET_B(net2074),
    .D(_1283_),
    .Q_N(_4715_),
    .Q(\logix.ram_r[299] ));
 sg13g2_dfrbp_1 \logix.ram_r[29]$_DFFE_PP_  (.CLK(net659),
    .RESET_B(net2075),
    .D(_1284_),
    .Q_N(_4714_),
    .Q(\logix.ram_r[29] ));
 sg13g2_dfrbp_1 \logix.ram_r[2]$_DFFE_PP_  (.CLK(net657),
    .RESET_B(net2076),
    .D(_1285_),
    .Q_N(_4713_),
    .Q(\logix.ram_r[2] ));
 sg13g2_dfrbp_1 \logix.ram_r[300]$_DFFE_PP_  (.CLK(net736),
    .RESET_B(net2077),
    .D(_1286_),
    .Q_N(_4712_),
    .Q(\logix.ram_r[300] ));
 sg13g2_dfrbp_1 \logix.ram_r[301]$_DFFE_PP_  (.CLK(net736),
    .RESET_B(net2078),
    .D(_1287_),
    .Q_N(_4711_),
    .Q(\logix.ram_r[301] ));
 sg13g2_dfrbp_1 \logix.ram_r[302]$_DFFE_PP_  (.CLK(net669),
    .RESET_B(net2079),
    .D(_1288_),
    .Q_N(_4710_),
    .Q(\logix.ram_r[302] ));
 sg13g2_dfrbp_1 \logix.ram_r[303]$_DFFE_PP_  (.CLK(net669),
    .RESET_B(net2080),
    .D(_1289_),
    .Q_N(_4709_),
    .Q(\logix.ram_r[303] ));
 sg13g2_dfrbp_1 \logix.ram_r[304]$_DFFE_PP_  (.CLK(net673),
    .RESET_B(net2081),
    .D(_1290_),
    .Q_N(_4708_),
    .Q(\logix.ram_r[304] ));
 sg13g2_dfrbp_1 \logix.ram_r[305]$_DFFE_PP_  (.CLK(net673),
    .RESET_B(net2082),
    .D(_1291_),
    .Q_N(_4707_),
    .Q(\logix.ram_r[305] ));
 sg13g2_dfrbp_1 \logix.ram_r[306]$_DFFE_PP_  (.CLK(net674),
    .RESET_B(net2083),
    .D(_1292_),
    .Q_N(_4706_),
    .Q(\logix.ram_r[306] ));
 sg13g2_dfrbp_1 \logix.ram_r[307]$_DFFE_PP_  (.CLK(net737),
    .RESET_B(net2084),
    .D(_1293_),
    .Q_N(_4705_),
    .Q(\logix.ram_r[307] ));
 sg13g2_dfrbp_1 \logix.ram_r[308]$_DFFE_PP_  (.CLK(net736),
    .RESET_B(net2085),
    .D(_1294_),
    .Q_N(_4704_),
    .Q(\logix.ram_r[308] ));
 sg13g2_dfrbp_1 \logix.ram_r[309]$_DFFE_PP_  (.CLK(net738),
    .RESET_B(net2086),
    .D(_1295_),
    .Q_N(_4703_),
    .Q(\logix.ram_r[309] ));
 sg13g2_dfrbp_1 \logix.ram_r[30]$_DFFE_PP_  (.CLK(net660),
    .RESET_B(net2087),
    .D(_1296_),
    .Q_N(_4702_),
    .Q(\logix.ram_r[30] ));
 sg13g2_dfrbp_1 \logix.ram_r[310]$_DFFE_PP_  (.CLK(net736),
    .RESET_B(net2088),
    .D(_1297_),
    .Q_N(_4701_),
    .Q(\logix.ram_r[310] ));
 sg13g2_dfrbp_1 \logix.ram_r[311]$_DFFE_PP_  (.CLK(net674),
    .RESET_B(net2089),
    .D(_1298_),
    .Q_N(_4700_),
    .Q(\logix.ram_r[311] ));
 sg13g2_dfrbp_1 \logix.ram_r[312]$_DFFE_PP_  (.CLK(net673),
    .RESET_B(net2090),
    .D(_1299_),
    .Q_N(_4699_),
    .Q(\logix.ram_r[312] ));
 sg13g2_dfrbp_1 \logix.ram_r[313]$_DFFE_PP_  (.CLK(net674),
    .RESET_B(net2091),
    .D(_1300_),
    .Q_N(_4698_),
    .Q(\logix.ram_r[313] ));
 sg13g2_dfrbp_1 \logix.ram_r[314]$_DFFE_PP_  (.CLK(net737),
    .RESET_B(net2092),
    .D(_1301_),
    .Q_N(_4697_),
    .Q(\logix.ram_r[314] ));
 sg13g2_dfrbp_1 \logix.ram_r[315]$_DFFE_PP_  (.CLK(net738),
    .RESET_B(net2093),
    .D(_1302_),
    .Q_N(_4696_),
    .Q(\logix.ram_r[315] ));
 sg13g2_dfrbp_1 \logix.ram_r[316]$_DFFE_PP_  (.CLK(net738),
    .RESET_B(net2094),
    .D(_1303_),
    .Q_N(_4695_),
    .Q(\logix.ram_r[316] ));
 sg13g2_dfrbp_1 \logix.ram_r[317]$_DFFE_PP_  (.CLK(net743),
    .RESET_B(net2095),
    .D(_1304_),
    .Q_N(_4694_),
    .Q(\logix.ram_r[317] ));
 sg13g2_dfrbp_1 \logix.ram_r[318]$_DFFE_PP_  (.CLK(net743),
    .RESET_B(net2096),
    .D(_1305_),
    .Q_N(_4693_),
    .Q(\logix.ram_r[318] ));
 sg13g2_dfrbp_1 \logix.ram_r[319]$_DFFE_PP_  (.CLK(net669),
    .RESET_B(net2097),
    .D(_1306_),
    .Q_N(_4692_),
    .Q(\logix.ram_r[319] ));
 sg13g2_dfrbp_1 \logix.ram_r[31]$_DFFE_PP_  (.CLK(net656),
    .RESET_B(net2098),
    .D(_1307_),
    .Q_N(_4691_),
    .Q(\logix.ram_r[31] ));
 sg13g2_dfrbp_1 \logix.ram_r[320]$_DFFE_PP_  (.CLK(net671),
    .RESET_B(net2099),
    .D(_1308_),
    .Q_N(_4690_),
    .Q(\logix.ram_r[320] ));
 sg13g2_dfrbp_1 \logix.ram_r[321]$_DFFE_PP_  (.CLK(net670),
    .RESET_B(net2100),
    .D(_1309_),
    .Q_N(_4689_),
    .Q(\logix.ram_r[321] ));
 sg13g2_dfrbp_1 \logix.ram_r[322]$_DFFE_PP_  (.CLK(net654),
    .RESET_B(net2101),
    .D(_1310_),
    .Q_N(_4688_),
    .Q(\logix.ram_r[322] ));
 sg13g2_dfrbp_1 \logix.ram_r[323]$_DFFE_PP_  (.CLK(net654),
    .RESET_B(net2102),
    .D(_1311_),
    .Q_N(_4687_),
    .Q(\logix.ram_r[323] ));
 sg13g2_dfrbp_1 \logix.ram_r[324]$_DFFE_PP_  (.CLK(net670),
    .RESET_B(net2103),
    .D(_1312_),
    .Q_N(_4686_),
    .Q(\logix.ram_r[324] ));
 sg13g2_dfrbp_1 \logix.ram_r[325]$_DFFE_PP_  (.CLK(net670),
    .RESET_B(net2104),
    .D(_1313_),
    .Q_N(_4685_),
    .Q(\logix.ram_r[325] ));
 sg13g2_dfrbp_1 \logix.ram_r[326]$_DFFE_PP_  (.CLK(net671),
    .RESET_B(net2105),
    .D(_1314_),
    .Q_N(_4684_),
    .Q(\logix.ram_r[326] ));
 sg13g2_dfrbp_1 \logix.ram_r[327]$_DFFE_PP_  (.CLK(net671),
    .RESET_B(net2106),
    .D(_1315_),
    .Q_N(_4683_),
    .Q(\logix.ram_r[327] ));
 sg13g2_dfrbp_1 \logix.ram_r[328]$_DFFE_PP_  (.CLK(net671),
    .RESET_B(net2107),
    .D(_1316_),
    .Q_N(_4682_),
    .Q(\logix.ram_r[328] ));
 sg13g2_dfrbp_1 \logix.ram_r[329]$_DFFE_PP_  (.CLK(net670),
    .RESET_B(net2108),
    .D(_1317_),
    .Q_N(_4681_),
    .Q(\logix.ram_r[329] ));
 sg13g2_dfrbp_1 \logix.ram_r[32]$_DFFE_PP_  (.CLK(net656),
    .RESET_B(net2109),
    .D(_1318_),
    .Q_N(_4680_),
    .Q(\logix.ram_r[32] ));
 sg13g2_dfrbp_1 \logix.ram_r[330]$_DFFE_PP_  (.CLK(net654),
    .RESET_B(net2110),
    .D(_1319_),
    .Q_N(_4679_),
    .Q(\logix.ram_r[330] ));
 sg13g2_dfrbp_1 \logix.ram_r[331]$_DFFE_PP_  (.CLK(net654),
    .RESET_B(net2111),
    .D(_1320_),
    .Q_N(_4678_),
    .Q(\logix.ram_r[331] ));
 sg13g2_dfrbp_1 \logix.ram_r[332]$_DFFE_PP_  (.CLK(net654),
    .RESET_B(net2112),
    .D(_1321_),
    .Q_N(_4677_),
    .Q(\logix.ram_r[332] ));
 sg13g2_dfrbp_1 \logix.ram_r[333]$_DFFE_PP_  (.CLK(net670),
    .RESET_B(net2113),
    .D(_1322_),
    .Q_N(_4676_),
    .Q(\logix.ram_r[333] ));
 sg13g2_dfrbp_1 \logix.ram_r[334]$_DFFE_PP_  (.CLK(net670),
    .RESET_B(net2114),
    .D(_1323_),
    .Q_N(_4675_),
    .Q(\logix.ram_r[334] ));
 sg13g2_dfrbp_1 \logix.ram_r[335]$_DFFE_PP_  (.CLK(net676),
    .RESET_B(net2115),
    .D(_1324_),
    .Q_N(_4674_),
    .Q(\logix.ram_r[335] ));
 sg13g2_dfrbp_1 \logix.ram_r[336]$_DFFE_PP_  (.CLK(net676),
    .RESET_B(net2116),
    .D(_1325_),
    .Q_N(_4673_),
    .Q(\logix.ram_r[336] ));
 sg13g2_dfrbp_1 \logix.ram_r[337]$_DFFE_PP_  (.CLK(net676),
    .RESET_B(net2117),
    .D(_1326_),
    .Q_N(_4672_),
    .Q(\logix.ram_r[337] ));
 sg13g2_dfrbp_1 \logix.ram_r[338]$_DFFE_PP_  (.CLK(net654),
    .RESET_B(net2118),
    .D(_1327_),
    .Q_N(_4671_),
    .Q(\logix.ram_r[338] ));
 sg13g2_dfrbp_1 \logix.ram_r[339]$_DFFE_PP_  (.CLK(net654),
    .RESET_B(net2119),
    .D(_1328_),
    .Q_N(_4670_),
    .Q(\logix.ram_r[339] ));
 sg13g2_dfrbp_1 \logix.ram_r[33]$_DFFE_PP_  (.CLK(net668),
    .RESET_B(net2120),
    .D(_1329_),
    .Q_N(_4669_),
    .Q(\logix.ram_r[33] ));
 sg13g2_dfrbp_1 \logix.ram_r[340]$_DFFE_PP_  (.CLK(net670),
    .RESET_B(net2121),
    .D(_1330_),
    .Q_N(_4668_),
    .Q(\logix.ram_r[340] ));
 sg13g2_dfrbp_1 \logix.ram_r[341]$_DFFE_PP_  (.CLK(net670),
    .RESET_B(net2122),
    .D(_1331_),
    .Q_N(_4667_),
    .Q(\logix.ram_r[341] ));
 sg13g2_dfrbp_1 \logix.ram_r[342]$_DFFE_PP_  (.CLK(net671),
    .RESET_B(net2123),
    .D(_1332_),
    .Q_N(_4666_),
    .Q(\logix.ram_r[342] ));
 sg13g2_dfrbp_1 \logix.ram_r[343]$_DFFE_PP_  (.CLK(net671),
    .RESET_B(net2124),
    .D(_1333_),
    .Q_N(_4665_),
    .Q(\logix.ram_r[343] ));
 sg13g2_dfrbp_1 \logix.ram_r[344]$_DFFE_PP_  (.CLK(net671),
    .RESET_B(net2125),
    .D(_1334_),
    .Q_N(_4664_),
    .Q(\logix.ram_r[344] ));
 sg13g2_dfrbp_1 \logix.ram_r[345]$_DFFE_PP_  (.CLK(net671),
    .RESET_B(net2126),
    .D(_1335_),
    .Q_N(_4663_),
    .Q(\logix.ram_r[345] ));
 sg13g2_dfrbp_1 \logix.ram_r[346]$_DFFE_PP_  (.CLK(net654),
    .RESET_B(net2127),
    .D(_1336_),
    .Q_N(_4662_),
    .Q(\logix.ram_r[346] ));
 sg13g2_dfrbp_1 \logix.ram_r[347]$_DFFE_PP_  (.CLK(net655),
    .RESET_B(net2128),
    .D(_1337_),
    .Q_N(_4661_),
    .Q(\logix.ram_r[347] ));
 sg13g2_dfrbp_1 \logix.ram_r[348]$_DFFE_PP_  (.CLK(net672),
    .RESET_B(net2129),
    .D(_1338_),
    .Q_N(_4660_),
    .Q(\logix.ram_r[348] ));
 sg13g2_dfrbp_1 \logix.ram_r[349]$_DFFE_PP_  (.CLK(net672),
    .RESET_B(net2130),
    .D(_1339_),
    .Q_N(_4659_),
    .Q(\logix.ram_r[349] ));
 sg13g2_dfrbp_1 \logix.ram_r[34]$_DFFE_PP_  (.CLK(net668),
    .RESET_B(net2131),
    .D(_1340_),
    .Q_N(_4658_),
    .Q(\logix.ram_r[34] ));
 sg13g2_dfrbp_1 \logix.ram_r[350]$_DFFE_PP_  (.CLK(net672),
    .RESET_B(net2132),
    .D(_1341_),
    .Q_N(_4657_),
    .Q(\logix.ram_r[350] ));
 sg13g2_dfrbp_1 \logix.ram_r[351]$_DFFE_PP_  (.CLK(net676),
    .RESET_B(net2133),
    .D(_1342_),
    .Q_N(_4656_),
    .Q(\logix.ram_r[351] ));
 sg13g2_dfrbp_1 \logix.ram_r[352]$_DFFE_PP_  (.CLK(net676),
    .RESET_B(net2134),
    .D(_1343_),
    .Q_N(_4655_),
    .Q(\logix.ram_r[352] ));
 sg13g2_dfrbp_1 \logix.ram_r[353]$_DFFE_PP_  (.CLK(net675),
    .RESET_B(net2135),
    .D(_1344_),
    .Q_N(_4654_),
    .Q(\logix.ram_r[353] ));
 sg13g2_dfrbp_1 \logix.ram_r[354]$_DFFE_PP_  (.CLK(net675),
    .RESET_B(net2136),
    .D(_1345_),
    .Q_N(_4653_),
    .Q(\logix.ram_r[354] ));
 sg13g2_dfrbp_1 \logix.ram_r[355]$_DFFE_PP_  (.CLK(net675),
    .RESET_B(net2137),
    .D(_1346_),
    .Q_N(_4652_),
    .Q(\logix.ram_r[355] ));
 sg13g2_dfrbp_1 \logix.ram_r[356]$_DFFE_PP_  (.CLK(net739),
    .RESET_B(net2138),
    .D(_1347_),
    .Q_N(_4651_),
    .Q(\logix.ram_r[356] ));
 sg13g2_dfrbp_1 \logix.ram_r[357]$_DFFE_PP_  (.CLK(net739),
    .RESET_B(net2139),
    .D(_1348_),
    .Q_N(_4650_),
    .Q(\logix.ram_r[357] ));
 sg13g2_dfrbp_1 \logix.ram_r[358]$_DFFE_PP_  (.CLK(net739),
    .RESET_B(net2140),
    .D(_1349_),
    .Q_N(_4649_),
    .Q(\logix.ram_r[358] ));
 sg13g2_dfrbp_1 \logix.ram_r[359]$_DFFE_PP_  (.CLK(net740),
    .RESET_B(net2141),
    .D(_1350_),
    .Q_N(_4648_),
    .Q(\logix.ram_r[359] ));
 sg13g2_dfrbp_1 \logix.ram_r[35]$_DFFE_PP_  (.CLK(net668),
    .RESET_B(net2142),
    .D(_1351_),
    .Q_N(_4647_),
    .Q(\logix.ram_r[35] ));
 sg13g2_dfrbp_1 \logix.ram_r[360]$_DFFE_PP_  (.CLK(net740),
    .RESET_B(net2143),
    .D(_1352_),
    .Q_N(_4646_),
    .Q(\logix.ram_r[360] ));
 sg13g2_dfrbp_1 \logix.ram_r[361]$_DFFE_PP_  (.CLK(net740),
    .RESET_B(net2144),
    .D(_1353_),
    .Q_N(_4645_),
    .Q(\logix.ram_r[361] ));
 sg13g2_dfrbp_1 \logix.ram_r[362]$_DFFE_PP_  (.CLK(net739),
    .RESET_B(net2145),
    .D(_1354_),
    .Q_N(_4644_),
    .Q(\logix.ram_r[362] ));
 sg13g2_dfrbp_1 \logix.ram_r[363]$_DFFE_PP_  (.CLK(net739),
    .RESET_B(net2146),
    .D(_1355_),
    .Q_N(_4643_),
    .Q(\logix.ram_r[363] ));
 sg13g2_dfrbp_1 \logix.ram_r[364]$_DFFE_PP_  (.CLK(net739),
    .RESET_B(net2147),
    .D(_1356_),
    .Q_N(_4642_),
    .Q(\logix.ram_r[364] ));
 sg13g2_dfrbp_1 \logix.ram_r[365]$_DFFE_PP_  (.CLK(net675),
    .RESET_B(net2148),
    .D(_1357_),
    .Q_N(_4641_),
    .Q(\logix.ram_r[365] ));
 sg13g2_dfrbp_1 \logix.ram_r[366]$_DFFE_PP_  (.CLK(net675),
    .RESET_B(net2149),
    .D(_1358_),
    .Q_N(_4640_),
    .Q(\logix.ram_r[366] ));
 sg13g2_dfrbp_1 \logix.ram_r[367]$_DFFE_PP_  (.CLK(net676),
    .RESET_B(net2150),
    .D(_1359_),
    .Q_N(_4639_),
    .Q(\logix.ram_r[367] ));
 sg13g2_dfrbp_1 \logix.ram_r[368]$_DFFE_PP_  (.CLK(net676),
    .RESET_B(net2151),
    .D(_1360_),
    .Q_N(_4638_),
    .Q(\logix.ram_r[368] ));
 sg13g2_dfrbp_1 \logix.ram_r[369]$_DFFE_PP_  (.CLK(net675),
    .RESET_B(net2152),
    .D(_1361_),
    .Q_N(_4637_),
    .Q(\logix.ram_r[369] ));
 sg13g2_dfrbp_1 \logix.ram_r[36]$_DFFE_PP_  (.CLK(net669),
    .RESET_B(net2153),
    .D(_1362_),
    .Q_N(_4636_),
    .Q(\logix.ram_r[36] ));
 sg13g2_dfrbp_1 \logix.ram_r[370]$_DFFE_PP_  (.CLK(net675),
    .RESET_B(net2154),
    .D(_1363_),
    .Q_N(_4635_),
    .Q(\logix.ram_r[370] ));
 sg13g2_dfrbp_1 \logix.ram_r[371]$_DFFE_PP_  (.CLK(net675),
    .RESET_B(net2155),
    .D(_1364_),
    .Q_N(_4634_),
    .Q(\logix.ram_r[371] ));
 sg13g2_dfrbp_1 \logix.ram_r[372]$_DFFE_PP_  (.CLK(net677),
    .RESET_B(net2156),
    .D(_1365_),
    .Q_N(_4633_),
    .Q(\logix.ram_r[372] ));
 sg13g2_dfrbp_1 \logix.ram_r[373]$_DFFE_PP_  (.CLK(net739),
    .RESET_B(net2157),
    .D(_1366_),
    .Q_N(_4632_),
    .Q(\logix.ram_r[373] ));
 sg13g2_dfrbp_1 \logix.ram_r[374]$_DFFE_PP_  (.CLK(net740),
    .RESET_B(net2158),
    .D(_1367_),
    .Q_N(_4631_),
    .Q(\logix.ram_r[374] ));
 sg13g2_dfrbp_1 \logix.ram_r[375]$_DFFE_PP_  (.CLK(net740),
    .RESET_B(net2159),
    .D(_1368_),
    .Q_N(_4630_),
    .Q(\logix.ram_r[375] ));
 sg13g2_dfrbp_1 \logix.ram_r[376]$_DFFE_PP_  (.CLK(net740),
    .RESET_B(net2160),
    .D(_1369_),
    .Q_N(_4629_),
    .Q(\logix.ram_r[376] ));
 sg13g2_dfrbp_1 \logix.ram_r[377]$_DFFE_PP_  (.CLK(net740),
    .RESET_B(net2161),
    .D(_1370_),
    .Q_N(_4628_),
    .Q(\logix.ram_r[377] ));
 sg13g2_dfrbp_1 \logix.ram_r[378]$_DFFE_PP_  (.CLK(net744),
    .RESET_B(net2162),
    .D(_1371_),
    .Q_N(_4627_),
    .Q(\logix.ram_r[378] ));
 sg13g2_dfrbp_1 \logix.ram_r[379]$_DFFE_PP_  (.CLK(net741),
    .RESET_B(net2163),
    .D(_1372_),
    .Q_N(_4626_),
    .Q(\logix.ram_r[379] ));
 sg13g2_dfrbp_1 \logix.ram_r[37]$_DFFE_PP_  (.CLK(net669),
    .RESET_B(net2164),
    .D(_1373_),
    .Q_N(_4625_),
    .Q(\logix.ram_r[37] ));
 sg13g2_dfrbp_1 \logix.ram_r[380]$_DFFE_PP_  (.CLK(net744),
    .RESET_B(net2165),
    .D(_1374_),
    .Q_N(_4624_),
    .Q(\logix.ram_r[380] ));
 sg13g2_dfrbp_1 \logix.ram_r[381]$_DFFE_PP_  (.CLK(net739),
    .RESET_B(net2166),
    .D(_1375_),
    .Q_N(_4623_),
    .Q(\logix.ram_r[381] ));
 sg13g2_dfrbp_1 \logix.ram_r[382]$_DFFE_PP_  (.CLK(net676),
    .RESET_B(net2167),
    .D(_1376_),
    .Q_N(_4622_),
    .Q(\logix.ram_r[382] ));
 sg13g2_dfrbp_1 \logix.ram_r[383]$_DFFE_PP_  (.CLK(net673),
    .RESET_B(net2168),
    .D(_1377_),
    .Q_N(_4621_),
    .Q(\logix.ram_r[383] ));
 sg13g2_dfrbp_1 \logix.ram_r[384]$_DFFE_PP_  (.CLK(net570),
    .RESET_B(net2169),
    .D(_1378_),
    .Q_N(_4620_),
    .Q(\logix.ram_r[384] ));
 sg13g2_dfrbp_1 \logix.ram_r[385]$_DFFE_PP_  (.CLK(net555),
    .RESET_B(net2170),
    .D(_1379_),
    .Q_N(_4619_),
    .Q(\logix.ram_r[385] ));
 sg13g2_dfrbp_1 \logix.ram_r[386]$_DFFE_PP_  (.CLK(net556),
    .RESET_B(net2171),
    .D(_1380_),
    .Q_N(_4618_),
    .Q(\logix.ram_r[386] ));
 sg13g2_dfrbp_1 \logix.ram_r[387]$_DFFE_PP_  (.CLK(net555),
    .RESET_B(net2172),
    .D(_1381_),
    .Q_N(_4617_),
    .Q(\logix.ram_r[387] ));
 sg13g2_dfrbp_1 \logix.ram_r[388]$_DFFE_PP_  (.CLK(net551),
    .RESET_B(net2173),
    .D(_1382_),
    .Q_N(_4616_),
    .Q(\logix.ram_r[388] ));
 sg13g2_dfrbp_1 \logix.ram_r[389]$_DFFE_PP_  (.CLK(net550),
    .RESET_B(net2174),
    .D(_1383_),
    .Q_N(_4615_),
    .Q(\logix.ram_r[389] ));
 sg13g2_dfrbp_1 \logix.ram_r[38]$_DFFE_PP_  (.CLK(net639),
    .RESET_B(net2175),
    .D(_1384_),
    .Q_N(_4614_),
    .Q(\logix.ram_r[38] ));
 sg13g2_dfrbp_1 \logix.ram_r[390]$_DFFE_PP_  (.CLK(net550),
    .RESET_B(net2176),
    .D(_1385_),
    .Q_N(_4613_),
    .Q(\logix.ram_r[390] ));
 sg13g2_dfrbp_1 \logix.ram_r[391]$_DFFE_PP_  (.CLK(net520),
    .RESET_B(net2177),
    .D(_1386_),
    .Q_N(_4612_),
    .Q(\logix.ram_r[391] ));
 sg13g2_dfrbp_1 \logix.ram_r[392]$_DFFE_PP_  (.CLK(net555),
    .RESET_B(net2178),
    .D(_1387_),
    .Q_N(_4611_),
    .Q(\logix.ram_r[392] ));
 sg13g2_dfrbp_1 \logix.ram_r[393]$_DFFE_PP_  (.CLK(net556),
    .RESET_B(net2179),
    .D(_1388_),
    .Q_N(_4610_),
    .Q(\logix.ram_r[393] ));
 sg13g2_dfrbp_1 \logix.ram_r[394]$_DFFE_PP_  (.CLK(net556),
    .RESET_B(net2180),
    .D(_1389_),
    .Q_N(_4609_),
    .Q(\logix.ram_r[394] ));
 sg13g2_dfrbp_1 \logix.ram_r[395]$_DFFE_PP_  (.CLK(net555),
    .RESET_B(net2181),
    .D(_1390_),
    .Q_N(_4608_),
    .Q(\logix.ram_r[395] ));
 sg13g2_dfrbp_1 \logix.ram_r[396]$_DFFE_PP_  (.CLK(net551),
    .RESET_B(net2182),
    .D(_1391_),
    .Q_N(_4607_),
    .Q(\logix.ram_r[396] ));
 sg13g2_dfrbp_1 \logix.ram_r[397]$_DFFE_PP_  (.CLK(net550),
    .RESET_B(net2183),
    .D(_1392_),
    .Q_N(_4606_),
    .Q(\logix.ram_r[397] ));
 sg13g2_dfrbp_1 \logix.ram_r[398]$_DFFE_PP_  (.CLK(net551),
    .RESET_B(net2184),
    .D(_1393_),
    .Q_N(_4605_),
    .Q(\logix.ram_r[398] ));
 sg13g2_dfrbp_1 \logix.ram_r[399]$_DFFE_PP_  (.CLK(net555),
    .RESET_B(net2185),
    .D(_1394_),
    .Q_N(_4604_),
    .Q(\logix.ram_r[399] ));
 sg13g2_dfrbp_1 \logix.ram_r[39]$_DFFE_PP_  (.CLK(net639),
    .RESET_B(net2186),
    .D(_1395_),
    .Q_N(_4603_),
    .Q(\logix.ram_r[39] ));
 sg13g2_dfrbp_1 \logix.ram_r[3]$_DFFE_PP_  (.CLK(net640),
    .RESET_B(net2187),
    .D(_1396_),
    .Q_N(_4602_),
    .Q(\logix.ram_r[3] ));
 sg13g2_dfrbp_1 \logix.ram_r[400]$_DFFE_PP_  (.CLK(net555),
    .RESET_B(net2188),
    .D(_1397_),
    .Q_N(_4601_),
    .Q(\logix.ram_r[400] ));
 sg13g2_dfrbp_1 \logix.ram_r[401]$_DFFE_PP_  (.CLK(net555),
    .RESET_B(net2189),
    .D(_1398_),
    .Q_N(_4600_),
    .Q(\logix.ram_r[401] ));
 sg13g2_dfrbp_1 \logix.ram_r[402]$_DFFE_PP_  (.CLK(net556),
    .RESET_B(net2190),
    .D(_1399_),
    .Q_N(_4599_),
    .Q(\logix.ram_r[402] ));
 sg13g2_dfrbp_1 \logix.ram_r[403]$_DFFE_PP_  (.CLK(net555),
    .RESET_B(net2191),
    .D(_1400_),
    .Q_N(_4598_),
    .Q(\logix.ram_r[403] ));
 sg13g2_dfrbp_1 \logix.ram_r[404]$_DFFE_PP_  (.CLK(net551),
    .RESET_B(net2192),
    .D(_1401_),
    .Q_N(_4597_),
    .Q(\logix.ram_r[404] ));
 sg13g2_dfrbp_1 \logix.ram_r[405]$_DFFE_PP_  (.CLK(net551),
    .RESET_B(net2193),
    .D(_1402_),
    .Q_N(_4596_),
    .Q(\logix.ram_r[405] ));
 sg13g2_dfrbp_1 \logix.ram_r[406]$_DFFE_PP_  (.CLK(net520),
    .RESET_B(net2194),
    .D(_1403_),
    .Q_N(_4595_),
    .Q(\logix.ram_r[406] ));
 sg13g2_dfrbp_1 \logix.ram_r[407]$_DFFE_PP_  (.CLK(net525),
    .RESET_B(net2195),
    .D(_1404_),
    .Q_N(_4594_),
    .Q(\logix.ram_r[407] ));
 sg13g2_dfrbp_1 \logix.ram_r[408]$_DFFE_PP_  (.CLK(net556),
    .RESET_B(net2196),
    .D(_1405_),
    .Q_N(_4593_),
    .Q(\logix.ram_r[408] ));
 sg13g2_dfrbp_1 \logix.ram_r[409]$_DFFE_PP_  (.CLK(net556),
    .RESET_B(net2197),
    .D(_1406_),
    .Q_N(_4592_),
    .Q(\logix.ram_r[409] ));
 sg13g2_dfrbp_1 \logix.ram_r[40]$_DFFE_PP_  (.CLK(net634),
    .RESET_B(net2198),
    .D(_1407_),
    .Q_N(_4591_),
    .Q(\logix.ram_r[40] ));
 sg13g2_dfrbp_1 \logix.ram_r[410]$_DFFE_PP_  (.CLK(net558),
    .RESET_B(net2199),
    .D(_1408_),
    .Q_N(_4590_),
    .Q(\logix.ram_r[410] ));
 sg13g2_dfrbp_1 \logix.ram_r[411]$_DFFE_PP_  (.CLK(net556),
    .RESET_B(net2200),
    .D(_1409_),
    .Q_N(_4589_),
    .Q(\logix.ram_r[411] ));
 sg13g2_dfrbp_1 \logix.ram_r[412]$_DFFE_PP_  (.CLK(net551),
    .RESET_B(net2201),
    .D(_1410_),
    .Q_N(_4588_),
    .Q(\logix.ram_r[412] ));
 sg13g2_dfrbp_1 \logix.ram_r[413]$_DFFE_PP_  (.CLK(net554),
    .RESET_B(net2202),
    .D(_1411_),
    .Q_N(_4587_),
    .Q(\logix.ram_r[413] ));
 sg13g2_dfrbp_1 \logix.ram_r[414]$_DFFE_PP_  (.CLK(net520),
    .RESET_B(net2203),
    .D(_1412_),
    .Q_N(_4586_),
    .Q(\logix.ram_r[414] ));
 sg13g2_dfrbp_1 \logix.ram_r[415]$_DFFE_PP_  (.CLK(net522),
    .RESET_B(net2204),
    .D(_1413_),
    .Q_N(_4585_),
    .Q(\logix.ram_r[415] ));
 sg13g2_dfrbp_1 \logix.ram_r[416]$_DFFE_PP_  (.CLK(net520),
    .RESET_B(net2205),
    .D(_1414_),
    .Q_N(_4584_),
    .Q(\logix.ram_r[416] ));
 sg13g2_dfrbp_1 \logix.ram_r[417]$_DFFE_PP_  (.CLK(net520),
    .RESET_B(net2206),
    .D(_1415_),
    .Q_N(_4583_),
    .Q(\logix.ram_r[417] ));
 sg13g2_dfrbp_1 \logix.ram_r[418]$_DFFE_PP_  (.CLK(net520),
    .RESET_B(net2207),
    .D(_1416_),
    .Q_N(_4582_),
    .Q(\logix.ram_r[418] ));
 sg13g2_dfrbp_1 \logix.ram_r[419]$_DFFE_PP_  (.CLK(net525),
    .RESET_B(net2208),
    .D(_1417_),
    .Q_N(_4581_),
    .Q(\logix.ram_r[419] ));
 sg13g2_dfrbp_1 \logix.ram_r[41]$_DFFE_PP_  (.CLK(net634),
    .RESET_B(net2209),
    .D(_1418_),
    .Q_N(_4580_),
    .Q(\logix.ram_r[41] ));
 sg13g2_dfrbp_1 \logix.ram_r[420]$_DFFE_PP_  (.CLK(net538),
    .RESET_B(net2210),
    .D(_1419_),
    .Q_N(_4579_),
    .Q(\logix.ram_r[420] ));
 sg13g2_dfrbp_1 \logix.ram_r[421]$_DFFE_PP_  (.CLK(net538),
    .RESET_B(net2211),
    .D(_1420_),
    .Q_N(_4578_),
    .Q(\logix.ram_r[421] ));
 sg13g2_dfrbp_1 \logix.ram_r[422]$_DFFE_PP_  (.CLK(net538),
    .RESET_B(net2212),
    .D(_1421_),
    .Q_N(_4577_),
    .Q(\logix.ram_r[422] ));
 sg13g2_dfrbp_1 \logix.ram_r[423]$_DFFE_PP_  (.CLK(net524),
    .RESET_B(net2213),
    .D(_1422_),
    .Q_N(_4576_),
    .Q(\logix.ram_r[423] ));
 sg13g2_dfrbp_1 \logix.ram_r[424]$_DFFE_PP_  (.CLK(net523),
    .RESET_B(net2214),
    .D(_1423_),
    .Q_N(_4575_),
    .Q(\logix.ram_r[424] ));
 sg13g2_dfrbp_1 \logix.ram_r[425]$_DFFE_PP_  (.CLK(net523),
    .RESET_B(net2215),
    .D(_1424_),
    .Q_N(_4574_),
    .Q(\logix.ram_r[425] ));
 sg13g2_dfrbp_1 \logix.ram_r[426]$_DFFE_PP_  (.CLK(net525),
    .RESET_B(net2216),
    .D(_1425_),
    .Q_N(_4573_),
    .Q(\logix.ram_r[426] ));
 sg13g2_dfrbp_1 \logix.ram_r[427]$_DFFE_PP_  (.CLK(net525),
    .RESET_B(net2217),
    .D(_1426_),
    .Q_N(_4572_),
    .Q(\logix.ram_r[427] ));
 sg13g2_dfrbp_1 \logix.ram_r[428]$_DFFE_PP_  (.CLK(net525),
    .RESET_B(net2218),
    .D(_1427_),
    .Q_N(_4571_),
    .Q(\logix.ram_r[428] ));
 sg13g2_dfrbp_1 \logix.ram_r[429]$_DFFE_PP_  (.CLK(net526),
    .RESET_B(net2219),
    .D(_1428_),
    .Q_N(_4570_),
    .Q(\logix.ram_r[429] ));
 sg13g2_dfrbp_1 \logix.ram_r[42]$_DFFE_PP_  (.CLK(net604),
    .RESET_B(net2220),
    .D(_1429_),
    .Q_N(_4569_),
    .Q(\logix.ram_r[42] ));
 sg13g2_dfrbp_1 \logix.ram_r[430]$_DFFE_PP_  (.CLK(net526),
    .RESET_B(net2221),
    .D(_1430_),
    .Q_N(_4568_),
    .Q(\logix.ram_r[430] ));
 sg13g2_dfrbp_1 \logix.ram_r[431]$_DFFE_PP_  (.CLK(net525),
    .RESET_B(net2222),
    .D(_1431_),
    .Q_N(_4567_),
    .Q(\logix.ram_r[431] ));
 sg13g2_dfrbp_1 \logix.ram_r[432]$_DFFE_PP_  (.CLK(net525),
    .RESET_B(net2223),
    .D(_1432_),
    .Q_N(_4566_),
    .Q(\logix.ram_r[432] ));
 sg13g2_dfrbp_1 \logix.ram_r[433]$_DFFE_PP_  (.CLK(net525),
    .RESET_B(net2224),
    .D(_1433_),
    .Q_N(_4565_),
    .Q(\logix.ram_r[433] ));
 sg13g2_dfrbp_1 \logix.ram_r[434]$_DFFE_PP_  (.CLK(net526),
    .RESET_B(net2225),
    .D(_1434_),
    .Q_N(_4564_),
    .Q(\logix.ram_r[434] ));
 sg13g2_dfrbp_1 \logix.ram_r[435]$_DFFE_PP_  (.CLK(net540),
    .RESET_B(net2226),
    .D(_1435_),
    .Q_N(_4563_),
    .Q(\logix.ram_r[435] ));
 sg13g2_dfrbp_1 \logix.ram_r[436]$_DFFE_PP_  (.CLK(net540),
    .RESET_B(net2227),
    .D(_1436_),
    .Q_N(_4562_),
    .Q(\logix.ram_r[436] ));
 sg13g2_dfrbp_1 \logix.ram_r[437]$_DFFE_PP_  (.CLK(net539),
    .RESET_B(net2228),
    .D(_1437_),
    .Q_N(_4561_),
    .Q(\logix.ram_r[437] ));
 sg13g2_dfrbp_1 \logix.ram_r[438]$_DFFE_PP_  (.CLK(net539),
    .RESET_B(net2229),
    .D(_1438_),
    .Q_N(_4560_),
    .Q(\logix.ram_r[438] ));
 sg13g2_dfrbp_1 \logix.ram_r[439]$_DFFE_PP_  (.CLK(net524),
    .RESET_B(net2230),
    .D(_1439_),
    .Q_N(_4559_),
    .Q(\logix.ram_r[439] ));
 sg13g2_dfrbp_1 \logix.ram_r[43]$_DFFE_PP_  (.CLK(net541),
    .RESET_B(net2231),
    .D(_1440_),
    .Q_N(_4558_),
    .Q(\logix.ram_r[43] ));
 sg13g2_dfrbp_1 \logix.ram_r[440]$_DFFE_PP_  (.CLK(net524),
    .RESET_B(net2232),
    .D(_1441_),
    .Q_N(_4557_),
    .Q(\logix.ram_r[440] ));
 sg13g2_dfrbp_1 \logix.ram_r[441]$_DFFE_PP_  (.CLK(net524),
    .RESET_B(net2233),
    .D(_1442_),
    .Q_N(_4556_),
    .Q(\logix.ram_r[441] ));
 sg13g2_dfrbp_1 \logix.ram_r[442]$_DFFE_PP_  (.CLK(net526),
    .RESET_B(net2234),
    .D(_1443_),
    .Q_N(_4555_),
    .Q(\logix.ram_r[442] ));
 sg13g2_dfrbp_1 \logix.ram_r[443]$_DFFE_PP_  (.CLK(net540),
    .RESET_B(net2235),
    .D(_1444_),
    .Q_N(_4554_),
    .Q(\logix.ram_r[443] ));
 sg13g2_dfrbp_1 \logix.ram_r[444]$_DFFE_PP_  (.CLK(net540),
    .RESET_B(net2236),
    .D(_1445_),
    .Q_N(_4553_),
    .Q(\logix.ram_r[444] ));
 sg13g2_dfrbp_1 \logix.ram_r[445]$_DFFE_PP_  (.CLK(net540),
    .RESET_B(net2237),
    .D(_1446_),
    .Q_N(_4552_),
    .Q(\logix.ram_r[445] ));
 sg13g2_dfrbp_1 \logix.ram_r[446]$_DFFE_PP_  (.CLK(net570),
    .RESET_B(net2238),
    .D(_1447_),
    .Q_N(_4551_),
    .Q(\logix.ram_r[446] ));
 sg13g2_dfrbp_1 \logix.ram_r[447]$_DFFE_PP_  (.CLK(net558),
    .RESET_B(net2239),
    .D(_1448_),
    .Q_N(_4550_),
    .Q(\logix.ram_r[447] ));
 sg13g2_dfrbp_1 \logix.ram_r[448]$_DFFE_PP_  (.CLK(net557),
    .RESET_B(net2240),
    .D(_1449_),
    .Q_N(_4549_),
    .Q(\logix.ram_r[448] ));
 sg13g2_dfrbp_1 \logix.ram_r[449]$_DFFE_PP_  (.CLK(net557),
    .RESET_B(net2241),
    .D(_1450_),
    .Q_N(_4548_),
    .Q(\logix.ram_r[449] ));
 sg13g2_dfrbp_1 \logix.ram_r[44]$_DFFE_PP_  (.CLK(net571),
    .RESET_B(net2242),
    .D(_1451_),
    .Q_N(_4547_),
    .Q(\logix.ram_r[44] ));
 sg13g2_dfrbp_1 \logix.ram_r[450]$_DFFE_PP_  (.CLK(net557),
    .RESET_B(net2243),
    .D(_1452_),
    .Q_N(_4546_),
    .Q(\logix.ram_r[450] ));
 sg13g2_dfrbp_1 \logix.ram_r[451]$_DFFE_PP_  (.CLK(net572),
    .RESET_B(net2244),
    .D(_1453_),
    .Q_N(_4545_),
    .Q(\logix.ram_r[451] ));
 sg13g2_dfrbp_1 \logix.ram_r[452]$_DFFE_PP_  (.CLK(net572),
    .RESET_B(net2245),
    .D(_1454_),
    .Q_N(_4544_),
    .Q(\logix.ram_r[452] ));
 sg13g2_dfrbp_1 \logix.ram_r[453]$_DFFE_PP_  (.CLK(net572),
    .RESET_B(net2246),
    .D(_1455_),
    .Q_N(_4543_),
    .Q(\logix.ram_r[453] ));
 sg13g2_dfrbp_1 \logix.ram_r[454]$_DFFE_PP_  (.CLK(net572),
    .RESET_B(net2247),
    .D(_1456_),
    .Q_N(_4542_),
    .Q(\logix.ram_r[454] ));
 sg13g2_dfrbp_1 \logix.ram_r[455]$_DFFE_PP_  (.CLK(net557),
    .RESET_B(net2248),
    .D(_1457_),
    .Q_N(_4541_),
    .Q(\logix.ram_r[455] ));
 sg13g2_dfrbp_1 \logix.ram_r[456]$_DFFE_PP_  (.CLK(net557),
    .RESET_B(net2249),
    .D(_1458_),
    .Q_N(_4540_),
    .Q(\logix.ram_r[456] ));
 sg13g2_dfrbp_1 \logix.ram_r[457]$_DFFE_PP_  (.CLK(net557),
    .RESET_B(net2250),
    .D(_1459_),
    .Q_N(_4539_),
    .Q(\logix.ram_r[457] ));
 sg13g2_dfrbp_1 \logix.ram_r[458]$_DFFE_PP_  (.CLK(net557),
    .RESET_B(net2251),
    .D(_1460_),
    .Q_N(_4538_),
    .Q(\logix.ram_r[458] ));
 sg13g2_dfrbp_1 \logix.ram_r[459]$_DFFE_PP_  (.CLK(net558),
    .RESET_B(net2252),
    .D(_1461_),
    .Q_N(_4537_),
    .Q(\logix.ram_r[459] ));
 sg13g2_dfrbp_1 \logix.ram_r[45]$_DFFE_PP_  (.CLK(net570),
    .RESET_B(net2253),
    .D(_1462_),
    .Q_N(_4536_),
    .Q(\logix.ram_r[45] ));
 sg13g2_dfrbp_1 \logix.ram_r[460]$_DFFE_PP_  (.CLK(net572),
    .RESET_B(net2254),
    .D(_1463_),
    .Q_N(_4535_),
    .Q(\logix.ram_r[460] ));
 sg13g2_dfrbp_1 \logix.ram_r[461]$_DFFE_PP_  (.CLK(net572),
    .RESET_B(net2255),
    .D(_1464_),
    .Q_N(_4534_),
    .Q(\logix.ram_r[461] ));
 sg13g2_dfrbp_1 \logix.ram_r[462]$_DFFE_PP_  (.CLK(net572),
    .RESET_B(net2256),
    .D(_1465_),
    .Q_N(_4533_),
    .Q(\logix.ram_r[462] ));
 sg13g2_dfrbp_1 \logix.ram_r[463]$_DFFE_PP_  (.CLK(net554),
    .RESET_B(net2257),
    .D(_1466_),
    .Q_N(_4532_),
    .Q(\logix.ram_r[463] ));
 sg13g2_dfrbp_1 \logix.ram_r[464]$_DFFE_PP_  (.CLK(net554),
    .RESET_B(net2258),
    .D(_1467_),
    .Q_N(_4531_),
    .Q(\logix.ram_r[464] ));
 sg13g2_dfrbp_1 \logix.ram_r[465]$_DFFE_PP_  (.CLK(net496),
    .RESET_B(net2259),
    .D(_1468_),
    .Q_N(_4530_),
    .Q(\logix.ram_r[465] ));
 sg13g2_dfrbp_1 \logix.ram_r[466]$_DFFE_PP_  (.CLK(net496),
    .RESET_B(net2260),
    .D(_1469_),
    .Q_N(_4529_),
    .Q(\logix.ram_r[466] ));
 sg13g2_dfrbp_1 \logix.ram_r[467]$_DFFE_PP_  (.CLK(net500),
    .RESET_B(net2261),
    .D(_1470_),
    .Q_N(_4528_),
    .Q(\logix.ram_r[467] ));
 sg13g2_dfrbp_1 \logix.ram_r[468]$_DFFE_PP_  (.CLK(net500),
    .RESET_B(net2262),
    .D(_1471_),
    .Q_N(_4527_),
    .Q(\logix.ram_r[468] ));
 sg13g2_dfrbp_1 \logix.ram_r[469]$_DFFE_PP_  (.CLK(net501),
    .RESET_B(net2263),
    .D(_1472_),
    .Q_N(_4526_),
    .Q(\logix.ram_r[469] ));
 sg13g2_dfrbp_1 \logix.ram_r[46]$_DFFE_PP_  (.CLK(net570),
    .RESET_B(net2264),
    .D(_1473_),
    .Q_N(_4525_),
    .Q(\logix.ram_r[46] ));
 sg13g2_dfrbp_1 \logix.ram_r[470]$_DFFE_PP_  (.CLK(net501),
    .RESET_B(net2265),
    .D(_1474_),
    .Q_N(_4524_),
    .Q(\logix.ram_r[470] ));
 sg13g2_dfrbp_1 \logix.ram_r[471]$_DFFE_PP_  (.CLK(net501),
    .RESET_B(net2266),
    .D(_1475_),
    .Q_N(_4523_),
    .Q(\logix.ram_r[471] ));
 sg13g2_dfrbp_1 \logix.ram_r[472]$_DFFE_PP_  (.CLK(net496),
    .RESET_B(net2267),
    .D(_1476_),
    .Q_N(_4522_),
    .Q(\logix.ram_r[472] ));
 sg13g2_dfrbp_1 \logix.ram_r[473]$_DFFE_PP_  (.CLK(net496),
    .RESET_B(net2268),
    .D(_1477_),
    .Q_N(_4521_),
    .Q(\logix.ram_r[473] ));
 sg13g2_dfrbp_1 \logix.ram_r[474]$_DFFE_PP_  (.CLK(net496),
    .RESET_B(net2269),
    .D(_1478_),
    .Q_N(_4520_),
    .Q(\logix.ram_r[474] ));
 sg13g2_dfrbp_1 \logix.ram_r[475]$_DFFE_PP_  (.CLK(net500),
    .RESET_B(net2270),
    .D(_1479_),
    .Q_N(_4519_),
    .Q(\logix.ram_r[475] ));
 sg13g2_dfrbp_1 \logix.ram_r[476]$_DFFE_PP_  (.CLK(net500),
    .RESET_B(net2271),
    .D(_1480_),
    .Q_N(_4518_),
    .Q(\logix.ram_r[476] ));
 sg13g2_dfrbp_1 \logix.ram_r[477]$_DFFE_PP_  (.CLK(net502),
    .RESET_B(net2272),
    .D(_1481_),
    .Q_N(_4517_),
    .Q(\logix.ram_r[477] ));
 sg13g2_dfrbp_1 \logix.ram_r[478]$_DFFE_PP_  (.CLK(net501),
    .RESET_B(net2273),
    .D(_1482_),
    .Q_N(_4516_),
    .Q(\logix.ram_r[478] ));
 sg13g2_dfrbp_1 \logix.ram_r[479]$_DFFE_PP_  (.CLK(net502),
    .RESET_B(net2274),
    .D(_1483_),
    .Q_N(_4515_),
    .Q(\logix.ram_r[479] ));
 sg13g2_dfrbp_1 \logix.ram_r[47]$_DFFE_PP_  (.CLK(net570),
    .RESET_B(net2275),
    .D(_1484_),
    .Q_N(_4514_),
    .Q(\logix.ram_r[47] ));
 sg13g2_dfrbp_1 \logix.ram_r[480]$_DFFE_PP_  (.CLK(net497),
    .RESET_B(net2276),
    .D(_1485_),
    .Q_N(_4513_),
    .Q(\logix.ram_r[480] ));
 sg13g2_dfrbp_1 \logix.ram_r[481]$_DFFE_PP_  (.CLK(net497),
    .RESET_B(net2277),
    .D(_1486_),
    .Q_N(_4512_),
    .Q(\logix.ram_r[481] ));
 sg13g2_dfrbp_1 \logix.ram_r[482]$_DFFE_PP_  (.CLK(net498),
    .RESET_B(net2278),
    .D(_1487_),
    .Q_N(_4511_),
    .Q(\logix.ram_r[482] ));
 sg13g2_dfrbp_1 \logix.ram_r[483]$_DFFE_PP_  (.CLK(net504),
    .RESET_B(net2279),
    .D(_1488_),
    .Q_N(_4510_),
    .Q(\logix.ram_r[483] ));
 sg13g2_dfrbp_1 \logix.ram_r[484]$_DFFE_PP_  (.CLK(net504),
    .RESET_B(net2280),
    .D(_1489_),
    .Q_N(_4509_),
    .Q(\logix.ram_r[484] ));
 sg13g2_dfrbp_1 \logix.ram_r[485]$_DFFE_PP_  (.CLK(net503),
    .RESET_B(net2281),
    .D(_1490_),
    .Q_N(_4508_),
    .Q(\logix.ram_r[485] ));
 sg13g2_dfrbp_1 \logix.ram_r[486]$_DFFE_PP_  (.CLK(net503),
    .RESET_B(net2282),
    .D(_1491_),
    .Q_N(_4507_),
    .Q(\logix.ram_r[486] ));
 sg13g2_dfrbp_1 \logix.ram_r[487]$_DFFE_PP_  (.CLK(net503),
    .RESET_B(net2283),
    .D(_1492_),
    .Q_N(_4506_),
    .Q(\logix.ram_r[487] ));
 sg13g2_dfrbp_1 \logix.ram_r[488]$_DFFE_PP_  (.CLK(net498),
    .RESET_B(net2284),
    .D(_1493_),
    .Q_N(_4505_),
    .Q(\logix.ram_r[488] ));
 sg13g2_dfrbp_1 \logix.ram_r[489]$_DFFE_PP_  (.CLK(net498),
    .RESET_B(net2285),
    .D(_1494_),
    .Q_N(_4504_),
    .Q(\logix.ram_r[489] ));
 sg13g2_dfrbp_1 \logix.ram_r[48]$_DFFE_PP_  (.CLK(net570),
    .RESET_B(net2286),
    .D(_1495_),
    .Q_N(_4503_),
    .Q(\logix.ram_r[48] ));
 sg13g2_dfrbp_1 \logix.ram_r[490]$_DFFE_PP_  (.CLK(net498),
    .RESET_B(net2287),
    .D(_1496_),
    .Q_N(_4502_),
    .Q(\logix.ram_r[490] ));
 sg13g2_dfrbp_1 \logix.ram_r[491]$_DFFE_PP_  (.CLK(net504),
    .RESET_B(net2288),
    .D(_1497_),
    .Q_N(_4501_),
    .Q(\logix.ram_r[491] ));
 sg13g2_dfrbp_1 \logix.ram_r[492]$_DFFE_PP_  (.CLK(net504),
    .RESET_B(net2289),
    .D(_1498_),
    .Q_N(_4500_),
    .Q(\logix.ram_r[492] ));
 sg13g2_dfrbp_1 \logix.ram_r[493]$_DFFE_PP_  (.CLK(net503),
    .RESET_B(net2290),
    .D(_1499_),
    .Q_N(_4499_),
    .Q(\logix.ram_r[493] ));
 sg13g2_dfrbp_1 \logix.ram_r[494]$_DFFE_PP_  (.CLK(net503),
    .RESET_B(net2291),
    .D(_1500_),
    .Q_N(_4498_),
    .Q(\logix.ram_r[494] ));
 sg13g2_dfrbp_1 \logix.ram_r[495]$_DFFE_PP_  (.CLK(net503),
    .RESET_B(net2292),
    .D(_1501_),
    .Q_N(_4497_),
    .Q(\logix.ram_r[495] ));
 sg13g2_dfrbp_1 \logix.ram_r[496]$_DFFE_PP_  (.CLK(net562),
    .RESET_B(net2293),
    .D(_1502_),
    .Q_N(_4496_),
    .Q(\logix.ram_r[496] ));
 sg13g2_dfrbp_1 \logix.ram_r[497]$_DFFE_PP_  (.CLK(net565),
    .RESET_B(net2294),
    .D(_1503_),
    .Q_N(_4495_),
    .Q(\logix.ram_r[497] ));
 sg13g2_dfrbp_1 \logix.ram_r[498]$_DFFE_PP_  (.CLK(net565),
    .RESET_B(net2295),
    .D(_1504_),
    .Q_N(_4494_),
    .Q(\logix.ram_r[498] ));
 sg13g2_dfrbp_1 \logix.ram_r[499]$_DFFE_PP_  (.CLK(net580),
    .RESET_B(net2296),
    .D(_1505_),
    .Q_N(_4493_),
    .Q(\logix.ram_r[499] ));
 sg13g2_dfrbp_1 \logix.ram_r[49]$_DFFE_PP_  (.CLK(net571),
    .RESET_B(net2297),
    .D(_1506_),
    .Q_N(_4492_),
    .Q(\logix.ram_r[49] ));
 sg13g2_dfrbp_1 \logix.ram_r[4]$_DFFE_PP_  (.CLK(net639),
    .RESET_B(net2298),
    .D(_1507_),
    .Q_N(_4491_),
    .Q(\logix.ram_r[4] ));
 sg13g2_dfrbp_1 \logix.ram_r[500]$_DFFE_PP_  (.CLK(net580),
    .RESET_B(net2299),
    .D(_1508_),
    .Q_N(_4490_),
    .Q(\logix.ram_r[500] ));
 sg13g2_dfrbp_1 \logix.ram_r[501]$_DFFE_PP_  (.CLK(net581),
    .RESET_B(net2300),
    .D(_1509_),
    .Q_N(_4489_),
    .Q(\logix.ram_r[501] ));
 sg13g2_dfrbp_1 \logix.ram_r[502]$_DFFE_PP_  (.CLK(net572),
    .RESET_B(net2301),
    .D(_1510_),
    .Q_N(_4488_),
    .Q(\logix.ram_r[502] ));
 sg13g2_dfrbp_1 \logix.ram_r[503]$_DFFE_PP_  (.CLK(net573),
    .RESET_B(net2302),
    .D(_1511_),
    .Q_N(_4487_),
    .Q(\logix.ram_r[503] ));
 sg13g2_dfrbp_1 \logix.ram_r[504]$_DFFE_PP_  (.CLK(net558),
    .RESET_B(net2303),
    .D(_1512_),
    .Q_N(_4486_),
    .Q(\logix.ram_r[504] ));
 sg13g2_dfrbp_1 \logix.ram_r[505]$_DFFE_PP_  (.CLK(net558),
    .RESET_B(net2304),
    .D(_1513_),
    .Q_N(_4485_),
    .Q(\logix.ram_r[505] ));
 sg13g2_dfrbp_1 \logix.ram_r[506]$_DFFE_PP_  (.CLK(net565),
    .RESET_B(net2305),
    .D(_1514_),
    .Q_N(_4484_),
    .Q(\logix.ram_r[506] ));
 sg13g2_dfrbp_1 \logix.ram_r[507]$_DFFE_PP_  (.CLK(net580),
    .RESET_B(net2306),
    .D(_1515_),
    .Q_N(_4483_),
    .Q(\logix.ram_r[507] ));
 sg13g2_dfrbp_1 \logix.ram_r[508]$_DFFE_PP_  (.CLK(net580),
    .RESET_B(net2307),
    .D(_1516_),
    .Q_N(_4482_),
    .Q(\logix.ram_r[508] ));
 sg13g2_dfrbp_1 \logix.ram_r[509]$_DFFE_PP_  (.CLK(net573),
    .RESET_B(net2308),
    .D(_1517_),
    .Q_N(_4481_),
    .Q(\logix.ram_r[509] ));
 sg13g2_dfrbp_1 \logix.ram_r[50]$_DFFE_PP_  (.CLK(net657),
    .RESET_B(net2309),
    .D(_1518_),
    .Q_N(_4480_),
    .Q(\logix.ram_r[50] ));
 sg13g2_dfrbp_1 \logix.ram_r[510]$_DFFE_PP_  (.CLK(net573),
    .RESET_B(net2310),
    .D(_1519_),
    .Q_N(_4479_),
    .Q(\logix.ram_r[510] ));
 sg13g2_dfrbp_1 \logix.ram_r[511]$_DFFE_PP_  (.CLK(net573),
    .RESET_B(net2311),
    .D(_1520_),
    .Q_N(_4478_),
    .Q(\logix.ram_r[511] ));
 sg13g2_dfrbp_1 \logix.ram_r[512]$_DFFE_PP_  (.CLK(net728),
    .RESET_B(net2312),
    .D(_1521_),
    .Q_N(_4477_),
    .Q(\logix.ram_r[512] ));
 sg13g2_dfrbp_1 \logix.ram_r[513]$_DFFE_PP_  (.CLK(net728),
    .RESET_B(net2313),
    .D(_1522_),
    .Q_N(_4476_),
    .Q(\logix.ram_r[513] ));
 sg13g2_dfrbp_1 \logix.ram_r[514]$_DFFE_PP_  (.CLK(net728),
    .RESET_B(net2314),
    .D(_1523_),
    .Q_N(_4475_),
    .Q(\logix.ram_r[514] ));
 sg13g2_dfrbp_1 \logix.ram_r[515]$_DFFE_PP_  (.CLK(net734),
    .RESET_B(net2315),
    .D(_1524_),
    .Q_N(_4474_),
    .Q(\logix.ram_r[515] ));
 sg13g2_dfrbp_1 \logix.ram_r[516]$_DFFE_PP_  (.CLK(net726),
    .RESET_B(net2316),
    .D(_1525_),
    .Q_N(_4473_),
    .Q(\logix.ram_r[516] ));
 sg13g2_dfrbp_1 \logix.ram_r[517]$_DFFE_PP_  (.CLK(net731),
    .RESET_B(net2317),
    .D(_1526_),
    .Q_N(_4472_),
    .Q(\logix.ram_r[517] ));
 sg13g2_dfrbp_1 \logix.ram_r[518]$_DFFE_PP_  (.CLK(net699),
    .RESET_B(net2318),
    .D(_1527_),
    .Q_N(_4471_),
    .Q(\logix.ram_r[518] ));
 sg13g2_dfrbp_1 \logix.ram_r[519]$_DFFE_PP_  (.CLK(net694),
    .RESET_B(net2319),
    .D(_1528_),
    .Q_N(_4470_),
    .Q(\logix.ram_r[519] ));
 sg13g2_dfrbp_1 \logix.ram_r[51]$_DFFE_PP_  (.CLK(net625),
    .RESET_B(net2320),
    .D(_1529_),
    .Q_N(_4469_),
    .Q(\logix.ram_r[51] ));
 sg13g2_dfrbp_1 \logix.ram_r[520]$_DFFE_PP_  (.CLK(net727),
    .RESET_B(net2321),
    .D(_1530_),
    .Q_N(_4468_),
    .Q(\logix.ram_r[520] ));
 sg13g2_dfrbp_1 \logix.ram_r[521]$_DFFE_PP_  (.CLK(net726),
    .RESET_B(net2322),
    .D(_1531_),
    .Q_N(_4467_),
    .Q(\logix.ram_r[521] ));
 sg13g2_dfrbp_1 \logix.ram_r[522]$_DFFE_PP_  (.CLK(net726),
    .RESET_B(net2323),
    .D(_1532_),
    .Q_N(_4466_),
    .Q(\logix.ram_r[522] ));
 sg13g2_dfrbp_1 \logix.ram_r[523]$_DFFE_PP_  (.CLK(net731),
    .RESET_B(net2324),
    .D(_1533_),
    .Q_N(_4465_),
    .Q(\logix.ram_r[523] ));
 sg13g2_dfrbp_1 \logix.ram_r[524]$_DFFE_PP_  (.CLK(net726),
    .RESET_B(net2325),
    .D(_1534_),
    .Q_N(_4464_),
    .Q(\logix.ram_r[524] ));
 sg13g2_dfrbp_1 \logix.ram_r[525]$_DFFE_PP_  (.CLK(net731),
    .RESET_B(net2326),
    .D(_1535_),
    .Q_N(_4463_),
    .Q(\logix.ram_r[525] ));
 sg13g2_dfrbp_1 \logix.ram_r[526]$_DFFE_PP_  (.CLK(net695),
    .RESET_B(net2327),
    .D(_1536_),
    .Q_N(_4462_),
    .Q(\logix.ram_r[526] ));
 sg13g2_dfrbp_1 \logix.ram_r[527]$_DFFE_PP_  (.CLK(net695),
    .RESET_B(net2328),
    .D(_1537_),
    .Q_N(_4461_),
    .Q(\logix.ram_r[527] ));
 sg13g2_dfrbp_1 \logix.ram_r[528]$_DFFE_PP_  (.CLK(net726),
    .RESET_B(net2329),
    .D(_1538_),
    .Q_N(_4460_),
    .Q(\logix.ram_r[528] ));
 sg13g2_dfrbp_1 \logix.ram_r[529]$_DFFE_PP_  (.CLK(net726),
    .RESET_B(net2330),
    .D(_1539_),
    .Q_N(_4459_),
    .Q(\logix.ram_r[529] ));
 sg13g2_dfrbp_1 \logix.ram_r[52]$_DFFE_PP_  (.CLK(net658),
    .RESET_B(net2331),
    .D(_1540_),
    .Q_N(_4458_),
    .Q(\logix.ram_r[52] ));
 sg13g2_dfrbp_1 \logix.ram_r[530]$_DFFE_PP_  (.CLK(net728),
    .RESET_B(net2332),
    .D(_1541_),
    .Q_N(_4457_),
    .Q(\logix.ram_r[530] ));
 sg13g2_dfrbp_1 \logix.ram_r[531]$_DFFE_PP_  (.CLK(net731),
    .RESET_B(net2333),
    .D(_1542_),
    .Q_N(_4456_),
    .Q(\logix.ram_r[531] ));
 sg13g2_dfrbp_1 \logix.ram_r[532]$_DFFE_PP_  (.CLK(net732),
    .RESET_B(net2334),
    .D(_1543_),
    .Q_N(_4455_),
    .Q(\logix.ram_r[532] ));
 sg13g2_dfrbp_1 \logix.ram_r[533]$_DFFE_PP_  (.CLK(net731),
    .RESET_B(net2335),
    .D(_1544_),
    .Q_N(_4454_),
    .Q(\logix.ram_r[533] ));
 sg13g2_dfrbp_1 \logix.ram_r[534]$_DFFE_PP_  (.CLK(net699),
    .RESET_B(net2336),
    .D(_1545_),
    .Q_N(_4453_),
    .Q(\logix.ram_r[534] ));
 sg13g2_dfrbp_1 \logix.ram_r[535]$_DFFE_PP_  (.CLK(net695),
    .RESET_B(net2337),
    .D(_1546_),
    .Q_N(_4452_),
    .Q(\logix.ram_r[535] ));
 sg13g2_dfrbp_1 \logix.ram_r[536]$_DFFE_PP_  (.CLK(net726),
    .RESET_B(net2338),
    .D(_1547_),
    .Q_N(_4451_),
    .Q(\logix.ram_r[536] ));
 sg13g2_dfrbp_1 \logix.ram_r[537]$_DFFE_PP_  (.CLK(net730),
    .RESET_B(net2339),
    .D(_1548_),
    .Q_N(_4450_),
    .Q(\logix.ram_r[537] ));
 sg13g2_dfrbp_1 \logix.ram_r[538]$_DFFE_PP_  (.CLK(net730),
    .RESET_B(net2340),
    .D(_1549_),
    .Q_N(_4449_),
    .Q(\logix.ram_r[538] ));
 sg13g2_dfrbp_1 \logix.ram_r[539]$_DFFE_PP_  (.CLK(net732),
    .RESET_B(net2341),
    .D(_1550_),
    .Q_N(_4448_),
    .Q(\logix.ram_r[539] ));
 sg13g2_dfrbp_1 \logix.ram_r[53]$_DFFE_PP_  (.CLK(net658),
    .RESET_B(net2342),
    .D(_1551_),
    .Q_N(_4447_),
    .Q(\logix.ram_r[53] ));
 sg13g2_dfrbp_1 \logix.ram_r[540]$_DFFE_PP_  (.CLK(net731),
    .RESET_B(net2343),
    .D(_1552_),
    .Q_N(_4446_),
    .Q(\logix.ram_r[540] ));
 sg13g2_dfrbp_1 \logix.ram_r[541]$_DFFE_PP_  (.CLK(net731),
    .RESET_B(net2344),
    .D(_1553_),
    .Q_N(_4445_),
    .Q(\logix.ram_r[541] ));
 sg13g2_dfrbp_1 \logix.ram_r[542]$_DFFE_PP_  (.CLK(net731),
    .RESET_B(net2345),
    .D(_1554_),
    .Q_N(_4444_),
    .Q(\logix.ram_r[542] ));
 sg13g2_dfrbp_1 \logix.ram_r[543]$_DFFE_PP_  (.CLK(net726),
    .RESET_B(net2346),
    .D(_1555_),
    .Q_N(_4443_),
    .Q(\logix.ram_r[543] ));
 sg13g2_dfrbp_1 \logix.ram_r[544]$_DFFE_PP_  (.CLK(net727),
    .RESET_B(net2347),
    .D(_1556_),
    .Q_N(_4442_),
    .Q(\logix.ram_r[544] ));
 sg13g2_dfrbp_1 \logix.ram_r[545]$_DFFE_PP_  (.CLK(net727),
    .RESET_B(net2348),
    .D(_1557_),
    .Q_N(_4441_),
    .Q(\logix.ram_r[545] ));
 sg13g2_dfrbp_1 \logix.ram_r[546]$_DFFE_PP_  (.CLK(net662),
    .RESET_B(net2349),
    .D(_1558_),
    .Q_N(_4440_),
    .Q(\logix.ram_r[546] ));
 sg13g2_dfrbp_1 \logix.ram_r[547]$_DFFE_PP_  (.CLK(net658),
    .RESET_B(net2350),
    .D(_1559_),
    .Q_N(_4439_),
    .Q(\logix.ram_r[547] ));
 sg13g2_dfrbp_1 \logix.ram_r[548]$_DFFE_PP_  (.CLK(net662),
    .RESET_B(net2351),
    .D(_1560_),
    .Q_N(_4438_),
    .Q(\logix.ram_r[548] ));
 sg13g2_dfrbp_1 \logix.ram_r[549]$_DFFE_PP_  (.CLK(net662),
    .RESET_B(net2352),
    .D(_1561_),
    .Q_N(_4437_),
    .Q(\logix.ram_r[549] ));
 sg13g2_dfrbp_1 \logix.ram_r[54]$_DFFE_PP_  (.CLK(net658),
    .RESET_B(net2353),
    .D(_1562_),
    .Q_N(_4436_),
    .Q(\logix.ram_r[54] ));
 sg13g2_dfrbp_1 \logix.ram_r[550]$_DFFE_PP_  (.CLK(net663),
    .RESET_B(net2354),
    .D(_1563_),
    .Q_N(_4435_),
    .Q(\logix.ram_r[550] ));
 sg13g2_dfrbp_1 \logix.ram_r[551]$_DFFE_PP_  (.CLK(net663),
    .RESET_B(net2355),
    .D(_1564_),
    .Q_N(_4434_),
    .Q(\logix.ram_r[551] ));
 sg13g2_dfrbp_1 \logix.ram_r[552]$_DFFE_PP_  (.CLK(net727),
    .RESET_B(net2356),
    .D(_1565_),
    .Q_N(_4433_),
    .Q(\logix.ram_r[552] ));
 sg13g2_dfrbp_1 \logix.ram_r[553]$_DFFE_PP_  (.CLK(net727),
    .RESET_B(net2357),
    .D(_1566_),
    .Q_N(_4432_),
    .Q(\logix.ram_r[553] ));
 sg13g2_dfrbp_1 \logix.ram_r[554]$_DFFE_PP_  (.CLK(net664),
    .RESET_B(net2358),
    .D(_1567_),
    .Q_N(_4431_),
    .Q(\logix.ram_r[554] ));
 sg13g2_dfrbp_1 \logix.ram_r[555]$_DFFE_PP_  (.CLK(net664),
    .RESET_B(net2359),
    .D(_1568_),
    .Q_N(_4430_),
    .Q(\logix.ram_r[555] ));
 sg13g2_dfrbp_1 \logix.ram_r[556]$_DFFE_PP_  (.CLK(net662),
    .RESET_B(net2360),
    .D(_1569_),
    .Q_N(_4429_),
    .Q(\logix.ram_r[556] ));
 sg13g2_dfrbp_1 \logix.ram_r[557]$_DFFE_PP_  (.CLK(net662),
    .RESET_B(net2361),
    .D(_1570_),
    .Q_N(_4428_),
    .Q(\logix.ram_r[557] ));
 sg13g2_dfrbp_1 \logix.ram_r[558]$_DFFE_PP_  (.CLK(net663),
    .RESET_B(net2362),
    .D(_1571_),
    .Q_N(_4427_),
    .Q(\logix.ram_r[558] ));
 sg13g2_dfrbp_1 \logix.ram_r[559]$_DFFE_PP_  (.CLK(net663),
    .RESET_B(net2363),
    .D(_1572_),
    .Q_N(_4426_),
    .Q(\logix.ram_r[559] ));
 sg13g2_dfrbp_1 \logix.ram_r[55]$_DFFE_PP_  (.CLK(net657),
    .RESET_B(net2364),
    .D(_1573_),
    .Q_N(_4425_),
    .Q(\logix.ram_r[55] ));
 sg13g2_dfrbp_1 \logix.ram_r[560]$_DFFE_PP_  (.CLK(net663),
    .RESET_B(net2365),
    .D(_1574_),
    .Q_N(_4424_),
    .Q(\logix.ram_r[560] ));
 sg13g2_dfrbp_1 \logix.ram_r[561]$_DFFE_PP_  (.CLK(net665),
    .RESET_B(net2366),
    .D(_1575_),
    .Q_N(_4423_),
    .Q(\logix.ram_r[561] ));
 sg13g2_dfrbp_1 \logix.ram_r[562]$_DFFE_PP_  (.CLK(net665),
    .RESET_B(net2367),
    .D(_1576_),
    .Q_N(_4422_),
    .Q(\logix.ram_r[562] ));
 sg13g2_dfrbp_1 \logix.ram_r[563]$_DFFE_PP_  (.CLK(net664),
    .RESET_B(net2368),
    .D(_1577_),
    .Q_N(_4421_),
    .Q(\logix.ram_r[563] ));
 sg13g2_dfrbp_1 \logix.ram_r[564]$_DFFE_PP_  (.CLK(net662),
    .RESET_B(net2369),
    .D(_1578_),
    .Q_N(_4420_),
    .Q(\logix.ram_r[564] ));
 sg13g2_dfrbp_1 \logix.ram_r[565]$_DFFE_PP_  (.CLK(net662),
    .RESET_B(net2370),
    .D(_1579_),
    .Q_N(_4419_),
    .Q(\logix.ram_r[565] ));
 sg13g2_dfrbp_1 \logix.ram_r[566]$_DFFE_PP_  (.CLK(net663),
    .RESET_B(net2371),
    .D(_1580_),
    .Q_N(_4418_),
    .Q(\logix.ram_r[566] ));
 sg13g2_dfrbp_1 \logix.ram_r[567]$_DFFE_PP_  (.CLK(net727),
    .RESET_B(net2372),
    .D(_1581_),
    .Q_N(_4417_),
    .Q(\logix.ram_r[567] ));
 sg13g2_dfrbp_1 \logix.ram_r[568]$_DFFE_PP_  (.CLK(net727),
    .RESET_B(net2373),
    .D(_1582_),
    .Q_N(_4416_),
    .Q(\logix.ram_r[568] ));
 sg13g2_dfrbp_1 \logix.ram_r[569]$_DFFE_PP_  (.CLK(net729),
    .RESET_B(net2374),
    .D(_1583_),
    .Q_N(_4415_),
    .Q(\logix.ram_r[569] ));
 sg13g2_dfrbp_1 \logix.ram_r[56]$_DFFE_PP_  (.CLK(net657),
    .RESET_B(net2375),
    .D(_1584_),
    .Q_N(_4414_),
    .Q(\logix.ram_r[56] ));
 sg13g2_dfrbp_1 \logix.ram_r[570]$_DFFE_PP_  (.CLK(net665),
    .RESET_B(net2376),
    .D(_1585_),
    .Q_N(_4413_),
    .Q(\logix.ram_r[570] ));
 sg13g2_dfrbp_1 \logix.ram_r[571]$_DFFE_PP_  (.CLK(net664),
    .RESET_B(net2377),
    .D(_1586_),
    .Q_N(_4412_),
    .Q(\logix.ram_r[571] ));
 sg13g2_dfrbp_1 \logix.ram_r[572]$_DFFE_PP_  (.CLK(net662),
    .RESET_B(net2378),
    .D(_1587_),
    .Q_N(_4411_),
    .Q(\logix.ram_r[572] ));
 sg13g2_dfrbp_1 \logix.ram_r[573]$_DFFE_PP_  (.CLK(net663),
    .RESET_B(net2379),
    .D(_1588_),
    .Q_N(_4410_),
    .Q(\logix.ram_r[573] ));
 sg13g2_dfrbp_1 \logix.ram_r[574]$_DFFE_PP_  (.CLK(net630),
    .RESET_B(net2380),
    .D(_1589_),
    .Q_N(_4409_),
    .Q(\logix.ram_r[574] ));
 sg13g2_dfrbp_1 \logix.ram_r[575]$_DFFE_PP_  (.CLK(net630),
    .RESET_B(net2381),
    .D(_1590_),
    .Q_N(_4408_),
    .Q(\logix.ram_r[575] ));
 sg13g2_dfrbp_1 \logix.ram_r[576]$_DFFE_PP_  (.CLK(net694),
    .RESET_B(net2382),
    .D(_1591_),
    .Q_N(_4407_),
    .Q(\logix.ram_r[576] ));
 sg13g2_dfrbp_1 \logix.ram_r[577]$_DFFE_PP_  (.CLK(net694),
    .RESET_B(net2383),
    .D(_1592_),
    .Q_N(_4406_),
    .Q(\logix.ram_r[577] ));
 sg13g2_dfrbp_1 \logix.ram_r[578]$_DFFE_PP_  (.CLK(net630),
    .RESET_B(net2384),
    .D(_1593_),
    .Q_N(_4405_),
    .Q(\logix.ram_r[578] ));
 sg13g2_dfrbp_1 \logix.ram_r[579]$_DFFE_PP_  (.CLK(net631),
    .RESET_B(net2385),
    .D(_1594_),
    .Q_N(_4404_),
    .Q(\logix.ram_r[579] ));
 sg13g2_dfrbp_1 \logix.ram_r[57]$_DFFE_PP_  (.CLK(net657),
    .RESET_B(net2386),
    .D(_1595_),
    .Q_N(_4403_),
    .Q(\logix.ram_r[57] ));
 sg13g2_dfrbp_1 \logix.ram_r[580]$_DFFE_PP_  (.CLK(net631),
    .RESET_B(net2387),
    .D(_1596_),
    .Q_N(_4402_),
    .Q(\logix.ram_r[580] ));
 sg13g2_dfrbp_1 \logix.ram_r[581]$_DFFE_PP_  (.CLK(net630),
    .RESET_B(net2388),
    .D(_1597_),
    .Q_N(_4401_),
    .Q(\logix.ram_r[581] ));
 sg13g2_dfrbp_1 \logix.ram_r[582]$_DFFE_PP_  (.CLK(net630),
    .RESET_B(net2389),
    .D(_1598_),
    .Q_N(_4400_),
    .Q(\logix.ram_r[582] ));
 sg13g2_dfrbp_1 \logix.ram_r[583]$_DFFE_PP_  (.CLK(net630),
    .RESET_B(net2390),
    .D(_1599_),
    .Q_N(_4399_),
    .Q(\logix.ram_r[583] ));
 sg13g2_dfrbp_1 \logix.ram_r[584]$_DFFE_PP_  (.CLK(net630),
    .RESET_B(net2391),
    .D(_1600_),
    .Q_N(_4398_),
    .Q(\logix.ram_r[584] ));
 sg13g2_dfrbp_1 \logix.ram_r[585]$_DFFE_PP_  (.CLK(net630),
    .RESET_B(net2392),
    .D(_1601_),
    .Q_N(_4397_),
    .Q(\logix.ram_r[585] ));
 sg13g2_dfrbp_1 \logix.ram_r[586]$_DFFE_PP_  (.CLK(net631),
    .RESET_B(net2393),
    .D(_1602_),
    .Q_N(_4396_),
    .Q(\logix.ram_r[586] ));
 sg13g2_dfrbp_1 \logix.ram_r[587]$_DFFE_PP_  (.CLK(net625),
    .RESET_B(net2394),
    .D(_1603_),
    .Q_N(_4395_),
    .Q(\logix.ram_r[587] ));
 sg13g2_dfrbp_1 \logix.ram_r[588]$_DFFE_PP_  (.CLK(net625),
    .RESET_B(net2395),
    .D(_1604_),
    .Q_N(_4394_),
    .Q(\logix.ram_r[588] ));
 sg13g2_dfrbp_1 \logix.ram_r[589]$_DFFE_PP_  (.CLK(net628),
    .RESET_B(net2396),
    .D(_1605_),
    .Q_N(_4393_),
    .Q(\logix.ram_r[589] ));
 sg13g2_dfrbp_1 \logix.ram_r[58]$_DFFE_PP_  (.CLK(net625),
    .RESET_B(net2397),
    .D(_1606_),
    .Q_N(_4392_),
    .Q(\logix.ram_r[58] ));
 sg13g2_dfrbp_1 \logix.ram_r[590]$_DFFE_PP_  (.CLK(net628),
    .RESET_B(net2398),
    .D(_1607_),
    .Q_N(_4391_),
    .Q(\logix.ram_r[590] ));
 sg13g2_dfrbp_1 \logix.ram_r[591]$_DFFE_PP_  (.CLK(net692),
    .RESET_B(net2399),
    .D(_1608_),
    .Q_N(_4390_),
    .Q(\logix.ram_r[591] ));
 sg13g2_dfrbp_1 \logix.ram_r[592]$_DFFE_PP_  (.CLK(net694),
    .RESET_B(net2400),
    .D(_1609_),
    .Q_N(_4389_),
    .Q(\logix.ram_r[592] ));
 sg13g2_dfrbp_1 \logix.ram_r[593]$_DFFE_PP_  (.CLK(net694),
    .RESET_B(net2401),
    .D(_1610_),
    .Q_N(_4388_),
    .Q(\logix.ram_r[593] ));
 sg13g2_dfrbp_1 \logix.ram_r[594]$_DFFE_PP_  (.CLK(net694),
    .RESET_B(net2402),
    .D(_1611_),
    .Q_N(_4387_),
    .Q(\logix.ram_r[594] ));
 sg13g2_dfrbp_1 \logix.ram_r[595]$_DFFE_PP_  (.CLK(net626),
    .RESET_B(net2403),
    .D(_1612_),
    .Q_N(_4386_),
    .Q(\logix.ram_r[595] ));
 sg13g2_dfrbp_1 \logix.ram_r[596]$_DFFE_PP_  (.CLK(net624),
    .RESET_B(net2404),
    .D(_1613_),
    .Q_N(_4385_),
    .Q(\logix.ram_r[596] ));
 sg13g2_dfrbp_1 \logix.ram_r[597]$_DFFE_PP_  (.CLK(net628),
    .RESET_B(net2405),
    .D(_1614_),
    .Q_N(_4384_),
    .Q(\logix.ram_r[597] ));
 sg13g2_dfrbp_1 \logix.ram_r[598]$_DFFE_PP_  (.CLK(net629),
    .RESET_B(net2406),
    .D(_1615_),
    .Q_N(_4383_),
    .Q(\logix.ram_r[598] ));
 sg13g2_dfrbp_1 \logix.ram_r[599]$_DFFE_PP_  (.CLK(net692),
    .RESET_B(net2407),
    .D(_1616_),
    .Q_N(_4382_),
    .Q(\logix.ram_r[599] ));
 sg13g2_dfrbp_1 \logix.ram_r[59]$_DFFE_PP_  (.CLK(net626),
    .RESET_B(net2408),
    .D(_1617_),
    .Q_N(_4381_),
    .Q(\logix.ram_r[59] ));
 sg13g2_dfrbp_1 \logix.ram_r[5]$_DFFE_PP_  (.CLK(net609),
    .RESET_B(net2409),
    .D(_1618_),
    .Q_N(_4380_),
    .Q(\logix.ram_r[5] ));
 sg13g2_dfrbp_1 \logix.ram_r[600]$_DFFE_PP_  (.CLK(net694),
    .RESET_B(net2410),
    .D(_1619_),
    .Q_N(_4379_),
    .Q(\logix.ram_r[600] ));
 sg13g2_dfrbp_1 \logix.ram_r[601]$_DFFE_PP_  (.CLK(net695),
    .RESET_B(net2411),
    .D(_1620_),
    .Q_N(_4378_),
    .Q(\logix.ram_r[601] ));
 sg13g2_dfrbp_1 \logix.ram_r[602]$_DFFE_PP_  (.CLK(net695),
    .RESET_B(net2412),
    .D(_1621_),
    .Q_N(_4377_),
    .Q(\logix.ram_r[602] ));
 sg13g2_dfrbp_1 \logix.ram_r[603]$_DFFE_PP_  (.CLK(net631),
    .RESET_B(net2413),
    .D(_1622_),
    .Q_N(_4376_),
    .Q(\logix.ram_r[603] ));
 sg13g2_dfrbp_1 \logix.ram_r[604]$_DFFE_PP_  (.CLK(net631),
    .RESET_B(net2414),
    .D(_1623_),
    .Q_N(_4375_),
    .Q(\logix.ram_r[604] ));
 sg13g2_dfrbp_1 \logix.ram_r[605]$_DFFE_PP_  (.CLK(net628),
    .RESET_B(net2415),
    .D(_1624_),
    .Q_N(_4374_),
    .Q(\logix.ram_r[605] ));
 sg13g2_dfrbp_1 \logix.ram_r[606]$_DFFE_PP_  (.CLK(net629),
    .RESET_B(net2416),
    .D(_1625_),
    .Q_N(_4373_),
    .Q(\logix.ram_r[606] ));
 sg13g2_dfrbp_1 \logix.ram_r[607]$_DFFE_PP_  (.CLK(net693),
    .RESET_B(net2417),
    .D(_1626_),
    .Q_N(_4372_),
    .Q(\logix.ram_r[607] ));
 sg13g2_dfrbp_1 \logix.ram_r[608]$_DFFE_PP_  (.CLK(net693),
    .RESET_B(net2418),
    .D(_1627_),
    .Q_N(_4371_),
    .Q(\logix.ram_r[608] ));
 sg13g2_dfrbp_1 \logix.ram_r[609]$_DFFE_PP_  (.CLK(net692),
    .RESET_B(net2419),
    .D(_1628_),
    .Q_N(_4370_),
    .Q(\logix.ram_r[609] ));
 sg13g2_dfrbp_1 \logix.ram_r[60]$_DFFE_PP_  (.CLK(net626),
    .RESET_B(net2420),
    .D(_1629_),
    .Q_N(_4369_),
    .Q(\logix.ram_r[60] ));
 sg13g2_dfrbp_1 \logix.ram_r[610]$_DFFE_PP_  (.CLK(net692),
    .RESET_B(net2421),
    .D(_1630_),
    .Q_N(_4368_),
    .Q(\logix.ram_r[610] ));
 sg13g2_dfrbp_1 \logix.ram_r[611]$_DFFE_PP_  (.CLK(net628),
    .RESET_B(net2422),
    .D(_1631_),
    .Q_N(_4367_),
    .Q(\logix.ram_r[611] ));
 sg13g2_dfrbp_1 \logix.ram_r[612]$_DFFE_PP_  (.CLK(net621),
    .RESET_B(net2423),
    .D(_1632_),
    .Q_N(_4366_),
    .Q(\logix.ram_r[612] ));
 sg13g2_dfrbp_1 \logix.ram_r[613]$_DFFE_PP_  (.CLK(net620),
    .RESET_B(net2424),
    .D(_1633_),
    .Q_N(_4365_),
    .Q(\logix.ram_r[613] ));
 sg13g2_dfrbp_1 \logix.ram_r[614]$_DFFE_PP_  (.CLK(net620),
    .RESET_B(net2425),
    .D(_1634_),
    .Q_N(_4364_),
    .Q(\logix.ram_r[614] ));
 sg13g2_dfrbp_1 \logix.ram_r[615]$_DFFE_PP_  (.CLK(net683),
    .RESET_B(net2426),
    .D(_1635_),
    .Q_N(_4363_),
    .Q(\logix.ram_r[615] ));
 sg13g2_dfrbp_1 \logix.ram_r[616]$_DFFE_PP_  (.CLK(net683),
    .RESET_B(net2427),
    .D(_1636_),
    .Q_N(_4362_),
    .Q(\logix.ram_r[616] ));
 sg13g2_dfrbp_1 \logix.ram_r[617]$_DFFE_PP_  (.CLK(net692),
    .RESET_B(net2428),
    .D(_1637_),
    .Q_N(_4361_),
    .Q(\logix.ram_r[617] ));
 sg13g2_dfrbp_1 \logix.ram_r[618]$_DFFE_PP_  (.CLK(net629),
    .RESET_B(net2429),
    .D(_1638_),
    .Q_N(_4360_),
    .Q(\logix.ram_r[618] ));
 sg13g2_dfrbp_1 \logix.ram_r[619]$_DFFE_PP_  (.CLK(net628),
    .RESET_B(net2430),
    .D(_1639_),
    .Q_N(_4359_),
    .Q(\logix.ram_r[619] ));
 sg13g2_dfrbp_1 \logix.ram_r[61]$_DFFE_PP_  (.CLK(net631),
    .RESET_B(net2431),
    .D(_1640_),
    .Q_N(_4358_),
    .Q(\logix.ram_r[61] ));
 sg13g2_dfrbp_1 \logix.ram_r[620]$_DFFE_PP_  (.CLK(net621),
    .RESET_B(net2432),
    .D(_1641_),
    .Q_N(_4357_),
    .Q(\logix.ram_r[620] ));
 sg13g2_dfrbp_1 \logix.ram_r[621]$_DFFE_PP_  (.CLK(net620),
    .RESET_B(net2433),
    .D(_1642_),
    .Q_N(_4356_),
    .Q(\logix.ram_r[621] ));
 sg13g2_dfrbp_1 \logix.ram_r[622]$_DFFE_PP_  (.CLK(net620),
    .RESET_B(net2434),
    .D(_1643_),
    .Q_N(_4355_),
    .Q(\logix.ram_r[622] ));
 sg13g2_dfrbp_1 \logix.ram_r[623]$_DFFE_PP_  (.CLK(net683),
    .RESET_B(net2435),
    .D(_1644_),
    .Q_N(_4354_),
    .Q(\logix.ram_r[623] ));
 sg13g2_dfrbp_1 \logix.ram_r[624]$_DFFE_PP_  (.CLK(net683),
    .RESET_B(net2436),
    .D(_1645_),
    .Q_N(_4353_),
    .Q(\logix.ram_r[624] ));
 sg13g2_dfrbp_1 \logix.ram_r[625]$_DFFE_PP_  (.CLK(net692),
    .RESET_B(net2437),
    .D(_1646_),
    .Q_N(_4352_),
    .Q(\logix.ram_r[625] ));
 sg13g2_dfrbp_1 \logix.ram_r[626]$_DFFE_PP_  (.CLK(net629),
    .RESET_B(net2438),
    .D(_1647_),
    .Q_N(_4351_),
    .Q(\logix.ram_r[626] ));
 sg13g2_dfrbp_1 \logix.ram_r[627]$_DFFE_PP_  (.CLK(net628),
    .RESET_B(net2439),
    .D(_1648_),
    .Q_N(_4350_),
    .Q(\logix.ram_r[627] ));
 sg13g2_dfrbp_1 \logix.ram_r[628]$_DFFE_PP_  (.CLK(net629),
    .RESET_B(net2440),
    .D(_1649_),
    .Q_N(_4349_),
    .Q(\logix.ram_r[628] ));
 sg13g2_dfrbp_1 \logix.ram_r[629]$_DFFE_PP_  (.CLK(net620),
    .RESET_B(net2441),
    .D(_1650_),
    .Q_N(_4348_),
    .Q(\logix.ram_r[629] ));
 sg13g2_dfrbp_1 \logix.ram_r[62]$_DFFE_PP_  (.CLK(net631),
    .RESET_B(net2442),
    .D(_1651_),
    .Q_N(_4347_),
    .Q(\logix.ram_r[62] ));
 sg13g2_dfrbp_1 \logix.ram_r[630]$_DFFE_PP_  (.CLK(net620),
    .RESET_B(net2443),
    .D(_1652_),
    .Q_N(_4346_),
    .Q(\logix.ram_r[630] ));
 sg13g2_dfrbp_1 \logix.ram_r[631]$_DFFE_PP_  (.CLK(net684),
    .RESET_B(net2444),
    .D(_1653_),
    .Q_N(_4345_),
    .Q(\logix.ram_r[631] ));
 sg13g2_dfrbp_1 \logix.ram_r[632]$_DFFE_PP_  (.CLK(net692),
    .RESET_B(net2445),
    .D(_1654_),
    .Q_N(_4344_),
    .Q(\logix.ram_r[632] ));
 sg13g2_dfrbp_1 \logix.ram_r[633]$_DFFE_PP_  (.CLK(net692),
    .RESET_B(net2446),
    .D(_1655_),
    .Q_N(_4343_),
    .Q(\logix.ram_r[633] ));
 sg13g2_dfrbp_1 \logix.ram_r[634]$_DFFE_PP_  (.CLK(net629),
    .RESET_B(net2447),
    .D(_1656_),
    .Q_N(_4342_),
    .Q(\logix.ram_r[634] ));
 sg13g2_dfrbp_1 \logix.ram_r[635]$_DFFE_PP_  (.CLK(net628),
    .RESET_B(net2448),
    .D(_1657_),
    .Q_N(_4341_),
    .Q(\logix.ram_r[635] ));
 sg13g2_dfrbp_1 \logix.ram_r[636]$_DFFE_PP_  (.CLK(net622),
    .RESET_B(net2449),
    .D(_1658_),
    .Q_N(_4340_),
    .Q(\logix.ram_r[636] ));
 sg13g2_dfrbp_1 \logix.ram_r[637]$_DFFE_PP_  (.CLK(net620),
    .RESET_B(net2450),
    .D(_1659_),
    .Q_N(_4339_),
    .Q(\logix.ram_r[637] ));
 sg13g2_dfrbp_1 \logix.ram_r[638]$_DFFE_PP_  (.CLK(net620),
    .RESET_B(net2451),
    .D(_1660_),
    .Q_N(_4338_),
    .Q(\logix.ram_r[638] ));
 sg13g2_dfrbp_1 \logix.ram_r[639]$_DFFE_PP_  (.CLK(net683),
    .RESET_B(net2452),
    .D(_1661_),
    .Q_N(_4337_),
    .Q(\logix.ram_r[639] ));
 sg13g2_dfrbp_1 \logix.ram_r[63]$_DFFE_PP_  (.CLK(net624),
    .RESET_B(net2453),
    .D(_1662_),
    .Q_N(_4336_),
    .Q(\logix.ram_r[63] ));
 sg13g2_dfrbp_1 \logix.ram_r[640]$_DFFE_PP_  (.CLK(net683),
    .RESET_B(net2454),
    .D(_1663_),
    .Q_N(_4335_),
    .Q(\logix.ram_r[640] ));
 sg13g2_dfrbp_1 \logix.ram_r[641]$_DFFE_PP_  (.CLK(net683),
    .RESET_B(net2455),
    .D(_1664_),
    .Q_N(_4334_),
    .Q(\logix.ram_r[641] ));
 sg13g2_dfrbp_1 \logix.ram_r[642]$_DFFE_PP_  (.CLK(net683),
    .RESET_B(net2456),
    .D(_1665_),
    .Q_N(_4333_),
    .Q(\logix.ram_r[642] ));
 sg13g2_dfrbp_1 \logix.ram_r[643]$_DFFE_PP_  (.CLK(net618),
    .RESET_B(net2457),
    .D(_1666_),
    .Q_N(_4332_),
    .Q(\logix.ram_r[643] ));
 sg13g2_dfrbp_1 \logix.ram_r[644]$_DFFE_PP_  (.CLK(net618),
    .RESET_B(net2458),
    .D(_1667_),
    .Q_N(_4331_),
    .Q(\logix.ram_r[644] ));
 sg13g2_dfrbp_1 \logix.ram_r[645]$_DFFE_PP_  (.CLK(net618),
    .RESET_B(net2459),
    .D(_1668_),
    .Q_N(_4330_),
    .Q(\logix.ram_r[645] ));
 sg13g2_dfrbp_1 \logix.ram_r[646]$_DFFE_PP_  (.CLK(net618),
    .RESET_B(net2460),
    .D(_1669_),
    .Q_N(_4329_),
    .Q(\logix.ram_r[646] ));
 sg13g2_dfrbp_1 \logix.ram_r[647]$_DFFE_PP_  (.CLK(net680),
    .RESET_B(net2461),
    .D(_1670_),
    .Q_N(_4328_),
    .Q(\logix.ram_r[647] ));
 sg13g2_dfrbp_1 \logix.ram_r[648]$_DFFE_PP_  (.CLK(net680),
    .RESET_B(net2462),
    .D(_1671_),
    .Q_N(_4327_),
    .Q(\logix.ram_r[648] ));
 sg13g2_dfrbp_1 \logix.ram_r[649]$_DFFE_PP_  (.CLK(net680),
    .RESET_B(net2463),
    .D(_1672_),
    .Q_N(_4326_),
    .Q(\logix.ram_r[649] ));
 sg13g2_dfrbp_1 \logix.ram_r[64]$_DFFE_PP_  (.CLK(net624),
    .RESET_B(net2464),
    .D(_1673_),
    .Q_N(_4325_),
    .Q(\logix.ram_r[64] ));
 sg13g2_dfrbp_1 \logix.ram_r[650]$_DFFE_PP_  (.CLK(net680),
    .RESET_B(net2465),
    .D(_1674_),
    .Q_N(_4324_),
    .Q(\logix.ram_r[650] ));
 sg13g2_dfrbp_1 \logix.ram_r[651]$_DFFE_PP_  (.CLK(net682),
    .RESET_B(net2466),
    .D(_1675_),
    .Q_N(_4323_),
    .Q(\logix.ram_r[651] ));
 sg13g2_dfrbp_1 \logix.ram_r[652]$_DFFE_PP_  (.CLK(net622),
    .RESET_B(net2467),
    .D(_1676_),
    .Q_N(_4322_),
    .Q(\logix.ram_r[652] ));
 sg13g2_dfrbp_1 \logix.ram_r[653]$_DFFE_PP_  (.CLK(net618),
    .RESET_B(net2468),
    .D(_1677_),
    .Q_N(_4321_),
    .Q(\logix.ram_r[653] ));
 sg13g2_dfrbp_1 \logix.ram_r[654]$_DFFE_PP_  (.CLK(net680),
    .RESET_B(net2469),
    .D(_1678_),
    .Q_N(_4320_),
    .Q(\logix.ram_r[654] ));
 sg13g2_dfrbp_1 \logix.ram_r[655]$_DFFE_PP_  (.CLK(net680),
    .RESET_B(net2470),
    .D(_1679_),
    .Q_N(_4319_),
    .Q(\logix.ram_r[655] ));
 sg13g2_dfrbp_1 \logix.ram_r[656]$_DFFE_PP_  (.CLK(net681),
    .RESET_B(net2471),
    .D(_1680_),
    .Q_N(_4318_),
    .Q(\logix.ram_r[656] ));
 sg13g2_dfrbp_1 \logix.ram_r[657]$_DFFE_PP_  (.CLK(net681),
    .RESET_B(net2472),
    .D(_1681_),
    .Q_N(_4317_),
    .Q(\logix.ram_r[657] ));
 sg13g2_dfrbp_1 \logix.ram_r[658]$_DFFE_PP_  (.CLK(net681),
    .RESET_B(net2473),
    .D(_1682_),
    .Q_N(_4316_),
    .Q(\logix.ram_r[658] ));
 sg13g2_dfrbp_1 \logix.ram_r[659]$_DFFE_PP_  (.CLK(net682),
    .RESET_B(net2474),
    .D(_1683_),
    .Q_N(_4315_),
    .Q(\logix.ram_r[659] ));
 sg13g2_dfrbp_1 \logix.ram_r[65]$_DFFE_PP_  (.CLK(net624),
    .RESET_B(net2475),
    .D(_1684_),
    .Q_N(_4314_),
    .Q(\logix.ram_r[65] ));
 sg13g2_dfrbp_1 \logix.ram_r[660]$_DFFE_PP_  (.CLK(net622),
    .RESET_B(net2476),
    .D(_1685_),
    .Q_N(_4313_),
    .Q(\logix.ram_r[660] ));
 sg13g2_dfrbp_1 \logix.ram_r[661]$_DFFE_PP_  (.CLK(net618),
    .RESET_B(net2477),
    .D(_1686_),
    .Q_N(_4312_),
    .Q(\logix.ram_r[661] ));
 sg13g2_dfrbp_1 \logix.ram_r[662]$_DFFE_PP_  (.CLK(net680),
    .RESET_B(net2478),
    .D(_1687_),
    .Q_N(_4311_),
    .Q(\logix.ram_r[662] ));
 sg13g2_dfrbp_1 \logix.ram_r[663]$_DFFE_PP_  (.CLK(net680),
    .RESET_B(net2479),
    .D(_1688_),
    .Q_N(_4310_),
    .Q(\logix.ram_r[663] ));
 sg13g2_dfrbp_1 \logix.ram_r[664]$_DFFE_PP_  (.CLK(net681),
    .RESET_B(net2480),
    .D(_1689_),
    .Q_N(_4309_),
    .Q(\logix.ram_r[664] ));
 sg13g2_dfrbp_1 \logix.ram_r[665]$_DFFE_PP_  (.CLK(net681),
    .RESET_B(net2481),
    .D(_1690_),
    .Q_N(_4308_),
    .Q(\logix.ram_r[665] ));
 sg13g2_dfrbp_1 \logix.ram_r[666]$_DFFE_PP_  (.CLK(net681),
    .RESET_B(net2482),
    .D(_1691_),
    .Q_N(_4307_),
    .Q(\logix.ram_r[666] ));
 sg13g2_dfrbp_1 \logix.ram_r[667]$_DFFE_PP_  (.CLK(net682),
    .RESET_B(net2483),
    .D(_1692_),
    .Q_N(_4306_),
    .Q(\logix.ram_r[667] ));
 sg13g2_dfrbp_1 \logix.ram_r[668]$_DFFE_PP_  (.CLK(net622),
    .RESET_B(net2484),
    .D(_1693_),
    .Q_N(_4305_),
    .Q(\logix.ram_r[668] ));
 sg13g2_dfrbp_1 \logix.ram_r[669]$_DFFE_PP_  (.CLK(net618),
    .RESET_B(net2485),
    .D(_1694_),
    .Q_N(_4304_),
    .Q(\logix.ram_r[669] ));
 sg13g2_dfrbp_1 \logix.ram_r[66]$_DFFE_PP_  (.CLK(net624),
    .RESET_B(net2486),
    .D(_1695_),
    .Q_N(_4303_),
    .Q(\logix.ram_r[66] ));
 sg13g2_dfrbp_1 \logix.ram_r[670]$_DFFE_PP_  (.CLK(net618),
    .RESET_B(net2487),
    .D(_1696_),
    .Q_N(_4302_),
    .Q(\logix.ram_r[670] ));
 sg13g2_dfrbp_1 \logix.ram_r[671]$_DFFE_PP_  (.CLK(net619),
    .RESET_B(net2488),
    .D(_1697_),
    .Q_N(_4301_),
    .Q(\logix.ram_r[671] ));
 sg13g2_dfrbp_1 \logix.ram_r[672]$_DFFE_PP_  (.CLK(net619),
    .RESET_B(net2489),
    .D(_1698_),
    .Q_N(_4300_),
    .Q(\logix.ram_r[672] ));
 sg13g2_dfrbp_1 \logix.ram_r[673]$_DFFE_PP_  (.CLK(net621),
    .RESET_B(net2490),
    .D(_1699_),
    .Q_N(_4299_),
    .Q(\logix.ram_r[673] ));
 sg13g2_dfrbp_1 \logix.ram_r[674]$_DFFE_PP_  (.CLK(net621),
    .RESET_B(net2491),
    .D(_1700_),
    .Q_N(_4298_),
    .Q(\logix.ram_r[674] ));
 sg13g2_dfrbp_1 \logix.ram_r[675]$_DFFE_PP_  (.CLK(net615),
    .RESET_B(net2492),
    .D(_1701_),
    .Q_N(_4297_),
    .Q(\logix.ram_r[675] ));
 sg13g2_dfrbp_1 \logix.ram_r[676]$_DFFE_PP_  (.CLK(net615),
    .RESET_B(net2493),
    .D(_1702_),
    .Q_N(_4296_),
    .Q(\logix.ram_r[676] ));
 sg13g2_dfrbp_1 \logix.ram_r[677]$_DFFE_PP_  (.CLK(net612),
    .RESET_B(net2494),
    .D(_1703_),
    .Q_N(_4295_),
    .Q(\logix.ram_r[677] ));
 sg13g2_dfrbp_1 \logix.ram_r[678]$_DFFE_PP_  (.CLK(net612),
    .RESET_B(net2495),
    .D(_1704_),
    .Q_N(_4294_),
    .Q(\logix.ram_r[678] ));
 sg13g2_dfrbp_1 \logix.ram_r[679]$_DFFE_PP_  (.CLK(net612),
    .RESET_B(net2496),
    .D(_1705_),
    .Q_N(_4293_),
    .Q(\logix.ram_r[679] ));
 sg13g2_dfrbp_1 \logix.ram_r[67]$_DFFE_PP_  (.CLK(net615),
    .RESET_B(net2497),
    .D(_1706_),
    .Q_N(_4292_),
    .Q(\logix.ram_r[67] ));
 sg13g2_dfrbp_1 \logix.ram_r[680]$_DFFE_PP_  (.CLK(net619),
    .RESET_B(net2498),
    .D(_1707_),
    .Q_N(_4291_),
    .Q(\logix.ram_r[680] ));
 sg13g2_dfrbp_1 \logix.ram_r[681]$_DFFE_PP_  (.CLK(net621),
    .RESET_B(net2499),
    .D(_1708_),
    .Q_N(_4290_),
    .Q(\logix.ram_r[681] ));
 sg13g2_dfrbp_1 \logix.ram_r[682]$_DFFE_PP_  (.CLK(net615),
    .RESET_B(net2500),
    .D(_1709_),
    .Q_N(_4289_),
    .Q(\logix.ram_r[682] ));
 sg13g2_dfrbp_1 \logix.ram_r[683]$_DFFE_PP_  (.CLK(net616),
    .RESET_B(net2501),
    .D(_1710_),
    .Q_N(_4288_),
    .Q(\logix.ram_r[683] ));
 sg13g2_dfrbp_1 \logix.ram_r[684]$_DFFE_PP_  (.CLK(net616),
    .RESET_B(net2502),
    .D(_1711_),
    .Q_N(_4287_),
    .Q(\logix.ram_r[684] ));
 sg13g2_dfrbp_1 \logix.ram_r[685]$_DFFE_PP_  (.CLK(net612),
    .RESET_B(net2503),
    .D(_1712_),
    .Q_N(_4286_),
    .Q(\logix.ram_r[685] ));
 sg13g2_dfrbp_1 \logix.ram_r[686]$_DFFE_PP_  (.CLK(net612),
    .RESET_B(net2504),
    .D(_1713_),
    .Q_N(_4285_),
    .Q(\logix.ram_r[686] ));
 sg13g2_dfrbp_1 \logix.ram_r[687]$_DFFE_PP_  (.CLK(net619),
    .RESET_B(net2505),
    .D(_1714_),
    .Q_N(_4284_),
    .Q(\logix.ram_r[687] ));
 sg13g2_dfrbp_1 \logix.ram_r[688]$_DFFE_PP_  (.CLK(net619),
    .RESET_B(net2506),
    .D(_1715_),
    .Q_N(_4283_),
    .Q(\logix.ram_r[688] ));
 sg13g2_dfrbp_1 \logix.ram_r[689]$_DFFE_PP_  (.CLK(net621),
    .RESET_B(net2507),
    .D(_1716_),
    .Q_N(_4282_),
    .Q(\logix.ram_r[689] ));
 sg13g2_dfrbp_1 \logix.ram_r[68]$_DFFE_PP_  (.CLK(net623),
    .RESET_B(net2508),
    .D(_1717_),
    .Q_N(_4281_),
    .Q(\logix.ram_r[68] ));
 sg13g2_dfrbp_1 \logix.ram_r[690]$_DFFE_PP_  (.CLK(net616),
    .RESET_B(net2509),
    .D(_1718_),
    .Q_N(_4280_),
    .Q(\logix.ram_r[690] ));
 sg13g2_dfrbp_1 \logix.ram_r[691]$_DFFE_PP_  (.CLK(net615),
    .RESET_B(net2510),
    .D(_1719_),
    .Q_N(_4279_),
    .Q(\logix.ram_r[691] ));
 sg13g2_dfrbp_1 \logix.ram_r[692]$_DFFE_PP_  (.CLK(net616),
    .RESET_B(net2511),
    .D(_1720_),
    .Q_N(_4278_),
    .Q(\logix.ram_r[692] ));
 sg13g2_dfrbp_1 \logix.ram_r[693]$_DFFE_PP_  (.CLK(net612),
    .RESET_B(net2512),
    .D(_1721_),
    .Q_N(_4277_),
    .Q(\logix.ram_r[693] ));
 sg13g2_dfrbp_1 \logix.ram_r[694]$_DFFE_PP_  (.CLK(net612),
    .RESET_B(net2513),
    .D(_1722_),
    .Q_N(_4276_),
    .Q(\logix.ram_r[694] ));
 sg13g2_dfrbp_1 \logix.ram_r[695]$_DFFE_PP_  (.CLK(net619),
    .RESET_B(net2514),
    .D(_1723_),
    .Q_N(_4275_),
    .Q(\logix.ram_r[695] ));
 sg13g2_dfrbp_1 \logix.ram_r[696]$_DFFE_PP_  (.CLK(net619),
    .RESET_B(net2515),
    .D(_1724_),
    .Q_N(_4274_),
    .Q(\logix.ram_r[696] ));
 sg13g2_dfrbp_1 \logix.ram_r[697]$_DFFE_PP_  (.CLK(net621),
    .RESET_B(net2516),
    .D(_1725_),
    .Q_N(_4273_),
    .Q(\logix.ram_r[697] ));
 sg13g2_dfrbp_1 \logix.ram_r[698]$_DFFE_PP_  (.CLK(net621),
    .RESET_B(net2517),
    .D(_1726_),
    .Q_N(_4272_),
    .Q(\logix.ram_r[698] ));
 sg13g2_dfrbp_1 \logix.ram_r[699]$_DFFE_PP_  (.CLK(net616),
    .RESET_B(net2518),
    .D(_1727_),
    .Q_N(_4271_),
    .Q(\logix.ram_r[699] ));
 sg13g2_dfrbp_1 \logix.ram_r[69]$_DFFE_PP_  (.CLK(net623),
    .RESET_B(net2519),
    .D(_1728_),
    .Q_N(_4270_),
    .Q(\logix.ram_r[69] ));
 sg13g2_dfrbp_1 \logix.ram_r[6]$_DFFE_PP_  (.CLK(net609),
    .RESET_B(net2520),
    .D(_1729_),
    .Q_N(_4269_),
    .Q(\logix.ram_r[6] ));
 sg13g2_dfrbp_1 \logix.ram_r[700]$_DFFE_PP_  (.CLK(net616),
    .RESET_B(net2521),
    .D(_1730_),
    .Q_N(_4268_),
    .Q(\logix.ram_r[700] ));
 sg13g2_dfrbp_1 \logix.ram_r[701]$_DFFE_PP_  (.CLK(net614),
    .RESET_B(net2522),
    .D(_1731_),
    .Q_N(_4267_),
    .Q(\logix.ram_r[701] ));
 sg13g2_dfrbp_1 \logix.ram_r[702]$_DFFE_PP_  (.CLK(net614),
    .RESET_B(net2523),
    .D(_1732_),
    .Q_N(_4266_),
    .Q(\logix.ram_r[702] ));
 sg13g2_dfrbp_1 \logix.ram_r[703]$_DFFE_PP_  (.CLK(net614),
    .RESET_B(net2524),
    .D(_1733_),
    .Q_N(_4265_),
    .Q(\logix.ram_r[703] ));
 sg13g2_dfrbp_1 \logix.ram_r[704]$_DFFE_PP_  (.CLK(net613),
    .RESET_B(net2525),
    .D(_1734_),
    .Q_N(_4264_),
    .Q(\logix.ram_r[704] ));
 sg13g2_dfrbp_1 \logix.ram_r[705]$_DFFE_PP_  (.CLK(net615),
    .RESET_B(net2526),
    .D(_1735_),
    .Q_N(_4263_),
    .Q(\logix.ram_r[705] ));
 sg13g2_dfrbp_1 \logix.ram_r[706]$_DFFE_PP_  (.CLK(net599),
    .RESET_B(net2527),
    .D(_1736_),
    .Q_N(_4262_),
    .Q(\logix.ram_r[706] ));
 sg13g2_dfrbp_1 \logix.ram_r[707]$_DFFE_PP_  (.CLK(net594),
    .RESET_B(net2528),
    .D(_1737_),
    .Q_N(_4261_),
    .Q(\logix.ram_r[707] ));
 sg13g2_dfrbp_1 \logix.ram_r[708]$_DFFE_PP_  (.CLK(net594),
    .RESET_B(net2529),
    .D(_1738_),
    .Q_N(_4260_),
    .Q(\logix.ram_r[708] ));
 sg13g2_dfrbp_1 \logix.ram_r[709]$_DFFE_PP_  (.CLK(net594),
    .RESET_B(net2530),
    .D(_1739_),
    .Q_N(_4259_),
    .Q(\logix.ram_r[709] ));
 sg13g2_dfrbp_1 \logix.ram_r[70]$_DFFE_PP_  (.CLK(net607),
    .RESET_B(net2531),
    .D(_1740_),
    .Q_N(_4258_),
    .Q(\logix.ram_r[70] ));
 sg13g2_dfrbp_1 \logix.ram_r[710]$_DFFE_PP_  (.CLK(net591),
    .RESET_B(net2532),
    .D(_1741_),
    .Q_N(_4257_),
    .Q(\logix.ram_r[710] ));
 sg13g2_dfrbp_1 \logix.ram_r[711]$_DFFE_PP_  (.CLK(net598),
    .RESET_B(net2533),
    .D(_1742_),
    .Q_N(_4256_),
    .Q(\logix.ram_r[711] ));
 sg13g2_dfrbp_1 \logix.ram_r[712]$_DFFE_PP_  (.CLK(net599),
    .RESET_B(net2534),
    .D(_1743_),
    .Q_N(_4255_),
    .Q(\logix.ram_r[712] ));
 sg13g2_dfrbp_1 \logix.ram_r[713]$_DFFE_PP_  (.CLK(net599),
    .RESET_B(net2535),
    .D(_1744_),
    .Q_N(_4254_),
    .Q(\logix.ram_r[713] ));
 sg13g2_dfrbp_1 \logix.ram_r[714]$_DFFE_PP_  (.CLK(net598),
    .RESET_B(net2536),
    .D(_1745_),
    .Q_N(_4253_),
    .Q(\logix.ram_r[714] ));
 sg13g2_dfrbp_1 \logix.ram_r[715]$_DFFE_PP_  (.CLK(net594),
    .RESET_B(net2537),
    .D(_1746_),
    .Q_N(_4252_),
    .Q(\logix.ram_r[715] ));
 sg13g2_dfrbp_1 \logix.ram_r[716]$_DFFE_PP_  (.CLK(net595),
    .RESET_B(net2538),
    .D(_1747_),
    .Q_N(_4251_),
    .Q(\logix.ram_r[716] ));
 sg13g2_dfrbp_1 \logix.ram_r[717]$_DFFE_PP_  (.CLK(net595),
    .RESET_B(net2539),
    .D(_1748_),
    .Q_N(_4250_),
    .Q(\logix.ram_r[717] ));
 sg13g2_dfrbp_1 \logix.ram_r[718]$_DFFE_PP_  (.CLK(net592),
    .RESET_B(net2540),
    .D(_1749_),
    .Q_N(_4249_),
    .Q(\logix.ram_r[718] ));
 sg13g2_dfrbp_1 \logix.ram_r[719]$_DFFE_PP_  (.CLK(net596),
    .RESET_B(net2541),
    .D(_1750_),
    .Q_N(_4248_),
    .Q(\logix.ram_r[719] ));
 sg13g2_dfrbp_1 \logix.ram_r[71]$_DFFE_PP_  (.CLK(net600),
    .RESET_B(net2542),
    .D(_1751_),
    .Q_N(_4247_),
    .Q(\logix.ram_r[71] ));
 sg13g2_dfrbp_1 \logix.ram_r[720]$_DFFE_PP_  (.CLK(net599),
    .RESET_B(net2543),
    .D(_1752_),
    .Q_N(_4246_),
    .Q(\logix.ram_r[720] ));
 sg13g2_dfrbp_1 \logix.ram_r[721]$_DFFE_PP_  (.CLK(net599),
    .RESET_B(net2544),
    .D(_1753_),
    .Q_N(_4245_),
    .Q(\logix.ram_r[721] ));
 sg13g2_dfrbp_1 \logix.ram_r[722]$_DFFE_PP_  (.CLK(net600),
    .RESET_B(net2545),
    .D(_1754_),
    .Q_N(_4244_),
    .Q(\logix.ram_r[722] ));
 sg13g2_dfrbp_1 \logix.ram_r[723]$_DFFE_PP_  (.CLK(net598),
    .RESET_B(net2546),
    .D(_1755_),
    .Q_N(_4243_),
    .Q(\logix.ram_r[723] ));
 sg13g2_dfrbp_1 \logix.ram_r[724]$_DFFE_PP_  (.CLK(net595),
    .RESET_B(net2547),
    .D(_1756_),
    .Q_N(_4242_),
    .Q(\logix.ram_r[724] ));
 sg13g2_dfrbp_1 \logix.ram_r[725]$_DFFE_PP_  (.CLK(net598),
    .RESET_B(net2548),
    .D(_1757_),
    .Q_N(_4241_),
    .Q(\logix.ram_r[725] ));
 sg13g2_dfrbp_1 \logix.ram_r[726]$_DFFE_PP_  (.CLK(net598),
    .RESET_B(net2549),
    .D(_1758_),
    .Q_N(_4240_),
    .Q(\logix.ram_r[726] ));
 sg13g2_dfrbp_1 \logix.ram_r[727]$_DFFE_PP_  (.CLK(net599),
    .RESET_B(net2550),
    .D(_1759_),
    .Q_N(_4239_),
    .Q(\logix.ram_r[727] ));
 sg13g2_dfrbp_1 \logix.ram_r[728]$_DFFE_PP_  (.CLK(net599),
    .RESET_B(net2551),
    .D(_1760_),
    .Q_N(_4238_),
    .Q(\logix.ram_r[728] ));
 sg13g2_dfrbp_1 \logix.ram_r[729]$_DFFE_PP_  (.CLK(net599),
    .RESET_B(net2552),
    .D(_1761_),
    .Q_N(_4237_),
    .Q(\logix.ram_r[729] ));
 sg13g2_dfrbp_1 \logix.ram_r[72]$_DFFE_PP_  (.CLK(net615),
    .RESET_B(net2553),
    .D(_1762_),
    .Q_N(_4236_),
    .Q(\logix.ram_r[72] ));
 sg13g2_dfrbp_1 \logix.ram_r[730]$_DFFE_PP_  (.CLK(net598),
    .RESET_B(net2554),
    .D(_1763_),
    .Q_N(_4235_),
    .Q(\logix.ram_r[730] ));
 sg13g2_dfrbp_1 \logix.ram_r[731]$_DFFE_PP_  (.CLK(net598),
    .RESET_B(net2555),
    .D(_1764_),
    .Q_N(_4234_),
    .Q(\logix.ram_r[731] ));
 sg13g2_dfrbp_1 \logix.ram_r[732]$_DFFE_PP_  (.CLK(net600),
    .RESET_B(net2556),
    .D(_1765_),
    .Q_N(_4233_),
    .Q(\logix.ram_r[732] ));
 sg13g2_dfrbp_1 \logix.ram_r[733]$_DFFE_PP_  (.CLK(net598),
    .RESET_B(net2557),
    .D(_1766_),
    .Q_N(_4232_),
    .Q(\logix.ram_r[733] ));
 sg13g2_dfrbp_1 \logix.ram_r[734]$_DFFE_PP_  (.CLK(net597),
    .RESET_B(net2558),
    .D(_1767_),
    .Q_N(_4231_),
    .Q(\logix.ram_r[734] ));
 sg13g2_dfrbp_1 \logix.ram_r[735]$_DFFE_PP_  (.CLK(net596),
    .RESET_B(net2559),
    .D(_1768_),
    .Q_N(_4230_),
    .Q(\logix.ram_r[735] ));
 sg13g2_dfrbp_1 \logix.ram_r[736]$_DFFE_PP_  (.CLK(net596),
    .RESET_B(net2560),
    .D(_1769_),
    .Q_N(_4229_),
    .Q(\logix.ram_r[736] ));
 sg13g2_dfrbp_1 \logix.ram_r[737]$_DFFE_PP_  (.CLK(net596),
    .RESET_B(net2561),
    .D(_1770_),
    .Q_N(_4228_),
    .Q(\logix.ram_r[737] ));
 sg13g2_dfrbp_1 \logix.ram_r[738]$_DFFE_PP_  (.CLK(net601),
    .RESET_B(net2562),
    .D(_1771_),
    .Q_N(_4227_),
    .Q(\logix.ram_r[738] ));
 sg13g2_dfrbp_1 \logix.ram_r[739]$_DFFE_PP_  (.CLK(net592),
    .RESET_B(net2563),
    .D(_1772_),
    .Q_N(_4226_),
    .Q(\logix.ram_r[739] ));
 sg13g2_dfrbp_1 \logix.ram_r[73]$_DFFE_PP_  (.CLK(net607),
    .RESET_B(net2564),
    .D(_1773_),
    .Q_N(_4225_),
    .Q(\logix.ram_r[73] ));
 sg13g2_dfrbp_1 \logix.ram_r[740]$_DFFE_PP_  (.CLK(net591),
    .RESET_B(net2565),
    .D(_1774_),
    .Q_N(_4224_),
    .Q(\logix.ram_r[740] ));
 sg13g2_dfrbp_1 \logix.ram_r[741]$_DFFE_PP_  (.CLK(net591),
    .RESET_B(net2566),
    .D(_1775_),
    .Q_N(_4223_),
    .Q(\logix.ram_r[741] ));
 sg13g2_dfrbp_1 \logix.ram_r[742]$_DFFE_PP_  (.CLK(net597),
    .RESET_B(net2567),
    .D(_1776_),
    .Q_N(_4222_),
    .Q(\logix.ram_r[742] ));
 sg13g2_dfrbp_1 \logix.ram_r[743]$_DFFE_PP_  (.CLK(net596),
    .RESET_B(net2568),
    .D(_1777_),
    .Q_N(_4221_),
    .Q(\logix.ram_r[743] ));
 sg13g2_dfrbp_1 \logix.ram_r[744]$_DFFE_PP_  (.CLK(net596),
    .RESET_B(net2569),
    .D(_1778_),
    .Q_N(_4220_),
    .Q(\logix.ram_r[744] ));
 sg13g2_dfrbp_1 \logix.ram_r[745]$_DFFE_PP_  (.CLK(net613),
    .RESET_B(net2570),
    .D(_1779_),
    .Q_N(_4219_),
    .Q(\logix.ram_r[745] ));
 sg13g2_dfrbp_1 \logix.ram_r[746]$_DFFE_PP_  (.CLK(net613),
    .RESET_B(net2571),
    .D(_1780_),
    .Q_N(_4218_),
    .Q(\logix.ram_r[746] ));
 sg13g2_dfrbp_1 \logix.ram_r[747]$_DFFE_PP_  (.CLK(net592),
    .RESET_B(net2572),
    .D(_1781_),
    .Q_N(_4217_),
    .Q(\logix.ram_r[747] ));
 sg13g2_dfrbp_1 \logix.ram_r[748]$_DFFE_PP_  (.CLK(net591),
    .RESET_B(net2573),
    .D(_1782_),
    .Q_N(_4216_),
    .Q(\logix.ram_r[748] ));
 sg13g2_dfrbp_1 \logix.ram_r[749]$_DFFE_PP_  (.CLK(net591),
    .RESET_B(net2574),
    .D(_1783_),
    .Q_N(_4215_),
    .Q(\logix.ram_r[749] ));
 sg13g2_dfrbp_1 \logix.ram_r[74]$_DFFE_PP_  (.CLK(net608),
    .RESET_B(net2575),
    .D(_1784_),
    .Q_N(_4214_),
    .Q(\logix.ram_r[74] ));
 sg13g2_dfrbp_1 \logix.ram_r[750]$_DFFE_PP_  (.CLK(net597),
    .RESET_B(net2576),
    .D(_1785_),
    .Q_N(_4213_),
    .Q(\logix.ram_r[750] ));
 sg13g2_dfrbp_1 \logix.ram_r[751]$_DFFE_PP_  (.CLK(net596),
    .RESET_B(net2577),
    .D(_1786_),
    .Q_N(_4212_),
    .Q(\logix.ram_r[751] ));
 sg13g2_dfrbp_1 \logix.ram_r[752]$_DFFE_PP_  (.CLK(net613),
    .RESET_B(net2578),
    .D(_1787_),
    .Q_N(_4211_),
    .Q(\logix.ram_r[752] ));
 sg13g2_dfrbp_1 \logix.ram_r[753]$_DFFE_PP_  (.CLK(net613),
    .RESET_B(net2579),
    .D(_1788_),
    .Q_N(_4210_),
    .Q(\logix.ram_r[753] ));
 sg13g2_dfrbp_1 \logix.ram_r[754]$_DFFE_PP_  (.CLK(net613),
    .RESET_B(net2580),
    .D(_1789_),
    .Q_N(_4209_),
    .Q(\logix.ram_r[754] ));
 sg13g2_dfrbp_1 \logix.ram_r[755]$_DFFE_PP_  (.CLK(net592),
    .RESET_B(net2581),
    .D(_1790_),
    .Q_N(_4208_),
    .Q(\logix.ram_r[755] ));
 sg13g2_dfrbp_1 \logix.ram_r[756]$_DFFE_PP_  (.CLK(net591),
    .RESET_B(net2582),
    .D(_1791_),
    .Q_N(_4207_),
    .Q(\logix.ram_r[756] ));
 sg13g2_dfrbp_1 \logix.ram_r[757]$_DFFE_PP_  (.CLK(net591),
    .RESET_B(net2583),
    .D(_1792_),
    .Q_N(_4206_),
    .Q(\logix.ram_r[757] ));
 sg13g2_dfrbp_1 \logix.ram_r[758]$_DFFE_PP_  (.CLK(net597),
    .RESET_B(net2584),
    .D(_1793_),
    .Q_N(_4205_),
    .Q(\logix.ram_r[758] ));
 sg13g2_dfrbp_1 \logix.ram_r[759]$_DFFE_PP_  (.CLK(net596),
    .RESET_B(net2585),
    .D(_1794_),
    .Q_N(_4204_),
    .Q(\logix.ram_r[759] ));
 sg13g2_dfrbp_1 \logix.ram_r[75]$_DFFE_PP_  (.CLK(net623),
    .RESET_B(net2586),
    .D(_1795_),
    .Q_N(_4203_),
    .Q(\logix.ram_r[75] ));
 sg13g2_dfrbp_1 \logix.ram_r[760]$_DFFE_PP_  (.CLK(net613),
    .RESET_B(net2587),
    .D(_1796_),
    .Q_N(_4202_),
    .Q(\logix.ram_r[760] ));
 sg13g2_dfrbp_1 \logix.ram_r[761]$_DFFE_PP_  (.CLK(net613),
    .RESET_B(net2588),
    .D(_1797_),
    .Q_N(_4201_),
    .Q(\logix.ram_r[761] ));
 sg13g2_dfrbp_1 \logix.ram_r[762]$_DFFE_PP_  (.CLK(net597),
    .RESET_B(net2589),
    .D(_1798_),
    .Q_N(_4200_),
    .Q(\logix.ram_r[762] ));
 sg13g2_dfrbp_1 \logix.ram_r[763]$_DFFE_PP_  (.CLK(net592),
    .RESET_B(net2590),
    .D(_1799_),
    .Q_N(_4199_),
    .Q(\logix.ram_r[763] ));
 sg13g2_dfrbp_1 \logix.ram_r[764]$_DFFE_PP_  (.CLK(net591),
    .RESET_B(net2591),
    .D(_1800_),
    .Q_N(_4198_),
    .Q(\logix.ram_r[764] ));
 sg13g2_dfrbp_1 \logix.ram_r[765]$_DFFE_PP_  (.CLK(net597),
    .RESET_B(net2592),
    .D(_1801_),
    .Q_N(_4197_),
    .Q(\logix.ram_r[765] ));
 sg13g2_dfrbp_1 \logix.ram_r[766]$_DFFE_PP_  (.CLK(net597),
    .RESET_B(net2593),
    .D(_1802_),
    .Q_N(_4196_),
    .Q(\logix.ram_r[766] ));
 sg13g2_dfrbp_1 \logix.ram_r[767]$_DFFE_PP_  (.CLK(net612),
    .RESET_B(net2594),
    .D(_1803_),
    .Q_N(_4195_),
    .Q(\logix.ram_r[767] ));
 sg13g2_dfrbp_1 \logix.ram_r[768]$_DFFE_PP_  (.CLK(net733),
    .RESET_B(net2595),
    .D(_1804_),
    .Q_N(_4194_),
    .Q(\logix.ram_r[768] ));
 sg13g2_dfrbp_1 \logix.ram_r[769]$_DFFE_PP_  (.CLK(net733),
    .RESET_B(net2596),
    .D(_1805_),
    .Q_N(_4193_),
    .Q(\logix.ram_r[769] ));
 sg13g2_dfrbp_1 \logix.ram_r[76]$_DFFE_PP_  (.CLK(net623),
    .RESET_B(net2597),
    .D(_1806_),
    .Q_N(_4192_),
    .Q(\logix.ram_r[76] ));
 sg13g2_dfrbp_1 \logix.ram_r[770]$_DFFE_PP_  (.CLK(net733),
    .RESET_B(net2598),
    .D(_1807_),
    .Q_N(_4191_),
    .Q(\logix.ram_r[770] ));
 sg13g2_dfrbp_1 \logix.ram_r[771]$_DFFE_PP_  (.CLK(net751),
    .RESET_B(net2599),
    .D(_1808_),
    .Q_N(_4190_),
    .Q(\logix.ram_r[771] ));
 sg13g2_dfrbp_1 \logix.ram_r[772]$_DFFE_PP_  (.CLK(net750),
    .RESET_B(net2600),
    .D(_1809_),
    .Q_N(_4189_),
    .Q(\logix.ram_r[772] ));
 sg13g2_dfrbp_1 \logix.ram_r[773]$_DFFE_PP_  (.CLK(net758),
    .RESET_B(net2601),
    .D(_1810_),
    .Q_N(_4188_),
    .Q(\logix.ram_r[773] ));
 sg13g2_dfrbp_1 \logix.ram_r[774]$_DFFE_PP_  (.CLK(net758),
    .RESET_B(net2602),
    .D(_1811_),
    .Q_N(_4187_),
    .Q(\logix.ram_r[774] ));
 sg13g2_dfrbp_1 \logix.ram_r[775]$_DFFE_PP_  (.CLK(net758),
    .RESET_B(net2603),
    .D(_1812_),
    .Q_N(_4186_),
    .Q(\logix.ram_r[775] ));
 sg13g2_dfrbp_1 \logix.ram_r[776]$_DFFE_PP_  (.CLK(net756),
    .RESET_B(net2604),
    .D(_1813_),
    .Q_N(_4185_),
    .Q(\logix.ram_r[776] ));
 sg13g2_dfrbp_1 \logix.ram_r[777]$_DFFE_PP_  (.CLK(net756),
    .RESET_B(net2605),
    .D(_1814_),
    .Q_N(_4184_),
    .Q(\logix.ram_r[777] ));
 sg13g2_dfrbp_1 \logix.ram_r[778]$_DFFE_PP_  (.CLK(net756),
    .RESET_B(net2606),
    .D(_1815_),
    .Q_N(_4183_),
    .Q(\logix.ram_r[778] ));
 sg13g2_dfrbp_1 \logix.ram_r[779]$_DFFE_PP_  (.CLK(net757),
    .RESET_B(net2607),
    .D(_1816_),
    .Q_N(_4182_),
    .Q(\logix.ram_r[779] ));
 sg13g2_dfrbp_1 \logix.ram_r[77]$_DFFE_PP_  (.CLK(net626),
    .RESET_B(net2608),
    .D(_1817_),
    .Q_N(_4181_),
    .Q(\logix.ram_r[77] ));
 sg13g2_dfrbp_1 \logix.ram_r[780]$_DFFE_PP_  (.CLK(net750),
    .RESET_B(net2609),
    .D(_1818_),
    .Q_N(_4180_),
    .Q(\logix.ram_r[780] ));
 sg13g2_dfrbp_1 \logix.ram_r[781]$_DFFE_PP_  (.CLK(net750),
    .RESET_B(net2610),
    .D(_1819_),
    .Q_N(_4179_),
    .Q(\logix.ram_r[781] ));
 sg13g2_dfrbp_1 \logix.ram_r[782]$_DFFE_PP_  (.CLK(net762),
    .RESET_B(net2611),
    .D(_1820_),
    .Q_N(_4178_),
    .Q(\logix.ram_r[782] ));
 sg13g2_dfrbp_1 \logix.ram_r[783]$_DFFE_PP_  (.CLK(net761),
    .RESET_B(net2612),
    .D(_1821_),
    .Q_N(_4177_),
    .Q(\logix.ram_r[783] ));
 sg13g2_dfrbp_1 \logix.ram_r[784]$_DFFE_PP_  (.CLK(net742),
    .RESET_B(net2613),
    .D(_1822_),
    .Q_N(_4176_),
    .Q(\logix.ram_r[784] ));
 sg13g2_dfrbp_1 \logix.ram_r[785]$_DFFE_PP_  (.CLK(net742),
    .RESET_B(net2614),
    .D(_1823_),
    .Q_N(_4175_),
    .Q(\logix.ram_r[785] ));
 sg13g2_dfrbp_1 \logix.ram_r[786]$_DFFE_PP_  (.CLK(net735),
    .RESET_B(net2615),
    .D(_1824_),
    .Q_N(_4174_),
    .Q(\logix.ram_r[786] ));
 sg13g2_dfrbp_1 \logix.ram_r[787]$_DFFE_PP_  (.CLK(net751),
    .RESET_B(net2616),
    .D(_1825_),
    .Q_N(_4173_),
    .Q(\logix.ram_r[787] ));
 sg13g2_dfrbp_1 \logix.ram_r[788]$_DFFE_PP_  (.CLK(net750),
    .RESET_B(net2617),
    .D(_1826_),
    .Q_N(_4172_),
    .Q(\logix.ram_r[788] ));
 sg13g2_dfrbp_1 \logix.ram_r[789]$_DFFE_PP_  (.CLK(net758),
    .RESET_B(net2618),
    .D(_1827_),
    .Q_N(_4171_),
    .Q(\logix.ram_r[789] ));
 sg13g2_dfrbp_1 \logix.ram_r[78]$_DFFE_PP_  (.CLK(net626),
    .RESET_B(net2619),
    .D(_1828_),
    .Q_N(_4170_),
    .Q(\logix.ram_r[78] ));
 sg13g2_dfrbp_1 \logix.ram_r[790]$_DFFE_PP_  (.CLK(net758),
    .RESET_B(net2620),
    .D(_1829_),
    .Q_N(_4169_),
    .Q(\logix.ram_r[790] ));
 sg13g2_dfrbp_1 \logix.ram_r[791]$_DFFE_PP_  (.CLK(net757),
    .RESET_B(net2621),
    .D(_1830_),
    .Q_N(_4168_),
    .Q(\logix.ram_r[791] ));
 sg13g2_dfrbp_1 \logix.ram_r[792]$_DFFE_PP_  (.CLK(net767),
    .RESET_B(net2622),
    .D(_1831_),
    .Q_N(_4167_),
    .Q(\logix.ram_r[792] ));
 sg13g2_dfrbp_1 \logix.ram_r[793]$_DFFE_PP_  (.CLK(net767),
    .RESET_B(net2623),
    .D(_1832_),
    .Q_N(_4166_),
    .Q(\logix.ram_r[793] ));
 sg13g2_dfrbp_1 \logix.ram_r[794]$_DFFE_PP_  (.CLK(net757),
    .RESET_B(net2624),
    .D(_1833_),
    .Q_N(_4165_),
    .Q(\logix.ram_r[794] ));
 sg13g2_dfrbp_1 \logix.ram_r[795]$_DFFE_PP_  (.CLK(net757),
    .RESET_B(net2625),
    .D(_1834_),
    .Q_N(_4164_),
    .Q(\logix.ram_r[795] ));
 sg13g2_dfrbp_1 \logix.ram_r[796]$_DFFE_PP_  (.CLK(net751),
    .RESET_B(net2626),
    .D(_1835_),
    .Q_N(_4163_),
    .Q(\logix.ram_r[796] ));
 sg13g2_dfrbp_1 \logix.ram_r[797]$_DFFE_PP_  (.CLK(net751),
    .RESET_B(net2627),
    .D(_1836_),
    .Q_N(_4162_),
    .Q(\logix.ram_r[797] ));
 sg13g2_dfrbp_1 \logix.ram_r[798]$_DFFE_PP_  (.CLK(net762),
    .RESET_B(net2628),
    .D(_1837_),
    .Q_N(_4161_),
    .Q(\logix.ram_r[798] ));
 sg13g2_dfrbp_1 \logix.ram_r[799]$_DFFE_PP_  (.CLK(net761),
    .RESET_B(net2629),
    .D(_1838_),
    .Q_N(_4160_),
    .Q(\logix.ram_r[799] ));
 sg13g2_dfrbp_1 \logix.ram_r[79]$_DFFE_PP_  (.CLK(net626),
    .RESET_B(net2630),
    .D(_1839_),
    .Q_N(_4159_),
    .Q(\logix.ram_r[79] ));
 sg13g2_dfrbp_1 \logix.ram_r[7]$_DFFE_PP_  (.CLK(net610),
    .RESET_B(net2631),
    .D(_1840_),
    .Q_N(_4158_),
    .Q(\logix.ram_r[7] ));
 sg13g2_dfrbp_1 \logix.ram_r[800]$_DFFE_PP_  (.CLK(net761),
    .RESET_B(net2632),
    .D(_1841_),
    .Q_N(_4157_),
    .Q(\logix.ram_r[800] ));
 sg13g2_dfrbp_1 \logix.ram_r[801]$_DFFE_PP_  (.CLK(net742),
    .RESET_B(net2633),
    .D(_1842_),
    .Q_N(_4156_),
    .Q(\logix.ram_r[801] ));
 sg13g2_dfrbp_1 \logix.ram_r[802]$_DFFE_PP_  (.CLK(net742),
    .RESET_B(net2634),
    .D(_1843_),
    .Q_N(_4155_),
    .Q(\logix.ram_r[802] ));
 sg13g2_dfrbp_1 \logix.ram_r[803]$_DFFE_PP_  (.CLK(net761),
    .RESET_B(net2635),
    .D(_1844_),
    .Q_N(_4154_),
    .Q(\logix.ram_r[803] ));
 sg13g2_dfrbp_1 \logix.ram_r[804]$_DFFE_PP_  (.CLK(net762),
    .RESET_B(net2636),
    .D(_1845_),
    .Q_N(_4153_),
    .Q(\logix.ram_r[804] ));
 sg13g2_dfrbp_1 \logix.ram_r[805]$_DFFE_PP_  (.CLK(net762),
    .RESET_B(net2637),
    .D(_1846_),
    .Q_N(_4152_),
    .Q(\logix.ram_r[805] ));
 sg13g2_dfrbp_1 \logix.ram_r[806]$_DFFE_PP_  (.CLK(net766),
    .RESET_B(net2638),
    .D(_1847_),
    .Q_N(_4151_),
    .Q(\logix.ram_r[806] ));
 sg13g2_dfrbp_1 \logix.ram_r[807]$_DFFE_PP_  (.CLK(net766),
    .RESET_B(net2639),
    .D(_1848_),
    .Q_N(_4150_),
    .Q(\logix.ram_r[807] ));
 sg13g2_dfrbp_1 \logix.ram_r[808]$_DFFE_PP_  (.CLK(net767),
    .RESET_B(net2640),
    .D(_1849_),
    .Q_N(_4149_),
    .Q(\logix.ram_r[808] ));
 sg13g2_dfrbp_1 \logix.ram_r[809]$_DFFE_PP_  (.CLK(net767),
    .RESET_B(net2641),
    .D(_1850_),
    .Q_N(_4148_),
    .Q(\logix.ram_r[809] ));
 sg13g2_dfrbp_1 \logix.ram_r[80]$_DFFE_PP_  (.CLK(net728),
    .RESET_B(net2642),
    .D(_1851_),
    .Q_N(_4147_),
    .Q(\logix.ram_r[80] ));
 sg13g2_dfrbp_1 \logix.ram_r[810]$_DFFE_PP_  (.CLK(net767),
    .RESET_B(net2643),
    .D(_1852_),
    .Q_N(_4146_),
    .Q(\logix.ram_r[810] ));
 sg13g2_dfrbp_1 \logix.ram_r[811]$_DFFE_PP_  (.CLK(net768),
    .RESET_B(net2644),
    .D(_1853_),
    .Q_N(_4145_),
    .Q(\logix.ram_r[811] ));
 sg13g2_dfrbp_1 \logix.ram_r[812]$_DFFE_PP_  (.CLK(net766),
    .RESET_B(net2645),
    .D(_1854_),
    .Q_N(_4144_),
    .Q(\logix.ram_r[812] ));
 sg13g2_dfrbp_1 \logix.ram_r[813]$_DFFE_PP_  (.CLK(net766),
    .RESET_B(net2646),
    .D(_1855_),
    .Q_N(_4143_),
    .Q(\logix.ram_r[813] ));
 sg13g2_dfrbp_1 \logix.ram_r[814]$_DFFE_PP_  (.CLK(net762),
    .RESET_B(net2647),
    .D(_1856_),
    .Q_N(_4142_),
    .Q(\logix.ram_r[814] ));
 sg13g2_dfrbp_1 \logix.ram_r[815]$_DFFE_PP_  (.CLK(net761),
    .RESET_B(net2648),
    .D(_1857_),
    .Q_N(_4141_),
    .Q(\logix.ram_r[815] ));
 sg13g2_dfrbp_1 \logix.ram_r[816]$_DFFE_PP_  (.CLK(net761),
    .RESET_B(net2649),
    .D(_1858_),
    .Q_N(_4140_),
    .Q(\logix.ram_r[816] ));
 sg13g2_dfrbp_1 \logix.ram_r[817]$_DFFE_PP_  (.CLK(net742),
    .RESET_B(net2650),
    .D(_1859_),
    .Q_N(_4139_),
    .Q(\logix.ram_r[817] ));
 sg13g2_dfrbp_1 \logix.ram_r[818]$_DFFE_PP_  (.CLK(net742),
    .RESET_B(net2651),
    .D(_1860_),
    .Q_N(_4138_),
    .Q(\logix.ram_r[818] ));
 sg13g2_dfrbp_1 \logix.ram_r[819]$_DFFE_PP_  (.CLK(net761),
    .RESET_B(net2652),
    .D(_1861_),
    .Q_N(_4137_),
    .Q(\logix.ram_r[819] ));
 sg13g2_dfrbp_1 \logix.ram_r[81]$_DFFE_PP_  (.CLK(net729),
    .RESET_B(net2653),
    .D(_1862_),
    .Q_N(_4136_),
    .Q(\logix.ram_r[81] ));
 sg13g2_dfrbp_1 \logix.ram_r[820]$_DFFE_PP_  (.CLK(net762),
    .RESET_B(net2654),
    .D(_1863_),
    .Q_N(_4135_),
    .Q(\logix.ram_r[820] ));
 sg13g2_dfrbp_1 \logix.ram_r[821]$_DFFE_PP_  (.CLK(net766),
    .RESET_B(net2655),
    .D(_1864_),
    .Q_N(_4134_),
    .Q(\logix.ram_r[821] ));
 sg13g2_dfrbp_1 \logix.ram_r[822]$_DFFE_PP_  (.CLK(net766),
    .RESET_B(net2656),
    .D(_1865_),
    .Q_N(_4133_),
    .Q(\logix.ram_r[822] ));
 sg13g2_dfrbp_1 \logix.ram_r[823]$_DFFE_PP_  (.CLK(net766),
    .RESET_B(net2657),
    .D(_1866_),
    .Q_N(_4132_),
    .Q(\logix.ram_r[823] ));
 sg13g2_dfrbp_1 \logix.ram_r[824]$_DFFE_PP_  (.CLK(net767),
    .RESET_B(net2658),
    .D(_1867_),
    .Q_N(_4131_),
    .Q(\logix.ram_r[824] ));
 sg13g2_dfrbp_1 \logix.ram_r[825]$_DFFE_PP_  (.CLK(net767),
    .RESET_B(net2659),
    .D(_1868_),
    .Q_N(_4130_),
    .Q(\logix.ram_r[825] ));
 sg13g2_dfrbp_1 \logix.ram_r[826]$_DFFE_PP_  (.CLK(net767),
    .RESET_B(net2660),
    .D(_1869_),
    .Q_N(_4129_),
    .Q(\logix.ram_r[826] ));
 sg13g2_dfrbp_1 \logix.ram_r[827]$_DFFE_PP_  (.CLK(net768),
    .RESET_B(net2661),
    .D(_1870_),
    .Q_N(_4128_),
    .Q(\logix.ram_r[827] ));
 sg13g2_dfrbp_1 \logix.ram_r[828]$_DFFE_PP_  (.CLK(net768),
    .RESET_B(net2662),
    .D(_1871_),
    .Q_N(_4127_),
    .Q(\logix.ram_r[828] ));
 sg13g2_dfrbp_1 \logix.ram_r[829]$_DFFE_PP_  (.CLK(net768),
    .RESET_B(net2663),
    .D(_1872_),
    .Q_N(_4126_),
    .Q(\logix.ram_r[829] ));
 sg13g2_dfrbp_1 \logix.ram_r[82]$_DFFE_PP_  (.CLK(net734),
    .RESET_B(net2664),
    .D(_1873_),
    .Q_N(_4125_),
    .Q(\logix.ram_r[82] ));
 sg13g2_dfrbp_1 \logix.ram_r[830]$_DFFE_PP_  (.CLK(net766),
    .RESET_B(net2665),
    .D(_1874_),
    .Q_N(_4124_),
    .Q(\logix.ram_r[830] ));
 sg13g2_dfrbp_1 \logix.ram_r[831]$_DFFE_PP_  (.CLK(net769),
    .RESET_B(net2666),
    .D(_1875_),
    .Q_N(_4123_),
    .Q(\logix.ram_r[831] ));
 sg13g2_dfrbp_1 \logix.ram_r[832]$_DFFE_PP_  (.CLK(net768),
    .RESET_B(net2667),
    .D(_1876_),
    .Q_N(_4122_),
    .Q(\logix.ram_r[832] ));
 sg13g2_dfrbp_1 \logix.ram_r[833]$_DFFE_PP_  (.CLK(net771),
    .RESET_B(net2668),
    .D(_1877_),
    .Q_N(_4121_),
    .Q(\logix.ram_r[833] ));
 sg13g2_dfrbp_1 \logix.ram_r[834]$_DFFE_PP_  (.CLK(net771),
    .RESET_B(net2669),
    .D(_1878_),
    .Q_N(_4120_),
    .Q(\logix.ram_r[834] ));
 sg13g2_dfrbp_1 \logix.ram_r[835]$_DFFE_PP_  (.CLK(net764),
    .RESET_B(net2670),
    .D(_1879_),
    .Q_N(_4119_),
    .Q(\logix.ram_r[835] ));
 sg13g2_dfrbp_1 \logix.ram_r[836]$_DFFE_PP_  (.CLK(net763),
    .RESET_B(net2671),
    .D(_1880_),
    .Q_N(_4118_),
    .Q(\logix.ram_r[836] ));
 sg13g2_dfrbp_1 \logix.ram_r[837]$_DFFE_PP_  (.CLK(net770),
    .RESET_B(net2672),
    .D(_1881_),
    .Q_N(_4117_),
    .Q(\logix.ram_r[837] ));
 sg13g2_dfrbp_1 \logix.ram_r[838]$_DFFE_PP_  (.CLK(net770),
    .RESET_B(net2673),
    .D(_1882_),
    .Q_N(_4116_),
    .Q(\logix.ram_r[838] ));
 sg13g2_dfrbp_1 \logix.ram_r[839]$_DFFE_PP_  (.CLK(net770),
    .RESET_B(net2674),
    .D(_1883_),
    .Q_N(_4115_),
    .Q(\logix.ram_r[839] ));
 sg13g2_dfrbp_1 \logix.ram_r[83]$_DFFE_PP_  (.CLK(net734),
    .RESET_B(net2675),
    .D(_1884_),
    .Q_N(_4114_),
    .Q(\logix.ram_r[83] ));
 sg13g2_dfrbp_1 \logix.ram_r[840]$_DFFE_PP_  (.CLK(net771),
    .RESET_B(net2676),
    .D(_1885_),
    .Q_N(_4113_),
    .Q(\logix.ram_r[840] ));
 sg13g2_dfrbp_1 \logix.ram_r[841]$_DFFE_PP_  (.CLK(net772),
    .RESET_B(net2677),
    .D(_1886_),
    .Q_N(_4112_),
    .Q(\logix.ram_r[841] ));
 sg13g2_dfrbp_1 \logix.ram_r[842]$_DFFE_PP_  (.CLK(net772),
    .RESET_B(net2678),
    .D(_1887_),
    .Q_N(_4111_),
    .Q(\logix.ram_r[842] ));
 sg13g2_dfrbp_1 \logix.ram_r[843]$_DFFE_PP_  (.CLK(net763),
    .RESET_B(net2679),
    .D(_1888_),
    .Q_N(_4110_),
    .Q(\logix.ram_r[843] ));
 sg13g2_dfrbp_1 \logix.ram_r[844]$_DFFE_PP_  (.CLK(net763),
    .RESET_B(net2680),
    .D(_1889_),
    .Q_N(_4109_),
    .Q(\logix.ram_r[844] ));
 sg13g2_dfrbp_1 \logix.ram_r[845]$_DFFE_PP_  (.CLK(net770),
    .RESET_B(net2681),
    .D(_1890_),
    .Q_N(_4108_),
    .Q(\logix.ram_r[845] ));
 sg13g2_dfrbp_1 \logix.ram_r[846]$_DFFE_PP_  (.CLK(net770),
    .RESET_B(net2682),
    .D(_1891_),
    .Q_N(_4107_),
    .Q(\logix.ram_r[846] ));
 sg13g2_dfrbp_1 \logix.ram_r[847]$_DFFE_PP_  (.CLK(net772),
    .RESET_B(net2683),
    .D(_1892_),
    .Q_N(_4106_),
    .Q(\logix.ram_r[847] ));
 sg13g2_dfrbp_1 \logix.ram_r[848]$_DFFE_PP_  (.CLK(net771),
    .RESET_B(net2684),
    .D(_1893_),
    .Q_N(_4105_),
    .Q(\logix.ram_r[848] ));
 sg13g2_dfrbp_1 \logix.ram_r[849]$_DFFE_PP_  (.CLK(net771),
    .RESET_B(net2685),
    .D(_1894_),
    .Q_N(_4104_),
    .Q(\logix.ram_r[849] ));
 sg13g2_dfrbp_1 \logix.ram_r[84]$_DFFE_PP_  (.CLK(net734),
    .RESET_B(net2686),
    .D(_1895_),
    .Q_N(_4103_),
    .Q(\logix.ram_r[84] ));
 sg13g2_dfrbp_1 \logix.ram_r[850]$_DFFE_PP_  (.CLK(net772),
    .RESET_B(net2687),
    .D(_1896_),
    .Q_N(_4102_),
    .Q(\logix.ram_r[850] ));
 sg13g2_dfrbp_1 \logix.ram_r[851]$_DFFE_PP_  (.CLK(net763),
    .RESET_B(net2688),
    .D(_1897_),
    .Q_N(_4101_),
    .Q(\logix.ram_r[851] ));
 sg13g2_dfrbp_1 \logix.ram_r[852]$_DFFE_PP_  (.CLK(net763),
    .RESET_B(net2689),
    .D(_1898_),
    .Q_N(_4100_),
    .Q(\logix.ram_r[852] ));
 sg13g2_dfrbp_1 \logix.ram_r[853]$_DFFE_PP_  (.CLK(net773),
    .RESET_B(net2690),
    .D(_1899_),
    .Q_N(_4099_),
    .Q(\logix.ram_r[853] ));
 sg13g2_dfrbp_1 \logix.ram_r[854]$_DFFE_PP_  (.CLK(net773),
    .RESET_B(net2691),
    .D(_1900_),
    .Q_N(_4098_),
    .Q(\logix.ram_r[854] ));
 sg13g2_dfrbp_1 \logix.ram_r[855]$_DFFE_PP_  (.CLK(net771),
    .RESET_B(net2692),
    .D(_1901_),
    .Q_N(_4097_),
    .Q(\logix.ram_r[855] ));
 sg13g2_dfrbp_1 \logix.ram_r[856]$_DFFE_PP_  (.CLK(net771),
    .RESET_B(net2693),
    .D(_1902_),
    .Q_N(_4096_),
    .Q(\logix.ram_r[856] ));
 sg13g2_dfrbp_1 \logix.ram_r[857]$_DFFE_PP_  (.CLK(net771),
    .RESET_B(net2694),
    .D(_1903_),
    .Q_N(_4095_),
    .Q(\logix.ram_r[857] ));
 sg13g2_dfrbp_1 \logix.ram_r[858]$_DFFE_PP_  (.CLK(net772),
    .RESET_B(net2695),
    .D(_1904_),
    .Q_N(_4094_),
    .Q(\logix.ram_r[858] ));
 sg13g2_dfrbp_1 \logix.ram_r[859]$_DFFE_PP_  (.CLK(net765),
    .RESET_B(net2696),
    .D(_1905_),
    .Q_N(_4093_),
    .Q(\logix.ram_r[859] ));
 sg13g2_dfrbp_1 \logix.ram_r[85]$_DFFE_PP_  (.CLK(net734),
    .RESET_B(net2697),
    .D(_1906_),
    .Q_N(_4092_),
    .Q(\logix.ram_r[85] ));
 sg13g2_dfrbp_1 \logix.ram_r[860]$_DFFE_PP_  (.CLK(net763),
    .RESET_B(net2698),
    .D(_1907_),
    .Q_N(_4091_),
    .Q(\logix.ram_r[860] ));
 sg13g2_dfrbp_1 \logix.ram_r[861]$_DFFE_PP_  (.CLK(net773),
    .RESET_B(net2699),
    .D(_1908_),
    .Q_N(_4090_),
    .Q(\logix.ram_r[861] ));
 sg13g2_dfrbp_1 \logix.ram_r[862]$_DFFE_PP_  (.CLK(net770),
    .RESET_B(net2700),
    .D(_1909_),
    .Q_N(_4089_),
    .Q(\logix.ram_r[862] ));
 sg13g2_dfrbp_1 \logix.ram_r[863]$_DFFE_PP_  (.CLK(net770),
    .RESET_B(net2701),
    .D(_1910_),
    .Q_N(_4088_),
    .Q(\logix.ram_r[863] ));
 sg13g2_dfrbp_1 \logix.ram_r[864]$_DFFE_PP_  (.CLK(net770),
    .RESET_B(net2702),
    .D(_1911_),
    .Q_N(_4087_),
    .Q(\logix.ram_r[864] ));
 sg13g2_dfrbp_1 \logix.ram_r[865]$_DFFE_PP_  (.CLK(net763),
    .RESET_B(net2703),
    .D(_1912_),
    .Q_N(_4086_),
    .Q(\logix.ram_r[865] ));
 sg13g2_dfrbp_1 \logix.ram_r[866]$_DFFE_PP_  (.CLK(net763),
    .RESET_B(net2704),
    .D(_1913_),
    .Q_N(_4085_),
    .Q(\logix.ram_r[866] ));
 sg13g2_dfrbp_1 \logix.ram_r[867]$_DFFE_PP_  (.CLK(net744),
    .RESET_B(net2705),
    .D(_1914_),
    .Q_N(_4084_),
    .Q(\logix.ram_r[867] ));
 sg13g2_dfrbp_1 \logix.ram_r[868]$_DFFE_PP_  (.CLK(net744),
    .RESET_B(net2706),
    .D(_1915_),
    .Q_N(_4083_),
    .Q(\logix.ram_r[868] ));
 sg13g2_dfrbp_1 \logix.ram_r[869]$_DFFE_PP_  (.CLK(net745),
    .RESET_B(net2707),
    .D(_1916_),
    .Q_N(_4082_),
    .Q(\logix.ram_r[869] ));
 sg13g2_dfrbp_1 \logix.ram_r[86]$_DFFE_PP_  (.CLK(net734),
    .RESET_B(net2708),
    .D(_1917_),
    .Q_N(_4081_),
    .Q(\logix.ram_r[86] ));
 sg13g2_dfrbp_1 \logix.ram_r[870]$_DFFE_PP_  (.CLK(net745),
    .RESET_B(net2709),
    .D(_1918_),
    .Q_N(_4080_),
    .Q(\logix.ram_r[870] ));
 sg13g2_dfrbp_1 \logix.ram_r[871]$_DFFE_PP_  (.CLK(net764),
    .RESET_B(net2710),
    .D(_1919_),
    .Q_N(_4079_),
    .Q(\logix.ram_r[871] ));
 sg13g2_dfrbp_1 \logix.ram_r[872]$_DFFE_PP_  (.CLK(net764),
    .RESET_B(net2711),
    .D(_1920_),
    .Q_N(_4078_),
    .Q(\logix.ram_r[872] ));
 sg13g2_dfrbp_1 \logix.ram_r[873]$_DFFE_PP_  (.CLK(net764),
    .RESET_B(net2712),
    .D(_1921_),
    .Q_N(_4077_),
    .Q(\logix.ram_r[873] ));
 sg13g2_dfrbp_1 \logix.ram_r[874]$_DFFE_PP_  (.CLK(net745),
    .RESET_B(net2713),
    .D(_1922_),
    .Q_N(_4076_),
    .Q(\logix.ram_r[874] ));
 sg13g2_dfrbp_1 \logix.ram_r[875]$_DFFE_PP_  (.CLK(net744),
    .RESET_B(net2714),
    .D(_1923_),
    .Q_N(_4075_),
    .Q(\logix.ram_r[875] ));
 sg13g2_dfrbp_1 \logix.ram_r[876]$_DFFE_PP_  (.CLK(net745),
    .RESET_B(net2715),
    .D(_1924_),
    .Q_N(_4074_),
    .Q(\logix.ram_r[876] ));
 sg13g2_dfrbp_1 \logix.ram_r[877]$_DFFE_PP_  (.CLK(net742),
    .RESET_B(net2716),
    .D(_1925_),
    .Q_N(_4073_),
    .Q(\logix.ram_r[877] ));
 sg13g2_dfrbp_1 \logix.ram_r[878]$_DFFE_PP_  (.CLK(net742),
    .RESET_B(net2717),
    .D(_1926_),
    .Q_N(_4072_),
    .Q(\logix.ram_r[878] ));
 sg13g2_dfrbp_1 \logix.ram_r[879]$_DFFE_PP_  (.CLK(net761),
    .RESET_B(net2718),
    .D(_1927_),
    .Q_N(_4071_),
    .Q(\logix.ram_r[879] ));
 sg13g2_dfrbp_1 \logix.ram_r[87]$_DFFE_PP_  (.CLK(net734),
    .RESET_B(net2719),
    .D(_1928_),
    .Q_N(_4070_),
    .Q(\logix.ram_r[87] ));
 sg13g2_dfrbp_1 \logix.ram_r[880]$_DFFE_PP_  (.CLK(net764),
    .RESET_B(net2720),
    .D(_1929_),
    .Q_N(_4069_),
    .Q(\logix.ram_r[880] ));
 sg13g2_dfrbp_1 \logix.ram_r[881]$_DFFE_PP_  (.CLK(net764),
    .RESET_B(net2721),
    .D(_1930_),
    .Q_N(_4068_),
    .Q(\logix.ram_r[881] ));
 sg13g2_dfrbp_1 \logix.ram_r[882]$_DFFE_PP_  (.CLK(net764),
    .RESET_B(net2722),
    .D(_1931_),
    .Q_N(_4067_),
    .Q(\logix.ram_r[882] ));
 sg13g2_dfrbp_1 \logix.ram_r[883]$_DFFE_PP_  (.CLK(net744),
    .RESET_B(net2723),
    .D(_1932_),
    .Q_N(_4066_),
    .Q(\logix.ram_r[883] ));
 sg13g2_dfrbp_1 \logix.ram_r[884]$_DFFE_PP_  (.CLK(net746),
    .RESET_B(net2724),
    .D(_1933_),
    .Q_N(_4065_),
    .Q(\logix.ram_r[884] ));
 sg13g2_dfrbp_1 \logix.ram_r[885]$_DFFE_PP_  (.CLK(net745),
    .RESET_B(net2725),
    .D(_1934_),
    .Q_N(_4064_),
    .Q(\logix.ram_r[885] ));
 sg13g2_dfrbp_1 \logix.ram_r[886]$_DFFE_PP_  (.CLK(net745),
    .RESET_B(net2726),
    .D(_1935_),
    .Q_N(_4063_),
    .Q(\logix.ram_r[886] ));
 sg13g2_dfrbp_1 \logix.ram_r[887]$_DFFE_PP_  (.CLK(net764),
    .RESET_B(net2727),
    .D(_1936_),
    .Q_N(_4062_),
    .Q(\logix.ram_r[887] ));
 sg13g2_dfrbp_1 \logix.ram_r[888]$_DFFE_PP_  (.CLK(net746),
    .RESET_B(net2728),
    .D(_1937_),
    .Q_N(_4061_),
    .Q(\logix.ram_r[888] ));
 sg13g2_dfrbp_1 \logix.ram_r[889]$_DFFE_PP_  (.CLK(net745),
    .RESET_B(net2729),
    .D(_1938_),
    .Q_N(_4060_),
    .Q(\logix.ram_r[889] ));
 sg13g2_dfrbp_1 \logix.ram_r[88]$_DFFE_PP_  (.CLK(net624),
    .RESET_B(net2730),
    .D(_1939_),
    .Q_N(_4059_),
    .Q(\logix.ram_r[88] ));
 sg13g2_dfrbp_1 \logix.ram_r[890]$_DFFE_PP_  (.CLK(net745),
    .RESET_B(net2731),
    .D(_1940_),
    .Q_N(_4058_),
    .Q(\logix.ram_r[890] ));
 sg13g2_dfrbp_1 \logix.ram_r[891]$_DFFE_PP_  (.CLK(net744),
    .RESET_B(net2732),
    .D(_1941_),
    .Q_N(_4057_),
    .Q(\logix.ram_r[891] ));
 sg13g2_dfrbp_1 \logix.ram_r[892]$_DFFE_PP_  (.CLK(net744),
    .RESET_B(net2733),
    .D(_1942_),
    .Q_N(_4056_),
    .Q(\logix.ram_r[892] ));
 sg13g2_dfrbp_1 \logix.ram_r[893]$_DFFE_PP_  (.CLK(net743),
    .RESET_B(net2734),
    .D(_1943_),
    .Q_N(_4055_),
    .Q(\logix.ram_r[893] ));
 sg13g2_dfrbp_1 \logix.ram_r[894]$_DFFE_PP_  (.CLK(net743),
    .RESET_B(net2735),
    .D(_1944_),
    .Q_N(_4054_),
    .Q(\logix.ram_r[894] ));
 sg13g2_dfrbp_1 \logix.ram_r[895]$_DFFE_PP_  (.CLK(net743),
    .RESET_B(net2736),
    .D(_1945_),
    .Q_N(_4053_),
    .Q(\logix.ram_r[895] ));
 sg13g2_dfrbp_1 \logix.ram_r[896]$_DFFE_PP_  (.CLK(net743),
    .RESET_B(net2737),
    .D(_1946_),
    .Q_N(_4052_),
    .Q(\logix.ram_r[896] ));
 sg13g2_dfrbp_1 \logix.ram_r[897]$_DFFE_PP_  (.CLK(net610),
    .RESET_B(net2738),
    .D(_1947_),
    .Q_N(_4051_),
    .Q(\logix.ram_r[897] ));
 sg13g2_dfrbp_1 \logix.ram_r[898]$_DFFE_PP_  (.CLK(net610),
    .RESET_B(net2739),
    .D(_1948_),
    .Q_N(_4050_),
    .Q(\logix.ram_r[898] ));
 sg13g2_dfrbp_1 \logix.ram_r[899]$_DFFE_PP_  (.CLK(net609),
    .RESET_B(net2740),
    .D(_1949_),
    .Q_N(_4049_),
    .Q(\logix.ram_r[899] ));
 sg13g2_dfrbp_1 \logix.ram_r[89]$_DFFE_PP_  (.CLK(net623),
    .RESET_B(net2741),
    .D(_1950_),
    .Q_N(_4048_),
    .Q(\logix.ram_r[89] ));
 sg13g2_dfrbp_1 \logix.ram_r[8]$_DFFE_PP_  (.CLK(net610),
    .RESET_B(net2742),
    .D(_1951_),
    .Q_N(_4047_),
    .Q(\logix.ram_r[8] ));
 sg13g2_dfrbp_1 \logix.ram_r[900]$_DFFE_PP_  (.CLK(net605),
    .RESET_B(net2743),
    .D(_1952_),
    .Q_N(_4046_),
    .Q(\logix.ram_r[900] ));
 sg13g2_dfrbp_1 \logix.ram_r[901]$_DFFE_PP_  (.CLK(net603),
    .RESET_B(net2744),
    .D(_1953_),
    .Q_N(_4045_),
    .Q(\logix.ram_r[901] ));
 sg13g2_dfrbp_1 \logix.ram_r[902]$_DFFE_PP_  (.CLK(net603),
    .RESET_B(net2745),
    .D(_1954_),
    .Q_N(_4044_),
    .Q(\logix.ram_r[902] ));
 sg13g2_dfrbp_1 \logix.ram_r[903]$_DFFE_PP_  (.CLK(net607),
    .RESET_B(net2746),
    .D(_1955_),
    .Q_N(_4043_),
    .Q(\logix.ram_r[903] ));
 sg13g2_dfrbp_1 \logix.ram_r[904]$_DFFE_PP_  (.CLK(net607),
    .RESET_B(net2747),
    .D(_1956_),
    .Q_N(_4042_),
    .Q(\logix.ram_r[904] ));
 sg13g2_dfrbp_1 \logix.ram_r[905]$_DFFE_PP_  (.CLK(net608),
    .RESET_B(net2748),
    .D(_1957_),
    .Q_N(_4041_),
    .Q(\logix.ram_r[905] ));
 sg13g2_dfrbp_1 \logix.ram_r[906]$_DFFE_PP_  (.CLK(net609),
    .RESET_B(net2749),
    .D(_1958_),
    .Q_N(_4040_),
    .Q(\logix.ram_r[906] ));
 sg13g2_dfrbp_1 \logix.ram_r[907]$_DFFE_PP_  (.CLK(net609),
    .RESET_B(net2750),
    .D(_1959_),
    .Q_N(_4039_),
    .Q(\logix.ram_r[907] ));
 sg13g2_dfrbp_1 \logix.ram_r[908]$_DFFE_PP_  (.CLK(net605),
    .RESET_B(net2751),
    .D(_1960_),
    .Q_N(_4038_),
    .Q(\logix.ram_r[908] ));
 sg13g2_dfrbp_1 \logix.ram_r[909]$_DFFE_PP_  (.CLK(net603),
    .RESET_B(net2752),
    .D(_1961_),
    .Q_N(_4037_),
    .Q(\logix.ram_r[909] ));
 sg13g2_dfrbp_1 \logix.ram_r[90]$_DFFE_PP_  (.CLK(net623),
    .RESET_B(net2753),
    .D(_1962_),
    .Q_N(_4036_),
    .Q(\logix.ram_r[90] ));
 sg13g2_dfrbp_1 \logix.ram_r[910]$_DFFE_PP_  (.CLK(net603),
    .RESET_B(net2754),
    .D(_1963_),
    .Q_N(_4035_),
    .Q(\logix.ram_r[910] ));
 sg13g2_dfrbp_1 \logix.ram_r[911]$_DFFE_PP_  (.CLK(net607),
    .RESET_B(net2755),
    .D(_1964_),
    .Q_N(_4034_),
    .Q(\logix.ram_r[911] ));
 sg13g2_dfrbp_1 \logix.ram_r[912]$_DFFE_PP_  (.CLK(net608),
    .RESET_B(net2756),
    .D(_1965_),
    .Q_N(_4033_),
    .Q(\logix.ram_r[912] ));
 sg13g2_dfrbp_1 \logix.ram_r[913]$_DFFE_PP_  (.CLK(net608),
    .RESET_B(net2757),
    .D(_1966_),
    .Q_N(_4032_),
    .Q(\logix.ram_r[913] ));
 sg13g2_dfrbp_1 \logix.ram_r[914]$_DFFE_PP_  (.CLK(net610),
    .RESET_B(net2758),
    .D(_1967_),
    .Q_N(_4031_),
    .Q(\logix.ram_r[914] ));
 sg13g2_dfrbp_1 \logix.ram_r[915]$_DFFE_PP_  (.CLK(net609),
    .RESET_B(net2759),
    .D(_1968_),
    .Q_N(_4030_),
    .Q(\logix.ram_r[915] ));
 sg13g2_dfrbp_1 \logix.ram_r[916]$_DFFE_PP_  (.CLK(net605),
    .RESET_B(net2760),
    .D(_1969_),
    .Q_N(_4029_),
    .Q(\logix.ram_r[916] ));
 sg13g2_dfrbp_1 \logix.ram_r[917]$_DFFE_PP_  (.CLK(net603),
    .RESET_B(net2761),
    .D(_1970_),
    .Q_N(_4028_),
    .Q(\logix.ram_r[917] ));
 sg13g2_dfrbp_1 \logix.ram_r[918]$_DFFE_PP_  (.CLK(net603),
    .RESET_B(net2762),
    .D(_1971_),
    .Q_N(_4027_),
    .Q(\logix.ram_r[918] ));
 sg13g2_dfrbp_1 \logix.ram_r[919]$_DFFE_PP_  (.CLK(net607),
    .RESET_B(net2763),
    .D(_1972_),
    .Q_N(_4026_),
    .Q(\logix.ram_r[919] ));
 sg13g2_dfrbp_1 \logix.ram_r[91]$_DFFE_PP_  (.CLK(net623),
    .RESET_B(net2764),
    .D(_1973_),
    .Q_N(_4025_),
    .Q(\logix.ram_r[91] ));
 sg13g2_dfrbp_1 \logix.ram_r[920]$_DFFE_PP_  (.CLK(net608),
    .RESET_B(net2765),
    .D(_1974_),
    .Q_N(_4024_),
    .Q(\logix.ram_r[920] ));
 sg13g2_dfrbp_1 \logix.ram_r[921]$_DFFE_PP_  (.CLK(net608),
    .RESET_B(net2766),
    .D(_1975_),
    .Q_N(_4023_),
    .Q(\logix.ram_r[921] ));
 sg13g2_dfrbp_1 \logix.ram_r[922]$_DFFE_PP_  (.CLK(net610),
    .RESET_B(net2767),
    .D(_1976_),
    .Q_N(_4022_),
    .Q(\logix.ram_r[922] ));
 sg13g2_dfrbp_1 \logix.ram_r[923]$_DFFE_PP_  (.CLK(net609),
    .RESET_B(net2768),
    .D(_1977_),
    .Q_N(_4021_),
    .Q(\logix.ram_r[923] ));
 sg13g2_dfrbp_1 \logix.ram_r[924]$_DFFE_PP_  (.CLK(net605),
    .RESET_B(net2769),
    .D(_1978_),
    .Q_N(_4020_),
    .Q(\logix.ram_r[924] ));
 sg13g2_dfrbp_1 \logix.ram_r[925]$_DFFE_PP_  (.CLK(net603),
    .RESET_B(net2770),
    .D(_1979_),
    .Q_N(_4019_),
    .Q(\logix.ram_r[925] ));
 sg13g2_dfrbp_1 \logix.ram_r[926]$_DFFE_PP_  (.CLK(net607),
    .RESET_B(net2771),
    .D(_1980_),
    .Q_N(_4018_),
    .Q(\logix.ram_r[926] ));
 sg13g2_dfrbp_1 \logix.ram_r[927]$_DFFE_PP_  (.CLK(net607),
    .RESET_B(net2772),
    .D(_1981_),
    .Q_N(_4017_),
    .Q(\logix.ram_r[927] ));
 sg13g2_dfrbp_1 \logix.ram_r[928]$_DFFE_PP_  (.CLK(net602),
    .RESET_B(net2773),
    .D(_1982_),
    .Q_N(_4016_),
    .Q(\logix.ram_r[928] ));
 sg13g2_dfrbp_1 \logix.ram_r[929]$_DFFE_PP_  (.CLK(net604),
    .RESET_B(net2774),
    .D(_1983_),
    .Q_N(_4015_),
    .Q(\logix.ram_r[929] ));
 sg13g2_dfrbp_1 \logix.ram_r[92]$_DFFE_PP_  (.CLK(net623),
    .RESET_B(net2775),
    .D(_1984_),
    .Q_N(_4014_),
    .Q(\logix.ram_r[92] ));
 sg13g2_dfrbp_1 \logix.ram_r[930]$_DFFE_PP_  (.CLK(net604),
    .RESET_B(net2776),
    .D(_1985_),
    .Q_N(_4013_),
    .Q(\logix.ram_r[930] ));
 sg13g2_dfrbp_1 \logix.ram_r[931]$_DFFE_PP_  (.CLK(net602),
    .RESET_B(net2777),
    .D(_1986_),
    .Q_N(_4012_),
    .Q(\logix.ram_r[931] ));
 sg13g2_dfrbp_1 \logix.ram_r[932]$_DFFE_PP_  (.CLK(net602),
    .RESET_B(net2778),
    .D(_1987_),
    .Q_N(_4011_),
    .Q(\logix.ram_r[932] ));
 sg13g2_dfrbp_1 \logix.ram_r[933]$_DFFE_PP_  (.CLK(net602),
    .RESET_B(net2779),
    .D(_1988_),
    .Q_N(_4010_),
    .Q(\logix.ram_r[933] ));
 sg13g2_dfrbp_1 \logix.ram_r[934]$_DFFE_PP_  (.CLK(net602),
    .RESET_B(net2780),
    .D(_1989_),
    .Q_N(_4009_),
    .Q(\logix.ram_r[934] ));
 sg13g2_dfrbp_1 \logix.ram_r[935]$_DFFE_PP_  (.CLK(net594),
    .RESET_B(net2781),
    .D(_1990_),
    .Q_N(_4008_),
    .Q(\logix.ram_r[935] ));
 sg13g2_dfrbp_1 \logix.ram_r[936]$_DFFE_PP_  (.CLK(net594),
    .RESET_B(net2782),
    .D(_1991_),
    .Q_N(_4007_),
    .Q(\logix.ram_r[936] ));
 sg13g2_dfrbp_1 \logix.ram_r[937]$_DFFE_PP_  (.CLK(net594),
    .RESET_B(net2783),
    .D(_1992_),
    .Q_N(_4006_),
    .Q(\logix.ram_r[937] ));
 sg13g2_dfrbp_1 \logix.ram_r[938]$_DFFE_PP_  (.CLK(net543),
    .RESET_B(net2784),
    .D(_1993_),
    .Q_N(_4005_),
    .Q(\logix.ram_r[938] ));
 sg13g2_dfrbp_1 \logix.ram_r[939]$_DFFE_PP_  (.CLK(net543),
    .RESET_B(net2785),
    .D(_1994_),
    .Q_N(_4004_),
    .Q(\logix.ram_r[939] ));
 sg13g2_dfrbp_1 \logix.ram_r[93]$_DFFE_PP_  (.CLK(net625),
    .RESET_B(net2786),
    .D(_1995_),
    .Q_N(_4003_),
    .Q(\logix.ram_r[93] ));
 sg13g2_dfrbp_1 \logix.ram_r[940]$_DFFE_PP_  (.CLK(net543),
    .RESET_B(net2787),
    .D(_1996_),
    .Q_N(_4002_),
    .Q(\logix.ram_r[940] ));
 sg13g2_dfrbp_1 \logix.ram_r[941]$_DFFE_PP_  (.CLK(net543),
    .RESET_B(net2788),
    .D(_1997_),
    .Q_N(_4001_),
    .Q(\logix.ram_r[941] ));
 sg13g2_dfrbp_1 \logix.ram_r[942]$_DFFE_PP_  (.CLK(net545),
    .RESET_B(net2789),
    .D(_1998_),
    .Q_N(_4000_),
    .Q(\logix.ram_r[942] ));
 sg13g2_dfrbp_1 \logix.ram_r[943]$_DFFE_PP_  (.CLK(net545),
    .RESET_B(net2790),
    .D(_1999_),
    .Q_N(_3999_),
    .Q(\logix.ram_r[943] ));
 sg13g2_dfrbp_1 \logix.ram_r[944]$_DFFE_PP_  (.CLK(net545),
    .RESET_B(net2791),
    .D(_2000_),
    .Q_N(_3998_),
    .Q(\logix.ram_r[944] ));
 sg13g2_dfrbp_1 \logix.ram_r[945]$_DFFE_PP_  (.CLK(net604),
    .RESET_B(net2792),
    .D(_2001_),
    .Q_N(_3997_),
    .Q(\logix.ram_r[945] ));
 sg13g2_dfrbp_1 \logix.ram_r[946]$_DFFE_PP_  (.CLK(net546),
    .RESET_B(net2793),
    .D(_2002_),
    .Q_N(_3996_),
    .Q(\logix.ram_r[946] ));
 sg13g2_dfrbp_1 \logix.ram_r[947]$_DFFE_PP_  (.CLK(net546),
    .RESET_B(net2794),
    .D(_2003_),
    .Q_N(_3995_),
    .Q(\logix.ram_r[947] ));
 sg13g2_dfrbp_1 \logix.ram_r[948]$_DFFE_PP_  (.CLK(net602),
    .RESET_B(net2795),
    .D(_2004_),
    .Q_N(_3994_),
    .Q(\logix.ram_r[948] ));
 sg13g2_dfrbp_1 \logix.ram_r[949]$_DFFE_PP_  (.CLK(net602),
    .RESET_B(net2796),
    .D(_2005_),
    .Q_N(_3993_),
    .Q(\logix.ram_r[949] ));
 sg13g2_dfrbp_1 \logix.ram_r[94]$_DFFE_PP_  (.CLK(net625),
    .RESET_B(net2797),
    .D(_2006_),
    .Q_N(_3992_),
    .Q(\logix.ram_r[94] ));
 sg13g2_dfrbp_1 \logix.ram_r[950]$_DFFE_PP_  (.CLK(net602),
    .RESET_B(net2798),
    .D(_2007_),
    .Q_N(_3991_),
    .Q(\logix.ram_r[950] ));
 sg13g2_dfrbp_1 \logix.ram_r[951]$_DFFE_PP_  (.CLK(net603),
    .RESET_B(net2799),
    .D(_2008_),
    .Q_N(_3990_),
    .Q(\logix.ram_r[951] ));
 sg13g2_dfrbp_1 \logix.ram_r[952]$_DFFE_PP_  (.CLK(net594),
    .RESET_B(net2800),
    .D(_2009_),
    .Q_N(_3989_),
    .Q(\logix.ram_r[952] ));
 sg13g2_dfrbp_1 \logix.ram_r[953]$_DFFE_PP_  (.CLK(net544),
    .RESET_B(net2801),
    .D(_2010_),
    .Q_N(_3988_),
    .Q(\logix.ram_r[953] ));
 sg13g2_dfrbp_1 \logix.ram_r[954]$_DFFE_PP_  (.CLK(net544),
    .RESET_B(net2802),
    .D(_2011_),
    .Q_N(_3987_),
    .Q(\logix.ram_r[954] ));
 sg13g2_dfrbp_1 \logix.ram_r[955]$_DFFE_PP_  (.CLK(net544),
    .RESET_B(net2803),
    .D(_2012_),
    .Q_N(_3986_),
    .Q(\logix.ram_r[955] ));
 sg13g2_dfrbp_1 \logix.ram_r[956]$_DFFE_PP_  (.CLK(net544),
    .RESET_B(net2804),
    .D(_2013_),
    .Q_N(_3985_),
    .Q(\logix.ram_r[956] ));
 sg13g2_dfrbp_1 \logix.ram_r[957]$_DFFE_PP_  (.CLK(net543),
    .RESET_B(net2805),
    .D(_2014_),
    .Q_N(_3984_),
    .Q(\logix.ram_r[957] ));
 sg13g2_dfrbp_1 \logix.ram_r[958]$_DFFE_PP_  (.CLK(net543),
    .RESET_B(net2806),
    .D(_2015_),
    .Q_N(_3983_),
    .Q(\logix.ram_r[958] ));
 sg13g2_dfrbp_1 \logix.ram_r[959]$_DFFE_PP_  (.CLK(net546),
    .RESET_B(net2807),
    .D(_2016_),
    .Q_N(_3982_),
    .Q(\logix.ram_r[959] ));
 sg13g2_dfrbp_1 \logix.ram_r[95]$_DFFE_PP_  (.CLK(net625),
    .RESET_B(net2808),
    .D(_2017_),
    .Q_N(_3981_),
    .Q(\logix.ram_r[95] ));
 sg13g2_dfrbp_1 \logix.ram_r[960]$_DFFE_PP_  (.CLK(net546),
    .RESET_B(net2809),
    .D(_2018_),
    .Q_N(_3980_),
    .Q(\logix.ram_r[960] ));
 sg13g2_dfrbp_1 \logix.ram_r[961]$_DFFE_PP_  (.CLK(net636),
    .RESET_B(net2810),
    .D(_2019_),
    .Q_N(_3979_),
    .Q(\logix.ram_r[961] ));
 sg13g2_dfrbp_1 \logix.ram_r[962]$_DFFE_PP_  (.CLK(net634),
    .RESET_B(net2811),
    .D(_2020_),
    .Q_N(_3978_),
    .Q(\logix.ram_r[962] ));
 sg13g2_dfrbp_1 \logix.ram_r[963]$_DFFE_PP_  (.CLK(net635),
    .RESET_B(net2812),
    .D(_2021_),
    .Q_N(_3977_),
    .Q(\logix.ram_r[963] ));
 sg13g2_dfrbp_1 \logix.ram_r[964]$_DFFE_PP_  (.CLK(net635),
    .RESET_B(net2813),
    .D(_2022_),
    .Q_N(_3976_),
    .Q(\logix.ram_r[964] ));
 sg13g2_dfrbp_1 \logix.ram_r[965]$_DFFE_PP_  (.CLK(net641),
    .RESET_B(net2814),
    .D(_2023_),
    .Q_N(_3975_),
    .Q(\logix.ram_r[965] ));
 sg13g2_dfrbp_1 \logix.ram_r[966]$_DFFE_PP_  (.CLK(net641),
    .RESET_B(net2815),
    .D(_2024_),
    .Q_N(_3974_),
    .Q(\logix.ram_r[966] ));
 sg13g2_dfrbp_1 \logix.ram_r[967]$_DFFE_PP_  (.CLK(net637),
    .RESET_B(net2816),
    .D(_2025_),
    .Q_N(_3973_),
    .Q(\logix.ram_r[967] ));
 sg13g2_dfrbp_1 \logix.ram_r[968]$_DFFE_PP_  (.CLK(net636),
    .RESET_B(net2817),
    .D(_2026_),
    .Q_N(_3972_),
    .Q(\logix.ram_r[968] ));
 sg13g2_dfrbp_1 \logix.ram_r[969]$_DFFE_PP_  (.CLK(net636),
    .RESET_B(net2818),
    .D(_2027_),
    .Q_N(_3971_),
    .Q(\logix.ram_r[969] ));
 sg13g2_dfrbp_1 \logix.ram_r[96]$_DFFE_PP_  (.CLK(net625),
    .RESET_B(net2819),
    .D(_2028_),
    .Q_N(_3970_),
    .Q(\logix.ram_r[96] ));
 sg13g2_dfrbp_1 \logix.ram_r[970]$_DFFE_PP_  (.CLK(net637),
    .RESET_B(net2820),
    .D(_2029_),
    .Q_N(_3969_),
    .Q(\logix.ram_r[970] ));
 sg13g2_dfrbp_1 \logix.ram_r[971]$_DFFE_PP_  (.CLK(net635),
    .RESET_B(net2821),
    .D(_2030_),
    .Q_N(_3968_),
    .Q(\logix.ram_r[971] ));
 sg13g2_dfrbp_1 \logix.ram_r[972]$_DFFE_PP_  (.CLK(net635),
    .RESET_B(net2822),
    .D(_2031_),
    .Q_N(_3967_),
    .Q(\logix.ram_r[972] ));
 sg13g2_dfrbp_1 \logix.ram_r[973]$_DFFE_PP_  (.CLK(net637),
    .RESET_B(net2823),
    .D(_2032_),
    .Q_N(_3966_),
    .Q(\logix.ram_r[973] ));
 sg13g2_dfrbp_1 \logix.ram_r[974]$_DFFE_PP_  (.CLK(net641),
    .RESET_B(net2824),
    .D(_2033_),
    .Q_N(_3965_),
    .Q(\logix.ram_r[974] ));
 sg13g2_dfrbp_1 \logix.ram_r[975]$_DFFE_PP_  (.CLK(net637),
    .RESET_B(net2825),
    .D(_2034_),
    .Q_N(_3964_),
    .Q(\logix.ram_r[975] ));
 sg13g2_dfrbp_1 \logix.ram_r[976]$_DFFE_PP_  (.CLK(net637),
    .RESET_B(net2826),
    .D(_2035_),
    .Q_N(_3963_),
    .Q(\logix.ram_r[976] ));
 sg13g2_dfrbp_1 \logix.ram_r[977]$_DFFE_PP_  (.CLK(net636),
    .RESET_B(net2827),
    .D(_2036_),
    .Q_N(_3962_),
    .Q(\logix.ram_r[977] ));
 sg13g2_dfrbp_1 \logix.ram_r[978]$_DFFE_PP_  (.CLK(net574),
    .RESET_B(net2828),
    .D(_2037_),
    .Q_N(_3961_),
    .Q(\logix.ram_r[978] ));
 sg13g2_dfrbp_1 \logix.ram_r[979]$_DFFE_PP_  (.CLK(net575),
    .RESET_B(net2829),
    .D(_2038_),
    .Q_N(_3960_),
    .Q(\logix.ram_r[979] ));
 sg13g2_dfrbp_1 \logix.ram_r[97]$_DFFE_PP_  (.CLK(net624),
    .RESET_B(net2830),
    .D(_2039_),
    .Q_N(_3959_),
    .Q(\logix.ram_r[97] ));
 sg13g2_dfrbp_1 \logix.ram_r[980]$_DFFE_PP_  (.CLK(net575),
    .RESET_B(net2831),
    .D(_2040_),
    .Q_N(_3958_),
    .Q(\logix.ram_r[980] ));
 sg13g2_dfrbp_1 \logix.ram_r[981]$_DFFE_PP_  (.CLK(net574),
    .RESET_B(net2832),
    .D(_2041_),
    .Q_N(_3957_),
    .Q(\logix.ram_r[981] ));
 sg13g2_dfrbp_1 \logix.ram_r[982]$_DFFE_PP_  (.CLK(net571),
    .RESET_B(net2833),
    .D(_2042_),
    .Q_N(_3956_),
    .Q(\logix.ram_r[982] ));
 sg13g2_dfrbp_1 \logix.ram_r[983]$_DFFE_PP_  (.CLK(net573),
    .RESET_B(net2834),
    .D(_2043_),
    .Q_N(_3955_),
    .Q(\logix.ram_r[983] ));
 sg13g2_dfrbp_1 \logix.ram_r[984]$_DFFE_PP_  (.CLK(net576),
    .RESET_B(net2835),
    .D(_2044_),
    .Q_N(_3954_),
    .Q(\logix.ram_r[984] ));
 sg13g2_dfrbp_1 \logix.ram_r[985]$_DFFE_PP_  (.CLK(net574),
    .RESET_B(net2836),
    .D(_2045_),
    .Q_N(_3953_),
    .Q(\logix.ram_r[985] ));
 sg13g2_dfrbp_1 \logix.ram_r[986]$_DFFE_PP_  (.CLK(net574),
    .RESET_B(net2837),
    .D(_2046_),
    .Q_N(_3952_),
    .Q(\logix.ram_r[986] ));
 sg13g2_dfrbp_1 \logix.ram_r[987]$_DFFE_PP_  (.CLK(net575),
    .RESET_B(net2838),
    .D(_2047_),
    .Q_N(_3951_),
    .Q(\logix.ram_r[987] ));
 sg13g2_dfrbp_1 \logix.ram_r[988]$_DFFE_PP_  (.CLK(net575),
    .RESET_B(net2839),
    .D(_2048_),
    .Q_N(_3950_),
    .Q(\logix.ram_r[988] ));
 sg13g2_dfrbp_1 \logix.ram_r[989]$_DFFE_PP_  (.CLK(net574),
    .RESET_B(net2840),
    .D(_2049_),
    .Q_N(_3949_),
    .Q(\logix.ram_r[989] ));
 sg13g2_dfrbp_1 \logix.ram_r[98]$_DFFE_PP_  (.CLK(net693),
    .RESET_B(net2841),
    .D(_2050_),
    .Q_N(_3948_),
    .Q(\logix.ram_r[98] ));
 sg13g2_dfrbp_1 \logix.ram_r[990]$_DFFE_PP_  (.CLK(net571),
    .RESET_B(net2842),
    .D(_2051_),
    .Q_N(_3947_),
    .Q(\logix.ram_r[990] ));
 sg13g2_dfrbp_1 \logix.ram_r[991]$_DFFE_PP_  (.CLK(net573),
    .RESET_B(net2843),
    .D(_2052_),
    .Q_N(_3946_),
    .Q(\logix.ram_r[991] ));
 sg13g2_dfrbp_1 \logix.ram_r[992]$_DFFE_PP_  (.CLK(net573),
    .RESET_B(net2844),
    .D(_2053_),
    .Q_N(_3945_),
    .Q(\logix.ram_r[992] ));
 sg13g2_dfrbp_1 \logix.ram_r[993]$_DFFE_PP_  (.CLK(net576),
    .RESET_B(net2845),
    .D(_2054_),
    .Q_N(_3944_),
    .Q(\logix.ram_r[993] ));
 sg13g2_dfrbp_1 \logix.ram_r[994]$_DFFE_PP_  (.CLK(net575),
    .RESET_B(net2846),
    .D(_2055_),
    .Q_N(_3943_),
    .Q(\logix.ram_r[994] ));
 sg13g2_dfrbp_1 \logix.ram_r[995]$_DFFE_PP_  (.CLK(net575),
    .RESET_B(net2847),
    .D(_2056_),
    .Q_N(_3942_),
    .Q(\logix.ram_r[995] ));
 sg13g2_dfrbp_1 \logix.ram_r[996]$_DFFE_PP_  (.CLK(net634),
    .RESET_B(net2848),
    .D(_2057_),
    .Q_N(_3941_),
    .Q(\logix.ram_r[996] ));
 sg13g2_dfrbp_1 \logix.ram_r[997]$_DFFE_PP_  (.CLK(net634),
    .RESET_B(net2849),
    .D(_2058_),
    .Q_N(_3940_),
    .Q(\logix.ram_r[997] ));
 sg13g2_dfrbp_1 \logix.ram_r[998]$_DFFE_PP_  (.CLK(net577),
    .RESET_B(net2850),
    .D(_2059_),
    .Q_N(_3939_),
    .Q(\logix.ram_r[998] ));
 sg13g2_dfrbp_1 \logix.ram_r[999]$_DFFE_PP_  (.CLK(net577),
    .RESET_B(net2851),
    .D(_2060_),
    .Q_N(_3938_),
    .Q(\logix.ram_r[999] ));
 sg13g2_dfrbp_1 \logix.ram_r[99]$_DFFE_PP_  (.CLK(net696),
    .RESET_B(net2852),
    .D(_2061_),
    .Q_N(_3937_),
    .Q(\logix.ram_r[99] ));
 sg13g2_dfrbp_1 \logix.ram_r[9]$_DFFE_PP_  (.CLK(net657),
    .RESET_B(net2853),
    .D(_2062_),
    .Q_N(_3936_),
    .Q(\logix.ram_r[9] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[5]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[6]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[7]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[2]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[3]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[4]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[5]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[6]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout22 (.X(net22),
    .A(_3051_));
 sg13g2_buf_2 fanout23 (.A(_3048_),
    .X(net23));
 sg13g2_buf_4 fanout24 (.X(net24),
    .A(_2742_));
 sg13g2_buf_4 fanout25 (.X(net25),
    .A(_2715_));
 sg13g2_buf_4 fanout26 (.X(net26),
    .A(_2700_));
 sg13g2_buf_2 fanout27 (.A(_2696_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_2684_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_2678_),
    .X(net29));
 sg13g2_buf_4 fanout30 (.X(net30),
    .A(_2661_));
 sg13g2_buf_2 fanout31 (.A(_2658_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_2624_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_2621_),
    .X(net33));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(_2619_));
 sg13g2_buf_2 fanout35 (.A(_2614_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_2554_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_2520_),
    .X(net37));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(_2492_));
 sg13g2_buf_2 fanout39 (.A(_2488_),
    .X(net39));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(_2467_));
 sg13g2_buf_2 fanout41 (.A(_2461_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_2440_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_2434_),
    .X(net43));
 sg13g2_buf_4 fanout44 (.X(net44),
    .A(_2421_));
 sg13g2_buf_4 fanout45 (.X(net45),
    .A(_2396_));
 sg13g2_buf_2 fanout46 (.A(_2390_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_2383_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2373_),
    .X(net48));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(_3032_));
 sg13g2_buf_2 fanout50 (.A(_3010_),
    .X(net50));
 sg13g2_buf_4 fanout51 (.X(net51),
    .A(_2997_));
 sg13g2_buf_4 fanout52 (.X(net52),
    .A(_2986_));
 sg13g2_buf_2 fanout53 (.A(_2973_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2967_),
    .X(net54));
 sg13g2_buf_4 fanout55 (.X(net55),
    .A(_2959_));
 sg13g2_buf_2 fanout56 (.A(_2955_),
    .X(net56));
 sg13g2_buf_4 fanout57 (.X(net57),
    .A(_2935_));
 sg13g2_buf_2 fanout58 (.A(_2900_),
    .X(net58));
 sg13g2_buf_4 fanout59 (.X(net59),
    .A(_2687_));
 sg13g2_buf_2 fanout60 (.A(_2681_),
    .X(net60));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(_2667_));
 sg13g2_buf_2 fanout62 (.A(_2663_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_2649_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_2641_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_2594_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_2582_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_2570_),
    .X(net67));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(_2568_));
 sg13g2_buf_2 fanout69 (.A(_2561_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_2547_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_2503_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_2499_));
 sg13g2_buf_2 fanout73 (.A(_2494_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2486_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_2482_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_2473_),
    .X(net76));
 sg13g2_buf_4 fanout77 (.X(net77),
    .A(_2466_));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(_2460_));
 sg13g2_buf_2 fanout79 (.A(_2445_),
    .X(net79));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_2420_));
 sg13g2_buf_2 fanout81 (.A(_2408_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_2353_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_2345_),
    .X(net83));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(_3056_));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_3053_));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(_3014_));
 sg13g2_buf_8 fanout87 (.A(_3013_),
    .X(net87));
 sg13g2_buf_8 fanout88 (.A(_2985_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_2984_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_2980_),
    .X(net90));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(_2965_));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(_2963_));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(_2938_));
 sg13g2_buf_8 fanout94 (.A(_2910_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_2879_),
    .X(net95));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(_2847_));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(_2808_));
 sg13g2_buf_2 fanout98 (.A(_2789_),
    .X(net98));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(_2785_));
 sg13g2_buf_8 fanout100 (.A(_2782_),
    .X(net100));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(_2758_));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(_2750_));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(_2744_));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(_2733_));
 sg13g2_buf_8 fanout105 (.A(_2721_),
    .X(net105));
 sg13g2_buf_8 fanout106 (.A(_2712_),
    .X(net106));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(_2702_));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(_2686_));
 sg13g2_buf_8 fanout109 (.A(_2664_),
    .X(net109));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_2654_));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(_2650_));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(_2648_));
 sg13g2_buf_2 fanout113 (.A(_2643_),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(_2640_));
 sg13g2_buf_8 fanout115 (.A(_2634_),
    .X(net115));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_2631_));
 sg13g2_buf_8 fanout117 (.A(_2630_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_2629_),
    .X(net118));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(_2616_));
 sg13g2_buf_2 fanout120 (.A(_2612_),
    .X(net120));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(_2609_));
 sg13g2_buf_8 fanout122 (.A(_2608_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_2605_),
    .X(net123));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(_2597_));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(_2595_));
 sg13g2_buf_2 fanout126 (.A(_2593_),
    .X(net126));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_2590_));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(_2588_));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(_2586_));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_2579_));
 sg13g2_buf_8 fanout131 (.A(_2577_),
    .X(net131));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(_2574_));
 sg13g2_buf_8 fanout133 (.A(_2573_),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(_2566_),
    .X(net134));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(_2564_));
 sg13g2_buf_8 fanout136 (.A(_2563_),
    .X(net136));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(_2558_));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(_2556_));
 sg13g2_buf_8 fanout139 (.A(_2555_),
    .X(net139));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(_2543_));
 sg13g2_buf_8 fanout141 (.A(_2540_),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(_2537_));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(_2534_));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(_2528_));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(_2524_));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(_2521_));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(_2512_));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(_2509_));
 sg13g2_buf_8 fanout149 (.A(_2508_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_2507_),
    .X(net150));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(_2497_));
 sg13g2_buf_8 fanout152 (.A(_2496_),
    .X(net152));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(_2489_));
 sg13g2_buf_2 fanout154 (.A(_2481_),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(_2477_),
    .X(net155));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(_2475_));
 sg13g2_buf_8 fanout157 (.A(_2474_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_2472_),
    .X(net158));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(_2469_));
 sg13g2_buf_8 fanout160 (.A(_2468_),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(_2463_),
    .X(net161));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(_2435_));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(_2427_));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(_2425_));
 sg13g2_buf_2 fanout165 (.A(_2423_),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(_2419_),
    .X(net166));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(_2417_));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(_2413_));
 sg13g2_buf_2 fanout169 (.A(_2412_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_2407_),
    .X(net170));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(_2392_));
 sg13g2_buf_8 fanout172 (.A(_2385_),
    .X(net172));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(_2375_));
 sg13g2_buf_2 fanout174 (.A(_2363_),
    .X(net174));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(_2355_));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(_2347_));
 sg13g2_buf_4 fanout177 (.X(net177),
    .A(_2338_));
 sg13g2_buf_8 fanout178 (.A(_2332_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_2327_),
    .X(net179));
 sg13g2_buf_8 fanout180 (.A(_2992_),
    .X(net180));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(_2990_));
 sg13g2_buf_8 fanout182 (.A(_2962_),
    .X(net182));
 sg13g2_buf_8 fanout183 (.A(_2957_),
    .X(net183));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(_2941_));
 sg13g2_buf_8 fanout185 (.A(_2937_),
    .X(net185));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(_2917_));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(_2800_));
 sg13g2_buf_2 fanout188 (.A(_2781_),
    .X(net188));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(_2736_));
 sg13g2_buf_4 fanout190 (.X(net190),
    .A(_2642_));
 sg13g2_buf_4 fanout191 (.X(net191),
    .A(_2615_));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(_2596_));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(_2587_));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(_2535_));
 sg13g2_buf_8 fanout195 (.A(_2527_),
    .X(net195));
 sg13g2_buf_8 fanout196 (.A(_2523_),
    .X(net196));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(_2516_));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(_2424_));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(_2414_));
 sg13g2_buf_8 fanout200 (.A(_2391_),
    .X(net200));
 sg13g2_buf_8 fanout201 (.A(_2384_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_2380_),
    .X(net202));
 sg13g2_buf_8 fanout203 (.A(_2374_),
    .X(net203));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(_2326_));
 sg13g2_buf_2 fanout205 (.A(_2978_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_2977_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_2378_),
    .X(net207));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(_2086_));
 sg13g2_buf_4 fanout209 (.X(net209),
    .A(_2085_));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(_2084_));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(_2083_));
 sg13g2_buf_4 fanout212 (.X(net212),
    .A(_2082_));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(_2081_));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(_2080_));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(_2078_));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(_2077_));
 sg13g2_buf_4 fanout217 (.X(net217),
    .A(_2076_));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(_2075_));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(_2074_));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(_2073_));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(_2072_));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(_2310_));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(_2309_));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(_2308_));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(_2307_));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(_2306_));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(_2305_));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(_2304_));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(_2303_));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(_2302_));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(_2301_));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(_2300_));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(_2299_));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(_2297_));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(_2296_));
 sg13g2_buf_4 fanout236 (.X(net236),
    .A(_2295_));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(_2294_));
 sg13g2_buf_4 fanout238 (.X(net238),
    .A(_2293_));
 sg13g2_buf_4 fanout239 (.X(net239),
    .A(_2292_));
 sg13g2_buf_4 fanout240 (.X(net240),
    .A(_2291_));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(_2289_));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(_2288_));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(_2287_));
 sg13g2_buf_4 fanout244 (.X(net244),
    .A(_2286_));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(_2285_));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(_2284_));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(_2283_));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(_2281_));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(_2280_));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(_2279_));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(_2278_));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(_2277_));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(_2276_));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(_2275_));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(_2273_));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(_2272_));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_2271_));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(_2270_));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(_2269_));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(_2268_));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_2267_));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(_2265_));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_2264_));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_2263_));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_2262_));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_2261_));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_2260_));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_2259_));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_2257_));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(_2256_));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_2255_));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(_2254_));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_2253_));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_2252_));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(_2251_));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(_2249_));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(_2248_));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(_2247_));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(_2246_));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(_2245_));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(_2244_));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(_2243_));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_2241_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_2240_));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_2239_));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(_2238_));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_2237_));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(_2236_));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(_2235_));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(_2233_));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(_2232_));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(_2231_));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(_2230_));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(_2229_));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(_2228_));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(_2227_));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(_2225_));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(_2224_));
 sg13g2_buf_4 fanout299 (.X(net299),
    .A(_2223_));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(_2222_));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(_2221_));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(_2220_));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(_2219_));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(_2217_));
 sg13g2_buf_4 fanout305 (.X(net305),
    .A(_2216_));
 sg13g2_buf_4 fanout306 (.X(net306),
    .A(_2215_));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(_2214_));
 sg13g2_buf_4 fanout308 (.X(net308),
    .A(_2213_));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(_2210_));
 sg13g2_buf_4 fanout310 (.X(net310),
    .A(_2203_));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(_2200_));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(_2199_));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(_2198_));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(_2197_));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(_2196_));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(_2195_));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(_2194_));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(_2192_));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(_2191_));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(_2190_));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(_2189_));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_2188_));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_2187_));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(_2186_));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_2184_));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_2183_));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(_2182_));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_2181_));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_2180_));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(_2179_));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(_2178_));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(_2176_));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_2175_));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(_2174_));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(_2173_));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(_2172_));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(_2171_));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(_2170_));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(_2168_));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(_2167_));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(_2166_));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(_2165_));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(_2164_));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(_2163_));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(_2162_));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(_2160_));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_2159_));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(_2158_));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(_2157_));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(_2156_));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(_2155_));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(_2154_));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(_2152_));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(_2151_));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(_2150_));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(_2149_));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(_2148_));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(_2147_));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(_2146_));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(_2143_));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(_2142_));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(_2141_));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(_2140_));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(_2139_));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(_2138_));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(_2137_));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(_2135_));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(_2134_));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(_2133_));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(_2132_));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(_2131_));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(_2130_));
 sg13g2_buf_4 fanout373 (.X(net373),
    .A(_2129_));
 sg13g2_buf_4 fanout374 (.X(net374),
    .A(_2127_));
 sg13g2_buf_4 fanout375 (.X(net375),
    .A(_2126_));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(_2125_));
 sg13g2_buf_4 fanout377 (.X(net377),
    .A(_2124_));
 sg13g2_buf_4 fanout378 (.X(net378),
    .A(_2123_));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(_2122_));
 sg13g2_buf_4 fanout380 (.X(net380),
    .A(_2121_));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(_2119_));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(_2118_));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(_2117_));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(_2116_));
 sg13g2_buf_4 fanout385 (.X(net385),
    .A(_2115_));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(_2114_));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(_2113_));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(_2111_));
 sg13g2_buf_4 fanout389 (.X(net389),
    .A(_2110_));
 sg13g2_buf_4 fanout390 (.X(net390),
    .A(_2109_));
 sg13g2_buf_4 fanout391 (.X(net391),
    .A(_2108_));
 sg13g2_buf_4 fanout392 (.X(net392),
    .A(_2107_));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(_2106_));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(_2105_));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(_2103_));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(_2102_));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_2101_));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(_2100_));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(_2099_));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(_2098_));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(_2097_));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(_2095_));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(_2094_));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(_2093_));
 sg13g2_buf_4 fanout405 (.X(net405),
    .A(_2092_));
 sg13g2_buf_4 fanout406 (.X(net406),
    .A(_2091_));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(_2090_));
 sg13g2_buf_4 fanout408 (.X(net408),
    .A(_2089_));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(_2069_));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(_2068_));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(_2067_));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_2066_));
 sg13g2_buf_2 fanout413 (.A(_2065_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(net417),
    .X(net414));
 sg13g2_buf_1 fanout415 (.A(net417),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(net417),
    .X(net416));
 sg13g2_buf_1 fanout417 (.A(net420),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(net419),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_1 fanout420 (.A(net438),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(net425),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(net425),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(net425),
    .X(net424));
 sg13g2_buf_1 fanout425 (.A(net438),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(net428),
    .X(net426));
 sg13g2_buf_1 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(net432),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(net431),
    .X(net429));
 sg13g2_buf_1 fanout430 (.A(net431),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_1 fanout432 (.A(net438),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(net437),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(net436),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_1 fanout437 (.A(net438),
    .X(net437));
 sg13g2_buf_1 fanout438 (.A(net461),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(net441),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(net441),
    .X(net440));
 sg13g2_buf_1 fanout441 (.A(net450),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(net444),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(net450),
    .X(net443));
 sg13g2_buf_1 fanout444 (.A(net450),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(net447),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_1 fanout447 (.A(net450),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net450),
    .X(net448));
 sg13g2_buf_1 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_1 fanout450 (.A(net461),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_1 fanout452 (.A(net455),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_1 fanout455 (.A(net461),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(net460),
    .X(net456));
 sg13g2_buf_1 fanout457 (.A(net460),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(net460),
    .X(net458));
 sg13g2_buf_1 fanout459 (.A(net460),
    .X(net459));
 sg13g2_buf_1 fanout460 (.A(net461),
    .X(net460));
 sg13g2_buf_1 fanout461 (.A(net506),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(net464),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_1 fanout464 (.A(net472),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(net466),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net472),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(net471),
    .X(net467));
 sg13g2_buf_1 fanout468 (.A(net471),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(net471),
    .X(net470));
 sg13g2_buf_1 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_1 fanout472 (.A(net506),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(net475),
    .X(net473));
 sg13g2_buf_1 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_1 fanout475 (.A(net479),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(net478),
    .X(net476));
 sg13g2_buf_1 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_1 fanout479 (.A(net485),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(net485),
    .X(net480));
 sg13g2_buf_1 fanout481 (.A(net485),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net484),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(net484),
    .X(net483));
 sg13g2_buf_1 fanout484 (.A(net485),
    .X(net484));
 sg13g2_buf_1 fanout485 (.A(net506),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(net487),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(net490),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(net490),
    .X(net489));
 sg13g2_buf_1 fanout490 (.A(net505),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(net494),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(net494),
    .X(net492));
 sg13g2_buf_1 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_1 fanout494 (.A(net505),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net499),
    .X(net495));
 sg13g2_buf_1 fanout496 (.A(net499),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net499),
    .X(net497));
 sg13g2_buf_1 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_1 fanout499 (.A(net505),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net502),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(net502),
    .X(net501));
 sg13g2_buf_1 fanout502 (.A(net505),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(net505),
    .X(net504));
 sg13g2_buf_1 fanout505 (.A(net506),
    .X(net505));
 sg13g2_buf_1 fanout506 (.A(net776),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net511),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net511),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(net511),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net517),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(net514),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_1 fanout514 (.A(net517),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(net517),
    .X(net515));
 sg13g2_buf_1 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_1 fanout517 (.A(net549),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(net522),
    .X(net518));
 sg13g2_buf_1 fanout519 (.A(net522),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(net521),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_1 fanout522 (.A(net549),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(net527),
    .X(net523));
 sg13g2_buf_1 fanout524 (.A(net527),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(net527),
    .X(net525));
 sg13g2_buf_1 fanout526 (.A(net527),
    .X(net526));
 sg13g2_buf_1 fanout527 (.A(net549),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net532),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(net532),
    .X(net530));
 sg13g2_buf_1 fanout531 (.A(net532),
    .X(net531));
 sg13g2_buf_1 fanout532 (.A(net548),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net535),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_1 fanout535 (.A(net548),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_1 fanout537 (.A(net548),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(net539),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(net542),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net542),
    .X(net540));
 sg13g2_buf_1 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_1 fanout542 (.A(net548),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net547),
    .X(net543));
 sg13g2_buf_1 fanout544 (.A(net547),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net547),
    .X(net545));
 sg13g2_buf_1 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_1 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_1 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_1 fanout549 (.A(net590),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net554),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net554),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_1 fanout554 (.A(net569),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(net556),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net558),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net569),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(net563),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net563),
    .X(net560));
 sg13g2_buf_1 fanout561 (.A(net563),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net563),
    .X(net562));
 sg13g2_buf_1 fanout563 (.A(net569),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net568),
    .X(net564));
 sg13g2_buf_1 fanout565 (.A(net568),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net568),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_1 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_1 fanout569 (.A(net590),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(net579),
    .X(net570));
 sg13g2_buf_1 fanout571 (.A(net579),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net579),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net578),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net578),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net578),
    .X(net576));
 sg13g2_buf_1 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_1 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_1 fanout579 (.A(net590),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net589),
    .X(net580));
 sg13g2_buf_1 fanout581 (.A(net589),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(net589),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net588),
    .X(net584));
 sg13g2_buf_1 fanout585 (.A(net588),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_1 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_1 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_1 fanout590 (.A(net776),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(net593),
    .X(net591));
 sg13g2_buf_1 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_1 fanout593 (.A(net595),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_1 fanout595 (.A(net601),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(net601),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net600),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_1 fanout600 (.A(net601),
    .X(net600));
 sg13g2_buf_1 fanout601 (.A(net633),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net606),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(net606),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(net606),
    .X(net604));
 sg13g2_buf_1 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_1 fanout606 (.A(net633),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(net611),
    .X(net607));
 sg13g2_buf_1 fanout608 (.A(net611),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(net611),
    .X(net609));
 sg13g2_buf_1 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_1 fanout611 (.A(net633),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(net614),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net617),
    .X(net613));
 sg13g2_buf_1 fanout614 (.A(net617),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net617),
    .X(net615));
 sg13g2_buf_1 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_1 fanout617 (.A(net633),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net622),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(net622),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_1 fanout622 (.A(net633),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(net627),
    .X(net623));
 sg13g2_buf_1 fanout624 (.A(net627),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(net627),
    .X(net625));
 sg13g2_buf_1 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_1 fanout627 (.A(net632),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(net632),
    .X(net628));
 sg13g2_buf_1 fanout629 (.A(net632),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(net632),
    .X(net631));
 sg13g2_buf_1 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_1 fanout633 (.A(net776),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net638),
    .X(net634));
 sg13g2_buf_1 fanout635 (.A(net638),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net638),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_1 fanout638 (.A(net644),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(net644),
    .X(net639));
 sg13g2_buf_1 fanout640 (.A(net644),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(net643),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_1 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_1 fanout644 (.A(net679),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(net650),
    .X(net645));
 sg13g2_buf_1 fanout646 (.A(net650),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(net650),
    .X(net648));
 sg13g2_buf_1 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_1 fanout650 (.A(net679),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(net656),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(net656),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(net655),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(net655),
    .X(net654));
 sg13g2_buf_1 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_1 fanout656 (.A(net679),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(net661),
    .X(net657));
 sg13g2_buf_1 fanout658 (.A(net661),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(net661),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_1 fanout661 (.A(net667),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(net667),
    .X(net662));
 sg13g2_buf_1 fanout663 (.A(net667),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net666),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net666),
    .X(net665));
 sg13g2_buf_1 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_1 fanout667 (.A(net679),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(net678),
    .X(net668));
 sg13g2_buf_1 fanout669 (.A(net678),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(net672),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_1 fanout672 (.A(net678),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(net677),
    .X(net673));
 sg13g2_buf_1 fanout674 (.A(net677),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(net677),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_1 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_1 fanout678 (.A(net679),
    .X(net678));
 sg13g2_buf_1 fanout679 (.A(net776),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(net682),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_1 fanout682 (.A(net685),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(net684),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(net685),
    .X(net684));
 sg13g2_buf_1 fanout685 (.A(net702),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(net688),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(net688),
    .X(net687));
 sg13g2_buf_1 fanout688 (.A(net691),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_1 fanout691 (.A(net702),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(net696),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(net696),
    .X(net694));
 sg13g2_buf_1 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_1 fanout696 (.A(net702),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net701),
    .X(net697));
 sg13g2_buf_1 fanout698 (.A(net701),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(net701),
    .X(net699));
 sg13g2_buf_1 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_1 fanout701 (.A(net702),
    .X(net701));
 sg13g2_buf_1 fanout702 (.A(net775),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net705),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_1 fanout705 (.A(net714),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(net714),
    .X(net706));
 sg13g2_buf_1 fanout707 (.A(net714),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(net709),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(net713),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(net712),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(net712),
    .X(net711));
 sg13g2_buf_1 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_1 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_1 fanout714 (.A(net775),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(net725),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(net725),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(net722),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net722),
    .X(net720));
 sg13g2_buf_1 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_1 fanout722 (.A(net725),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(net725),
    .X(net724));
 sg13g2_buf_1 fanout725 (.A(net775),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(net730),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(net729),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net730),
    .X(net729));
 sg13g2_buf_1 fanout730 (.A(net747),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(net732),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net735),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(net735),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(net735),
    .X(net734));
 sg13g2_buf_1 fanout735 (.A(net747),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(net738),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(net741),
    .X(net737));
 sg13g2_buf_1 fanout738 (.A(net741),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(net740),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(net741),
    .X(net740));
 sg13g2_buf_1 fanout741 (.A(net747),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_1 fanout743 (.A(net747),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(net746),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_1 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_1 fanout747 (.A(net775),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(net760),
    .X(net748));
 sg13g2_buf_1 fanout749 (.A(net760),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(net751),
    .X(net750));
 sg13g2_buf_1 fanout751 (.A(net760),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(net755),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(net755),
    .X(net753));
 sg13g2_buf_1 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_1 fanout755 (.A(net759),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(net759),
    .X(net756));
 sg13g2_buf_1 fanout757 (.A(net759),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_1 fanout759 (.A(net760),
    .X(net759));
 sg13g2_buf_1 fanout760 (.A(net774),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(net765),
    .X(net761));
 sg13g2_buf_1 fanout762 (.A(net765),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net765),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_1 fanout765 (.A(net774),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(net769),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(net769),
    .X(net767));
 sg13g2_buf_1 fanout768 (.A(net769),
    .X(net768));
 sg13g2_buf_1 fanout769 (.A(net774),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(net773),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(net773),
    .X(net771));
 sg13g2_buf_1 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_1 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_1 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_1 fanout775 (.A(net776),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(net9),
    .X(net776));
 sg13g2_tielo _9937__777 (.L_LO(net777));
 sg13g2_tielo _9938__778 (.L_LO(net778));
 sg13g2_tielo _9939__779 (.L_LO(net779));
 sg13g2_tielo _9940__780 (.L_LO(net780));
 sg13g2_tielo _9941__781 (.L_LO(net781));
 sg13g2_tielo _9945__782 (.L_LO(net782));
 sg13g2_tielo _9946__783 (.L_LO(net783));
 sg13g2_tielo _9947__784 (.L_LO(net784));
 sg13g2_tielo _9948__785 (.L_LO(net785));
 sg13g2_tielo _9949__786 (.L_LO(net786));
 sg13g2_tiehi _9943__788 (.L_HI(net788));
 sg13g2_tiehi _9944__789 (.L_HI(net789));
 sg13g2_tiehi \logix.feedback_r[0]$_DFF_P__790  (.L_HI(net790));
 sg13g2_tiehi \logix.feedback_r[1]$_DFF_P__791  (.L_HI(net791));
 sg13g2_tiehi \logix.feedback_r[2]$_DFF_P__792  (.L_HI(net792));
 sg13g2_tiehi \logix.feedback_r[3]$_DFF_P__793  (.L_HI(net793));
 sg13g2_tiehi \logix.feedback_r[4]$_DFF_P__794  (.L_HI(net794));
 sg13g2_tiehi \logix.feedback_r[5]$_DFF_P__795  (.L_HI(net795));
 sg13g2_tiehi \logix.feedback_r[6]$_DFF_P__796  (.L_HI(net796));
 sg13g2_tiehi \logix.feedback_r[7]$_DFF_P__797  (.L_HI(net797));
 sg13g2_tiehi \logix.ram_r[0]$_DFFE_PP__798  (.L_HI(net798));
 sg13g2_tiehi \logix.ram_r[1000]$_DFFE_PP__799  (.L_HI(net799));
 sg13g2_tiehi \logix.ram_r[1001]$_DFFE_PP__800  (.L_HI(net800));
 sg13g2_tiehi \logix.ram_r[1002]$_DFFE_PP__801  (.L_HI(net801));
 sg13g2_tiehi \logix.ram_r[1003]$_DFFE_PP__802  (.L_HI(net802));
 sg13g2_tiehi \logix.ram_r[1004]$_DFFE_PP__803  (.L_HI(net803));
 sg13g2_tiehi \logix.ram_r[1005]$_DFFE_PP__804  (.L_HI(net804));
 sg13g2_tiehi \logix.ram_r[1006]$_DFFE_PP__805  (.L_HI(net805));
 sg13g2_tiehi \logix.ram_r[1007]$_DFFE_PP__806  (.L_HI(net806));
 sg13g2_tiehi \logix.ram_r[1008]$_DFFE_PP__807  (.L_HI(net807));
 sg13g2_tiehi \logix.ram_r[1009]$_DFFE_PP__808  (.L_HI(net808));
 sg13g2_tiehi \logix.ram_r[100]$_DFFE_PP__809  (.L_HI(net809));
 sg13g2_tiehi \logix.ram_r[1010]$_DFFE_PP__810  (.L_HI(net810));
 sg13g2_tiehi \logix.ram_r[1011]$_DFFE_PP__811  (.L_HI(net811));
 sg13g2_tiehi \logix.ram_r[1012]$_DFFE_PP__812  (.L_HI(net812));
 sg13g2_tiehi \logix.ram_r[1013]$_DFFE_PP__813  (.L_HI(net813));
 sg13g2_tiehi \logix.ram_r[1014]$_DFFE_PP__814  (.L_HI(net814));
 sg13g2_tiehi \logix.ram_r[1015]$_DFFE_PP__815  (.L_HI(net815));
 sg13g2_tiehi \logix.ram_r[1016]$_DFFE_PP__816  (.L_HI(net816));
 sg13g2_tiehi \logix.ram_r[1017]$_DFFE_PP__817  (.L_HI(net817));
 sg13g2_tiehi \logix.ram_r[1018]$_DFFE_PP__818  (.L_HI(net818));
 sg13g2_tiehi \logix.ram_r[1019]$_DFFE_PP__819  (.L_HI(net819));
 sg13g2_tiehi \logix.ram_r[101]$_DFFE_PP__820  (.L_HI(net820));
 sg13g2_tiehi \logix.ram_r[1020]$_DFFE_PP__821  (.L_HI(net821));
 sg13g2_tiehi \logix.ram_r[1021]$_DFFE_PP__822  (.L_HI(net822));
 sg13g2_tiehi \logix.ram_r[1022]$_DFFE_PP__823  (.L_HI(net823));
 sg13g2_tiehi \logix.ram_r[1023]$_DFFE_PP__824  (.L_HI(net824));
 sg13g2_tiehi \logix.ram_r[1024]$_DFFE_PP__825  (.L_HI(net825));
 sg13g2_tiehi \logix.ram_r[1025]$_DFFE_PP__826  (.L_HI(net826));
 sg13g2_tiehi \logix.ram_r[1026]$_DFFE_PP__827  (.L_HI(net827));
 sg13g2_tiehi \logix.ram_r[1027]$_DFFE_PP__828  (.L_HI(net828));
 sg13g2_tiehi \logix.ram_r[1028]$_DFFE_PP__829  (.L_HI(net829));
 sg13g2_tiehi \logix.ram_r[1029]$_DFFE_PP__830  (.L_HI(net830));
 sg13g2_tiehi \logix.ram_r[102]$_DFFE_PP__831  (.L_HI(net831));
 sg13g2_tiehi \logix.ram_r[1030]$_DFFE_PP__832  (.L_HI(net832));
 sg13g2_tiehi \logix.ram_r[1031]$_DFFE_PP__833  (.L_HI(net833));
 sg13g2_tiehi \logix.ram_r[1032]$_DFFE_PP__834  (.L_HI(net834));
 sg13g2_tiehi \logix.ram_r[1033]$_DFFE_PP__835  (.L_HI(net835));
 sg13g2_tiehi \logix.ram_r[1034]$_DFFE_PP__836  (.L_HI(net836));
 sg13g2_tiehi \logix.ram_r[1035]$_DFFE_PP__837  (.L_HI(net837));
 sg13g2_tiehi \logix.ram_r[1036]$_DFFE_PP__838  (.L_HI(net838));
 sg13g2_tiehi \logix.ram_r[1037]$_DFFE_PP__839  (.L_HI(net839));
 sg13g2_tiehi \logix.ram_r[1038]$_DFFE_PP__840  (.L_HI(net840));
 sg13g2_tiehi \logix.ram_r[1039]$_DFFE_PP__841  (.L_HI(net841));
 sg13g2_tiehi \logix.ram_r[103]$_DFFE_PP__842  (.L_HI(net842));
 sg13g2_tiehi \logix.ram_r[1040]$_DFFE_PP__843  (.L_HI(net843));
 sg13g2_tiehi \logix.ram_r[1041]$_DFFE_PP__844  (.L_HI(net844));
 sg13g2_tiehi \logix.ram_r[1042]$_DFFE_PP__845  (.L_HI(net845));
 sg13g2_tiehi \logix.ram_r[1043]$_DFFE_PP__846  (.L_HI(net846));
 sg13g2_tiehi \logix.ram_r[1044]$_DFFE_PP__847  (.L_HI(net847));
 sg13g2_tiehi \logix.ram_r[1045]$_DFFE_PP__848  (.L_HI(net848));
 sg13g2_tiehi \logix.ram_r[1046]$_DFFE_PP__849  (.L_HI(net849));
 sg13g2_tiehi \logix.ram_r[1047]$_DFFE_PP__850  (.L_HI(net850));
 sg13g2_tiehi \logix.ram_r[1048]$_DFFE_PP__851  (.L_HI(net851));
 sg13g2_tiehi \logix.ram_r[1049]$_DFFE_PP__852  (.L_HI(net852));
 sg13g2_tiehi \logix.ram_r[104]$_DFFE_PP__853  (.L_HI(net853));
 sg13g2_tiehi \logix.ram_r[1050]$_DFFE_PP__854  (.L_HI(net854));
 sg13g2_tiehi \logix.ram_r[1051]$_DFFE_PP__855  (.L_HI(net855));
 sg13g2_tiehi \logix.ram_r[1052]$_DFFE_PP__856  (.L_HI(net856));
 sg13g2_tiehi \logix.ram_r[1053]$_DFFE_PP__857  (.L_HI(net857));
 sg13g2_tiehi \logix.ram_r[1054]$_DFFE_PP__858  (.L_HI(net858));
 sg13g2_tiehi \logix.ram_r[1055]$_DFFE_PP__859  (.L_HI(net859));
 sg13g2_tiehi \logix.ram_r[1056]$_DFFE_PP__860  (.L_HI(net860));
 sg13g2_tiehi \logix.ram_r[1057]$_DFFE_PP__861  (.L_HI(net861));
 sg13g2_tiehi \logix.ram_r[1058]$_DFFE_PP__862  (.L_HI(net862));
 sg13g2_tiehi \logix.ram_r[1059]$_DFFE_PP__863  (.L_HI(net863));
 sg13g2_tiehi \logix.ram_r[105]$_DFFE_PP__864  (.L_HI(net864));
 sg13g2_tiehi \logix.ram_r[1060]$_DFFE_PP__865  (.L_HI(net865));
 sg13g2_tiehi \logix.ram_r[1061]$_DFFE_PP__866  (.L_HI(net866));
 sg13g2_tiehi \logix.ram_r[1062]$_DFFE_PP__867  (.L_HI(net867));
 sg13g2_tiehi \logix.ram_r[1063]$_DFFE_PP__868  (.L_HI(net868));
 sg13g2_tiehi \logix.ram_r[1064]$_DFFE_PP__869  (.L_HI(net869));
 sg13g2_tiehi \logix.ram_r[1065]$_DFFE_PP__870  (.L_HI(net870));
 sg13g2_tiehi \logix.ram_r[1066]$_DFFE_PP__871  (.L_HI(net871));
 sg13g2_tiehi \logix.ram_r[1067]$_DFFE_PP__872  (.L_HI(net872));
 sg13g2_tiehi \logix.ram_r[1068]$_DFFE_PP__873  (.L_HI(net873));
 sg13g2_tiehi \logix.ram_r[1069]$_DFFE_PP__874  (.L_HI(net874));
 sg13g2_tiehi \logix.ram_r[106]$_DFFE_PP__875  (.L_HI(net875));
 sg13g2_tiehi \logix.ram_r[1070]$_DFFE_PP__876  (.L_HI(net876));
 sg13g2_tiehi \logix.ram_r[1071]$_DFFE_PP__877  (.L_HI(net877));
 sg13g2_tiehi \logix.ram_r[1072]$_DFFE_PP__878  (.L_HI(net878));
 sg13g2_tiehi \logix.ram_r[1073]$_DFFE_PP__879  (.L_HI(net879));
 sg13g2_tiehi \logix.ram_r[1074]$_DFFE_PP__880  (.L_HI(net880));
 sg13g2_tiehi \logix.ram_r[1075]$_DFFE_PP__881  (.L_HI(net881));
 sg13g2_tiehi \logix.ram_r[1076]$_DFFE_PP__882  (.L_HI(net882));
 sg13g2_tiehi \logix.ram_r[1077]$_DFFE_PP__883  (.L_HI(net883));
 sg13g2_tiehi \logix.ram_r[1078]$_DFFE_PP__884  (.L_HI(net884));
 sg13g2_tiehi \logix.ram_r[1079]$_DFFE_PP__885  (.L_HI(net885));
 sg13g2_tiehi \logix.ram_r[107]$_DFFE_PP__886  (.L_HI(net886));
 sg13g2_tiehi \logix.ram_r[1080]$_DFFE_PP__887  (.L_HI(net887));
 sg13g2_tiehi \logix.ram_r[1081]$_DFFE_PP__888  (.L_HI(net888));
 sg13g2_tiehi \logix.ram_r[1082]$_DFFE_PP__889  (.L_HI(net889));
 sg13g2_tiehi \logix.ram_r[1083]$_DFFE_PP__890  (.L_HI(net890));
 sg13g2_tiehi \logix.ram_r[1084]$_DFFE_PP__891  (.L_HI(net891));
 sg13g2_tiehi \logix.ram_r[1085]$_DFFE_PP__892  (.L_HI(net892));
 sg13g2_tiehi \logix.ram_r[1086]$_DFFE_PP__893  (.L_HI(net893));
 sg13g2_tiehi \logix.ram_r[1087]$_DFFE_PP__894  (.L_HI(net894));
 sg13g2_tiehi \logix.ram_r[1088]$_DFFE_PP__895  (.L_HI(net895));
 sg13g2_tiehi \logix.ram_r[1089]$_DFFE_PP__896  (.L_HI(net896));
 sg13g2_tiehi \logix.ram_r[108]$_DFFE_PP__897  (.L_HI(net897));
 sg13g2_tiehi \logix.ram_r[1090]$_DFFE_PP__898  (.L_HI(net898));
 sg13g2_tiehi \logix.ram_r[1091]$_DFFE_PP__899  (.L_HI(net899));
 sg13g2_tiehi \logix.ram_r[1092]$_DFFE_PP__900  (.L_HI(net900));
 sg13g2_tiehi \logix.ram_r[1093]$_DFFE_PP__901  (.L_HI(net901));
 sg13g2_tiehi \logix.ram_r[1094]$_DFFE_PP__902  (.L_HI(net902));
 sg13g2_tiehi \logix.ram_r[1095]$_DFFE_PP__903  (.L_HI(net903));
 sg13g2_tiehi \logix.ram_r[1096]$_DFFE_PP__904  (.L_HI(net904));
 sg13g2_tiehi \logix.ram_r[1097]$_DFFE_PP__905  (.L_HI(net905));
 sg13g2_tiehi \logix.ram_r[1098]$_DFFE_PP__906  (.L_HI(net906));
 sg13g2_tiehi \logix.ram_r[1099]$_DFFE_PP__907  (.L_HI(net907));
 sg13g2_tiehi \logix.ram_r[109]$_DFFE_PP__908  (.L_HI(net908));
 sg13g2_tiehi \logix.ram_r[10]$_DFFE_PP__909  (.L_HI(net909));
 sg13g2_tiehi \logix.ram_r[1100]$_DFFE_PP__910  (.L_HI(net910));
 sg13g2_tiehi \logix.ram_r[1101]$_DFFE_PP__911  (.L_HI(net911));
 sg13g2_tiehi \logix.ram_r[1102]$_DFFE_PP__912  (.L_HI(net912));
 sg13g2_tiehi \logix.ram_r[1103]$_DFFE_PP__913  (.L_HI(net913));
 sg13g2_tiehi \logix.ram_r[1104]$_DFFE_PP__914  (.L_HI(net914));
 sg13g2_tiehi \logix.ram_r[1105]$_DFFE_PP__915  (.L_HI(net915));
 sg13g2_tiehi \logix.ram_r[1106]$_DFFE_PP__916  (.L_HI(net916));
 sg13g2_tiehi \logix.ram_r[1107]$_DFFE_PP__917  (.L_HI(net917));
 sg13g2_tiehi \logix.ram_r[1108]$_DFFE_PP__918  (.L_HI(net918));
 sg13g2_tiehi \logix.ram_r[1109]$_DFFE_PP__919  (.L_HI(net919));
 sg13g2_tiehi \logix.ram_r[110]$_DFFE_PP__920  (.L_HI(net920));
 sg13g2_tiehi \logix.ram_r[1110]$_DFFE_PP__921  (.L_HI(net921));
 sg13g2_tiehi \logix.ram_r[1111]$_DFFE_PP__922  (.L_HI(net922));
 sg13g2_tiehi \logix.ram_r[1112]$_DFFE_PP__923  (.L_HI(net923));
 sg13g2_tiehi \logix.ram_r[1113]$_DFFE_PP__924  (.L_HI(net924));
 sg13g2_tiehi \logix.ram_r[1114]$_DFFE_PP__925  (.L_HI(net925));
 sg13g2_tiehi \logix.ram_r[1115]$_DFFE_PP__926  (.L_HI(net926));
 sg13g2_tiehi \logix.ram_r[1116]$_DFFE_PP__927  (.L_HI(net927));
 sg13g2_tiehi \logix.ram_r[1117]$_DFFE_PP__928  (.L_HI(net928));
 sg13g2_tiehi \logix.ram_r[1118]$_DFFE_PP__929  (.L_HI(net929));
 sg13g2_tiehi \logix.ram_r[1119]$_DFFE_PP__930  (.L_HI(net930));
 sg13g2_tiehi \logix.ram_r[111]$_DFFE_PP__931  (.L_HI(net931));
 sg13g2_tiehi \logix.ram_r[1120]$_DFFE_PP__932  (.L_HI(net932));
 sg13g2_tiehi \logix.ram_r[1121]$_DFFE_PP__933  (.L_HI(net933));
 sg13g2_tiehi \logix.ram_r[1122]$_DFFE_PP__934  (.L_HI(net934));
 sg13g2_tiehi \logix.ram_r[1123]$_DFFE_PP__935  (.L_HI(net935));
 sg13g2_tiehi \logix.ram_r[1124]$_DFFE_PP__936  (.L_HI(net936));
 sg13g2_tiehi \logix.ram_r[1125]$_DFFE_PP__937  (.L_HI(net937));
 sg13g2_tiehi \logix.ram_r[1126]$_DFFE_PP__938  (.L_HI(net938));
 sg13g2_tiehi \logix.ram_r[1127]$_DFFE_PP__939  (.L_HI(net939));
 sg13g2_tiehi \logix.ram_r[1128]$_DFFE_PP__940  (.L_HI(net940));
 sg13g2_tiehi \logix.ram_r[1129]$_DFFE_PP__941  (.L_HI(net941));
 sg13g2_tiehi \logix.ram_r[112]$_DFFE_PP__942  (.L_HI(net942));
 sg13g2_tiehi \logix.ram_r[1130]$_DFFE_PP__943  (.L_HI(net943));
 sg13g2_tiehi \logix.ram_r[1131]$_DFFE_PP__944  (.L_HI(net944));
 sg13g2_tiehi \logix.ram_r[1132]$_DFFE_PP__945  (.L_HI(net945));
 sg13g2_tiehi \logix.ram_r[1133]$_DFFE_PP__946  (.L_HI(net946));
 sg13g2_tiehi \logix.ram_r[1134]$_DFFE_PP__947  (.L_HI(net947));
 sg13g2_tiehi \logix.ram_r[1135]$_DFFE_PP__948  (.L_HI(net948));
 sg13g2_tiehi \logix.ram_r[1136]$_DFFE_PP__949  (.L_HI(net949));
 sg13g2_tiehi \logix.ram_r[1137]$_DFFE_PP__950  (.L_HI(net950));
 sg13g2_tiehi \logix.ram_r[1138]$_DFFE_PP__951  (.L_HI(net951));
 sg13g2_tiehi \logix.ram_r[1139]$_DFFE_PP__952  (.L_HI(net952));
 sg13g2_tiehi \logix.ram_r[113]$_DFFE_PP__953  (.L_HI(net953));
 sg13g2_tiehi \logix.ram_r[1140]$_DFFE_PP__954  (.L_HI(net954));
 sg13g2_tiehi \logix.ram_r[1141]$_DFFE_PP__955  (.L_HI(net955));
 sg13g2_tiehi \logix.ram_r[1142]$_DFFE_PP__956  (.L_HI(net956));
 sg13g2_tiehi \logix.ram_r[1143]$_DFFE_PP__957  (.L_HI(net957));
 sg13g2_tiehi \logix.ram_r[1144]$_DFFE_PP__958  (.L_HI(net958));
 sg13g2_tiehi \logix.ram_r[1145]$_DFFE_PP__959  (.L_HI(net959));
 sg13g2_tiehi \logix.ram_r[1146]$_DFFE_PP__960  (.L_HI(net960));
 sg13g2_tiehi \logix.ram_r[1147]$_DFFE_PP__961  (.L_HI(net961));
 sg13g2_tiehi \logix.ram_r[1148]$_DFFE_PP__962  (.L_HI(net962));
 sg13g2_tiehi \logix.ram_r[1149]$_DFFE_PP__963  (.L_HI(net963));
 sg13g2_tiehi \logix.ram_r[114]$_DFFE_PP__964  (.L_HI(net964));
 sg13g2_tiehi \logix.ram_r[1150]$_DFFE_PP__965  (.L_HI(net965));
 sg13g2_tiehi \logix.ram_r[1151]$_DFFE_PP__966  (.L_HI(net966));
 sg13g2_tiehi \logix.ram_r[1152]$_DFFE_PP__967  (.L_HI(net967));
 sg13g2_tiehi \logix.ram_r[1153]$_DFFE_PP__968  (.L_HI(net968));
 sg13g2_tiehi \logix.ram_r[1154]$_DFFE_PP__969  (.L_HI(net969));
 sg13g2_tiehi \logix.ram_r[1155]$_DFFE_PP__970  (.L_HI(net970));
 sg13g2_tiehi \logix.ram_r[1156]$_DFFE_PP__971  (.L_HI(net971));
 sg13g2_tiehi \logix.ram_r[1157]$_DFFE_PP__972  (.L_HI(net972));
 sg13g2_tiehi \logix.ram_r[1158]$_DFFE_PP__973  (.L_HI(net973));
 sg13g2_tiehi \logix.ram_r[1159]$_DFFE_PP__974  (.L_HI(net974));
 sg13g2_tiehi \logix.ram_r[115]$_DFFE_PP__975  (.L_HI(net975));
 sg13g2_tiehi \logix.ram_r[1160]$_DFFE_PP__976  (.L_HI(net976));
 sg13g2_tiehi \logix.ram_r[1161]$_DFFE_PP__977  (.L_HI(net977));
 sg13g2_tiehi \logix.ram_r[1162]$_DFFE_PP__978  (.L_HI(net978));
 sg13g2_tiehi \logix.ram_r[1163]$_DFFE_PP__979  (.L_HI(net979));
 sg13g2_tiehi \logix.ram_r[1164]$_DFFE_PP__980  (.L_HI(net980));
 sg13g2_tiehi \logix.ram_r[1165]$_DFFE_PP__981  (.L_HI(net981));
 sg13g2_tiehi \logix.ram_r[1166]$_DFFE_PP__982  (.L_HI(net982));
 sg13g2_tiehi \logix.ram_r[1167]$_DFFE_PP__983  (.L_HI(net983));
 sg13g2_tiehi \logix.ram_r[1168]$_DFFE_PP__984  (.L_HI(net984));
 sg13g2_tiehi \logix.ram_r[1169]$_DFFE_PP__985  (.L_HI(net985));
 sg13g2_tiehi \logix.ram_r[116]$_DFFE_PP__986  (.L_HI(net986));
 sg13g2_tiehi \logix.ram_r[1170]$_DFFE_PP__987  (.L_HI(net987));
 sg13g2_tiehi \logix.ram_r[1171]$_DFFE_PP__988  (.L_HI(net988));
 sg13g2_tiehi \logix.ram_r[1172]$_DFFE_PP__989  (.L_HI(net989));
 sg13g2_tiehi \logix.ram_r[1173]$_DFFE_PP__990  (.L_HI(net990));
 sg13g2_tiehi \logix.ram_r[1174]$_DFFE_PP__991  (.L_HI(net991));
 sg13g2_tiehi \logix.ram_r[1175]$_DFFE_PP__992  (.L_HI(net992));
 sg13g2_tiehi \logix.ram_r[1176]$_DFFE_PP__993  (.L_HI(net993));
 sg13g2_tiehi \logix.ram_r[1177]$_DFFE_PP__994  (.L_HI(net994));
 sg13g2_tiehi \logix.ram_r[1178]$_DFFE_PP__995  (.L_HI(net995));
 sg13g2_tiehi \logix.ram_r[1179]$_DFFE_PP__996  (.L_HI(net996));
 sg13g2_tiehi \logix.ram_r[117]$_DFFE_PP__997  (.L_HI(net997));
 sg13g2_tiehi \logix.ram_r[1180]$_DFFE_PP__998  (.L_HI(net998));
 sg13g2_tiehi \logix.ram_r[1181]$_DFFE_PP__999  (.L_HI(net999));
 sg13g2_tiehi \logix.ram_r[1182]$_DFFE_PP__1000  (.L_HI(net1000));
 sg13g2_tiehi \logix.ram_r[1183]$_DFFE_PP__1001  (.L_HI(net1001));
 sg13g2_tiehi \logix.ram_r[1184]$_DFFE_PP__1002  (.L_HI(net1002));
 sg13g2_tiehi \logix.ram_r[1185]$_DFFE_PP__1003  (.L_HI(net1003));
 sg13g2_tiehi \logix.ram_r[1186]$_DFFE_PP__1004  (.L_HI(net1004));
 sg13g2_tiehi \logix.ram_r[1187]$_DFFE_PP__1005  (.L_HI(net1005));
 sg13g2_tiehi \logix.ram_r[1188]$_DFFE_PP__1006  (.L_HI(net1006));
 sg13g2_tiehi \logix.ram_r[1189]$_DFFE_PP__1007  (.L_HI(net1007));
 sg13g2_tiehi \logix.ram_r[118]$_DFFE_PP__1008  (.L_HI(net1008));
 sg13g2_tiehi \logix.ram_r[1190]$_DFFE_PP__1009  (.L_HI(net1009));
 sg13g2_tiehi \logix.ram_r[1191]$_DFFE_PP__1010  (.L_HI(net1010));
 sg13g2_tiehi \logix.ram_r[1192]$_DFFE_PP__1011  (.L_HI(net1011));
 sg13g2_tiehi \logix.ram_r[1193]$_DFFE_PP__1012  (.L_HI(net1012));
 sg13g2_tiehi \logix.ram_r[1194]$_DFFE_PP__1013  (.L_HI(net1013));
 sg13g2_tiehi \logix.ram_r[1195]$_DFFE_PP__1014  (.L_HI(net1014));
 sg13g2_tiehi \logix.ram_r[1196]$_DFFE_PP__1015  (.L_HI(net1015));
 sg13g2_tiehi \logix.ram_r[1197]$_DFFE_PP__1016  (.L_HI(net1016));
 sg13g2_tiehi \logix.ram_r[1198]$_DFFE_PP__1017  (.L_HI(net1017));
 sg13g2_tiehi \logix.ram_r[1199]$_DFFE_PP__1018  (.L_HI(net1018));
 sg13g2_tiehi \logix.ram_r[119]$_DFFE_PP__1019  (.L_HI(net1019));
 sg13g2_tiehi \logix.ram_r[11]$_DFFE_PP__1020  (.L_HI(net1020));
 sg13g2_tiehi \logix.ram_r[1200]$_DFFE_PP__1021  (.L_HI(net1021));
 sg13g2_tiehi \logix.ram_r[1201]$_DFFE_PP__1022  (.L_HI(net1022));
 sg13g2_tiehi \logix.ram_r[1202]$_DFFE_PP__1023  (.L_HI(net1023));
 sg13g2_tiehi \logix.ram_r[1203]$_DFFE_PP__1024  (.L_HI(net1024));
 sg13g2_tiehi \logix.ram_r[1204]$_DFFE_PP__1025  (.L_HI(net1025));
 sg13g2_tiehi \logix.ram_r[1205]$_DFFE_PP__1026  (.L_HI(net1026));
 sg13g2_tiehi \logix.ram_r[1206]$_DFFE_PP__1027  (.L_HI(net1027));
 sg13g2_tiehi \logix.ram_r[1207]$_DFFE_PP__1028  (.L_HI(net1028));
 sg13g2_tiehi \logix.ram_r[1208]$_DFFE_PP__1029  (.L_HI(net1029));
 sg13g2_tiehi \logix.ram_r[1209]$_DFFE_PP__1030  (.L_HI(net1030));
 sg13g2_tiehi \logix.ram_r[120]$_DFFE_PP__1031  (.L_HI(net1031));
 sg13g2_tiehi \logix.ram_r[1210]$_DFFE_PP__1032  (.L_HI(net1032));
 sg13g2_tiehi \logix.ram_r[1211]$_DFFE_PP__1033  (.L_HI(net1033));
 sg13g2_tiehi \logix.ram_r[1212]$_DFFE_PP__1034  (.L_HI(net1034));
 sg13g2_tiehi \logix.ram_r[1213]$_DFFE_PP__1035  (.L_HI(net1035));
 sg13g2_tiehi \logix.ram_r[1214]$_DFFE_PP__1036  (.L_HI(net1036));
 sg13g2_tiehi \logix.ram_r[1215]$_DFFE_PP__1037  (.L_HI(net1037));
 sg13g2_tiehi \logix.ram_r[1216]$_DFFE_PP__1038  (.L_HI(net1038));
 sg13g2_tiehi \logix.ram_r[1217]$_DFFE_PP__1039  (.L_HI(net1039));
 sg13g2_tiehi \logix.ram_r[1218]$_DFFE_PP__1040  (.L_HI(net1040));
 sg13g2_tiehi \logix.ram_r[1219]$_DFFE_PP__1041  (.L_HI(net1041));
 sg13g2_tiehi \logix.ram_r[121]$_DFFE_PP__1042  (.L_HI(net1042));
 sg13g2_tiehi \logix.ram_r[1220]$_DFFE_PP__1043  (.L_HI(net1043));
 sg13g2_tiehi \logix.ram_r[1221]$_DFFE_PP__1044  (.L_HI(net1044));
 sg13g2_tiehi \logix.ram_r[1222]$_DFFE_PP__1045  (.L_HI(net1045));
 sg13g2_tiehi \logix.ram_r[1223]$_DFFE_PP__1046  (.L_HI(net1046));
 sg13g2_tiehi \logix.ram_r[1224]$_DFFE_PP__1047  (.L_HI(net1047));
 sg13g2_tiehi \logix.ram_r[1225]$_DFFE_PP__1048  (.L_HI(net1048));
 sg13g2_tiehi \logix.ram_r[1226]$_DFFE_PP__1049  (.L_HI(net1049));
 sg13g2_tiehi \logix.ram_r[1227]$_DFFE_PP__1050  (.L_HI(net1050));
 sg13g2_tiehi \logix.ram_r[1228]$_DFFE_PP__1051  (.L_HI(net1051));
 sg13g2_tiehi \logix.ram_r[1229]$_DFFE_PP__1052  (.L_HI(net1052));
 sg13g2_tiehi \logix.ram_r[122]$_DFFE_PP__1053  (.L_HI(net1053));
 sg13g2_tiehi \logix.ram_r[1230]$_DFFE_PP__1054  (.L_HI(net1054));
 sg13g2_tiehi \logix.ram_r[1231]$_DFFE_PP__1055  (.L_HI(net1055));
 sg13g2_tiehi \logix.ram_r[1232]$_DFFE_PP__1056  (.L_HI(net1056));
 sg13g2_tiehi \logix.ram_r[1233]$_DFFE_PP__1057  (.L_HI(net1057));
 sg13g2_tiehi \logix.ram_r[1234]$_DFFE_PP__1058  (.L_HI(net1058));
 sg13g2_tiehi \logix.ram_r[1235]$_DFFE_PP__1059  (.L_HI(net1059));
 sg13g2_tiehi \logix.ram_r[1236]$_DFFE_PP__1060  (.L_HI(net1060));
 sg13g2_tiehi \logix.ram_r[1237]$_DFFE_PP__1061  (.L_HI(net1061));
 sg13g2_tiehi \logix.ram_r[1238]$_DFFE_PP__1062  (.L_HI(net1062));
 sg13g2_tiehi \logix.ram_r[1239]$_DFFE_PP__1063  (.L_HI(net1063));
 sg13g2_tiehi \logix.ram_r[123]$_DFFE_PP__1064  (.L_HI(net1064));
 sg13g2_tiehi \logix.ram_r[1240]$_DFFE_PP__1065  (.L_HI(net1065));
 sg13g2_tiehi \logix.ram_r[1241]$_DFFE_PP__1066  (.L_HI(net1066));
 sg13g2_tiehi \logix.ram_r[1242]$_DFFE_PP__1067  (.L_HI(net1067));
 sg13g2_tiehi \logix.ram_r[1243]$_DFFE_PP__1068  (.L_HI(net1068));
 sg13g2_tiehi \logix.ram_r[1244]$_DFFE_PP__1069  (.L_HI(net1069));
 sg13g2_tiehi \logix.ram_r[1245]$_DFFE_PP__1070  (.L_HI(net1070));
 sg13g2_tiehi \logix.ram_r[1246]$_DFFE_PP__1071  (.L_HI(net1071));
 sg13g2_tiehi \logix.ram_r[1247]$_DFFE_PP__1072  (.L_HI(net1072));
 sg13g2_tiehi \logix.ram_r[1248]$_DFFE_PP__1073  (.L_HI(net1073));
 sg13g2_tiehi \logix.ram_r[1249]$_DFFE_PP__1074  (.L_HI(net1074));
 sg13g2_tiehi \logix.ram_r[124]$_DFFE_PP__1075  (.L_HI(net1075));
 sg13g2_tiehi \logix.ram_r[1250]$_DFFE_PP__1076  (.L_HI(net1076));
 sg13g2_tiehi \logix.ram_r[1251]$_DFFE_PP__1077  (.L_HI(net1077));
 sg13g2_tiehi \logix.ram_r[1252]$_DFFE_PP__1078  (.L_HI(net1078));
 sg13g2_tiehi \logix.ram_r[1253]$_DFFE_PP__1079  (.L_HI(net1079));
 sg13g2_tiehi \logix.ram_r[1254]$_DFFE_PP__1080  (.L_HI(net1080));
 sg13g2_tiehi \logix.ram_r[1255]$_DFFE_PP__1081  (.L_HI(net1081));
 sg13g2_tiehi \logix.ram_r[1256]$_DFFE_PP__1082  (.L_HI(net1082));
 sg13g2_tiehi \logix.ram_r[1257]$_DFFE_PP__1083  (.L_HI(net1083));
 sg13g2_tiehi \logix.ram_r[1258]$_DFFE_PP__1084  (.L_HI(net1084));
 sg13g2_tiehi \logix.ram_r[1259]$_DFFE_PP__1085  (.L_HI(net1085));
 sg13g2_tiehi \logix.ram_r[125]$_DFFE_PP__1086  (.L_HI(net1086));
 sg13g2_tiehi \logix.ram_r[1260]$_DFFE_PP__1087  (.L_HI(net1087));
 sg13g2_tiehi \logix.ram_r[1261]$_DFFE_PP__1088  (.L_HI(net1088));
 sg13g2_tiehi \logix.ram_r[1262]$_DFFE_PP__1089  (.L_HI(net1089));
 sg13g2_tiehi \logix.ram_r[1263]$_DFFE_PP__1090  (.L_HI(net1090));
 sg13g2_tiehi \logix.ram_r[1264]$_DFFE_PP__1091  (.L_HI(net1091));
 sg13g2_tiehi \logix.ram_r[1265]$_DFFE_PP__1092  (.L_HI(net1092));
 sg13g2_tiehi \logix.ram_r[1266]$_DFFE_PP__1093  (.L_HI(net1093));
 sg13g2_tiehi \logix.ram_r[1267]$_DFFE_PP__1094  (.L_HI(net1094));
 sg13g2_tiehi \logix.ram_r[1268]$_DFFE_PP__1095  (.L_HI(net1095));
 sg13g2_tiehi \logix.ram_r[1269]$_DFFE_PP__1096  (.L_HI(net1096));
 sg13g2_tiehi \logix.ram_r[126]$_DFFE_PP__1097  (.L_HI(net1097));
 sg13g2_tiehi \logix.ram_r[1270]$_DFFE_PP__1098  (.L_HI(net1098));
 sg13g2_tiehi \logix.ram_r[1271]$_DFFE_PP__1099  (.L_HI(net1099));
 sg13g2_tiehi \logix.ram_r[1272]$_DFFE_PP__1100  (.L_HI(net1100));
 sg13g2_tiehi \logix.ram_r[1273]$_DFFE_PP__1101  (.L_HI(net1101));
 sg13g2_tiehi \logix.ram_r[1274]$_DFFE_PP__1102  (.L_HI(net1102));
 sg13g2_tiehi \logix.ram_r[1275]$_DFFE_PP__1103  (.L_HI(net1103));
 sg13g2_tiehi \logix.ram_r[1276]$_DFFE_PP__1104  (.L_HI(net1104));
 sg13g2_tiehi \logix.ram_r[1277]$_DFFE_PP__1105  (.L_HI(net1105));
 sg13g2_tiehi \logix.ram_r[1278]$_DFFE_PP__1106  (.L_HI(net1106));
 sg13g2_tiehi \logix.ram_r[1279]$_DFFE_PP__1107  (.L_HI(net1107));
 sg13g2_tiehi \logix.ram_r[127]$_DFFE_PP__1108  (.L_HI(net1108));
 sg13g2_tiehi \logix.ram_r[1280]$_DFFE_PP__1109  (.L_HI(net1109));
 sg13g2_tiehi \logix.ram_r[1281]$_DFFE_PP__1110  (.L_HI(net1110));
 sg13g2_tiehi \logix.ram_r[1282]$_DFFE_PP__1111  (.L_HI(net1111));
 sg13g2_tiehi \logix.ram_r[1283]$_DFFE_PP__1112  (.L_HI(net1112));
 sg13g2_tiehi \logix.ram_r[1284]$_DFFE_PP__1113  (.L_HI(net1113));
 sg13g2_tiehi \logix.ram_r[1285]$_DFFE_PP__1114  (.L_HI(net1114));
 sg13g2_tiehi \logix.ram_r[1286]$_DFFE_PP__1115  (.L_HI(net1115));
 sg13g2_tiehi \logix.ram_r[1287]$_DFFE_PP__1116  (.L_HI(net1116));
 sg13g2_tiehi \logix.ram_r[1288]$_DFFE_PP__1117  (.L_HI(net1117));
 sg13g2_tiehi \logix.ram_r[1289]$_DFFE_PP__1118  (.L_HI(net1118));
 sg13g2_tiehi \logix.ram_r[128]$_DFFE_PP__1119  (.L_HI(net1119));
 sg13g2_tiehi \logix.ram_r[1290]$_DFFE_PP__1120  (.L_HI(net1120));
 sg13g2_tiehi \logix.ram_r[1291]$_DFFE_PP__1121  (.L_HI(net1121));
 sg13g2_tiehi \logix.ram_r[1292]$_DFFE_PP__1122  (.L_HI(net1122));
 sg13g2_tiehi \logix.ram_r[1293]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \logix.ram_r[1294]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \logix.ram_r[1295]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \logix.ram_r[1296]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \logix.ram_r[1297]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \logix.ram_r[1298]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \logix.ram_r[1299]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \logix.ram_r[129]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \logix.ram_r[12]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \logix.ram_r[1300]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \logix.ram_r[1301]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \logix.ram_r[1302]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \logix.ram_r[1303]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \logix.ram_r[1304]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \logix.ram_r[1305]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \logix.ram_r[1306]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \logix.ram_r[1307]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \logix.ram_r[1308]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \logix.ram_r[1309]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \logix.ram_r[130]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \logix.ram_r[1310]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \logix.ram_r[1311]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \logix.ram_r[1312]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \logix.ram_r[1313]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \logix.ram_r[1314]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \logix.ram_r[1315]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \logix.ram_r[1316]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \logix.ram_r[1317]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \logix.ram_r[1318]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \logix.ram_r[1319]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \logix.ram_r[131]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \logix.ram_r[1320]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \logix.ram_r[1321]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \logix.ram_r[1322]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \logix.ram_r[1323]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \logix.ram_r[1324]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \logix.ram_r[1325]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \logix.ram_r[1326]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \logix.ram_r[1327]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \logix.ram_r[1328]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \logix.ram_r[1329]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \logix.ram_r[132]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \logix.ram_r[1330]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \logix.ram_r[1331]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \logix.ram_r[1332]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \logix.ram_r[1333]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \logix.ram_r[1334]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \logix.ram_r[1335]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \logix.ram_r[1336]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \logix.ram_r[1337]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \logix.ram_r[1338]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \logix.ram_r[1339]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \logix.ram_r[133]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \logix.ram_r[1340]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \logix.ram_r[1341]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \logix.ram_r[1342]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \logix.ram_r[1343]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \logix.ram_r[1344]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \logix.ram_r[1345]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \logix.ram_r[1346]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \logix.ram_r[1347]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \logix.ram_r[1348]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \logix.ram_r[1349]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \logix.ram_r[134]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \logix.ram_r[1350]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \logix.ram_r[1351]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \logix.ram_r[1352]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \logix.ram_r[1353]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \logix.ram_r[1354]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \logix.ram_r[1355]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \logix.ram_r[1356]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \logix.ram_r[1357]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \logix.ram_r[1358]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \logix.ram_r[1359]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \logix.ram_r[135]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \logix.ram_r[1360]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \logix.ram_r[1361]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \logix.ram_r[1362]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \logix.ram_r[1363]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \logix.ram_r[1364]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \logix.ram_r[1365]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \logix.ram_r[1366]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \logix.ram_r[1367]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \logix.ram_r[1368]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \logix.ram_r[1369]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \logix.ram_r[136]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \logix.ram_r[1370]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \logix.ram_r[1371]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \logix.ram_r[1372]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \logix.ram_r[1373]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \logix.ram_r[1374]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \logix.ram_r[1375]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \logix.ram_r[1376]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \logix.ram_r[1377]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \logix.ram_r[1378]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \logix.ram_r[1379]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \logix.ram_r[137]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \logix.ram_r[1380]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \logix.ram_r[1381]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \logix.ram_r[1382]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \logix.ram_r[1383]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \logix.ram_r[1384]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \logix.ram_r[1385]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \logix.ram_r[1386]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \logix.ram_r[1387]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \logix.ram_r[1388]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \logix.ram_r[1389]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \logix.ram_r[138]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \logix.ram_r[1390]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \logix.ram_r[1391]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \logix.ram_r[1392]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \logix.ram_r[1393]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \logix.ram_r[1394]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \logix.ram_r[1395]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \logix.ram_r[1396]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \logix.ram_r[1397]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \logix.ram_r[1398]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \logix.ram_r[1399]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \logix.ram_r[139]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \logix.ram_r[13]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \logix.ram_r[1400]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \logix.ram_r[1401]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \logix.ram_r[1402]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \logix.ram_r[1403]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \logix.ram_r[1404]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \logix.ram_r[1405]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \logix.ram_r[1406]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \logix.ram_r[1407]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \logix.ram_r[1408]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \logix.ram_r[1409]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \logix.ram_r[140]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \logix.ram_r[1410]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \logix.ram_r[1411]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \logix.ram_r[1412]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \logix.ram_r[1413]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \logix.ram_r[1414]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \logix.ram_r[1415]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \logix.ram_r[1416]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \logix.ram_r[1417]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \logix.ram_r[1418]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \logix.ram_r[1419]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \logix.ram_r[141]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \logix.ram_r[1420]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \logix.ram_r[1421]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \logix.ram_r[1422]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \logix.ram_r[1423]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \logix.ram_r[1424]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \logix.ram_r[1425]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \logix.ram_r[1426]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \logix.ram_r[1427]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \logix.ram_r[1428]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \logix.ram_r[1429]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \logix.ram_r[142]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \logix.ram_r[1430]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \logix.ram_r[1431]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \logix.ram_r[1432]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \logix.ram_r[1433]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \logix.ram_r[1434]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \logix.ram_r[1435]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \logix.ram_r[1436]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \logix.ram_r[1437]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \logix.ram_r[1438]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \logix.ram_r[1439]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \logix.ram_r[143]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \logix.ram_r[1440]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \logix.ram_r[1441]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \logix.ram_r[1442]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \logix.ram_r[1443]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \logix.ram_r[1444]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \logix.ram_r[1445]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \logix.ram_r[1446]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \logix.ram_r[1447]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \logix.ram_r[1448]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \logix.ram_r[1449]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \logix.ram_r[144]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \logix.ram_r[1450]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \logix.ram_r[1451]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \logix.ram_r[1452]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \logix.ram_r[1453]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \logix.ram_r[1454]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \logix.ram_r[1455]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \logix.ram_r[1456]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \logix.ram_r[1457]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \logix.ram_r[1458]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \logix.ram_r[1459]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \logix.ram_r[145]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \logix.ram_r[1460]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \logix.ram_r[1461]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \logix.ram_r[1462]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \logix.ram_r[1463]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \logix.ram_r[1464]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \logix.ram_r[1465]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \logix.ram_r[1466]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \logix.ram_r[1467]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \logix.ram_r[1468]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \logix.ram_r[1469]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \logix.ram_r[146]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \logix.ram_r[1470]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \logix.ram_r[1471]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \logix.ram_r[1472]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \logix.ram_r[1473]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \logix.ram_r[1474]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \logix.ram_r[1475]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \logix.ram_r[1476]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \logix.ram_r[1477]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \logix.ram_r[1478]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \logix.ram_r[1479]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \logix.ram_r[147]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \logix.ram_r[1480]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \logix.ram_r[1481]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \logix.ram_r[1482]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \logix.ram_r[1483]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \logix.ram_r[1484]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \logix.ram_r[1485]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \logix.ram_r[1486]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \logix.ram_r[1487]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \logix.ram_r[1488]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \logix.ram_r[1489]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \logix.ram_r[148]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \logix.ram_r[1490]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \logix.ram_r[1491]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \logix.ram_r[1492]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \logix.ram_r[1493]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \logix.ram_r[1494]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \logix.ram_r[1495]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \logix.ram_r[1496]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \logix.ram_r[1497]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \logix.ram_r[1498]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \logix.ram_r[1499]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \logix.ram_r[149]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \logix.ram_r[14]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \logix.ram_r[1500]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \logix.ram_r[1501]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \logix.ram_r[1502]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \logix.ram_r[1503]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \logix.ram_r[1504]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \logix.ram_r[1505]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \logix.ram_r[1506]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \logix.ram_r[1507]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \logix.ram_r[1508]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \logix.ram_r[1509]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \logix.ram_r[150]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \logix.ram_r[1510]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \logix.ram_r[1511]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \logix.ram_r[1512]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \logix.ram_r[1513]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \logix.ram_r[1514]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \logix.ram_r[1515]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \logix.ram_r[1516]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \logix.ram_r[1517]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \logix.ram_r[1518]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \logix.ram_r[1519]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \logix.ram_r[151]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \logix.ram_r[1520]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \logix.ram_r[1521]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \logix.ram_r[1522]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \logix.ram_r[1523]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \logix.ram_r[1524]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \logix.ram_r[1525]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \logix.ram_r[1526]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \logix.ram_r[1527]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \logix.ram_r[1528]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \logix.ram_r[1529]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \logix.ram_r[152]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \logix.ram_r[1530]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \logix.ram_r[1531]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \logix.ram_r[1532]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \logix.ram_r[1533]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \logix.ram_r[1534]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \logix.ram_r[1535]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \logix.ram_r[1536]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \logix.ram_r[1537]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \logix.ram_r[1538]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \logix.ram_r[1539]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \logix.ram_r[153]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \logix.ram_r[1540]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \logix.ram_r[1541]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \logix.ram_r[1542]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \logix.ram_r[1543]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \logix.ram_r[1544]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \logix.ram_r[1545]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \logix.ram_r[1546]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \logix.ram_r[1547]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \logix.ram_r[1548]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \logix.ram_r[1549]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \logix.ram_r[154]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \logix.ram_r[1550]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \logix.ram_r[1551]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \logix.ram_r[1552]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \logix.ram_r[1553]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \logix.ram_r[1554]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \logix.ram_r[1555]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \logix.ram_r[1556]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \logix.ram_r[1557]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \logix.ram_r[1558]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \logix.ram_r[1559]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \logix.ram_r[155]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \logix.ram_r[1560]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \logix.ram_r[1561]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \logix.ram_r[1562]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \logix.ram_r[1563]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \logix.ram_r[1564]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \logix.ram_r[1565]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \logix.ram_r[1566]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \logix.ram_r[1567]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \logix.ram_r[1568]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \logix.ram_r[1569]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \logix.ram_r[156]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \logix.ram_r[1570]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \logix.ram_r[1571]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \logix.ram_r[1572]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \logix.ram_r[1573]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \logix.ram_r[1574]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \logix.ram_r[1575]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \logix.ram_r[1576]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \logix.ram_r[1577]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \logix.ram_r[1578]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \logix.ram_r[1579]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \logix.ram_r[157]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \logix.ram_r[1580]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \logix.ram_r[1581]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \logix.ram_r[1582]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \logix.ram_r[1583]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \logix.ram_r[1584]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \logix.ram_r[1585]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \logix.ram_r[1586]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \logix.ram_r[1587]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \logix.ram_r[1588]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \logix.ram_r[1589]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \logix.ram_r[158]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \logix.ram_r[1590]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \logix.ram_r[1591]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \logix.ram_r[1592]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \logix.ram_r[1593]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \logix.ram_r[1594]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \logix.ram_r[1595]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \logix.ram_r[1596]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \logix.ram_r[1597]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \logix.ram_r[1598]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \logix.ram_r[1599]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \logix.ram_r[159]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \logix.ram_r[15]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \logix.ram_r[1600]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \logix.ram_r[1601]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \logix.ram_r[1602]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \logix.ram_r[1603]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \logix.ram_r[1604]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \logix.ram_r[1605]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \logix.ram_r[1606]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \logix.ram_r[1607]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \logix.ram_r[1608]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \logix.ram_r[1609]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \logix.ram_r[160]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \logix.ram_r[1610]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \logix.ram_r[1611]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \logix.ram_r[1612]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \logix.ram_r[1613]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \logix.ram_r[1614]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \logix.ram_r[1615]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \logix.ram_r[1616]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \logix.ram_r[1617]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \logix.ram_r[1618]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \logix.ram_r[1619]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \logix.ram_r[161]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \logix.ram_r[1620]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \logix.ram_r[1621]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \logix.ram_r[1622]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \logix.ram_r[1623]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \logix.ram_r[1624]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \logix.ram_r[1625]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \logix.ram_r[1626]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \logix.ram_r[1627]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \logix.ram_r[1628]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \logix.ram_r[1629]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \logix.ram_r[162]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \logix.ram_r[1630]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \logix.ram_r[1631]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \logix.ram_r[1632]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \logix.ram_r[1633]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \logix.ram_r[1634]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \logix.ram_r[1635]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \logix.ram_r[1636]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \logix.ram_r[1637]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \logix.ram_r[1638]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \logix.ram_r[1639]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \logix.ram_r[163]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \logix.ram_r[1640]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \logix.ram_r[1641]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \logix.ram_r[1642]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \logix.ram_r[1643]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \logix.ram_r[1644]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \logix.ram_r[1645]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \logix.ram_r[1646]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \logix.ram_r[1647]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \logix.ram_r[1648]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \logix.ram_r[1649]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \logix.ram_r[164]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \logix.ram_r[1650]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \logix.ram_r[1651]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \logix.ram_r[1652]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \logix.ram_r[1653]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \logix.ram_r[1654]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \logix.ram_r[1655]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \logix.ram_r[1656]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \logix.ram_r[1657]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \logix.ram_r[1658]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \logix.ram_r[1659]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \logix.ram_r[165]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \logix.ram_r[1660]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \logix.ram_r[1661]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \logix.ram_r[1662]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \logix.ram_r[1663]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \logix.ram_r[1664]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \logix.ram_r[1665]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \logix.ram_r[1666]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \logix.ram_r[1667]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \logix.ram_r[1668]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \logix.ram_r[1669]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \logix.ram_r[166]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \logix.ram_r[1670]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \logix.ram_r[1671]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \logix.ram_r[1672]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \logix.ram_r[1673]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \logix.ram_r[1674]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \logix.ram_r[1675]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \logix.ram_r[1676]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \logix.ram_r[1677]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \logix.ram_r[1678]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \logix.ram_r[1679]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \logix.ram_r[167]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \logix.ram_r[1680]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \logix.ram_r[1681]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \logix.ram_r[1682]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \logix.ram_r[1683]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \logix.ram_r[1684]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \logix.ram_r[1685]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \logix.ram_r[1686]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \logix.ram_r[1687]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \logix.ram_r[1688]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \logix.ram_r[1689]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \logix.ram_r[168]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \logix.ram_r[1690]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \logix.ram_r[1691]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \logix.ram_r[1692]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \logix.ram_r[1693]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \logix.ram_r[1694]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \logix.ram_r[1695]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \logix.ram_r[1696]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \logix.ram_r[1697]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \logix.ram_r[1698]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \logix.ram_r[1699]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \logix.ram_r[169]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \logix.ram_r[16]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \logix.ram_r[1700]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \logix.ram_r[1701]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \logix.ram_r[1702]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \logix.ram_r[1703]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \logix.ram_r[1704]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \logix.ram_r[1705]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \logix.ram_r[1706]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \logix.ram_r[1707]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \logix.ram_r[1708]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \logix.ram_r[1709]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \logix.ram_r[170]$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \logix.ram_r[1710]$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \logix.ram_r[1711]$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \logix.ram_r[1712]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \logix.ram_r[1713]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \logix.ram_r[1714]$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \logix.ram_r[1715]$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \logix.ram_r[1716]$_DFFE_PP__1593  (.L_HI(net1593));
 sg13g2_tiehi \logix.ram_r[1717]$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \logix.ram_r[1718]$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \logix.ram_r[1719]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \logix.ram_r[171]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \logix.ram_r[1720]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \logix.ram_r[1721]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \logix.ram_r[1722]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \logix.ram_r[1723]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \logix.ram_r[1724]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \logix.ram_r[1725]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \logix.ram_r[1726]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \logix.ram_r[1727]$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \logix.ram_r[1728]$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \logix.ram_r[1729]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \logix.ram_r[172]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \logix.ram_r[1730]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \logix.ram_r[1731]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \logix.ram_r[1732]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \logix.ram_r[1733]$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \logix.ram_r[1734]$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \logix.ram_r[1735]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \logix.ram_r[1736]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \logix.ram_r[1737]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \logix.ram_r[1738]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \logix.ram_r[1739]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \logix.ram_r[173]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \logix.ram_r[1740]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \logix.ram_r[1741]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \logix.ram_r[1742]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \logix.ram_r[1743]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \logix.ram_r[1744]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \logix.ram_r[1745]$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \logix.ram_r[1746]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \logix.ram_r[1747]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \logix.ram_r[1748]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \logix.ram_r[1749]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \logix.ram_r[174]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \logix.ram_r[1750]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \logix.ram_r[1751]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \logix.ram_r[1752]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \logix.ram_r[1753]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \logix.ram_r[1754]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \logix.ram_r[1755]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \logix.ram_r[1756]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \logix.ram_r[1757]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \logix.ram_r[1758]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \logix.ram_r[1759]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \logix.ram_r[175]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \logix.ram_r[1760]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \logix.ram_r[1761]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \logix.ram_r[1762]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \logix.ram_r[1763]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \logix.ram_r[1764]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \logix.ram_r[1765]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \logix.ram_r[1766]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \logix.ram_r[1767]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \logix.ram_r[1768]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \logix.ram_r[1769]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \logix.ram_r[176]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \logix.ram_r[1770]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \logix.ram_r[1771]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \logix.ram_r[1772]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \logix.ram_r[1773]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \logix.ram_r[1774]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \logix.ram_r[1775]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \logix.ram_r[1776]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \logix.ram_r[1777]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \logix.ram_r[1778]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \logix.ram_r[1779]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \logix.ram_r[177]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \logix.ram_r[1780]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \logix.ram_r[1781]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \logix.ram_r[1782]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \logix.ram_r[1783]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \logix.ram_r[1784]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \logix.ram_r[1785]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \logix.ram_r[1786]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \logix.ram_r[1787]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \logix.ram_r[1788]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \logix.ram_r[1789]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \logix.ram_r[178]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \logix.ram_r[1790]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \logix.ram_r[1791]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \logix.ram_r[1792]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \logix.ram_r[1793]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \logix.ram_r[1794]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \logix.ram_r[1795]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \logix.ram_r[1796]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \logix.ram_r[1797]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \logix.ram_r[1798]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \logix.ram_r[1799]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \logix.ram_r[179]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \logix.ram_r[17]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \logix.ram_r[1800]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \logix.ram_r[1801]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \logix.ram_r[1802]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \logix.ram_r[1803]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \logix.ram_r[1804]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \logix.ram_r[1805]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \logix.ram_r[1806]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \logix.ram_r[1807]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \logix.ram_r[1808]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \logix.ram_r[1809]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \logix.ram_r[180]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \logix.ram_r[1810]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \logix.ram_r[1811]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \logix.ram_r[1812]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \logix.ram_r[1813]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \logix.ram_r[1814]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \logix.ram_r[1815]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \logix.ram_r[1816]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \logix.ram_r[1817]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \logix.ram_r[1818]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \logix.ram_r[1819]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \logix.ram_r[181]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \logix.ram_r[1820]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \logix.ram_r[1821]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \logix.ram_r[1822]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \logix.ram_r[1823]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \logix.ram_r[1824]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \logix.ram_r[1825]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \logix.ram_r[1826]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \logix.ram_r[1827]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \logix.ram_r[1828]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \logix.ram_r[1829]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \logix.ram_r[182]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \logix.ram_r[1830]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \logix.ram_r[1831]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \logix.ram_r[1832]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \logix.ram_r[1833]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \logix.ram_r[1834]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \logix.ram_r[1835]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \logix.ram_r[1836]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \logix.ram_r[1837]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \logix.ram_r[1838]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \logix.ram_r[1839]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \logix.ram_r[183]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \logix.ram_r[1840]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \logix.ram_r[1841]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \logix.ram_r[1842]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \logix.ram_r[1843]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \logix.ram_r[1844]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \logix.ram_r[1845]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \logix.ram_r[1846]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \logix.ram_r[1847]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \logix.ram_r[1848]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \logix.ram_r[1849]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \logix.ram_r[184]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \logix.ram_r[1850]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \logix.ram_r[1851]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \logix.ram_r[1852]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \logix.ram_r[1853]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \logix.ram_r[1854]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \logix.ram_r[1855]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \logix.ram_r[1856]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \logix.ram_r[1857]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \logix.ram_r[1858]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \logix.ram_r[1859]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \logix.ram_r[185]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \logix.ram_r[1860]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \logix.ram_r[1861]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \logix.ram_r[1862]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \logix.ram_r[1863]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \logix.ram_r[1864]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \logix.ram_r[1865]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \logix.ram_r[1866]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \logix.ram_r[1867]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \logix.ram_r[1868]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \logix.ram_r[1869]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \logix.ram_r[186]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \logix.ram_r[1870]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \logix.ram_r[1871]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \logix.ram_r[1872]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \logix.ram_r[1873]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \logix.ram_r[1874]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \logix.ram_r[1875]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \logix.ram_r[1876]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \logix.ram_r[1877]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \logix.ram_r[1878]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \logix.ram_r[1879]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \logix.ram_r[187]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \logix.ram_r[1880]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \logix.ram_r[1881]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \logix.ram_r[1882]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \logix.ram_r[1883]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \logix.ram_r[1884]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \logix.ram_r[1885]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \logix.ram_r[1886]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \logix.ram_r[1887]$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \logix.ram_r[1888]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \logix.ram_r[1889]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \logix.ram_r[188]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \logix.ram_r[1890]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \logix.ram_r[1891]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \logix.ram_r[1892]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \logix.ram_r[1893]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \logix.ram_r[1894]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \logix.ram_r[1895]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \logix.ram_r[1896]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \logix.ram_r[1897]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \logix.ram_r[1898]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \logix.ram_r[1899]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \logix.ram_r[189]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \logix.ram_r[18]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \logix.ram_r[1900]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \logix.ram_r[1901]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \logix.ram_r[1902]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \logix.ram_r[1903]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \logix.ram_r[1904]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \logix.ram_r[1905]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \logix.ram_r[1906]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \logix.ram_r[1907]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \logix.ram_r[1908]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \logix.ram_r[1909]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \logix.ram_r[190]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \logix.ram_r[1910]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \logix.ram_r[1911]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \logix.ram_r[1912]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \logix.ram_r[1913]$_DFFE_PP__1812  (.L_HI(net1812));
 sg13g2_tiehi \logix.ram_r[1914]$_DFFE_PP__1813  (.L_HI(net1813));
 sg13g2_tiehi \logix.ram_r[1915]$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \logix.ram_r[1916]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \logix.ram_r[1917]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \logix.ram_r[1918]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \logix.ram_r[1919]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \logix.ram_r[191]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \logix.ram_r[1920]$_DFFE_PP__1820  (.L_HI(net1820));
 sg13g2_tiehi \logix.ram_r[1921]$_DFFE_PP__1821  (.L_HI(net1821));
 sg13g2_tiehi \logix.ram_r[1922]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \logix.ram_r[1923]$_DFFE_PP__1823  (.L_HI(net1823));
 sg13g2_tiehi \logix.ram_r[1924]$_DFFE_PP__1824  (.L_HI(net1824));
 sg13g2_tiehi \logix.ram_r[1925]$_DFFE_PP__1825  (.L_HI(net1825));
 sg13g2_tiehi \logix.ram_r[1926]$_DFFE_PP__1826  (.L_HI(net1826));
 sg13g2_tiehi \logix.ram_r[1927]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \logix.ram_r[1928]$_DFFE_PP__1828  (.L_HI(net1828));
 sg13g2_tiehi \logix.ram_r[1929]$_DFFE_PP__1829  (.L_HI(net1829));
 sg13g2_tiehi \logix.ram_r[192]$_DFFE_PP__1830  (.L_HI(net1830));
 sg13g2_tiehi \logix.ram_r[1930]$_DFFE_PP__1831  (.L_HI(net1831));
 sg13g2_tiehi \logix.ram_r[1931]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \logix.ram_r[1932]$_DFFE_PP__1833  (.L_HI(net1833));
 sg13g2_tiehi \logix.ram_r[1933]$_DFFE_PP__1834  (.L_HI(net1834));
 sg13g2_tiehi \logix.ram_r[1934]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \logix.ram_r[1935]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \logix.ram_r[1936]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \logix.ram_r[1937]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \logix.ram_r[1938]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \logix.ram_r[1939]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \logix.ram_r[193]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \logix.ram_r[1940]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \logix.ram_r[1941]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \logix.ram_r[1942]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \logix.ram_r[1943]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \logix.ram_r[1944]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \logix.ram_r[1945]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \logix.ram_r[1946]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \logix.ram_r[1947]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \logix.ram_r[1948]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \logix.ram_r[1949]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \logix.ram_r[194]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \logix.ram_r[1950]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \logix.ram_r[1951]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \logix.ram_r[1952]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \logix.ram_r[1953]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \logix.ram_r[1954]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \logix.ram_r[1955]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \logix.ram_r[1956]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \logix.ram_r[1957]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \logix.ram_r[1958]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \logix.ram_r[1959]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \logix.ram_r[195]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \logix.ram_r[1960]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \logix.ram_r[1961]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \logix.ram_r[1962]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \logix.ram_r[1963]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \logix.ram_r[1964]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \logix.ram_r[1965]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \logix.ram_r[1966]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \logix.ram_r[1967]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \logix.ram_r[1968]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \logix.ram_r[1969]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \logix.ram_r[196]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \logix.ram_r[1970]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \logix.ram_r[1971]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \logix.ram_r[1972]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \logix.ram_r[1973]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \logix.ram_r[1974]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \logix.ram_r[1975]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \logix.ram_r[1976]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \logix.ram_r[1977]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \logix.ram_r[1978]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \logix.ram_r[1979]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \logix.ram_r[197]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \logix.ram_r[1980]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \logix.ram_r[1981]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \logix.ram_r[1982]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \logix.ram_r[1983]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \logix.ram_r[1984]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \logix.ram_r[1985]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \logix.ram_r[1986]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \logix.ram_r[1987]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \logix.ram_r[1988]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \logix.ram_r[1989]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \logix.ram_r[198]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \logix.ram_r[1990]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \logix.ram_r[1991]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \logix.ram_r[1992]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \logix.ram_r[1993]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \logix.ram_r[1994]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \logix.ram_r[1995]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \logix.ram_r[1996]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \logix.ram_r[1997]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \logix.ram_r[1998]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \logix.ram_r[1999]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \logix.ram_r[199]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \logix.ram_r[19]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \logix.ram_r[1]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \logix.ram_r[2000]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \logix.ram_r[2001]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \logix.ram_r[2002]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \logix.ram_r[2003]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \logix.ram_r[2004]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \logix.ram_r[2005]$_DFFE_PP__1915  (.L_HI(net1915));
 sg13g2_tiehi \logix.ram_r[2006]$_DFFE_PP__1916  (.L_HI(net1916));
 sg13g2_tiehi \logix.ram_r[2007]$_DFFE_PP__1917  (.L_HI(net1917));
 sg13g2_tiehi \logix.ram_r[2008]$_DFFE_PP__1918  (.L_HI(net1918));
 sg13g2_tiehi \logix.ram_r[2009]$_DFFE_PP__1919  (.L_HI(net1919));
 sg13g2_tiehi \logix.ram_r[200]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \logix.ram_r[2010]$_DFFE_PP__1921  (.L_HI(net1921));
 sg13g2_tiehi \logix.ram_r[2011]$_DFFE_PP__1922  (.L_HI(net1922));
 sg13g2_tiehi \logix.ram_r[2012]$_DFFE_PP__1923  (.L_HI(net1923));
 sg13g2_tiehi \logix.ram_r[2013]$_DFFE_PP__1924  (.L_HI(net1924));
 sg13g2_tiehi \logix.ram_r[2014]$_DFFE_PP__1925  (.L_HI(net1925));
 sg13g2_tiehi \logix.ram_r[2015]$_DFFE_PP__1926  (.L_HI(net1926));
 sg13g2_tiehi \logix.ram_r[2016]$_DFFE_PP__1927  (.L_HI(net1927));
 sg13g2_tiehi \logix.ram_r[2017]$_DFFE_PP__1928  (.L_HI(net1928));
 sg13g2_tiehi \logix.ram_r[2018]$_DFFE_PP__1929  (.L_HI(net1929));
 sg13g2_tiehi \logix.ram_r[2019]$_DFFE_PP__1930  (.L_HI(net1930));
 sg13g2_tiehi \logix.ram_r[201]$_DFFE_PP__1931  (.L_HI(net1931));
 sg13g2_tiehi \logix.ram_r[2020]$_DFFE_PP__1932  (.L_HI(net1932));
 sg13g2_tiehi \logix.ram_r[2021]$_DFFE_PP__1933  (.L_HI(net1933));
 sg13g2_tiehi \logix.ram_r[2022]$_DFFE_PP__1934  (.L_HI(net1934));
 sg13g2_tiehi \logix.ram_r[2023]$_DFFE_PP__1935  (.L_HI(net1935));
 sg13g2_tiehi \logix.ram_r[2024]$_DFFE_PP__1936  (.L_HI(net1936));
 sg13g2_tiehi \logix.ram_r[2025]$_DFFE_PP__1937  (.L_HI(net1937));
 sg13g2_tiehi \logix.ram_r[2026]$_DFFE_PP__1938  (.L_HI(net1938));
 sg13g2_tiehi \logix.ram_r[2027]$_DFFE_PP__1939  (.L_HI(net1939));
 sg13g2_tiehi \logix.ram_r[2028]$_DFFE_PP__1940  (.L_HI(net1940));
 sg13g2_tiehi \logix.ram_r[2029]$_DFFE_PP__1941  (.L_HI(net1941));
 sg13g2_tiehi \logix.ram_r[202]$_DFFE_PP__1942  (.L_HI(net1942));
 sg13g2_tiehi \logix.ram_r[2030]$_DFFE_PP__1943  (.L_HI(net1943));
 sg13g2_tiehi \logix.ram_r[2031]$_DFFE_PP__1944  (.L_HI(net1944));
 sg13g2_tiehi \logix.ram_r[2032]$_DFFE_PP__1945  (.L_HI(net1945));
 sg13g2_tiehi \logix.ram_r[2033]$_DFFE_PP__1946  (.L_HI(net1946));
 sg13g2_tiehi \logix.ram_r[2034]$_DFFE_PP__1947  (.L_HI(net1947));
 sg13g2_tiehi \logix.ram_r[2035]$_DFFE_PP__1948  (.L_HI(net1948));
 sg13g2_tiehi \logix.ram_r[2036]$_DFFE_PP__1949  (.L_HI(net1949));
 sg13g2_tiehi \logix.ram_r[2037]$_DFFE_PP__1950  (.L_HI(net1950));
 sg13g2_tiehi \logix.ram_r[2038]$_DFFE_PP__1951  (.L_HI(net1951));
 sg13g2_tiehi \logix.ram_r[2039]$_DFFE_PP__1952  (.L_HI(net1952));
 sg13g2_tiehi \logix.ram_r[203]$_DFFE_PP__1953  (.L_HI(net1953));
 sg13g2_tiehi \logix.ram_r[2040]$_DFFE_PP__1954  (.L_HI(net1954));
 sg13g2_tiehi \logix.ram_r[2041]$_DFFE_PP__1955  (.L_HI(net1955));
 sg13g2_tiehi \logix.ram_r[2042]$_DFFE_PP__1956  (.L_HI(net1956));
 sg13g2_tiehi \logix.ram_r[2043]$_DFFE_PP__1957  (.L_HI(net1957));
 sg13g2_tiehi \logix.ram_r[2044]$_DFFE_PP__1958  (.L_HI(net1958));
 sg13g2_tiehi \logix.ram_r[2045]$_DFFE_PP__1959  (.L_HI(net1959));
 sg13g2_tiehi \logix.ram_r[2046]$_DFFE_PP__1960  (.L_HI(net1960));
 sg13g2_tiehi \logix.ram_r[2047]$_DFFE_PP__1961  (.L_HI(net1961));
 sg13g2_tiehi \logix.ram_r[2048]$_DFFE_PP__1962  (.L_HI(net1962));
 sg13g2_tiehi \logix.ram_r[2049]$_DFFE_PP__1963  (.L_HI(net1963));
 sg13g2_tiehi \logix.ram_r[204]$_DFFE_PP__1964  (.L_HI(net1964));
 sg13g2_tiehi \logix.ram_r[2050]$_DFFE_PP__1965  (.L_HI(net1965));
 sg13g2_tiehi \logix.ram_r[2051]$_DFFE_PP__1966  (.L_HI(net1966));
 sg13g2_tiehi \logix.ram_r[2052]$_DFFE_PP__1967  (.L_HI(net1967));
 sg13g2_tiehi \logix.ram_r[2053]$_DFFE_PP__1968  (.L_HI(net1968));
 sg13g2_tiehi \logix.ram_r[2054]$_DFFE_PP__1969  (.L_HI(net1969));
 sg13g2_tiehi \logix.ram_r[2055]$_DFFE_PP__1970  (.L_HI(net1970));
 sg13g2_tiehi \logix.ram_r[205]$_DFFE_PP__1971  (.L_HI(net1971));
 sg13g2_tiehi \logix.ram_r[206]$_DFFE_PP__1972  (.L_HI(net1972));
 sg13g2_tiehi \logix.ram_r[207]$_DFFE_PP__1973  (.L_HI(net1973));
 sg13g2_tiehi \logix.ram_r[208]$_DFFE_PP__1974  (.L_HI(net1974));
 sg13g2_tiehi \logix.ram_r[209]$_DFFE_PP__1975  (.L_HI(net1975));
 sg13g2_tiehi \logix.ram_r[20]$_DFFE_PP__1976  (.L_HI(net1976));
 sg13g2_tiehi \logix.ram_r[210]$_DFFE_PP__1977  (.L_HI(net1977));
 sg13g2_tiehi \logix.ram_r[211]$_DFFE_PP__1978  (.L_HI(net1978));
 sg13g2_tiehi \logix.ram_r[212]$_DFFE_PP__1979  (.L_HI(net1979));
 sg13g2_tiehi \logix.ram_r[213]$_DFFE_PP__1980  (.L_HI(net1980));
 sg13g2_tiehi \logix.ram_r[214]$_DFFE_PP__1981  (.L_HI(net1981));
 sg13g2_tiehi \logix.ram_r[215]$_DFFE_PP__1982  (.L_HI(net1982));
 sg13g2_tiehi \logix.ram_r[216]$_DFFE_PP__1983  (.L_HI(net1983));
 sg13g2_tiehi \logix.ram_r[217]$_DFFE_PP__1984  (.L_HI(net1984));
 sg13g2_tiehi \logix.ram_r[218]$_DFFE_PP__1985  (.L_HI(net1985));
 sg13g2_tiehi \logix.ram_r[219]$_DFFE_PP__1986  (.L_HI(net1986));
 sg13g2_tiehi \logix.ram_r[21]$_DFFE_PP__1987  (.L_HI(net1987));
 sg13g2_tiehi \logix.ram_r[220]$_DFFE_PP__1988  (.L_HI(net1988));
 sg13g2_tiehi \logix.ram_r[221]$_DFFE_PP__1989  (.L_HI(net1989));
 sg13g2_tiehi \logix.ram_r[222]$_DFFE_PP__1990  (.L_HI(net1990));
 sg13g2_tiehi \logix.ram_r[223]$_DFFE_PP__1991  (.L_HI(net1991));
 sg13g2_tiehi \logix.ram_r[224]$_DFFE_PP__1992  (.L_HI(net1992));
 sg13g2_tiehi \logix.ram_r[225]$_DFFE_PP__1993  (.L_HI(net1993));
 sg13g2_tiehi \logix.ram_r[226]$_DFFE_PP__1994  (.L_HI(net1994));
 sg13g2_tiehi \logix.ram_r[227]$_DFFE_PP__1995  (.L_HI(net1995));
 sg13g2_tiehi \logix.ram_r[228]$_DFFE_PP__1996  (.L_HI(net1996));
 sg13g2_tiehi \logix.ram_r[229]$_DFFE_PP__1997  (.L_HI(net1997));
 sg13g2_tiehi \logix.ram_r[22]$_DFFE_PP__1998  (.L_HI(net1998));
 sg13g2_tiehi \logix.ram_r[230]$_DFFE_PP__1999  (.L_HI(net1999));
 sg13g2_tiehi \logix.ram_r[231]$_DFFE_PP__2000  (.L_HI(net2000));
 sg13g2_tiehi \logix.ram_r[232]$_DFFE_PP__2001  (.L_HI(net2001));
 sg13g2_tiehi \logix.ram_r[233]$_DFFE_PP__2002  (.L_HI(net2002));
 sg13g2_tiehi \logix.ram_r[234]$_DFFE_PP__2003  (.L_HI(net2003));
 sg13g2_tiehi \logix.ram_r[235]$_DFFE_PP__2004  (.L_HI(net2004));
 sg13g2_tiehi \logix.ram_r[236]$_DFFE_PP__2005  (.L_HI(net2005));
 sg13g2_tiehi \logix.ram_r[237]$_DFFE_PP__2006  (.L_HI(net2006));
 sg13g2_tiehi \logix.ram_r[238]$_DFFE_PP__2007  (.L_HI(net2007));
 sg13g2_tiehi \logix.ram_r[239]$_DFFE_PP__2008  (.L_HI(net2008));
 sg13g2_tiehi \logix.ram_r[23]$_DFFE_PP__2009  (.L_HI(net2009));
 sg13g2_tiehi \logix.ram_r[240]$_DFFE_PP__2010  (.L_HI(net2010));
 sg13g2_tiehi \logix.ram_r[241]$_DFFE_PP__2011  (.L_HI(net2011));
 sg13g2_tiehi \logix.ram_r[242]$_DFFE_PP__2012  (.L_HI(net2012));
 sg13g2_tiehi \logix.ram_r[243]$_DFFE_PP__2013  (.L_HI(net2013));
 sg13g2_tiehi \logix.ram_r[244]$_DFFE_PP__2014  (.L_HI(net2014));
 sg13g2_tiehi \logix.ram_r[245]$_DFFE_PP__2015  (.L_HI(net2015));
 sg13g2_tiehi \logix.ram_r[246]$_DFFE_PP__2016  (.L_HI(net2016));
 sg13g2_tiehi \logix.ram_r[247]$_DFFE_PP__2017  (.L_HI(net2017));
 sg13g2_tiehi \logix.ram_r[248]$_DFFE_PP__2018  (.L_HI(net2018));
 sg13g2_tiehi \logix.ram_r[249]$_DFFE_PP__2019  (.L_HI(net2019));
 sg13g2_tiehi \logix.ram_r[24]$_DFFE_PP__2020  (.L_HI(net2020));
 sg13g2_tiehi \logix.ram_r[250]$_DFFE_PP__2021  (.L_HI(net2021));
 sg13g2_tiehi \logix.ram_r[251]$_DFFE_PP__2022  (.L_HI(net2022));
 sg13g2_tiehi \logix.ram_r[252]$_DFFE_PP__2023  (.L_HI(net2023));
 sg13g2_tiehi \logix.ram_r[253]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \logix.ram_r[254]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \logix.ram_r[255]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \logix.ram_r[256]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \logix.ram_r[257]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \logix.ram_r[258]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \logix.ram_r[259]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \logix.ram_r[25]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \logix.ram_r[260]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \logix.ram_r[261]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \logix.ram_r[262]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \logix.ram_r[263]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \logix.ram_r[264]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \logix.ram_r[265]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \logix.ram_r[266]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \logix.ram_r[267]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \logix.ram_r[268]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \logix.ram_r[269]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \logix.ram_r[26]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \logix.ram_r[270]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \logix.ram_r[271]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \logix.ram_r[272]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \logix.ram_r[273]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \logix.ram_r[274]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \logix.ram_r[275]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \logix.ram_r[276]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \logix.ram_r[277]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \logix.ram_r[278]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \logix.ram_r[279]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \logix.ram_r[27]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \logix.ram_r[280]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \logix.ram_r[281]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \logix.ram_r[282]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \logix.ram_r[283]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \logix.ram_r[284]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \logix.ram_r[285]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \logix.ram_r[286]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \logix.ram_r[287]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \logix.ram_r[288]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \logix.ram_r[289]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \logix.ram_r[28]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \logix.ram_r[290]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \logix.ram_r[291]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \logix.ram_r[292]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \logix.ram_r[293]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \logix.ram_r[294]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \logix.ram_r[295]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \logix.ram_r[296]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \logix.ram_r[297]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \logix.ram_r[298]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \logix.ram_r[299]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \logix.ram_r[29]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \logix.ram_r[2]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \logix.ram_r[300]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \logix.ram_r[301]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \logix.ram_r[302]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \logix.ram_r[303]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \logix.ram_r[304]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \logix.ram_r[305]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \logix.ram_r[306]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \logix.ram_r[307]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \logix.ram_r[308]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \logix.ram_r[309]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \logix.ram_r[30]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \logix.ram_r[310]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \logix.ram_r[311]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \logix.ram_r[312]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \logix.ram_r[313]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \logix.ram_r[314]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \logix.ram_r[315]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \logix.ram_r[316]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \logix.ram_r[317]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \logix.ram_r[318]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \logix.ram_r[319]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \logix.ram_r[31]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \logix.ram_r[320]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \logix.ram_r[321]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \logix.ram_r[322]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \logix.ram_r[323]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \logix.ram_r[324]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \logix.ram_r[325]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \logix.ram_r[326]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \logix.ram_r[327]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \logix.ram_r[328]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \logix.ram_r[329]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \logix.ram_r[32]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \logix.ram_r[330]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \logix.ram_r[331]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \logix.ram_r[332]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \logix.ram_r[333]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \logix.ram_r[334]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \logix.ram_r[335]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \logix.ram_r[336]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \logix.ram_r[337]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \logix.ram_r[338]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \logix.ram_r[339]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \logix.ram_r[33]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \logix.ram_r[340]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \logix.ram_r[341]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \logix.ram_r[342]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \logix.ram_r[343]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \logix.ram_r[344]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \logix.ram_r[345]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \logix.ram_r[346]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \logix.ram_r[347]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \logix.ram_r[348]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \logix.ram_r[349]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \logix.ram_r[34]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \logix.ram_r[350]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \logix.ram_r[351]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \logix.ram_r[352]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \logix.ram_r[353]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \logix.ram_r[354]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \logix.ram_r[355]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \logix.ram_r[356]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \logix.ram_r[357]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \logix.ram_r[358]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \logix.ram_r[359]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \logix.ram_r[35]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \logix.ram_r[360]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \logix.ram_r[361]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \logix.ram_r[362]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \logix.ram_r[363]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \logix.ram_r[364]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \logix.ram_r[365]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \logix.ram_r[366]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \logix.ram_r[367]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \logix.ram_r[368]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \logix.ram_r[369]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \logix.ram_r[36]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \logix.ram_r[370]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \logix.ram_r[371]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \logix.ram_r[372]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \logix.ram_r[373]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \logix.ram_r[374]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \logix.ram_r[375]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \logix.ram_r[376]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \logix.ram_r[377]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \logix.ram_r[378]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \logix.ram_r[379]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \logix.ram_r[37]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \logix.ram_r[380]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \logix.ram_r[381]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \logix.ram_r[382]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \logix.ram_r[383]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \logix.ram_r[384]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \logix.ram_r[385]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \logix.ram_r[386]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \logix.ram_r[387]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \logix.ram_r[388]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \logix.ram_r[389]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \logix.ram_r[38]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \logix.ram_r[390]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \logix.ram_r[391]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \logix.ram_r[392]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \logix.ram_r[393]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \logix.ram_r[394]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \logix.ram_r[395]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \logix.ram_r[396]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \logix.ram_r[397]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \logix.ram_r[398]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \logix.ram_r[399]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \logix.ram_r[39]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \logix.ram_r[3]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \logix.ram_r[400]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \logix.ram_r[401]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \logix.ram_r[402]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \logix.ram_r[403]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \logix.ram_r[404]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \logix.ram_r[405]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \logix.ram_r[406]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \logix.ram_r[407]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \logix.ram_r[408]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \logix.ram_r[409]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \logix.ram_r[40]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \logix.ram_r[410]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \logix.ram_r[411]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \logix.ram_r[412]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \logix.ram_r[413]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \logix.ram_r[414]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \logix.ram_r[415]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \logix.ram_r[416]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \logix.ram_r[417]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \logix.ram_r[418]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \logix.ram_r[419]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \logix.ram_r[41]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \logix.ram_r[420]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \logix.ram_r[421]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \logix.ram_r[422]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \logix.ram_r[423]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \logix.ram_r[424]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \logix.ram_r[425]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \logix.ram_r[426]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \logix.ram_r[427]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \logix.ram_r[428]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \logix.ram_r[429]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \logix.ram_r[42]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \logix.ram_r[430]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \logix.ram_r[431]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \logix.ram_r[432]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \logix.ram_r[433]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \logix.ram_r[434]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \logix.ram_r[435]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \logix.ram_r[436]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \logix.ram_r[437]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \logix.ram_r[438]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \logix.ram_r[439]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \logix.ram_r[43]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \logix.ram_r[440]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \logix.ram_r[441]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \logix.ram_r[442]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \logix.ram_r[443]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \logix.ram_r[444]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \logix.ram_r[445]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \logix.ram_r[446]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \logix.ram_r[447]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \logix.ram_r[448]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \logix.ram_r[449]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \logix.ram_r[44]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \logix.ram_r[450]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \logix.ram_r[451]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \logix.ram_r[452]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \logix.ram_r[453]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \logix.ram_r[454]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \logix.ram_r[455]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \logix.ram_r[456]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \logix.ram_r[457]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \logix.ram_r[458]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \logix.ram_r[459]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \logix.ram_r[45]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \logix.ram_r[460]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \logix.ram_r[461]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \logix.ram_r[462]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \logix.ram_r[463]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \logix.ram_r[464]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \logix.ram_r[465]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \logix.ram_r[466]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \logix.ram_r[467]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \logix.ram_r[468]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \logix.ram_r[469]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \logix.ram_r[46]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \logix.ram_r[470]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \logix.ram_r[471]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \logix.ram_r[472]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \logix.ram_r[473]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \logix.ram_r[474]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \logix.ram_r[475]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \logix.ram_r[476]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \logix.ram_r[477]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \logix.ram_r[478]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \logix.ram_r[479]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \logix.ram_r[47]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \logix.ram_r[480]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \logix.ram_r[481]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \logix.ram_r[482]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \logix.ram_r[483]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \logix.ram_r[484]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \logix.ram_r[485]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \logix.ram_r[486]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \logix.ram_r[487]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \logix.ram_r[488]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \logix.ram_r[489]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \logix.ram_r[48]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \logix.ram_r[490]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \logix.ram_r[491]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \logix.ram_r[492]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \logix.ram_r[493]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \logix.ram_r[494]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \logix.ram_r[495]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \logix.ram_r[496]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \logix.ram_r[497]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \logix.ram_r[498]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \logix.ram_r[499]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \logix.ram_r[49]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \logix.ram_r[4]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \logix.ram_r[500]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \logix.ram_r[501]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \logix.ram_r[502]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \logix.ram_r[503]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \logix.ram_r[504]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \logix.ram_r[505]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \logix.ram_r[506]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \logix.ram_r[507]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \logix.ram_r[508]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \logix.ram_r[509]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \logix.ram_r[50]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \logix.ram_r[510]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \logix.ram_r[511]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \logix.ram_r[512]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \logix.ram_r[513]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \logix.ram_r[514]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \logix.ram_r[515]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \logix.ram_r[516]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \logix.ram_r[517]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \logix.ram_r[518]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \logix.ram_r[519]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \logix.ram_r[51]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \logix.ram_r[520]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \logix.ram_r[521]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \logix.ram_r[522]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \logix.ram_r[523]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \logix.ram_r[524]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \logix.ram_r[525]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \logix.ram_r[526]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \logix.ram_r[527]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \logix.ram_r[528]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \logix.ram_r[529]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \logix.ram_r[52]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \logix.ram_r[530]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \logix.ram_r[531]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \logix.ram_r[532]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \logix.ram_r[533]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \logix.ram_r[534]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \logix.ram_r[535]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \logix.ram_r[536]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \logix.ram_r[537]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \logix.ram_r[538]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \logix.ram_r[539]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \logix.ram_r[53]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \logix.ram_r[540]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \logix.ram_r[541]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \logix.ram_r[542]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \logix.ram_r[543]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \logix.ram_r[544]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \logix.ram_r[545]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \logix.ram_r[546]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \logix.ram_r[547]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \logix.ram_r[548]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \logix.ram_r[549]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \logix.ram_r[54]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \logix.ram_r[550]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \logix.ram_r[551]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \logix.ram_r[552]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \logix.ram_r[553]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \logix.ram_r[554]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \logix.ram_r[555]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \logix.ram_r[556]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \logix.ram_r[557]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \logix.ram_r[558]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \logix.ram_r[559]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \logix.ram_r[55]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \logix.ram_r[560]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \logix.ram_r[561]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \logix.ram_r[562]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \logix.ram_r[563]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \logix.ram_r[564]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \logix.ram_r[565]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \logix.ram_r[566]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \logix.ram_r[567]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \logix.ram_r[568]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \logix.ram_r[569]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \logix.ram_r[56]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \logix.ram_r[570]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \logix.ram_r[571]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \logix.ram_r[572]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \logix.ram_r[573]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \logix.ram_r[574]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \logix.ram_r[575]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \logix.ram_r[576]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \logix.ram_r[577]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \logix.ram_r[578]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \logix.ram_r[579]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \logix.ram_r[57]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \logix.ram_r[580]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \logix.ram_r[581]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \logix.ram_r[582]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \logix.ram_r[583]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \logix.ram_r[584]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \logix.ram_r[585]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \logix.ram_r[586]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \logix.ram_r[587]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \logix.ram_r[588]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \logix.ram_r[589]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \logix.ram_r[58]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \logix.ram_r[590]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \logix.ram_r[591]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \logix.ram_r[592]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \logix.ram_r[593]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \logix.ram_r[594]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \logix.ram_r[595]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \logix.ram_r[596]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \logix.ram_r[597]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \logix.ram_r[598]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \logix.ram_r[599]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \logix.ram_r[59]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \logix.ram_r[5]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \logix.ram_r[600]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \logix.ram_r[601]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \logix.ram_r[602]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \logix.ram_r[603]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \logix.ram_r[604]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \logix.ram_r[605]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \logix.ram_r[606]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \logix.ram_r[607]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \logix.ram_r[608]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \logix.ram_r[609]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \logix.ram_r[60]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \logix.ram_r[610]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \logix.ram_r[611]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \logix.ram_r[612]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \logix.ram_r[613]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \logix.ram_r[614]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \logix.ram_r[615]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \logix.ram_r[616]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \logix.ram_r[617]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \logix.ram_r[618]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \logix.ram_r[619]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \logix.ram_r[61]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \logix.ram_r[620]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \logix.ram_r[621]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \logix.ram_r[622]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \logix.ram_r[623]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \logix.ram_r[624]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \logix.ram_r[625]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \logix.ram_r[626]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \logix.ram_r[627]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \logix.ram_r[628]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \logix.ram_r[629]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \logix.ram_r[62]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \logix.ram_r[630]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \logix.ram_r[631]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \logix.ram_r[632]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \logix.ram_r[633]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \logix.ram_r[634]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \logix.ram_r[635]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \logix.ram_r[636]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \logix.ram_r[637]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \logix.ram_r[638]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \logix.ram_r[639]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \logix.ram_r[63]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \logix.ram_r[640]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \logix.ram_r[641]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \logix.ram_r[642]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \logix.ram_r[643]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \logix.ram_r[644]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \logix.ram_r[645]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \logix.ram_r[646]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \logix.ram_r[647]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \logix.ram_r[648]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \logix.ram_r[649]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \logix.ram_r[64]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \logix.ram_r[650]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \logix.ram_r[651]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \logix.ram_r[652]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \logix.ram_r[653]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \logix.ram_r[654]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \logix.ram_r[655]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \logix.ram_r[656]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \logix.ram_r[657]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \logix.ram_r[658]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \logix.ram_r[659]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \logix.ram_r[65]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \logix.ram_r[660]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \logix.ram_r[661]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \logix.ram_r[662]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \logix.ram_r[663]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \logix.ram_r[664]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \logix.ram_r[665]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \logix.ram_r[666]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \logix.ram_r[667]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \logix.ram_r[668]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \logix.ram_r[669]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \logix.ram_r[66]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \logix.ram_r[670]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \logix.ram_r[671]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \logix.ram_r[672]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \logix.ram_r[673]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \logix.ram_r[674]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \logix.ram_r[675]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \logix.ram_r[676]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \logix.ram_r[677]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \logix.ram_r[678]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \logix.ram_r[679]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \logix.ram_r[67]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \logix.ram_r[680]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \logix.ram_r[681]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \logix.ram_r[682]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \logix.ram_r[683]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \logix.ram_r[684]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \logix.ram_r[685]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \logix.ram_r[686]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \logix.ram_r[687]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \logix.ram_r[688]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \logix.ram_r[689]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \logix.ram_r[68]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \logix.ram_r[690]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \logix.ram_r[691]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \logix.ram_r[692]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \logix.ram_r[693]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \logix.ram_r[694]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \logix.ram_r[695]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \logix.ram_r[696]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \logix.ram_r[697]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \logix.ram_r[698]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \logix.ram_r[699]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \logix.ram_r[69]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \logix.ram_r[6]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \logix.ram_r[700]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \logix.ram_r[701]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \logix.ram_r[702]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \logix.ram_r[703]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \logix.ram_r[704]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \logix.ram_r[705]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \logix.ram_r[706]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \logix.ram_r[707]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \logix.ram_r[708]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \logix.ram_r[709]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \logix.ram_r[70]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \logix.ram_r[710]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \logix.ram_r[711]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \logix.ram_r[712]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \logix.ram_r[713]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \logix.ram_r[714]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \logix.ram_r[715]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \logix.ram_r[716]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \logix.ram_r[717]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \logix.ram_r[718]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \logix.ram_r[719]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \logix.ram_r[71]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \logix.ram_r[720]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \logix.ram_r[721]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \logix.ram_r[722]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \logix.ram_r[723]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \logix.ram_r[724]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \logix.ram_r[725]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \logix.ram_r[726]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \logix.ram_r[727]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \logix.ram_r[728]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \logix.ram_r[729]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \logix.ram_r[72]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \logix.ram_r[730]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \logix.ram_r[731]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \logix.ram_r[732]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \logix.ram_r[733]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \logix.ram_r[734]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \logix.ram_r[735]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \logix.ram_r[736]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \logix.ram_r[737]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \logix.ram_r[738]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \logix.ram_r[739]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \logix.ram_r[73]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \logix.ram_r[740]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \logix.ram_r[741]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \logix.ram_r[742]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \logix.ram_r[743]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \logix.ram_r[744]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \logix.ram_r[745]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \logix.ram_r[746]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \logix.ram_r[747]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \logix.ram_r[748]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \logix.ram_r[749]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \logix.ram_r[74]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \logix.ram_r[750]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \logix.ram_r[751]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \logix.ram_r[752]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \logix.ram_r[753]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \logix.ram_r[754]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \logix.ram_r[755]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \logix.ram_r[756]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \logix.ram_r[757]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \logix.ram_r[758]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \logix.ram_r[759]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \logix.ram_r[75]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \logix.ram_r[760]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \logix.ram_r[761]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \logix.ram_r[762]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \logix.ram_r[763]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \logix.ram_r[764]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \logix.ram_r[765]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \logix.ram_r[766]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \logix.ram_r[767]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \logix.ram_r[768]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \logix.ram_r[769]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \logix.ram_r[76]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \logix.ram_r[770]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \logix.ram_r[771]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \logix.ram_r[772]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \logix.ram_r[773]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \logix.ram_r[774]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \logix.ram_r[775]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \logix.ram_r[776]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \logix.ram_r[777]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \logix.ram_r[778]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \logix.ram_r[779]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \logix.ram_r[77]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \logix.ram_r[780]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \logix.ram_r[781]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \logix.ram_r[782]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \logix.ram_r[783]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \logix.ram_r[784]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \logix.ram_r[785]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \logix.ram_r[786]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \logix.ram_r[787]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \logix.ram_r[788]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \logix.ram_r[789]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \logix.ram_r[78]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \logix.ram_r[790]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \logix.ram_r[791]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \logix.ram_r[792]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \logix.ram_r[793]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \logix.ram_r[794]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \logix.ram_r[795]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \logix.ram_r[796]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \logix.ram_r[797]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \logix.ram_r[798]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \logix.ram_r[799]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \logix.ram_r[79]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \logix.ram_r[7]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \logix.ram_r[800]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \logix.ram_r[801]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \logix.ram_r[802]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \logix.ram_r[803]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \logix.ram_r[804]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \logix.ram_r[805]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \logix.ram_r[806]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \logix.ram_r[807]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \logix.ram_r[808]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \logix.ram_r[809]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \logix.ram_r[80]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \logix.ram_r[810]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \logix.ram_r[811]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \logix.ram_r[812]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \logix.ram_r[813]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \logix.ram_r[814]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \logix.ram_r[815]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \logix.ram_r[816]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \logix.ram_r[817]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \logix.ram_r[818]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \logix.ram_r[819]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \logix.ram_r[81]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \logix.ram_r[820]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \logix.ram_r[821]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \logix.ram_r[822]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \logix.ram_r[823]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \logix.ram_r[824]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \logix.ram_r[825]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \logix.ram_r[826]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \logix.ram_r[827]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \logix.ram_r[828]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \logix.ram_r[829]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \logix.ram_r[82]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \logix.ram_r[830]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \logix.ram_r[831]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \logix.ram_r[832]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \logix.ram_r[833]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \logix.ram_r[834]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \logix.ram_r[835]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \logix.ram_r[836]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \logix.ram_r[837]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \logix.ram_r[838]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \logix.ram_r[839]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \logix.ram_r[83]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \logix.ram_r[840]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \logix.ram_r[841]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \logix.ram_r[842]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \logix.ram_r[843]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \logix.ram_r[844]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \logix.ram_r[845]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \logix.ram_r[846]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \logix.ram_r[847]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \logix.ram_r[848]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \logix.ram_r[849]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \logix.ram_r[84]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \logix.ram_r[850]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \logix.ram_r[851]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \logix.ram_r[852]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \logix.ram_r[853]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \logix.ram_r[854]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \logix.ram_r[855]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \logix.ram_r[856]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \logix.ram_r[857]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \logix.ram_r[858]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \logix.ram_r[859]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \logix.ram_r[85]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \logix.ram_r[860]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \logix.ram_r[861]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \logix.ram_r[862]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \logix.ram_r[863]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \logix.ram_r[864]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \logix.ram_r[865]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \logix.ram_r[866]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \logix.ram_r[867]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \logix.ram_r[868]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \logix.ram_r[869]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \logix.ram_r[86]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \logix.ram_r[870]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \logix.ram_r[871]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \logix.ram_r[872]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \logix.ram_r[873]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \logix.ram_r[874]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \logix.ram_r[875]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \logix.ram_r[876]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \logix.ram_r[877]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \logix.ram_r[878]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \logix.ram_r[879]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \logix.ram_r[87]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \logix.ram_r[880]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \logix.ram_r[881]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \logix.ram_r[882]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \logix.ram_r[883]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \logix.ram_r[884]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \logix.ram_r[885]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \logix.ram_r[886]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \logix.ram_r[887]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \logix.ram_r[888]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \logix.ram_r[889]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \logix.ram_r[88]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \logix.ram_r[890]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \logix.ram_r[891]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \logix.ram_r[892]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \logix.ram_r[893]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \logix.ram_r[894]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \logix.ram_r[895]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \logix.ram_r[896]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \logix.ram_r[897]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \logix.ram_r[898]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \logix.ram_r[899]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \logix.ram_r[89]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \logix.ram_r[8]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \logix.ram_r[900]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \logix.ram_r[901]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \logix.ram_r[902]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \logix.ram_r[903]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \logix.ram_r[904]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \logix.ram_r[905]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \logix.ram_r[906]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \logix.ram_r[907]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \logix.ram_r[908]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \logix.ram_r[909]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \logix.ram_r[90]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \logix.ram_r[910]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \logix.ram_r[911]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \logix.ram_r[912]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \logix.ram_r[913]$_DFFE_PP__2757  (.L_HI(net2757));
 sg13g2_tiehi \logix.ram_r[914]$_DFFE_PP__2758  (.L_HI(net2758));
 sg13g2_tiehi \logix.ram_r[915]$_DFFE_PP__2759  (.L_HI(net2759));
 sg13g2_tiehi \logix.ram_r[916]$_DFFE_PP__2760  (.L_HI(net2760));
 sg13g2_tiehi \logix.ram_r[917]$_DFFE_PP__2761  (.L_HI(net2761));
 sg13g2_tiehi \logix.ram_r[918]$_DFFE_PP__2762  (.L_HI(net2762));
 sg13g2_tiehi \logix.ram_r[919]$_DFFE_PP__2763  (.L_HI(net2763));
 sg13g2_tiehi \logix.ram_r[91]$_DFFE_PP__2764  (.L_HI(net2764));
 sg13g2_tiehi \logix.ram_r[920]$_DFFE_PP__2765  (.L_HI(net2765));
 sg13g2_tiehi \logix.ram_r[921]$_DFFE_PP__2766  (.L_HI(net2766));
 sg13g2_tiehi \logix.ram_r[922]$_DFFE_PP__2767  (.L_HI(net2767));
 sg13g2_tiehi \logix.ram_r[923]$_DFFE_PP__2768  (.L_HI(net2768));
 sg13g2_tiehi \logix.ram_r[924]$_DFFE_PP__2769  (.L_HI(net2769));
 sg13g2_tiehi \logix.ram_r[925]$_DFFE_PP__2770  (.L_HI(net2770));
 sg13g2_tiehi \logix.ram_r[926]$_DFFE_PP__2771  (.L_HI(net2771));
 sg13g2_tiehi \logix.ram_r[927]$_DFFE_PP__2772  (.L_HI(net2772));
 sg13g2_tiehi \logix.ram_r[928]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \logix.ram_r[929]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \logix.ram_r[92]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \logix.ram_r[930]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \logix.ram_r[931]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \logix.ram_r[932]$_DFFE_PP__2778  (.L_HI(net2778));
 sg13g2_tiehi \logix.ram_r[933]$_DFFE_PP__2779  (.L_HI(net2779));
 sg13g2_tiehi \logix.ram_r[934]$_DFFE_PP__2780  (.L_HI(net2780));
 sg13g2_tiehi \logix.ram_r[935]$_DFFE_PP__2781  (.L_HI(net2781));
 sg13g2_tiehi \logix.ram_r[936]$_DFFE_PP__2782  (.L_HI(net2782));
 sg13g2_tiehi \logix.ram_r[937]$_DFFE_PP__2783  (.L_HI(net2783));
 sg13g2_tiehi \logix.ram_r[938]$_DFFE_PP__2784  (.L_HI(net2784));
 sg13g2_tiehi \logix.ram_r[939]$_DFFE_PP__2785  (.L_HI(net2785));
 sg13g2_tiehi \logix.ram_r[93]$_DFFE_PP__2786  (.L_HI(net2786));
 sg13g2_tiehi \logix.ram_r[940]$_DFFE_PP__2787  (.L_HI(net2787));
 sg13g2_tiehi \logix.ram_r[941]$_DFFE_PP__2788  (.L_HI(net2788));
 sg13g2_tiehi \logix.ram_r[942]$_DFFE_PP__2789  (.L_HI(net2789));
 sg13g2_tiehi \logix.ram_r[943]$_DFFE_PP__2790  (.L_HI(net2790));
 sg13g2_tiehi \logix.ram_r[944]$_DFFE_PP__2791  (.L_HI(net2791));
 sg13g2_tiehi \logix.ram_r[945]$_DFFE_PP__2792  (.L_HI(net2792));
 sg13g2_tiehi \logix.ram_r[946]$_DFFE_PP__2793  (.L_HI(net2793));
 sg13g2_tiehi \logix.ram_r[947]$_DFFE_PP__2794  (.L_HI(net2794));
 sg13g2_tiehi \logix.ram_r[948]$_DFFE_PP__2795  (.L_HI(net2795));
 sg13g2_tiehi \logix.ram_r[949]$_DFFE_PP__2796  (.L_HI(net2796));
 sg13g2_tiehi \logix.ram_r[94]$_DFFE_PP__2797  (.L_HI(net2797));
 sg13g2_tiehi \logix.ram_r[950]$_DFFE_PP__2798  (.L_HI(net2798));
 sg13g2_tiehi \logix.ram_r[951]$_DFFE_PP__2799  (.L_HI(net2799));
 sg13g2_tiehi \logix.ram_r[952]$_DFFE_PP__2800  (.L_HI(net2800));
 sg13g2_tiehi \logix.ram_r[953]$_DFFE_PP__2801  (.L_HI(net2801));
 sg13g2_tiehi \logix.ram_r[954]$_DFFE_PP__2802  (.L_HI(net2802));
 sg13g2_tiehi \logix.ram_r[955]$_DFFE_PP__2803  (.L_HI(net2803));
 sg13g2_tiehi \logix.ram_r[956]$_DFFE_PP__2804  (.L_HI(net2804));
 sg13g2_tiehi \logix.ram_r[957]$_DFFE_PP__2805  (.L_HI(net2805));
 sg13g2_tiehi \logix.ram_r[958]$_DFFE_PP__2806  (.L_HI(net2806));
 sg13g2_tiehi \logix.ram_r[959]$_DFFE_PP__2807  (.L_HI(net2807));
 sg13g2_tiehi \logix.ram_r[95]$_DFFE_PP__2808  (.L_HI(net2808));
 sg13g2_tiehi \logix.ram_r[960]$_DFFE_PP__2809  (.L_HI(net2809));
 sg13g2_tiehi \logix.ram_r[961]$_DFFE_PP__2810  (.L_HI(net2810));
 sg13g2_tiehi \logix.ram_r[962]$_DFFE_PP__2811  (.L_HI(net2811));
 sg13g2_tiehi \logix.ram_r[963]$_DFFE_PP__2812  (.L_HI(net2812));
 sg13g2_tiehi \logix.ram_r[964]$_DFFE_PP__2813  (.L_HI(net2813));
 sg13g2_tiehi \logix.ram_r[965]$_DFFE_PP__2814  (.L_HI(net2814));
 sg13g2_tiehi \logix.ram_r[966]$_DFFE_PP__2815  (.L_HI(net2815));
 sg13g2_tiehi \logix.ram_r[967]$_DFFE_PP__2816  (.L_HI(net2816));
 sg13g2_tiehi \logix.ram_r[968]$_DFFE_PP__2817  (.L_HI(net2817));
 sg13g2_tiehi \logix.ram_r[969]$_DFFE_PP__2818  (.L_HI(net2818));
 sg13g2_tiehi \logix.ram_r[96]$_DFFE_PP__2819  (.L_HI(net2819));
 sg13g2_tiehi \logix.ram_r[970]$_DFFE_PP__2820  (.L_HI(net2820));
 sg13g2_tiehi \logix.ram_r[971]$_DFFE_PP__2821  (.L_HI(net2821));
 sg13g2_tiehi \logix.ram_r[972]$_DFFE_PP__2822  (.L_HI(net2822));
 sg13g2_tiehi \logix.ram_r[973]$_DFFE_PP__2823  (.L_HI(net2823));
 sg13g2_tiehi \logix.ram_r[974]$_DFFE_PP__2824  (.L_HI(net2824));
 sg13g2_tiehi \logix.ram_r[975]$_DFFE_PP__2825  (.L_HI(net2825));
 sg13g2_tiehi \logix.ram_r[976]$_DFFE_PP__2826  (.L_HI(net2826));
 sg13g2_tiehi \logix.ram_r[977]$_DFFE_PP__2827  (.L_HI(net2827));
 sg13g2_tiehi \logix.ram_r[978]$_DFFE_PP__2828  (.L_HI(net2828));
 sg13g2_tiehi \logix.ram_r[979]$_DFFE_PP__2829  (.L_HI(net2829));
 sg13g2_tiehi \logix.ram_r[97]$_DFFE_PP__2830  (.L_HI(net2830));
 sg13g2_tiehi \logix.ram_r[980]$_DFFE_PP__2831  (.L_HI(net2831));
 sg13g2_tiehi \logix.ram_r[981]$_DFFE_PP__2832  (.L_HI(net2832));
 sg13g2_tiehi \logix.ram_r[982]$_DFFE_PP__2833  (.L_HI(net2833));
 sg13g2_tiehi \logix.ram_r[983]$_DFFE_PP__2834  (.L_HI(net2834));
 sg13g2_tiehi \logix.ram_r[984]$_DFFE_PP__2835  (.L_HI(net2835));
 sg13g2_tiehi \logix.ram_r[985]$_DFFE_PP__2836  (.L_HI(net2836));
 sg13g2_tiehi \logix.ram_r[986]$_DFFE_PP__2837  (.L_HI(net2837));
 sg13g2_tiehi \logix.ram_r[987]$_DFFE_PP__2838  (.L_HI(net2838));
 sg13g2_tiehi \logix.ram_r[988]$_DFFE_PP__2839  (.L_HI(net2839));
 sg13g2_tiehi \logix.ram_r[989]$_DFFE_PP__2840  (.L_HI(net2840));
 sg13g2_tiehi \logix.ram_r[98]$_DFFE_PP__2841  (.L_HI(net2841));
 sg13g2_tiehi \logix.ram_r[990]$_DFFE_PP__2842  (.L_HI(net2842));
 sg13g2_tiehi \logix.ram_r[991]$_DFFE_PP__2843  (.L_HI(net2843));
 sg13g2_tiehi \logix.ram_r[992]$_DFFE_PP__2844  (.L_HI(net2844));
 sg13g2_tiehi \logix.ram_r[993]$_DFFE_PP__2845  (.L_HI(net2845));
 sg13g2_tiehi \logix.ram_r[994]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \logix.ram_r[995]$_DFFE_PP__2847  (.L_HI(net2847));
 sg13g2_tiehi \logix.ram_r[996]$_DFFE_PP__2848  (.L_HI(net2848));
 sg13g2_tiehi \logix.ram_r[997]$_DFFE_PP__2849  (.L_HI(net2849));
 sg13g2_tiehi \logix.ram_r[998]$_DFFE_PP__2850  (.L_HI(net2850));
 sg13g2_tiehi \logix.ram_r[999]$_DFFE_PP__2851  (.L_HI(net2851));
 sg13g2_tiehi \logix.ram_r[99]$_DFFE_PP__2852  (.L_HI(net2852));
 sg13g2_tiehi \logix.ram_r[9]$_DFFE_PP__2853  (.L_HI(net2853));
 sg13g2_buf_4 clkbuf_1_0__f_clk (.X(clknet_1_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_1_1__f_clk (.X(clknet_1_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_2064_));
 sg13g2_antennanp ANTENNA_2 (.A(_2064_));
 sg13g2_antennanp ANTENNA_3 (.A(_2064_));
 sg13g2_antennanp ANTENNA_4 (.A(_2064_));
 sg13g2_antennanp ANTENNA_5 (.A(_2064_));
 sg13g2_antennanp ANTENNA_6 (.A(_2064_));
 sg13g2_antennanp ANTENNA_7 (.A(_2064_));
 sg13g2_antennanp ANTENNA_8 (.A(_2064_));
 sg13g2_antennanp ANTENNA_9 (.A(_2201_));
 sg13g2_antennanp ANTENNA_10 (.A(_2201_));
 sg13g2_antennanp ANTENNA_11 (.A(_2201_));
 sg13g2_antennanp ANTENNA_12 (.A(_2201_));
 sg13g2_antennanp ANTENNA_13 (.A(_2201_));
 sg13g2_antennanp ANTENNA_14 (.A(_2201_));
 sg13g2_antennanp ANTENNA_15 (.A(_2201_));
 sg13g2_antennanp ANTENNA_16 (.A(_2344_));
 sg13g2_antennanp ANTENNA_17 (.A(_2344_));
 sg13g2_antennanp ANTENNA_18 (.A(_2344_));
 sg13g2_antennanp ANTENNA_19 (.A(_2344_));
 sg13g2_antennanp ANTENNA_20 (.A(_2344_));
 sg13g2_antennanp ANTENNA_21 (.A(_2344_));
 sg13g2_antennanp ANTENNA_22 (.A(_2344_));
 sg13g2_antennanp ANTENNA_23 (.A(_2353_));
 sg13g2_antennanp ANTENNA_24 (.A(_2353_));
 sg13g2_antennanp ANTENNA_25 (.A(_2353_));
 sg13g2_antennanp ANTENNA_26 (.A(_2353_));
 sg13g2_antennanp ANTENNA_27 (.A(_2378_));
 sg13g2_antennanp ANTENNA_28 (.A(_2378_));
 sg13g2_antennanp ANTENNA_29 (.A(_2378_));
 sg13g2_antennanp ANTENNA_30 (.A(_2378_));
 sg13g2_antennanp ANTENNA_31 (.A(_2378_));
 sg13g2_antennanp ANTENNA_32 (.A(_2378_));
 sg13g2_antennanp ANTENNA_33 (.A(_2378_));
 sg13g2_antennanp ANTENNA_34 (.A(_2378_));
 sg13g2_antennanp ANTENNA_35 (.A(_2378_));
 sg13g2_antennanp ANTENNA_36 (.A(_2378_));
 sg13g2_antennanp ANTENNA_37 (.A(_2401_));
 sg13g2_antennanp ANTENNA_38 (.A(_2401_));
 sg13g2_antennanp ANTENNA_39 (.A(_2411_));
 sg13g2_antennanp ANTENNA_40 (.A(_2411_));
 sg13g2_antennanp ANTENNA_41 (.A(_2411_));
 sg13g2_antennanp ANTENNA_42 (.A(_2411_));
 sg13g2_antennanp ANTENNA_43 (.A(_2411_));
 sg13g2_antennanp ANTENNA_44 (.A(_2411_));
 sg13g2_antennanp ANTENNA_45 (.A(_2411_));
 sg13g2_antennanp ANTENNA_46 (.A(_2443_));
 sg13g2_antennanp ANTENNA_47 (.A(_2443_));
 sg13g2_antennanp ANTENNA_48 (.A(_2458_));
 sg13g2_antennanp ANTENNA_49 (.A(_2458_));
 sg13g2_antennanp ANTENNA_50 (.A(_2458_));
 sg13g2_antennanp ANTENNA_51 (.A(_2458_));
 sg13g2_antennanp ANTENNA_52 (.A(_2458_));
 sg13g2_antennanp ANTENNA_53 (.A(_2458_));
 sg13g2_antennanp ANTENNA_54 (.A(_2458_));
 sg13g2_antennanp ANTENNA_55 (.A(_2458_));
 sg13g2_antennanp ANTENNA_56 (.A(_2473_));
 sg13g2_antennanp ANTENNA_57 (.A(_2473_));
 sg13g2_antennanp ANTENNA_58 (.A(_2473_));
 sg13g2_antennanp ANTENNA_59 (.A(_2488_));
 sg13g2_antennanp ANTENNA_60 (.A(_2488_));
 sg13g2_antennanp ANTENNA_61 (.A(_2488_));
 sg13g2_antennanp ANTENNA_62 (.A(_2494_));
 sg13g2_antennanp ANTENNA_63 (.A(_2494_));
 sg13g2_antennanp ANTENNA_64 (.A(_2494_));
 sg13g2_antennanp ANTENNA_65 (.A(_2494_));
 sg13g2_antennanp ANTENNA_66 (.A(_2550_));
 sg13g2_antennanp ANTENNA_67 (.A(_2550_));
 sg13g2_antennanp ANTENNA_68 (.A(_2588_));
 sg13g2_antennanp ANTENNA_69 (.A(_2588_));
 sg13g2_antennanp ANTENNA_70 (.A(_2588_));
 sg13g2_antennanp ANTENNA_71 (.A(_2588_));
 sg13g2_antennanp ANTENNA_72 (.A(_2596_));
 sg13g2_antennanp ANTENNA_73 (.A(_2596_));
 sg13g2_antennanp ANTENNA_74 (.A(_2596_));
 sg13g2_antennanp ANTENNA_75 (.A(_2596_));
 sg13g2_antennanp ANTENNA_76 (.A(_2598_));
 sg13g2_antennanp ANTENNA_77 (.A(_2612_));
 sg13g2_antennanp ANTENNA_78 (.A(_2612_));
 sg13g2_antennanp ANTENNA_79 (.A(_2612_));
 sg13g2_antennanp ANTENNA_80 (.A(_2624_));
 sg13g2_antennanp ANTENNA_81 (.A(_2624_));
 sg13g2_antennanp ANTENNA_82 (.A(_2624_));
 sg13g2_antennanp ANTENNA_83 (.A(_2711_));
 sg13g2_antennanp ANTENNA_84 (.A(_2762_));
 sg13g2_antennanp ANTENNA_85 (.A(_2878_));
 sg13g2_antennanp ANTENNA_86 (.A(_2906_));
 sg13g2_antennanp ANTENNA_87 (.A(_2941_));
 sg13g2_antennanp ANTENNA_88 (.A(_2941_));
 sg13g2_antennanp ANTENNA_89 (.A(_2941_));
 sg13g2_antennanp ANTENNA_90 (.A(_2955_));
 sg13g2_antennanp ANTENNA_91 (.A(_2955_));
 sg13g2_antennanp ANTENNA_92 (.A(_2955_));
 sg13g2_antennanp ANTENNA_93 (.A(_2977_));
 sg13g2_antennanp ANTENNA_94 (.A(_2977_));
 sg13g2_antennanp ANTENNA_95 (.A(_2977_));
 sg13g2_antennanp ANTENNA_96 (.A(_2978_));
 sg13g2_antennanp ANTENNA_97 (.A(_2978_));
 sg13g2_antennanp ANTENNA_98 (.A(_2978_));
 sg13g2_antennanp ANTENNA_99 (.A(_2990_));
 sg13g2_antennanp ANTENNA_100 (.A(_2990_));
 sg13g2_antennanp ANTENNA_101 (.A(_2990_));
 sg13g2_antennanp ANTENNA_102 (.A(_2990_));
 sg13g2_antennanp ANTENNA_103 (.A(_3003_));
 sg13g2_antennanp ANTENNA_104 (.A(_3021_));
 sg13g2_antennanp ANTENNA_105 (.A(_3046_));
 sg13g2_antennanp ANTENNA_106 (.A(_3046_));
 sg13g2_antennanp ANTENNA_107 (.A(_3053_));
 sg13g2_antennanp ANTENNA_108 (.A(_3053_));
 sg13g2_antennanp ANTENNA_109 (.A(_3053_));
 sg13g2_antennanp ANTENNA_110 (.A(_3079_));
 sg13g2_antennanp ANTENNA_111 (.A(_3098_));
 sg13g2_antennanp ANTENNA_112 (.A(_3130_));
 sg13g2_antennanp ANTENNA_113 (.A(_3130_));
 sg13g2_antennanp ANTENNA_114 (.A(_3141_));
 sg13g2_antennanp ANTENNA_115 (.A(_3213_));
 sg13g2_antennanp ANTENNA_116 (.A(_3213_));
 sg13g2_antennanp ANTENNA_117 (.A(_3221_));
 sg13g2_antennanp ANTENNA_118 (.A(_3221_));
 sg13g2_antennanp ANTENNA_119 (.A(_3228_));
 sg13g2_antennanp ANTENNA_120 (.A(_3241_));
 sg13g2_antennanp ANTENNA_121 (.A(_3259_));
 sg13g2_antennanp ANTENNA_122 (.A(_3294_));
 sg13g2_antennanp ANTENNA_123 (.A(_3299_));
 sg13g2_antennanp ANTENNA_124 (.A(_3333_));
 sg13g2_antennanp ANTENNA_125 (.A(_3333_));
 sg13g2_antennanp ANTENNA_126 (.A(_3348_));
 sg13g2_antennanp ANTENNA_127 (.A(_3372_));
 sg13g2_antennanp ANTENNA_128 (.A(_3472_));
 sg13g2_antennanp ANTENNA_129 (.A(_3522_));
 sg13g2_antennanp ANTENNA_130 (.A(_3614_));
 sg13g2_antennanp ANTENNA_131 (.A(_3640_));
 sg13g2_antennanp ANTENNA_132 (.A(_3751_));
 sg13g2_antennanp ANTENNA_133 (.A(_3751_));
 sg13g2_antennanp ANTENNA_134 (.A(_3835_));
 sg13g2_antennanp ANTENNA_135 (.A(_3858_));
 sg13g2_antennanp ANTENNA_136 (.A(_3871_));
 sg13g2_antennanp ANTENNA_137 (.A(_3891_));
 sg13g2_antennanp ANTENNA_138 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_139 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_140 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_141 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_142 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_143 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_144 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_145 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_146 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_147 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_148 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_149 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_150 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_151 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_152 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_153 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_154 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_155 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_156 (.A(net10));
 sg13g2_antennanp ANTENNA_157 (.A(net14));
 sg13g2_antennanp ANTENNA_158 (.A(net14));
 sg13g2_antennanp ANTENNA_159 (.A(net14));
 sg13g2_antennanp ANTENNA_160 (.A(net14));
 sg13g2_antennanp ANTENNA_161 (.A(net14));
 sg13g2_antennanp ANTENNA_162 (.A(net14));
 sg13g2_antennanp ANTENNA_163 (.A(net14));
 sg13g2_antennanp ANTENNA_164 (.A(net14));
 sg13g2_antennanp ANTENNA_165 (.A(net15));
 sg13g2_antennanp ANTENNA_166 (.A(net15));
 sg13g2_antennanp ANTENNA_167 (.A(net17));
 sg13g2_antennanp ANTENNA_168 (.A(net17));
 sg13g2_antennanp ANTENNA_169 (.A(net17));
 sg13g2_antennanp ANTENNA_170 (.A(net18));
 sg13g2_antennanp ANTENNA_171 (.A(net18));
 sg13g2_antennanp ANTENNA_172 (.A(net18));
 sg13g2_antennanp ANTENNA_173 (.A(net19));
 sg13g2_antennanp ANTENNA_174 (.A(net19));
 sg13g2_antennanp ANTENNA_175 (.A(net19));
 sg13g2_antennanp ANTENNA_176 (.A(net20));
 sg13g2_antennanp ANTENNA_177 (.A(net20));
 sg13g2_antennanp ANTENNA_178 (.A(net20));
 sg13g2_antennanp ANTENNA_179 (.A(net20));
 sg13g2_antennanp ANTENNA_180 (.A(net21));
 sg13g2_antennanp ANTENNA_181 (.A(net21));
 sg13g2_antennanp ANTENNA_182 (.A(net21));
 sg13g2_antennanp ANTENNA_183 (.A(net21));
 sg13g2_antennanp ANTENNA_184 (.A(net21));
 sg13g2_antennanp ANTENNA_185 (.A(net21));
 sg13g2_antennanp ANTENNA_186 (.A(net21));
 sg13g2_antennanp ANTENNA_187 (.A(net21));
 sg13g2_antennanp ANTENNA_188 (.A(net23));
 sg13g2_antennanp ANTENNA_189 (.A(net23));
 sg13g2_antennanp ANTENNA_190 (.A(net23));
 sg13g2_antennanp ANTENNA_191 (.A(net23));
 sg13g2_antennanp ANTENNA_192 (.A(net23));
 sg13g2_antennanp ANTENNA_193 (.A(net23));
 sg13g2_antennanp ANTENNA_194 (.A(net23));
 sg13g2_antennanp ANTENNA_195 (.A(net23));
 sg13g2_antennanp ANTENNA_196 (.A(net27));
 sg13g2_antennanp ANTENNA_197 (.A(net27));
 sg13g2_antennanp ANTENNA_198 (.A(net27));
 sg13g2_antennanp ANTENNA_199 (.A(net27));
 sg13g2_antennanp ANTENNA_200 (.A(net27));
 sg13g2_antennanp ANTENNA_201 (.A(net27));
 sg13g2_antennanp ANTENNA_202 (.A(net27));
 sg13g2_antennanp ANTENNA_203 (.A(net27));
 sg13g2_antennanp ANTENNA_204 (.A(net27));
 sg13g2_antennanp ANTENNA_205 (.A(net45));
 sg13g2_antennanp ANTENNA_206 (.A(net45));
 sg13g2_antennanp ANTENNA_207 (.A(net45));
 sg13g2_antennanp ANTENNA_208 (.A(net45));
 sg13g2_antennanp ANTENNA_209 (.A(net45));
 sg13g2_antennanp ANTENNA_210 (.A(net45));
 sg13g2_antennanp ANTENNA_211 (.A(net45));
 sg13g2_antennanp ANTENNA_212 (.A(net45));
 sg13g2_antennanp ANTENNA_213 (.A(net61));
 sg13g2_antennanp ANTENNA_214 (.A(net61));
 sg13g2_antennanp ANTENNA_215 (.A(net61));
 sg13g2_antennanp ANTENNA_216 (.A(net61));
 sg13g2_antennanp ANTENNA_217 (.A(net61));
 sg13g2_antennanp ANTENNA_218 (.A(net61));
 sg13g2_antennanp ANTENNA_219 (.A(net61));
 sg13g2_antennanp ANTENNA_220 (.A(net61));
 sg13g2_antennanp ANTENNA_221 (.A(net73));
 sg13g2_antennanp ANTENNA_222 (.A(net73));
 sg13g2_antennanp ANTENNA_223 (.A(net73));
 sg13g2_antennanp ANTENNA_224 (.A(net73));
 sg13g2_antennanp ANTENNA_225 (.A(net73));
 sg13g2_antennanp ANTENNA_226 (.A(net73));
 sg13g2_antennanp ANTENNA_227 (.A(net73));
 sg13g2_antennanp ANTENNA_228 (.A(net73));
 sg13g2_antennanp ANTENNA_229 (.A(net73));
 sg13g2_antennanp ANTENNA_230 (.A(net74));
 sg13g2_antennanp ANTENNA_231 (.A(net74));
 sg13g2_antennanp ANTENNA_232 (.A(net74));
 sg13g2_antennanp ANTENNA_233 (.A(net74));
 sg13g2_antennanp ANTENNA_234 (.A(net74));
 sg13g2_antennanp ANTENNA_235 (.A(net74));
 sg13g2_antennanp ANTENNA_236 (.A(net74));
 sg13g2_antennanp ANTENNA_237 (.A(net74));
 sg13g2_antennanp ANTENNA_238 (.A(net74));
 sg13g2_antennanp ANTENNA_239 (.A(net79));
 sg13g2_antennanp ANTENNA_240 (.A(net79));
 sg13g2_antennanp ANTENNA_241 (.A(net79));
 sg13g2_antennanp ANTENNA_242 (.A(net79));
 sg13g2_antennanp ANTENNA_243 (.A(net79));
 sg13g2_antennanp ANTENNA_244 (.A(net79));
 sg13g2_antennanp ANTENNA_245 (.A(net79));
 sg13g2_antennanp ANTENNA_246 (.A(net79));
 sg13g2_antennanp ANTENNA_247 (.A(net79));
 sg13g2_antennanp ANTENNA_248 (.A(net79));
 sg13g2_antennanp ANTENNA_249 (.A(net79));
 sg13g2_antennanp ANTENNA_250 (.A(net79));
 sg13g2_antennanp ANTENNA_251 (.A(net79));
 sg13g2_antennanp ANTENNA_252 (.A(net84));
 sg13g2_antennanp ANTENNA_253 (.A(net84));
 sg13g2_antennanp ANTENNA_254 (.A(net84));
 sg13g2_antennanp ANTENNA_255 (.A(net84));
 sg13g2_antennanp ANTENNA_256 (.A(net84));
 sg13g2_antennanp ANTENNA_257 (.A(net84));
 sg13g2_antennanp ANTENNA_258 (.A(net84));
 sg13g2_antennanp ANTENNA_259 (.A(net84));
 sg13g2_antennanp ANTENNA_260 (.A(net84));
 sg13g2_antennanp ANTENNA_261 (.A(net85));
 sg13g2_antennanp ANTENNA_262 (.A(net85));
 sg13g2_antennanp ANTENNA_263 (.A(net85));
 sg13g2_antennanp ANTENNA_264 (.A(net85));
 sg13g2_antennanp ANTENNA_265 (.A(net85));
 sg13g2_antennanp ANTENNA_266 (.A(net85));
 sg13g2_antennanp ANTENNA_267 (.A(net85));
 sg13g2_antennanp ANTENNA_268 (.A(net85));
 sg13g2_antennanp ANTENNA_269 (.A(net85));
 sg13g2_antennanp ANTENNA_270 (.A(net90));
 sg13g2_antennanp ANTENNA_271 (.A(net90));
 sg13g2_antennanp ANTENNA_272 (.A(net90));
 sg13g2_antennanp ANTENNA_273 (.A(net90));
 sg13g2_antennanp ANTENNA_274 (.A(net90));
 sg13g2_antennanp ANTENNA_275 (.A(net90));
 sg13g2_antennanp ANTENNA_276 (.A(net90));
 sg13g2_antennanp ANTENNA_277 (.A(net90));
 sg13g2_antennanp ANTENNA_278 (.A(net90));
 sg13g2_antennanp ANTENNA_279 (.A(net92));
 sg13g2_antennanp ANTENNA_280 (.A(net92));
 sg13g2_antennanp ANTENNA_281 (.A(net92));
 sg13g2_antennanp ANTENNA_282 (.A(net92));
 sg13g2_antennanp ANTENNA_283 (.A(net92));
 sg13g2_antennanp ANTENNA_284 (.A(net92));
 sg13g2_antennanp ANTENNA_285 (.A(net92));
 sg13g2_antennanp ANTENNA_286 (.A(net92));
 sg13g2_antennanp ANTENNA_287 (.A(net92));
 sg13g2_antennanp ANTENNA_288 (.A(net95));
 sg13g2_antennanp ANTENNA_289 (.A(net95));
 sg13g2_antennanp ANTENNA_290 (.A(net95));
 sg13g2_antennanp ANTENNA_291 (.A(net95));
 sg13g2_antennanp ANTENNA_292 (.A(net95));
 sg13g2_antennanp ANTENNA_293 (.A(net95));
 sg13g2_antennanp ANTENNA_294 (.A(net95));
 sg13g2_antennanp ANTENNA_295 (.A(net95));
 sg13g2_antennanp ANTENNA_296 (.A(net95));
 sg13g2_antennanp ANTENNA_297 (.A(net140));
 sg13g2_antennanp ANTENNA_298 (.A(net140));
 sg13g2_antennanp ANTENNA_299 (.A(net140));
 sg13g2_antennanp ANTENNA_300 (.A(net140));
 sg13g2_antennanp ANTENNA_301 (.A(net140));
 sg13g2_antennanp ANTENNA_302 (.A(net140));
 sg13g2_antennanp ANTENNA_303 (.A(net140));
 sg13g2_antennanp ANTENNA_304 (.A(net140));
 sg13g2_antennanp ANTENNA_305 (.A(net140));
 sg13g2_antennanp ANTENNA_306 (.A(net153));
 sg13g2_antennanp ANTENNA_307 (.A(net153));
 sg13g2_antennanp ANTENNA_308 (.A(net153));
 sg13g2_antennanp ANTENNA_309 (.A(net153));
 sg13g2_antennanp ANTENNA_310 (.A(net153));
 sg13g2_antennanp ANTENNA_311 (.A(net153));
 sg13g2_antennanp ANTENNA_312 (.A(net153));
 sg13g2_antennanp ANTENNA_313 (.A(net153));
 sg13g2_antennanp ANTENNA_314 (.A(net153));
 sg13g2_antennanp ANTENNA_315 (.A(net162));
 sg13g2_antennanp ANTENNA_316 (.A(net162));
 sg13g2_antennanp ANTENNA_317 (.A(net162));
 sg13g2_antennanp ANTENNA_318 (.A(net162));
 sg13g2_antennanp ANTENNA_319 (.A(net162));
 sg13g2_antennanp ANTENNA_320 (.A(net162));
 sg13g2_antennanp ANTENNA_321 (.A(net162));
 sg13g2_antennanp ANTENNA_322 (.A(net162));
 sg13g2_antennanp ANTENNA_323 (.A(net162));
 sg13g2_antennanp ANTENNA_324 (.A(net162));
 sg13g2_antennanp ANTENNA_325 (.A(net162));
 sg13g2_antennanp ANTENNA_326 (.A(net162));
 sg13g2_antennanp ANTENNA_327 (.A(net163));
 sg13g2_antennanp ANTENNA_328 (.A(net163));
 sg13g2_antennanp ANTENNA_329 (.A(net163));
 sg13g2_antennanp ANTENNA_330 (.A(net163));
 sg13g2_antennanp ANTENNA_331 (.A(net163));
 sg13g2_antennanp ANTENNA_332 (.A(net163));
 sg13g2_antennanp ANTENNA_333 (.A(net163));
 sg13g2_antennanp ANTENNA_334 (.A(net163));
 sg13g2_antennanp ANTENNA_335 (.A(net163));
 sg13g2_antennanp ANTENNA_336 (.A(net174));
 sg13g2_antennanp ANTENNA_337 (.A(net174));
 sg13g2_antennanp ANTENNA_338 (.A(net174));
 sg13g2_antennanp ANTENNA_339 (.A(net174));
 sg13g2_antennanp ANTENNA_340 (.A(net174));
 sg13g2_antennanp ANTENNA_341 (.A(net174));
 sg13g2_antennanp ANTENNA_342 (.A(net174));
 sg13g2_antennanp ANTENNA_343 (.A(net174));
 sg13g2_antennanp ANTENNA_344 (.A(net174));
 sg13g2_antennanp ANTENNA_345 (.A(net174));
 sg13g2_antennanp ANTENNA_346 (.A(net174));
 sg13g2_antennanp ANTENNA_347 (.A(net174));
 sg13g2_antennanp ANTENNA_348 (.A(net174));
 sg13g2_antennanp ANTENNA_349 (.A(net181));
 sg13g2_antennanp ANTENNA_350 (.A(net181));
 sg13g2_antennanp ANTENNA_351 (.A(net181));
 sg13g2_antennanp ANTENNA_352 (.A(net181));
 sg13g2_antennanp ANTENNA_353 (.A(net181));
 sg13g2_antennanp ANTENNA_354 (.A(net181));
 sg13g2_antennanp ANTENNA_355 (.A(net181));
 sg13g2_antennanp ANTENNA_356 (.A(net181));
 sg13g2_antennanp ANTENNA_357 (.A(net184));
 sg13g2_antennanp ANTENNA_358 (.A(net184));
 sg13g2_antennanp ANTENNA_359 (.A(net184));
 sg13g2_antennanp ANTENNA_360 (.A(net184));
 sg13g2_antennanp ANTENNA_361 (.A(net184));
 sg13g2_antennanp ANTENNA_362 (.A(net184));
 sg13g2_antennanp ANTENNA_363 (.A(net184));
 sg13g2_antennanp ANTENNA_364 (.A(net184));
 sg13g2_antennanp ANTENNA_365 (.A(net184));
 sg13g2_antennanp ANTENNA_366 (.A(net192));
 sg13g2_antennanp ANTENNA_367 (.A(net192));
 sg13g2_antennanp ANTENNA_368 (.A(net192));
 sg13g2_antennanp ANTENNA_369 (.A(net192));
 sg13g2_antennanp ANTENNA_370 (.A(net192));
 sg13g2_antennanp ANTENNA_371 (.A(net192));
 sg13g2_antennanp ANTENNA_372 (.A(net192));
 sg13g2_antennanp ANTENNA_373 (.A(net192));
 sg13g2_antennanp ANTENNA_374 (.A(net192));
 sg13g2_antennanp ANTENNA_375 (.A(net192));
 sg13g2_antennanp ANTENNA_376 (.A(net192));
 sg13g2_antennanp ANTENNA_377 (.A(net192));
 sg13g2_antennanp ANTENNA_378 (.A(net192));
 sg13g2_antennanp ANTENNA_379 (.A(net192));
 sg13g2_antennanp ANTENNA_380 (.A(net192));
 sg13g2_antennanp ANTENNA_381 (.A(net192));
 sg13g2_antennanp ANTENNA_382 (.A(net192));
 sg13g2_antennanp ANTENNA_383 (.A(net192));
 sg13g2_antennanp ANTENNA_384 (.A(net202));
 sg13g2_antennanp ANTENNA_385 (.A(net202));
 sg13g2_antennanp ANTENNA_386 (.A(net202));
 sg13g2_antennanp ANTENNA_387 (.A(net202));
 sg13g2_antennanp ANTENNA_388 (.A(net202));
 sg13g2_antennanp ANTENNA_389 (.A(net202));
 sg13g2_antennanp ANTENNA_390 (.A(net202));
 sg13g2_antennanp ANTENNA_391 (.A(net202));
 sg13g2_antennanp ANTENNA_392 (.A(net202));
 sg13g2_antennanp ANTENNA_393 (.A(net205));
 sg13g2_antennanp ANTENNA_394 (.A(net205));
 sg13g2_antennanp ANTENNA_395 (.A(net205));
 sg13g2_antennanp ANTENNA_396 (.A(net205));
 sg13g2_antennanp ANTENNA_397 (.A(net205));
 sg13g2_antennanp ANTENNA_398 (.A(net205));
 sg13g2_antennanp ANTENNA_399 (.A(net205));
 sg13g2_antennanp ANTENNA_400 (.A(net205));
 sg13g2_antennanp ANTENNA_401 (.A(net205));
 sg13g2_antennanp ANTENNA_402 (.A(net206));
 sg13g2_antennanp ANTENNA_403 (.A(net206));
 sg13g2_antennanp ANTENNA_404 (.A(net206));
 sg13g2_antennanp ANTENNA_405 (.A(net206));
 sg13g2_antennanp ANTENNA_406 (.A(net206));
 sg13g2_antennanp ANTENNA_407 (.A(net206));
 sg13g2_antennanp ANTENNA_408 (.A(net206));
 sg13g2_antennanp ANTENNA_409 (.A(net206));
 sg13g2_antennanp ANTENNA_410 (.A(net206));
 sg13g2_antennanp ANTENNA_411 (.A(net207));
 sg13g2_antennanp ANTENNA_412 (.A(net207));
 sg13g2_antennanp ANTENNA_413 (.A(net207));
 sg13g2_antennanp ANTENNA_414 (.A(net207));
 sg13g2_antennanp ANTENNA_415 (.A(net207));
 sg13g2_antennanp ANTENNA_416 (.A(net207));
 sg13g2_antennanp ANTENNA_417 (.A(net207));
 sg13g2_antennanp ANTENNA_418 (.A(net207));
 sg13g2_antennanp ANTENNA_419 (.A(net207));
 sg13g2_antennanp ANTENNA_420 (.A(_2064_));
 sg13g2_antennanp ANTENNA_421 (.A(_2064_));
 sg13g2_antennanp ANTENNA_422 (.A(_2064_));
 sg13g2_antennanp ANTENNA_423 (.A(_2064_));
 sg13g2_antennanp ANTENNA_424 (.A(_2064_));
 sg13g2_antennanp ANTENNA_425 (.A(_2064_));
 sg13g2_antennanp ANTENNA_426 (.A(_2064_));
 sg13g2_antennanp ANTENNA_427 (.A(_2064_));
 sg13g2_antennanp ANTENNA_428 (.A(_2201_));
 sg13g2_antennanp ANTENNA_429 (.A(_2201_));
 sg13g2_antennanp ANTENNA_430 (.A(_2201_));
 sg13g2_antennanp ANTENNA_431 (.A(_2201_));
 sg13g2_antennanp ANTENNA_432 (.A(_2201_));
 sg13g2_antennanp ANTENNA_433 (.A(_2201_));
 sg13g2_antennanp ANTENNA_434 (.A(_2201_));
 sg13g2_antennanp ANTENNA_435 (.A(_2201_));
 sg13g2_antennanp ANTENNA_436 (.A(_2344_));
 sg13g2_antennanp ANTENNA_437 (.A(_2344_));
 sg13g2_antennanp ANTENNA_438 (.A(_2344_));
 sg13g2_antennanp ANTENNA_439 (.A(_2344_));
 sg13g2_antennanp ANTENNA_440 (.A(_2344_));
 sg13g2_antennanp ANTENNA_441 (.A(_2344_));
 sg13g2_antennanp ANTENNA_442 (.A(_2344_));
 sg13g2_antennanp ANTENNA_443 (.A(_2353_));
 sg13g2_antennanp ANTENNA_444 (.A(_2353_));
 sg13g2_antennanp ANTENNA_445 (.A(_2353_));
 sg13g2_antennanp ANTENNA_446 (.A(_2353_));
 sg13g2_antennanp ANTENNA_447 (.A(_2378_));
 sg13g2_antennanp ANTENNA_448 (.A(_2378_));
 sg13g2_antennanp ANTENNA_449 (.A(_2378_));
 sg13g2_antennanp ANTENNA_450 (.A(_2378_));
 sg13g2_antennanp ANTENNA_451 (.A(_2378_));
 sg13g2_antennanp ANTENNA_452 (.A(_2378_));
 sg13g2_antennanp ANTENNA_453 (.A(_2378_));
 sg13g2_antennanp ANTENNA_454 (.A(_2378_));
 sg13g2_antennanp ANTENNA_455 (.A(_2378_));
 sg13g2_antennanp ANTENNA_456 (.A(_2378_));
 sg13g2_antennanp ANTENNA_457 (.A(_2401_));
 sg13g2_antennanp ANTENNA_458 (.A(_2411_));
 sg13g2_antennanp ANTENNA_459 (.A(_2411_));
 sg13g2_antennanp ANTENNA_460 (.A(_2411_));
 sg13g2_antennanp ANTENNA_461 (.A(_2411_));
 sg13g2_antennanp ANTENNA_462 (.A(_2411_));
 sg13g2_antennanp ANTENNA_463 (.A(_2411_));
 sg13g2_antennanp ANTENNA_464 (.A(_2411_));
 sg13g2_antennanp ANTENNA_465 (.A(_2433_));
 sg13g2_antennanp ANTENNA_466 (.A(_2433_));
 sg13g2_antennanp ANTENNA_467 (.A(_2433_));
 sg13g2_antennanp ANTENNA_468 (.A(_2433_));
 sg13g2_antennanp ANTENNA_469 (.A(_2433_));
 sg13g2_antennanp ANTENNA_470 (.A(_2433_));
 sg13g2_antennanp ANTENNA_471 (.A(_2433_));
 sg13g2_antennanp ANTENNA_472 (.A(_2433_));
 sg13g2_antennanp ANTENNA_473 (.A(_2433_));
 sg13g2_antennanp ANTENNA_474 (.A(_2433_));
 sg13g2_antennanp ANTENNA_475 (.A(_2433_));
 sg13g2_antennanp ANTENNA_476 (.A(_2433_));
 sg13g2_antennanp ANTENNA_477 (.A(_2443_));
 sg13g2_antennanp ANTENNA_478 (.A(_2443_));
 sg13g2_antennanp ANTENNA_479 (.A(_2461_));
 sg13g2_antennanp ANTENNA_480 (.A(_2461_));
 sg13g2_antennanp ANTENNA_481 (.A(_2461_));
 sg13g2_antennanp ANTENNA_482 (.A(_2473_));
 sg13g2_antennanp ANTENNA_483 (.A(_2473_));
 sg13g2_antennanp ANTENNA_484 (.A(_2473_));
 sg13g2_antennanp ANTENNA_485 (.A(_2488_));
 sg13g2_antennanp ANTENNA_486 (.A(_2488_));
 sg13g2_antennanp ANTENNA_487 (.A(_2488_));
 sg13g2_antennanp ANTENNA_488 (.A(_2488_));
 sg13g2_antennanp ANTENNA_489 (.A(_2488_));
 sg13g2_antennanp ANTENNA_490 (.A(_2488_));
 sg13g2_antennanp ANTENNA_491 (.A(_2568_));
 sg13g2_antennanp ANTENNA_492 (.A(_2568_));
 sg13g2_antennanp ANTENNA_493 (.A(_2568_));
 sg13g2_antennanp ANTENNA_494 (.A(_2588_));
 sg13g2_antennanp ANTENNA_495 (.A(_2588_));
 sg13g2_antennanp ANTENNA_496 (.A(_2588_));
 sg13g2_antennanp ANTENNA_497 (.A(_2596_));
 sg13g2_antennanp ANTENNA_498 (.A(_2596_));
 sg13g2_antennanp ANTENNA_499 (.A(_2596_));
 sg13g2_antennanp ANTENNA_500 (.A(_2596_));
 sg13g2_antennanp ANTENNA_501 (.A(_2598_));
 sg13g2_antennanp ANTENNA_502 (.A(_2612_));
 sg13g2_antennanp ANTENNA_503 (.A(_2612_));
 sg13g2_antennanp ANTENNA_504 (.A(_2612_));
 sg13g2_antennanp ANTENNA_505 (.A(_2711_));
 sg13g2_antennanp ANTENNA_506 (.A(_2762_));
 sg13g2_antennanp ANTENNA_507 (.A(_2762_));
 sg13g2_antennanp ANTENNA_508 (.A(_2870_));
 sg13g2_antennanp ANTENNA_509 (.A(_2878_));
 sg13g2_antennanp ANTENNA_510 (.A(_2955_));
 sg13g2_antennanp ANTENNA_511 (.A(_2955_));
 sg13g2_antennanp ANTENNA_512 (.A(_2955_));
 sg13g2_antennanp ANTENNA_513 (.A(_2977_));
 sg13g2_antennanp ANTENNA_514 (.A(_2977_));
 sg13g2_antennanp ANTENNA_515 (.A(_2977_));
 sg13g2_antennanp ANTENNA_516 (.A(_2978_));
 sg13g2_antennanp ANTENNA_517 (.A(_2978_));
 sg13g2_antennanp ANTENNA_518 (.A(_2978_));
 sg13g2_antennanp ANTENNA_519 (.A(_2978_));
 sg13g2_antennanp ANTENNA_520 (.A(_2990_));
 sg13g2_antennanp ANTENNA_521 (.A(_2990_));
 sg13g2_antennanp ANTENNA_522 (.A(_2990_));
 sg13g2_antennanp ANTENNA_523 (.A(_2990_));
 sg13g2_antennanp ANTENNA_524 (.A(_3003_));
 sg13g2_antennanp ANTENNA_525 (.A(_3021_));
 sg13g2_antennanp ANTENNA_526 (.A(_3046_));
 sg13g2_antennanp ANTENNA_527 (.A(_3046_));
 sg13g2_antennanp ANTENNA_528 (.A(_3056_));
 sg13g2_antennanp ANTENNA_529 (.A(_3056_));
 sg13g2_antennanp ANTENNA_530 (.A(_3056_));
 sg13g2_antennanp ANTENNA_531 (.A(_3056_));
 sg13g2_antennanp ANTENNA_532 (.A(_3079_));
 sg13g2_antennanp ANTENNA_533 (.A(_3098_));
 sg13g2_antennanp ANTENNA_534 (.A(_3098_));
 sg13g2_antennanp ANTENNA_535 (.A(_3130_));
 sg13g2_antennanp ANTENNA_536 (.A(_3221_));
 sg13g2_antennanp ANTENNA_537 (.A(_3221_));
 sg13g2_antennanp ANTENNA_538 (.A(_3228_));
 sg13g2_antennanp ANTENNA_539 (.A(_3241_));
 sg13g2_antennanp ANTENNA_540 (.A(_3259_));
 sg13g2_antennanp ANTENNA_541 (.A(_3294_));
 sg13g2_antennanp ANTENNA_542 (.A(_3299_));
 sg13g2_antennanp ANTENNA_543 (.A(_3333_));
 sg13g2_antennanp ANTENNA_544 (.A(_3348_));
 sg13g2_antennanp ANTENNA_545 (.A(_3372_));
 sg13g2_antennanp ANTENNA_546 (.A(_3472_));
 sg13g2_antennanp ANTENNA_547 (.A(_3522_));
 sg13g2_antennanp ANTENNA_548 (.A(_3614_));
 sg13g2_antennanp ANTENNA_549 (.A(_3640_));
 sg13g2_antennanp ANTENNA_550 (.A(_3835_));
 sg13g2_antennanp ANTENNA_551 (.A(_3835_));
 sg13g2_antennanp ANTENNA_552 (.A(_3858_));
 sg13g2_antennanp ANTENNA_553 (.A(_3871_));
 sg13g2_antennanp ANTENNA_554 (.A(_3891_));
 sg13g2_antennanp ANTENNA_555 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_556 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_557 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_558 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_559 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_560 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_561 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_562 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_563 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_564 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_565 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_566 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_567 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_568 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_569 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_570 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_571 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_572 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_573 (.A(net10));
 sg13g2_antennanp ANTENNA_574 (.A(net14));
 sg13g2_antennanp ANTENNA_575 (.A(net14));
 sg13g2_antennanp ANTENNA_576 (.A(net14));
 sg13g2_antennanp ANTENNA_577 (.A(net15));
 sg13g2_antennanp ANTENNA_578 (.A(net15));
 sg13g2_antennanp ANTENNA_579 (.A(net15));
 sg13g2_antennanp ANTENNA_580 (.A(net23));
 sg13g2_antennanp ANTENNA_581 (.A(net23));
 sg13g2_antennanp ANTENNA_582 (.A(net23));
 sg13g2_antennanp ANTENNA_583 (.A(net23));
 sg13g2_antennanp ANTENNA_584 (.A(net23));
 sg13g2_antennanp ANTENNA_585 (.A(net23));
 sg13g2_antennanp ANTENNA_586 (.A(net23));
 sg13g2_antennanp ANTENNA_587 (.A(net23));
 sg13g2_antennanp ANTENNA_588 (.A(net61));
 sg13g2_antennanp ANTENNA_589 (.A(net61));
 sg13g2_antennanp ANTENNA_590 (.A(net61));
 sg13g2_antennanp ANTENNA_591 (.A(net61));
 sg13g2_antennanp ANTENNA_592 (.A(net61));
 sg13g2_antennanp ANTENNA_593 (.A(net61));
 sg13g2_antennanp ANTENNA_594 (.A(net61));
 sg13g2_antennanp ANTENNA_595 (.A(net61));
 sg13g2_antennanp ANTENNA_596 (.A(net68));
 sg13g2_antennanp ANTENNA_597 (.A(net68));
 sg13g2_antennanp ANTENNA_598 (.A(net68));
 sg13g2_antennanp ANTENNA_599 (.A(net68));
 sg13g2_antennanp ANTENNA_600 (.A(net68));
 sg13g2_antennanp ANTENNA_601 (.A(net68));
 sg13g2_antennanp ANTENNA_602 (.A(net68));
 sg13g2_antennanp ANTENNA_603 (.A(net68));
 sg13g2_antennanp ANTENNA_604 (.A(net68));
 sg13g2_antennanp ANTENNA_605 (.A(net69));
 sg13g2_antennanp ANTENNA_606 (.A(net69));
 sg13g2_antennanp ANTENNA_607 (.A(net69));
 sg13g2_antennanp ANTENNA_608 (.A(net69));
 sg13g2_antennanp ANTENNA_609 (.A(net69));
 sg13g2_antennanp ANTENNA_610 (.A(net69));
 sg13g2_antennanp ANTENNA_611 (.A(net69));
 sg13g2_antennanp ANTENNA_612 (.A(net69));
 sg13g2_antennanp ANTENNA_613 (.A(net69));
 sg13g2_antennanp ANTENNA_614 (.A(net73));
 sg13g2_antennanp ANTENNA_615 (.A(net73));
 sg13g2_antennanp ANTENNA_616 (.A(net73));
 sg13g2_antennanp ANTENNA_617 (.A(net73));
 sg13g2_antennanp ANTENNA_618 (.A(net73));
 sg13g2_antennanp ANTENNA_619 (.A(net73));
 sg13g2_antennanp ANTENNA_620 (.A(net73));
 sg13g2_antennanp ANTENNA_621 (.A(net73));
 sg13g2_antennanp ANTENNA_622 (.A(net73));
 sg13g2_antennanp ANTENNA_623 (.A(net74));
 sg13g2_antennanp ANTENNA_624 (.A(net74));
 sg13g2_antennanp ANTENNA_625 (.A(net74));
 sg13g2_antennanp ANTENNA_626 (.A(net74));
 sg13g2_antennanp ANTENNA_627 (.A(net74));
 sg13g2_antennanp ANTENNA_628 (.A(net74));
 sg13g2_antennanp ANTENNA_629 (.A(net74));
 sg13g2_antennanp ANTENNA_630 (.A(net74));
 sg13g2_antennanp ANTENNA_631 (.A(net74));
 sg13g2_antennanp ANTENNA_632 (.A(net79));
 sg13g2_antennanp ANTENNA_633 (.A(net79));
 sg13g2_antennanp ANTENNA_634 (.A(net79));
 sg13g2_antennanp ANTENNA_635 (.A(net79));
 sg13g2_antennanp ANTENNA_636 (.A(net79));
 sg13g2_antennanp ANTENNA_637 (.A(net79));
 sg13g2_antennanp ANTENNA_638 (.A(net79));
 sg13g2_antennanp ANTENNA_639 (.A(net79));
 sg13g2_antennanp ANTENNA_640 (.A(net79));
 sg13g2_antennanp ANTENNA_641 (.A(net85));
 sg13g2_antennanp ANTENNA_642 (.A(net85));
 sg13g2_antennanp ANTENNA_643 (.A(net85));
 sg13g2_antennanp ANTENNA_644 (.A(net85));
 sg13g2_antennanp ANTENNA_645 (.A(net85));
 sg13g2_antennanp ANTENNA_646 (.A(net85));
 sg13g2_antennanp ANTENNA_647 (.A(net85));
 sg13g2_antennanp ANTENNA_648 (.A(net85));
 sg13g2_antennanp ANTENNA_649 (.A(net85));
 sg13g2_antennanp ANTENNA_650 (.A(net92));
 sg13g2_antennanp ANTENNA_651 (.A(net92));
 sg13g2_antennanp ANTENNA_652 (.A(net92));
 sg13g2_antennanp ANTENNA_653 (.A(net92));
 sg13g2_antennanp ANTENNA_654 (.A(net92));
 sg13g2_antennanp ANTENNA_655 (.A(net92));
 sg13g2_antennanp ANTENNA_656 (.A(net92));
 sg13g2_antennanp ANTENNA_657 (.A(net92));
 sg13g2_antennanp ANTENNA_658 (.A(net93));
 sg13g2_antennanp ANTENNA_659 (.A(net93));
 sg13g2_antennanp ANTENNA_660 (.A(net93));
 sg13g2_antennanp ANTENNA_661 (.A(net93));
 sg13g2_antennanp ANTENNA_662 (.A(net93));
 sg13g2_antennanp ANTENNA_663 (.A(net93));
 sg13g2_antennanp ANTENNA_664 (.A(net93));
 sg13g2_antennanp ANTENNA_665 (.A(net93));
 sg13g2_antennanp ANTENNA_666 (.A(net93));
 sg13g2_antennanp ANTENNA_667 (.A(net163));
 sg13g2_antennanp ANTENNA_668 (.A(net163));
 sg13g2_antennanp ANTENNA_669 (.A(net163));
 sg13g2_antennanp ANTENNA_670 (.A(net163));
 sg13g2_antennanp ANTENNA_671 (.A(net163));
 sg13g2_antennanp ANTENNA_672 (.A(net163));
 sg13g2_antennanp ANTENNA_673 (.A(net163));
 sg13g2_antennanp ANTENNA_674 (.A(net163));
 sg13g2_antennanp ANTENNA_675 (.A(net174));
 sg13g2_antennanp ANTENNA_676 (.A(net174));
 sg13g2_antennanp ANTENNA_677 (.A(net174));
 sg13g2_antennanp ANTENNA_678 (.A(net174));
 sg13g2_antennanp ANTENNA_679 (.A(net174));
 sg13g2_antennanp ANTENNA_680 (.A(net174));
 sg13g2_antennanp ANTENNA_681 (.A(net174));
 sg13g2_antennanp ANTENNA_682 (.A(net174));
 sg13g2_antennanp ANTENNA_683 (.A(net174));
 sg13g2_antennanp ANTENNA_684 (.A(net184));
 sg13g2_antennanp ANTENNA_685 (.A(net184));
 sg13g2_antennanp ANTENNA_686 (.A(net184));
 sg13g2_antennanp ANTENNA_687 (.A(net184));
 sg13g2_antennanp ANTENNA_688 (.A(net184));
 sg13g2_antennanp ANTENNA_689 (.A(net184));
 sg13g2_antennanp ANTENNA_690 (.A(net184));
 sg13g2_antennanp ANTENNA_691 (.A(net184));
 sg13g2_antennanp ANTENNA_692 (.A(net184));
 sg13g2_antennanp ANTENNA_693 (.A(net184));
 sg13g2_antennanp ANTENNA_694 (.A(net184));
 sg13g2_antennanp ANTENNA_695 (.A(net184));
 sg13g2_antennanp ANTENNA_696 (.A(net184));
 sg13g2_antennanp ANTENNA_697 (.A(net184));
 sg13g2_antennanp ANTENNA_698 (.A(net192));
 sg13g2_antennanp ANTENNA_699 (.A(net192));
 sg13g2_antennanp ANTENNA_700 (.A(net192));
 sg13g2_antennanp ANTENNA_701 (.A(net192));
 sg13g2_antennanp ANTENNA_702 (.A(net192));
 sg13g2_antennanp ANTENNA_703 (.A(net192));
 sg13g2_antennanp ANTENNA_704 (.A(net192));
 sg13g2_antennanp ANTENNA_705 (.A(net192));
 sg13g2_antennanp ANTENNA_706 (.A(net192));
 sg13g2_antennanp ANTENNA_707 (.A(net192));
 sg13g2_antennanp ANTENNA_708 (.A(net192));
 sg13g2_antennanp ANTENNA_709 (.A(net192));
 sg13g2_antennanp ANTENNA_710 (.A(net192));
 sg13g2_antennanp ANTENNA_711 (.A(net192));
 sg13g2_antennanp ANTENNA_712 (.A(net202));
 sg13g2_antennanp ANTENNA_713 (.A(net202));
 sg13g2_antennanp ANTENNA_714 (.A(net202));
 sg13g2_antennanp ANTENNA_715 (.A(net202));
 sg13g2_antennanp ANTENNA_716 (.A(net202));
 sg13g2_antennanp ANTENNA_717 (.A(net202));
 sg13g2_antennanp ANTENNA_718 (.A(net202));
 sg13g2_antennanp ANTENNA_719 (.A(net202));
 sg13g2_antennanp ANTENNA_720 (.A(net202));
 sg13g2_antennanp ANTENNA_721 (.A(net205));
 sg13g2_antennanp ANTENNA_722 (.A(net205));
 sg13g2_antennanp ANTENNA_723 (.A(net205));
 sg13g2_antennanp ANTENNA_724 (.A(net205));
 sg13g2_antennanp ANTENNA_725 (.A(net205));
 sg13g2_antennanp ANTENNA_726 (.A(net205));
 sg13g2_antennanp ANTENNA_727 (.A(net205));
 sg13g2_antennanp ANTENNA_728 (.A(net205));
 sg13g2_antennanp ANTENNA_729 (.A(net205));
 sg13g2_antennanp ANTENNA_730 (.A(net206));
 sg13g2_antennanp ANTENNA_731 (.A(net206));
 sg13g2_antennanp ANTENNA_732 (.A(net206));
 sg13g2_antennanp ANTENNA_733 (.A(net206));
 sg13g2_antennanp ANTENNA_734 (.A(net206));
 sg13g2_antennanp ANTENNA_735 (.A(net206));
 sg13g2_antennanp ANTENNA_736 (.A(net206));
 sg13g2_antennanp ANTENNA_737 (.A(net206));
 sg13g2_antennanp ANTENNA_738 (.A(net206));
 sg13g2_antennanp ANTENNA_739 (.A(_2064_));
 sg13g2_antennanp ANTENNA_740 (.A(_2064_));
 sg13g2_antennanp ANTENNA_741 (.A(_2064_));
 sg13g2_antennanp ANTENNA_742 (.A(_2064_));
 sg13g2_antennanp ANTENNA_743 (.A(_2064_));
 sg13g2_antennanp ANTENNA_744 (.A(_2064_));
 sg13g2_antennanp ANTENNA_745 (.A(_2064_));
 sg13g2_antennanp ANTENNA_746 (.A(_2064_));
 sg13g2_antennanp ANTENNA_747 (.A(_2201_));
 sg13g2_antennanp ANTENNA_748 (.A(_2201_));
 sg13g2_antennanp ANTENNA_749 (.A(_2201_));
 sg13g2_antennanp ANTENNA_750 (.A(_2201_));
 sg13g2_antennanp ANTENNA_751 (.A(_2201_));
 sg13g2_antennanp ANTENNA_752 (.A(_2201_));
 sg13g2_antennanp ANTENNA_753 (.A(_2201_));
 sg13g2_antennanp ANTENNA_754 (.A(_2344_));
 sg13g2_antennanp ANTENNA_755 (.A(_2344_));
 sg13g2_antennanp ANTENNA_756 (.A(_2344_));
 sg13g2_antennanp ANTENNA_757 (.A(_2344_));
 sg13g2_antennanp ANTENNA_758 (.A(_2344_));
 sg13g2_antennanp ANTENNA_759 (.A(_2344_));
 sg13g2_antennanp ANTENNA_760 (.A(_2344_));
 sg13g2_antennanp ANTENNA_761 (.A(_2353_));
 sg13g2_antennanp ANTENNA_762 (.A(_2353_));
 sg13g2_antennanp ANTENNA_763 (.A(_2353_));
 sg13g2_antennanp ANTENNA_764 (.A(_2353_));
 sg13g2_antennanp ANTENNA_765 (.A(_2378_));
 sg13g2_antennanp ANTENNA_766 (.A(_2378_));
 sg13g2_antennanp ANTENNA_767 (.A(_2378_));
 sg13g2_antennanp ANTENNA_768 (.A(_2378_));
 sg13g2_antennanp ANTENNA_769 (.A(_2378_));
 sg13g2_antennanp ANTENNA_770 (.A(_2378_));
 sg13g2_antennanp ANTENNA_771 (.A(_2378_));
 sg13g2_antennanp ANTENNA_772 (.A(_2378_));
 sg13g2_antennanp ANTENNA_773 (.A(_2378_));
 sg13g2_antennanp ANTENNA_774 (.A(_2378_));
 sg13g2_antennanp ANTENNA_775 (.A(_2380_));
 sg13g2_antennanp ANTENNA_776 (.A(_2380_));
 sg13g2_antennanp ANTENNA_777 (.A(_2380_));
 sg13g2_antennanp ANTENNA_778 (.A(_2380_));
 sg13g2_antennanp ANTENNA_779 (.A(_2401_));
 sg13g2_antennanp ANTENNA_780 (.A(_2443_));
 sg13g2_antennanp ANTENNA_781 (.A(_2443_));
 sg13g2_antennanp ANTENNA_782 (.A(_2461_));
 sg13g2_antennanp ANTENNA_783 (.A(_2461_));
 sg13g2_antennanp ANTENNA_784 (.A(_2461_));
 sg13g2_antennanp ANTENNA_785 (.A(_2488_));
 sg13g2_antennanp ANTENNA_786 (.A(_2488_));
 sg13g2_antennanp ANTENNA_787 (.A(_2488_));
 sg13g2_antennanp ANTENNA_788 (.A(_2488_));
 sg13g2_antennanp ANTENNA_789 (.A(_2488_));
 sg13g2_antennanp ANTENNA_790 (.A(_2488_));
 sg13g2_antennanp ANTENNA_791 (.A(_2568_));
 sg13g2_antennanp ANTENNA_792 (.A(_2568_));
 sg13g2_antennanp ANTENNA_793 (.A(_2568_));
 sg13g2_antennanp ANTENNA_794 (.A(_2588_));
 sg13g2_antennanp ANTENNA_795 (.A(_2588_));
 sg13g2_antennanp ANTENNA_796 (.A(_2588_));
 sg13g2_antennanp ANTENNA_797 (.A(_2596_));
 sg13g2_antennanp ANTENNA_798 (.A(_2596_));
 sg13g2_antennanp ANTENNA_799 (.A(_2596_));
 sg13g2_antennanp ANTENNA_800 (.A(_2596_));
 sg13g2_antennanp ANTENNA_801 (.A(_2598_));
 sg13g2_antennanp ANTENNA_802 (.A(_2711_));
 sg13g2_antennanp ANTENNA_803 (.A(_2762_));
 sg13g2_antennanp ANTENNA_804 (.A(_2762_));
 sg13g2_antennanp ANTENNA_805 (.A(_2870_));
 sg13g2_antennanp ANTENNA_806 (.A(_2878_));
 sg13g2_antennanp ANTENNA_807 (.A(_2955_));
 sg13g2_antennanp ANTENNA_808 (.A(_2955_));
 sg13g2_antennanp ANTENNA_809 (.A(_2955_));
 sg13g2_antennanp ANTENNA_810 (.A(_2977_));
 sg13g2_antennanp ANTENNA_811 (.A(_2977_));
 sg13g2_antennanp ANTENNA_812 (.A(_2977_));
 sg13g2_antennanp ANTENNA_813 (.A(_2978_));
 sg13g2_antennanp ANTENNA_814 (.A(_2978_));
 sg13g2_antennanp ANTENNA_815 (.A(_2978_));
 sg13g2_antennanp ANTENNA_816 (.A(_2978_));
 sg13g2_antennanp ANTENNA_817 (.A(_2990_));
 sg13g2_antennanp ANTENNA_818 (.A(_2990_));
 sg13g2_antennanp ANTENNA_819 (.A(_2990_));
 sg13g2_antennanp ANTENNA_820 (.A(_2990_));
 sg13g2_antennanp ANTENNA_821 (.A(_3003_));
 sg13g2_antennanp ANTENNA_822 (.A(_3021_));
 sg13g2_antennanp ANTENNA_823 (.A(_3046_));
 sg13g2_antennanp ANTENNA_824 (.A(_3046_));
 sg13g2_antennanp ANTENNA_825 (.A(_3079_));
 sg13g2_antennanp ANTENNA_826 (.A(_3098_));
 sg13g2_antennanp ANTENNA_827 (.A(_3098_));
 sg13g2_antennanp ANTENNA_828 (.A(_3130_));
 sg13g2_antennanp ANTENNA_829 (.A(_3221_));
 sg13g2_antennanp ANTENNA_830 (.A(_3221_));
 sg13g2_antennanp ANTENNA_831 (.A(_3228_));
 sg13g2_antennanp ANTENNA_832 (.A(_3241_));
 sg13g2_antennanp ANTENNA_833 (.A(_3259_));
 sg13g2_antennanp ANTENNA_834 (.A(_3294_));
 sg13g2_antennanp ANTENNA_835 (.A(_3299_));
 sg13g2_antennanp ANTENNA_836 (.A(_3333_));
 sg13g2_antennanp ANTENNA_837 (.A(_3348_));
 sg13g2_antennanp ANTENNA_838 (.A(_3372_));
 sg13g2_antennanp ANTENNA_839 (.A(_3472_));
 sg13g2_antennanp ANTENNA_840 (.A(_3522_));
 sg13g2_antennanp ANTENNA_841 (.A(_3614_));
 sg13g2_antennanp ANTENNA_842 (.A(_3640_));
 sg13g2_antennanp ANTENNA_843 (.A(_3835_));
 sg13g2_antennanp ANTENNA_844 (.A(_3835_));
 sg13g2_antennanp ANTENNA_845 (.A(_3858_));
 sg13g2_antennanp ANTENNA_846 (.A(_3871_));
 sg13g2_antennanp ANTENNA_847 (.A(_3891_));
 sg13g2_antennanp ANTENNA_848 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_849 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_850 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_851 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_852 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_853 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_854 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_855 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_856 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_857 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_858 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_859 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_860 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_861 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_862 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_863 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_864 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_865 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_866 (.A(net10));
 sg13g2_antennanp ANTENNA_867 (.A(net15));
 sg13g2_antennanp ANTENNA_868 (.A(net15));
 sg13g2_antennanp ANTENNA_869 (.A(net15));
 sg13g2_antennanp ANTENNA_870 (.A(net17));
 sg13g2_antennanp ANTENNA_871 (.A(net17));
 sg13g2_antennanp ANTENNA_872 (.A(net17));
 sg13g2_antennanp ANTENNA_873 (.A(net21));
 sg13g2_antennanp ANTENNA_874 (.A(net21));
 sg13g2_antennanp ANTENNA_875 (.A(net21));
 sg13g2_antennanp ANTENNA_876 (.A(net21));
 sg13g2_antennanp ANTENNA_877 (.A(net21));
 sg13g2_antennanp ANTENNA_878 (.A(net21));
 sg13g2_antennanp ANTENNA_879 (.A(net21));
 sg13g2_antennanp ANTENNA_880 (.A(net21));
 sg13g2_antennanp ANTENNA_881 (.A(net23));
 sg13g2_antennanp ANTENNA_882 (.A(net23));
 sg13g2_antennanp ANTENNA_883 (.A(net23));
 sg13g2_antennanp ANTENNA_884 (.A(net23));
 sg13g2_antennanp ANTENNA_885 (.A(net23));
 sg13g2_antennanp ANTENNA_886 (.A(net23));
 sg13g2_antennanp ANTENNA_887 (.A(net23));
 sg13g2_antennanp ANTENNA_888 (.A(net23));
 sg13g2_antennanp ANTENNA_889 (.A(net61));
 sg13g2_antennanp ANTENNA_890 (.A(net61));
 sg13g2_antennanp ANTENNA_891 (.A(net61));
 sg13g2_antennanp ANTENNA_892 (.A(net61));
 sg13g2_antennanp ANTENNA_893 (.A(net61));
 sg13g2_antennanp ANTENNA_894 (.A(net61));
 sg13g2_antennanp ANTENNA_895 (.A(net61));
 sg13g2_antennanp ANTENNA_896 (.A(net61));
 sg13g2_antennanp ANTENNA_897 (.A(net68));
 sg13g2_antennanp ANTENNA_898 (.A(net68));
 sg13g2_antennanp ANTENNA_899 (.A(net68));
 sg13g2_antennanp ANTENNA_900 (.A(net68));
 sg13g2_antennanp ANTENNA_901 (.A(net68));
 sg13g2_antennanp ANTENNA_902 (.A(net68));
 sg13g2_antennanp ANTENNA_903 (.A(net68));
 sg13g2_antennanp ANTENNA_904 (.A(net68));
 sg13g2_antennanp ANTENNA_905 (.A(net68));
 sg13g2_antennanp ANTENNA_906 (.A(net70));
 sg13g2_antennanp ANTENNA_907 (.A(net70));
 sg13g2_antennanp ANTENNA_908 (.A(net70));
 sg13g2_antennanp ANTENNA_909 (.A(net70));
 sg13g2_antennanp ANTENNA_910 (.A(net70));
 sg13g2_antennanp ANTENNA_911 (.A(net70));
 sg13g2_antennanp ANTENNA_912 (.A(net70));
 sg13g2_antennanp ANTENNA_913 (.A(net70));
 sg13g2_antennanp ANTENNA_914 (.A(net70));
 sg13g2_antennanp ANTENNA_915 (.A(net73));
 sg13g2_antennanp ANTENNA_916 (.A(net73));
 sg13g2_antennanp ANTENNA_917 (.A(net73));
 sg13g2_antennanp ANTENNA_918 (.A(net73));
 sg13g2_antennanp ANTENNA_919 (.A(net73));
 sg13g2_antennanp ANTENNA_920 (.A(net73));
 sg13g2_antennanp ANTENNA_921 (.A(net73));
 sg13g2_antennanp ANTENNA_922 (.A(net73));
 sg13g2_antennanp ANTENNA_923 (.A(net73));
 sg13g2_antennanp ANTENNA_924 (.A(net74));
 sg13g2_antennanp ANTENNA_925 (.A(net74));
 sg13g2_antennanp ANTENNA_926 (.A(net74));
 sg13g2_antennanp ANTENNA_927 (.A(net74));
 sg13g2_antennanp ANTENNA_928 (.A(net74));
 sg13g2_antennanp ANTENNA_929 (.A(net74));
 sg13g2_antennanp ANTENNA_930 (.A(net74));
 sg13g2_antennanp ANTENNA_931 (.A(net74));
 sg13g2_antennanp ANTENNA_932 (.A(net74));
 sg13g2_antennanp ANTENNA_933 (.A(net79));
 sg13g2_antennanp ANTENNA_934 (.A(net79));
 sg13g2_antennanp ANTENNA_935 (.A(net79));
 sg13g2_antennanp ANTENNA_936 (.A(net79));
 sg13g2_antennanp ANTENNA_937 (.A(net79));
 sg13g2_antennanp ANTENNA_938 (.A(net79));
 sg13g2_antennanp ANTENNA_939 (.A(net79));
 sg13g2_antennanp ANTENNA_940 (.A(net79));
 sg13g2_antennanp ANTENNA_941 (.A(net79));
 sg13g2_antennanp ANTENNA_942 (.A(net85));
 sg13g2_antennanp ANTENNA_943 (.A(net85));
 sg13g2_antennanp ANTENNA_944 (.A(net85));
 sg13g2_antennanp ANTENNA_945 (.A(net85));
 sg13g2_antennanp ANTENNA_946 (.A(net85));
 sg13g2_antennanp ANTENNA_947 (.A(net85));
 sg13g2_antennanp ANTENNA_948 (.A(net85));
 sg13g2_antennanp ANTENNA_949 (.A(net85));
 sg13g2_antennanp ANTENNA_950 (.A(net85));
 sg13g2_antennanp ANTENNA_951 (.A(net92));
 sg13g2_antennanp ANTENNA_952 (.A(net92));
 sg13g2_antennanp ANTENNA_953 (.A(net92));
 sg13g2_antennanp ANTENNA_954 (.A(net92));
 sg13g2_antennanp ANTENNA_955 (.A(net92));
 sg13g2_antennanp ANTENNA_956 (.A(net92));
 sg13g2_antennanp ANTENNA_957 (.A(net92));
 sg13g2_antennanp ANTENNA_958 (.A(net92));
 sg13g2_antennanp ANTENNA_959 (.A(net163));
 sg13g2_antennanp ANTENNA_960 (.A(net163));
 sg13g2_antennanp ANTENNA_961 (.A(net163));
 sg13g2_antennanp ANTENNA_962 (.A(net163));
 sg13g2_antennanp ANTENNA_963 (.A(net163));
 sg13g2_antennanp ANTENNA_964 (.A(net163));
 sg13g2_antennanp ANTENNA_965 (.A(net163));
 sg13g2_antennanp ANTENNA_966 (.A(net163));
 sg13g2_antennanp ANTENNA_967 (.A(net163));
 sg13g2_antennanp ANTENNA_968 (.A(net174));
 sg13g2_antennanp ANTENNA_969 (.A(net174));
 sg13g2_antennanp ANTENNA_970 (.A(net174));
 sg13g2_antennanp ANTENNA_971 (.A(net174));
 sg13g2_antennanp ANTENNA_972 (.A(net174));
 sg13g2_antennanp ANTENNA_973 (.A(net174));
 sg13g2_antennanp ANTENNA_974 (.A(net174));
 sg13g2_antennanp ANTENNA_975 (.A(net174));
 sg13g2_antennanp ANTENNA_976 (.A(net184));
 sg13g2_antennanp ANTENNA_977 (.A(net184));
 sg13g2_antennanp ANTENNA_978 (.A(net184));
 sg13g2_antennanp ANTENNA_979 (.A(net184));
 sg13g2_antennanp ANTENNA_980 (.A(net184));
 sg13g2_antennanp ANTENNA_981 (.A(net184));
 sg13g2_antennanp ANTENNA_982 (.A(net184));
 sg13g2_antennanp ANTENNA_983 (.A(net184));
 sg13g2_antennanp ANTENNA_984 (.A(net184));
 sg13g2_antennanp ANTENNA_985 (.A(net184));
 sg13g2_antennanp ANTENNA_986 (.A(net184));
 sg13g2_antennanp ANTENNA_987 (.A(net184));
 sg13g2_antennanp ANTENNA_988 (.A(net184));
 sg13g2_antennanp ANTENNA_989 (.A(net202));
 sg13g2_antennanp ANTENNA_990 (.A(net202));
 sg13g2_antennanp ANTENNA_991 (.A(net202));
 sg13g2_antennanp ANTENNA_992 (.A(net202));
 sg13g2_antennanp ANTENNA_993 (.A(net202));
 sg13g2_antennanp ANTENNA_994 (.A(net202));
 sg13g2_antennanp ANTENNA_995 (.A(net202));
 sg13g2_antennanp ANTENNA_996 (.A(net202));
 sg13g2_antennanp ANTENNA_997 (.A(net202));
 sg13g2_antennanp ANTENNA_998 (.A(net205));
 sg13g2_antennanp ANTENNA_999 (.A(net205));
 sg13g2_antennanp ANTENNA_1000 (.A(net205));
 sg13g2_antennanp ANTENNA_1001 (.A(net205));
 sg13g2_antennanp ANTENNA_1002 (.A(net205));
 sg13g2_antennanp ANTENNA_1003 (.A(net205));
 sg13g2_antennanp ANTENNA_1004 (.A(net205));
 sg13g2_antennanp ANTENNA_1005 (.A(net205));
 sg13g2_antennanp ANTENNA_1006 (.A(net205));
 sg13g2_antennanp ANTENNA_1007 (.A(net206));
 sg13g2_antennanp ANTENNA_1008 (.A(net206));
 sg13g2_antennanp ANTENNA_1009 (.A(net206));
 sg13g2_antennanp ANTENNA_1010 (.A(net206));
 sg13g2_antennanp ANTENNA_1011 (.A(net206));
 sg13g2_antennanp ANTENNA_1012 (.A(net206));
 sg13g2_antennanp ANTENNA_1013 (.A(net206));
 sg13g2_antennanp ANTENNA_1014 (.A(net206));
 sg13g2_antennanp ANTENNA_1015 (.A(net206));
 sg13g2_antennanp ANTENNA_1016 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1017 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1018 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1019 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1020 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1021 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1022 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1023 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1024 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1025 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1026 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1027 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1028 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1029 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1030 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1031 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1032 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1033 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1034 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1035 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1036 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1037 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1038 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1039 (.A(_2353_));
 sg13g2_antennanp ANTENNA_1040 (.A(_2353_));
 sg13g2_antennanp ANTENNA_1041 (.A(_2353_));
 sg13g2_antennanp ANTENNA_1042 (.A(_2353_));
 sg13g2_antennanp ANTENNA_1043 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1044 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1045 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1046 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1047 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1048 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1049 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1050 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1051 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1052 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1053 (.A(_2380_));
 sg13g2_antennanp ANTENNA_1054 (.A(_2380_));
 sg13g2_antennanp ANTENNA_1055 (.A(_2380_));
 sg13g2_antennanp ANTENNA_1056 (.A(_2380_));
 sg13g2_antennanp ANTENNA_1057 (.A(_2401_));
 sg13g2_antennanp ANTENNA_1058 (.A(_2443_));
 sg13g2_antennanp ANTENNA_1059 (.A(_2443_));
 sg13g2_antennanp ANTENNA_1060 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1061 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1062 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1063 (.A(_2488_));
 sg13g2_antennanp ANTENNA_1064 (.A(_2488_));
 sg13g2_antennanp ANTENNA_1065 (.A(_2488_));
 sg13g2_antennanp ANTENNA_1066 (.A(_2568_));
 sg13g2_antennanp ANTENNA_1067 (.A(_2568_));
 sg13g2_antennanp ANTENNA_1068 (.A(_2568_));
 sg13g2_antennanp ANTENNA_1069 (.A(_2588_));
 sg13g2_antennanp ANTENNA_1070 (.A(_2588_));
 sg13g2_antennanp ANTENNA_1071 (.A(_2588_));
 sg13g2_antennanp ANTENNA_1072 (.A(_2596_));
 sg13g2_antennanp ANTENNA_1073 (.A(_2596_));
 sg13g2_antennanp ANTENNA_1074 (.A(_2596_));
 sg13g2_antennanp ANTENNA_1075 (.A(_2596_));
 sg13g2_antennanp ANTENNA_1076 (.A(_2598_));
 sg13g2_antennanp ANTENNA_1077 (.A(_2711_));
 sg13g2_antennanp ANTENNA_1078 (.A(_2762_));
 sg13g2_antennanp ANTENNA_1079 (.A(_2762_));
 sg13g2_antennanp ANTENNA_1080 (.A(_2870_));
 sg13g2_antennanp ANTENNA_1081 (.A(_2878_));
 sg13g2_antennanp ANTENNA_1082 (.A(_2955_));
 sg13g2_antennanp ANTENNA_1083 (.A(_2955_));
 sg13g2_antennanp ANTENNA_1084 (.A(_2955_));
 sg13g2_antennanp ANTENNA_1085 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1086 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1087 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1088 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1089 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1090 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1091 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1092 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1093 (.A(_2990_));
 sg13g2_antennanp ANTENNA_1094 (.A(_2990_));
 sg13g2_antennanp ANTENNA_1095 (.A(_2990_));
 sg13g2_antennanp ANTENNA_1096 (.A(_2990_));
 sg13g2_antennanp ANTENNA_1097 (.A(_3003_));
 sg13g2_antennanp ANTENNA_1098 (.A(_3003_));
 sg13g2_antennanp ANTENNA_1099 (.A(_3021_));
 sg13g2_antennanp ANTENNA_1100 (.A(_3046_));
 sg13g2_antennanp ANTENNA_1101 (.A(_3046_));
 sg13g2_antennanp ANTENNA_1102 (.A(_3046_));
 sg13g2_antennanp ANTENNA_1103 (.A(_3079_));
 sg13g2_antennanp ANTENNA_1104 (.A(_3098_));
 sg13g2_antennanp ANTENNA_1105 (.A(_3098_));
 sg13g2_antennanp ANTENNA_1106 (.A(_3130_));
 sg13g2_antennanp ANTENNA_1107 (.A(_3213_));
 sg13g2_antennanp ANTENNA_1108 (.A(_3221_));
 sg13g2_antennanp ANTENNA_1109 (.A(_3221_));
 sg13g2_antennanp ANTENNA_1110 (.A(_3228_));
 sg13g2_antennanp ANTENNA_1111 (.A(_3241_));
 sg13g2_antennanp ANTENNA_1112 (.A(_3259_));
 sg13g2_antennanp ANTENNA_1113 (.A(_3294_));
 sg13g2_antennanp ANTENNA_1114 (.A(_3299_));
 sg13g2_antennanp ANTENNA_1115 (.A(_3333_));
 sg13g2_antennanp ANTENNA_1116 (.A(_3348_));
 sg13g2_antennanp ANTENNA_1117 (.A(_3472_));
 sg13g2_antennanp ANTENNA_1118 (.A(_3522_));
 sg13g2_antennanp ANTENNA_1119 (.A(_3614_));
 sg13g2_antennanp ANTENNA_1120 (.A(_3640_));
 sg13g2_antennanp ANTENNA_1121 (.A(_3835_));
 sg13g2_antennanp ANTENNA_1122 (.A(_3835_));
 sg13g2_antennanp ANTENNA_1123 (.A(_3871_));
 sg13g2_antennanp ANTENNA_1124 (.A(_3891_));
 sg13g2_antennanp ANTENNA_1125 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1126 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1127 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1128 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1129 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1130 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1131 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1132 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1133 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1134 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1135 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_1136 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_1137 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_1138 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_1139 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_1140 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_1141 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_1142 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_1143 (.A(net15));
 sg13g2_antennanp ANTENNA_1144 (.A(net15));
 sg13g2_antennanp ANTENNA_1145 (.A(net15));
 sg13g2_antennanp ANTENNA_1146 (.A(net17));
 sg13g2_antennanp ANTENNA_1147 (.A(net17));
 sg13g2_antennanp ANTENNA_1148 (.A(net17));
 sg13g2_antennanp ANTENNA_1149 (.A(net23));
 sg13g2_antennanp ANTENNA_1150 (.A(net23));
 sg13g2_antennanp ANTENNA_1151 (.A(net23));
 sg13g2_antennanp ANTENNA_1152 (.A(net23));
 sg13g2_antennanp ANTENNA_1153 (.A(net23));
 sg13g2_antennanp ANTENNA_1154 (.A(net23));
 sg13g2_antennanp ANTENNA_1155 (.A(net23));
 sg13g2_antennanp ANTENNA_1156 (.A(net23));
 sg13g2_antennanp ANTENNA_1157 (.A(net43));
 sg13g2_antennanp ANTENNA_1158 (.A(net43));
 sg13g2_antennanp ANTENNA_1159 (.A(net43));
 sg13g2_antennanp ANTENNA_1160 (.A(net43));
 sg13g2_antennanp ANTENNA_1161 (.A(net43));
 sg13g2_antennanp ANTENNA_1162 (.A(net43));
 sg13g2_antennanp ANTENNA_1163 (.A(net43));
 sg13g2_antennanp ANTENNA_1164 (.A(net43));
 sg13g2_antennanp ANTENNA_1165 (.A(net61));
 sg13g2_antennanp ANTENNA_1166 (.A(net61));
 sg13g2_antennanp ANTENNA_1167 (.A(net61));
 sg13g2_antennanp ANTENNA_1168 (.A(net61));
 sg13g2_antennanp ANTENNA_1169 (.A(net61));
 sg13g2_antennanp ANTENNA_1170 (.A(net61));
 sg13g2_antennanp ANTENNA_1171 (.A(net61));
 sg13g2_antennanp ANTENNA_1172 (.A(net61));
 sg13g2_antennanp ANTENNA_1173 (.A(net68));
 sg13g2_antennanp ANTENNA_1174 (.A(net68));
 sg13g2_antennanp ANTENNA_1175 (.A(net68));
 sg13g2_antennanp ANTENNA_1176 (.A(net68));
 sg13g2_antennanp ANTENNA_1177 (.A(net68));
 sg13g2_antennanp ANTENNA_1178 (.A(net68));
 sg13g2_antennanp ANTENNA_1179 (.A(net68));
 sg13g2_antennanp ANTENNA_1180 (.A(net68));
 sg13g2_antennanp ANTENNA_1181 (.A(net68));
 sg13g2_antennanp ANTENNA_1182 (.A(net70));
 sg13g2_antennanp ANTENNA_1183 (.A(net70));
 sg13g2_antennanp ANTENNA_1184 (.A(net70));
 sg13g2_antennanp ANTENNA_1185 (.A(net70));
 sg13g2_antennanp ANTENNA_1186 (.A(net70));
 sg13g2_antennanp ANTENNA_1187 (.A(net70));
 sg13g2_antennanp ANTENNA_1188 (.A(net70));
 sg13g2_antennanp ANTENNA_1189 (.A(net70));
 sg13g2_antennanp ANTENNA_1190 (.A(net70));
 sg13g2_antennanp ANTENNA_1191 (.A(net73));
 sg13g2_antennanp ANTENNA_1192 (.A(net73));
 sg13g2_antennanp ANTENNA_1193 (.A(net73));
 sg13g2_antennanp ANTENNA_1194 (.A(net73));
 sg13g2_antennanp ANTENNA_1195 (.A(net73));
 sg13g2_antennanp ANTENNA_1196 (.A(net73));
 sg13g2_antennanp ANTENNA_1197 (.A(net73));
 sg13g2_antennanp ANTENNA_1198 (.A(net73));
 sg13g2_antennanp ANTENNA_1199 (.A(net73));
 sg13g2_antennanp ANTENNA_1200 (.A(net74));
 sg13g2_antennanp ANTENNA_1201 (.A(net74));
 sg13g2_antennanp ANTENNA_1202 (.A(net74));
 sg13g2_antennanp ANTENNA_1203 (.A(net74));
 sg13g2_antennanp ANTENNA_1204 (.A(net74));
 sg13g2_antennanp ANTENNA_1205 (.A(net74));
 sg13g2_antennanp ANTENNA_1206 (.A(net74));
 sg13g2_antennanp ANTENNA_1207 (.A(net74));
 sg13g2_antennanp ANTENNA_1208 (.A(net74));
 sg13g2_antennanp ANTENNA_1209 (.A(net79));
 sg13g2_antennanp ANTENNA_1210 (.A(net79));
 sg13g2_antennanp ANTENNA_1211 (.A(net79));
 sg13g2_antennanp ANTENNA_1212 (.A(net79));
 sg13g2_antennanp ANTENNA_1213 (.A(net79));
 sg13g2_antennanp ANTENNA_1214 (.A(net79));
 sg13g2_antennanp ANTENNA_1215 (.A(net79));
 sg13g2_antennanp ANTENNA_1216 (.A(net79));
 sg13g2_antennanp ANTENNA_1217 (.A(net79));
 sg13g2_antennanp ANTENNA_1218 (.A(net85));
 sg13g2_antennanp ANTENNA_1219 (.A(net85));
 sg13g2_antennanp ANTENNA_1220 (.A(net85));
 sg13g2_antennanp ANTENNA_1221 (.A(net85));
 sg13g2_antennanp ANTENNA_1222 (.A(net85));
 sg13g2_antennanp ANTENNA_1223 (.A(net85));
 sg13g2_antennanp ANTENNA_1224 (.A(net85));
 sg13g2_antennanp ANTENNA_1225 (.A(net85));
 sg13g2_antennanp ANTENNA_1226 (.A(net85));
 sg13g2_antennanp ANTENNA_1227 (.A(net92));
 sg13g2_antennanp ANTENNA_1228 (.A(net92));
 sg13g2_antennanp ANTENNA_1229 (.A(net92));
 sg13g2_antennanp ANTENNA_1230 (.A(net92));
 sg13g2_antennanp ANTENNA_1231 (.A(net92));
 sg13g2_antennanp ANTENNA_1232 (.A(net92));
 sg13g2_antennanp ANTENNA_1233 (.A(net92));
 sg13g2_antennanp ANTENNA_1234 (.A(net92));
 sg13g2_antennanp ANTENNA_1235 (.A(net163));
 sg13g2_antennanp ANTENNA_1236 (.A(net163));
 sg13g2_antennanp ANTENNA_1237 (.A(net163));
 sg13g2_antennanp ANTENNA_1238 (.A(net163));
 sg13g2_antennanp ANTENNA_1239 (.A(net163));
 sg13g2_antennanp ANTENNA_1240 (.A(net163));
 sg13g2_antennanp ANTENNA_1241 (.A(net163));
 sg13g2_antennanp ANTENNA_1242 (.A(net163));
 sg13g2_antennanp ANTENNA_1243 (.A(net163));
 sg13g2_antennanp ANTENNA_1244 (.A(net174));
 sg13g2_antennanp ANTENNA_1245 (.A(net174));
 sg13g2_antennanp ANTENNA_1246 (.A(net174));
 sg13g2_antennanp ANTENNA_1247 (.A(net174));
 sg13g2_antennanp ANTENNA_1248 (.A(net174));
 sg13g2_antennanp ANTENNA_1249 (.A(net174));
 sg13g2_antennanp ANTENNA_1250 (.A(net174));
 sg13g2_antennanp ANTENNA_1251 (.A(net174));
 sg13g2_antennanp ANTENNA_1252 (.A(net184));
 sg13g2_antennanp ANTENNA_1253 (.A(net184));
 sg13g2_antennanp ANTENNA_1254 (.A(net184));
 sg13g2_antennanp ANTENNA_1255 (.A(net184));
 sg13g2_antennanp ANTENNA_1256 (.A(net184));
 sg13g2_antennanp ANTENNA_1257 (.A(net184));
 sg13g2_antennanp ANTENNA_1258 (.A(net184));
 sg13g2_antennanp ANTENNA_1259 (.A(net184));
 sg13g2_antennanp ANTENNA_1260 (.A(net184));
 sg13g2_antennanp ANTENNA_1261 (.A(net184));
 sg13g2_antennanp ANTENNA_1262 (.A(net184));
 sg13g2_antennanp ANTENNA_1263 (.A(net184));
 sg13g2_antennanp ANTENNA_1264 (.A(net184));
 sg13g2_antennanp ANTENNA_1265 (.A(net184));
 sg13g2_antennanp ANTENNA_1266 (.A(net184));
 sg13g2_antennanp ANTENNA_1267 (.A(net184));
 sg13g2_antennanp ANTENNA_1268 (.A(net184));
 sg13g2_antennanp ANTENNA_1269 (.A(net202));
 sg13g2_antennanp ANTENNA_1270 (.A(net202));
 sg13g2_antennanp ANTENNA_1271 (.A(net202));
 sg13g2_antennanp ANTENNA_1272 (.A(net202));
 sg13g2_antennanp ANTENNA_1273 (.A(net202));
 sg13g2_antennanp ANTENNA_1274 (.A(net202));
 sg13g2_antennanp ANTENNA_1275 (.A(net202));
 sg13g2_antennanp ANTENNA_1276 (.A(net202));
 sg13g2_antennanp ANTENNA_1277 (.A(net202));
 sg13g2_antennanp ANTENNA_1278 (.A(net205));
 sg13g2_antennanp ANTENNA_1279 (.A(net205));
 sg13g2_antennanp ANTENNA_1280 (.A(net205));
 sg13g2_antennanp ANTENNA_1281 (.A(net205));
 sg13g2_antennanp ANTENNA_1282 (.A(net205));
 sg13g2_antennanp ANTENNA_1283 (.A(net205));
 sg13g2_antennanp ANTENNA_1284 (.A(net205));
 sg13g2_antennanp ANTENNA_1285 (.A(net205));
 sg13g2_antennanp ANTENNA_1286 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1287 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1288 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1289 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1290 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1291 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1292 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1293 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1294 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1295 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1296 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1297 (.A(_2064_));
 sg13g2_antennanp ANTENNA_1298 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1299 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1300 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1301 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1302 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1303 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1304 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1305 (.A(_2201_));
 sg13g2_antennanp ANTENNA_1306 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1307 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1308 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1309 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1310 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1311 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1312 (.A(_2344_));
 sg13g2_antennanp ANTENNA_1313 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1314 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1315 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1316 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1317 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1318 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1319 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1320 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1321 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1322 (.A(_2378_));
 sg13g2_antennanp ANTENNA_1323 (.A(_2380_));
 sg13g2_antennanp ANTENNA_1324 (.A(_2380_));
 sg13g2_antennanp ANTENNA_1325 (.A(_2380_));
 sg13g2_antennanp ANTENNA_1326 (.A(_2380_));
 sg13g2_antennanp ANTENNA_1327 (.A(_2401_));
 sg13g2_antennanp ANTENNA_1328 (.A(_2401_));
 sg13g2_antennanp ANTENNA_1329 (.A(_2443_));
 sg13g2_antennanp ANTENNA_1330 (.A(_2443_));
 sg13g2_antennanp ANTENNA_1331 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1332 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1333 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1334 (.A(_2473_));
 sg13g2_antennanp ANTENNA_1335 (.A(_2473_));
 sg13g2_antennanp ANTENNA_1336 (.A(_2473_));
 sg13g2_antennanp ANTENNA_1337 (.A(_2488_));
 sg13g2_antennanp ANTENNA_1338 (.A(_2488_));
 sg13g2_antennanp ANTENNA_1339 (.A(_2488_));
 sg13g2_antennanp ANTENNA_1340 (.A(_2488_));
 sg13g2_antennanp ANTENNA_1341 (.A(_2568_));
 sg13g2_antennanp ANTENNA_1342 (.A(_2568_));
 sg13g2_antennanp ANTENNA_1343 (.A(_2568_));
 sg13g2_antennanp ANTENNA_1344 (.A(_2588_));
 sg13g2_antennanp ANTENNA_1345 (.A(_2588_));
 sg13g2_antennanp ANTENNA_1346 (.A(_2588_));
 sg13g2_antennanp ANTENNA_1347 (.A(_2596_));
 sg13g2_antennanp ANTENNA_1348 (.A(_2596_));
 sg13g2_antennanp ANTENNA_1349 (.A(_2596_));
 sg13g2_antennanp ANTENNA_1350 (.A(_2596_));
 sg13g2_antennanp ANTENNA_1351 (.A(_2711_));
 sg13g2_antennanp ANTENNA_1352 (.A(_2762_));
 sg13g2_antennanp ANTENNA_1353 (.A(_2870_));
 sg13g2_antennanp ANTENNA_1354 (.A(_2878_));
 sg13g2_antennanp ANTENNA_1355 (.A(_2955_));
 sg13g2_antennanp ANTENNA_1356 (.A(_2955_));
 sg13g2_antennanp ANTENNA_1357 (.A(_2955_));
 sg13g2_antennanp ANTENNA_1358 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1359 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1360 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1361 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1362 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1363 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1364 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1365 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1366 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1367 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1368 (.A(_2978_));
 sg13g2_antennanp ANTENNA_1369 (.A(_2990_));
 sg13g2_antennanp ANTENNA_1370 (.A(_2990_));
 sg13g2_antennanp ANTENNA_1371 (.A(_2990_));
 sg13g2_antennanp ANTENNA_1372 (.A(_2990_));
 sg13g2_antennanp ANTENNA_1373 (.A(_3003_));
 sg13g2_antennanp ANTENNA_1374 (.A(_3021_));
 sg13g2_antennanp ANTENNA_1375 (.A(_3046_));
 sg13g2_antennanp ANTENNA_1376 (.A(_3046_));
 sg13g2_antennanp ANTENNA_1377 (.A(_3079_));
 sg13g2_antennanp ANTENNA_1378 (.A(_3098_));
 sg13g2_antennanp ANTENNA_1379 (.A(_3098_));
 sg13g2_antennanp ANTENNA_1380 (.A(_3130_));
 sg13g2_antennanp ANTENNA_1381 (.A(_3213_));
 sg13g2_antennanp ANTENNA_1382 (.A(_3221_));
 sg13g2_antennanp ANTENNA_1383 (.A(_3221_));
 sg13g2_antennanp ANTENNA_1384 (.A(_3228_));
 sg13g2_antennanp ANTENNA_1385 (.A(_3241_));
 sg13g2_antennanp ANTENNA_1386 (.A(_3259_));
 sg13g2_antennanp ANTENNA_1387 (.A(_3294_));
 sg13g2_antennanp ANTENNA_1388 (.A(_3299_));
 sg13g2_antennanp ANTENNA_1389 (.A(_3333_));
 sg13g2_antennanp ANTENNA_1390 (.A(_3348_));
 sg13g2_antennanp ANTENNA_1391 (.A(_3472_));
 sg13g2_antennanp ANTENNA_1392 (.A(_3522_));
 sg13g2_antennanp ANTENNA_1393 (.A(_3614_));
 sg13g2_antennanp ANTENNA_1394 (.A(_3640_));
 sg13g2_antennanp ANTENNA_1395 (.A(_3835_));
 sg13g2_antennanp ANTENNA_1396 (.A(_3835_));
 sg13g2_antennanp ANTENNA_1397 (.A(_3871_));
 sg13g2_antennanp ANTENNA_1398 (.A(_3891_));
 sg13g2_antennanp ANTENNA_1399 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1400 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1401 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1402 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1403 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1404 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1405 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1406 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1407 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1408 (.A(\logix.ram_r[1280] ));
 sg13g2_antennanp ANTENNA_1409 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_1410 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_1411 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_1412 (.A(\logix.ram_r[1408] ));
 sg13g2_antennanp ANTENNA_1413 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_1414 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_1415 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_1416 (.A(\logix.ram_r[383] ));
 sg13g2_antennanp ANTENNA_1417 (.A(net61));
 sg13g2_antennanp ANTENNA_1418 (.A(net61));
 sg13g2_antennanp ANTENNA_1419 (.A(net61));
 sg13g2_antennanp ANTENNA_1420 (.A(net61));
 sg13g2_antennanp ANTENNA_1421 (.A(net61));
 sg13g2_antennanp ANTENNA_1422 (.A(net61));
 sg13g2_antennanp ANTENNA_1423 (.A(net61));
 sg13g2_antennanp ANTENNA_1424 (.A(net61));
 sg13g2_antennanp ANTENNA_1425 (.A(net68));
 sg13g2_antennanp ANTENNA_1426 (.A(net68));
 sg13g2_antennanp ANTENNA_1427 (.A(net68));
 sg13g2_antennanp ANTENNA_1428 (.A(net68));
 sg13g2_antennanp ANTENNA_1429 (.A(net68));
 sg13g2_antennanp ANTENNA_1430 (.A(net68));
 sg13g2_antennanp ANTENNA_1431 (.A(net68));
 sg13g2_antennanp ANTENNA_1432 (.A(net68));
 sg13g2_antennanp ANTENNA_1433 (.A(net68));
 sg13g2_antennanp ANTENNA_1434 (.A(net70));
 sg13g2_antennanp ANTENNA_1435 (.A(net70));
 sg13g2_antennanp ANTENNA_1436 (.A(net70));
 sg13g2_antennanp ANTENNA_1437 (.A(net70));
 sg13g2_antennanp ANTENNA_1438 (.A(net70));
 sg13g2_antennanp ANTENNA_1439 (.A(net70));
 sg13g2_antennanp ANTENNA_1440 (.A(net70));
 sg13g2_antennanp ANTENNA_1441 (.A(net70));
 sg13g2_antennanp ANTENNA_1442 (.A(net70));
 sg13g2_antennanp ANTENNA_1443 (.A(net73));
 sg13g2_antennanp ANTENNA_1444 (.A(net73));
 sg13g2_antennanp ANTENNA_1445 (.A(net73));
 sg13g2_antennanp ANTENNA_1446 (.A(net73));
 sg13g2_antennanp ANTENNA_1447 (.A(net73));
 sg13g2_antennanp ANTENNA_1448 (.A(net73));
 sg13g2_antennanp ANTENNA_1449 (.A(net73));
 sg13g2_antennanp ANTENNA_1450 (.A(net73));
 sg13g2_antennanp ANTENNA_1451 (.A(net73));
 sg13g2_antennanp ANTENNA_1452 (.A(net74));
 sg13g2_antennanp ANTENNA_1453 (.A(net74));
 sg13g2_antennanp ANTENNA_1454 (.A(net74));
 sg13g2_antennanp ANTENNA_1455 (.A(net74));
 sg13g2_antennanp ANTENNA_1456 (.A(net74));
 sg13g2_antennanp ANTENNA_1457 (.A(net74));
 sg13g2_antennanp ANTENNA_1458 (.A(net74));
 sg13g2_antennanp ANTENNA_1459 (.A(net74));
 sg13g2_antennanp ANTENNA_1460 (.A(net74));
 sg13g2_antennanp ANTENNA_1461 (.A(net79));
 sg13g2_antennanp ANTENNA_1462 (.A(net79));
 sg13g2_antennanp ANTENNA_1463 (.A(net79));
 sg13g2_antennanp ANTENNA_1464 (.A(net79));
 sg13g2_antennanp ANTENNA_1465 (.A(net79));
 sg13g2_antennanp ANTENNA_1466 (.A(net79));
 sg13g2_antennanp ANTENNA_1467 (.A(net79));
 sg13g2_antennanp ANTENNA_1468 (.A(net79));
 sg13g2_antennanp ANTENNA_1469 (.A(net79));
 sg13g2_antennanp ANTENNA_1470 (.A(net85));
 sg13g2_antennanp ANTENNA_1471 (.A(net85));
 sg13g2_antennanp ANTENNA_1472 (.A(net85));
 sg13g2_antennanp ANTENNA_1473 (.A(net85));
 sg13g2_antennanp ANTENNA_1474 (.A(net85));
 sg13g2_antennanp ANTENNA_1475 (.A(net85));
 sg13g2_antennanp ANTENNA_1476 (.A(net85));
 sg13g2_antennanp ANTENNA_1477 (.A(net85));
 sg13g2_antennanp ANTENNA_1478 (.A(net85));
 sg13g2_antennanp ANTENNA_1479 (.A(net92));
 sg13g2_antennanp ANTENNA_1480 (.A(net92));
 sg13g2_antennanp ANTENNA_1481 (.A(net92));
 sg13g2_antennanp ANTENNA_1482 (.A(net92));
 sg13g2_antennanp ANTENNA_1483 (.A(net92));
 sg13g2_antennanp ANTENNA_1484 (.A(net92));
 sg13g2_antennanp ANTENNA_1485 (.A(net92));
 sg13g2_antennanp ANTENNA_1486 (.A(net92));
 sg13g2_antennanp ANTENNA_1487 (.A(net163));
 sg13g2_antennanp ANTENNA_1488 (.A(net163));
 sg13g2_antennanp ANTENNA_1489 (.A(net163));
 sg13g2_antennanp ANTENNA_1490 (.A(net163));
 sg13g2_antennanp ANTENNA_1491 (.A(net163));
 sg13g2_antennanp ANTENNA_1492 (.A(net163));
 sg13g2_antennanp ANTENNA_1493 (.A(net163));
 sg13g2_antennanp ANTENNA_1494 (.A(net163));
 sg13g2_antennanp ANTENNA_1495 (.A(net184));
 sg13g2_antennanp ANTENNA_1496 (.A(net184));
 sg13g2_antennanp ANTENNA_1497 (.A(net184));
 sg13g2_antennanp ANTENNA_1498 (.A(net184));
 sg13g2_antennanp ANTENNA_1499 (.A(net184));
 sg13g2_antennanp ANTENNA_1500 (.A(net184));
 sg13g2_antennanp ANTENNA_1501 (.A(net184));
 sg13g2_antennanp ANTENNA_1502 (.A(net184));
 sg13g2_antennanp ANTENNA_1503 (.A(net184));
 sg13g2_antennanp ANTENNA_1504 (.A(net202));
 sg13g2_antennanp ANTENNA_1505 (.A(net202));
 sg13g2_antennanp ANTENNA_1506 (.A(net202));
 sg13g2_antennanp ANTENNA_1507 (.A(net202));
 sg13g2_antennanp ANTENNA_1508 (.A(net202));
 sg13g2_antennanp ANTENNA_1509 (.A(net202));
 sg13g2_antennanp ANTENNA_1510 (.A(net202));
 sg13g2_antennanp ANTENNA_1511 (.A(net202));
 sg13g2_antennanp ANTENNA_1512 (.A(net202));
 sg13g2_antennanp ANTENNA_1513 (.A(net205));
 sg13g2_antennanp ANTENNA_1514 (.A(net205));
 sg13g2_antennanp ANTENNA_1515 (.A(net205));
 sg13g2_antennanp ANTENNA_1516 (.A(net205));
 sg13g2_antennanp ANTENNA_1517 (.A(net205));
 sg13g2_antennanp ANTENNA_1518 (.A(net205));
 sg13g2_antennanp ANTENNA_1519 (.A(net205));
 sg13g2_antennanp ANTENNA_1520 (.A(net205));
 sg13g2_antennanp ANTENNA_1521 (.A(net207));
 sg13g2_antennanp ANTENNA_1522 (.A(net207));
 sg13g2_antennanp ANTENNA_1523 (.A(net207));
 sg13g2_antennanp ANTENNA_1524 (.A(net207));
 sg13g2_antennanp ANTENNA_1525 (.A(net207));
 sg13g2_antennanp ANTENNA_1526 (.A(net207));
 sg13g2_antennanp ANTENNA_1527 (.A(net207));
 sg13g2_antennanp ANTENNA_1528 (.A(net207));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_fill_1 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_67 ();
 sg13g2_decap_8 FILLER_0_74 ();
 sg13g2_decap_8 FILLER_0_81 ();
 sg13g2_fill_2 FILLER_0_88 ();
 sg13g2_fill_1 FILLER_0_90 ();
 sg13g2_decap_8 FILLER_0_95 ();
 sg13g2_decap_8 FILLER_0_102 ();
 sg13g2_decap_4 FILLER_0_109 ();
 sg13g2_fill_1 FILLER_0_113 ();
 sg13g2_fill_1 FILLER_0_124 ();
 sg13g2_decap_8 FILLER_0_129 ();
 sg13g2_decap_8 FILLER_0_136 ();
 sg13g2_decap_8 FILLER_0_143 ();
 sg13g2_decap_8 FILLER_0_150 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_fill_2 FILLER_0_164 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_fill_1 FILLER_0_206 ();
 sg13g2_fill_2 FILLER_0_217 ();
 sg13g2_fill_1 FILLER_0_219 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_fill_2 FILLER_0_257 ();
 sg13g2_fill_1 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_4 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_8 FILLER_0_321 ();
 sg13g2_decap_8 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_4 FILLER_0_342 ();
 sg13g2_fill_1 FILLER_0_346 ();
 sg13g2_fill_1 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_fill_2 FILLER_0_397 ();
 sg13g2_fill_1 FILLER_0_399 ();
 sg13g2_fill_1 FILLER_0_430 ();
 sg13g2_decap_8 FILLER_0_435 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_fill_1 FILLER_0_449 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_4 FILLER_0_483 ();
 sg13g2_fill_2 FILLER_0_487 ();
 sg13g2_decap_8 FILLER_0_515 ();
 sg13g2_decap_8 FILLER_0_522 ();
 sg13g2_decap_8 FILLER_0_529 ();
 sg13g2_decap_8 FILLER_0_536 ();
 sg13g2_fill_2 FILLER_0_543 ();
 sg13g2_fill_1 FILLER_0_545 ();
 sg13g2_decap_8 FILLER_0_576 ();
 sg13g2_decap_8 FILLER_0_583 ();
 sg13g2_decap_8 FILLER_0_590 ();
 sg13g2_decap_4 FILLER_0_597 ();
 sg13g2_fill_1 FILLER_0_601 ();
 sg13g2_decap_8 FILLER_0_628 ();
 sg13g2_decap_8 FILLER_0_635 ();
 sg13g2_decap_4 FILLER_0_642 ();
 sg13g2_fill_1 FILLER_0_646 ();
 sg13g2_fill_1 FILLER_0_651 ();
 sg13g2_decap_4 FILLER_0_656 ();
 sg13g2_fill_1 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_695 ();
 sg13g2_decap_8 FILLER_0_702 ();
 sg13g2_decap_8 FILLER_0_709 ();
 sg13g2_decap_8 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_723 ();
 sg13g2_decap_8 FILLER_0_730 ();
 sg13g2_fill_2 FILLER_0_737 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_fill_1 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_797 ();
 sg13g2_decap_8 FILLER_0_804 ();
 sg13g2_decap_8 FILLER_0_811 ();
 sg13g2_decap_8 FILLER_0_818 ();
 sg13g2_fill_1 FILLER_0_825 ();
 sg13g2_decap_4 FILLER_0_834 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_4 FILLER_0_889 ();
 sg13g2_fill_2 FILLER_0_893 ();
 sg13g2_decap_8 FILLER_0_921 ();
 sg13g2_decap_8 FILLER_0_928 ();
 sg13g2_decap_8 FILLER_0_935 ();
 sg13g2_decap_8 FILLER_0_942 ();
 sg13g2_fill_2 FILLER_0_949 ();
 sg13g2_fill_1 FILLER_0_951 ();
 sg13g2_decap_8 FILLER_0_982 ();
 sg13g2_decap_8 FILLER_0_989 ();
 sg13g2_decap_4 FILLER_0_996 ();
 sg13g2_decap_8 FILLER_0_1036 ();
 sg13g2_decap_8 FILLER_0_1043 ();
 sg13g2_decap_8 FILLER_0_1050 ();
 sg13g2_decap_4 FILLER_0_1057 ();
 sg13g2_fill_1 FILLER_0_1061 ();
 sg13g2_decap_8 FILLER_0_1088 ();
 sg13g2_decap_4 FILLER_0_1095 ();
 sg13g2_fill_2 FILLER_0_1099 ();
 sg13g2_fill_2 FILLER_0_1111 ();
 sg13g2_fill_1 FILLER_0_1113 ();
 sg13g2_decap_8 FILLER_0_1124 ();
 sg13g2_decap_8 FILLER_0_1131 ();
 sg13g2_decap_8 FILLER_0_1138 ();
 sg13g2_decap_8 FILLER_0_1145 ();
 sg13g2_decap_8 FILLER_0_1152 ();
 sg13g2_decap_8 FILLER_0_1159 ();
 sg13g2_decap_8 FILLER_0_1166 ();
 sg13g2_decap_8 FILLER_0_1173 ();
 sg13g2_decap_8 FILLER_0_1180 ();
 sg13g2_decap_8 FILLER_0_1187 ();
 sg13g2_fill_2 FILLER_0_1194 ();
 sg13g2_decap_4 FILLER_0_1222 ();
 sg13g2_fill_1 FILLER_0_1226 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_4 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1268 ();
 sg13g2_decap_8 FILLER_0_1275 ();
 sg13g2_decap_8 FILLER_0_1282 ();
 sg13g2_decap_4 FILLER_0_1289 ();
 sg13g2_decap_8 FILLER_0_1297 ();
 sg13g2_decap_8 FILLER_0_1304 ();
 sg13g2_decap_8 FILLER_0_1311 ();
 sg13g2_fill_1 FILLER_0_1318 ();
 sg13g2_decap_4 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1331 ();
 sg13g2_decap_8 FILLER_0_1338 ();
 sg13g2_decap_8 FILLER_0_1345 ();
 sg13g2_decap_8 FILLER_0_1352 ();
 sg13g2_decap_8 FILLER_0_1359 ();
 sg13g2_decap_8 FILLER_0_1366 ();
 sg13g2_decap_4 FILLER_0_1373 ();
 sg13g2_fill_2 FILLER_0_1377 ();
 sg13g2_decap_8 FILLER_0_1405 ();
 sg13g2_decap_8 FILLER_0_1412 ();
 sg13g2_decap_8 FILLER_0_1419 ();
 sg13g2_decap_8 FILLER_0_1426 ();
 sg13g2_decap_8 FILLER_0_1433 ();
 sg13g2_decap_4 FILLER_0_1440 ();
 sg13g2_fill_1 FILLER_0_1444 ();
 sg13g2_decap_8 FILLER_0_1466 ();
 sg13g2_decap_8 FILLER_0_1473 ();
 sg13g2_decap_8 FILLER_0_1480 ();
 sg13g2_decap_8 FILLER_0_1487 ();
 sg13g2_decap_8 FILLER_0_1494 ();
 sg13g2_decap_8 FILLER_0_1501 ();
 sg13g2_decap_8 FILLER_0_1508 ();
 sg13g2_fill_2 FILLER_0_1515 ();
 sg13g2_fill_1 FILLER_0_1517 ();
 sg13g2_decap_8 FILLER_0_1544 ();
 sg13g2_decap_8 FILLER_0_1551 ();
 sg13g2_decap_8 FILLER_0_1558 ();
 sg13g2_decap_8 FILLER_0_1565 ();
 sg13g2_fill_1 FILLER_0_1572 ();
 sg13g2_decap_8 FILLER_0_1599 ();
 sg13g2_fill_2 FILLER_0_1606 ();
 sg13g2_fill_1 FILLER_0_1608 ();
 sg13g2_decap_8 FILLER_0_1635 ();
 sg13g2_decap_8 FILLER_0_1642 ();
 sg13g2_decap_4 FILLER_0_1649 ();
 sg13g2_fill_2 FILLER_0_1653 ();
 sg13g2_decap_8 FILLER_0_1665 ();
 sg13g2_decap_8 FILLER_0_1672 ();
 sg13g2_decap_8 FILLER_0_1679 ();
 sg13g2_decap_8 FILLER_0_1686 ();
 sg13g2_decap_8 FILLER_0_1693 ();
 sg13g2_decap_8 FILLER_0_1700 ();
 sg13g2_decap_8 FILLER_0_1707 ();
 sg13g2_decap_8 FILLER_0_1714 ();
 sg13g2_decap_8 FILLER_0_1721 ();
 sg13g2_decap_8 FILLER_0_1728 ();
 sg13g2_decap_8 FILLER_0_1735 ();
 sg13g2_decap_8 FILLER_0_1742 ();
 sg13g2_decap_8 FILLER_0_1749 ();
 sg13g2_decap_8 FILLER_0_1756 ();
 sg13g2_decap_8 FILLER_0_1763 ();
 sg13g2_decap_4 FILLER_0_1770 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_fill_1 FILLER_1_21 ();
 sg13g2_fill_2 FILLER_1_36 ();
 sg13g2_fill_1 FILLER_1_38 ();
 sg13g2_decap_4 FILLER_1_79 ();
 sg13g2_fill_1 FILLER_1_83 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_4 FILLER_1_168 ();
 sg13g2_fill_1 FILLER_1_172 ();
 sg13g2_fill_2 FILLER_1_223 ();
 sg13g2_fill_2 FILLER_1_235 ();
 sg13g2_decap_4 FILLER_1_267 ();
 sg13g2_fill_2 FILLER_1_271 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_fill_2 FILLER_1_331 ();
 sg13g2_fill_1 FILLER_1_347 ();
 sg13g2_fill_1 FILLER_1_374 ();
 sg13g2_fill_1 FILLER_1_401 ();
 sg13g2_fill_2 FILLER_1_412 ();
 sg13g2_decap_8 FILLER_1_486 ();
 sg13g2_fill_1 FILLER_1_493 ();
 sg13g2_decap_8 FILLER_1_528 ();
 sg13g2_decap_8 FILLER_1_535 ();
 sg13g2_fill_2 FILLER_1_542 ();
 sg13g2_fill_1 FILLER_1_544 ();
 sg13g2_decap_4 FILLER_1_549 ();
 sg13g2_decap_4 FILLER_1_599 ();
 sg13g2_decap_8 FILLER_1_617 ();
 sg13g2_decap_8 FILLER_1_624 ();
 sg13g2_decap_8 FILLER_1_631 ();
 sg13g2_fill_2 FILLER_1_638 ();
 sg13g2_fill_1 FILLER_1_666 ();
 sg13g2_decap_8 FILLER_1_703 ();
 sg13g2_decap_8 FILLER_1_710 ();
 sg13g2_decap_8 FILLER_1_717 ();
 sg13g2_decap_8 FILLER_1_724 ();
 sg13g2_fill_2 FILLER_1_761 ();
 sg13g2_fill_1 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_794 ();
 sg13g2_decap_8 FILLER_1_801 ();
 sg13g2_fill_1 FILLER_1_808 ();
 sg13g2_fill_2 FILLER_1_845 ();
 sg13g2_fill_2 FILLER_1_851 ();
 sg13g2_fill_1 FILLER_1_853 ();
 sg13g2_fill_1 FILLER_1_880 ();
 sg13g2_fill_2 FILLER_1_891 ();
 sg13g2_fill_1 FILLER_1_893 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_fill_2 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_4 FILLER_1_994 ();
 sg13g2_fill_2 FILLER_1_998 ();
 sg13g2_decap_8 FILLER_1_1030 ();
 sg13g2_fill_1 FILLER_1_1037 ();
 sg13g2_decap_4 FILLER_1_1046 ();
 sg13g2_fill_1 FILLER_1_1050 ();
 sg13g2_fill_1 FILLER_1_1091 ();
 sg13g2_fill_2 FILLER_1_1154 ();
 sg13g2_fill_1 FILLER_1_1156 ();
 sg13g2_decap_4 FILLER_1_1213 ();
 sg13g2_decap_8 FILLER_1_1243 ();
 sg13g2_decap_8 FILLER_1_1250 ();
 sg13g2_fill_2 FILLER_1_1283 ();
 sg13g2_fill_1 FILLER_1_1285 ();
 sg13g2_fill_1 FILLER_1_1312 ();
 sg13g2_decap_8 FILLER_1_1339 ();
 sg13g2_fill_1 FILLER_1_1346 ();
 sg13g2_decap_8 FILLER_1_1403 ();
 sg13g2_decap_4 FILLER_1_1410 ();
 sg13g2_fill_2 FILLER_1_1444 ();
 sg13g2_fill_1 FILLER_1_1446 ();
 sg13g2_fill_2 FILLER_1_1539 ();
 sg13g2_fill_2 FILLER_1_1601 ();
 sg13g2_decap_8 FILLER_1_1639 ();
 sg13g2_decap_8 FILLER_1_1646 ();
 sg13g2_fill_2 FILLER_1_1653 ();
 sg13g2_decap_4 FILLER_1_1659 ();
 sg13g2_fill_2 FILLER_1_1689 ();
 sg13g2_decap_8 FILLER_1_1727 ();
 sg13g2_decap_8 FILLER_1_1734 ();
 sg13g2_decap_8 FILLER_1_1741 ();
 sg13g2_decap_8 FILLER_1_1748 ();
 sg13g2_decap_8 FILLER_1_1755 ();
 sg13g2_decap_8 FILLER_1_1762 ();
 sg13g2_decap_4 FILLER_1_1769 ();
 sg13g2_fill_1 FILLER_1_1773 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_fill_2 FILLER_2_40 ();
 sg13g2_fill_1 FILLER_2_42 ();
 sg13g2_decap_4 FILLER_2_73 ();
 sg13g2_fill_2 FILLER_2_113 ();
 sg13g2_decap_8 FILLER_2_145 ();
 sg13g2_decap_4 FILLER_2_152 ();
 sg13g2_fill_1 FILLER_2_156 ();
 sg13g2_fill_1 FILLER_2_161 ();
 sg13g2_fill_2 FILLER_2_192 ();
 sg13g2_decap_4 FILLER_2_224 ();
 sg13g2_fill_2 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_260 ();
 sg13g2_decap_8 FILLER_2_267 ();
 sg13g2_decap_4 FILLER_2_274 ();
 sg13g2_fill_1 FILLER_2_278 ();
 sg13g2_fill_2 FILLER_2_289 ();
 sg13g2_fill_2 FILLER_2_317 ();
 sg13g2_fill_1 FILLER_2_319 ();
 sg13g2_fill_1 FILLER_2_324 ();
 sg13g2_decap_4 FILLER_2_351 ();
 sg13g2_fill_1 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_decap_4 FILLER_2_429 ();
 sg13g2_fill_1 FILLER_2_433 ();
 sg13g2_decap_4 FILLER_2_500 ();
 sg13g2_decap_4 FILLER_2_508 ();
 sg13g2_fill_2 FILLER_2_564 ();
 sg13g2_decap_4 FILLER_2_576 ();
 sg13g2_decap_4 FILLER_2_606 ();
 sg13g2_fill_1 FILLER_2_610 ();
 sg13g2_fill_2 FILLER_2_641 ();
 sg13g2_decap_4 FILLER_2_669 ();
 sg13g2_fill_2 FILLER_2_673 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_4 FILLER_2_718 ();
 sg13g2_fill_1 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_fill_2 FILLER_2_849 ();
 sg13g2_fill_1 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_4 FILLER_2_928 ();
 sg13g2_fill_2 FILLER_2_932 ();
 sg13g2_fill_2 FILLER_2_1030 ();
 sg13g2_fill_1 FILLER_2_1108 ();
 sg13g2_decap_8 FILLER_2_1143 ();
 sg13g2_fill_2 FILLER_2_1150 ();
 sg13g2_fill_1 FILLER_2_1152 ();
 sg13g2_fill_2 FILLER_2_1193 ();
 sg13g2_decap_8 FILLER_2_1205 ();
 sg13g2_decap_8 FILLER_2_1212 ();
 sg13g2_fill_1 FILLER_2_1219 ();
 sg13g2_fill_1 FILLER_2_1357 ();
 sg13g2_fill_1 FILLER_2_1362 ();
 sg13g2_fill_2 FILLER_2_1373 ();
 sg13g2_fill_2 FILLER_2_1385 ();
 sg13g2_fill_2 FILLER_2_1391 ();
 sg13g2_decap_8 FILLER_2_1397 ();
 sg13g2_decap_8 FILLER_2_1404 ();
 sg13g2_decap_8 FILLER_2_1411 ();
 sg13g2_decap_4 FILLER_2_1418 ();
 sg13g2_decap_4 FILLER_2_1436 ();
 sg13g2_fill_1 FILLER_2_1440 ();
 sg13g2_fill_1 FILLER_2_1549 ();
 sg13g2_decap_8 FILLER_2_1573 ();
 sg13g2_fill_1 FILLER_2_1580 ();
 sg13g2_fill_2 FILLER_2_1595 ();
 sg13g2_fill_1 FILLER_2_1597 ();
 sg13g2_fill_1 FILLER_2_1616 ();
 sg13g2_fill_2 FILLER_2_1699 ();
 sg13g2_decap_8 FILLER_2_1715 ();
 sg13g2_decap_8 FILLER_2_1722 ();
 sg13g2_decap_8 FILLER_2_1729 ();
 sg13g2_decap_8 FILLER_2_1736 ();
 sg13g2_decap_8 FILLER_2_1743 ();
 sg13g2_decap_8 FILLER_2_1750 ();
 sg13g2_decap_8 FILLER_2_1757 ();
 sg13g2_decap_8 FILLER_2_1764 ();
 sg13g2_fill_2 FILLER_2_1771 ();
 sg13g2_fill_1 FILLER_2_1773 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_12 ();
 sg13g2_fill_2 FILLER_3_43 ();
 sg13g2_fill_1 FILLER_3_45 ();
 sg13g2_decap_4 FILLER_3_63 ();
 sg13g2_fill_1 FILLER_3_77 ();
 sg13g2_decap_4 FILLER_3_82 ();
 sg13g2_fill_2 FILLER_3_86 ();
 sg13g2_fill_1 FILLER_3_98 ();
 sg13g2_fill_2 FILLER_3_125 ();
 sg13g2_fill_2 FILLER_3_131 ();
 sg13g2_fill_2 FILLER_3_159 ();
 sg13g2_fill_2 FILLER_3_191 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_4 FILLER_3_228 ();
 sg13g2_fill_2 FILLER_3_232 ();
 sg13g2_fill_1 FILLER_3_264 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_fill_1 FILLER_3_386 ();
 sg13g2_fill_1 FILLER_3_391 ();
 sg13g2_fill_1 FILLER_3_402 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_fill_2 FILLER_3_485 ();
 sg13g2_fill_2 FILLER_3_517 ();
 sg13g2_decap_8 FILLER_3_529 ();
 sg13g2_decap_8 FILLER_3_536 ();
 sg13g2_decap_4 FILLER_3_543 ();
 sg13g2_fill_1 FILLER_3_547 ();
 sg13g2_decap_8 FILLER_3_603 ();
 sg13g2_fill_2 FILLER_3_610 ();
 sg13g2_fill_1 FILLER_3_612 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_709 ();
 sg13g2_decap_8 FILLER_3_716 ();
 sg13g2_decap_8 FILLER_3_723 ();
 sg13g2_fill_1 FILLER_3_775 ();
 sg13g2_fill_2 FILLER_3_786 ();
 sg13g2_fill_1 FILLER_3_792 ();
 sg13g2_fill_1 FILLER_3_819 ();
 sg13g2_decap_4 FILLER_3_876 ();
 sg13g2_decap_8 FILLER_3_890 ();
 sg13g2_fill_2 FILLER_3_901 ();
 sg13g2_fill_1 FILLER_3_903 ();
 sg13g2_decap_8 FILLER_3_908 ();
 sg13g2_decap_8 FILLER_3_928 ();
 sg13g2_fill_2 FILLER_3_935 ();
 sg13g2_fill_1 FILLER_3_937 ();
 sg13g2_fill_1 FILLER_3_948 ();
 sg13g2_fill_1 FILLER_3_975 ();
 sg13g2_fill_2 FILLER_3_986 ();
 sg13g2_fill_1 FILLER_3_1009 ();
 sg13g2_fill_2 FILLER_3_1020 ();
 sg13g2_fill_2 FILLER_3_1026 ();
 sg13g2_fill_1 FILLER_3_1028 ();
 sg13g2_decap_4 FILLER_3_1064 ();
 sg13g2_fill_1 FILLER_3_1068 ();
 sg13g2_fill_1 FILLER_3_1073 ();
 sg13g2_fill_2 FILLER_3_1095 ();
 sg13g2_fill_1 FILLER_3_1097 ();
 sg13g2_fill_2 FILLER_3_1163 ();
 sg13g2_fill_1 FILLER_3_1169 ();
 sg13g2_decap_8 FILLER_3_1174 ();
 sg13g2_fill_2 FILLER_3_1195 ();
 sg13g2_fill_1 FILLER_3_1197 ();
 sg13g2_decap_8 FILLER_3_1202 ();
 sg13g2_fill_2 FILLER_3_1209 ();
 sg13g2_decap_8 FILLER_3_1221 ();
 sg13g2_decap_4 FILLER_3_1228 ();
 sg13g2_fill_1 FILLER_3_1232 ();
 sg13g2_decap_8 FILLER_3_1237 ();
 sg13g2_decap_4 FILLER_3_1244 ();
 sg13g2_fill_2 FILLER_3_1248 ();
 sg13g2_fill_2 FILLER_3_1254 ();
 sg13g2_fill_2 FILLER_3_1308 ();
 sg13g2_fill_1 FILLER_3_1310 ();
 sg13g2_fill_2 FILLER_3_1383 ();
 sg13g2_decap_8 FILLER_3_1389 ();
 sg13g2_decap_8 FILLER_3_1396 ();
 sg13g2_decap_8 FILLER_3_1403 ();
 sg13g2_decap_8 FILLER_3_1410 ();
 sg13g2_fill_2 FILLER_3_1417 ();
 sg13g2_fill_1 FILLER_3_1445 ();
 sg13g2_fill_1 FILLER_3_1482 ();
 sg13g2_fill_2 FILLER_3_1513 ();
 sg13g2_fill_1 FILLER_3_1515 ();
 sg13g2_decap_4 FILLER_3_1524 ();
 sg13g2_fill_2 FILLER_3_1528 ();
 sg13g2_decap_8 FILLER_3_1584 ();
 sg13g2_decap_8 FILLER_3_1591 ();
 sg13g2_fill_2 FILLER_3_1598 ();
 sg13g2_fill_1 FILLER_3_1600 ();
 sg13g2_decap_8 FILLER_3_1647 ();
 sg13g2_decap_4 FILLER_3_1654 ();
 sg13g2_fill_1 FILLER_3_1658 ();
 sg13g2_decap_4 FILLER_3_1699 ();
 sg13g2_fill_2 FILLER_3_1703 ();
 sg13g2_decap_8 FILLER_3_1735 ();
 sg13g2_decap_8 FILLER_3_1742 ();
 sg13g2_decap_8 FILLER_3_1749 ();
 sg13g2_decap_8 FILLER_3_1756 ();
 sg13g2_decap_8 FILLER_3_1763 ();
 sg13g2_decap_4 FILLER_3_1770 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_24 ();
 sg13g2_fill_1 FILLER_4_26 ();
 sg13g2_decap_4 FILLER_4_37 ();
 sg13g2_fill_2 FILLER_4_41 ();
 sg13g2_fill_2 FILLER_4_53 ();
 sg13g2_fill_1 FILLER_4_55 ();
 sg13g2_fill_2 FILLER_4_113 ();
 sg13g2_fill_2 FILLER_4_125 ();
 sg13g2_decap_8 FILLER_4_148 ();
 sg13g2_decap_8 FILLER_4_155 ();
 sg13g2_fill_2 FILLER_4_172 ();
 sg13g2_fill_1 FILLER_4_174 ();
 sg13g2_decap_4 FILLER_4_221 ();
 sg13g2_fill_2 FILLER_4_225 ();
 sg13g2_fill_1 FILLER_4_247 ();
 sg13g2_fill_2 FILLER_4_283 ();
 sg13g2_fill_2 FILLER_4_295 ();
 sg13g2_fill_1 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_fill_2 FILLER_4_326 ();
 sg13g2_fill_1 FILLER_4_328 ();
 sg13g2_fill_1 FILLER_4_343 ();
 sg13g2_fill_2 FILLER_4_368 ();
 sg13g2_fill_1 FILLER_4_370 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_fill_1 FILLER_4_388 ();
 sg13g2_fill_1 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_404 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_2 FILLER_4_439 ();
 sg13g2_fill_1 FILLER_4_441 ();
 sg13g2_fill_1 FILLER_4_446 ();
 sg13g2_fill_2 FILLER_4_468 ();
 sg13g2_fill_2 FILLER_4_474 ();
 sg13g2_fill_2 FILLER_4_486 ();
 sg13g2_fill_1 FILLER_4_488 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_fill_2 FILLER_4_553 ();
 sg13g2_fill_1 FILLER_4_555 ();
 sg13g2_fill_1 FILLER_4_596 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_fill_2 FILLER_4_630 ();
 sg13g2_fill_2 FILLER_4_662 ();
 sg13g2_decap_8 FILLER_4_759 ();
 sg13g2_decap_8 FILLER_4_766 ();
 sg13g2_fill_2 FILLER_4_773 ();
 sg13g2_fill_2 FILLER_4_783 ();
 sg13g2_decap_8 FILLER_4_815 ();
 sg13g2_decap_4 FILLER_4_822 ();
 sg13g2_fill_2 FILLER_4_840 ();
 sg13g2_fill_2 FILLER_4_852 ();
 sg13g2_fill_2 FILLER_4_858 ();
 sg13g2_fill_1 FILLER_4_860 ();
 sg13g2_fill_2 FILLER_4_865 ();
 sg13g2_fill_1 FILLER_4_867 ();
 sg13g2_decap_8 FILLER_4_889 ();
 sg13g2_decap_8 FILLER_4_896 ();
 sg13g2_decap_8 FILLER_4_903 ();
 sg13g2_decap_8 FILLER_4_910 ();
 sg13g2_decap_8 FILLER_4_917 ();
 sg13g2_decap_8 FILLER_4_924 ();
 sg13g2_decap_8 FILLER_4_977 ();
 sg13g2_decap_4 FILLER_4_984 ();
 sg13g2_fill_1 FILLER_4_988 ();
 sg13g2_decap_4 FILLER_4_1029 ();
 sg13g2_decap_8 FILLER_4_1059 ();
 sg13g2_decap_8 FILLER_4_1066 ();
 sg13g2_decap_8 FILLER_4_1073 ();
 sg13g2_decap_8 FILLER_4_1080 ();
 sg13g2_fill_2 FILLER_4_1087 ();
 sg13g2_fill_1 FILLER_4_1089 ();
 sg13g2_decap_8 FILLER_4_1136 ();
 sg13g2_decap_8 FILLER_4_1143 ();
 sg13g2_fill_2 FILLER_4_1150 ();
 sg13g2_fill_1 FILLER_4_1152 ();
 sg13g2_fill_2 FILLER_4_1215 ();
 sg13g2_decap_8 FILLER_4_1243 ();
 sg13g2_decap_8 FILLER_4_1250 ();
 sg13g2_fill_1 FILLER_4_1257 ();
 sg13g2_fill_2 FILLER_4_1262 ();
 sg13g2_fill_1 FILLER_4_1264 ();
 sg13g2_fill_2 FILLER_4_1275 ();
 sg13g2_fill_2 FILLER_4_1313 ();
 sg13g2_fill_1 FILLER_4_1315 ();
 sg13g2_fill_2 FILLER_4_1330 ();
 sg13g2_fill_1 FILLER_4_1332 ();
 sg13g2_fill_2 FILLER_4_1369 ();
 sg13g2_fill_1 FILLER_4_1371 ();
 sg13g2_decap_8 FILLER_4_1398 ();
 sg13g2_fill_1 FILLER_4_1405 ();
 sg13g2_decap_4 FILLER_4_1432 ();
 sg13g2_decap_8 FILLER_4_1446 ();
 sg13g2_fill_2 FILLER_4_1463 ();
 sg13g2_fill_1 FILLER_4_1465 ();
 sg13g2_fill_2 FILLER_4_1506 ();
 sg13g2_fill_1 FILLER_4_1508 ();
 sg13g2_fill_2 FILLER_4_1535 ();
 sg13g2_decap_8 FILLER_4_1577 ();
 sg13g2_decap_8 FILLER_4_1584 ();
 sg13g2_decap_4 FILLER_4_1591 ();
 sg13g2_fill_2 FILLER_4_1595 ();
 sg13g2_fill_1 FILLER_4_1654 ();
 sg13g2_fill_2 FILLER_4_1679 ();
 sg13g2_fill_1 FILLER_4_1681 ();
 sg13g2_fill_2 FILLER_4_1703 ();
 sg13g2_decap_8 FILLER_4_1731 ();
 sg13g2_decap_8 FILLER_4_1738 ();
 sg13g2_decap_8 FILLER_4_1745 ();
 sg13g2_decap_8 FILLER_4_1752 ();
 sg13g2_decap_8 FILLER_4_1759 ();
 sg13g2_decap_8 FILLER_4_1766 ();
 sg13g2_fill_1 FILLER_4_1773 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_4 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_25 ();
 sg13g2_fill_1 FILLER_5_30 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_fill_2 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_86 ();
 sg13g2_fill_1 FILLER_5_117 ();
 sg13g2_decap_8 FILLER_5_139 ();
 sg13g2_fill_1 FILLER_5_146 ();
 sg13g2_decap_8 FILLER_5_157 ();
 sg13g2_decap_8 FILLER_5_164 ();
 sg13g2_decap_8 FILLER_5_171 ();
 sg13g2_decap_8 FILLER_5_178 ();
 sg13g2_decap_8 FILLER_5_225 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_fill_1 FILLER_5_239 ();
 sg13g2_decap_8 FILLER_5_243 ();
 sg13g2_decap_8 FILLER_5_250 ();
 sg13g2_decap_8 FILLER_5_257 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_decap_4 FILLER_5_271 ();
 sg13g2_fill_2 FILLER_5_275 ();
 sg13g2_fill_1 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_4 FILLER_5_355 ();
 sg13g2_fill_2 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_5_430 ();
 sg13g2_decap_8 FILLER_5_437 ();
 sg13g2_decap_8 FILLER_5_444 ();
 sg13g2_decap_8 FILLER_5_451 ();
 sg13g2_decap_8 FILLER_5_458 ();
 sg13g2_decap_8 FILLER_5_465 ();
 sg13g2_fill_1 FILLER_5_482 ();
 sg13g2_decap_8 FILLER_5_491 ();
 sg13g2_fill_1 FILLER_5_498 ();
 sg13g2_fill_2 FILLER_5_503 ();
 sg13g2_fill_2 FILLER_5_515 ();
 sg13g2_fill_1 FILLER_5_517 ();
 sg13g2_decap_4 FILLER_5_544 ();
 sg13g2_fill_2 FILLER_5_548 ();
 sg13g2_fill_2 FILLER_5_575 ();
 sg13g2_fill_1 FILLER_5_603 ();
 sg13g2_decap_8 FILLER_5_608 ();
 sg13g2_decap_8 FILLER_5_615 ();
 sg13g2_decap_8 FILLER_5_622 ();
 sg13g2_fill_1 FILLER_5_633 ();
 sg13g2_decap_4 FILLER_5_654 ();
 sg13g2_decap_8 FILLER_5_668 ();
 sg13g2_fill_2 FILLER_5_675 ();
 sg13g2_fill_1 FILLER_5_677 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_4 FILLER_5_728 ();
 sg13g2_fill_2 FILLER_5_772 ();
 sg13g2_decap_4 FILLER_5_807 ();
 sg13g2_fill_1 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_fill_1 FILLER_5_865 ();
 sg13g2_decap_8 FILLER_5_921 ();
 sg13g2_decap_8 FILLER_5_928 ();
 sg13g2_fill_2 FILLER_5_935 ();
 sg13g2_decap_4 FILLER_5_941 ();
 sg13g2_fill_2 FILLER_5_945 ();
 sg13g2_fill_1 FILLER_5_982 ();
 sg13g2_fill_1 FILLER_5_1009 ();
 sg13g2_decap_8 FILLER_5_1014 ();
 sg13g2_decap_4 FILLER_5_1021 ();
 sg13g2_fill_1 FILLER_5_1025 ();
 sg13g2_fill_1 FILLER_5_1036 ();
 sg13g2_decap_8 FILLER_5_1041 ();
 sg13g2_decap_8 FILLER_5_1048 ();
 sg13g2_decap_4 FILLER_5_1055 ();
 sg13g2_fill_1 FILLER_5_1059 ();
 sg13g2_decap_8 FILLER_5_1096 ();
 sg13g2_decap_4 FILLER_5_1103 ();
 sg13g2_decap_8 FILLER_5_1111 ();
 sg13g2_decap_8 FILLER_5_1118 ();
 sg13g2_decap_8 FILLER_5_1125 ();
 sg13g2_decap_8 FILLER_5_1132 ();
 sg13g2_decap_8 FILLER_5_1139 ();
 sg13g2_decap_8 FILLER_5_1146 ();
 sg13g2_decap_8 FILLER_5_1167 ();
 sg13g2_decap_8 FILLER_5_1174 ();
 sg13g2_decap_8 FILLER_5_1181 ();
 sg13g2_decap_8 FILLER_5_1188 ();
 sg13g2_fill_2 FILLER_5_1195 ();
 sg13g2_fill_1 FILLER_5_1197 ();
 sg13g2_decap_8 FILLER_5_1238 ();
 sg13g2_decap_8 FILLER_5_1245 ();
 sg13g2_decap_4 FILLER_5_1252 ();
 sg13g2_fill_1 FILLER_5_1256 ();
 sg13g2_fill_1 FILLER_5_1308 ();
 sg13g2_decap_8 FILLER_5_1313 ();
 sg13g2_fill_1 FILLER_5_1320 ();
 sg13g2_decap_4 FILLER_5_1342 ();
 sg13g2_fill_2 FILLER_5_1346 ();
 sg13g2_decap_4 FILLER_5_1352 ();
 sg13g2_fill_1 FILLER_5_1356 ();
 sg13g2_decap_8 FILLER_5_1378 ();
 sg13g2_decap_8 FILLER_5_1385 ();
 sg13g2_decap_8 FILLER_5_1392 ();
 sg13g2_fill_2 FILLER_5_1399 ();
 sg13g2_fill_1 FILLER_5_1401 ();
 sg13g2_decap_4 FILLER_5_1406 ();
 sg13g2_fill_1 FILLER_5_1410 ();
 sg13g2_decap_8 FILLER_5_1425 ();
 sg13g2_decap_8 FILLER_5_1458 ();
 sg13g2_decap_8 FILLER_5_1465 ();
 sg13g2_decap_4 FILLER_5_1472 ();
 sg13g2_decap_4 FILLER_5_1480 ();
 sg13g2_fill_2 FILLER_5_1484 ();
 sg13g2_decap_8 FILLER_5_1509 ();
 sg13g2_decap_8 FILLER_5_1516 ();
 sg13g2_decap_8 FILLER_5_1523 ();
 sg13g2_decap_8 FILLER_5_1530 ();
 sg13g2_decap_8 FILLER_5_1537 ();
 sg13g2_decap_4 FILLER_5_1544 ();
 sg13g2_fill_1 FILLER_5_1548 ();
 sg13g2_fill_1 FILLER_5_1552 ();
 sg13g2_decap_8 FILLER_5_1589 ();
 sg13g2_decap_8 FILLER_5_1596 ();
 sg13g2_decap_8 FILLER_5_1603 ();
 sg13g2_decap_8 FILLER_5_1654 ();
 sg13g2_fill_1 FILLER_5_1661 ();
 sg13g2_decap_8 FILLER_5_1687 ();
 sg13g2_fill_2 FILLER_5_1694 ();
 sg13g2_fill_2 FILLER_5_1706 ();
 sg13g2_fill_1 FILLER_5_1708 ();
 sg13g2_decap_4 FILLER_5_1713 ();
 sg13g2_fill_2 FILLER_5_1717 ();
 sg13g2_fill_1 FILLER_5_1739 ();
 sg13g2_decap_8 FILLER_5_1766 ();
 sg13g2_fill_1 FILLER_5_1773 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_45 ();
 sg13g2_fill_1 FILLER_6_79 ();
 sg13g2_decap_4 FILLER_6_90 ();
 sg13g2_fill_1 FILLER_6_94 ();
 sg13g2_fill_2 FILLER_6_99 ();
 sg13g2_fill_1 FILLER_6_101 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_178 ();
 sg13g2_fill_2 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_187 ();
 sg13g2_fill_2 FILLER_6_192 ();
 sg13g2_fill_1 FILLER_6_194 ();
 sg13g2_fill_2 FILLER_6_205 ();
 sg13g2_fill_1 FILLER_6_207 ();
 sg13g2_decap_4 FILLER_6_212 ();
 sg13g2_fill_1 FILLER_6_216 ();
 sg13g2_fill_1 FILLER_6_227 ();
 sg13g2_decap_4 FILLER_6_232 ();
 sg13g2_decap_4 FILLER_6_261 ();
 sg13g2_fill_1 FILLER_6_265 ();
 sg13g2_decap_8 FILLER_6_292 ();
 sg13g2_fill_2 FILLER_6_299 ();
 sg13g2_fill_1 FILLER_6_301 ();
 sg13g2_fill_2 FILLER_6_328 ();
 sg13g2_fill_1 FILLER_6_330 ();
 sg13g2_decap_4 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_fill_2 FILLER_6_389 ();
 sg13g2_fill_2 FILLER_6_416 ();
 sg13g2_fill_1 FILLER_6_418 ();
 sg13g2_decap_8 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_6_436 ();
 sg13g2_decap_8 FILLER_6_443 ();
 sg13g2_decap_4 FILLER_6_450 ();
 sg13g2_fill_2 FILLER_6_454 ();
 sg13g2_fill_1 FILLER_6_460 ();
 sg13g2_fill_1 FILLER_6_471 ();
 sg13g2_fill_1 FILLER_6_482 ();
 sg13g2_fill_1 FILLER_6_530 ();
 sg13g2_decap_8 FILLER_6_535 ();
 sg13g2_decap_8 FILLER_6_542 ();
 sg13g2_decap_8 FILLER_6_549 ();
 sg13g2_fill_2 FILLER_6_556 ();
 sg13g2_fill_1 FILLER_6_558 ();
 sg13g2_fill_2 FILLER_6_572 ();
 sg13g2_decap_4 FILLER_6_599 ();
 sg13g2_fill_2 FILLER_6_603 ();
 sg13g2_fill_2 FILLER_6_609 ();
 sg13g2_fill_1 FILLER_6_611 ();
 sg13g2_fill_2 FILLER_6_648 ();
 sg13g2_fill_1 FILLER_6_650 ();
 sg13g2_fill_2 FILLER_6_655 ();
 sg13g2_fill_2 FILLER_6_667 ();
 sg13g2_fill_1 FILLER_6_669 ();
 sg13g2_fill_2 FILLER_6_691 ();
 sg13g2_fill_1 FILLER_6_693 ();
 sg13g2_fill_2 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_710 ();
 sg13g2_decap_4 FILLER_6_717 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_4 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_810 ();
 sg13g2_fill_2 FILLER_6_817 ();
 sg13g2_fill_1 FILLER_6_819 ();
 sg13g2_decap_4 FILLER_6_882 ();
 sg13g2_decap_8 FILLER_6_922 ();
 sg13g2_decap_8 FILLER_6_929 ();
 sg13g2_decap_8 FILLER_6_936 ();
 sg13g2_fill_1 FILLER_6_943 ();
 sg13g2_fill_1 FILLER_6_970 ();
 sg13g2_fill_1 FILLER_6_981 ();
 sg13g2_fill_1 FILLER_6_992 ();
 sg13g2_fill_1 FILLER_6_997 ();
 sg13g2_decap_8 FILLER_6_1008 ();
 sg13g2_decap_4 FILLER_6_1015 ();
 sg13g2_fill_1 FILLER_6_1019 ();
 sg13g2_decap_8 FILLER_6_1028 ();
 sg13g2_decap_8 FILLER_6_1035 ();
 sg13g2_decap_8 FILLER_6_1042 ();
 sg13g2_decap_8 FILLER_6_1049 ();
 sg13g2_fill_1 FILLER_6_1082 ();
 sg13g2_fill_2 FILLER_6_1109 ();
 sg13g2_decap_8 FILLER_6_1121 ();
 sg13g2_decap_8 FILLER_6_1128 ();
 sg13g2_decap_8 FILLER_6_1135 ();
 sg13g2_decap_8 FILLER_6_1142 ();
 sg13g2_decap_8 FILLER_6_1149 ();
 sg13g2_fill_2 FILLER_6_1156 ();
 sg13g2_fill_1 FILLER_6_1158 ();
 sg13g2_fill_1 FILLER_6_1224 ();
 sg13g2_fill_2 FILLER_6_1229 ();
 sg13g2_fill_1 FILLER_6_1231 ();
 sg13g2_decap_8 FILLER_6_1236 ();
 sg13g2_decap_8 FILLER_6_1243 ();
 sg13g2_decap_8 FILLER_6_1250 ();
 sg13g2_decap_8 FILLER_6_1257 ();
 sg13g2_decap_4 FILLER_6_1264 ();
 sg13g2_fill_2 FILLER_6_1268 ();
 sg13g2_decap_8 FILLER_6_1304 ();
 sg13g2_decap_8 FILLER_6_1311 ();
 sg13g2_decap_8 FILLER_6_1318 ();
 sg13g2_decap_8 FILLER_6_1325 ();
 sg13g2_decap_8 FILLER_6_1368 ();
 sg13g2_fill_2 FILLER_6_1375 ();
 sg13g2_decap_8 FILLER_6_1381 ();
 sg13g2_decap_8 FILLER_6_1388 ();
 sg13g2_decap_8 FILLER_6_1445 ();
 sg13g2_fill_2 FILLER_6_1452 ();
 sg13g2_decap_8 FILLER_6_1464 ();
 sg13g2_decap_8 FILLER_6_1471 ();
 sg13g2_decap_8 FILLER_6_1478 ();
 sg13g2_fill_2 FILLER_6_1493 ();
 sg13g2_fill_1 FILLER_6_1495 ();
 sg13g2_fill_2 FILLER_6_1517 ();
 sg13g2_decap_4 FILLER_6_1523 ();
 sg13g2_decap_8 FILLER_6_1537 ();
 sg13g2_fill_1 FILLER_6_1544 ();
 sg13g2_decap_8 FILLER_6_1584 ();
 sg13g2_decap_8 FILLER_6_1591 ();
 sg13g2_decap_4 FILLER_6_1598 ();
 sg13g2_decap_4 FILLER_6_1623 ();
 sg13g2_fill_2 FILLER_6_1627 ();
 sg13g2_decap_8 FILLER_6_1643 ();
 sg13g2_decap_8 FILLER_6_1650 ();
 sg13g2_decap_8 FILLER_6_1657 ();
 sg13g2_fill_2 FILLER_6_1664 ();
 sg13g2_fill_1 FILLER_6_1738 ();
 sg13g2_decap_8 FILLER_6_1765 ();
 sg13g2_fill_2 FILLER_6_1772 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_44 ();
 sg13g2_fill_1 FILLER_7_55 ();
 sg13g2_decap_8 FILLER_7_78 ();
 sg13g2_decap_8 FILLER_7_85 ();
 sg13g2_decap_4 FILLER_7_92 ();
 sg13g2_fill_2 FILLER_7_96 ();
 sg13g2_fill_2 FILLER_7_107 ();
 sg13g2_decap_4 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_247 ();
 sg13g2_fill_1 FILLER_7_280 ();
 sg13g2_decap_4 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_338 ();
 sg13g2_fill_2 FILLER_7_345 ();
 sg13g2_fill_1 FILLER_7_347 ();
 sg13g2_decap_4 FILLER_7_378 ();
 sg13g2_fill_1 FILLER_7_382 ();
 sg13g2_decap_4 FILLER_7_396 ();
 sg13g2_fill_2 FILLER_7_400 ();
 sg13g2_decap_4 FILLER_7_436 ();
 sg13g2_fill_1 FILLER_7_454 ();
 sg13g2_fill_1 FILLER_7_481 ();
 sg13g2_fill_1 FILLER_7_508 ();
 sg13g2_decap_4 FILLER_7_530 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_fill_1 FILLER_7_581 ();
 sg13g2_fill_1 FILLER_7_594 ();
 sg13g2_fill_2 FILLER_7_641 ();
 sg13g2_fill_1 FILLER_7_643 ();
 sg13g2_fill_2 FILLER_7_696 ();
 sg13g2_fill_1 FILLER_7_698 ();
 sg13g2_decap_4 FILLER_7_703 ();
 sg13g2_fill_1 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_4 FILLER_7_728 ();
 sg13g2_fill_2 FILLER_7_732 ();
 sg13g2_fill_2 FILLER_7_764 ();
 sg13g2_fill_1 FILLER_7_766 ();
 sg13g2_fill_1 FILLER_7_777 ();
 sg13g2_fill_1 FILLER_7_799 ();
 sg13g2_fill_1 FILLER_7_826 ();
 sg13g2_fill_1 FILLER_7_853 ();
 sg13g2_fill_1 FILLER_7_858 ();
 sg13g2_fill_2 FILLER_7_869 ();
 sg13g2_decap_4 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_889 ();
 sg13g2_fill_2 FILLER_7_900 ();
 sg13g2_fill_1 FILLER_7_902 ();
 sg13g2_decap_8 FILLER_7_907 ();
 sg13g2_decap_8 FILLER_7_914 ();
 sg13g2_decap_8 FILLER_7_921 ();
 sg13g2_decap_8 FILLER_7_928 ();
 sg13g2_fill_1 FILLER_7_935 ();
 sg13g2_decap_4 FILLER_7_972 ();
 sg13g2_fill_2 FILLER_7_1002 ();
 sg13g2_fill_2 FILLER_7_1035 ();
 sg13g2_fill_1 FILLER_7_1067 ();
 sg13g2_fill_1 FILLER_7_1072 ();
 sg13g2_fill_1 FILLER_7_1083 ();
 sg13g2_fill_1 FILLER_7_1088 ();
 sg13g2_fill_2 FILLER_7_1093 ();
 sg13g2_fill_2 FILLER_7_1173 ();
 sg13g2_decap_8 FILLER_7_1248 ();
 sg13g2_decap_8 FILLER_7_1255 ();
 sg13g2_fill_2 FILLER_7_1262 ();
 sg13g2_fill_1 FILLER_7_1264 ();
 sg13g2_decap_8 FILLER_7_1295 ();
 sg13g2_fill_2 FILLER_7_1302 ();
 sg13g2_fill_2 FILLER_7_1358 ();
 sg13g2_decap_8 FILLER_7_1396 ();
 sg13g2_fill_1 FILLER_7_1403 ();
 sg13g2_decap_4 FILLER_7_1491 ();
 sg13g2_decap_4 FILLER_7_1505 ();
 sg13g2_fill_2 FILLER_7_1535 ();
 sg13g2_fill_1 FILLER_7_1537 ();
 sg13g2_fill_2 FILLER_7_1564 ();
 sg13g2_fill_1 FILLER_7_1566 ();
 sg13g2_decap_8 FILLER_7_1593 ();
 sg13g2_fill_2 FILLER_7_1600 ();
 sg13g2_fill_1 FILLER_7_1602 ();
 sg13g2_fill_2 FILLER_7_1665 ();
 sg13g2_fill_1 FILLER_7_1667 ();
 sg13g2_decap_8 FILLER_7_1678 ();
 sg13g2_fill_2 FILLER_7_1689 ();
 sg13g2_fill_1 FILLER_7_1695 ();
 sg13g2_fill_2 FILLER_7_1706 ();
 sg13g2_fill_2 FILLER_7_1738 ();
 sg13g2_fill_1 FILLER_7_1740 ();
 sg13g2_fill_1 FILLER_7_1749 ();
 sg13g2_decap_8 FILLER_7_1754 ();
 sg13g2_decap_8 FILLER_7_1761 ();
 sg13g2_decap_4 FILLER_7_1768 ();
 sg13g2_fill_2 FILLER_7_1772 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_fill_1 FILLER_8_52 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_4 FILLER_8_84 ();
 sg13g2_fill_1 FILLER_8_118 ();
 sg13g2_fill_1 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_158 ();
 sg13g2_fill_1 FILLER_8_163 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_fill_1 FILLER_8_175 ();
 sg13g2_fill_2 FILLER_8_186 ();
 sg13g2_decap_4 FILLER_8_209 ();
 sg13g2_fill_2 FILLER_8_277 ();
 sg13g2_fill_1 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_325 ();
 sg13g2_fill_1 FILLER_8_332 ();
 sg13g2_fill_2 FILLER_8_354 ();
 sg13g2_fill_1 FILLER_8_356 ();
 sg13g2_fill_1 FILLER_8_367 ();
 sg13g2_fill_2 FILLER_8_394 ();
 sg13g2_fill_1 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_fill_1 FILLER_8_430 ();
 sg13g2_decap_4 FILLER_8_492 ();
 sg13g2_fill_1 FILLER_8_500 ();
 sg13g2_fill_1 FILLER_8_505 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_4 FILLER_8_543 ();
 sg13g2_fill_2 FILLER_8_547 ();
 sg13g2_fill_1 FILLER_8_584 ();
 sg13g2_fill_1 FILLER_8_591 ();
 sg13g2_fill_2 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_722 ();
 sg13g2_decap_8 FILLER_8_729 ();
 sg13g2_decap_4 FILLER_8_736 ();
 sg13g2_fill_2 FILLER_8_740 ();
 sg13g2_fill_1 FILLER_8_746 ();
 sg13g2_fill_1 FILLER_8_757 ();
 sg13g2_fill_2 FILLER_8_768 ();
 sg13g2_fill_1 FILLER_8_774 ();
 sg13g2_fill_2 FILLER_8_801 ();
 sg13g2_fill_2 FILLER_8_813 ();
 sg13g2_fill_2 FILLER_8_836 ();
 sg13g2_decap_8 FILLER_8_885 ();
 sg13g2_decap_8 FILLER_8_892 ();
 sg13g2_decap_4 FILLER_8_899 ();
 sg13g2_fill_1 FILLER_8_920 ();
 sg13g2_decap_8 FILLER_8_934 ();
 sg13g2_fill_1 FILLER_8_941 ();
 sg13g2_fill_2 FILLER_8_982 ();
 sg13g2_fill_1 FILLER_8_984 ();
 sg13g2_fill_2 FILLER_8_999 ();
 sg13g2_fill_1 FILLER_8_1001 ();
 sg13g2_decap_4 FILLER_8_1016 ();
 sg13g2_fill_2 FILLER_8_1020 ();
 sg13g2_decap_4 FILLER_8_1026 ();
 sg13g2_fill_2 FILLER_8_1030 ();
 sg13g2_fill_1 FILLER_8_1042 ();
 sg13g2_fill_2 FILLER_8_1056 ();
 sg13g2_decap_4 FILLER_8_1066 ();
 sg13g2_fill_2 FILLER_8_1070 ();
 sg13g2_fill_1 FILLER_8_1082 ();
 sg13g2_fill_2 FILLER_8_1086 ();
 sg13g2_fill_1 FILLER_8_1101 ();
 sg13g2_fill_2 FILLER_8_1109 ();
 sg13g2_fill_1 FILLER_8_1111 ();
 sg13g2_fill_1 FILLER_8_1142 ();
 sg13g2_fill_1 FILLER_8_1169 ();
 sg13g2_decap_4 FILLER_8_1180 ();
 sg13g2_fill_2 FILLER_8_1184 ();
 sg13g2_fill_1 FILLER_8_1190 ();
 sg13g2_decap_8 FILLER_8_1243 ();
 sg13g2_fill_2 FILLER_8_1258 ();
 sg13g2_fill_1 FILLER_8_1260 ();
 sg13g2_fill_1 FILLER_8_1307 ();
 sg13g2_decap_8 FILLER_8_1354 ();
 sg13g2_decap_4 FILLER_8_1361 ();
 sg13g2_decap_8 FILLER_8_1401 ();
 sg13g2_decap_8 FILLER_8_1408 ();
 sg13g2_decap_4 FILLER_8_1415 ();
 sg13g2_fill_1 FILLER_8_1459 ();
 sg13g2_fill_2 FILLER_8_1494 ();
 sg13g2_fill_1 FILLER_8_1496 ();
 sg13g2_decap_4 FILLER_8_1593 ();
 sg13g2_fill_2 FILLER_8_1597 ();
 sg13g2_fill_1 FILLER_8_1635 ();
 sg13g2_fill_2 FILLER_8_1644 ();
 sg13g2_fill_2 FILLER_8_1650 ();
 sg13g2_fill_2 FILLER_8_1662 ();
 sg13g2_fill_2 FILLER_8_1668 ();
 sg13g2_fill_2 FILLER_8_1675 ();
 sg13g2_fill_1 FILLER_8_1677 ();
 sg13g2_fill_2 FILLER_8_1704 ();
 sg13g2_fill_1 FILLER_8_1706 ();
 sg13g2_fill_2 FILLER_8_1733 ();
 sg13g2_decap_8 FILLER_8_1739 ();
 sg13g2_decap_8 FILLER_8_1746 ();
 sg13g2_decap_8 FILLER_8_1753 ();
 sg13g2_decap_8 FILLER_8_1760 ();
 sg13g2_decap_8 FILLER_8_1767 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_11 ();
 sg13g2_fill_1 FILLER_9_64 ();
 sg13g2_decap_4 FILLER_9_79 ();
 sg13g2_fill_1 FILLER_9_129 ();
 sg13g2_decap_8 FILLER_9_134 ();
 sg13g2_fill_1 FILLER_9_141 ();
 sg13g2_decap_8 FILLER_9_163 ();
 sg13g2_decap_4 FILLER_9_170 ();
 sg13g2_fill_2 FILLER_9_174 ();
 sg13g2_fill_1 FILLER_9_180 ();
 sg13g2_fill_2 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_235 ();
 sg13g2_fill_2 FILLER_9_246 ();
 sg13g2_fill_2 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_fill_2 FILLER_9_308 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_decap_8 FILLER_9_332 ();
 sg13g2_decap_8 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_346 ();
 sg13g2_fill_1 FILLER_9_348 ();
 sg13g2_fill_1 FILLER_9_401 ();
 sg13g2_fill_2 FILLER_9_433 ();
 sg13g2_fill_2 FILLER_9_443 ();
 sg13g2_fill_2 FILLER_9_486 ();
 sg13g2_fill_1 FILLER_9_488 ();
 sg13g2_fill_1 FILLER_9_519 ();
 sg13g2_fill_1 FILLER_9_538 ();
 sg13g2_fill_1 FILLER_9_591 ();
 sg13g2_fill_1 FILLER_9_598 ();
 sg13g2_decap_8 FILLER_9_716 ();
 sg13g2_decap_8 FILLER_9_723 ();
 sg13g2_decap_8 FILLER_9_730 ();
 sg13g2_fill_2 FILLER_9_737 ();
 sg13g2_fill_1 FILLER_9_748 ();
 sg13g2_fill_2 FILLER_9_779 ();
 sg13g2_decap_4 FILLER_9_791 ();
 sg13g2_fill_2 FILLER_9_795 ();
 sg13g2_fill_1 FILLER_9_823 ();
 sg13g2_decap_8 FILLER_9_843 ();
 sg13g2_decap_8 FILLER_9_850 ();
 sg13g2_decap_8 FILLER_9_857 ();
 sg13g2_fill_2 FILLER_9_864 ();
 sg13g2_fill_1 FILLER_9_866 ();
 sg13g2_decap_8 FILLER_9_879 ();
 sg13g2_decap_8 FILLER_9_886 ();
 sg13g2_decap_8 FILLER_9_893 ();
 sg13g2_decap_4 FILLER_9_900 ();
 sg13g2_decap_4 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_934 ();
 sg13g2_decap_4 FILLER_9_941 ();
 sg13g2_fill_2 FILLER_9_945 ();
 sg13g2_fill_2 FILLER_9_951 ();
 sg13g2_fill_2 FILLER_9_957 ();
 sg13g2_fill_2 FILLER_9_980 ();
 sg13g2_decap_4 FILLER_9_986 ();
 sg13g2_fill_1 FILLER_9_1014 ();
 sg13g2_fill_2 FILLER_9_1041 ();
 sg13g2_fill_1 FILLER_9_1049 ();
 sg13g2_fill_2 FILLER_9_1071 ();
 sg13g2_fill_1 FILLER_9_1073 ();
 sg13g2_fill_1 FILLER_9_1086 ();
 sg13g2_decap_8 FILLER_9_1098 ();
 sg13g2_fill_1 FILLER_9_1105 ();
 sg13g2_decap_4 FILLER_9_1111 ();
 sg13g2_fill_1 FILLER_9_1115 ();
 sg13g2_fill_2 FILLER_9_1148 ();
 sg13g2_fill_2 FILLER_9_1154 ();
 sg13g2_fill_2 FILLER_9_1166 ();
 sg13g2_fill_1 FILLER_9_1168 ();
 sg13g2_fill_2 FILLER_9_1173 ();
 sg13g2_decap_4 FILLER_9_1194 ();
 sg13g2_fill_2 FILLER_9_1198 ();
 sg13g2_decap_4 FILLER_9_1204 ();
 sg13g2_fill_2 FILLER_9_1208 ();
 sg13g2_decap_4 FILLER_9_1220 ();
 sg13g2_fill_1 FILLER_9_1224 ();
 sg13g2_fill_2 FILLER_9_1229 ();
 sg13g2_decap_8 FILLER_9_1241 ();
 sg13g2_decap_4 FILLER_9_1248 ();
 sg13g2_fill_1 FILLER_9_1252 ();
 sg13g2_decap_8 FILLER_9_1298 ();
 sg13g2_fill_2 FILLER_9_1305 ();
 sg13g2_fill_1 FILLER_9_1307 ();
 sg13g2_fill_1 FILLER_9_1361 ();
 sg13g2_decap_8 FILLER_9_1402 ();
 sg13g2_decap_8 FILLER_9_1409 ();
 sg13g2_decap_8 FILLER_9_1416 ();
 sg13g2_fill_2 FILLER_9_1423 ();
 sg13g2_fill_2 FILLER_9_1465 ();
 sg13g2_decap_4 FILLER_9_1493 ();
 sg13g2_fill_2 FILLER_9_1497 ();
 sg13g2_fill_2 FILLER_9_1545 ();
 sg13g2_fill_1 FILLER_9_1547 ();
 sg13g2_fill_1 FILLER_9_1556 ();
 sg13g2_fill_2 FILLER_9_1588 ();
 sg13g2_decap_4 FILLER_9_1611 ();
 sg13g2_fill_2 FILLER_9_1624 ();
 sg13g2_fill_1 FILLER_9_1626 ();
 sg13g2_decap_4 FILLER_9_1641 ();
 sg13g2_decap_8 FILLER_9_1649 ();
 sg13g2_fill_1 FILLER_9_1656 ();
 sg13g2_decap_8 FILLER_9_1724 ();
 sg13g2_decap_8 FILLER_9_1731 ();
 sg13g2_decap_8 FILLER_9_1738 ();
 sg13g2_decap_8 FILLER_9_1745 ();
 sg13g2_decap_8 FILLER_9_1752 ();
 sg13g2_decap_8 FILLER_9_1759 ();
 sg13g2_decap_8 FILLER_9_1766 ();
 sg13g2_fill_1 FILLER_9_1773 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_9 ();
 sg13g2_fill_1 FILLER_10_66 ();
 sg13g2_fill_1 FILLER_10_93 ();
 sg13g2_fill_1 FILLER_10_119 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_139 ();
 sg13g2_decap_8 FILLER_10_146 ();
 sg13g2_decap_8 FILLER_10_153 ();
 sg13g2_decap_8 FILLER_10_160 ();
 sg13g2_decap_8 FILLER_10_167 ();
 sg13g2_fill_2 FILLER_10_174 ();
 sg13g2_fill_2 FILLER_10_201 ();
 sg13g2_fill_2 FILLER_10_219 ();
 sg13g2_fill_2 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_294 ();
 sg13g2_fill_1 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_318 ();
 sg13g2_decap_4 FILLER_10_325 ();
 sg13g2_fill_1 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_372 ();
 sg13g2_fill_1 FILLER_10_374 ();
 sg13g2_decap_4 FILLER_10_390 ();
 sg13g2_fill_1 FILLER_10_399 ();
 sg13g2_decap_4 FILLER_10_432 ();
 sg13g2_fill_1 FILLER_10_436 ();
 sg13g2_fill_1 FILLER_10_448 ();
 sg13g2_decap_4 FILLER_10_471 ();
 sg13g2_decap_4 FILLER_10_479 ();
 sg13g2_fill_2 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_523 ();
 sg13g2_decap_8 FILLER_10_530 ();
 sg13g2_decap_8 FILLER_10_537 ();
 sg13g2_decap_8 FILLER_10_544 ();
 sg13g2_fill_2 FILLER_10_551 ();
 sg13g2_fill_1 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_558 ();
 sg13g2_fill_2 FILLER_10_565 ();
 sg13g2_fill_1 FILLER_10_567 ();
 sg13g2_fill_1 FILLER_10_596 ();
 sg13g2_fill_1 FILLER_10_611 ();
 sg13g2_fill_1 FILLER_10_618 ();
 sg13g2_fill_1 FILLER_10_634 ();
 sg13g2_fill_2 FILLER_10_649 ();
 sg13g2_decap_8 FILLER_10_660 ();
 sg13g2_decap_8 FILLER_10_667 ();
 sg13g2_fill_2 FILLER_10_674 ();
 sg13g2_fill_1 FILLER_10_676 ();
 sg13g2_decap_8 FILLER_10_716 ();
 sg13g2_fill_1 FILLER_10_723 ();
 sg13g2_fill_1 FILLER_10_744 ();
 sg13g2_fill_2 FILLER_10_762 ();
 sg13g2_decap_4 FILLER_10_798 ();
 sg13g2_fill_1 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_4 FILLER_10_814 ();
 sg13g2_fill_2 FILLER_10_818 ();
 sg13g2_decap_8 FILLER_10_825 ();
 sg13g2_decap_8 FILLER_10_832 ();
 sg13g2_fill_1 FILLER_10_839 ();
 sg13g2_decap_4 FILLER_10_870 ();
 sg13g2_fill_1 FILLER_10_874 ();
 sg13g2_decap_8 FILLER_10_896 ();
 sg13g2_fill_1 FILLER_10_929 ();
 sg13g2_decap_4 FILLER_10_943 ();
 sg13g2_fill_1 FILLER_10_951 ();
 sg13g2_decap_8 FILLER_10_996 ();
 sg13g2_fill_2 FILLER_10_1003 ();
 sg13g2_fill_1 FILLER_10_1005 ();
 sg13g2_fill_1 FILLER_10_1073 ();
 sg13g2_fill_1 FILLER_10_1080 ();
 sg13g2_decap_8 FILLER_10_1100 ();
 sg13g2_decap_4 FILLER_10_1107 ();
 sg13g2_fill_1 FILLER_10_1111 ();
 sg13g2_decap_8 FILLER_10_1126 ();
 sg13g2_decap_8 FILLER_10_1133 ();
 sg13g2_decap_8 FILLER_10_1140 ();
 sg13g2_decap_4 FILLER_10_1147 ();
 sg13g2_fill_1 FILLER_10_1151 ();
 sg13g2_decap_8 FILLER_10_1188 ();
 sg13g2_decap_4 FILLER_10_1195 ();
 sg13g2_fill_2 FILLER_10_1199 ();
 sg13g2_decap_8 FILLER_10_1204 ();
 sg13g2_decap_8 FILLER_10_1211 ();
 sg13g2_fill_1 FILLER_10_1280 ();
 sg13g2_decap_4 FILLER_10_1295 ();
 sg13g2_fill_2 FILLER_10_1299 ();
 sg13g2_decap_8 FILLER_10_1314 ();
 sg13g2_fill_2 FILLER_10_1376 ();
 sg13g2_decap_8 FILLER_10_1404 ();
 sg13g2_decap_8 FILLER_10_1411 ();
 sg13g2_decap_8 FILLER_10_1418 ();
 sg13g2_decap_8 FILLER_10_1425 ();
 sg13g2_decap_8 FILLER_10_1432 ();
 sg13g2_decap_4 FILLER_10_1439 ();
 sg13g2_fill_2 FILLER_10_1443 ();
 sg13g2_decap_8 FILLER_10_1449 ();
 sg13g2_decap_4 FILLER_10_1456 ();
 sg13g2_fill_1 FILLER_10_1460 ();
 sg13g2_decap_4 FILLER_10_1479 ();
 sg13g2_fill_1 FILLER_10_1483 ();
 sg13g2_decap_8 FILLER_10_1489 ();
 sg13g2_fill_2 FILLER_10_1496 ();
 sg13g2_fill_2 FILLER_10_1506 ();
 sg13g2_decap_8 FILLER_10_1538 ();
 sg13g2_fill_2 FILLER_10_1545 ();
 sg13g2_fill_1 FILLER_10_1547 ();
 sg13g2_decap_4 FILLER_10_1574 ();
 sg13g2_fill_1 FILLER_10_1578 ();
 sg13g2_fill_1 FILLER_10_1583 ();
 sg13g2_decap_8 FILLER_10_1588 ();
 sg13g2_decap_8 FILLER_10_1595 ();
 sg13g2_decap_8 FILLER_10_1602 ();
 sg13g2_decap_8 FILLER_10_1609 ();
 sg13g2_decap_8 FILLER_10_1616 ();
 sg13g2_fill_2 FILLER_10_1623 ();
 sg13g2_fill_2 FILLER_10_1635 ();
 sg13g2_decap_8 FILLER_10_1663 ();
 sg13g2_decap_4 FILLER_10_1670 ();
 sg13g2_fill_1 FILLER_10_1674 ();
 sg13g2_decap_4 FILLER_10_1685 ();
 sg13g2_fill_2 FILLER_10_1689 ();
 sg13g2_decap_4 FILLER_10_1717 ();
 sg13g2_fill_1 FILLER_10_1721 ();
 sg13g2_decap_8 FILLER_10_1726 ();
 sg13g2_decap_8 FILLER_10_1733 ();
 sg13g2_decap_8 FILLER_10_1740 ();
 sg13g2_decap_8 FILLER_10_1747 ();
 sg13g2_decap_8 FILLER_10_1754 ();
 sg13g2_decap_8 FILLER_10_1761 ();
 sg13g2_decap_4 FILLER_10_1768 ();
 sg13g2_fill_2 FILLER_10_1772 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_fill_2 FILLER_11_57 ();
 sg13g2_fill_1 FILLER_11_59 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_145 ();
 sg13g2_fill_2 FILLER_11_156 ();
 sg13g2_decap_8 FILLER_11_162 ();
 sg13g2_decap_4 FILLER_11_169 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_fill_2 FILLER_11_238 ();
 sg13g2_fill_1 FILLER_11_240 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_fill_1 FILLER_11_252 ();
 sg13g2_fill_1 FILLER_11_278 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_fill_1 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_decap_8 FILLER_11_407 ();
 sg13g2_fill_2 FILLER_11_418 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_4 FILLER_11_441 ();
 sg13g2_fill_1 FILLER_11_445 ();
 sg13g2_fill_1 FILLER_11_486 ();
 sg13g2_decap_4 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_537 ();
 sg13g2_fill_2 FILLER_11_544 ();
 sg13g2_fill_1 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_555 ();
 sg13g2_fill_2 FILLER_11_562 ();
 sg13g2_fill_1 FILLER_11_564 ();
 sg13g2_fill_1 FILLER_11_574 ();
 sg13g2_fill_1 FILLER_11_584 ();
 sg13g2_fill_1 FILLER_11_589 ();
 sg13g2_decap_4 FILLER_11_595 ();
 sg13g2_fill_2 FILLER_11_608 ();
 sg13g2_fill_1 FILLER_11_610 ();
 sg13g2_fill_1 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_664 ();
 sg13g2_decap_8 FILLER_11_671 ();
 sg13g2_decap_4 FILLER_11_678 ();
 sg13g2_decap_4 FILLER_11_686 ();
 sg13g2_fill_2 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_698 ();
 sg13g2_decap_4 FILLER_11_720 ();
 sg13g2_fill_2 FILLER_11_784 ();
 sg13g2_fill_1 FILLER_11_786 ();
 sg13g2_decap_8 FILLER_11_817 ();
 sg13g2_decap_8 FILLER_11_824 ();
 sg13g2_decap_4 FILLER_11_831 ();
 sg13g2_fill_2 FILLER_11_835 ();
 sg13g2_fill_2 FILLER_11_850 ();
 sg13g2_fill_1 FILLER_11_852 ();
 sg13g2_decap_8 FILLER_11_863 ();
 sg13g2_decap_8 FILLER_11_870 ();
 sg13g2_decap_8 FILLER_11_877 ();
 sg13g2_decap_8 FILLER_11_884 ();
 sg13g2_decap_8 FILLER_11_891 ();
 sg13g2_decap_8 FILLER_11_898 ();
 sg13g2_decap_8 FILLER_11_905 ();
 sg13g2_decap_8 FILLER_11_912 ();
 sg13g2_decap_8 FILLER_11_919 ();
 sg13g2_decap_8 FILLER_11_926 ();
 sg13g2_decap_8 FILLER_11_933 ();
 sg13g2_decap_8 FILLER_11_940 ();
 sg13g2_decap_8 FILLER_11_947 ();
 sg13g2_fill_2 FILLER_11_954 ();
 sg13g2_decap_8 FILLER_11_964 ();
 sg13g2_decap_4 FILLER_11_971 ();
 sg13g2_fill_2 FILLER_11_975 ();
 sg13g2_fill_2 FILLER_11_1106 ();
 sg13g2_decap_8 FILLER_11_1112 ();
 sg13g2_fill_2 FILLER_11_1119 ();
 sg13g2_decap_4 FILLER_11_1133 ();
 sg13g2_decap_4 FILLER_11_1171 ();
 sg13g2_fill_1 FILLER_11_1175 ();
 sg13g2_decap_4 FILLER_11_1189 ();
 sg13g2_fill_2 FILLER_11_1193 ();
 sg13g2_fill_2 FILLER_11_1214 ();
 sg13g2_fill_1 FILLER_11_1216 ();
 sg13g2_fill_1 FILLER_11_1227 ();
 sg13g2_fill_1 FILLER_11_1232 ();
 sg13g2_fill_1 FILLER_11_1237 ();
 sg13g2_fill_2 FILLER_11_1259 ();
 sg13g2_fill_1 FILLER_11_1266 ();
 sg13g2_fill_2 FILLER_11_1288 ();
 sg13g2_decap_4 FILLER_11_1320 ();
 sg13g2_fill_1 FILLER_11_1324 ();
 sg13g2_decap_8 FILLER_11_1351 ();
 sg13g2_decap_8 FILLER_11_1358 ();
 sg13g2_decap_8 FILLER_11_1365 ();
 sg13g2_decap_8 FILLER_11_1372 ();
 sg13g2_decap_4 FILLER_11_1379 ();
 sg13g2_fill_2 FILLER_11_1383 ();
 sg13g2_fill_2 FILLER_11_1389 ();
 sg13g2_decap_4 FILLER_11_1395 ();
 sg13g2_decap_4 FILLER_11_1409 ();
 sg13g2_decap_8 FILLER_11_1439 ();
 sg13g2_decap_8 FILLER_11_1446 ();
 sg13g2_decap_8 FILLER_11_1463 ();
 sg13g2_fill_1 FILLER_11_1470 ();
 sg13g2_decap_4 FILLER_11_1507 ();
 sg13g2_fill_2 FILLER_11_1511 ();
 sg13g2_decap_8 FILLER_11_1527 ();
 sg13g2_decap_8 FILLER_11_1534 ();
 sg13g2_decap_8 FILLER_11_1541 ();
 sg13g2_decap_8 FILLER_11_1548 ();
 sg13g2_decap_8 FILLER_11_1555 ();
 sg13g2_fill_2 FILLER_11_1562 ();
 sg13g2_decap_8 FILLER_11_1568 ();
 sg13g2_decap_8 FILLER_11_1575 ();
 sg13g2_decap_8 FILLER_11_1582 ();
 sg13g2_decap_8 FILLER_11_1589 ();
 sg13g2_decap_8 FILLER_11_1596 ();
 sg13g2_decap_8 FILLER_11_1603 ();
 sg13g2_decap_8 FILLER_11_1610 ();
 sg13g2_fill_2 FILLER_11_1617 ();
 sg13g2_decap_8 FILLER_11_1739 ();
 sg13g2_decap_8 FILLER_11_1746 ();
 sg13g2_decap_8 FILLER_11_1753 ();
 sg13g2_decap_8 FILLER_11_1760 ();
 sg13g2_decap_8 FILLER_11_1767 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_48 ();
 sg13g2_fill_2 FILLER_12_55 ();
 sg13g2_fill_1 FILLER_12_57 ();
 sg13g2_fill_2 FILLER_12_98 ();
 sg13g2_fill_2 FILLER_12_110 ();
 sg13g2_fill_1 FILLER_12_138 ();
 sg13g2_fill_2 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_fill_2 FILLER_12_176 ();
 sg13g2_fill_1 FILLER_12_178 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_fill_2 FILLER_12_196 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_4 FILLER_12_242 ();
 sg13g2_fill_1 FILLER_12_246 ();
 sg13g2_decap_8 FILLER_12_250 ();
 sg13g2_decap_8 FILLER_12_257 ();
 sg13g2_decap_4 FILLER_12_264 ();
 sg13g2_fill_2 FILLER_12_268 ();
 sg13g2_fill_2 FILLER_12_284 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_fill_1 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_fill_1 FILLER_12_379 ();
 sg13g2_decap_4 FILLER_12_416 ();
 sg13g2_fill_2 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_429 ();
 sg13g2_fill_1 FILLER_12_431 ();
 sg13g2_fill_1 FILLER_12_464 ();
 sg13g2_fill_2 FILLER_12_501 ();
 sg13g2_fill_2 FILLER_12_555 ();
 sg13g2_fill_2 FILLER_12_561 ();
 sg13g2_fill_1 FILLER_12_589 ();
 sg13g2_fill_2 FILLER_12_611 ();
 sg13g2_fill_1 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_664 ();
 sg13g2_decap_8 FILLER_12_671 ();
 sg13g2_decap_8 FILLER_12_678 ();
 sg13g2_decap_8 FILLER_12_685 ();
 sg13g2_decap_4 FILLER_12_698 ();
 sg13g2_fill_2 FILLER_12_702 ();
 sg13g2_fill_1 FILLER_12_710 ();
 sg13g2_fill_1 FILLER_12_715 ();
 sg13g2_fill_2 FILLER_12_726 ();
 sg13g2_fill_1 FILLER_12_754 ();
 sg13g2_fill_2 FILLER_12_765 ();
 sg13g2_fill_2 FILLER_12_773 ();
 sg13g2_fill_2 FILLER_12_793 ();
 sg13g2_fill_2 FILLER_12_821 ();
 sg13g2_decap_8 FILLER_12_827 ();
 sg13g2_decap_8 FILLER_12_834 ();
 sg13g2_decap_8 FILLER_12_841 ();
 sg13g2_decap_8 FILLER_12_848 ();
 sg13g2_decap_8 FILLER_12_855 ();
 sg13g2_decap_8 FILLER_12_862 ();
 sg13g2_decap_8 FILLER_12_869 ();
 sg13g2_decap_8 FILLER_12_876 ();
 sg13g2_decap_8 FILLER_12_883 ();
 sg13g2_decap_8 FILLER_12_890 ();
 sg13g2_fill_2 FILLER_12_897 ();
 sg13g2_decap_4 FILLER_12_924 ();
 sg13g2_fill_2 FILLER_12_928 ();
 sg13g2_decap_4 FILLER_12_943 ();
 sg13g2_fill_1 FILLER_12_947 ();
 sg13g2_fill_2 FILLER_12_982 ();
 sg13g2_fill_1 FILLER_12_984 ();
 sg13g2_decap_4 FILLER_12_1006 ();
 sg13g2_fill_1 FILLER_12_1010 ();
 sg13g2_decap_4 FILLER_12_1021 ();
 sg13g2_fill_1 FILLER_12_1025 ();
 sg13g2_fill_2 FILLER_12_1030 ();
 sg13g2_fill_1 FILLER_12_1032 ();
 sg13g2_decap_8 FILLER_12_1037 ();
 sg13g2_fill_2 FILLER_12_1044 ();
 sg13g2_fill_1 FILLER_12_1046 ();
 sg13g2_fill_1 FILLER_12_1057 ();
 sg13g2_fill_1 FILLER_12_1062 ();
 sg13g2_fill_2 FILLER_12_1089 ();
 sg13g2_fill_1 FILLER_12_1091 ();
 sg13g2_decap_8 FILLER_12_1127 ();
 sg13g2_fill_2 FILLER_12_1164 ();
 sg13g2_fill_2 FILLER_12_1196 ();
 sg13g2_fill_1 FILLER_12_1204 ();
 sg13g2_fill_2 FILLER_12_1261 ();
 sg13g2_fill_1 FILLER_12_1263 ();
 sg13g2_decap_8 FILLER_12_1289 ();
 sg13g2_decap_8 FILLER_12_1296 ();
 sg13g2_decap_8 FILLER_12_1303 ();
 sg13g2_decap_8 FILLER_12_1310 ();
 sg13g2_decap_4 FILLER_12_1317 ();
 sg13g2_fill_2 FILLER_12_1321 ();
 sg13g2_decap_8 FILLER_12_1363 ();
 sg13g2_decap_8 FILLER_12_1370 ();
 sg13g2_fill_2 FILLER_12_1377 ();
 sg13g2_fill_1 FILLER_12_1379 ();
 sg13g2_fill_2 FILLER_12_1427 ();
 sg13g2_fill_2 FILLER_12_1455 ();
 sg13g2_fill_1 FILLER_12_1457 ();
 sg13g2_fill_2 FILLER_12_1484 ();
 sg13g2_fill_1 FILLER_12_1486 ();
 sg13g2_decap_4 FILLER_12_1491 ();
 sg13g2_fill_1 FILLER_12_1495 ();
 sg13g2_fill_1 FILLER_12_1510 ();
 sg13g2_decap_8 FILLER_12_1560 ();
 sg13g2_decap_8 FILLER_12_1567 ();
 sg13g2_fill_1 FILLER_12_1574 ();
 sg13g2_decap_4 FILLER_12_1588 ();
 sg13g2_fill_1 FILLER_12_1592 ();
 sg13g2_decap_4 FILLER_12_1597 ();
 sg13g2_fill_2 FILLER_12_1601 ();
 sg13g2_decap_8 FILLER_12_1611 ();
 sg13g2_decap_4 FILLER_12_1618 ();
 sg13g2_fill_1 FILLER_12_1622 ();
 sg13g2_decap_4 FILLER_12_1628 ();
 sg13g2_fill_2 FILLER_12_1632 ();
 sg13g2_fill_1 FILLER_12_1678 ();
 sg13g2_decap_8 FILLER_12_1715 ();
 sg13g2_decap_8 FILLER_12_1722 ();
 sg13g2_decap_8 FILLER_12_1729 ();
 sg13g2_decap_8 FILLER_12_1736 ();
 sg13g2_decap_4 FILLER_12_1743 ();
 sg13g2_fill_1 FILLER_12_1747 ();
 sg13g2_decap_8 FILLER_12_1752 ();
 sg13g2_decap_8 FILLER_12_1759 ();
 sg13g2_decap_8 FILLER_12_1766 ();
 sg13g2_fill_1 FILLER_12_1773 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_16 ();
 sg13g2_decap_8 FILLER_13_47 ();
 sg13g2_fill_2 FILLER_13_54 ();
 sg13g2_decap_8 FILLER_13_87 ();
 sg13g2_decap_4 FILLER_13_94 ();
 sg13g2_fill_2 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_104 ();
 sg13g2_decap_8 FILLER_13_111 ();
 sg13g2_decap_8 FILLER_13_118 ();
 sg13g2_decap_8 FILLER_13_125 ();
 sg13g2_decap_8 FILLER_13_132 ();
 sg13g2_decap_8 FILLER_13_139 ();
 sg13g2_fill_1 FILLER_13_146 ();
 sg13g2_fill_1 FILLER_13_157 ();
 sg13g2_fill_2 FILLER_13_218 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_4 FILLER_13_238 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_decap_8 FILLER_13_262 ();
 sg13g2_decap_8 FILLER_13_269 ();
 sg13g2_fill_1 FILLER_13_276 ();
 sg13g2_fill_2 FILLER_13_303 ();
 sg13g2_fill_1 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_fill_1 FILLER_13_339 ();
 sg13g2_fill_2 FILLER_13_344 ();
 sg13g2_decap_4 FILLER_13_350 ();
 sg13g2_decap_4 FILLER_13_364 ();
 sg13g2_decap_4 FILLER_13_394 ();
 sg13g2_fill_2 FILLER_13_408 ();
 sg13g2_decap_4 FILLER_13_440 ();
 sg13g2_fill_1 FILLER_13_444 ();
 sg13g2_fill_1 FILLER_13_464 ();
 sg13g2_fill_2 FILLER_13_469 ();
 sg13g2_fill_1 FILLER_13_507 ();
 sg13g2_fill_2 FILLER_13_520 ();
 sg13g2_fill_1 FILLER_13_522 ();
 sg13g2_fill_2 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_fill_2 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_fill_2 FILLER_13_672 ();
 sg13g2_fill_1 FILLER_13_674 ();
 sg13g2_decap_4 FILLER_13_738 ();
 sg13g2_fill_2 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_fill_1 FILLER_13_777 ();
 sg13g2_decap_4 FILLER_13_788 ();
 sg13g2_decap_4 FILLER_13_800 ();
 sg13g2_fill_1 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_867 ();
 sg13g2_decap_8 FILLER_13_874 ();
 sg13g2_decap_8 FILLER_13_881 ();
 sg13g2_decap_8 FILLER_13_888 ();
 sg13g2_decap_8 FILLER_13_895 ();
 sg13g2_decap_8 FILLER_13_902 ();
 sg13g2_decap_4 FILLER_13_909 ();
 sg13g2_fill_1 FILLER_13_913 ();
 sg13g2_decap_8 FILLER_13_927 ();
 sg13g2_decap_8 FILLER_13_934 ();
 sg13g2_decap_4 FILLER_13_941 ();
 sg13g2_fill_1 FILLER_13_945 ();
 sg13g2_decap_4 FILLER_13_982 ();
 sg13g2_decap_8 FILLER_13_990 ();
 sg13g2_fill_2 FILLER_13_1049 ();
 sg13g2_decap_8 FILLER_13_1061 ();
 sg13g2_fill_1 FILLER_13_1073 ();
 sg13g2_fill_1 FILLER_13_1078 ();
 sg13g2_fill_2 FILLER_13_1113 ();
 sg13g2_fill_1 FILLER_13_1120 ();
 sg13g2_decap_8 FILLER_13_1124 ();
 sg13g2_decap_4 FILLER_13_1131 ();
 sg13g2_decap_8 FILLER_13_1265 ();
 sg13g2_fill_1 FILLER_13_1272 ();
 sg13g2_decap_8 FILLER_13_1279 ();
 sg13g2_decap_8 FILLER_13_1286 ();
 sg13g2_fill_2 FILLER_13_1293 ();
 sg13g2_fill_1 FILLER_13_1295 ();
 sg13g2_decap_4 FILLER_13_1326 ();
 sg13g2_fill_1 FILLER_13_1330 ();
 sg13g2_fill_2 FILLER_13_1408 ();
 sg13g2_fill_2 FILLER_13_1420 ();
 sg13g2_decap_4 FILLER_13_1440 ();
 sg13g2_decap_8 FILLER_13_1555 ();
 sg13g2_decap_8 FILLER_13_1562 ();
 sg13g2_decap_8 FILLER_13_1569 ();
 sg13g2_decap_8 FILLER_13_1646 ();
 sg13g2_fill_1 FILLER_13_1653 ();
 sg13g2_decap_4 FILLER_13_1658 ();
 sg13g2_fill_2 FILLER_13_1662 ();
 sg13g2_decap_4 FILLER_13_1695 ();
 sg13g2_decap_8 FILLER_13_1703 ();
 sg13g2_decap_8 FILLER_13_1710 ();
 sg13g2_decap_8 FILLER_13_1717 ();
 sg13g2_decap_8 FILLER_13_1724 ();
 sg13g2_decap_8 FILLER_13_1767 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_23 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_65 ();
 sg13g2_decap_8 FILLER_14_71 ();
 sg13g2_fill_2 FILLER_14_78 ();
 sg13g2_fill_1 FILLER_14_80 ();
 sg13g2_decap_8 FILLER_14_111 ();
 sg13g2_decap_8 FILLER_14_118 ();
 sg13g2_decap_4 FILLER_14_125 ();
 sg13g2_decap_4 FILLER_14_133 ();
 sg13g2_fill_2 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_152 ();
 sg13g2_decap_4 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_decap_8 FILLER_14_219 ();
 sg13g2_fill_2 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_228 ();
 sg13g2_fill_2 FILLER_14_239 ();
 sg13g2_fill_1 FILLER_14_241 ();
 sg13g2_fill_1 FILLER_14_268 ();
 sg13g2_fill_1 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_fill_2 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_fill_2 FILLER_14_298 ();
 sg13g2_decap_4 FILLER_14_336 ();
 sg13g2_decap_4 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_414 ();
 sg13g2_decap_4 FILLER_14_447 ();
 sg13g2_fill_1 FILLER_14_451 ();
 sg13g2_fill_2 FILLER_14_456 ();
 sg13g2_decap_4 FILLER_14_461 ();
 sg13g2_fill_2 FILLER_14_465 ();
 sg13g2_fill_2 FILLER_14_501 ();
 sg13g2_fill_2 FILLER_14_537 ();
 sg13g2_fill_1 FILLER_14_539 ();
 sg13g2_fill_1 FILLER_14_567 ();
 sg13g2_fill_2 FILLER_14_633 ();
 sg13g2_fill_2 FILLER_14_651 ();
 sg13g2_fill_1 FILLER_14_653 ();
 sg13g2_decap_8 FILLER_14_668 ();
 sg13g2_decap_4 FILLER_14_675 ();
 sg13g2_fill_1 FILLER_14_719 ();
 sg13g2_fill_1 FILLER_14_730 ();
 sg13g2_fill_1 FILLER_14_752 ();
 sg13g2_decap_4 FILLER_14_774 ();
 sg13g2_decap_4 FILLER_14_782 ();
 sg13g2_decap_4 FILLER_14_806 ();
 sg13g2_decap_8 FILLER_14_862 ();
 sg13g2_decap_8 FILLER_14_869 ();
 sg13g2_decap_8 FILLER_14_876 ();
 sg13g2_decap_8 FILLER_14_883 ();
 sg13g2_decap_8 FILLER_14_890 ();
 sg13g2_decap_4 FILLER_14_897 ();
 sg13g2_decap_8 FILLER_14_914 ();
 sg13g2_fill_2 FILLER_14_921 ();
 sg13g2_fill_1 FILLER_14_923 ();
 sg13g2_decap_4 FILLER_14_937 ();
 sg13g2_fill_1 FILLER_14_941 ();
 sg13g2_decap_8 FILLER_14_979 ();
 sg13g2_fill_2 FILLER_14_986 ();
 sg13g2_decap_8 FILLER_14_1022 ();
 sg13g2_decap_8 FILLER_14_1029 ();
 sg13g2_decap_8 FILLER_14_1036 ();
 sg13g2_decap_8 FILLER_14_1043 ();
 sg13g2_decap_8 FILLER_14_1064 ();
 sg13g2_fill_2 FILLER_14_1071 ();
 sg13g2_fill_1 FILLER_14_1073 ();
 sg13g2_fill_2 FILLER_14_1084 ();
 sg13g2_fill_1 FILLER_14_1086 ();
 sg13g2_decap_8 FILLER_14_1113 ();
 sg13g2_decap_8 FILLER_14_1120 ();
 sg13g2_decap_8 FILLER_14_1131 ();
 sg13g2_fill_2 FILLER_14_1138 ();
 sg13g2_fill_2 FILLER_14_1181 ();
 sg13g2_fill_2 FILLER_14_1189 ();
 sg13g2_fill_1 FILLER_14_1210 ();
 sg13g2_fill_2 FILLER_14_1236 ();
 sg13g2_fill_1 FILLER_14_1248 ();
 sg13g2_decap_8 FILLER_14_1253 ();
 sg13g2_decap_8 FILLER_14_1260 ();
 sg13g2_decap_4 FILLER_14_1267 ();
 sg13g2_fill_2 FILLER_14_1271 ();
 sg13g2_decap_8 FILLER_14_1276 ();
 sg13g2_decap_8 FILLER_14_1283 ();
 sg13g2_decap_8 FILLER_14_1361 ();
 sg13g2_decap_8 FILLER_14_1368 ();
 sg13g2_decap_8 FILLER_14_1375 ();
 sg13g2_decap_8 FILLER_14_1382 ();
 sg13g2_fill_2 FILLER_14_1407 ();
 sg13g2_decap_8 FILLER_14_1435 ();
 sg13g2_fill_2 FILLER_14_1452 ();
 sg13g2_decap_4 FILLER_14_1458 ();
 sg13g2_fill_2 FILLER_14_1462 ();
 sg13g2_fill_2 FILLER_14_1474 ();
 sg13g2_fill_1 FILLER_14_1532 ();
 sg13g2_fill_1 FILLER_14_1564 ();
 sg13g2_fill_2 FILLER_14_1644 ();
 sg13g2_fill_1 FILLER_14_1646 ();
 sg13g2_decap_8 FILLER_14_1673 ();
 sg13g2_fill_2 FILLER_14_1680 ();
 sg13g2_fill_1 FILLER_14_1682 ();
 sg13g2_decap_8 FILLER_14_1687 ();
 sg13g2_decap_8 FILLER_14_1694 ();
 sg13g2_fill_2 FILLER_14_1701 ();
 sg13g2_fill_1 FILLER_14_1703 ();
 sg13g2_decap_4 FILLER_14_1725 ();
 sg13g2_fill_2 FILLER_14_1729 ();
 sg13g2_decap_8 FILLER_14_1767 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_fill_2 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_fill_1 FILLER_15_69 ();
 sg13g2_decap_4 FILLER_15_106 ();
 sg13g2_fill_2 FILLER_15_110 ();
 sg13g2_fill_1 FILLER_15_184 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_fill_2 FILLER_15_295 ();
 sg13g2_fill_1 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_4 FILLER_15_455 ();
 sg13g2_fill_1 FILLER_15_459 ();
 sg13g2_decap_4 FILLER_15_464 ();
 sg13g2_fill_2 FILLER_15_468 ();
 sg13g2_decap_8 FILLER_15_482 ();
 sg13g2_fill_2 FILLER_15_489 ();
 sg13g2_fill_1 FILLER_15_499 ();
 sg13g2_fill_2 FILLER_15_561 ();
 sg13g2_fill_1 FILLER_15_563 ();
 sg13g2_fill_2 FILLER_15_570 ();
 sg13g2_fill_1 FILLER_15_572 ();
 sg13g2_fill_2 FILLER_15_633 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_fill_1 FILLER_15_669 ();
 sg13g2_decap_4 FILLER_15_678 ();
 sg13g2_fill_2 FILLER_15_682 ();
 sg13g2_decap_8 FILLER_15_715 ();
 sg13g2_decap_8 FILLER_15_722 ();
 sg13g2_decap_4 FILLER_15_729 ();
 sg13g2_fill_2 FILLER_15_733 ();
 sg13g2_decap_4 FILLER_15_765 ();
 sg13g2_fill_1 FILLER_15_795 ();
 sg13g2_decap_4 FILLER_15_843 ();
 sg13g2_decap_8 FILLER_15_855 ();
 sg13g2_decap_8 FILLER_15_862 ();
 sg13g2_fill_2 FILLER_15_869 ();
 sg13g2_fill_2 FILLER_15_892 ();
 sg13g2_fill_1 FILLER_15_894 ();
 sg13g2_decap_4 FILLER_15_920 ();
 sg13g2_fill_1 FILLER_15_924 ();
 sg13g2_decap_8 FILLER_15_981 ();
 sg13g2_fill_2 FILLER_15_988 ();
 sg13g2_decap_8 FILLER_15_1014 ();
 sg13g2_fill_2 FILLER_15_1031 ();
 sg13g2_fill_1 FILLER_15_1033 ();
 sg13g2_fill_2 FILLER_15_1038 ();
 sg13g2_fill_1 FILLER_15_1040 ();
 sg13g2_fill_2 FILLER_15_1051 ();
 sg13g2_fill_2 FILLER_15_1079 ();
 sg13g2_fill_2 FILLER_15_1137 ();
 sg13g2_decap_4 FILLER_15_1149 ();
 sg13g2_fill_1 FILLER_15_1186 ();
 sg13g2_decap_8 FILLER_15_1254 ();
 sg13g2_decap_8 FILLER_15_1261 ();
 sg13g2_decap_8 FILLER_15_1268 ();
 sg13g2_decap_4 FILLER_15_1275 ();
 sg13g2_decap_4 FILLER_15_1315 ();
 sg13g2_fill_2 FILLER_15_1319 ();
 sg13g2_decap_8 FILLER_15_1331 ();
 sg13g2_decap_4 FILLER_15_1338 ();
 sg13g2_decap_8 FILLER_15_1350 ();
 sg13g2_decap_8 FILLER_15_1357 ();
 sg13g2_decap_8 FILLER_15_1364 ();
 sg13g2_decap_8 FILLER_15_1371 ();
 sg13g2_decap_4 FILLER_15_1378 ();
 sg13g2_fill_1 FILLER_15_1382 ();
 sg13g2_fill_2 FILLER_15_1409 ();
 sg13g2_fill_1 FILLER_15_1415 ();
 sg13g2_decap_4 FILLER_15_1447 ();
 sg13g2_fill_1 FILLER_15_1503 ();
 sg13g2_fill_1 FILLER_15_1511 ();
 sg13g2_fill_2 FILLER_15_1515 ();
 sg13g2_fill_1 FILLER_15_1517 ();
 sg13g2_fill_2 FILLER_15_1575 ();
 sg13g2_fill_1 FILLER_15_1577 ();
 sg13g2_decap_4 FILLER_15_1599 ();
 sg13g2_fill_1 FILLER_15_1603 ();
 sg13g2_fill_2 FILLER_15_1614 ();
 sg13g2_fill_2 FILLER_15_1642 ();
 sg13g2_fill_2 FILLER_15_1654 ();
 sg13g2_fill_1 FILLER_15_1656 ();
 sg13g2_fill_2 FILLER_15_1661 ();
 sg13g2_fill_1 FILLER_15_1663 ();
 sg13g2_fill_2 FILLER_15_1674 ();
 sg13g2_decap_8 FILLER_15_1757 ();
 sg13g2_decap_8 FILLER_15_1764 ();
 sg13g2_fill_2 FILLER_15_1771 ();
 sg13g2_fill_1 FILLER_15_1773 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_fill_2 FILLER_16_10 ();
 sg13g2_decap_8 FILLER_16_38 ();
 sg13g2_decap_4 FILLER_16_48 ();
 sg13g2_fill_1 FILLER_16_52 ();
 sg13g2_decap_4 FILLER_16_77 ();
 sg13g2_fill_1 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_99 ();
 sg13g2_fill_2 FILLER_16_106 ();
 sg13g2_decap_8 FILLER_16_148 ();
 sg13g2_fill_2 FILLER_16_155 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_1 FILLER_16_167 ();
 sg13g2_decap_4 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_fill_2 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_205 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_fill_1 FILLER_16_297 ();
 sg13g2_decap_4 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_362 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_fill_1 FILLER_16_383 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_fill_1 FILLER_16_413 ();
 sg13g2_fill_2 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_424 ();
 sg13g2_fill_2 FILLER_16_451 ();
 sg13g2_decap_8 FILLER_16_461 ();
 sg13g2_decap_8 FILLER_16_468 ();
 sg13g2_fill_2 FILLER_16_475 ();
 sg13g2_fill_1 FILLER_16_477 ();
 sg13g2_decap_8 FILLER_16_492 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_fill_2 FILLER_16_506 ();
 sg13g2_fill_1 FILLER_16_508 ();
 sg13g2_fill_1 FILLER_16_527 ();
 sg13g2_decap_8 FILLER_16_554 ();
 sg13g2_decap_8 FILLER_16_561 ();
 sg13g2_decap_8 FILLER_16_568 ();
 sg13g2_fill_1 FILLER_16_620 ();
 sg13g2_fill_2 FILLER_16_642 ();
 sg13g2_fill_1 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_652 ();
 sg13g2_fill_2 FILLER_16_659 ();
 sg13g2_decap_4 FILLER_16_682 ();
 sg13g2_fill_2 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_4 FILLER_16_746 ();
 sg13g2_fill_1 FILLER_16_750 ();
 sg13g2_fill_1 FILLER_16_777 ();
 sg13g2_fill_2 FILLER_16_783 ();
 sg13g2_fill_1 FILLER_16_816 ();
 sg13g2_decap_4 FILLER_16_821 ();
 sg13g2_fill_1 FILLER_16_825 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_decap_4 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_16_888 ();
 sg13g2_fill_2 FILLER_16_895 ();
 sg13g2_decap_8 FILLER_16_936 ();
 sg13g2_fill_2 FILLER_16_943 ();
 sg13g2_decap_8 FILLER_16_981 ();
 sg13g2_decap_8 FILLER_16_988 ();
 sg13g2_decap_4 FILLER_16_995 ();
 sg13g2_fill_2 FILLER_16_999 ();
 sg13g2_fill_1 FILLER_16_1057 ();
 sg13g2_fill_2 FILLER_16_1130 ();
 sg13g2_fill_1 FILLER_16_1158 ();
 sg13g2_fill_2 FILLER_16_1211 ();
 sg13g2_fill_1 FILLER_16_1216 ();
 sg13g2_decap_8 FILLER_16_1221 ();
 sg13g2_fill_2 FILLER_16_1264 ();
 sg13g2_fill_1 FILLER_16_1266 ();
 sg13g2_fill_2 FILLER_16_1271 ();
 sg13g2_fill_1 FILLER_16_1273 ();
 sg13g2_fill_2 FILLER_16_1284 ();
 sg13g2_decap_8 FILLER_16_1290 ();
 sg13g2_fill_2 FILLER_16_1327 ();
 sg13g2_decap_8 FILLER_16_1369 ();
 sg13g2_decap_8 FILLER_16_1376 ();
 sg13g2_decap_8 FILLER_16_1383 ();
 sg13g2_decap_8 FILLER_16_1404 ();
 sg13g2_decap_8 FILLER_16_1411 ();
 sg13g2_decap_8 FILLER_16_1418 ();
 sg13g2_decap_8 FILLER_16_1425 ();
 sg13g2_decap_8 FILLER_16_1432 ();
 sg13g2_fill_2 FILLER_16_1439 ();
 sg13g2_decap_4 FILLER_16_1451 ();
 sg13g2_fill_1 FILLER_16_1511 ();
 sg13g2_fill_1 FILLER_16_1541 ();
 sg13g2_fill_2 FILLER_16_1568 ();
 sg13g2_fill_1 FILLER_16_1570 ();
 sg13g2_fill_2 FILLER_16_1617 ();
 sg13g2_fill_1 FILLER_16_1619 ();
 sg13g2_decap_8 FILLER_16_1672 ();
 sg13g2_decap_8 FILLER_16_1679 ();
 sg13g2_fill_1 FILLER_16_1686 ();
 sg13g2_decap_8 FILLER_16_1691 ();
 sg13g2_decap_4 FILLER_16_1698 ();
 sg13g2_fill_2 FILLER_16_1702 ();
 sg13g2_fill_1 FILLER_16_1740 ();
 sg13g2_decap_8 FILLER_16_1767 ();
 sg13g2_decap_8 FILLER_17_26 ();
 sg13g2_fill_2 FILLER_17_33 ();
 sg13g2_fill_2 FILLER_17_66 ();
 sg13g2_fill_2 FILLER_17_94 ();
 sg13g2_decap_8 FILLER_17_117 ();
 sg13g2_decap_8 FILLER_17_124 ();
 sg13g2_decap_8 FILLER_17_131 ();
 sg13g2_decap_8 FILLER_17_138 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_209 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_313 ();
 sg13g2_fill_1 FILLER_17_320 ();
 sg13g2_decap_4 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_fill_1 FILLER_17_346 ();
 sg13g2_fill_2 FILLER_17_357 ();
 sg13g2_fill_2 FILLER_17_367 ();
 sg13g2_fill_1 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_fill_2 FILLER_17_403 ();
 sg13g2_fill_1 FILLER_17_431 ();
 sg13g2_fill_1 FILLER_17_436 ();
 sg13g2_fill_2 FILLER_17_447 ();
 sg13g2_decap_8 FILLER_17_453 ();
 sg13g2_fill_1 FILLER_17_460 ();
 sg13g2_fill_2 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_489 ();
 sg13g2_decap_8 FILLER_17_496 ();
 sg13g2_decap_4 FILLER_17_503 ();
 sg13g2_decap_4 FILLER_17_520 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_fill_1 FILLER_17_567 ();
 sg13g2_decap_4 FILLER_17_581 ();
 sg13g2_fill_2 FILLER_17_585 ();
 sg13g2_fill_1 FILLER_17_601 ();
 sg13g2_fill_2 FILLER_17_630 ();
 sg13g2_decap_4 FILLER_17_663 ();
 sg13g2_fill_2 FILLER_17_667 ();
 sg13g2_fill_1 FILLER_17_677 ();
 sg13g2_fill_1 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_713 ();
 sg13g2_fill_2 FILLER_17_720 ();
 sg13g2_fill_2 FILLER_17_748 ();
 sg13g2_fill_1 FILLER_17_750 ();
 sg13g2_decap_8 FILLER_17_809 ();
 sg13g2_decap_8 FILLER_17_816 ();
 sg13g2_decap_8 FILLER_17_823 ();
 sg13g2_decap_4 FILLER_17_830 ();
 sg13g2_fill_2 FILLER_17_834 ();
 sg13g2_decap_8 FILLER_17_849 ();
 sg13g2_decap_8 FILLER_17_856 ();
 sg13g2_decap_8 FILLER_17_863 ();
 sg13g2_decap_4 FILLER_17_870 ();
 sg13g2_fill_1 FILLER_17_874 ();
 sg13g2_decap_8 FILLER_17_888 ();
 sg13g2_fill_2 FILLER_17_895 ();
 sg13g2_fill_1 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_924 ();
 sg13g2_fill_2 FILLER_17_931 ();
 sg13g2_fill_1 FILLER_17_933 ();
 sg13g2_decap_8 FILLER_17_984 ();
 sg13g2_fill_2 FILLER_17_991 ();
 sg13g2_fill_2 FILLER_17_1003 ();
 sg13g2_fill_1 FILLER_17_1005 ();
 sg13g2_fill_2 FILLER_17_1010 ();
 sg13g2_fill_2 FILLER_17_1022 ();
 sg13g2_fill_1 FILLER_17_1024 ();
 sg13g2_decap_4 FILLER_17_1051 ();
 sg13g2_fill_2 FILLER_17_1055 ();
 sg13g2_decap_8 FILLER_17_1091 ();
 sg13g2_fill_2 FILLER_17_1098 ();
 sg13g2_fill_1 FILLER_17_1158 ();
 sg13g2_fill_1 FILLER_17_1169 ();
 sg13g2_fill_2 FILLER_17_1231 ();
 sg13g2_fill_1 FILLER_17_1233 ();
 sg13g2_decap_4 FILLER_17_1238 ();
 sg13g2_fill_2 FILLER_17_1242 ();
 sg13g2_fill_2 FILLER_17_1248 ();
 sg13g2_decap_8 FILLER_17_1317 ();
 sg13g2_fill_1 FILLER_17_1324 ();
 sg13g2_decap_8 FILLER_17_1365 ();
 sg13g2_decap_8 FILLER_17_1372 ();
 sg13g2_decap_8 FILLER_17_1379 ();
 sg13g2_decap_8 FILLER_17_1386 ();
 sg13g2_decap_4 FILLER_17_1393 ();
 sg13g2_fill_1 FILLER_17_1397 ();
 sg13g2_decap_8 FILLER_17_1448 ();
 sg13g2_decap_4 FILLER_17_1455 ();
 sg13g2_decap_8 FILLER_17_1469 ();
 sg13g2_fill_2 FILLER_17_1476 ();
 sg13g2_fill_1 FILLER_17_1478 ();
 sg13g2_fill_1 FILLER_17_1490 ();
 sg13g2_fill_1 FILLER_17_1501 ();
 sg13g2_fill_1 FILLER_17_1531 ();
 sg13g2_fill_1 FILLER_17_1535 ();
 sg13g2_fill_1 FILLER_17_1562 ();
 sg13g2_fill_1 FILLER_17_1588 ();
 sg13g2_fill_2 FILLER_17_1610 ();
 sg13g2_fill_1 FILLER_17_1642 ();
 sg13g2_decap_8 FILLER_17_1647 ();
 sg13g2_decap_8 FILLER_17_1654 ();
 sg13g2_decap_4 FILLER_17_1661 ();
 sg13g2_decap_4 FILLER_17_1675 ();
 sg13g2_fill_1 FILLER_17_1679 ();
 sg13g2_fill_2 FILLER_17_1745 ();
 sg13g2_fill_1 FILLER_17_1747 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_198 ();
 sg13g2_fill_2 FILLER_18_301 ();
 sg13g2_fill_1 FILLER_18_303 ();
 sg13g2_decap_4 FILLER_18_318 ();
 sg13g2_decap_4 FILLER_18_369 ();
 sg13g2_decap_4 FILLER_18_387 ();
 sg13g2_fill_1 FILLER_18_391 ();
 sg13g2_decap_4 FILLER_18_475 ();
 sg13g2_fill_1 FILLER_18_479 ();
 sg13g2_decap_8 FILLER_18_506 ();
 sg13g2_fill_2 FILLER_18_513 ();
 sg13g2_fill_2 FILLER_18_530 ();
 sg13g2_fill_1 FILLER_18_532 ();
 sg13g2_fill_1 FILLER_18_564 ();
 sg13g2_fill_2 FILLER_18_569 ();
 sg13g2_fill_1 FILLER_18_577 ();
 sg13g2_fill_2 FILLER_18_590 ();
 sg13g2_fill_2 FILLER_18_618 ();
 sg13g2_fill_1 FILLER_18_620 ();
 sg13g2_fill_1 FILLER_18_634 ();
 sg13g2_fill_2 FILLER_18_639 ();
 sg13g2_fill_2 FILLER_18_677 ();
 sg13g2_fill_1 FILLER_18_679 ();
 sg13g2_fill_1 FILLER_18_751 ();
 sg13g2_decap_8 FILLER_18_758 ();
 sg13g2_fill_2 FILLER_18_765 ();
 sg13g2_fill_1 FILLER_18_767 ();
 sg13g2_fill_2 FILLER_18_804 ();
 sg13g2_decap_8 FILLER_18_810 ();
 sg13g2_decap_8 FILLER_18_817 ();
 sg13g2_fill_1 FILLER_18_824 ();
 sg13g2_fill_2 FILLER_18_859 ();
 sg13g2_decap_4 FILLER_18_874 ();
 sg13g2_fill_2 FILLER_18_878 ();
 sg13g2_decap_4 FILLER_18_906 ();
 sg13g2_fill_1 FILLER_18_910 ();
 sg13g2_decap_8 FILLER_18_916 ();
 sg13g2_decap_8 FILLER_18_923 ();
 sg13g2_decap_8 FILLER_18_930 ();
 sg13g2_decap_8 FILLER_18_937 ();
 sg13g2_decap_4 FILLER_18_944 ();
 sg13g2_fill_1 FILLER_18_948 ();
 sg13g2_fill_2 FILLER_18_953 ();
 sg13g2_fill_1 FILLER_18_955 ();
 sg13g2_decap_4 FILLER_18_1002 ();
 sg13g2_fill_2 FILLER_18_1016 ();
 sg13g2_fill_1 FILLER_18_1018 ();
 sg13g2_fill_2 FILLER_18_1053 ();
 sg13g2_decap_8 FILLER_18_1063 ();
 sg13g2_fill_2 FILLER_18_1070 ();
 sg13g2_fill_2 FILLER_18_1076 ();
 sg13g2_fill_2 FILLER_18_1088 ();
 sg13g2_fill_2 FILLER_18_1094 ();
 sg13g2_fill_1 FILLER_18_1096 ();
 sg13g2_fill_1 FILLER_18_1110 ();
 sg13g2_decap_8 FILLER_18_1116 ();
 sg13g2_decap_4 FILLER_18_1123 ();
 sg13g2_fill_1 FILLER_18_1127 ();
 sg13g2_decap_4 FILLER_18_1134 ();
 sg13g2_fill_2 FILLER_18_1142 ();
 sg13g2_fill_2 FILLER_18_1165 ();
 sg13g2_fill_2 FILLER_18_1229 ();
 sg13g2_fill_2 FILLER_18_1241 ();
 sg13g2_fill_1 FILLER_18_1243 ();
 sg13g2_decap_4 FILLER_18_1249 ();
 sg13g2_fill_1 FILLER_18_1253 ();
 sg13g2_fill_2 FILLER_18_1265 ();
 sg13g2_fill_1 FILLER_18_1267 ();
 sg13g2_decap_8 FILLER_18_1304 ();
 sg13g2_decap_8 FILLER_18_1311 ();
 sg13g2_decap_8 FILLER_18_1318 ();
 sg13g2_fill_2 FILLER_18_1325 ();
 sg13g2_fill_1 FILLER_18_1337 ();
 sg13g2_fill_2 FILLER_18_1359 ();
 sg13g2_fill_1 FILLER_18_1387 ();
 sg13g2_fill_2 FILLER_18_1414 ();
 sg13g2_fill_1 FILLER_18_1456 ();
 sg13g2_fill_1 FILLER_18_1493 ();
 sg13g2_fill_1 FILLER_18_1511 ();
 sg13g2_fill_2 FILLER_18_1527 ();
 sg13g2_decap_8 FILLER_18_1570 ();
 sg13g2_decap_8 FILLER_18_1577 ();
 sg13g2_decap_8 FILLER_18_1584 ();
 sg13g2_fill_2 FILLER_18_1591 ();
 sg13g2_fill_1 FILLER_18_1593 ();
 sg13g2_decap_8 FILLER_18_1598 ();
 sg13g2_fill_2 FILLER_18_1605 ();
 sg13g2_decap_8 FILLER_18_1637 ();
 sg13g2_decap_8 FILLER_18_1644 ();
 sg13g2_decap_8 FILLER_18_1651 ();
 sg13g2_decap_4 FILLER_18_1658 ();
 sg13g2_fill_2 FILLER_18_1662 ();
 sg13g2_fill_1 FILLER_18_1669 ();
 sg13g2_fill_2 FILLER_18_1700 ();
 sg13g2_fill_1 FILLER_18_1702 ();
 sg13g2_fill_2 FILLER_18_1713 ();
 sg13g2_decap_4 FILLER_18_1739 ();
 sg13g2_fill_2 FILLER_18_1753 ();
 sg13g2_fill_1 FILLER_18_1755 ();
 sg13g2_decap_8 FILLER_18_1760 ();
 sg13g2_decap_8 FILLER_18_1767 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_12 ();
 sg13g2_fill_1 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_25 ();
 sg13g2_decap_4 FILLER_19_37 ();
 sg13g2_fill_2 FILLER_19_59 ();
 sg13g2_fill_2 FILLER_19_71 ();
 sg13g2_fill_2 FILLER_19_97 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_120 ();
 sg13g2_fill_2 FILLER_19_148 ();
 sg13g2_fill_1 FILLER_19_150 ();
 sg13g2_decap_4 FILLER_19_177 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_187 ();
 sg13g2_fill_2 FILLER_19_194 ();
 sg13g2_fill_2 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_fill_2 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_4 FILLER_19_377 ();
 sg13g2_fill_1 FILLER_19_381 ();
 sg13g2_fill_2 FILLER_19_447 ();
 sg13g2_fill_1 FILLER_19_449 ();
 sg13g2_fill_1 FILLER_19_476 ();
 sg13g2_decap_4 FILLER_19_491 ();
 sg13g2_decap_8 FILLER_19_499 ();
 sg13g2_decap_4 FILLER_19_506 ();
 sg13g2_fill_1 FILLER_19_510 ();
 sg13g2_fill_1 FILLER_19_537 ();
 sg13g2_fill_1 FILLER_19_542 ();
 sg13g2_fill_2 FILLER_19_547 ();
 sg13g2_fill_1 FILLER_19_570 ();
 sg13g2_fill_2 FILLER_19_577 ();
 sg13g2_fill_1 FILLER_19_595 ();
 sg13g2_fill_2 FILLER_19_632 ();
 sg13g2_fill_1 FILLER_19_634 ();
 sg13g2_fill_2 FILLER_19_654 ();
 sg13g2_decap_8 FILLER_19_660 ();
 sg13g2_decap_8 FILLER_19_667 ();
 sg13g2_fill_2 FILLER_19_674 ();
 sg13g2_fill_1 FILLER_19_710 ();
 sg13g2_fill_1 FILLER_19_715 ();
 sg13g2_fill_2 FILLER_19_774 ();
 sg13g2_fill_1 FILLER_19_776 ();
 sg13g2_fill_2 FILLER_19_782 ();
 sg13g2_fill_1 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_825 ();
 sg13g2_decap_4 FILLER_19_832 ();
 sg13g2_fill_2 FILLER_19_836 ();
 sg13g2_fill_2 FILLER_19_851 ();
 sg13g2_fill_1 FILLER_19_853 ();
 sg13g2_decap_4 FILLER_19_867 ();
 sg13g2_fill_2 FILLER_19_871 ();
 sg13g2_decap_4 FILLER_19_900 ();
 sg13g2_fill_1 FILLER_19_908 ();
 sg13g2_decap_8 FILLER_19_945 ();
 sg13g2_fill_2 FILLER_19_952 ();
 sg13g2_decap_8 FILLER_19_1054 ();
 sg13g2_decap_8 FILLER_19_1061 ();
 sg13g2_decap_8 FILLER_19_1068 ();
 sg13g2_fill_2 FILLER_19_1075 ();
 sg13g2_fill_1 FILLER_19_1103 ();
 sg13g2_decap_8 FILLER_19_1112 ();
 sg13g2_fill_1 FILLER_19_1119 ();
 sg13g2_fill_1 FILLER_19_1146 ();
 sg13g2_fill_1 FILLER_19_1177 ();
 sg13g2_fill_2 FILLER_19_1215 ();
 sg13g2_decap_4 FILLER_19_1254 ();
 sg13g2_fill_1 FILLER_19_1258 ();
 sg13g2_fill_1 FILLER_19_1269 ();
 sg13g2_fill_1 FILLER_19_1275 ();
 sg13g2_fill_1 FILLER_19_1280 ();
 sg13g2_fill_1 FILLER_19_1302 ();
 sg13g2_decap_4 FILLER_19_1355 ();
 sg13g2_fill_1 FILLER_19_1359 ();
 sg13g2_fill_2 FILLER_19_1369 ();
 sg13g2_fill_1 FILLER_19_1371 ();
 sg13g2_fill_2 FILLER_19_1376 ();
 sg13g2_decap_8 FILLER_19_1467 ();
 sg13g2_decap_4 FILLER_19_1474 ();
 sg13g2_fill_1 FILLER_19_1478 ();
 sg13g2_fill_2 FILLER_19_1493 ();
 sg13g2_fill_2 FILLER_19_1498 ();
 sg13g2_fill_1 FILLER_19_1541 ();
 sg13g2_fill_1 FILLER_19_1552 ();
 sg13g2_decap_4 FILLER_19_1579 ();
 sg13g2_decap_8 FILLER_19_1587 ();
 sg13g2_decap_8 FILLER_19_1594 ();
 sg13g2_decap_8 FILLER_19_1601 ();
 sg13g2_fill_2 FILLER_19_1608 ();
 sg13g2_fill_1 FILLER_19_1610 ();
 sg13g2_fill_2 FILLER_19_1649 ();
 sg13g2_fill_2 FILLER_19_1655 ();
 sg13g2_fill_1 FILLER_19_1657 ();
 sg13g2_decap_4 FILLER_19_1668 ();
 sg13g2_fill_2 FILLER_19_1672 ();
 sg13g2_decap_8 FILLER_19_1684 ();
 sg13g2_decap_4 FILLER_19_1691 ();
 sg13g2_decap_8 FILLER_19_1716 ();
 sg13g2_decap_8 FILLER_19_1723 ();
 sg13g2_decap_8 FILLER_19_1730 ();
 sg13g2_decap_8 FILLER_19_1767 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_4 FILLER_20_61 ();
 sg13g2_fill_2 FILLER_20_65 ();
 sg13g2_fill_1 FILLER_20_83 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_fill_2 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_146 ();
 sg13g2_fill_1 FILLER_20_157 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_230 ();
 sg13g2_decap_4 FILLER_20_294 ();
 sg13g2_fill_2 FILLER_20_298 ();
 sg13g2_fill_2 FILLER_20_340 ();
 sg13g2_fill_1 FILLER_20_342 ();
 sg13g2_fill_2 FILLER_20_383 ();
 sg13g2_decap_4 FILLER_20_395 ();
 sg13g2_decap_4 FILLER_20_409 ();
 sg13g2_fill_1 FILLER_20_423 ();
 sg13g2_fill_2 FILLER_20_450 ();
 sg13g2_fill_1 FILLER_20_452 ();
 sg13g2_decap_8 FILLER_20_478 ();
 sg13g2_decap_4 FILLER_20_485 ();
 sg13g2_fill_2 FILLER_20_515 ();
 sg13g2_fill_1 FILLER_20_517 ();
 sg13g2_decap_4 FILLER_20_522 ();
 sg13g2_fill_1 FILLER_20_526 ();
 sg13g2_fill_1 FILLER_20_537 ();
 sg13g2_fill_2 FILLER_20_564 ();
 sg13g2_fill_2 FILLER_20_576 ();
 sg13g2_fill_1 FILLER_20_578 ();
 sg13g2_fill_1 FILLER_20_591 ();
 sg13g2_fill_1 FILLER_20_597 ();
 sg13g2_fill_2 FILLER_20_606 ();
 sg13g2_fill_1 FILLER_20_608 ();
 sg13g2_decap_8 FILLER_20_621 ();
 sg13g2_fill_2 FILLER_20_628 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_4 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_673 ();
 sg13g2_decap_8 FILLER_20_680 ();
 sg13g2_decap_8 FILLER_20_691 ();
 sg13g2_decap_4 FILLER_20_698 ();
 sg13g2_fill_2 FILLER_20_702 ();
 sg13g2_decap_8 FILLER_20_718 ();
 sg13g2_fill_1 FILLER_20_725 ();
 sg13g2_fill_1 FILLER_20_776 ();
 sg13g2_decap_8 FILLER_20_803 ();
 sg13g2_decap_8 FILLER_20_810 ();
 sg13g2_fill_2 FILLER_20_817 ();
 sg13g2_fill_1 FILLER_20_844 ();
 sg13g2_fill_2 FILLER_20_858 ();
 sg13g2_decap_4 FILLER_20_890 ();
 sg13g2_fill_1 FILLER_20_894 ();
 sg13g2_decap_4 FILLER_20_931 ();
 sg13g2_decap_8 FILLER_20_939 ();
 sg13g2_decap_8 FILLER_20_946 ();
 sg13g2_fill_2 FILLER_20_953 ();
 sg13g2_fill_1 FILLER_20_999 ();
 sg13g2_decap_8 FILLER_20_1005 ();
 sg13g2_fill_2 FILLER_20_1012 ();
 sg13g2_decap_4 FILLER_20_1035 ();
 sg13g2_fill_1 FILLER_20_1039 ();
 sg13g2_fill_1 FILLER_20_1044 ();
 sg13g2_fill_2 FILLER_20_1057 ();
 sg13g2_decap_4 FILLER_20_1066 ();
 sg13g2_fill_2 FILLER_20_1096 ();
 sg13g2_fill_2 FILLER_20_1124 ();
 sg13g2_fill_1 FILLER_20_1126 ();
 sg13g2_fill_2 FILLER_20_1137 ();
 sg13g2_fill_1 FILLER_20_1139 ();
 sg13g2_fill_2 FILLER_20_1150 ();
 sg13g2_fill_2 FILLER_20_1160 ();
 sg13g2_fill_1 FILLER_20_1162 ();
 sg13g2_fill_1 FILLER_20_1200 ();
 sg13g2_fill_2 FILLER_20_1217 ();
 sg13g2_fill_1 FILLER_20_1229 ();
 sg13g2_fill_1 FILLER_20_1260 ();
 sg13g2_fill_1 FILLER_20_1313 ();
 sg13g2_decap_4 FILLER_20_1318 ();
 sg13g2_fill_2 FILLER_20_1322 ();
 sg13g2_decap_8 FILLER_20_1364 ();
 sg13g2_decap_8 FILLER_20_1371 ();
 sg13g2_decap_8 FILLER_20_1378 ();
 sg13g2_decap_4 FILLER_20_1385 ();
 sg13g2_fill_1 FILLER_20_1389 ();
 sg13g2_fill_1 FILLER_20_1435 ();
 sg13g2_decap_8 FILLER_20_1472 ();
 sg13g2_decap_8 FILLER_20_1479 ();
 sg13g2_fill_1 FILLER_20_1498 ();
 sg13g2_fill_1 FILLER_20_1528 ();
 sg13g2_fill_2 FILLER_20_1540 ();
 sg13g2_decap_4 FILLER_20_1553 ();
 sg13g2_decap_4 FILLER_20_1562 ();
 sg13g2_decap_8 FILLER_20_1602 ();
 sg13g2_fill_1 FILLER_20_1609 ();
 sg13g2_fill_2 FILLER_20_1618 ();
 sg13g2_decap_8 FILLER_20_1672 ();
 sg13g2_fill_1 FILLER_20_1679 ();
 sg13g2_decap_8 FILLER_20_1706 ();
 sg13g2_fill_2 FILLER_20_1713 ();
 sg13g2_fill_1 FILLER_20_1725 ();
 sg13g2_fill_1 FILLER_20_1752 ();
 sg13g2_decap_8 FILLER_20_1757 ();
 sg13g2_decap_8 FILLER_20_1764 ();
 sg13g2_fill_2 FILLER_20_1771 ();
 sg13g2_fill_1 FILLER_20_1773 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_9 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_16 ();
 sg13g2_fill_2 FILLER_21_47 ();
 sg13g2_fill_2 FILLER_21_59 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_fill_1 FILLER_21_78 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_114 ();
 sg13g2_decap_8 FILLER_21_121 ();
 sg13g2_decap_4 FILLER_21_128 ();
 sg13g2_fill_1 FILLER_21_132 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_4 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_decap_4 FILLER_21_190 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_decap_4 FILLER_21_206 ();
 sg13g2_fill_1 FILLER_21_210 ();
 sg13g2_decap_4 FILLER_21_215 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_fill_2 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_333 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_387 ();
 sg13g2_fill_2 FILLER_21_415 ();
 sg13g2_decap_4 FILLER_21_447 ();
 sg13g2_fill_2 FILLER_21_460 ();
 sg13g2_decap_4 FILLER_21_488 ();
 sg13g2_decap_4 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_509 ();
 sg13g2_decap_8 FILLER_21_516 ();
 sg13g2_decap_8 FILLER_21_523 ();
 sg13g2_fill_2 FILLER_21_530 ();
 sg13g2_decap_8 FILLER_21_542 ();
 sg13g2_decap_4 FILLER_21_549 ();
 sg13g2_fill_1 FILLER_21_553 ();
 sg13g2_fill_2 FILLER_21_600 ();
 sg13g2_decap_4 FILLER_21_632 ();
 sg13g2_fill_1 FILLER_21_639 ();
 sg13g2_decap_8 FILLER_21_666 ();
 sg13g2_decap_8 FILLER_21_673 ();
 sg13g2_decap_8 FILLER_21_680 ();
 sg13g2_decap_4 FILLER_21_687 ();
 sg13g2_fill_2 FILLER_21_727 ();
 sg13g2_fill_1 FILLER_21_729 ();
 sg13g2_decap_4 FILLER_21_736 ();
 sg13g2_decap_4 FILLER_21_776 ();
 sg13g2_fill_2 FILLER_21_780 ();
 sg13g2_decap_8 FILLER_21_790 ();
 sg13g2_decap_8 FILLER_21_797 ();
 sg13g2_fill_1 FILLER_21_804 ();
 sg13g2_decap_8 FILLER_21_813 ();
 sg13g2_decap_8 FILLER_21_820 ();
 sg13g2_decap_8 FILLER_21_827 ();
 sg13g2_decap_8 FILLER_21_834 ();
 sg13g2_decap_8 FILLER_21_841 ();
 sg13g2_decap_8 FILLER_21_848 ();
 sg13g2_fill_2 FILLER_21_855 ();
 sg13g2_decap_4 FILLER_21_877 ();
 sg13g2_fill_1 FILLER_21_907 ();
 sg13g2_fill_1 FILLER_21_928 ();
 sg13g2_decap_8 FILLER_21_941 ();
 sg13g2_decap_4 FILLER_21_948 ();
 sg13g2_fill_2 FILLER_21_952 ();
 sg13g2_decap_8 FILLER_21_958 ();
 sg13g2_decap_8 FILLER_21_965 ();
 sg13g2_decap_8 FILLER_21_972 ();
 sg13g2_decap_8 FILLER_21_979 ();
 sg13g2_decap_4 FILLER_21_986 ();
 sg13g2_fill_1 FILLER_21_990 ();
 sg13g2_decap_8 FILLER_21_995 ();
 sg13g2_decap_8 FILLER_21_1002 ();
 sg13g2_decap_8 FILLER_21_1009 ();
 sg13g2_decap_8 FILLER_21_1016 ();
 sg13g2_fill_2 FILLER_21_1023 ();
 sg13g2_decap_8 FILLER_21_1034 ();
 sg13g2_fill_1 FILLER_21_1041 ();
 sg13g2_fill_1 FILLER_21_1053 ();
 sg13g2_decap_8 FILLER_21_1058 ();
 sg13g2_decap_4 FILLER_21_1065 ();
 sg13g2_fill_1 FILLER_21_1079 ();
 sg13g2_decap_4 FILLER_21_1108 ();
 sg13g2_decap_4 FILLER_21_1116 ();
 sg13g2_fill_2 FILLER_21_1124 ();
 sg13g2_fill_2 FILLER_21_1165 ();
 sg13g2_fill_1 FILLER_21_1167 ();
 sg13g2_fill_1 FILLER_21_1197 ();
 sg13g2_fill_1 FILLER_21_1216 ();
 sg13g2_fill_2 FILLER_21_1292 ();
 sg13g2_fill_1 FILLER_21_1294 ();
 sg13g2_decap_8 FILLER_21_1309 ();
 sg13g2_decap_8 FILLER_21_1316 ();
 sg13g2_decap_8 FILLER_21_1323 ();
 sg13g2_fill_2 FILLER_21_1330 ();
 sg13g2_fill_1 FILLER_21_1342 ();
 sg13g2_fill_2 FILLER_21_1384 ();
 sg13g2_fill_2 FILLER_21_1402 ();
 sg13g2_decap_4 FILLER_21_1433 ();
 sg13g2_fill_1 FILLER_21_1437 ();
 sg13g2_fill_2 FILLER_21_1446 ();
 sg13g2_fill_2 FILLER_21_1457 ();
 sg13g2_fill_1 FILLER_21_1459 ();
 sg13g2_fill_1 FILLER_21_1491 ();
 sg13g2_fill_1 FILLER_21_1498 ();
 sg13g2_fill_1 FILLER_21_1504 ();
 sg13g2_fill_2 FILLER_21_1515 ();
 sg13g2_fill_1 FILLER_21_1517 ();
 sg13g2_decap_4 FILLER_21_1523 ();
 sg13g2_fill_1 FILLER_21_1527 ();
 sg13g2_decap_8 FILLER_21_1546 ();
 sg13g2_decap_8 FILLER_21_1553 ();
 sg13g2_fill_2 FILLER_21_1560 ();
 sg13g2_fill_2 FILLER_21_1587 ();
 sg13g2_fill_1 FILLER_21_1589 ();
 sg13g2_fill_2 FILLER_21_1595 ();
 sg13g2_fill_1 FILLER_21_1597 ();
 sg13g2_fill_1 FILLER_21_1608 ();
 sg13g2_fill_1 FILLER_21_1635 ();
 sg13g2_fill_1 FILLER_21_1662 ();
 sg13g2_decap_8 FILLER_21_1759 ();
 sg13g2_decap_8 FILLER_21_1766 ();
 sg13g2_fill_1 FILLER_21_1773 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_40 ();
 sg13g2_fill_2 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_82 ();
 sg13g2_fill_1 FILLER_22_115 ();
 sg13g2_fill_2 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_290 ();
 sg13g2_decap_8 FILLER_22_297 ();
 sg13g2_decap_8 FILLER_22_304 ();
 sg13g2_decap_8 FILLER_22_311 ();
 sg13g2_decap_8 FILLER_22_318 ();
 sg13g2_decap_4 FILLER_22_325 ();
 sg13g2_fill_1 FILLER_22_329 ();
 sg13g2_decap_4 FILLER_22_334 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_decap_8 FILLER_22_438 ();
 sg13g2_decap_8 FILLER_22_445 ();
 sg13g2_decap_4 FILLER_22_452 ();
 sg13g2_fill_2 FILLER_22_521 ();
 sg13g2_fill_1 FILLER_22_533 ();
 sg13g2_fill_2 FILLER_22_570 ();
 sg13g2_fill_2 FILLER_22_598 ();
 sg13g2_fill_1 FILLER_22_600 ();
 sg13g2_fill_2 FILLER_22_655 ();
 sg13g2_fill_2 FILLER_22_688 ();
 sg13g2_fill_1 FILLER_22_726 ();
 sg13g2_fill_2 FILLER_22_735 ();
 sg13g2_fill_1 FILLER_22_758 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_775 ();
 sg13g2_decap_8 FILLER_22_782 ();
 sg13g2_fill_1 FILLER_22_789 ();
 sg13g2_decap_8 FILLER_22_803 ();
 sg13g2_fill_1 FILLER_22_853 ();
 sg13g2_fill_1 FILLER_22_864 ();
 sg13g2_fill_1 FILLER_22_869 ();
 sg13g2_fill_1 FILLER_22_880 ();
 sg13g2_fill_1 FILLER_22_891 ();
 sg13g2_decap_8 FILLER_22_938 ();
 sg13g2_decap_8 FILLER_22_1001 ();
 sg13g2_fill_1 FILLER_22_1012 ();
 sg13g2_decap_8 FILLER_22_1039 ();
 sg13g2_decap_8 FILLER_22_1046 ();
 sg13g2_decap_8 FILLER_22_1053 ();
 sg13g2_fill_2 FILLER_22_1060 ();
 sg13g2_fill_1 FILLER_22_1062 ();
 sg13g2_decap_8 FILLER_22_1103 ();
 sg13g2_fill_2 FILLER_22_1110 ();
 sg13g2_decap_4 FILLER_22_1122 ();
 sg13g2_fill_1 FILLER_22_1169 ();
 sg13g2_decap_4 FILLER_22_1185 ();
 sg13g2_decap_4 FILLER_22_1202 ();
 sg13g2_decap_4 FILLER_22_1232 ();
 sg13g2_fill_2 FILLER_22_1246 ();
 sg13g2_decap_8 FILLER_22_1276 ();
 sg13g2_decap_8 FILLER_22_1283 ();
 sg13g2_decap_4 FILLER_22_1290 ();
 sg13g2_fill_1 FILLER_22_1294 ();
 sg13g2_fill_2 FILLER_22_1305 ();
 sg13g2_decap_4 FILLER_22_1317 ();
 sg13g2_fill_1 FILLER_22_1321 ();
 sg13g2_decap_8 FILLER_22_1326 ();
 sg13g2_decap_4 FILLER_22_1354 ();
 sg13g2_fill_2 FILLER_22_1358 ();
 sg13g2_decap_8 FILLER_22_1364 ();
 sg13g2_decap_8 FILLER_22_1375 ();
 sg13g2_decap_8 FILLER_22_1382 ();
 sg13g2_fill_1 FILLER_22_1401 ();
 sg13g2_fill_2 FILLER_22_1432 ();
 sg13g2_fill_1 FILLER_22_1434 ();
 sg13g2_decap_4 FILLER_22_1445 ();
 sg13g2_fill_2 FILLER_22_1479 ();
 sg13g2_fill_1 FILLER_22_1507 ();
 sg13g2_fill_2 FILLER_22_1516 ();
 sg13g2_fill_1 FILLER_22_1518 ();
 sg13g2_decap_8 FILLER_22_1573 ();
 sg13g2_decap_8 FILLER_22_1580 ();
 sg13g2_decap_4 FILLER_22_1587 ();
 sg13g2_fill_2 FILLER_22_1591 ();
 sg13g2_fill_1 FILLER_22_1611 ();
 sg13g2_fill_2 FILLER_22_1626 ();
 sg13g2_decap_8 FILLER_22_1632 ();
 sg13g2_fill_1 FILLER_22_1639 ();
 sg13g2_decap_4 FILLER_22_1648 ();
 sg13g2_fill_1 FILLER_22_1726 ();
 sg13g2_decap_8 FILLER_22_1767 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_27 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_113 ();
 sg13g2_fill_1 FILLER_23_141 ();
 sg13g2_fill_1 FILLER_23_168 ();
 sg13g2_fill_1 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_200 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_264 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_fill_2 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_decap_8 FILLER_23_407 ();
 sg13g2_decap_4 FILLER_23_414 ();
 sg13g2_fill_1 FILLER_23_418 ();
 sg13g2_decap_4 FILLER_23_423 ();
 sg13g2_fill_1 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_432 ();
 sg13g2_decap_4 FILLER_23_439 ();
 sg13g2_fill_2 FILLER_23_443 ();
 sg13g2_decap_4 FILLER_23_473 ();
 sg13g2_fill_2 FILLER_23_477 ();
 sg13g2_fill_1 FILLER_23_517 ();
 sg13g2_fill_2 FILLER_23_539 ();
 sg13g2_fill_1 FILLER_23_545 ();
 sg13g2_decap_4 FILLER_23_563 ();
 sg13g2_fill_1 FILLER_23_567 ();
 sg13g2_fill_2 FILLER_23_578 ();
 sg13g2_fill_1 FILLER_23_642 ();
 sg13g2_decap_4 FILLER_23_656 ();
 sg13g2_fill_2 FILLER_23_660 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_fill_2 FILLER_23_679 ();
 sg13g2_decap_4 FILLER_23_742 ();
 sg13g2_fill_1 FILLER_23_746 ();
 sg13g2_fill_1 FILLER_23_751 ();
 sg13g2_fill_2 FILLER_23_761 ();
 sg13g2_fill_2 FILLER_23_796 ();
 sg13g2_decap_4 FILLER_23_811 ();
 sg13g2_fill_1 FILLER_23_815 ();
 sg13g2_decap_4 FILLER_23_829 ();
 sg13g2_fill_2 FILLER_23_843 ();
 sg13g2_fill_2 FILLER_23_871 ();
 sg13g2_decap_8 FILLER_23_899 ();
 sg13g2_fill_2 FILLER_23_906 ();
 sg13g2_fill_2 FILLER_23_911 ();
 sg13g2_decap_8 FILLER_23_953 ();
 sg13g2_fill_1 FILLER_23_964 ();
 sg13g2_decap_8 FILLER_23_991 ();
 sg13g2_decap_4 FILLER_23_998 ();
 sg13g2_fill_1 FILLER_23_1002 ();
 sg13g2_decap_8 FILLER_23_1059 ();
 sg13g2_fill_1 FILLER_23_1066 ();
 sg13g2_decap_8 FILLER_23_1071 ();
 sg13g2_decap_4 FILLER_23_1082 ();
 sg13g2_fill_2 FILLER_23_1086 ();
 sg13g2_fill_2 FILLER_23_1140 ();
 sg13g2_fill_1 FILLER_23_1142 ();
 sg13g2_decap_8 FILLER_23_1194 ();
 sg13g2_decap_4 FILLER_23_1201 ();
 sg13g2_fill_1 FILLER_23_1205 ();
 sg13g2_fill_1 FILLER_23_1242 ();
 sg13g2_fill_1 FILLER_23_1253 ();
 sg13g2_fill_2 FILLER_23_1262 ();
 sg13g2_fill_1 FILLER_23_1314 ();
 sg13g2_decap_8 FILLER_23_1351 ();
 sg13g2_decap_8 FILLER_23_1358 ();
 sg13g2_fill_2 FILLER_23_1365 ();
 sg13g2_decap_8 FILLER_23_1371 ();
 sg13g2_fill_2 FILLER_23_1378 ();
 sg13g2_fill_1 FILLER_23_1380 ();
 sg13g2_fill_2 FILLER_23_1394 ();
 sg13g2_decap_4 FILLER_23_1422 ();
 sg13g2_decap_8 FILLER_23_1436 ();
 sg13g2_decap_8 FILLER_23_1469 ();
 sg13g2_decap_8 FILLER_23_1476 ();
 sg13g2_decap_8 FILLER_23_1483 ();
 sg13g2_decap_4 FILLER_23_1494 ();
 sg13g2_fill_1 FILLER_23_1498 ();
 sg13g2_fill_2 FILLER_23_1509 ();
 sg13g2_fill_2 FILLER_23_1537 ();
 sg13g2_fill_1 FILLER_23_1539 ();
 sg13g2_fill_1 FILLER_23_1566 ();
 sg13g2_fill_2 FILLER_23_1571 ();
 sg13g2_fill_1 FILLER_23_1573 ();
 sg13g2_decap_8 FILLER_23_1624 ();
 sg13g2_decap_8 FILLER_23_1631 ();
 sg13g2_decap_8 FILLER_23_1638 ();
 sg13g2_decap_8 FILLER_23_1645 ();
 sg13g2_decap_8 FILLER_23_1652 ();
 sg13g2_decap_8 FILLER_23_1659 ();
 sg13g2_decap_8 FILLER_23_1666 ();
 sg13g2_decap_4 FILLER_23_1673 ();
 sg13g2_fill_2 FILLER_23_1677 ();
 sg13g2_fill_1 FILLER_23_1689 ();
 sg13g2_decap_4 FILLER_23_1694 ();
 sg13g2_decap_8 FILLER_23_1702 ();
 sg13g2_decap_4 FILLER_23_1709 ();
 sg13g2_fill_2 FILLER_23_1713 ();
 sg13g2_decap_8 FILLER_23_1725 ();
 sg13g2_decap_8 FILLER_23_1732 ();
 sg13g2_decap_8 FILLER_23_1739 ();
 sg13g2_decap_8 FILLER_23_1746 ();
 sg13g2_decap_8 FILLER_23_1753 ();
 sg13g2_decap_8 FILLER_23_1760 ();
 sg13g2_decap_8 FILLER_23_1767 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_9 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_132 ();
 sg13g2_decap_4 FILLER_24_146 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_1 FILLER_24_201 ();
 sg13g2_fill_2 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_268 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_fill_2 FILLER_24_303 ();
 sg13g2_decap_4 FILLER_24_318 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_337 ();
 sg13g2_fill_1 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_365 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_415 ();
 sg13g2_decap_8 FILLER_24_422 ();
 sg13g2_decap_8 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_24_436 ();
 sg13g2_decap_8 FILLER_24_443 ();
 sg13g2_decap_8 FILLER_24_450 ();
 sg13g2_decap_8 FILLER_24_457 ();
 sg13g2_decap_4 FILLER_24_464 ();
 sg13g2_fill_1 FILLER_24_468 ();
 sg13g2_decap_4 FILLER_24_482 ();
 sg13g2_fill_2 FILLER_24_486 ();
 sg13g2_decap_4 FILLER_24_498 ();
 sg13g2_fill_2 FILLER_24_528 ();
 sg13g2_decap_4 FILLER_24_551 ();
 sg13g2_fill_2 FILLER_24_568 ();
 sg13g2_fill_1 FILLER_24_570 ();
 sg13g2_decap_8 FILLER_24_601 ();
 sg13g2_decap_8 FILLER_24_608 ();
 sg13g2_fill_2 FILLER_24_615 ();
 sg13g2_fill_1 FILLER_24_617 ();
 sg13g2_fill_2 FILLER_24_625 ();
 sg13g2_decap_8 FILLER_24_646 ();
 sg13g2_decap_8 FILLER_24_653 ();
 sg13g2_decap_8 FILLER_24_660 ();
 sg13g2_decap_8 FILLER_24_667 ();
 sg13g2_decap_4 FILLER_24_674 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_fill_1 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_741 ();
 sg13g2_fill_2 FILLER_24_748 ();
 sg13g2_fill_1 FILLER_24_750 ();
 sg13g2_decap_4 FILLER_24_756 ();
 sg13g2_decap_4 FILLER_24_764 ();
 sg13g2_fill_2 FILLER_24_768 ();
 sg13g2_fill_1 FILLER_24_775 ();
 sg13g2_decap_4 FILLER_24_789 ();
 sg13g2_fill_2 FILLER_24_806 ();
 sg13g2_fill_1 FILLER_24_808 ();
 sg13g2_decap_8 FILLER_24_822 ();
 sg13g2_decap_4 FILLER_24_829 ();
 sg13g2_fill_1 FILLER_24_833 ();
 sg13g2_fill_2 FILLER_24_844 ();
 sg13g2_fill_1 FILLER_24_846 ();
 sg13g2_decap_4 FILLER_24_860 ();
 sg13g2_fill_1 FILLER_24_864 ();
 sg13g2_decap_8 FILLER_24_895 ();
 sg13g2_fill_2 FILLER_24_902 ();
 sg13g2_fill_1 FILLER_24_904 ();
 sg13g2_decap_4 FILLER_24_938 ();
 sg13g2_fill_2 FILLER_24_942 ();
 sg13g2_decap_4 FILLER_24_952 ();
 sg13g2_fill_2 FILLER_24_1038 ();
 sg13g2_fill_2 FILLER_24_1044 ();
 sg13g2_fill_1 FILLER_24_1046 ();
 sg13g2_decap_8 FILLER_24_1073 ();
 sg13g2_decap_8 FILLER_24_1080 ();
 sg13g2_decap_8 FILLER_24_1087 ();
 sg13g2_fill_2 FILLER_24_1094 ();
 sg13g2_fill_1 FILLER_24_1122 ();
 sg13g2_fill_1 FILLER_24_1127 ();
 sg13g2_fill_1 FILLER_24_1149 ();
 sg13g2_fill_2 FILLER_24_1168 ();
 sg13g2_fill_2 FILLER_24_1206 ();
 sg13g2_fill_1 FILLER_24_1208 ();
 sg13g2_fill_1 FILLER_24_1217 ();
 sg13g2_fill_2 FILLER_24_1222 ();
 sg13g2_fill_2 FILLER_24_1234 ();
 sg13g2_decap_8 FILLER_24_1292 ();
 sg13g2_decap_8 FILLER_24_1299 ();
 sg13g2_decap_4 FILLER_24_1306 ();
 sg13g2_fill_1 FILLER_24_1310 ();
 sg13g2_fill_2 FILLER_24_1347 ();
 sg13g2_fill_1 FILLER_24_1349 ();
 sg13g2_decap_8 FILLER_24_1376 ();
 sg13g2_decap_4 FILLER_24_1383 ();
 sg13g2_fill_1 FILLER_24_1387 ();
 sg13g2_decap_8 FILLER_24_1412 ();
 sg13g2_decap_4 FILLER_24_1419 ();
 sg13g2_fill_2 FILLER_24_1423 ();
 sg13g2_decap_8 FILLER_24_1455 ();
 sg13g2_decap_8 FILLER_24_1462 ();
 sg13g2_decap_8 FILLER_24_1469 ();
 sg13g2_decap_8 FILLER_24_1476 ();
 sg13g2_decap_8 FILLER_24_1483 ();
 sg13g2_decap_4 FILLER_24_1490 ();
 sg13g2_fill_1 FILLER_24_1515 ();
 sg13g2_fill_1 FILLER_24_1520 ();
 sg13g2_fill_2 FILLER_24_1531 ();
 sg13g2_fill_1 FILLER_24_1537 ();
 sg13g2_fill_1 FILLER_24_1543 ();
 sg13g2_fill_1 FILLER_24_1548 ();
 sg13g2_fill_2 FILLER_24_1559 ();
 sg13g2_decap_4 FILLER_24_1587 ();
 sg13g2_decap_4 FILLER_24_1617 ();
 sg13g2_fill_2 FILLER_24_1621 ();
 sg13g2_decap_8 FILLER_24_1631 ();
 sg13g2_decap_8 FILLER_24_1638 ();
 sg13g2_decap_8 FILLER_24_1645 ();
 sg13g2_fill_1 FILLER_24_1652 ();
 sg13g2_fill_2 FILLER_24_1663 ();
 sg13g2_fill_1 FILLER_24_1665 ();
 sg13g2_decap_8 FILLER_24_1702 ();
 sg13g2_decap_8 FILLER_24_1709 ();
 sg13g2_decap_8 FILLER_24_1716 ();
 sg13g2_decap_8 FILLER_24_1723 ();
 sg13g2_decap_4 FILLER_24_1730 ();
 sg13g2_fill_2 FILLER_24_1734 ();
 sg13g2_fill_1 FILLER_24_1740 ();
 sg13g2_decap_8 FILLER_24_1767 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_22 ();
 sg13g2_fill_1 FILLER_25_48 ();
 sg13g2_decap_4 FILLER_25_53 ();
 sg13g2_fill_2 FILLER_25_67 ();
 sg13g2_fill_2 FILLER_25_89 ();
 sg13g2_fill_2 FILLER_25_127 ();
 sg13g2_fill_1 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_174 ();
 sg13g2_decap_8 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_201 ();
 sg13g2_decap_8 FILLER_25_212 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_decap_4 FILLER_25_226 ();
 sg13g2_fill_1 FILLER_25_230 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_4 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_fill_2 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_4 FILLER_25_331 ();
 sg13g2_fill_1 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_414 ();
 sg13g2_decap_8 FILLER_25_421 ();
 sg13g2_decap_8 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_25_435 ();
 sg13g2_decap_8 FILLER_25_442 ();
 sg13g2_decap_8 FILLER_25_449 ();
 sg13g2_decap_8 FILLER_25_456 ();
 sg13g2_decap_8 FILLER_25_463 ();
 sg13g2_fill_2 FILLER_25_470 ();
 sg13g2_fill_2 FILLER_25_498 ();
 sg13g2_decap_8 FILLER_25_531 ();
 sg13g2_decap_4 FILLER_25_538 ();
 sg13g2_fill_2 FILLER_25_542 ();
 sg13g2_decap_4 FILLER_25_570 ();
 sg13g2_fill_1 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_589 ();
 sg13g2_fill_1 FILLER_25_596 ();
 sg13g2_decap_8 FILLER_25_607 ();
 sg13g2_decap_8 FILLER_25_614 ();
 sg13g2_decap_4 FILLER_25_621 ();
 sg13g2_fill_2 FILLER_25_625 ();
 sg13g2_decap_4 FILLER_25_630 ();
 sg13g2_fill_1 FILLER_25_634 ();
 sg13g2_decap_8 FILLER_25_643 ();
 sg13g2_decap_4 FILLER_25_650 ();
 sg13g2_decap_8 FILLER_25_664 ();
 sg13g2_decap_8 FILLER_25_671 ();
 sg13g2_decap_8 FILLER_25_678 ();
 sg13g2_decap_8 FILLER_25_685 ();
 sg13g2_decap_8 FILLER_25_692 ();
 sg13g2_decap_8 FILLER_25_699 ();
 sg13g2_fill_2 FILLER_25_706 ();
 sg13g2_decap_4 FILLER_25_712 ();
 sg13g2_fill_1 FILLER_25_716 ();
 sg13g2_decap_8 FILLER_25_740 ();
 sg13g2_decap_4 FILLER_25_757 ();
 sg13g2_fill_1 FILLER_25_765 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_fill_2 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_801 ();
 sg13g2_decap_8 FILLER_25_808 ();
 sg13g2_fill_2 FILLER_25_815 ();
 sg13g2_fill_1 FILLER_25_817 ();
 sg13g2_decap_4 FILLER_25_831 ();
 sg13g2_fill_1 FILLER_25_838 ();
 sg13g2_decap_8 FILLER_25_856 ();
 sg13g2_decap_4 FILLER_25_863 ();
 sg13g2_fill_2 FILLER_25_867 ();
 sg13g2_fill_1 FILLER_25_879 ();
 sg13g2_fill_2 FILLER_25_884 ();
 sg13g2_decap_8 FILLER_25_890 ();
 sg13g2_fill_2 FILLER_25_941 ();
 sg13g2_fill_1 FILLER_25_973 ();
 sg13g2_fill_1 FILLER_25_1004 ();
 sg13g2_decap_8 FILLER_25_1015 ();
 sg13g2_fill_2 FILLER_25_1022 ();
 sg13g2_decap_8 FILLER_25_1028 ();
 sg13g2_decap_8 FILLER_25_1035 ();
 sg13g2_fill_1 FILLER_25_1042 ();
 sg13g2_fill_2 FILLER_25_1057 ();
 sg13g2_decap_8 FILLER_25_1076 ();
 sg13g2_decap_8 FILLER_25_1083 ();
 sg13g2_decap_4 FILLER_25_1090 ();
 sg13g2_fill_2 FILLER_25_1094 ();
 sg13g2_decap_4 FILLER_25_1100 ();
 sg13g2_fill_1 FILLER_25_1120 ();
 sg13g2_fill_2 FILLER_25_1151 ();
 sg13g2_decap_8 FILLER_25_1202 ();
 sg13g2_decap_4 FILLER_25_1209 ();
 sg13g2_fill_1 FILLER_25_1234 ();
 sg13g2_fill_2 FILLER_25_1261 ();
 sg13g2_fill_2 FILLER_25_1273 ();
 sg13g2_fill_2 FILLER_25_1279 ();
 sg13g2_decap_8 FILLER_25_1285 ();
 sg13g2_decap_4 FILLER_25_1292 ();
 sg13g2_decap_8 FILLER_25_1300 ();
 sg13g2_fill_2 FILLER_25_1307 ();
 sg13g2_fill_1 FILLER_25_1309 ();
 sg13g2_fill_2 FILLER_25_1340 ();
 sg13g2_fill_1 FILLER_25_1342 ();
 sg13g2_decap_8 FILLER_25_1383 ();
 sg13g2_fill_1 FILLER_25_1390 ();
 sg13g2_decap_8 FILLER_25_1395 ();
 sg13g2_decap_8 FILLER_25_1402 ();
 sg13g2_decap_8 FILLER_25_1409 ();
 sg13g2_decap_8 FILLER_25_1416 ();
 sg13g2_decap_8 FILLER_25_1423 ();
 sg13g2_decap_4 FILLER_25_1434 ();
 sg13g2_fill_2 FILLER_25_1438 ();
 sg13g2_decap_8 FILLER_25_1461 ();
 sg13g2_fill_2 FILLER_25_1468 ();
 sg13g2_decap_8 FILLER_25_1480 ();
 sg13g2_fill_2 FILLER_25_1487 ();
 sg13g2_decap_4 FILLER_25_1525 ();
 sg13g2_fill_2 FILLER_25_1529 ();
 sg13g2_decap_8 FILLER_25_1567 ();
 sg13g2_decap_8 FILLER_25_1574 ();
 sg13g2_fill_1 FILLER_25_1581 ();
 sg13g2_decap_8 FILLER_25_1586 ();
 sg13g2_decap_4 FILLER_25_1593 ();
 sg13g2_fill_2 FILLER_25_1597 ();
 sg13g2_decap_8 FILLER_25_1629 ();
 sg13g2_decap_8 FILLER_25_1636 ();
 sg13g2_decap_4 FILLER_25_1643 ();
 sg13g2_fill_2 FILLER_25_1673 ();
 sg13g2_fill_1 FILLER_25_1727 ();
 sg13g2_fill_2 FILLER_25_1768 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_44 ();
 sg13g2_decap_8 FILLER_26_51 ();
 sg13g2_decap_8 FILLER_26_58 ();
 sg13g2_decap_8 FILLER_26_65 ();
 sg13g2_decap_4 FILLER_26_72 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_decap_4 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_96 ();
 sg13g2_decap_8 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_108 ();
 sg13g2_decap_8 FILLER_26_115 ();
 sg13g2_fill_2 FILLER_26_122 ();
 sg13g2_fill_1 FILLER_26_124 ();
 sg13g2_decap_4 FILLER_26_138 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_fill_1 FILLER_26_243 ();
 sg13g2_fill_2 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_decap_8 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_331 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_decap_4 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_365 ();
 sg13g2_fill_2 FILLER_26_393 ();
 sg13g2_fill_1 FILLER_26_395 ();
 sg13g2_fill_2 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_424 ();
 sg13g2_fill_2 FILLER_26_451 ();
 sg13g2_fill_1 FILLER_26_453 ();
 sg13g2_fill_2 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_496 ();
 sg13g2_decap_8 FILLER_26_503 ();
 sg13g2_decap_8 FILLER_26_510 ();
 sg13g2_decap_8 FILLER_26_517 ();
 sg13g2_decap_8 FILLER_26_524 ();
 sg13g2_decap_8 FILLER_26_531 ();
 sg13g2_decap_8 FILLER_26_538 ();
 sg13g2_fill_2 FILLER_26_545 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_fill_2 FILLER_26_595 ();
 sg13g2_fill_1 FILLER_26_597 ();
 sg13g2_decap_8 FILLER_26_624 ();
 sg13g2_decap_8 FILLER_26_661 ();
 sg13g2_decap_8 FILLER_26_682 ();
 sg13g2_decap_8 FILLER_26_689 ();
 sg13g2_fill_1 FILLER_26_696 ();
 sg13g2_decap_8 FILLER_26_788 ();
 sg13g2_decap_8 FILLER_26_795 ();
 sg13g2_decap_8 FILLER_26_802 ();
 sg13g2_decap_8 FILLER_26_809 ();
 sg13g2_decap_4 FILLER_26_816 ();
 sg13g2_fill_2 FILLER_26_820 ();
 sg13g2_fill_1 FILLER_26_857 ();
 sg13g2_decap_8 FILLER_26_905 ();
 sg13g2_decap_8 FILLER_26_912 ();
 sg13g2_decap_4 FILLER_26_919 ();
 sg13g2_fill_1 FILLER_26_923 ();
 sg13g2_decap_8 FILLER_26_934 ();
 sg13g2_decap_8 FILLER_26_941 ();
 sg13g2_decap_4 FILLER_26_948 ();
 sg13g2_fill_1 FILLER_26_952 ();
 sg13g2_fill_2 FILLER_26_1002 ();
 sg13g2_fill_2 FILLER_26_1014 ();
 sg13g2_decap_8 FILLER_26_1078 ();
 sg13g2_fill_1 FILLER_26_1085 ();
 sg13g2_fill_1 FILLER_26_1104 ();
 sg13g2_decap_8 FILLER_26_1115 ();
 sg13g2_fill_2 FILLER_26_1122 ();
 sg13g2_fill_1 FILLER_26_1124 ();
 sg13g2_fill_1 FILLER_26_1135 ();
 sg13g2_fill_1 FILLER_26_1146 ();
 sg13g2_fill_2 FILLER_26_1153 ();
 sg13g2_fill_1 FILLER_26_1155 ();
 sg13g2_decap_8 FILLER_26_1180 ();
 sg13g2_decap_4 FILLER_26_1187 ();
 sg13g2_fill_1 FILLER_26_1191 ();
 sg13g2_decap_4 FILLER_26_1218 ();
 sg13g2_fill_1 FILLER_26_1222 ();
 sg13g2_fill_2 FILLER_26_1244 ();
 sg13g2_fill_1 FILLER_26_1250 ();
 sg13g2_decap_8 FILLER_26_1259 ();
 sg13g2_decap_8 FILLER_26_1266 ();
 sg13g2_decap_8 FILLER_26_1273 ();
 sg13g2_decap_8 FILLER_26_1280 ();
 sg13g2_fill_2 FILLER_26_1287 ();
 sg13g2_decap_8 FILLER_26_1315 ();
 sg13g2_fill_2 FILLER_26_1322 ();
 sg13g2_fill_2 FILLER_26_1345 ();
 sg13g2_fill_1 FILLER_26_1347 ();
 sg13g2_decap_8 FILLER_26_1374 ();
 sg13g2_fill_2 FILLER_26_1381 ();
 sg13g2_fill_1 FILLER_26_1383 ();
 sg13g2_decap_8 FILLER_26_1414 ();
 sg13g2_decap_8 FILLER_26_1421 ();
 sg13g2_decap_8 FILLER_26_1428 ();
 sg13g2_decap_8 FILLER_26_1435 ();
 sg13g2_decap_4 FILLER_26_1514 ();
 sg13g2_fill_1 FILLER_26_1518 ();
 sg13g2_decap_8 FILLER_26_1523 ();
 sg13g2_decap_8 FILLER_26_1530 ();
 sg13g2_fill_1 FILLER_26_1537 ();
 sg13g2_fill_2 FILLER_26_1584 ();
 sg13g2_decap_8 FILLER_26_1616 ();
 sg13g2_decap_8 FILLER_26_1623 ();
 sg13g2_decap_4 FILLER_26_1630 ();
 sg13g2_fill_2 FILLER_26_1690 ();
 sg13g2_fill_1 FILLER_26_1692 ();
 sg13g2_decap_8 FILLER_26_1765 ();
 sg13g2_fill_2 FILLER_26_1772 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_18 ();
 sg13g2_decap_8 FILLER_27_24 ();
 sg13g2_fill_2 FILLER_27_31 ();
 sg13g2_fill_1 FILLER_27_43 ();
 sg13g2_decap_8 FILLER_27_96 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_decap_8 FILLER_27_110 ();
 sg13g2_fill_1 FILLER_27_117 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_151 ();
 sg13g2_decap_8 FILLER_27_157 ();
 sg13g2_decap_8 FILLER_27_164 ();
 sg13g2_decap_4 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_fill_1 FILLER_27_255 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_decap_4 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_fill_2 FILLER_27_288 ();
 sg13g2_decap_4 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_fill_2 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_fill_1 FILLER_27_404 ();
 sg13g2_fill_2 FILLER_27_409 ();
 sg13g2_fill_1 FILLER_27_415 ();
 sg13g2_fill_2 FILLER_27_442 ();
 sg13g2_fill_2 FILLER_27_454 ();
 sg13g2_decap_8 FILLER_27_486 ();
 sg13g2_decap_8 FILLER_27_493 ();
 sg13g2_decap_4 FILLER_27_500 ();
 sg13g2_fill_1 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_541 ();
 sg13g2_decap_4 FILLER_27_548 ();
 sg13g2_fill_2 FILLER_27_552 ();
 sg13g2_fill_2 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_582 ();
 sg13g2_fill_2 FILLER_27_589 ();
 sg13g2_fill_1 FILLER_27_595 ();
 sg13g2_fill_2 FILLER_27_640 ();
 sg13g2_decap_8 FILLER_27_652 ();
 sg13g2_decap_4 FILLER_27_663 ();
 sg13g2_decap_8 FILLER_27_697 ();
 sg13g2_decap_8 FILLER_27_704 ();
 sg13g2_decap_8 FILLER_27_711 ();
 sg13g2_fill_1 FILLER_27_718 ();
 sg13g2_decap_4 FILLER_27_753 ();
 sg13g2_decap_8 FILLER_27_793 ();
 sg13g2_fill_2 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_fill_2 FILLER_27_814 ();
 sg13g2_fill_1 FILLER_27_816 ();
 sg13g2_decap_8 FILLER_27_867 ();
 sg13g2_fill_2 FILLER_27_874 ();
 sg13g2_fill_1 FILLER_27_907 ();
 sg13g2_fill_1 FILLER_27_922 ();
 sg13g2_decap_8 FILLER_27_949 ();
 sg13g2_decap_4 FILLER_27_982 ();
 sg13g2_fill_1 FILLER_27_986 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_decap_4 FILLER_27_1024 ();
 sg13g2_fill_2 FILLER_27_1028 ();
 sg13g2_decap_8 FILLER_27_1102 ();
 sg13g2_fill_1 FILLER_27_1109 ();
 sg13g2_decap_8 FILLER_27_1136 ();
 sg13g2_fill_1 FILLER_27_1143 ();
 sg13g2_fill_1 FILLER_27_1171 ();
 sg13g2_decap_8 FILLER_27_1202 ();
 sg13g2_decap_8 FILLER_27_1209 ();
 sg13g2_decap_8 FILLER_27_1216 ();
 sg13g2_decap_8 FILLER_27_1223 ();
 sg13g2_decap_4 FILLER_27_1230 ();
 sg13g2_fill_1 FILLER_27_1234 ();
 sg13g2_decap_8 FILLER_27_1259 ();
 sg13g2_decap_4 FILLER_27_1266 ();
 sg13g2_fill_1 FILLER_27_1270 ();
 sg13g2_decap_8 FILLER_27_1301 ();
 sg13g2_decap_8 FILLER_27_1308 ();
 sg13g2_decap_8 FILLER_27_1315 ();
 sg13g2_decap_8 FILLER_27_1322 ();
 sg13g2_fill_2 FILLER_27_1338 ();
 sg13g2_fill_1 FILLER_27_1340 ();
 sg13g2_fill_2 FILLER_27_1351 ();
 sg13g2_fill_1 FILLER_27_1353 ();
 sg13g2_decap_8 FILLER_27_1358 ();
 sg13g2_decap_4 FILLER_27_1365 ();
 sg13g2_fill_2 FILLER_27_1369 ();
 sg13g2_decap_4 FILLER_27_1421 ();
 sg13g2_decap_4 FILLER_27_1435 ();
 sg13g2_fill_2 FILLER_27_1460 ();
 sg13g2_fill_1 FILLER_27_1462 ();
 sg13g2_decap_8 FILLER_27_1467 ();
 sg13g2_fill_2 FILLER_27_1474 ();
 sg13g2_fill_1 FILLER_27_1476 ();
 sg13g2_decap_8 FILLER_27_1524 ();
 sg13g2_decap_8 FILLER_27_1531 ();
 sg13g2_fill_1 FILLER_27_1538 ();
 sg13g2_fill_2 FILLER_27_1575 ();
 sg13g2_fill_1 FILLER_27_1577 ();
 sg13g2_fill_2 FILLER_27_1588 ();
 sg13g2_decap_8 FILLER_27_1594 ();
 sg13g2_decap_8 FILLER_27_1601 ();
 sg13g2_decap_8 FILLER_27_1608 ();
 sg13g2_decap_8 FILLER_27_1615 ();
 sg13g2_decap_8 FILLER_27_1622 ();
 sg13g2_decap_8 FILLER_27_1629 ();
 sg13g2_fill_2 FILLER_27_1636 ();
 sg13g2_fill_1 FILLER_27_1638 ();
 sg13g2_fill_1 FILLER_27_1678 ();
 sg13g2_fill_1 FILLER_27_1683 ();
 sg13g2_fill_2 FILLER_27_1704 ();
 sg13g2_fill_1 FILLER_27_1706 ();
 sg13g2_fill_1 FILLER_27_1711 ();
 sg13g2_fill_1 FILLER_27_1716 ();
 sg13g2_fill_1 FILLER_27_1727 ();
 sg13g2_decap_4 FILLER_27_1738 ();
 sg13g2_fill_1 FILLER_27_1742 ();
 sg13g2_decap_8 FILLER_27_1747 ();
 sg13g2_decap_8 FILLER_27_1754 ();
 sg13g2_decap_8 FILLER_27_1761 ();
 sg13g2_decap_4 FILLER_27_1768 ();
 sg13g2_fill_2 FILLER_27_1772 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_59 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_75 ();
 sg13g2_decap_4 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_165 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_229 ();
 sg13g2_decap_8 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_250 ();
 sg13g2_fill_2 FILLER_28_257 ();
 sg13g2_decap_4 FILLER_28_263 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_decap_4 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_309 ();
 sg13g2_decap_8 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_decap_4 FILLER_28_348 ();
 sg13g2_fill_1 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_fill_2 FILLER_28_390 ();
 sg13g2_fill_1 FILLER_28_392 ();
 sg13g2_fill_2 FILLER_28_419 ();
 sg13g2_fill_1 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_488 ();
 sg13g2_decap_4 FILLER_28_511 ();
 sg13g2_fill_1 FILLER_28_515 ();
 sg13g2_decap_8 FILLER_28_546 ();
 sg13g2_decap_8 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_560 ();
 sg13g2_decap_8 FILLER_28_567 ();
 sg13g2_decap_8 FILLER_28_574 ();
 sg13g2_fill_1 FILLER_28_604 ();
 sg13g2_decap_8 FILLER_28_615 ();
 sg13g2_fill_2 FILLER_28_622 ();
 sg13g2_fill_2 FILLER_28_706 ();
 sg13g2_fill_1 FILLER_28_708 ();
 sg13g2_decap_8 FILLER_28_715 ();
 sg13g2_decap_4 FILLER_28_722 ();
 sg13g2_decap_8 FILLER_28_740 ();
 sg13g2_decap_8 FILLER_28_747 ();
 sg13g2_decap_8 FILLER_28_754 ();
 sg13g2_fill_1 FILLER_28_771 ();
 sg13g2_fill_1 FILLER_28_806 ();
 sg13g2_fill_2 FILLER_28_833 ();
 sg13g2_fill_2 FILLER_28_858 ();
 sg13g2_fill_1 FILLER_28_916 ();
 sg13g2_decap_4 FILLER_28_921 ();
 sg13g2_fill_2 FILLER_28_925 ();
 sg13g2_decap_8 FILLER_28_935 ();
 sg13g2_fill_1 FILLER_28_942 ();
 sg13g2_fill_2 FILLER_28_947 ();
 sg13g2_fill_2 FILLER_28_962 ();
 sg13g2_fill_1 FILLER_28_964 ();
 sg13g2_fill_2 FILLER_28_975 ();
 sg13g2_fill_1 FILLER_28_977 ();
 sg13g2_fill_2 FILLER_28_1004 ();
 sg13g2_fill_1 FILLER_28_1032 ();
 sg13g2_fill_2 FILLER_28_1038 ();
 sg13g2_fill_1 FILLER_28_1061 ();
 sg13g2_fill_2 FILLER_28_1066 ();
 sg13g2_fill_1 FILLER_28_1068 ();
 sg13g2_decap_8 FILLER_28_1077 ();
 sg13g2_fill_1 FILLER_28_1084 ();
 sg13g2_decap_4 FILLER_28_1089 ();
 sg13g2_fill_2 FILLER_28_1093 ();
 sg13g2_decap_4 FILLER_28_1101 ();
 sg13g2_fill_1 FILLER_28_1105 ();
 sg13g2_fill_1 FILLER_28_1161 ();
 sg13g2_decap_8 FILLER_28_1188 ();
 sg13g2_decap_8 FILLER_28_1195 ();
 sg13g2_decap_4 FILLER_28_1202 ();
 sg13g2_fill_2 FILLER_28_1206 ();
 sg13g2_fill_1 FILLER_28_1243 ();
 sg13g2_fill_1 FILLER_28_1254 ();
 sg13g2_decap_4 FILLER_28_1295 ();
 sg13g2_decap_8 FILLER_28_1303 ();
 sg13g2_fill_2 FILLER_28_1346 ();
 sg13g2_decap_8 FILLER_28_1374 ();
 sg13g2_fill_2 FILLER_28_1381 ();
 sg13g2_fill_1 FILLER_28_1383 ();
 sg13g2_fill_2 FILLER_28_1394 ();
 sg13g2_decap_4 FILLER_28_1422 ();
 sg13g2_decap_8 FILLER_28_1461 ();
 sg13g2_decap_8 FILLER_28_1468 ();
 sg13g2_fill_2 FILLER_28_1475 ();
 sg13g2_fill_1 FILLER_28_1477 ();
 sg13g2_fill_1 FILLER_28_1491 ();
 sg13g2_decap_8 FILLER_28_1532 ();
 sg13g2_decap_8 FILLER_28_1539 ();
 sg13g2_fill_2 FILLER_28_1546 ();
 sg13g2_decap_8 FILLER_28_1604 ();
 sg13g2_fill_2 FILLER_28_1611 ();
 sg13g2_decap_8 FILLER_28_1617 ();
 sg13g2_decap_8 FILLER_28_1624 ();
 sg13g2_decap_8 FILLER_28_1631 ();
 sg13g2_decap_8 FILLER_28_1638 ();
 sg13g2_decap_4 FILLER_28_1645 ();
 sg13g2_fill_2 FILLER_28_1649 ();
 sg13g2_decap_4 FILLER_28_1696 ();
 sg13g2_fill_2 FILLER_28_1700 ();
 sg13g2_decap_4 FILLER_28_1706 ();
 sg13g2_fill_2 FILLER_28_1710 ();
 sg13g2_decap_4 FILLER_28_1720 ();
 sg13g2_fill_2 FILLER_28_1724 ();
 sg13g2_decap_8 FILLER_28_1762 ();
 sg13g2_decap_4 FILLER_28_1769 ();
 sg13g2_fill_1 FILLER_28_1773 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_4 ();
 sg13g2_fill_2 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_37 ();
 sg13g2_fill_2 FILLER_29_54 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_83 ();
 sg13g2_decap_4 FILLER_29_131 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_decap_4 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_234 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_decap_4 FILLER_29_246 ();
 sg13g2_fill_2 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_260 ();
 sg13g2_decap_8 FILLER_29_267 ();
 sg13g2_decap_8 FILLER_29_274 ();
 sg13g2_decap_8 FILLER_29_281 ();
 sg13g2_fill_2 FILLER_29_288 ();
 sg13g2_fill_1 FILLER_29_290 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_decap_4 FILLER_29_330 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_2 FILLER_29_397 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_410 ();
 sg13g2_decap_4 FILLER_29_425 ();
 sg13g2_fill_2 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_29_448 ();
 sg13g2_fill_1 FILLER_29_460 ();
 sg13g2_decap_8 FILLER_29_496 ();
 sg13g2_decap_8 FILLER_29_503 ();
 sg13g2_fill_1 FILLER_29_524 ();
 sg13g2_decap_8 FILLER_29_565 ();
 sg13g2_decap_8 FILLER_29_572 ();
 sg13g2_decap_8 FILLER_29_579 ();
 sg13g2_fill_1 FILLER_29_616 ();
 sg13g2_decap_4 FILLER_29_653 ();
 sg13g2_fill_1 FILLER_29_657 ();
 sg13g2_fill_2 FILLER_29_693 ();
 sg13g2_fill_2 FILLER_29_734 ();
 sg13g2_decap_8 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_787 ();
 sg13g2_decap_4 FILLER_29_794 ();
 sg13g2_fill_2 FILLER_29_798 ();
 sg13g2_fill_2 FILLER_29_805 ();
 sg13g2_fill_1 FILLER_29_859 ();
 sg13g2_fill_1 FILLER_29_922 ();
 sg13g2_fill_2 FILLER_29_942 ();
 sg13g2_decap_8 FILLER_29_948 ();
 sg13g2_decap_4 FILLER_29_955 ();
 sg13g2_fill_1 FILLER_29_959 ();
 sg13g2_fill_2 FILLER_29_1018 ();
 sg13g2_decap_8 FILLER_29_1030 ();
 sg13g2_decap_8 FILLER_29_1037 ();
 sg13g2_fill_2 FILLER_29_1044 ();
 sg13g2_fill_1 FILLER_29_1046 ();
 sg13g2_fill_1 FILLER_29_1091 ();
 sg13g2_fill_1 FILLER_29_1179 ();
 sg13g2_decap_8 FILLER_29_1184 ();
 sg13g2_decap_8 FILLER_29_1191 ();
 sg13g2_decap_4 FILLER_29_1198 ();
 sg13g2_fill_2 FILLER_29_1202 ();
 sg13g2_decap_4 FILLER_29_1214 ();
 sg13g2_fill_1 FILLER_29_1218 ();
 sg13g2_decap_8 FILLER_29_1358 ();
 sg13g2_decap_4 FILLER_29_1365 ();
 sg13g2_fill_1 FILLER_29_1369 ();
 sg13g2_decap_8 FILLER_29_1375 ();
 sg13g2_decap_4 FILLER_29_1396 ();
 sg13g2_fill_1 FILLER_29_1400 ();
 sg13g2_decap_8 FILLER_29_1441 ();
 sg13g2_decap_8 FILLER_29_1448 ();
 sg13g2_fill_1 FILLER_29_1455 ();
 sg13g2_fill_1 FILLER_29_1482 ();
 sg13g2_decap_8 FILLER_29_1487 ();
 sg13g2_decap_4 FILLER_29_1494 ();
 sg13g2_fill_2 FILLER_29_1512 ();
 sg13g2_fill_2 FILLER_29_1518 ();
 sg13g2_fill_1 FILLER_29_1520 ();
 sg13g2_fill_2 FILLER_29_1551 ();
 sg13g2_fill_2 FILLER_29_1577 ();
 sg13g2_decap_8 FILLER_29_1631 ();
 sg13g2_decap_4 FILLER_29_1638 ();
 sg13g2_fill_2 FILLER_29_1642 ();
 sg13g2_fill_1 FILLER_29_1648 ();
 sg13g2_decap_4 FILLER_29_1680 ();
 sg13g2_fill_1 FILLER_29_1684 ();
 sg13g2_decap_4 FILLER_29_1721 ();
 sg13g2_fill_2 FILLER_29_1761 ();
 sg13g2_fill_1 FILLER_29_1763 ();
 sg13g2_decap_4 FILLER_29_1768 ();
 sg13g2_fill_2 FILLER_29_1772 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_17 ();
 sg13g2_decap_4 FILLER_30_24 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_62 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_225 ();
 sg13g2_decap_8 FILLER_30_253 ();
 sg13g2_decap_8 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_281 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_decap_4 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_2 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_314 ();
 sg13g2_decap_4 FILLER_30_351 ();
 sg13g2_fill_2 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_30_416 ();
 sg13g2_decap_8 FILLER_30_423 ();
 sg13g2_fill_1 FILLER_30_430 ();
 sg13g2_decap_8 FILLER_30_459 ();
 sg13g2_fill_2 FILLER_30_466 ();
 sg13g2_fill_1 FILLER_30_468 ();
 sg13g2_fill_2 FILLER_30_473 ();
 sg13g2_decap_8 FILLER_30_506 ();
 sg13g2_decap_4 FILLER_30_513 ();
 sg13g2_fill_2 FILLER_30_517 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_decap_4 FILLER_30_539 ();
 sg13g2_fill_2 FILLER_30_543 ();
 sg13g2_decap_8 FILLER_30_562 ();
 sg13g2_fill_1 FILLER_30_569 ();
 sg13g2_decap_4 FILLER_30_578 ();
 sg13g2_fill_1 FILLER_30_588 ();
 sg13g2_fill_1 FILLER_30_594 ();
 sg13g2_fill_1 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_638 ();
 sg13g2_decap_8 FILLER_30_655 ();
 sg13g2_fill_1 FILLER_30_662 ();
 sg13g2_fill_1 FILLER_30_667 ();
 sg13g2_fill_1 FILLER_30_723 ();
 sg13g2_fill_2 FILLER_30_727 ();
 sg13g2_fill_1 FILLER_30_743 ();
 sg13g2_fill_2 FILLER_30_748 ();
 sg13g2_decap_8 FILLER_30_786 ();
 sg13g2_decap_8 FILLER_30_793 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_fill_1 FILLER_30_807 ();
 sg13g2_fill_1 FILLER_30_834 ();
 sg13g2_fill_2 FILLER_30_851 ();
 sg13g2_fill_2 FILLER_30_879 ();
 sg13g2_fill_2 FILLER_30_884 ();
 sg13g2_fill_2 FILLER_30_915 ();
 sg13g2_fill_1 FILLER_30_943 ();
 sg13g2_fill_1 FILLER_30_949 ();
 sg13g2_fill_1 FILLER_30_955 ();
 sg13g2_fill_2 FILLER_30_1006 ();
 sg13g2_decap_8 FILLER_30_1038 ();
 sg13g2_decap_8 FILLER_30_1045 ();
 sg13g2_fill_1 FILLER_30_1052 ();
 sg13g2_fill_2 FILLER_30_1102 ();
 sg13g2_fill_2 FILLER_30_1117 ();
 sg13g2_fill_1 FILLER_30_1122 ();
 sg13g2_fill_1 FILLER_30_1132 ();
 sg13g2_fill_2 FILLER_30_1137 ();
 sg13g2_fill_1 FILLER_30_1142 ();
 sg13g2_fill_2 FILLER_30_1150 ();
 sg13g2_decap_8 FILLER_30_1175 ();
 sg13g2_decap_8 FILLER_30_1182 ();
 sg13g2_fill_2 FILLER_30_1189 ();
 sg13g2_fill_2 FILLER_30_1195 ();
 sg13g2_fill_1 FILLER_30_1197 ();
 sg13g2_fill_2 FILLER_30_1251 ();
 sg13g2_decap_8 FILLER_30_1304 ();
 sg13g2_fill_2 FILLER_30_1311 ();
 sg13g2_fill_1 FILLER_30_1313 ();
 sg13g2_fill_1 FILLER_30_1338 ();
 sg13g2_decap_8 FILLER_30_1365 ();
 sg13g2_decap_8 FILLER_30_1372 ();
 sg13g2_fill_2 FILLER_30_1379 ();
 sg13g2_fill_1 FILLER_30_1381 ();
 sg13g2_fill_1 FILLER_30_1426 ();
 sg13g2_fill_1 FILLER_30_1458 ();
 sg13g2_fill_1 FILLER_30_1469 ();
 sg13g2_decap_8 FILLER_30_1474 ();
 sg13g2_decap_8 FILLER_30_1481 ();
 sg13g2_fill_1 FILLER_30_1488 ();
 sg13g2_decap_8 FILLER_30_1499 ();
 sg13g2_fill_2 FILLER_30_1523 ();
 sg13g2_fill_1 FILLER_30_1545 ();
 sg13g2_fill_2 FILLER_30_1551 ();
 sg13g2_fill_2 FILLER_30_1563 ();
 sg13g2_fill_2 FILLER_30_1570 ();
 sg13g2_fill_2 FILLER_30_1594 ();
 sg13g2_fill_2 FILLER_30_1666 ();
 sg13g2_fill_1 FILLER_30_1668 ();
 sg13g2_decap_8 FILLER_30_1761 ();
 sg13g2_decap_4 FILLER_30_1768 ();
 sg13g2_fill_2 FILLER_30_1772 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_44 ();
 sg13g2_fill_1 FILLER_31_46 ();
 sg13g2_decap_4 FILLER_31_50 ();
 sg13g2_fill_1 FILLER_31_54 ();
 sg13g2_decap_8 FILLER_31_86 ();
 sg13g2_decap_8 FILLER_31_97 ();
 sg13g2_decap_8 FILLER_31_104 ();
 sg13g2_fill_1 FILLER_31_111 ();
 sg13g2_fill_1 FILLER_31_116 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_142 ();
 sg13g2_fill_1 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_fill_1 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_289 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_4 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_397 ();
 sg13g2_fill_1 FILLER_31_424 ();
 sg13g2_decap_4 FILLER_31_440 ();
 sg13g2_decap_8 FILLER_31_480 ();
 sg13g2_fill_1 FILLER_31_487 ();
 sg13g2_fill_1 FILLER_31_509 ();
 sg13g2_decap_8 FILLER_31_514 ();
 sg13g2_decap_8 FILLER_31_521 ();
 sg13g2_decap_8 FILLER_31_528 ();
 sg13g2_decap_8 FILLER_31_535 ();
 sg13g2_decap_8 FILLER_31_542 ();
 sg13g2_decap_8 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_556 ();
 sg13g2_decap_4 FILLER_31_563 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_fill_1 FILLER_31_595 ();
 sg13g2_fill_2 FILLER_31_604 ();
 sg13g2_fill_1 FILLER_31_606 ();
 sg13g2_fill_2 FILLER_31_611 ();
 sg13g2_fill_1 FILLER_31_613 ();
 sg13g2_decap_8 FILLER_31_650 ();
 sg13g2_fill_1 FILLER_31_657 ();
 sg13g2_decap_4 FILLER_31_668 ();
 sg13g2_fill_2 FILLER_31_672 ();
 sg13g2_fill_1 FILLER_31_682 ();
 sg13g2_decap_8 FILLER_31_779 ();
 sg13g2_decap_8 FILLER_31_786 ();
 sg13g2_decap_8 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_800 ();
 sg13g2_decap_8 FILLER_31_807 ();
 sg13g2_decap_4 FILLER_31_818 ();
 sg13g2_fill_1 FILLER_31_862 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_8 FILLER_31_952 ();
 sg13g2_fill_1 FILLER_31_959 ();
 sg13g2_fill_1 FILLER_31_964 ();
 sg13g2_fill_1 FILLER_31_975 ();
 sg13g2_fill_1 FILLER_31_997 ();
 sg13g2_fill_2 FILLER_31_1002 ();
 sg13g2_fill_2 FILLER_31_1044 ();
 sg13g2_decap_4 FILLER_31_1081 ();
 sg13g2_fill_2 FILLER_31_1085 ();
 sg13g2_fill_2 FILLER_31_1099 ();
 sg13g2_fill_2 FILLER_31_1137 ();
 sg13g2_decap_8 FILLER_31_1163 ();
 sg13g2_decap_8 FILLER_31_1170 ();
 sg13g2_decap_8 FILLER_31_1177 ();
 sg13g2_fill_2 FILLER_31_1184 ();
 sg13g2_fill_1 FILLER_31_1186 ();
 sg13g2_decap_4 FILLER_31_1257 ();
 sg13g2_fill_2 FILLER_31_1334 ();
 sg13g2_fill_1 FILLER_31_1336 ();
 sg13g2_decap_8 FILLER_31_1371 ();
 sg13g2_decap_4 FILLER_31_1378 ();
 sg13g2_fill_1 FILLER_31_1382 ();
 sg13g2_fill_2 FILLER_31_1411 ();
 sg13g2_fill_2 FILLER_31_1438 ();
 sg13g2_fill_2 FILLER_31_1466 ();
 sg13g2_fill_2 FILLER_31_1472 ();
 sg13g2_fill_1 FILLER_31_1474 ();
 sg13g2_fill_1 FILLER_31_1501 ();
 sg13g2_fill_2 FILLER_31_1528 ();
 sg13g2_fill_1 FILLER_31_1530 ();
 sg13g2_fill_1 FILLER_31_1562 ();
 sg13g2_decap_8 FILLER_31_1629 ();
 sg13g2_decap_8 FILLER_31_1636 ();
 sg13g2_fill_2 FILLER_31_1651 ();
 sg13g2_fill_1 FILLER_31_1653 ();
 sg13g2_fill_1 FILLER_31_1658 ();
 sg13g2_fill_2 FILLER_31_1739 ();
 sg13g2_decap_8 FILLER_31_1767 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_43 ();
 sg13g2_decap_8 FILLER_32_68 ();
 sg13g2_decap_8 FILLER_32_101 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_fill_2 FILLER_32_165 ();
 sg13g2_decap_4 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_289 ();
 sg13g2_decap_8 FILLER_32_300 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_2 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_341 ();
 sg13g2_decap_4 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_357 ();
 sg13g2_decap_4 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_421 ();
 sg13g2_fill_1 FILLER_32_448 ();
 sg13g2_fill_2 FILLER_32_479 ();
 sg13g2_fill_1 FILLER_32_481 ();
 sg13g2_decap_8 FILLER_32_529 ();
 sg13g2_fill_1 FILLER_32_536 ();
 sg13g2_decap_8 FILLER_32_592 ();
 sg13g2_decap_4 FILLER_32_672 ();
 sg13g2_fill_2 FILLER_32_676 ();
 sg13g2_fill_2 FILLER_32_749 ();
 sg13g2_fill_1 FILLER_32_751 ();
 sg13g2_fill_1 FILLER_32_761 ();
 sg13g2_decap_4 FILLER_32_766 ();
 sg13g2_fill_1 FILLER_32_770 ();
 sg13g2_fill_2 FILLER_32_776 ();
 sg13g2_fill_1 FILLER_32_778 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_4 FILLER_32_791 ();
 sg13g2_fill_2 FILLER_32_795 ();
 sg13g2_decap_8 FILLER_32_802 ();
 sg13g2_fill_1 FILLER_32_809 ();
 sg13g2_fill_2 FILLER_32_814 ();
 sg13g2_decap_4 FILLER_32_842 ();
 sg13g2_decap_4 FILLER_32_856 ();
 sg13g2_decap_8 FILLER_32_864 ();
 sg13g2_decap_8 FILLER_32_930 ();
 sg13g2_decap_8 FILLER_32_937 ();
 sg13g2_decap_8 FILLER_32_944 ();
 sg13g2_fill_2 FILLER_32_951 ();
 sg13g2_fill_1 FILLER_32_953 ();
 sg13g2_fill_1 FILLER_32_994 ();
 sg13g2_fill_2 FILLER_32_1008 ();
 sg13g2_fill_2 FILLER_32_1031 ();
 sg13g2_decap_8 FILLER_32_1039 ();
 sg13g2_fill_2 FILLER_32_1050 ();
 sg13g2_decap_8 FILLER_32_1078 ();
 sg13g2_decap_8 FILLER_32_1085 ();
 sg13g2_fill_2 FILLER_32_1147 ();
 sg13g2_fill_2 FILLER_32_1180 ();
 sg13g2_fill_1 FILLER_32_1182 ();
 sg13g2_fill_2 FILLER_32_1192 ();
 sg13g2_fill_1 FILLER_32_1275 ();
 sg13g2_fill_2 FILLER_32_1288 ();
 sg13g2_fill_1 FILLER_32_1300 ();
 sg13g2_fill_2 FILLER_32_1327 ();
 sg13g2_fill_1 FILLER_32_1329 ();
 sg13g2_decap_4 FILLER_32_1350 ();
 sg13g2_fill_1 FILLER_32_1354 ();
 sg13g2_fill_2 FILLER_32_1369 ();
 sg13g2_fill_1 FILLER_32_1371 ();
 sg13g2_decap_4 FILLER_32_1414 ();
 sg13g2_fill_1 FILLER_32_1418 ();
 sg13g2_fill_2 FILLER_32_1429 ();
 sg13g2_fill_1 FILLER_32_1431 ();
 sg13g2_decap_8 FILLER_32_1436 ();
 sg13g2_decap_8 FILLER_32_1443 ();
 sg13g2_decap_8 FILLER_32_1460 ();
 sg13g2_fill_2 FILLER_32_1467 ();
 sg13g2_fill_1 FILLER_32_1469 ();
 sg13g2_decap_4 FILLER_32_1478 ();
 sg13g2_fill_1 FILLER_32_1482 ();
 sg13g2_fill_2 FILLER_32_1495 ();
 sg13g2_fill_1 FILLER_32_1497 ();
 sg13g2_fill_1 FILLER_32_1508 ();
 sg13g2_fill_1 FILLER_32_1513 ();
 sg13g2_fill_2 FILLER_32_1550 ();
 sg13g2_fill_2 FILLER_32_1560 ();
 sg13g2_decap_4 FILLER_32_1598 ();
 sg13g2_fill_1 FILLER_32_1602 ();
 sg13g2_fill_2 FILLER_32_1639 ();
 sg13g2_fill_1 FILLER_32_1641 ();
 sg13g2_fill_1 FILLER_32_1652 ();
 sg13g2_fill_2 FILLER_32_1673 ();
 sg13g2_fill_1 FILLER_32_1675 ();
 sg13g2_decap_4 FILLER_32_1686 ();
 sg13g2_fill_1 FILLER_32_1690 ();
 sg13g2_fill_1 FILLER_32_1695 ();
 sg13g2_decap_8 FILLER_32_1705 ();
 sg13g2_decap_8 FILLER_32_1712 ();
 sg13g2_decap_8 FILLER_32_1719 ();
 sg13g2_fill_2 FILLER_32_1726 ();
 sg13g2_decap_4 FILLER_32_1768 ();
 sg13g2_fill_2 FILLER_32_1772 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_23 ();
 sg13g2_fill_2 FILLER_33_50 ();
 sg13g2_fill_2 FILLER_33_62 ();
 sg13g2_fill_2 FILLER_33_90 ();
 sg13g2_fill_1 FILLER_33_92 ();
 sg13g2_decap_4 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_133 ();
 sg13g2_decap_4 FILLER_33_183 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_284 ();
 sg13g2_fill_1 FILLER_33_286 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_fill_1 FILLER_33_411 ();
 sg13g2_fill_1 FILLER_33_448 ();
 sg13g2_fill_1 FILLER_33_459 ();
 sg13g2_fill_1 FILLER_33_464 ();
 sg13g2_fill_1 FILLER_33_507 ();
 sg13g2_fill_1 FILLER_33_534 ();
 sg13g2_fill_2 FILLER_33_571 ();
 sg13g2_fill_1 FILLER_33_579 ();
 sg13g2_fill_2 FILLER_33_606 ();
 sg13g2_fill_1 FILLER_33_640 ();
 sg13g2_fill_2 FILLER_33_728 ();
 sg13g2_decap_4 FILLER_33_766 ();
 sg13g2_fill_1 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_4 FILLER_33_811 ();
 sg13g2_fill_1 FILLER_33_815 ();
 sg13g2_fill_1 FILLER_33_852 ();
 sg13g2_decap_8 FILLER_33_899 ();
 sg13g2_fill_2 FILLER_33_932 ();
 sg13g2_fill_1 FILLER_33_934 ();
 sg13g2_decap_8 FILLER_33_943 ();
 sg13g2_decap_8 FILLER_33_950 ();
 sg13g2_decap_4 FILLER_33_957 ();
 sg13g2_decap_8 FILLER_33_997 ();
 sg13g2_decap_8 FILLER_33_1004 ();
 sg13g2_decap_4 FILLER_33_1011 ();
 sg13g2_fill_1 FILLER_33_1015 ();
 sg13g2_decap_8 FILLER_33_1084 ();
 sg13g2_fill_2 FILLER_33_1091 ();
 sg13g2_fill_2 FILLER_33_1152 ();
 sg13g2_fill_1 FILLER_33_1212 ();
 sg13g2_fill_1 FILLER_33_1223 ();
 sg13g2_fill_1 FILLER_33_1261 ();
 sg13g2_fill_1 FILLER_33_1268 ();
 sg13g2_fill_2 FILLER_33_1282 ();
 sg13g2_fill_2 FILLER_33_1288 ();
 sg13g2_decap_8 FILLER_33_1295 ();
 sg13g2_fill_1 FILLER_33_1302 ();
 sg13g2_decap_8 FILLER_33_1311 ();
 sg13g2_fill_2 FILLER_33_1318 ();
 sg13g2_decap_4 FILLER_33_1341 ();
 sg13g2_fill_1 FILLER_33_1345 ();
 sg13g2_decap_8 FILLER_33_1372 ();
 sg13g2_fill_2 FILLER_33_1379 ();
 sg13g2_fill_1 FILLER_33_1381 ();
 sg13g2_decap_8 FILLER_33_1395 ();
 sg13g2_fill_2 FILLER_33_1402 ();
 sg13g2_fill_1 FILLER_33_1404 ();
 sg13g2_decap_8 FILLER_33_1431 ();
 sg13g2_decap_4 FILLER_33_1438 ();
 sg13g2_fill_1 FILLER_33_1446 ();
 sg13g2_decap_8 FILLER_33_1473 ();
 sg13g2_fill_1 FILLER_33_1480 ();
 sg13g2_decap_8 FILLER_33_1495 ();
 sg13g2_fill_2 FILLER_33_1538 ();
 sg13g2_fill_2 FILLER_33_1575 ();
 sg13g2_fill_1 FILLER_33_1603 ();
 sg13g2_decap_4 FILLER_33_1640 ();
 sg13g2_fill_1 FILLER_33_1668 ();
 sg13g2_decap_8 FILLER_33_1673 ();
 sg13g2_decap_8 FILLER_33_1680 ();
 sg13g2_decap_8 FILLER_33_1708 ();
 sg13g2_fill_2 FILLER_33_1715 ();
 sg13g2_fill_1 FILLER_33_1717 ();
 sg13g2_decap_8 FILLER_33_1728 ();
 sg13g2_fill_2 FILLER_33_1761 ();
 sg13g2_fill_1 FILLER_33_1763 ();
 sg13g2_decap_4 FILLER_33_1768 ();
 sg13g2_fill_2 FILLER_33_1772 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_fill_1 FILLER_34_45 ();
 sg13g2_decap_8 FILLER_34_90 ();
 sg13g2_decap_4 FILLER_34_97 ();
 sg13g2_decap_4 FILLER_34_115 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_decap_4 FILLER_34_156 ();
 sg13g2_fill_2 FILLER_34_160 ();
 sg13g2_decap_4 FILLER_34_171 ();
 sg13g2_fill_2 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_191 ();
 sg13g2_fill_2 FILLER_34_198 ();
 sg13g2_decap_4 FILLER_34_212 ();
 sg13g2_fill_2 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_260 ();
 sg13g2_decap_8 FILLER_34_288 ();
 sg13g2_decap_8 FILLER_34_295 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_330 ();
 sg13g2_decap_8 FILLER_34_337 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_2 FILLER_34_457 ();
 sg13g2_fill_1 FILLER_34_514 ();
 sg13g2_decap_4 FILLER_34_532 ();
 sg13g2_decap_4 FILLER_34_546 ();
 sg13g2_decap_8 FILLER_34_554 ();
 sg13g2_decap_8 FILLER_34_561 ();
 sg13g2_decap_4 FILLER_34_568 ();
 sg13g2_decap_4 FILLER_34_577 ();
 sg13g2_fill_1 FILLER_34_602 ();
 sg13g2_fill_1 FILLER_34_613 ();
 sg13g2_fill_2 FILLER_34_617 ();
 sg13g2_fill_1 FILLER_34_626 ();
 sg13g2_fill_2 FILLER_34_653 ();
 sg13g2_fill_1 FILLER_34_655 ();
 sg13g2_fill_1 FILLER_34_671 ();
 sg13g2_fill_1 FILLER_34_678 ();
 sg13g2_decap_8 FILLER_34_689 ();
 sg13g2_fill_2 FILLER_34_696 ();
 sg13g2_fill_1 FILLER_34_710 ();
 sg13g2_fill_1 FILLER_34_733 ();
 sg13g2_decap_8 FILLER_34_765 ();
 sg13g2_decap_4 FILLER_34_785 ();
 sg13g2_fill_1 FILLER_34_789 ();
 sg13g2_decap_4 FILLER_34_799 ();
 sg13g2_fill_1 FILLER_34_803 ();
 sg13g2_decap_4 FILLER_34_827 ();
 sg13g2_decap_8 FILLER_34_835 ();
 sg13g2_fill_1 FILLER_34_873 ();
 sg13g2_decap_4 FILLER_34_930 ();
 sg13g2_fill_1 FILLER_34_934 ();
 sg13g2_decap_4 FILLER_34_948 ();
 sg13g2_fill_1 FILLER_34_999 ();
 sg13g2_fill_1 FILLER_34_1026 ();
 sg13g2_fill_1 FILLER_34_1032 ();
 sg13g2_decap_4 FILLER_34_1043 ();
 sg13g2_fill_1 FILLER_34_1047 ();
 sg13g2_decap_8 FILLER_34_1078 ();
 sg13g2_fill_2 FILLER_34_1085 ();
 sg13g2_decap_4 FILLER_34_1093 ();
 sg13g2_decap_8 FILLER_34_1118 ();
 sg13g2_fill_1 FILLER_34_1125 ();
 sg13g2_decap_4 FILLER_34_1129 ();
 sg13g2_fill_1 FILLER_34_1133 ();
 sg13g2_fill_1 FILLER_34_1144 ();
 sg13g2_fill_2 FILLER_34_1156 ();
 sg13g2_fill_2 FILLER_34_1189 ();
 sg13g2_fill_1 FILLER_34_1195 ();
 sg13g2_decap_8 FILLER_34_1254 ();
 sg13g2_fill_1 FILLER_34_1261 ();
 sg13g2_decap_8 FILLER_34_1265 ();
 sg13g2_decap_4 FILLER_34_1272 ();
 sg13g2_fill_1 FILLER_34_1284 ();
 sg13g2_decap_4 FILLER_34_1288 ();
 sg13g2_fill_1 FILLER_34_1292 ();
 sg13g2_decap_8 FILLER_34_1391 ();
 sg13g2_decap_8 FILLER_34_1398 ();
 sg13g2_fill_2 FILLER_34_1405 ();
 sg13g2_fill_2 FILLER_34_1463 ();
 sg13g2_fill_1 FILLER_34_1465 ();
 sg13g2_decap_8 FILLER_34_1502 ();
 sg13g2_decap_8 FILLER_34_1509 ();
 sg13g2_decap_4 FILLER_34_1516 ();
 sg13g2_fill_1 FILLER_34_1520 ();
 sg13g2_fill_1 FILLER_34_1557 ();
 sg13g2_fill_2 FILLER_34_1626 ();
 sg13g2_fill_1 FILLER_34_1628 ();
 sg13g2_decap_8 FILLER_34_1633 ();
 sg13g2_decap_4 FILLER_34_1640 ();
 sg13g2_decap_4 FILLER_34_1680 ();
 sg13g2_fill_1 FILLER_34_1684 ();
 sg13g2_fill_2 FILLER_34_1689 ();
 sg13g2_fill_2 FILLER_34_1717 ();
 sg13g2_fill_1 FILLER_34_1719 ();
 sg13g2_fill_2 FILLER_34_1730 ();
 sg13g2_fill_1 FILLER_34_1732 ();
 sg13g2_decap_8 FILLER_34_1763 ();
 sg13g2_decap_4 FILLER_34_1770 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_14 ();
 sg13g2_decap_4 FILLER_35_22 ();
 sg13g2_fill_2 FILLER_35_26 ();
 sg13g2_fill_1 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_45 ();
 sg13g2_decap_8 FILLER_35_57 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_decap_8 FILLER_35_69 ();
 sg13g2_decap_8 FILLER_35_76 ();
 sg13g2_decap_8 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_90 ();
 sg13g2_fill_1 FILLER_35_92 ();
 sg13g2_decap_8 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_113 ();
 sg13g2_decap_8 FILLER_35_151 ();
 sg13g2_decap_8 FILLER_35_158 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_decap_4 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_224 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_fill_2 FILLER_35_359 ();
 sg13g2_fill_1 FILLER_35_361 ();
 sg13g2_decap_4 FILLER_35_380 ();
 sg13g2_fill_2 FILLER_35_384 ();
 sg13g2_fill_2 FILLER_35_452 ();
 sg13g2_fill_2 FILLER_35_460 ();
 sg13g2_decap_8 FILLER_35_499 ();
 sg13g2_decap_8 FILLER_35_506 ();
 sg13g2_decap_8 FILLER_35_513 ();
 sg13g2_decap_4 FILLER_35_520 ();
 sg13g2_fill_1 FILLER_35_524 ();
 sg13g2_fill_2 FILLER_35_530 ();
 sg13g2_fill_1 FILLER_35_532 ();
 sg13g2_fill_1 FILLER_35_573 ();
 sg13g2_fill_2 FILLER_35_584 ();
 sg13g2_decap_4 FILLER_35_591 ();
 sg13g2_fill_1 FILLER_35_609 ();
 sg13g2_fill_2 FILLER_35_645 ();
 sg13g2_fill_1 FILLER_35_647 ();
 sg13g2_fill_1 FILLER_35_674 ();
 sg13g2_fill_2 FILLER_35_699 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_fill_2 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_771 ();
 sg13g2_decap_8 FILLER_35_778 ();
 sg13g2_decap_4 FILLER_35_785 ();
 sg13g2_fill_1 FILLER_35_789 ();
 sg13g2_decap_4 FILLER_35_794 ();
 sg13g2_fill_2 FILLER_35_798 ();
 sg13g2_fill_2 FILLER_35_806 ();
 sg13g2_decap_4 FILLER_35_852 ();
 sg13g2_decap_4 FILLER_35_860 ();
 sg13g2_fill_2 FILLER_35_864 ();
 sg13g2_decap_4 FILLER_35_922 ();
 sg13g2_fill_2 FILLER_35_926 ();
 sg13g2_fill_2 FILLER_35_933 ();
 sg13g2_fill_1 FILLER_35_935 ();
 sg13g2_decap_8 FILLER_35_941 ();
 sg13g2_fill_1 FILLER_35_948 ();
 sg13g2_fill_1 FILLER_35_959 ();
 sg13g2_fill_2 FILLER_35_964 ();
 sg13g2_fill_1 FILLER_35_966 ();
 sg13g2_decap_4 FILLER_35_979 ();
 sg13g2_fill_1 FILLER_35_1009 ();
 sg13g2_decap_4 FILLER_35_1028 ();
 sg13g2_fill_1 FILLER_35_1032 ();
 sg13g2_decap_4 FILLER_35_1039 ();
 sg13g2_fill_2 FILLER_35_1043 ();
 sg13g2_fill_1 FILLER_35_1050 ();
 sg13g2_fill_1 FILLER_35_1061 ();
 sg13g2_decap_8 FILLER_35_1070 ();
 sg13g2_decap_4 FILLER_35_1077 ();
 sg13g2_fill_1 FILLER_35_1081 ();
 sg13g2_decap_4 FILLER_35_1143 ();
 sg13g2_fill_1 FILLER_35_1147 ();
 sg13g2_decap_4 FILLER_35_1157 ();
 sg13g2_fill_1 FILLER_35_1161 ();
 sg13g2_fill_2 FILLER_35_1196 ();
 sg13g2_decap_8 FILLER_35_1253 ();
 sg13g2_decap_8 FILLER_35_1260 ();
 sg13g2_decap_4 FILLER_35_1267 ();
 sg13g2_fill_2 FILLER_35_1271 ();
 sg13g2_decap_4 FILLER_35_1277 ();
 sg13g2_fill_1 FILLER_35_1281 ();
 sg13g2_decap_4 FILLER_35_1328 ();
 sg13g2_fill_1 FILLER_35_1332 ();
 sg13g2_fill_2 FILLER_35_1348 ();
 sg13g2_fill_1 FILLER_35_1354 ();
 sg13g2_decap_8 FILLER_35_1395 ();
 sg13g2_decap_8 FILLER_35_1402 ();
 sg13g2_decap_8 FILLER_35_1409 ();
 sg13g2_fill_2 FILLER_35_1416 ();
 sg13g2_decap_4 FILLER_35_1422 ();
 sg13g2_decap_8 FILLER_35_1450 ();
 sg13g2_decap_4 FILLER_35_1457 ();
 sg13g2_fill_1 FILLER_35_1461 ();
 sg13g2_decap_8 FILLER_35_1488 ();
 sg13g2_decap_8 FILLER_35_1521 ();
 sg13g2_decap_4 FILLER_35_1528 ();
 sg13g2_fill_1 FILLER_35_1532 ();
 sg13g2_fill_2 FILLER_35_1537 ();
 sg13g2_fill_1 FILLER_35_1542 ();
 sg13g2_fill_1 FILLER_35_1588 ();
 sg13g2_decap_8 FILLER_35_1619 ();
 sg13g2_decap_8 FILLER_35_1626 ();
 sg13g2_decap_8 FILLER_35_1633 ();
 sg13g2_fill_2 FILLER_35_1680 ();
 sg13g2_fill_1 FILLER_35_1682 ();
 sg13g2_decap_4 FILLER_35_1769 ();
 sg13g2_fill_1 FILLER_35_1773 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_40 ();
 sg13g2_decap_8 FILLER_36_55 ();
 sg13g2_decap_8 FILLER_36_72 ();
 sg13g2_fill_2 FILLER_36_79 ();
 sg13g2_decap_8 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_decap_4 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_decap_4 FILLER_36_130 ();
 sg13g2_fill_2 FILLER_36_134 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_4 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_165 ();
 sg13g2_fill_2 FILLER_36_191 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_204 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_decap_4 FILLER_36_321 ();
 sg13g2_fill_2 FILLER_36_325 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_fill_2 FILLER_36_387 ();
 sg13g2_fill_2 FILLER_36_413 ();
 sg13g2_fill_1 FILLER_36_415 ();
 sg13g2_fill_2 FILLER_36_452 ();
 sg13g2_fill_2 FILLER_36_460 ();
 sg13g2_decap_8 FILLER_36_508 ();
 sg13g2_decap_8 FILLER_36_523 ();
 sg13g2_fill_1 FILLER_36_530 ();
 sg13g2_fill_2 FILLER_36_567 ();
 sg13g2_decap_8 FILLER_36_636 ();
 sg13g2_decap_4 FILLER_36_653 ();
 sg13g2_fill_2 FILLER_36_657 ();
 sg13g2_fill_1 FILLER_36_669 ();
 sg13g2_fill_2 FILLER_36_688 ();
 sg13g2_fill_1 FILLER_36_690 ();
 sg13g2_fill_1 FILLER_36_694 ();
 sg13g2_fill_1 FILLER_36_705 ();
 sg13g2_decap_8 FILLER_36_750 ();
 sg13g2_decap_8 FILLER_36_757 ();
 sg13g2_decap_8 FILLER_36_764 ();
 sg13g2_fill_1 FILLER_36_797 ();
 sg13g2_fill_2 FILLER_36_844 ();
 sg13g2_fill_1 FILLER_36_846 ();
 sg13g2_decap_4 FILLER_36_855 ();
 sg13g2_fill_1 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_882 ();
 sg13g2_fill_1 FILLER_36_889 ();
 sg13g2_fill_1 FILLER_36_894 ();
 sg13g2_decap_4 FILLER_36_905 ();
 sg13g2_fill_2 FILLER_36_909 ();
 sg13g2_decap_8 FILLER_36_915 ();
 sg13g2_decap_8 FILLER_36_922 ();
 sg13g2_decap_8 FILLER_36_929 ();
 sg13g2_decap_8 FILLER_36_946 ();
 sg13g2_decap_8 FILLER_36_953 ();
 sg13g2_decap_8 FILLER_36_960 ();
 sg13g2_decap_8 FILLER_36_967 ();
 sg13g2_fill_2 FILLER_36_974 ();
 sg13g2_fill_1 FILLER_36_976 ();
 sg13g2_fill_1 FILLER_36_995 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_4 FILLER_36_1015 ();
 sg13g2_fill_2 FILLER_36_1019 ();
 sg13g2_fill_2 FILLER_36_1026 ();
 sg13g2_decap_8 FILLER_36_1052 ();
 sg13g2_fill_2 FILLER_36_1059 ();
 sg13g2_fill_1 FILLER_36_1061 ();
 sg13g2_fill_1 FILLER_36_1074 ();
 sg13g2_decap_4 FILLER_36_1107 ();
 sg13g2_fill_1 FILLER_36_1115 ();
 sg13g2_decap_4 FILLER_36_1121 ();
 sg13g2_fill_2 FILLER_36_1125 ();
 sg13g2_fill_2 FILLER_36_1136 ();
 sg13g2_fill_1 FILLER_36_1138 ();
 sg13g2_decap_4 FILLER_36_1149 ();
 sg13g2_decap_4 FILLER_36_1157 ();
 sg13g2_fill_1 FILLER_36_1171 ();
 sg13g2_fill_2 FILLER_36_1262 ();
 sg13g2_fill_2 FILLER_36_1290 ();
 sg13g2_decap_4 FILLER_36_1296 ();
 sg13g2_fill_2 FILLER_36_1318 ();
 sg13g2_fill_1 FILLER_36_1320 ();
 sg13g2_fill_1 FILLER_36_1354 ();
 sg13g2_decap_8 FILLER_36_1359 ();
 sg13g2_decap_4 FILLER_36_1366 ();
 sg13g2_fill_1 FILLER_36_1378 ();
 sg13g2_decap_8 FILLER_36_1400 ();
 sg13g2_decap_8 FILLER_36_1407 ();
 sg13g2_decap_8 FILLER_36_1414 ();
 sg13g2_fill_1 FILLER_36_1421 ();
 sg13g2_decap_8 FILLER_36_1430 ();
 sg13g2_decap_8 FILLER_36_1437 ();
 sg13g2_decap_8 FILLER_36_1444 ();
 sg13g2_decap_8 FILLER_36_1451 ();
 sg13g2_decap_8 FILLER_36_1458 ();
 sg13g2_decap_4 FILLER_36_1465 ();
 sg13g2_fill_1 FILLER_36_1469 ();
 sg13g2_decap_8 FILLER_36_1483 ();
 sg13g2_fill_2 FILLER_36_1500 ();
 sg13g2_fill_1 FILLER_36_1502 ();
 sg13g2_fill_2 FILLER_36_1507 ();
 sg13g2_fill_1 FILLER_36_1509 ();
 sg13g2_fill_2 FILLER_36_1520 ();
 sg13g2_fill_1 FILLER_36_1522 ();
 sg13g2_fill_2 FILLER_36_1533 ();
 sg13g2_fill_1 FILLER_36_1535 ();
 sg13g2_fill_2 FILLER_36_1545 ();
 sg13g2_decap_4 FILLER_36_1607 ();
 sg13g2_fill_2 FILLER_36_1637 ();
 sg13g2_fill_1 FILLER_36_1639 ();
 sg13g2_fill_2 FILLER_36_1648 ();
 sg13g2_fill_1 FILLER_36_1650 ();
 sg13g2_decap_4 FILLER_36_1692 ();
 sg13g2_fill_2 FILLER_36_1696 ();
 sg13g2_fill_2 FILLER_36_1723 ();
 sg13g2_fill_2 FILLER_36_1735 ();
 sg13g2_decap_8 FILLER_36_1763 ();
 sg13g2_decap_4 FILLER_36_1770 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_13 ();
 sg13g2_fill_2 FILLER_37_40 ();
 sg13g2_fill_2 FILLER_37_108 ();
 sg13g2_fill_1 FILLER_37_136 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_decap_4 FILLER_37_184 ();
 sg13g2_decap_8 FILLER_37_219 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_fill_2 FILLER_37_290 ();
 sg13g2_decap_4 FILLER_37_302 ();
 sg13g2_decap_4 FILLER_37_336 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_decap_4 FILLER_37_345 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_decap_4 FILLER_37_397 ();
 sg13g2_fill_1 FILLER_37_401 ();
 sg13g2_decap_8 FILLER_37_414 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_decap_4 FILLER_37_428 ();
 sg13g2_fill_2 FILLER_37_481 ();
 sg13g2_fill_1 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_fill_2 FILLER_37_546 ();
 sg13g2_fill_1 FILLER_37_548 ();
 sg13g2_decap_8 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_fill_2 FILLER_37_567 ();
 sg13g2_decap_4 FILLER_37_572 ();
 sg13g2_fill_2 FILLER_37_576 ();
 sg13g2_decap_4 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_635 ();
 sg13g2_fill_2 FILLER_37_678 ();
 sg13g2_decap_8 FILLER_37_706 ();
 sg13g2_decap_8 FILLER_37_713 ();
 sg13g2_decap_4 FILLER_37_759 ();
 sg13g2_decap_4 FILLER_37_767 ();
 sg13g2_fill_2 FILLER_37_771 ();
 sg13g2_fill_1 FILLER_37_802 ();
 sg13g2_fill_2 FILLER_37_840 ();
 sg13g2_fill_2 FILLER_37_847 ();
 sg13g2_fill_1 FILLER_37_849 ();
 sg13g2_fill_2 FILLER_37_855 ();
 sg13g2_fill_2 FILLER_37_867 ();
 sg13g2_fill_1 FILLER_37_885 ();
 sg13g2_fill_1 FILLER_37_893 ();
 sg13g2_decap_8 FILLER_37_907 ();
 sg13g2_decap_8 FILLER_37_914 ();
 sg13g2_decap_8 FILLER_37_967 ();
 sg13g2_fill_2 FILLER_37_974 ();
 sg13g2_fill_1 FILLER_37_976 ();
 sg13g2_decap_8 FILLER_37_981 ();
 sg13g2_fill_2 FILLER_37_988 ();
 sg13g2_decap_8 FILLER_37_1003 ();
 sg13g2_decap_8 FILLER_37_1010 ();
 sg13g2_fill_1 FILLER_37_1017 ();
 sg13g2_fill_2 FILLER_37_1022 ();
 sg13g2_fill_2 FILLER_37_1028 ();
 sg13g2_decap_4 FILLER_37_1064 ();
 sg13g2_fill_2 FILLER_37_1072 ();
 sg13g2_fill_1 FILLER_37_1092 ();
 sg13g2_fill_1 FILLER_37_1106 ();
 sg13g2_fill_1 FILLER_37_1115 ();
 sg13g2_decap_8 FILLER_37_1137 ();
 sg13g2_fill_2 FILLER_37_1144 ();
 sg13g2_fill_2 FILLER_37_1176 ();
 sg13g2_fill_1 FILLER_37_1178 ();
 sg13g2_fill_1 FILLER_37_1217 ();
 sg13g2_fill_1 FILLER_37_1226 ();
 sg13g2_fill_1 FILLER_37_1257 ();
 sg13g2_fill_1 FILLER_37_1263 ();
 sg13g2_decap_4 FILLER_37_1305 ();
 sg13g2_fill_1 FILLER_37_1309 ();
 sg13g2_fill_2 FILLER_37_1336 ();
 sg13g2_fill_1 FILLER_37_1344 ();
 sg13g2_decap_4 FILLER_37_1371 ();
 sg13g2_fill_2 FILLER_37_1405 ();
 sg13g2_fill_2 FILLER_37_1433 ();
 sg13g2_decap_4 FILLER_37_1445 ();
 sg13g2_fill_1 FILLER_37_1449 ();
 sg13g2_decap_8 FILLER_37_1454 ();
 sg13g2_decap_4 FILLER_37_1461 ();
 sg13g2_fill_1 FILLER_37_1465 ();
 sg13g2_fill_2 FILLER_37_1476 ();
 sg13g2_fill_1 FILLER_37_1503 ();
 sg13g2_fill_2 FILLER_37_1530 ();
 sg13g2_fill_2 FILLER_37_1559 ();
 sg13g2_decap_8 FILLER_37_1571 ();
 sg13g2_fill_2 FILLER_37_1578 ();
 sg13g2_fill_1 FILLER_37_1580 ();
 sg13g2_decap_8 FILLER_37_1601 ();
 sg13g2_fill_2 FILLER_37_1608 ();
 sg13g2_fill_1 FILLER_37_1610 ();
 sg13g2_decap_8 FILLER_37_1641 ();
 sg13g2_decap_4 FILLER_37_1648 ();
 sg13g2_fill_1 FILLER_37_1652 ();
 sg13g2_fill_2 FILLER_37_1724 ();
 sg13g2_fill_1 FILLER_37_1731 ();
 sg13g2_decap_8 FILLER_37_1736 ();
 sg13g2_fill_2 FILLER_37_1743 ();
 sg13g2_decap_8 FILLER_37_1749 ();
 sg13g2_decap_8 FILLER_37_1756 ();
 sg13g2_decap_8 FILLER_37_1763 ();
 sg13g2_decap_4 FILLER_37_1770 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_4 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_80 ();
 sg13g2_fill_1 FILLER_38_92 ();
 sg13g2_fill_2 FILLER_38_103 ();
 sg13g2_fill_2 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_fill_1 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_267 ();
 sg13g2_decap_4 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_fill_1 FILLER_38_396 ();
 sg13g2_fill_1 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_409 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_4 FILLER_38_434 ();
 sg13g2_fill_2 FILLER_38_448 ();
 sg13g2_decap_4 FILLER_38_476 ();
 sg13g2_fill_2 FILLER_38_499 ();
 sg13g2_fill_1 FILLER_38_501 ();
 sg13g2_decap_8 FILLER_38_507 ();
 sg13g2_decap_8 FILLER_38_514 ();
 sg13g2_fill_1 FILLER_38_521 ();
 sg13g2_decap_8 FILLER_38_548 ();
 sg13g2_decap_8 FILLER_38_555 ();
 sg13g2_fill_1 FILLER_38_562 ();
 sg13g2_fill_1 FILLER_38_584 ();
 sg13g2_fill_1 FILLER_38_589 ();
 sg13g2_fill_1 FILLER_38_596 ();
 sg13g2_fill_1 FILLER_38_607 ();
 sg13g2_fill_1 FILLER_38_673 ();
 sg13g2_decap_4 FILLER_38_710 ();
 sg13g2_fill_2 FILLER_38_714 ();
 sg13g2_fill_1 FILLER_38_720 ();
 sg13g2_decap_4 FILLER_38_751 ();
 sg13g2_fill_2 FILLER_38_755 ();
 sg13g2_fill_2 FILLER_38_783 ();
 sg13g2_fill_1 FILLER_38_806 ();
 sg13g2_fill_2 FILLER_38_817 ();
 sg13g2_fill_2 FILLER_38_829 ();
 sg13g2_fill_1 FILLER_38_831 ();
 sg13g2_decap_8 FILLER_38_902 ();
 sg13g2_decap_8 FILLER_38_909 ();
 sg13g2_decap_8 FILLER_38_916 ();
 sg13g2_fill_1 FILLER_38_923 ();
 sg13g2_decap_8 FILLER_38_954 ();
 sg13g2_decap_4 FILLER_38_961 ();
 sg13g2_fill_1 FILLER_38_975 ();
 sg13g2_fill_1 FILLER_38_1038 ();
 sg13g2_fill_2 FILLER_38_1088 ();
 sg13g2_fill_2 FILLER_38_1123 ();
 sg13g2_fill_1 FILLER_38_1125 ();
 sg13g2_fill_2 FILLER_38_1166 ();
 sg13g2_fill_1 FILLER_38_1168 ();
 sg13g2_decap_8 FILLER_38_1179 ();
 sg13g2_fill_1 FILLER_38_1186 ();
 sg13g2_fill_1 FILLER_38_1209 ();
 sg13g2_fill_2 FILLER_38_1249 ();
 sg13g2_fill_1 FILLER_38_1251 ();
 sg13g2_fill_2 FILLER_38_1263 ();
 sg13g2_decap_8 FILLER_38_1270 ();
 sg13g2_decap_8 FILLER_38_1277 ();
 sg13g2_decap_8 FILLER_38_1284 ();
 sg13g2_decap_8 FILLER_38_1291 ();
 sg13g2_fill_1 FILLER_38_1298 ();
 sg13g2_fill_2 FILLER_38_1335 ();
 sg13g2_fill_1 FILLER_38_1337 ();
 sg13g2_fill_2 FILLER_38_1346 ();
 sg13g2_fill_1 FILLER_38_1353 ();
 sg13g2_fill_1 FILLER_38_1358 ();
 sg13g2_fill_1 FILLER_38_1363 ();
 sg13g2_fill_2 FILLER_38_1374 ();
 sg13g2_fill_1 FILLER_38_1376 ();
 sg13g2_decap_8 FILLER_38_1499 ();
 sg13g2_decap_8 FILLER_38_1506 ();
 sg13g2_fill_2 FILLER_38_1513 ();
 sg13g2_decap_8 FILLER_38_1519 ();
 sg13g2_fill_2 FILLER_38_1526 ();
 sg13g2_fill_1 FILLER_38_1532 ();
 sg13g2_fill_2 FILLER_38_1543 ();
 sg13g2_fill_1 FILLER_38_1545 ();
 sg13g2_fill_1 FILLER_38_1577 ();
 sg13g2_fill_2 FILLER_38_1644 ();
 sg13g2_fill_1 FILLER_38_1646 ();
 sg13g2_decap_8 FILLER_38_1673 ();
 sg13g2_decap_8 FILLER_38_1680 ();
 sg13g2_decap_8 FILLER_38_1687 ();
 sg13g2_decap_8 FILLER_38_1698 ();
 sg13g2_decap_8 FILLER_38_1705 ();
 sg13g2_decap_8 FILLER_38_1712 ();
 sg13g2_decap_4 FILLER_38_1719 ();
 sg13g2_fill_2 FILLER_38_1723 ();
 sg13g2_decap_8 FILLER_38_1751 ();
 sg13g2_decap_8 FILLER_38_1758 ();
 sg13g2_decap_8 FILLER_38_1765 ();
 sg13g2_fill_2 FILLER_38_1772 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_57 ();
 sg13g2_decap_4 FILLER_39_69 ();
 sg13g2_decap_4 FILLER_39_83 ();
 sg13g2_fill_2 FILLER_39_91 ();
 sg13g2_fill_1 FILLER_39_93 ();
 sg13g2_fill_2 FILLER_39_150 ();
 sg13g2_fill_2 FILLER_39_252 ();
 sg13g2_decap_4 FILLER_39_279 ();
 sg13g2_fill_1 FILLER_39_286 ();
 sg13g2_fill_2 FILLER_39_307 ();
 sg13g2_fill_2 FILLER_39_322 ();
 sg13g2_fill_1 FILLER_39_328 ();
 sg13g2_fill_1 FILLER_39_339 ();
 sg13g2_fill_1 FILLER_39_348 ();
 sg13g2_decap_4 FILLER_39_367 ();
 sg13g2_fill_1 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_fill_1 FILLER_39_401 ();
 sg13g2_fill_2 FILLER_39_406 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_decap_8 FILLER_39_466 ();
 sg13g2_decap_8 FILLER_39_473 ();
 sg13g2_decap_4 FILLER_39_480 ();
 sg13g2_fill_2 FILLER_39_484 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_decap_8 FILLER_39_497 ();
 sg13g2_fill_1 FILLER_39_504 ();
 sg13g2_decap_8 FILLER_39_509 ();
 sg13g2_decap_8 FILLER_39_520 ();
 sg13g2_fill_2 FILLER_39_527 ();
 sg13g2_fill_1 FILLER_39_529 ();
 sg13g2_fill_1 FILLER_39_534 ();
 sg13g2_fill_2 FILLER_39_556 ();
 sg13g2_fill_1 FILLER_39_632 ();
 sg13g2_fill_2 FILLER_39_641 ();
 sg13g2_fill_2 FILLER_39_647 ();
 sg13g2_fill_1 FILLER_39_672 ();
 sg13g2_decap_4 FILLER_39_698 ();
 sg13g2_fill_2 FILLER_39_702 ();
 sg13g2_fill_2 FILLER_39_709 ();
 sg13g2_fill_2 FILLER_39_751 ();
 sg13g2_fill_2 FILLER_39_763 ();
 sg13g2_fill_2 FILLER_39_775 ();
 sg13g2_decap_4 FILLER_39_781 ();
 sg13g2_fill_2 FILLER_39_789 ();
 sg13g2_decap_4 FILLER_39_801 ();
 sg13g2_decap_4 FILLER_39_837 ();
 sg13g2_fill_1 FILLER_39_849 ();
 sg13g2_fill_2 FILLER_39_894 ();
 sg13g2_fill_2 FILLER_39_958 ();
 sg13g2_decap_8 FILLER_39_996 ();
 sg13g2_decap_8 FILLER_39_1003 ();
 sg13g2_fill_1 FILLER_39_1010 ();
 sg13g2_fill_1 FILLER_39_1042 ();
 sg13g2_fill_1 FILLER_39_1068 ();
 sg13g2_fill_1 FILLER_39_1073 ();
 sg13g2_fill_2 FILLER_39_1079 ();
 sg13g2_decap_8 FILLER_39_1099 ();
 sg13g2_decap_8 FILLER_39_1106 ();
 sg13g2_decap_8 FILLER_39_1113 ();
 sg13g2_fill_2 FILLER_39_1120 ();
 sg13g2_decap_8 FILLER_39_1169 ();
 sg13g2_decap_4 FILLER_39_1176 ();
 sg13g2_fill_1 FILLER_39_1184 ();
 sg13g2_fill_1 FILLER_39_1189 ();
 sg13g2_fill_2 FILLER_39_1194 ();
 sg13g2_decap_8 FILLER_39_1230 ();
 sg13g2_decap_8 FILLER_39_1237 ();
 sg13g2_decap_8 FILLER_39_1244 ();
 sg13g2_decap_8 FILLER_39_1251 ();
 sg13g2_fill_2 FILLER_39_1258 ();
 sg13g2_fill_1 FILLER_39_1260 ();
 sg13g2_decap_8 FILLER_39_1273 ();
 sg13g2_fill_2 FILLER_39_1290 ();
 sg13g2_fill_1 FILLER_39_1292 ();
 sg13g2_decap_8 FILLER_39_1297 ();
 sg13g2_fill_1 FILLER_39_1304 ();
 sg13g2_decap_8 FILLER_39_1315 ();
 sg13g2_decap_4 FILLER_39_1322 ();
 sg13g2_decap_8 FILLER_39_1330 ();
 sg13g2_decap_8 FILLER_39_1337 ();
 sg13g2_decap_8 FILLER_39_1344 ();
 sg13g2_decap_8 FILLER_39_1351 ();
 sg13g2_fill_2 FILLER_39_1358 ();
 sg13g2_decap_4 FILLER_39_1391 ();
 sg13g2_fill_2 FILLER_39_1399 ();
 sg13g2_fill_2 FILLER_39_1411 ();
 sg13g2_decap_4 FILLER_39_1423 ();
 sg13g2_fill_1 FILLER_39_1432 ();
 sg13g2_decap_8 FILLER_39_1488 ();
 sg13g2_decap_4 FILLER_39_1495 ();
 sg13g2_decap_8 FILLER_39_1503 ();
 sg13g2_fill_2 FILLER_39_1510 ();
 sg13g2_fill_1 FILLER_39_1512 ();
 sg13g2_decap_4 FILLER_39_1518 ();
 sg13g2_fill_2 FILLER_39_1526 ();
 sg13g2_fill_1 FILLER_39_1528 ();
 sg13g2_fill_1 FILLER_39_1534 ();
 sg13g2_decap_8 FILLER_39_1540 ();
 sg13g2_fill_1 FILLER_39_1552 ();
 sg13g2_fill_1 FILLER_39_1557 ();
 sg13g2_fill_1 FILLER_39_1562 ();
 sg13g2_fill_1 FILLER_39_1568 ();
 sg13g2_decap_8 FILLER_39_1636 ();
 sg13g2_decap_4 FILLER_39_1643 ();
 sg13g2_fill_2 FILLER_39_1647 ();
 sg13g2_decap_8 FILLER_39_1653 ();
 sg13g2_decap_8 FILLER_39_1660 ();
 sg13g2_decap_8 FILLER_39_1667 ();
 sg13g2_decap_8 FILLER_39_1674 ();
 sg13g2_fill_2 FILLER_39_1681 ();
 sg13g2_decap_8 FILLER_39_1704 ();
 sg13g2_decap_8 FILLER_39_1711 ();
 sg13g2_decap_4 FILLER_39_1718 ();
 sg13g2_decap_8 FILLER_39_1736 ();
 sg13g2_decap_8 FILLER_39_1743 ();
 sg13g2_decap_8 FILLER_39_1750 ();
 sg13g2_decap_8 FILLER_39_1757 ();
 sg13g2_decap_8 FILLER_39_1764 ();
 sg13g2_fill_2 FILLER_39_1771 ();
 sg13g2_fill_1 FILLER_39_1773 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_9 ();
 sg13g2_fill_1 FILLER_40_19 ();
 sg13g2_fill_1 FILLER_40_24 ();
 sg13g2_decap_8 FILLER_40_86 ();
 sg13g2_decap_4 FILLER_40_93 ();
 sg13g2_fill_1 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_201 ();
 sg13g2_decap_8 FILLER_40_207 ();
 sg13g2_fill_2 FILLER_40_214 ();
 sg13g2_fill_1 FILLER_40_216 ();
 sg13g2_fill_1 FILLER_40_221 ();
 sg13g2_decap_8 FILLER_40_226 ();
 sg13g2_decap_4 FILLER_40_233 ();
 sg13g2_fill_1 FILLER_40_237 ();
 sg13g2_fill_1 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_270 ();
 sg13g2_fill_2 FILLER_40_281 ();
 sg13g2_fill_2 FILLER_40_333 ();
 sg13g2_fill_1 FILLER_40_369 ();
 sg13g2_decap_4 FILLER_40_383 ();
 sg13g2_fill_1 FILLER_40_391 ();
 sg13g2_decap_8 FILLER_40_405 ();
 sg13g2_decap_4 FILLER_40_412 ();
 sg13g2_fill_2 FILLER_40_416 ();
 sg13g2_fill_2 FILLER_40_428 ();
 sg13g2_fill_1 FILLER_40_430 ();
 sg13g2_decap_8 FILLER_40_439 ();
 sg13g2_decap_8 FILLER_40_446 ();
 sg13g2_decap_8 FILLER_40_453 ();
 sg13g2_decap_8 FILLER_40_460 ();
 sg13g2_decap_4 FILLER_40_467 ();
 sg13g2_fill_2 FILLER_40_575 ();
 sg13g2_fill_1 FILLER_40_577 ();
 sg13g2_decap_8 FILLER_40_582 ();
 sg13g2_decap_8 FILLER_40_594 ();
 sg13g2_decap_8 FILLER_40_601 ();
 sg13g2_decap_8 FILLER_40_608 ();
 sg13g2_fill_2 FILLER_40_627 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_4 FILLER_40_644 ();
 sg13g2_fill_2 FILLER_40_648 ();
 sg13g2_fill_2 FILLER_40_658 ();
 sg13g2_fill_1 FILLER_40_665 ();
 sg13g2_fill_2 FILLER_40_676 ();
 sg13g2_decap_4 FILLER_40_686 ();
 sg13g2_fill_2 FILLER_40_690 ();
 sg13g2_decap_4 FILLER_40_696 ();
 sg13g2_decap_8 FILLER_40_705 ();
 sg13g2_fill_1 FILLER_40_712 ();
 sg13g2_decap_8 FILLER_40_723 ();
 sg13g2_fill_1 FILLER_40_730 ();
 sg13g2_fill_2 FILLER_40_827 ();
 sg13g2_decap_4 FILLER_40_847 ();
 sg13g2_fill_2 FILLER_40_864 ();
 sg13g2_decap_8 FILLER_40_870 ();
 sg13g2_decap_8 FILLER_40_877 ();
 sg13g2_decap_8 FILLER_40_884 ();
 sg13g2_fill_1 FILLER_40_891 ();
 sg13g2_decap_4 FILLER_40_905 ();
 sg13g2_fill_2 FILLER_40_909 ();
 sg13g2_fill_1 FILLER_40_916 ();
 sg13g2_fill_1 FILLER_40_921 ();
 sg13g2_decap_8 FILLER_40_932 ();
 sg13g2_fill_1 FILLER_40_939 ();
 sg13g2_decap_4 FILLER_40_944 ();
 sg13g2_decap_4 FILLER_40_960 ();
 sg13g2_decap_4 FILLER_40_1016 ();
 sg13g2_fill_1 FILLER_40_1020 ();
 sg13g2_decap_8 FILLER_40_1061 ();
 sg13g2_decap_4 FILLER_40_1068 ();
 sg13g2_fill_2 FILLER_40_1072 ();
 sg13g2_fill_1 FILLER_40_1080 ();
 sg13g2_decap_8 FILLER_40_1088 ();
 sg13g2_decap_8 FILLER_40_1095 ();
 sg13g2_decap_8 FILLER_40_1102 ();
 sg13g2_fill_2 FILLER_40_1109 ();
 sg13g2_fill_1 FILLER_40_1132 ();
 sg13g2_fill_1 FILLER_40_1154 ();
 sg13g2_decap_8 FILLER_40_1189 ();
 sg13g2_fill_2 FILLER_40_1196 ();
 sg13g2_fill_2 FILLER_40_1208 ();
 sg13g2_decap_8 FILLER_40_1225 ();
 sg13g2_decap_4 FILLER_40_1251 ();
 sg13g2_fill_1 FILLER_40_1255 ();
 sg13g2_fill_2 FILLER_40_1282 ();
 sg13g2_fill_1 FILLER_40_1284 ();
 sg13g2_fill_2 FILLER_40_1337 ();
 sg13g2_decap_8 FILLER_40_1345 ();
 sg13g2_fill_2 FILLER_40_1352 ();
 sg13g2_fill_1 FILLER_40_1354 ();
 sg13g2_decap_4 FILLER_40_1359 ();
 sg13g2_fill_1 FILLER_40_1363 ();
 sg13g2_decap_8 FILLER_40_1395 ();
 sg13g2_decap_8 FILLER_40_1402 ();
 sg13g2_decap_8 FILLER_40_1409 ();
 sg13g2_fill_1 FILLER_40_1446 ();
 sg13g2_fill_2 FILLER_40_1473 ();
 sg13g2_decap_8 FILLER_40_1479 ();
 sg13g2_decap_8 FILLER_40_1486 ();
 sg13g2_fill_2 FILLER_40_1493 ();
 sg13g2_fill_2 FILLER_40_1499 ();
 sg13g2_fill_1 FILLER_40_1501 ();
 sg13g2_decap_4 FILLER_40_1506 ();
 sg13g2_fill_2 FILLER_40_1510 ();
 sg13g2_decap_4 FILLER_40_1518 ();
 sg13g2_fill_1 FILLER_40_1522 ();
 sg13g2_decap_8 FILLER_40_1528 ();
 sg13g2_decap_4 FILLER_40_1535 ();
 sg13g2_fill_2 FILLER_40_1539 ();
 sg13g2_fill_2 FILLER_40_1553 ();
 sg13g2_fill_1 FILLER_40_1555 ();
 sg13g2_decap_8 FILLER_40_1562 ();
 sg13g2_decap_8 FILLER_40_1569 ();
 sg13g2_decap_8 FILLER_40_1576 ();
 sg13g2_fill_2 FILLER_40_1583 ();
 sg13g2_decap_8 FILLER_40_1593 ();
 sg13g2_decap_8 FILLER_40_1600 ();
 sg13g2_decap_8 FILLER_40_1607 ();
 sg13g2_fill_2 FILLER_40_1614 ();
 sg13g2_fill_1 FILLER_40_1616 ();
 sg13g2_decap_4 FILLER_40_1621 ();
 sg13g2_decap_8 FILLER_40_1629 ();
 sg13g2_decap_4 FILLER_40_1636 ();
 sg13g2_decap_8 FILLER_40_1673 ();
 sg13g2_decap_4 FILLER_40_1680 ();
 sg13g2_fill_1 FILLER_40_1684 ();
 sg13g2_fill_1 FILLER_40_1773 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_45 ();
 sg13g2_decap_8 FILLER_41_76 ();
 sg13g2_decap_8 FILLER_41_83 ();
 sg13g2_fill_2 FILLER_41_90 ();
 sg13g2_decap_8 FILLER_41_102 ();
 sg13g2_decap_8 FILLER_41_131 ();
 sg13g2_decap_4 FILLER_41_138 ();
 sg13g2_fill_2 FILLER_41_142 ();
 sg13g2_fill_2 FILLER_41_169 ();
 sg13g2_fill_1 FILLER_41_171 ();
 sg13g2_decap_4 FILLER_41_178 ();
 sg13g2_fill_1 FILLER_41_182 ();
 sg13g2_fill_2 FILLER_41_218 ();
 sg13g2_fill_2 FILLER_41_224 ();
 sg13g2_fill_1 FILLER_41_226 ();
 sg13g2_decap_8 FILLER_41_240 ();
 sg13g2_decap_4 FILLER_41_260 ();
 sg13g2_fill_1 FILLER_41_264 ();
 sg13g2_fill_1 FILLER_41_291 ();
 sg13g2_fill_1 FILLER_41_328 ();
 sg13g2_fill_2 FILLER_41_355 ();
 sg13g2_decap_4 FILLER_41_365 ();
 sg13g2_fill_2 FILLER_41_369 ();
 sg13g2_fill_2 FILLER_41_397 ();
 sg13g2_decap_8 FILLER_41_404 ();
 sg13g2_fill_2 FILLER_41_411 ();
 sg13g2_fill_1 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_450 ();
 sg13g2_decap_8 FILLER_41_457 ();
 sg13g2_decap_8 FILLER_41_464 ();
 sg13g2_decap_8 FILLER_41_471 ();
 sg13g2_fill_2 FILLER_41_478 ();
 sg13g2_fill_1 FILLER_41_530 ();
 sg13g2_decap_4 FILLER_41_587 ();
 sg13g2_fill_1 FILLER_41_635 ();
 sg13g2_fill_2 FILLER_41_644 ();
 sg13g2_decap_4 FILLER_41_660 ();
 sg13g2_fill_1 FILLER_41_664 ();
 sg13g2_decap_4 FILLER_41_669 ();
 sg13g2_fill_1 FILLER_41_673 ();
 sg13g2_decap_4 FILLER_41_708 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_decap_8 FILLER_41_759 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_decap_4 FILLER_41_773 ();
 sg13g2_fill_1 FILLER_41_777 ();
 sg13g2_fill_2 FILLER_41_787 ();
 sg13g2_fill_1 FILLER_41_789 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_decap_8 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_decap_4 FILLER_41_875 ();
 sg13g2_decap_4 FILLER_41_892 ();
 sg13g2_fill_2 FILLER_41_896 ();
 sg13g2_decap_8 FILLER_41_934 ();
 sg13g2_decap_8 FILLER_41_941 ();
 sg13g2_decap_8 FILLER_41_948 ();
 sg13g2_decap_8 FILLER_41_955 ();
 sg13g2_fill_1 FILLER_41_962 ();
 sg13g2_fill_1 FILLER_41_968 ();
 sg13g2_fill_1 FILLER_41_973 ();
 sg13g2_fill_2 FILLER_41_984 ();
 sg13g2_fill_2 FILLER_41_991 ();
 sg13g2_decap_8 FILLER_41_1005 ();
 sg13g2_decap_8 FILLER_41_1012 ();
 sg13g2_fill_2 FILLER_41_1019 ();
 sg13g2_fill_1 FILLER_41_1021 ();
 sg13g2_decap_4 FILLER_41_1036 ();
 sg13g2_decap_8 FILLER_41_1088 ();
 sg13g2_decap_8 FILLER_41_1095 ();
 sg13g2_fill_1 FILLER_41_1102 ();
 sg13g2_fill_1 FILLER_41_1158 ();
 sg13g2_decap_8 FILLER_41_1189 ();
 sg13g2_decap_8 FILLER_41_1196 ();
 sg13g2_decap_8 FILLER_41_1203 ();
 sg13g2_decap_8 FILLER_41_1210 ();
 sg13g2_decap_4 FILLER_41_1217 ();
 sg13g2_fill_1 FILLER_41_1221 ();
 sg13g2_decap_4 FILLER_41_1232 ();
 sg13g2_decap_4 FILLER_41_1245 ();
 sg13g2_fill_1 FILLER_41_1249 ();
 sg13g2_decap_4 FILLER_41_1260 ();
 sg13g2_decap_8 FILLER_41_1268 ();
 sg13g2_fill_2 FILLER_41_1275 ();
 sg13g2_fill_1 FILLER_41_1277 ();
 sg13g2_decap_8 FILLER_41_1299 ();
 sg13g2_decap_4 FILLER_41_1306 ();
 sg13g2_fill_2 FILLER_41_1310 ();
 sg13g2_decap_8 FILLER_41_1320 ();
 sg13g2_decap_8 FILLER_41_1327 ();
 sg13g2_decap_8 FILLER_41_1334 ();
 sg13g2_decap_8 FILLER_41_1341 ();
 sg13g2_decap_4 FILLER_41_1348 ();
 sg13g2_fill_1 FILLER_41_1352 ();
 sg13g2_fill_2 FILLER_41_1363 ();
 sg13g2_fill_1 FILLER_41_1365 ();
 sg13g2_decap_4 FILLER_41_1376 ();
 sg13g2_fill_1 FILLER_41_1380 ();
 sg13g2_decap_4 FILLER_41_1407 ();
 sg13g2_fill_1 FILLER_41_1411 ();
 sg13g2_fill_2 FILLER_41_1422 ();
 sg13g2_fill_1 FILLER_41_1424 ();
 sg13g2_decap_4 FILLER_41_1429 ();
 sg13g2_fill_2 FILLER_41_1433 ();
 sg13g2_fill_2 FILLER_41_1496 ();
 sg13g2_fill_1 FILLER_41_1498 ();
 sg13g2_fill_2 FILLER_41_1504 ();
 sg13g2_fill_1 FILLER_41_1506 ();
 sg13g2_decap_8 FILLER_41_1511 ();
 sg13g2_decap_4 FILLER_41_1518 ();
 sg13g2_fill_2 FILLER_41_1522 ();
 sg13g2_decap_8 FILLER_41_1545 ();
 sg13g2_decap_4 FILLER_41_1552 ();
 sg13g2_fill_2 FILLER_41_1556 ();
 sg13g2_decap_8 FILLER_41_1562 ();
 sg13g2_fill_1 FILLER_41_1569 ();
 sg13g2_decap_8 FILLER_41_1576 ();
 sg13g2_fill_1 FILLER_41_1583 ();
 sg13g2_decap_8 FILLER_41_1594 ();
 sg13g2_decap_4 FILLER_41_1601 ();
 sg13g2_fill_2 FILLER_41_1605 ();
 sg13g2_decap_8 FILLER_41_1615 ();
 sg13g2_decap_8 FILLER_41_1622 ();
 sg13g2_decap_4 FILLER_41_1629 ();
 sg13g2_fill_1 FILLER_41_1633 ();
 sg13g2_decap_8 FILLER_41_1670 ();
 sg13g2_fill_2 FILLER_41_1677 ();
 sg13g2_fill_1 FILLER_41_1679 ();
 sg13g2_fill_2 FILLER_41_1734 ();
 sg13g2_decap_8 FILLER_41_1766 ();
 sg13g2_fill_1 FILLER_41_1773 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_4 FILLER_42_14 ();
 sg13g2_fill_2 FILLER_42_28 ();
 sg13g2_fill_1 FILLER_42_30 ();
 sg13g2_fill_2 FILLER_42_35 ();
 sg13g2_fill_1 FILLER_42_47 ();
 sg13g2_fill_2 FILLER_42_54 ();
 sg13g2_fill_1 FILLER_42_76 ();
 sg13g2_decap_4 FILLER_42_81 ();
 sg13g2_fill_2 FILLER_42_100 ();
 sg13g2_fill_2 FILLER_42_140 ();
 sg13g2_fill_1 FILLER_42_142 ();
 sg13g2_fill_2 FILLER_42_204 ();
 sg13g2_fill_2 FILLER_42_241 ();
 sg13g2_decap_8 FILLER_42_247 ();
 sg13g2_fill_2 FILLER_42_254 ();
 sg13g2_fill_1 FILLER_42_256 ();
 sg13g2_fill_2 FILLER_42_261 ();
 sg13g2_decap_4 FILLER_42_269 ();
 sg13g2_decap_4 FILLER_42_277 ();
 sg13g2_decap_4 FILLER_42_307 ();
 sg13g2_fill_2 FILLER_42_315 ();
 sg13g2_fill_1 FILLER_42_317 ();
 sg13g2_decap_4 FILLER_42_322 ();
 sg13g2_fill_2 FILLER_42_326 ();
 sg13g2_fill_2 FILLER_42_338 ();
 sg13g2_decap_8 FILLER_42_348 ();
 sg13g2_decap_8 FILLER_42_355 ();
 sg13g2_decap_4 FILLER_42_362 ();
 sg13g2_fill_2 FILLER_42_366 ();
 sg13g2_fill_1 FILLER_42_381 ();
 sg13g2_fill_2 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_452 ();
 sg13g2_decap_8 FILLER_42_459 ();
 sg13g2_decap_4 FILLER_42_466 ();
 sg13g2_decap_4 FILLER_42_510 ();
 sg13g2_fill_2 FILLER_42_541 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_564 ();
 sg13g2_decap_8 FILLER_42_628 ();
 sg13g2_fill_1 FILLER_42_635 ();
 sg13g2_fill_2 FILLER_42_714 ();
 sg13g2_decap_8 FILLER_42_750 ();
 sg13g2_decap_8 FILLER_42_757 ();
 sg13g2_decap_8 FILLER_42_764 ();
 sg13g2_decap_8 FILLER_42_771 ();
 sg13g2_fill_2 FILLER_42_778 ();
 sg13g2_fill_2 FILLER_42_806 ();
 sg13g2_fill_2 FILLER_42_812 ();
 sg13g2_fill_1 FILLER_42_814 ();
 sg13g2_decap_8 FILLER_42_819 ();
 sg13g2_decap_4 FILLER_42_826 ();
 sg13g2_fill_1 FILLER_42_830 ();
 sg13g2_fill_2 FILLER_42_841 ();
 sg13g2_fill_1 FILLER_42_843 ();
 sg13g2_decap_8 FILLER_42_870 ();
 sg13g2_decap_8 FILLER_42_877 ();
 sg13g2_decap_8 FILLER_42_884 ();
 sg13g2_decap_4 FILLER_42_891 ();
 sg13g2_fill_1 FILLER_42_895 ();
 sg13g2_decap_8 FILLER_42_930 ();
 sg13g2_decap_8 FILLER_42_937 ();
 sg13g2_decap_4 FILLER_42_944 ();
 sg13g2_decap_8 FILLER_42_952 ();
 sg13g2_fill_1 FILLER_42_959 ();
 sg13g2_decap_4 FILLER_42_970 ();
 sg13g2_fill_1 FILLER_42_974 ();
 sg13g2_decap_4 FILLER_42_979 ();
 sg13g2_decap_8 FILLER_42_993 ();
 sg13g2_decap_8 FILLER_42_1000 ();
 sg13g2_decap_8 FILLER_42_1007 ();
 sg13g2_decap_8 FILLER_42_1014 ();
 sg13g2_decap_4 FILLER_42_1021 ();
 sg13g2_fill_1 FILLER_42_1025 ();
 sg13g2_decap_8 FILLER_42_1052 ();
 sg13g2_decap_4 FILLER_42_1059 ();
 sg13g2_fill_1 FILLER_42_1063 ();
 sg13g2_decap_8 FILLER_42_1085 ();
 sg13g2_fill_1 FILLER_42_1092 ();
 sg13g2_decap_8 FILLER_42_1101 ();
 sg13g2_decap_8 FILLER_42_1160 ();
 sg13g2_fill_1 FILLER_42_1167 ();
 sg13g2_decap_8 FILLER_42_1194 ();
 sg13g2_decap_8 FILLER_42_1201 ();
 sg13g2_decap_8 FILLER_42_1208 ();
 sg13g2_fill_1 FILLER_42_1215 ();
 sg13g2_fill_2 FILLER_42_1220 ();
 sg13g2_fill_1 FILLER_42_1222 ();
 sg13g2_decap_4 FILLER_42_1270 ();
 sg13g2_decap_8 FILLER_42_1321 ();
 sg13g2_decap_8 FILLER_42_1328 ();
 sg13g2_decap_8 FILLER_42_1335 ();
 sg13g2_decap_8 FILLER_42_1342 ();
 sg13g2_decap_4 FILLER_42_1349 ();
 sg13g2_fill_2 FILLER_42_1379 ();
 sg13g2_fill_2 FILLER_42_1407 ();
 sg13g2_decap_8 FILLER_42_1445 ();
 sg13g2_fill_2 FILLER_42_1452 ();
 sg13g2_fill_1 FILLER_42_1454 ();
 sg13g2_fill_2 FILLER_42_1472 ();
 sg13g2_fill_1 FILLER_42_1493 ();
 sg13g2_decap_8 FILLER_42_1502 ();
 sg13g2_fill_1 FILLER_42_1509 ();
 sg13g2_fill_2 FILLER_42_1524 ();
 sg13g2_fill_1 FILLER_42_1526 ();
 sg13g2_fill_1 FILLER_42_1553 ();
 sg13g2_fill_2 FILLER_42_1559 ();
 sg13g2_fill_1 FILLER_42_1561 ();
 sg13g2_decap_4 FILLER_42_1628 ();
 sg13g2_fill_2 FILLER_42_1632 ();
 sg13g2_decap_4 FILLER_42_1642 ();
 sg13g2_fill_2 FILLER_42_1650 ();
 sg13g2_fill_2 FILLER_42_1761 ();
 sg13g2_decap_8 FILLER_42_1767 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_9 ();
 sg13g2_fill_1 FILLER_43_36 ();
 sg13g2_fill_1 FILLER_43_47 ();
 sg13g2_fill_1 FILLER_43_90 ();
 sg13g2_fill_1 FILLER_43_101 ();
 sg13g2_fill_1 FILLER_43_112 ();
 sg13g2_fill_2 FILLER_43_117 ();
 sg13g2_fill_2 FILLER_43_123 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_fill_1 FILLER_43_166 ();
 sg13g2_decap_4 FILLER_43_210 ();
 sg13g2_fill_1 FILLER_43_214 ();
 sg13g2_decap_4 FILLER_43_219 ();
 sg13g2_fill_2 FILLER_43_223 ();
 sg13g2_fill_2 FILLER_43_261 ();
 sg13g2_decap_8 FILLER_43_268 ();
 sg13g2_decap_8 FILLER_43_275 ();
 sg13g2_decap_4 FILLER_43_282 ();
 sg13g2_fill_2 FILLER_43_286 ();
 sg13g2_decap_8 FILLER_43_338 ();
 sg13g2_decap_8 FILLER_43_345 ();
 sg13g2_decap_8 FILLER_43_352 ();
 sg13g2_decap_8 FILLER_43_359 ();
 sg13g2_decap_8 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_373 ();
 sg13g2_decap_8 FILLER_43_412 ();
 sg13g2_fill_2 FILLER_43_419 ();
 sg13g2_decap_8 FILLER_43_457 ();
 sg13g2_decap_8 FILLER_43_464 ();
 sg13g2_fill_2 FILLER_43_471 ();
 sg13g2_fill_1 FILLER_43_473 ();
 sg13g2_decap_8 FILLER_43_478 ();
 sg13g2_fill_2 FILLER_43_485 ();
 sg13g2_fill_1 FILLER_43_487 ();
 sg13g2_decap_8 FILLER_43_548 ();
 sg13g2_decap_8 FILLER_43_555 ();
 sg13g2_decap_8 FILLER_43_562 ();
 sg13g2_decap_8 FILLER_43_569 ();
 sg13g2_decap_4 FILLER_43_576 ();
 sg13g2_fill_1 FILLER_43_580 ();
 sg13g2_decap_8 FILLER_43_607 ();
 sg13g2_fill_2 FILLER_43_614 ();
 sg13g2_decap_8 FILLER_43_673 ();
 sg13g2_decap_8 FILLER_43_680 ();
 sg13g2_fill_2 FILLER_43_687 ();
 sg13g2_fill_1 FILLER_43_689 ();
 sg13g2_fill_2 FILLER_43_695 ();
 sg13g2_decap_4 FILLER_43_701 ();
 sg13g2_fill_2 FILLER_43_757 ();
 sg13g2_decap_4 FILLER_43_785 ();
 sg13g2_fill_1 FILLER_43_793 ();
 sg13g2_decap_8 FILLER_43_804 ();
 sg13g2_fill_1 FILLER_43_811 ();
 sg13g2_fill_1 FILLER_43_843 ();
 sg13g2_decap_8 FILLER_43_870 ();
 sg13g2_decap_8 FILLER_43_877 ();
 sg13g2_decap_8 FILLER_43_884 ();
 sg13g2_decap_8 FILLER_43_891 ();
 sg13g2_decap_4 FILLER_43_898 ();
 sg13g2_fill_2 FILLER_43_902 ();
 sg13g2_decap_4 FILLER_43_914 ();
 sg13g2_decap_8 FILLER_43_922 ();
 sg13g2_fill_1 FILLER_43_929 ();
 sg13g2_fill_2 FILLER_43_966 ();
 sg13g2_fill_2 FILLER_43_998 ();
 sg13g2_fill_1 FILLER_43_1000 ();
 sg13g2_decap_4 FILLER_43_1008 ();
 sg13g2_fill_2 FILLER_43_1012 ();
 sg13g2_fill_2 FILLER_43_1050 ();
 sg13g2_decap_4 FILLER_43_1062 ();
 sg13g2_fill_2 FILLER_43_1066 ();
 sg13g2_decap_8 FILLER_43_1089 ();
 sg13g2_fill_1 FILLER_43_1096 ();
 sg13g2_decap_8 FILLER_43_1202 ();
 sg13g2_fill_2 FILLER_43_1209 ();
 sg13g2_decap_4 FILLER_43_1261 ();
 sg13g2_fill_2 FILLER_43_1265 ();
 sg13g2_decap_4 FILLER_43_1277 ();
 sg13g2_fill_2 FILLER_43_1285 ();
 sg13g2_decap_8 FILLER_43_1343 ();
 sg13g2_decap_8 FILLER_43_1350 ();
 sg13g2_fill_2 FILLER_43_1357 ();
 sg13g2_decap_8 FILLER_43_1401 ();
 sg13g2_decap_4 FILLER_43_1408 ();
 sg13g2_fill_2 FILLER_43_1412 ();
 sg13g2_decap_8 FILLER_43_1461 ();
 sg13g2_decap_8 FILLER_43_1468 ();
 sg13g2_fill_2 FILLER_43_1475 ();
 sg13g2_fill_1 FILLER_43_1477 ();
 sg13g2_decap_8 FILLER_43_1484 ();
 sg13g2_fill_1 FILLER_43_1568 ();
 sg13g2_decap_4 FILLER_43_1609 ();
 sg13g2_fill_1 FILLER_43_1613 ();
 sg13g2_decap_8 FILLER_43_1624 ();
 sg13g2_decap_4 FILLER_43_1631 ();
 sg13g2_fill_1 FILLER_43_1635 ();
 sg13g2_decap_8 FILLER_43_1676 ();
 sg13g2_decap_8 FILLER_43_1683 ();
 sg13g2_decap_4 FILLER_43_1690 ();
 sg13g2_fill_1 FILLER_43_1694 ();
 sg13g2_decap_8 FILLER_43_1699 ();
 sg13g2_fill_2 FILLER_43_1706 ();
 sg13g2_fill_1 FILLER_43_1708 ();
 sg13g2_decap_4 FILLER_43_1719 ();
 sg13g2_fill_2 FILLER_43_1723 ();
 sg13g2_decap_8 FILLER_43_1759 ();
 sg13g2_decap_8 FILLER_43_1766 ();
 sg13g2_fill_1 FILLER_43_1773 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_95 ();
 sg13g2_decap_4 FILLER_44_107 ();
 sg13g2_fill_2 FILLER_44_137 ();
 sg13g2_decap_8 FILLER_44_149 ();
 sg13g2_fill_1 FILLER_44_156 ();
 sg13g2_fill_2 FILLER_44_215 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_fill_1 FILLER_44_223 ();
 sg13g2_fill_2 FILLER_44_242 ();
 sg13g2_fill_2 FILLER_44_274 ();
 sg13g2_fill_1 FILLER_44_276 ();
 sg13g2_fill_1 FILLER_44_303 ();
 sg13g2_decap_8 FILLER_44_330 ();
 sg13g2_fill_2 FILLER_44_337 ();
 sg13g2_decap_4 FILLER_44_349 ();
 sg13g2_fill_2 FILLER_44_353 ();
 sg13g2_fill_2 FILLER_44_363 ();
 sg13g2_fill_1 FILLER_44_365 ();
 sg13g2_decap_8 FILLER_44_372 ();
 sg13g2_decap_8 FILLER_44_379 ();
 sg13g2_decap_8 FILLER_44_386 ();
 sg13g2_decap_4 FILLER_44_393 ();
 sg13g2_fill_2 FILLER_44_397 ();
 sg13g2_decap_8 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_410 ();
 sg13g2_decap_8 FILLER_44_417 ();
 sg13g2_decap_8 FILLER_44_424 ();
 sg13g2_fill_2 FILLER_44_431 ();
 sg13g2_fill_1 FILLER_44_437 ();
 sg13g2_decap_8 FILLER_44_474 ();
 sg13g2_decap_8 FILLER_44_481 ();
 sg13g2_decap_4 FILLER_44_488 ();
 sg13g2_fill_1 FILLER_44_492 ();
 sg13g2_decap_4 FILLER_44_520 ();
 sg13g2_fill_2 FILLER_44_524 ();
 sg13g2_decap_8 FILLER_44_556 ();
 sg13g2_decap_8 FILLER_44_563 ();
 sg13g2_decap_8 FILLER_44_570 ();
 sg13g2_decap_8 FILLER_44_577 ();
 sg13g2_fill_2 FILLER_44_584 ();
 sg13g2_fill_1 FILLER_44_590 ();
 sg13g2_fill_2 FILLER_44_595 ();
 sg13g2_fill_1 FILLER_44_633 ();
 sg13g2_fill_1 FILLER_44_639 ();
 sg13g2_decap_8 FILLER_44_657 ();
 sg13g2_decap_8 FILLER_44_664 ();
 sg13g2_decap_8 FILLER_44_671 ();
 sg13g2_decap_8 FILLER_44_678 ();
 sg13g2_fill_2 FILLER_44_685 ();
 sg13g2_fill_1 FILLER_44_687 ();
 sg13g2_decap_4 FILLER_44_693 ();
 sg13g2_fill_1 FILLER_44_697 ();
 sg13g2_fill_1 FILLER_44_702 ();
 sg13g2_decap_8 FILLER_44_733 ();
 sg13g2_fill_1 FILLER_44_740 ();
 sg13g2_decap_4 FILLER_44_745 ();
 sg13g2_fill_1 FILLER_44_767 ();
 sg13g2_decap_4 FILLER_44_772 ();
 sg13g2_decap_8 FILLER_44_802 ();
 sg13g2_decap_4 FILLER_44_809 ();
 sg13g2_fill_1 FILLER_44_813 ();
 sg13g2_decap_8 FILLER_44_874 ();
 sg13g2_fill_1 FILLER_44_881 ();
 sg13g2_fill_2 FILLER_44_918 ();
 sg13g2_fill_1 FILLER_44_920 ();
 sg13g2_fill_1 FILLER_44_924 ();
 sg13g2_fill_1 FILLER_44_938 ();
 sg13g2_decap_4 FILLER_44_948 ();
 sg13g2_fill_1 FILLER_44_971 ();
 sg13g2_fill_2 FILLER_44_982 ();
 sg13g2_fill_1 FILLER_44_984 ();
 sg13g2_fill_1 FILLER_44_1060 ();
 sg13g2_decap_8 FILLER_44_1082 ();
 sg13g2_decap_8 FILLER_44_1089 ();
 sg13g2_decap_4 FILLER_44_1096 ();
 sg13g2_fill_1 FILLER_44_1110 ();
 sg13g2_fill_2 FILLER_44_1115 ();
 sg13g2_fill_1 FILLER_44_1127 ();
 sg13g2_fill_1 FILLER_44_1132 ();
 sg13g2_decap_8 FILLER_44_1146 ();
 sg13g2_fill_2 FILLER_44_1153 ();
 sg13g2_decap_8 FILLER_44_1165 ();
 sg13g2_decap_8 FILLER_44_1172 ();
 sg13g2_fill_1 FILLER_44_1179 ();
 sg13g2_decap_8 FILLER_44_1188 ();
 sg13g2_fill_2 FILLER_44_1195 ();
 sg13g2_fill_1 FILLER_44_1197 ();
 sg13g2_fill_2 FILLER_44_1249 ();
 sg13g2_fill_2 FILLER_44_1277 ();
 sg13g2_fill_2 FILLER_44_1289 ();
 sg13g2_fill_1 FILLER_44_1291 ();
 sg13g2_fill_2 FILLER_44_1302 ();
 sg13g2_fill_1 FILLER_44_1304 ();
 sg13g2_decap_8 FILLER_44_1335 ();
 sg13g2_decap_8 FILLER_44_1342 ();
 sg13g2_decap_8 FILLER_44_1349 ();
 sg13g2_decap_8 FILLER_44_1356 ();
 sg13g2_decap_8 FILLER_44_1363 ();
 sg13g2_fill_1 FILLER_44_1370 ();
 sg13g2_decap_8 FILLER_44_1391 ();
 sg13g2_fill_2 FILLER_44_1398 ();
 sg13g2_fill_1 FILLER_44_1400 ();
 sg13g2_fill_2 FILLER_44_1454 ();
 sg13g2_decap_8 FILLER_44_1482 ();
 sg13g2_decap_4 FILLER_44_1489 ();
 sg13g2_fill_1 FILLER_44_1493 ();
 sg13g2_decap_4 FILLER_44_1544 ();
 sg13g2_fill_2 FILLER_44_1548 ();
 sg13g2_decap_4 FILLER_44_1554 ();
 sg13g2_fill_1 FILLER_44_1558 ();
 sg13g2_fill_1 FILLER_44_1580 ();
 sg13g2_fill_1 FILLER_44_1585 ();
 sg13g2_fill_1 FILLER_44_1590 ();
 sg13g2_fill_1 FILLER_44_1682 ();
 sg13g2_fill_2 FILLER_44_1693 ();
 sg13g2_fill_2 FILLER_44_1716 ();
 sg13g2_fill_2 FILLER_44_1723 ();
 sg13g2_fill_1 FILLER_44_1725 ();
 sg13g2_decap_8 FILLER_44_1766 ();
 sg13g2_fill_1 FILLER_44_1773 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_9 ();
 sg13g2_fill_1 FILLER_45_36 ();
 sg13g2_fill_1 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_74 ();
 sg13g2_fill_2 FILLER_45_90 ();
 sg13g2_fill_1 FILLER_45_92 ();
 sg13g2_fill_2 FILLER_45_97 ();
 sg13g2_fill_1 FILLER_45_99 ();
 sg13g2_decap_4 FILLER_45_170 ();
 sg13g2_fill_2 FILLER_45_174 ();
 sg13g2_fill_2 FILLER_45_179 ();
 sg13g2_fill_2 FILLER_45_231 ();
 sg13g2_fill_1 FILLER_45_233 ();
 sg13g2_decap_8 FILLER_45_237 ();
 sg13g2_decap_8 FILLER_45_244 ();
 sg13g2_decap_4 FILLER_45_251 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_fill_1 FILLER_45_294 ();
 sg13g2_fill_2 FILLER_45_321 ();
 sg13g2_decap_8 FILLER_45_387 ();
 sg13g2_decap_8 FILLER_45_394 ();
 sg13g2_decap_4 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_405 ();
 sg13g2_decap_8 FILLER_45_419 ();
 sg13g2_decap_8 FILLER_45_426 ();
 sg13g2_fill_1 FILLER_45_447 ();
 sg13g2_fill_1 FILLER_45_474 ();
 sg13g2_decap_8 FILLER_45_479 ();
 sg13g2_decap_4 FILLER_45_486 ();
 sg13g2_fill_1 FILLER_45_490 ();
 sg13g2_fill_2 FILLER_45_501 ();
 sg13g2_fill_1 FILLER_45_503 ();
 sg13g2_fill_1 FILLER_45_591 ();
 sg13g2_fill_2 FILLER_45_618 ();
 sg13g2_fill_2 FILLER_45_624 ();
 sg13g2_fill_2 FILLER_45_647 ();
 sg13g2_fill_1 FILLER_45_649 ();
 sg13g2_decap_8 FILLER_45_680 ();
 sg13g2_decap_8 FILLER_45_687 ();
 sg13g2_fill_2 FILLER_45_694 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_fill_2 FILLER_45_746 ();
 sg13g2_fill_1 FILLER_45_748 ();
 sg13g2_fill_1 FILLER_45_760 ();
 sg13g2_fill_2 FILLER_45_814 ();
 sg13g2_fill_2 FILLER_45_868 ();
 sg13g2_decap_4 FILLER_45_874 ();
 sg13g2_decap_4 FILLER_45_914 ();
 sg13g2_fill_2 FILLER_45_926 ();
 sg13g2_decap_4 FILLER_45_944 ();
 sg13g2_fill_1 FILLER_45_948 ();
 sg13g2_decap_8 FILLER_45_963 ();
 sg13g2_decap_4 FILLER_45_970 ();
 sg13g2_fill_2 FILLER_45_974 ();
 sg13g2_fill_1 FILLER_45_981 ();
 sg13g2_fill_2 FILLER_45_1006 ();
 sg13g2_fill_1 FILLER_45_1008 ();
 sg13g2_fill_2 FILLER_45_1035 ();
 sg13g2_decap_8 FILLER_45_1073 ();
 sg13g2_decap_8 FILLER_45_1080 ();
 sg13g2_decap_4 FILLER_45_1087 ();
 sg13g2_decap_8 FILLER_45_1112 ();
 sg13g2_decap_4 FILLER_45_1119 ();
 sg13g2_fill_2 FILLER_45_1133 ();
 sg13g2_decap_8 FILLER_45_1187 ();
 sg13g2_decap_8 FILLER_45_1194 ();
 sg13g2_fill_2 FILLER_45_1201 ();
 sg13g2_decap_8 FILLER_45_1213 ();
 sg13g2_fill_2 FILLER_45_1220 ();
 sg13g2_fill_1 FILLER_45_1272 ();
 sg13g2_fill_2 FILLER_45_1299 ();
 sg13g2_decap_4 FILLER_45_1311 ();
 sg13g2_fill_1 FILLER_45_1325 ();
 sg13g2_fill_2 FILLER_45_1352 ();
 sg13g2_fill_2 FILLER_45_1362 ();
 sg13g2_fill_1 FILLER_45_1364 ();
 sg13g2_fill_2 FILLER_45_1411 ();
 sg13g2_fill_1 FILLER_45_1413 ();
 sg13g2_fill_2 FILLER_45_1424 ();
 sg13g2_fill_1 FILLER_45_1426 ();
 sg13g2_fill_2 FILLER_45_1431 ();
 sg13g2_fill_1 FILLER_45_1433 ();
 sg13g2_decap_8 FILLER_45_1474 ();
 sg13g2_decap_8 FILLER_45_1481 ();
 sg13g2_decap_8 FILLER_45_1488 ();
 sg13g2_fill_2 FILLER_45_1495 ();
 sg13g2_fill_1 FILLER_45_1497 ();
 sg13g2_decap_4 FILLER_45_1516 ();
 sg13g2_decap_8 FILLER_45_1566 ();
 sg13g2_fill_1 FILLER_45_1573 ();
 sg13g2_fill_1 FILLER_45_1586 ();
 sg13g2_decap_4 FILLER_45_1631 ();
 sg13g2_decap_8 FILLER_45_1643 ();
 sg13g2_decap_8 FILLER_45_1650 ();
 sg13g2_decap_4 FILLER_45_1657 ();
 sg13g2_fill_2 FILLER_45_1661 ();
 sg13g2_decap_8 FILLER_45_1667 ();
 sg13g2_decap_8 FILLER_45_1674 ();
 sg13g2_decap_4 FILLER_45_1681 ();
 sg13g2_fill_2 FILLER_45_1685 ();
 sg13g2_decap_8 FILLER_45_1713 ();
 sg13g2_fill_2 FILLER_45_1720 ();
 sg13g2_fill_1 FILLER_45_1722 ();
 sg13g2_decap_8 FILLER_45_1741 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_18 ();
 sg13g2_fill_1 FILLER_46_20 ();
 sg13g2_fill_1 FILLER_46_25 ();
 sg13g2_decap_8 FILLER_46_30 ();
 sg13g2_decap_8 FILLER_46_37 ();
 sg13g2_fill_2 FILLER_46_44 ();
 sg13g2_decap_8 FILLER_46_53 ();
 sg13g2_decap_8 FILLER_46_60 ();
 sg13g2_decap_8 FILLER_46_67 ();
 sg13g2_decap_8 FILLER_46_74 ();
 sg13g2_decap_4 FILLER_46_81 ();
 sg13g2_fill_2 FILLER_46_85 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_fill_1 FILLER_46_154 ();
 sg13g2_decap_4 FILLER_46_181 ();
 sg13g2_decap_8 FILLER_46_223 ();
 sg13g2_fill_1 FILLER_46_230 ();
 sg13g2_decap_4 FILLER_46_291 ();
 sg13g2_fill_1 FILLER_46_295 ();
 sg13g2_decap_8 FILLER_46_299 ();
 sg13g2_decap_4 FILLER_46_306 ();
 sg13g2_decap_4 FILLER_46_369 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_4 FILLER_46_413 ();
 sg13g2_decap_4 FILLER_46_427 ();
 sg13g2_decap_4 FILLER_46_444 ();
 sg13g2_fill_2 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_505 ();
 sg13g2_fill_2 FILLER_46_512 ();
 sg13g2_fill_1 FILLER_46_514 ();
 sg13g2_fill_2 FILLER_46_541 ();
 sg13g2_fill_2 FILLER_46_553 ();
 sg13g2_fill_1 FILLER_46_555 ();
 sg13g2_fill_2 FILLER_46_566 ();
 sg13g2_fill_1 FILLER_46_568 ();
 sg13g2_fill_2 FILLER_46_595 ();
 sg13g2_fill_2 FILLER_46_678 ();
 sg13g2_fill_1 FILLER_46_695 ();
 sg13g2_fill_2 FILLER_46_706 ();
 sg13g2_decap_8 FILLER_46_734 ();
 sg13g2_decap_8 FILLER_46_741 ();
 sg13g2_decap_4 FILLER_46_748 ();
 sg13g2_fill_2 FILLER_46_752 ();
 sg13g2_decap_8 FILLER_46_758 ();
 sg13g2_fill_2 FILLER_46_765 ();
 sg13g2_fill_1 FILLER_46_767 ();
 sg13g2_decap_8 FILLER_46_778 ();
 sg13g2_decap_8 FILLER_46_789 ();
 sg13g2_decap_8 FILLER_46_796 ();
 sg13g2_decap_8 FILLER_46_803 ();
 sg13g2_fill_1 FILLER_46_810 ();
 sg13g2_fill_1 FILLER_46_815 ();
 sg13g2_fill_1 FILLER_46_842 ();
 sg13g2_fill_2 FILLER_46_847 ();
 sg13g2_fill_2 FILLER_46_859 ();
 sg13g2_fill_1 FILLER_46_917 ();
 sg13g2_fill_1 FILLER_46_926 ();
 sg13g2_fill_2 FILLER_46_944 ();
 sg13g2_fill_1 FILLER_46_946 ();
 sg13g2_decap_4 FILLER_46_955 ();
 sg13g2_decap_8 FILLER_46_963 ();
 sg13g2_fill_1 FILLER_46_970 ();
 sg13g2_decap_4 FILLER_46_981 ();
 sg13g2_fill_1 FILLER_46_985 ();
 sg13g2_fill_1 FILLER_46_994 ();
 sg13g2_fill_2 FILLER_46_1005 ();
 sg13g2_fill_1 FILLER_46_1017 ();
 sg13g2_fill_2 FILLER_46_1022 ();
 sg13g2_decap_4 FILLER_46_1028 ();
 sg13g2_fill_2 FILLER_46_1032 ();
 sg13g2_decap_4 FILLER_46_1038 ();
 sg13g2_fill_1 FILLER_46_1042 ();
 sg13g2_fill_2 FILLER_46_1053 ();
 sg13g2_fill_1 FILLER_46_1055 ();
 sg13g2_fill_2 FILLER_46_1082 ();
 sg13g2_decap_4 FILLER_46_1114 ();
 sg13g2_fill_2 FILLER_46_1118 ();
 sg13g2_decap_8 FILLER_46_1145 ();
 sg13g2_decap_8 FILLER_46_1152 ();
 sg13g2_fill_2 FILLER_46_1159 ();
 sg13g2_fill_1 FILLER_46_1161 ();
 sg13g2_fill_1 FILLER_46_1166 ();
 sg13g2_decap_8 FILLER_46_1200 ();
 sg13g2_decap_8 FILLER_46_1207 ();
 sg13g2_decap_4 FILLER_46_1214 ();
 sg13g2_fill_2 FILLER_46_1218 ();
 sg13g2_decap_8 FILLER_46_1246 ();
 sg13g2_fill_1 FILLER_46_1274 ();
 sg13g2_decap_8 FILLER_46_1345 ();
 sg13g2_decap_8 FILLER_46_1352 ();
 sg13g2_decap_4 FILLER_46_1402 ();
 sg13g2_fill_1 FILLER_46_1406 ();
 sg13g2_decap_8 FILLER_46_1417 ();
 sg13g2_fill_1 FILLER_46_1428 ();
 sg13g2_fill_2 FILLER_46_1450 ();
 sg13g2_decap_8 FILLER_46_1466 ();
 sg13g2_decap_8 FILLER_46_1473 ();
 sg13g2_decap_8 FILLER_46_1480 ();
 sg13g2_decap_8 FILLER_46_1487 ();
 sg13g2_fill_1 FILLER_46_1494 ();
 sg13g2_decap_4 FILLER_46_1521 ();
 sg13g2_fill_2 FILLER_46_1525 ();
 sg13g2_fill_2 FILLER_46_1535 ();
 sg13g2_decap_4 FILLER_46_1541 ();
 sg13g2_fill_2 FILLER_46_1549 ();
 sg13g2_decap_8 FILLER_46_1616 ();
 sg13g2_decap_8 FILLER_46_1623 ();
 sg13g2_fill_2 FILLER_46_1630 ();
 sg13g2_fill_1 FILLER_46_1632 ();
 sg13g2_decap_8 FILLER_46_1669 ();
 sg13g2_fill_1 FILLER_46_1676 ();
 sg13g2_decap_8 FILLER_46_1713 ();
 sg13g2_decap_4 FILLER_46_1720 ();
 sg13g2_fill_2 FILLER_46_1734 ();
 sg13g2_decap_8 FILLER_46_1762 ();
 sg13g2_decap_4 FILLER_46_1769 ();
 sg13g2_fill_1 FILLER_46_1773 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_11 ();
 sg13g2_decap_8 FILLER_47_39 ();
 sg13g2_decap_8 FILLER_47_46 ();
 sg13g2_decap_8 FILLER_47_53 ();
 sg13g2_decap_8 FILLER_47_60 ();
 sg13g2_fill_1 FILLER_47_67 ();
 sg13g2_decap_8 FILLER_47_72 ();
 sg13g2_decap_8 FILLER_47_79 ();
 sg13g2_decap_8 FILLER_47_86 ();
 sg13g2_decap_8 FILLER_47_93 ();
 sg13g2_decap_8 FILLER_47_100 ();
 sg13g2_decap_8 FILLER_47_107 ();
 sg13g2_decap_8 FILLER_47_114 ();
 sg13g2_decap_8 FILLER_47_121 ();
 sg13g2_decap_8 FILLER_47_128 ();
 sg13g2_decap_8 FILLER_47_135 ();
 sg13g2_decap_4 FILLER_47_142 ();
 sg13g2_fill_1 FILLER_47_146 ();
 sg13g2_decap_4 FILLER_47_155 ();
 sg13g2_fill_2 FILLER_47_159 ();
 sg13g2_decap_4 FILLER_47_165 ();
 sg13g2_fill_1 FILLER_47_169 ();
 sg13g2_fill_2 FILLER_47_192 ();
 sg13g2_fill_1 FILLER_47_198 ();
 sg13g2_decap_8 FILLER_47_229 ();
 sg13g2_decap_8 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_243 ();
 sg13g2_decap_4 FILLER_47_254 ();
 sg13g2_fill_1 FILLER_47_263 ();
 sg13g2_fill_2 FILLER_47_274 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_fill_1 FILLER_47_282 ();
 sg13g2_fill_2 FILLER_47_293 ();
 sg13g2_fill_1 FILLER_47_295 ();
 sg13g2_decap_4 FILLER_47_368 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_decap_4 FILLER_47_387 ();
 sg13g2_fill_1 FILLER_47_391 ();
 sg13g2_fill_1 FILLER_47_446 ();
 sg13g2_fill_2 FILLER_47_462 ();
 sg13g2_fill_1 FILLER_47_464 ();
 sg13g2_fill_2 FILLER_47_491 ();
 sg13g2_fill_2 FILLER_47_496 ();
 sg13g2_fill_1 FILLER_47_498 ();
 sg13g2_fill_2 FILLER_47_507 ();
 sg13g2_fill_1 FILLER_47_509 ();
 sg13g2_decap_8 FILLER_47_534 ();
 sg13g2_fill_1 FILLER_47_541 ();
 sg13g2_fill_2 FILLER_47_552 ();
 sg13g2_fill_2 FILLER_47_580 ();
 sg13g2_decap_4 FILLER_47_586 ();
 sg13g2_decap_4 FILLER_47_598 ();
 sg13g2_fill_2 FILLER_47_612 ();
 sg13g2_fill_1 FILLER_47_624 ();
 sg13g2_fill_2 FILLER_47_629 ();
 sg13g2_fill_1 FILLER_47_631 ();
 sg13g2_fill_2 FILLER_47_658 ();
 sg13g2_fill_1 FILLER_47_660 ();
 sg13g2_fill_1 FILLER_47_681 ();
 sg13g2_fill_2 FILLER_47_710 ();
 sg13g2_fill_2 FILLER_47_716 ();
 sg13g2_fill_1 FILLER_47_718 ();
 sg13g2_decap_8 FILLER_47_723 ();
 sg13g2_decap_8 FILLER_47_730 ();
 sg13g2_decap_8 FILLER_47_737 ();
 sg13g2_fill_2 FILLER_47_757 ();
 sg13g2_fill_2 FILLER_47_785 ();
 sg13g2_decap_8 FILLER_47_842 ();
 sg13g2_fill_2 FILLER_47_857 ();
 sg13g2_fill_1 FILLER_47_859 ();
 sg13g2_fill_2 FILLER_47_886 ();
 sg13g2_decap_4 FILLER_47_902 ();
 sg13g2_decap_4 FILLER_47_916 ();
 sg13g2_fill_1 FILLER_47_920 ();
 sg13g2_fill_2 FILLER_47_924 ();
 sg13g2_fill_1 FILLER_47_926 ();
 sg13g2_decap_4 FILLER_47_935 ();
 sg13g2_decap_8 FILLER_47_942 ();
 sg13g2_fill_1 FILLER_47_949 ();
 sg13g2_decap_8 FILLER_47_992 ();
 sg13g2_decap_8 FILLER_47_999 ();
 sg13g2_decap_8 FILLER_47_1006 ();
 sg13g2_decap_8 FILLER_47_1013 ();
 sg13g2_fill_2 FILLER_47_1020 ();
 sg13g2_fill_1 FILLER_47_1022 ();
 sg13g2_decap_8 FILLER_47_1028 ();
 sg13g2_fill_1 FILLER_47_1035 ();
 sg13g2_decap_4 FILLER_47_1040 ();
 sg13g2_decap_4 FILLER_47_1058 ();
 sg13g2_fill_2 FILLER_47_1062 ();
 sg13g2_decap_8 FILLER_47_1068 ();
 sg13g2_decap_4 FILLER_47_1075 ();
 sg13g2_fill_2 FILLER_47_1079 ();
 sg13g2_decap_8 FILLER_47_1091 ();
 sg13g2_fill_1 FILLER_47_1098 ();
 sg13g2_fill_2 FILLER_47_1135 ();
 sg13g2_fill_1 FILLER_47_1137 ();
 sg13g2_decap_4 FILLER_47_1159 ();
 sg13g2_fill_1 FILLER_47_1163 ();
 sg13g2_fill_1 FILLER_47_1193 ();
 sg13g2_decap_4 FILLER_47_1218 ();
 sg13g2_fill_2 FILLER_47_1252 ();
 sg13g2_fill_2 FILLER_47_1280 ();
 sg13g2_decap_4 FILLER_47_1286 ();
 sg13g2_fill_2 FILLER_47_1290 ();
 sg13g2_decap_8 FILLER_47_1296 ();
 sg13g2_fill_1 FILLER_47_1303 ();
 sg13g2_decap_8 FILLER_47_1328 ();
 sg13g2_decap_8 FILLER_47_1335 ();
 sg13g2_decap_8 FILLER_47_1342 ();
 sg13g2_decap_8 FILLER_47_1349 ();
 sg13g2_decap_4 FILLER_47_1356 ();
 sg13g2_fill_1 FILLER_47_1360 ();
 sg13g2_fill_2 FILLER_47_1371 ();
 sg13g2_decap_4 FILLER_47_1404 ();
 sg13g2_fill_2 FILLER_47_1418 ();
 sg13g2_fill_1 FILLER_47_1420 ();
 sg13g2_decap_8 FILLER_47_1473 ();
 sg13g2_decap_8 FILLER_47_1524 ();
 sg13g2_decap_8 FILLER_47_1571 ();
 sg13g2_decap_8 FILLER_47_1578 ();
 sg13g2_fill_2 FILLER_47_1585 ();
 sg13g2_fill_1 FILLER_47_1587 ();
 sg13g2_decap_8 FILLER_47_1628 ();
 sg13g2_decap_8 FILLER_47_1635 ();
 sg13g2_decap_8 FILLER_47_1642 ();
 sg13g2_fill_2 FILLER_47_1649 ();
 sg13g2_decap_8 FILLER_47_1655 ();
 sg13g2_fill_2 FILLER_47_1662 ();
 sg13g2_fill_1 FILLER_47_1664 ();
 sg13g2_decap_8 FILLER_47_1675 ();
 sg13g2_fill_2 FILLER_47_1682 ();
 sg13g2_fill_1 FILLER_47_1684 ();
 sg13g2_decap_8 FILLER_47_1703 ();
 sg13g2_fill_2 FILLER_47_1745 ();
 sg13g2_fill_1 FILLER_47_1747 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_48_7 ();
 sg13g2_fill_2 FILLER_48_11 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_56 ();
 sg13g2_fill_1 FILLER_48_58 ();
 sg13g2_fill_1 FILLER_48_115 ();
 sg13g2_fill_1 FILLER_48_142 ();
 sg13g2_decap_4 FILLER_48_153 ();
 sg13g2_fill_1 FILLER_48_157 ();
 sg13g2_fill_2 FILLER_48_174 ();
 sg13g2_fill_2 FILLER_48_185 ();
 sg13g2_decap_8 FILLER_48_228 ();
 sg13g2_decap_8 FILLER_48_235 ();
 sg13g2_decap_8 FILLER_48_242 ();
 sg13g2_decap_8 FILLER_48_249 ();
 sg13g2_decap_4 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_270 ();
 sg13g2_fill_2 FILLER_48_297 ();
 sg13g2_fill_2 FILLER_48_303 ();
 sg13g2_fill_2 FILLER_48_310 ();
 sg13g2_fill_2 FILLER_48_358 ();
 sg13g2_fill_1 FILLER_48_360 ();
 sg13g2_fill_1 FILLER_48_414 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_fill_2 FILLER_48_455 ();
 sg13g2_fill_1 FILLER_48_457 ();
 sg13g2_fill_2 FILLER_48_472 ();
 sg13g2_fill_2 FILLER_48_482 ();
 sg13g2_fill_2 FILLER_48_498 ();
 sg13g2_fill_1 FILLER_48_500 ();
 sg13g2_decap_8 FILLER_48_506 ();
 sg13g2_decap_8 FILLER_48_513 ();
 sg13g2_fill_1 FILLER_48_520 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_fill_2 FILLER_48_546 ();
 sg13g2_fill_1 FILLER_48_548 ();
 sg13g2_decap_4 FILLER_48_588 ();
 sg13g2_fill_2 FILLER_48_592 ();
 sg13g2_decap_4 FILLER_48_598 ();
 sg13g2_fill_1 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_643 ();
 sg13g2_decap_8 FILLER_48_650 ();
 sg13g2_fill_2 FILLER_48_675 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_739 ();
 sg13g2_decap_4 FILLER_48_746 ();
 sg13g2_fill_1 FILLER_48_750 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_fill_2 FILLER_48_798 ();
 sg13g2_decap_4 FILLER_48_804 ();
 sg13g2_fill_2 FILLER_48_808 ();
 sg13g2_fill_2 FILLER_48_856 ();
 sg13g2_fill_2 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_880 ();
 sg13g2_fill_1 FILLER_48_887 ();
 sg13g2_decap_4 FILLER_48_914 ();
 sg13g2_fill_1 FILLER_48_918 ();
 sg13g2_decap_8 FILLER_48_924 ();
 sg13g2_decap_4 FILLER_48_931 ();
 sg13g2_decap_4 FILLER_48_949 ();
 sg13g2_decap_8 FILLER_48_1005 ();
 sg13g2_decap_8 FILLER_48_1012 ();
 sg13g2_decap_8 FILLER_48_1019 ();
 sg13g2_fill_1 FILLER_48_1026 ();
 sg13g2_fill_2 FILLER_48_1079 ();
 sg13g2_fill_1 FILLER_48_1081 ();
 sg13g2_fill_1 FILLER_48_1092 ();
 sg13g2_fill_2 FILLER_48_1128 ();
 sg13g2_fill_1 FILLER_48_1130 ();
 sg13g2_decap_4 FILLER_48_1157 ();
 sg13g2_fill_2 FILLER_48_1161 ();
 sg13g2_decap_4 FILLER_48_1187 ();
 sg13g2_decap_8 FILLER_48_1201 ();
 sg13g2_fill_2 FILLER_48_1208 ();
 sg13g2_fill_1 FILLER_48_1240 ();
 sg13g2_decap_8 FILLER_48_1278 ();
 sg13g2_decap_4 FILLER_48_1285 ();
 sg13g2_fill_2 FILLER_48_1289 ();
 sg13g2_decap_8 FILLER_48_1346 ();
 sg13g2_fill_2 FILLER_48_1387 ();
 sg13g2_fill_1 FILLER_48_1389 ();
 sg13g2_fill_2 FILLER_48_1452 ();
 sg13g2_fill_1 FILLER_48_1454 ();
 sg13g2_decap_8 FILLER_48_1459 ();
 sg13g2_fill_2 FILLER_48_1466 ();
 sg13g2_fill_1 FILLER_48_1468 ();
 sg13g2_fill_1 FILLER_48_1482 ();
 sg13g2_decap_8 FILLER_48_1513 ();
 sg13g2_decap_8 FILLER_48_1520 ();
 sg13g2_fill_2 FILLER_48_1527 ();
 sg13g2_fill_1 FILLER_48_1529 ();
 sg13g2_fill_2 FILLER_48_1587 ();
 sg13g2_fill_2 FILLER_48_1645 ();
 sg13g2_fill_1 FILLER_48_1647 ();
 sg13g2_fill_1 FILLER_48_1674 ();
 sg13g2_fill_2 FILLER_48_1679 ();
 sg13g2_decap_4 FILLER_48_1686 ();
 sg13g2_fill_1 FILLER_48_1690 ();
 sg13g2_decap_4 FILLER_48_1717 ();
 sg13g2_fill_1 FILLER_48_1721 ();
 sg13g2_decap_8 FILLER_48_1762 ();
 sg13g2_decap_4 FILLER_48_1769 ();
 sg13g2_fill_1 FILLER_48_1773 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_92 ();
 sg13g2_decap_8 FILLER_49_99 ();
 sg13g2_fill_2 FILLER_49_106 ();
 sg13g2_fill_1 FILLER_49_108 ();
 sg13g2_fill_2 FILLER_49_119 ();
 sg13g2_fill_2 FILLER_49_147 ();
 sg13g2_decap_4 FILLER_49_185 ();
 sg13g2_fill_2 FILLER_49_189 ();
 sg13g2_fill_2 FILLER_49_201 ();
 sg13g2_fill_2 FILLER_49_229 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_4 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_283 ();
 sg13g2_decap_8 FILLER_49_290 ();
 sg13g2_decap_8 FILLER_49_297 ();
 sg13g2_fill_2 FILLER_49_304 ();
 sg13g2_decap_8 FILLER_49_316 ();
 sg13g2_fill_2 FILLER_49_323 ();
 sg13g2_decap_4 FILLER_49_335 ();
 sg13g2_fill_2 FILLER_49_343 ();
 sg13g2_fill_2 FILLER_49_357 ();
 sg13g2_fill_1 FILLER_49_398 ();
 sg13g2_fill_1 FILLER_49_410 ();
 sg13g2_fill_2 FILLER_49_421 ();
 sg13g2_decap_4 FILLER_49_452 ();
 sg13g2_fill_2 FILLER_49_456 ();
 sg13g2_decap_4 FILLER_49_499 ();
 sg13g2_fill_1 FILLER_49_503 ();
 sg13g2_decap_4 FILLER_49_513 ();
 sg13g2_fill_2 FILLER_49_517 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_540 ();
 sg13g2_decap_8 FILLER_49_547 ();
 sg13g2_fill_1 FILLER_49_554 ();
 sg13g2_fill_2 FILLER_49_581 ();
 sg13g2_fill_2 FILLER_49_596 ();
 sg13g2_decap_8 FILLER_49_628 ();
 sg13g2_decap_8 FILLER_49_635 ();
 sg13g2_decap_8 FILLER_49_642 ();
 sg13g2_decap_4 FILLER_49_649 ();
 sg13g2_fill_2 FILLER_49_653 ();
 sg13g2_fill_2 FILLER_49_708 ();
 sg13g2_fill_2 FILLER_49_720 ();
 sg13g2_decap_8 FILLER_49_727 ();
 sg13g2_decap_8 FILLER_49_734 ();
 sg13g2_decap_8 FILLER_49_741 ();
 sg13g2_decap_4 FILLER_49_758 ();
 sg13g2_fill_1 FILLER_49_762 ();
 sg13g2_decap_8 FILLER_49_767 ();
 sg13g2_decap_8 FILLER_49_774 ();
 sg13g2_decap_8 FILLER_49_781 ();
 sg13g2_decap_4 FILLER_49_788 ();
 sg13g2_fill_1 FILLER_49_792 ();
 sg13g2_fill_1 FILLER_49_797 ();
 sg13g2_fill_1 FILLER_49_824 ();
 sg13g2_fill_1 FILLER_49_835 ();
 sg13g2_fill_2 FILLER_49_862 ();
 sg13g2_fill_1 FILLER_49_868 ();
 sg13g2_fill_2 FILLER_49_879 ();
 sg13g2_fill_2 FILLER_49_891 ();
 sg13g2_fill_2 FILLER_49_897 ();
 sg13g2_fill_1 FILLER_49_899 ();
 sg13g2_fill_1 FILLER_49_904 ();
 sg13g2_decap_4 FILLER_49_975 ();
 sg13g2_decap_8 FILLER_49_1013 ();
 sg13g2_fill_1 FILLER_49_1020 ();
 sg13g2_fill_2 FILLER_49_1051 ();
 sg13g2_fill_1 FILLER_49_1053 ();
 sg13g2_decap_8 FILLER_49_1084 ();
 sg13g2_decap_8 FILLER_49_1091 ();
 sg13g2_fill_2 FILLER_49_1098 ();
 sg13g2_fill_1 FILLER_49_1100 ();
 sg13g2_decap_8 FILLER_49_1105 ();
 sg13g2_decap_8 FILLER_49_1112 ();
 sg13g2_decap_4 FILLER_49_1119 ();
 sg13g2_fill_2 FILLER_49_1123 ();
 sg13g2_decap_8 FILLER_49_1139 ();
 sg13g2_decap_8 FILLER_49_1146 ();
 sg13g2_decap_8 FILLER_49_1153 ();
 sg13g2_decap_8 FILLER_49_1160 ();
 sg13g2_decap_4 FILLER_49_1167 ();
 sg13g2_fill_1 FILLER_49_1171 ();
 sg13g2_fill_2 FILLER_49_1236 ();
 sg13g2_fill_1 FILLER_49_1238 ();
 sg13g2_decap_4 FILLER_49_1274 ();
 sg13g2_decap_8 FILLER_49_1288 ();
 sg13g2_fill_1 FILLER_49_1295 ();
 sg13g2_decap_8 FILLER_49_1348 ();
 sg13g2_fill_2 FILLER_49_1368 ();
 sg13g2_fill_1 FILLER_49_1396 ();
 sg13g2_fill_1 FILLER_49_1401 ();
 sg13g2_decap_4 FILLER_49_1437 ();
 sg13g2_fill_2 FILLER_49_1441 ();
 sg13g2_decap_8 FILLER_49_1447 ();
 sg13g2_decap_8 FILLER_49_1454 ();
 sg13g2_fill_2 FILLER_49_1461 ();
 sg13g2_fill_1 FILLER_49_1463 ();
 sg13g2_decap_8 FILLER_49_1510 ();
 sg13g2_decap_8 FILLER_49_1517 ();
 sg13g2_fill_1 FILLER_49_1524 ();
 sg13g2_fill_1 FILLER_49_1537 ();
 sg13g2_decap_4 FILLER_49_1551 ();
 sg13g2_fill_1 FILLER_49_1585 ();
 sg13g2_decap_8 FILLER_49_1596 ();
 sg13g2_decap_8 FILLER_49_1603 ();
 sg13g2_fill_2 FILLER_49_1610 ();
 sg13g2_fill_1 FILLER_49_1612 ();
 sg13g2_decap_4 FILLER_49_1623 ();
 sg13g2_fill_1 FILLER_49_1627 ();
 sg13g2_decap_8 FILLER_49_1632 ();
 sg13g2_decap_4 FILLER_49_1639 ();
 sg13g2_decap_4 FILLER_49_1653 ();
 sg13g2_decap_8 FILLER_49_1661 ();
 sg13g2_fill_2 FILLER_49_1668 ();
 sg13g2_fill_1 FILLER_49_1670 ();
 sg13g2_decap_8 FILLER_49_1701 ();
 sg13g2_decap_8 FILLER_49_1708 ();
 sg13g2_decap_4 FILLER_49_1715 ();
 sg13g2_fill_2 FILLER_49_1719 ();
 sg13g2_fill_1 FILLER_49_1735 ();
 sg13g2_decap_8 FILLER_49_1766 ();
 sg13g2_fill_1 FILLER_49_1773 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_5 ();
 sg13g2_fill_1 FILLER_50_10 ();
 sg13g2_fill_2 FILLER_50_41 ();
 sg13g2_decap_4 FILLER_50_62 ();
 sg13g2_fill_2 FILLER_50_66 ();
 sg13g2_decap_4 FILLER_50_98 ();
 sg13g2_fill_2 FILLER_50_150 ();
 sg13g2_fill_1 FILLER_50_152 ();
 sg13g2_fill_2 FILLER_50_193 ();
 sg13g2_fill_1 FILLER_50_195 ();
 sg13g2_fill_2 FILLER_50_226 ();
 sg13g2_decap_8 FILLER_50_232 ();
 sg13g2_decap_8 FILLER_50_239 ();
 sg13g2_decap_8 FILLER_50_246 ();
 sg13g2_fill_2 FILLER_50_253 ();
 sg13g2_decap_8 FILLER_50_281 ();
 sg13g2_decap_8 FILLER_50_288 ();
 sg13g2_fill_2 FILLER_50_305 ();
 sg13g2_decap_8 FILLER_50_333 ();
 sg13g2_decap_8 FILLER_50_376 ();
 sg13g2_decap_8 FILLER_50_383 ();
 sg13g2_fill_1 FILLER_50_390 ();
 sg13g2_fill_2 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_50_458 ();
 sg13g2_decap_8 FILLER_50_465 ();
 sg13g2_decap_4 FILLER_50_472 ();
 sg13g2_decap_4 FILLER_50_489 ();
 sg13g2_fill_1 FILLER_50_493 ();
 sg13g2_decap_4 FILLER_50_497 ();
 sg13g2_fill_1 FILLER_50_501 ();
 sg13g2_decap_8 FILLER_50_554 ();
 sg13g2_fill_1 FILLER_50_561 ();
 sg13g2_decap_8 FILLER_50_566 ();
 sg13g2_decap_4 FILLER_50_573 ();
 sg13g2_fill_1 FILLER_50_582 ();
 sg13g2_decap_8 FILLER_50_589 ();
 sg13g2_decap_8 FILLER_50_596 ();
 sg13g2_fill_1 FILLER_50_603 ();
 sg13g2_decap_8 FILLER_50_630 ();
 sg13g2_fill_1 FILLER_50_637 ();
 sg13g2_fill_1 FILLER_50_698 ();
 sg13g2_decap_4 FILLER_50_712 ();
 sg13g2_fill_2 FILLER_50_716 ();
 sg13g2_decap_8 FILLER_50_761 ();
 sg13g2_fill_1 FILLER_50_778 ();
 sg13g2_fill_2 FILLER_50_789 ();
 sg13g2_decap_4 FILLER_50_817 ();
 sg13g2_fill_2 FILLER_50_844 ();
 sg13g2_fill_1 FILLER_50_854 ();
 sg13g2_fill_2 FILLER_50_886 ();
 sg13g2_fill_1 FILLER_50_888 ();
 sg13g2_fill_1 FILLER_50_925 ();
 sg13g2_fill_1 FILLER_50_930 ();
 sg13g2_fill_1 FILLER_50_957 ();
 sg13g2_fill_1 FILLER_50_985 ();
 sg13g2_fill_1 FILLER_50_1012 ();
 sg13g2_decap_8 FILLER_50_1021 ();
 sg13g2_fill_1 FILLER_50_1028 ();
 sg13g2_fill_2 FILLER_50_1043 ();
 sg13g2_decap_8 FILLER_50_1055 ();
 sg13g2_decap_4 FILLER_50_1062 ();
 sg13g2_fill_1 FILLER_50_1066 ();
 sg13g2_decap_8 FILLER_50_1071 ();
 sg13g2_fill_2 FILLER_50_1078 ();
 sg13g2_fill_1 FILLER_50_1090 ();
 sg13g2_decap_8 FILLER_50_1117 ();
 sg13g2_decap_8 FILLER_50_1124 ();
 sg13g2_fill_2 FILLER_50_1131 ();
 sg13g2_fill_1 FILLER_50_1133 ();
 sg13g2_decap_4 FILLER_50_1138 ();
 sg13g2_fill_2 FILLER_50_1142 ();
 sg13g2_decap_8 FILLER_50_1174 ();
 sg13g2_decap_4 FILLER_50_1181 ();
 sg13g2_fill_1 FILLER_50_1185 ();
 sg13g2_decap_4 FILLER_50_1190 ();
 sg13g2_fill_1 FILLER_50_1194 ();
 sg13g2_fill_2 FILLER_50_1203 ();
 sg13g2_fill_1 FILLER_50_1241 ();
 sg13g2_fill_2 FILLER_50_1278 ();
 sg13g2_decap_8 FILLER_50_1310 ();
 sg13g2_fill_1 FILLER_50_1317 ();
 sg13g2_decap_4 FILLER_50_1344 ();
 sg13g2_decap_8 FILLER_50_1352 ();
 sg13g2_decap_8 FILLER_50_1359 ();
 sg13g2_decap_8 FILLER_50_1366 ();
 sg13g2_fill_1 FILLER_50_1373 ();
 sg13g2_decap_4 FILLER_50_1388 ();
 sg13g2_fill_1 FILLER_50_1392 ();
 sg13g2_fill_1 FILLER_50_1403 ();
 sg13g2_fill_2 FILLER_50_1430 ();
 sg13g2_fill_1 FILLER_50_1432 ();
 sg13g2_fill_1 FILLER_50_1469 ();
 sg13g2_fill_2 FILLER_50_1506 ();
 sg13g2_fill_1 FILLER_50_1508 ();
 sg13g2_decap_4 FILLER_50_1519 ();
 sg13g2_fill_2 FILLER_50_1523 ();
 sg13g2_fill_2 FILLER_50_1546 ();
 sg13g2_fill_2 FILLER_50_1569 ();
 sg13g2_fill_1 FILLER_50_1571 ();
 sg13g2_fill_1 FILLER_50_1582 ();
 sg13g2_fill_2 FILLER_50_1609 ();
 sg13g2_decap_8 FILLER_50_1662 ();
 sg13g2_decap_4 FILLER_50_1669 ();
 sg13g2_fill_2 FILLER_50_1683 ();
 sg13g2_decap_4 FILLER_50_1706 ();
 sg13g2_fill_2 FILLER_50_1710 ();
 sg13g2_decap_8 FILLER_50_1758 ();
 sg13g2_decap_8 FILLER_50_1765 ();
 sg13g2_fill_2 FILLER_50_1772 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_7 ();
 sg13g2_fill_1 FILLER_51_9 ();
 sg13g2_decap_8 FILLER_51_30 ();
 sg13g2_decap_8 FILLER_51_37 ();
 sg13g2_fill_2 FILLER_51_44 ();
 sg13g2_fill_1 FILLER_51_46 ();
 sg13g2_decap_8 FILLER_51_57 ();
 sg13g2_fill_2 FILLER_51_64 ();
 sg13g2_fill_2 FILLER_51_89 ();
 sg13g2_decap_4 FILLER_51_95 ();
 sg13g2_fill_2 FILLER_51_109 ();
 sg13g2_fill_1 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_120 ();
 sg13g2_fill_1 FILLER_51_122 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_fill_2 FILLER_51_154 ();
 sg13g2_fill_1 FILLER_51_156 ();
 sg13g2_fill_2 FILLER_51_187 ();
 sg13g2_fill_1 FILLER_51_189 ();
 sg13g2_decap_4 FILLER_51_217 ();
 sg13g2_decap_8 FILLER_51_247 ();
 sg13g2_decap_4 FILLER_51_254 ();
 sg13g2_fill_2 FILLER_51_258 ();
 sg13g2_fill_1 FILLER_51_268 ();
 sg13g2_fill_2 FILLER_51_279 ();
 sg13g2_fill_2 FILLER_51_285 ();
 sg13g2_fill_2 FILLER_51_313 ();
 sg13g2_fill_1 FILLER_51_325 ();
 sg13g2_fill_1 FILLER_51_374 ();
 sg13g2_decap_8 FILLER_51_415 ();
 sg13g2_fill_1 FILLER_51_422 ();
 sg13g2_fill_1 FILLER_51_433 ();
 sg13g2_decap_8 FILLER_51_442 ();
 sg13g2_decap_8 FILLER_51_485 ();
 sg13g2_fill_2 FILLER_51_502 ();
 sg13g2_fill_1 FILLER_51_504 ();
 sg13g2_decap_8 FILLER_51_545 ();
 sg13g2_decap_8 FILLER_51_552 ();
 sg13g2_decap_8 FILLER_51_559 ();
 sg13g2_decap_8 FILLER_51_566 ();
 sg13g2_fill_2 FILLER_51_573 ();
 sg13g2_decap_4 FILLER_51_625 ();
 sg13g2_fill_2 FILLER_51_629 ();
 sg13g2_fill_1 FILLER_51_641 ();
 sg13g2_fill_1 FILLER_51_668 ();
 sg13g2_fill_2 FILLER_51_719 ();
 sg13g2_decap_8 FILLER_51_725 ();
 sg13g2_decap_8 FILLER_51_732 ();
 sg13g2_fill_2 FILLER_51_739 ();
 sg13g2_fill_1 FILLER_51_741 ();
 sg13g2_fill_1 FILLER_51_804 ();
 sg13g2_fill_1 FILLER_51_809 ();
 sg13g2_fill_1 FILLER_51_820 ();
 sg13g2_decap_4 FILLER_51_837 ();
 sg13g2_fill_2 FILLER_51_841 ();
 sg13g2_decap_8 FILLER_51_847 ();
 sg13g2_decap_8 FILLER_51_854 ();
 sg13g2_decap_4 FILLER_51_861 ();
 sg13g2_fill_1 FILLER_51_865 ();
 sg13g2_decap_8 FILLER_51_870 ();
 sg13g2_decap_4 FILLER_51_877 ();
 sg13g2_fill_2 FILLER_51_881 ();
 sg13g2_fill_2 FILLER_51_886 ();
 sg13g2_fill_2 FILLER_51_924 ();
 sg13g2_fill_2 FILLER_51_930 ();
 sg13g2_fill_1 FILLER_51_932 ();
 sg13g2_fill_1 FILLER_51_937 ();
 sg13g2_decap_8 FILLER_51_948 ();
 sg13g2_decap_4 FILLER_51_975 ();
 sg13g2_fill_1 FILLER_51_979 ();
 sg13g2_decap_8 FILLER_51_1010 ();
 sg13g2_decap_8 FILLER_51_1017 ();
 sg13g2_fill_1 FILLER_51_1024 ();
 sg13g2_decap_8 FILLER_51_1059 ();
 sg13g2_fill_2 FILLER_51_1066 ();
 sg13g2_fill_1 FILLER_51_1068 ();
 sg13g2_fill_2 FILLER_51_1109 ();
 sg13g2_fill_1 FILLER_51_1121 ();
 sg13g2_fill_2 FILLER_51_1158 ();
 sg13g2_decap_8 FILLER_51_1186 ();
 sg13g2_decap_8 FILLER_51_1193 ();
 sg13g2_fill_1 FILLER_51_1200 ();
 sg13g2_decap_8 FILLER_51_1205 ();
 sg13g2_fill_2 FILLER_51_1248 ();
 sg13g2_fill_2 FILLER_51_1254 ();
 sg13g2_fill_1 FILLER_51_1256 ();
 sg13g2_fill_2 FILLER_51_1283 ();
 sg13g2_fill_1 FILLER_51_1285 ();
 sg13g2_fill_2 FILLER_51_1290 ();
 sg13g2_fill_2 FILLER_51_1338 ();
 sg13g2_fill_1 FILLER_51_1366 ();
 sg13g2_decap_8 FILLER_51_1403 ();
 sg13g2_fill_2 FILLER_51_1410 ();
 sg13g2_fill_1 FILLER_51_1412 ();
 sg13g2_fill_1 FILLER_51_1417 ();
 sg13g2_decap_8 FILLER_51_1484 ();
 sg13g2_decap_8 FILLER_51_1491 ();
 sg13g2_decap_4 FILLER_51_1508 ();
 sg13g2_fill_2 FILLER_51_1512 ();
 sg13g2_fill_2 FILLER_51_1540 ();
 sg13g2_decap_4 FILLER_51_1572 ();
 sg13g2_decap_4 FILLER_51_1612 ();
 sg13g2_fill_2 FILLER_51_1616 ();
 sg13g2_decap_4 FILLER_51_1622 ();
 sg13g2_fill_1 FILLER_51_1626 ();
 sg13g2_fill_2 FILLER_51_1663 ();
 sg13g2_fill_1 FILLER_51_1665 ();
 sg13g2_decap_8 FILLER_51_1706 ();
 sg13g2_decap_4 FILLER_51_1713 ();
 sg13g2_fill_1 FILLER_51_1717 ();
 sg13g2_decap_8 FILLER_51_1758 ();
 sg13g2_decap_8 FILLER_51_1765 ();
 sg13g2_fill_2 FILLER_51_1772 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_11 ();
 sg13g2_fill_1 FILLER_52_20 ();
 sg13g2_fill_1 FILLER_52_47 ();
 sg13g2_fill_1 FILLER_52_58 ();
 sg13g2_fill_2 FILLER_52_95 ();
 sg13g2_decap_8 FILLER_52_107 ();
 sg13g2_decap_4 FILLER_52_114 ();
 sg13g2_fill_1 FILLER_52_154 ();
 sg13g2_decap_4 FILLER_52_169 ();
 sg13g2_fill_1 FILLER_52_173 ();
 sg13g2_decap_4 FILLER_52_263 ();
 sg13g2_decap_8 FILLER_52_277 ();
 sg13g2_fill_1 FILLER_52_284 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_decap_4 FILLER_52_317 ();
 sg13g2_decap_8 FILLER_52_329 ();
 sg13g2_fill_2 FILLER_52_336 ();
 sg13g2_decap_4 FILLER_52_342 ();
 sg13g2_decap_8 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_4 FILLER_52_364 ();
 sg13g2_fill_2 FILLER_52_368 ();
 sg13g2_fill_2 FILLER_52_383 ();
 sg13g2_fill_2 FILLER_52_389 ();
 sg13g2_decap_8 FILLER_52_425 ();
 sg13g2_decap_8 FILLER_52_432 ();
 sg13g2_decap_8 FILLER_52_439 ();
 sg13g2_decap_8 FILLER_52_446 ();
 sg13g2_decap_4 FILLER_52_453 ();
 sg13g2_fill_1 FILLER_52_471 ();
 sg13g2_decap_8 FILLER_52_502 ();
 sg13g2_fill_2 FILLER_52_509 ();
 sg13g2_decap_4 FILLER_52_521 ();
 sg13g2_fill_1 FILLER_52_525 ();
 sg13g2_decap_8 FILLER_52_566 ();
 sg13g2_decap_8 FILLER_52_573 ();
 sg13g2_fill_1 FILLER_52_580 ();
 sg13g2_fill_2 FILLER_52_591 ();
 sg13g2_fill_1 FILLER_52_593 ();
 sg13g2_decap_4 FILLER_52_601 ();
 sg13g2_fill_2 FILLER_52_605 ();
 sg13g2_fill_2 FILLER_52_612 ();
 sg13g2_fill_1 FILLER_52_614 ();
 sg13g2_decap_4 FILLER_52_641 ();
 sg13g2_fill_2 FILLER_52_645 ();
 sg13g2_decap_4 FILLER_52_683 ();
 sg13g2_fill_1 FILLER_52_687 ();
 sg13g2_fill_2 FILLER_52_698 ();
 sg13g2_decap_8 FILLER_52_730 ();
 sg13g2_decap_8 FILLER_52_737 ();
 sg13g2_decap_4 FILLER_52_744 ();
 sg13g2_fill_1 FILLER_52_748 ();
 sg13g2_fill_2 FILLER_52_783 ();
 sg13g2_fill_1 FILLER_52_785 ();
 sg13g2_decap_4 FILLER_52_796 ();
 sg13g2_fill_2 FILLER_52_800 ();
 sg13g2_decap_8 FILLER_52_806 ();
 sg13g2_fill_2 FILLER_52_813 ();
 sg13g2_fill_2 FILLER_52_831 ();
 sg13g2_decap_4 FILLER_52_867 ();
 sg13g2_decap_4 FILLER_52_875 ();
 sg13g2_decap_8 FILLER_52_889 ();
 sg13g2_decap_8 FILLER_52_896 ();
 sg13g2_decap_8 FILLER_52_903 ();
 sg13g2_fill_2 FILLER_52_990 ();
 sg13g2_decap_8 FILLER_52_996 ();
 sg13g2_decap_8 FILLER_52_1003 ();
 sg13g2_decap_8 FILLER_52_1010 ();
 sg13g2_decap_4 FILLER_52_1017 ();
 sg13g2_fill_2 FILLER_52_1021 ();
 sg13g2_fill_2 FILLER_52_1033 ();
 sg13g2_fill_1 FILLER_52_1035 ();
 sg13g2_fill_2 FILLER_52_1062 ();
 sg13g2_fill_2 FILLER_52_1084 ();
 sg13g2_fill_1 FILLER_52_1086 ();
 sg13g2_decap_4 FILLER_52_1091 ();
 sg13g2_fill_1 FILLER_52_1095 ();
 sg13g2_decap_8 FILLER_52_1122 ();
 sg13g2_fill_2 FILLER_52_1129 ();
 sg13g2_fill_2 FILLER_52_1145 ();
 sg13g2_fill_1 FILLER_52_1147 ();
 sg13g2_fill_2 FILLER_52_1197 ();
 sg13g2_fill_1 FILLER_52_1199 ();
 sg13g2_decap_4 FILLER_52_1210 ();
 sg13g2_decap_8 FILLER_52_1218 ();
 sg13g2_decap_4 FILLER_52_1225 ();
 sg13g2_fill_1 FILLER_52_1229 ();
 sg13g2_decap_8 FILLER_52_1234 ();
 sg13g2_decap_8 FILLER_52_1241 ();
 sg13g2_fill_1 FILLER_52_1248 ();
 sg13g2_decap_4 FILLER_52_1259 ();
 sg13g2_fill_1 FILLER_52_1263 ();
 sg13g2_decap_8 FILLER_52_1272 ();
 sg13g2_decap_8 FILLER_52_1279 ();
 sg13g2_decap_8 FILLER_52_1286 ();
 sg13g2_decap_8 FILLER_52_1293 ();
 sg13g2_decap_8 FILLER_52_1300 ();
 sg13g2_fill_2 FILLER_52_1321 ();
 sg13g2_fill_1 FILLER_52_1323 ();
 sg13g2_decap_4 FILLER_52_1328 ();
 sg13g2_decap_8 FILLER_52_1340 ();
 sg13g2_fill_1 FILLER_52_1347 ();
 sg13g2_fill_2 FILLER_52_1393 ();
 sg13g2_decap_4 FILLER_52_1431 ();
 sg13g2_decap_8 FILLER_52_1439 ();
 sg13g2_fill_2 FILLER_52_1446 ();
 sg13g2_decap_8 FILLER_52_1452 ();
 sg13g2_decap_8 FILLER_52_1459 ();
 sg13g2_fill_2 FILLER_52_1466 ();
 sg13g2_decap_4 FILLER_52_1508 ();
 sg13g2_fill_2 FILLER_52_1512 ();
 sg13g2_decap_8 FILLER_52_1540 ();
 sg13g2_decap_4 FILLER_52_1547 ();
 sg13g2_fill_1 FILLER_52_1551 ();
 sg13g2_decap_8 FILLER_52_1562 ();
 sg13g2_decap_4 FILLER_52_1569 ();
 sg13g2_fill_1 FILLER_52_1573 ();
 sg13g2_fill_2 FILLER_52_1584 ();
 sg13g2_decap_8 FILLER_52_1616 ();
 sg13g2_decap_8 FILLER_52_1623 ();
 sg13g2_decap_8 FILLER_52_1630 ();
 sg13g2_decap_4 FILLER_52_1637 ();
 sg13g2_fill_2 FILLER_52_1641 ();
 sg13g2_decap_8 FILLER_52_1647 ();
 sg13g2_decap_8 FILLER_52_1654 ();
 sg13g2_decap_4 FILLER_52_1661 ();
 sg13g2_fill_1 FILLER_52_1665 ();
 sg13g2_decap_8 FILLER_52_1692 ();
 sg13g2_fill_1 FILLER_52_1699 ();
 sg13g2_decap_8 FILLER_52_1726 ();
 sg13g2_decap_8 FILLER_52_1767 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_18 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_fill_2 FILLER_53_115 ();
 sg13g2_fill_1 FILLER_53_117 ();
 sg13g2_decap_4 FILLER_53_131 ();
 sg13g2_decap_8 FILLER_53_161 ();
 sg13g2_decap_4 FILLER_53_168 ();
 sg13g2_fill_2 FILLER_53_172 ();
 sg13g2_fill_2 FILLER_53_184 ();
 sg13g2_fill_1 FILLER_53_186 ();
 sg13g2_decap_4 FILLER_53_200 ();
 sg13g2_fill_1 FILLER_53_204 ();
 sg13g2_decap_4 FILLER_53_229 ();
 sg13g2_fill_2 FILLER_53_233 ();
 sg13g2_decap_8 FILLER_53_240 ();
 sg13g2_decap_8 FILLER_53_247 ();
 sg13g2_decap_8 FILLER_53_254 ();
 sg13g2_decap_8 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_268 ();
 sg13g2_fill_1 FILLER_53_310 ();
 sg13g2_decap_8 FILLER_53_321 ();
 sg13g2_decap_8 FILLER_53_328 ();
 sg13g2_decap_8 FILLER_53_335 ();
 sg13g2_decap_8 FILLER_53_342 ();
 sg13g2_fill_2 FILLER_53_349 ();
 sg13g2_decap_4 FILLER_53_355 ();
 sg13g2_fill_1 FILLER_53_389 ();
 sg13g2_fill_2 FILLER_53_398 ();
 sg13g2_decap_8 FILLER_53_487 ();
 sg13g2_decap_8 FILLER_53_494 ();
 sg13g2_decap_4 FILLER_53_501 ();
 sg13g2_fill_1 FILLER_53_505 ();
 sg13g2_decap_8 FILLER_53_542 ();
 sg13g2_decap_8 FILLER_53_549 ();
 sg13g2_decap_8 FILLER_53_556 ();
 sg13g2_fill_1 FILLER_53_563 ();
 sg13g2_fill_1 FILLER_53_568 ();
 sg13g2_fill_1 FILLER_53_579 ();
 sg13g2_fill_1 FILLER_53_584 ();
 sg13g2_fill_2 FILLER_53_611 ();
 sg13g2_decap_8 FILLER_53_681 ();
 sg13g2_fill_2 FILLER_53_688 ();
 sg13g2_fill_2 FILLER_53_698 ();
 sg13g2_fill_1 FILLER_53_700 ();
 sg13g2_decap_8 FILLER_53_737 ();
 sg13g2_decap_8 FILLER_53_744 ();
 sg13g2_fill_2 FILLER_53_751 ();
 sg13g2_fill_1 FILLER_53_753 ();
 sg13g2_fill_2 FILLER_53_778 ();
 sg13g2_fill_1 FILLER_53_780 ();
 sg13g2_decap_4 FILLER_53_807 ();
 sg13g2_decap_4 FILLER_53_815 ();
 sg13g2_fill_2 FILLER_53_828 ();
 sg13g2_fill_1 FILLER_53_830 ();
 sg13g2_fill_1 FILLER_53_867 ();
 sg13g2_fill_1 FILLER_53_874 ();
 sg13g2_fill_2 FILLER_53_879 ();
 sg13g2_fill_2 FILLER_53_886 ();
 sg13g2_fill_2 FILLER_53_898 ();
 sg13g2_fill_1 FILLER_53_900 ();
 sg13g2_fill_2 FILLER_53_921 ();
 sg13g2_fill_1 FILLER_53_933 ();
 sg13g2_fill_2 FILLER_53_979 ();
 sg13g2_fill_2 FILLER_53_991 ();
 sg13g2_fill_1 FILLER_53_993 ();
 sg13g2_fill_2 FILLER_53_1020 ();
 sg13g2_fill_1 FILLER_53_1062 ();
 sg13g2_fill_1 FILLER_53_1073 ();
 sg13g2_fill_1 FILLER_53_1110 ();
 sg13g2_fill_2 FILLER_53_1121 ();
 sg13g2_decap_8 FILLER_53_1133 ();
 sg13g2_decap_8 FILLER_53_1140 ();
 sg13g2_decap_8 FILLER_53_1147 ();
 sg13g2_decap_8 FILLER_53_1154 ();
 sg13g2_decap_8 FILLER_53_1161 ();
 sg13g2_decap_8 FILLER_53_1168 ();
 sg13g2_decap_8 FILLER_53_1179 ();
 sg13g2_fill_2 FILLER_53_1186 ();
 sg13g2_decap_8 FILLER_53_1214 ();
 sg13g2_fill_2 FILLER_53_1221 ();
 sg13g2_fill_1 FILLER_53_1223 ();
 sg13g2_decap_4 FILLER_53_1232 ();
 sg13g2_fill_1 FILLER_53_1236 ();
 sg13g2_decap_8 FILLER_53_1263 ();
 sg13g2_fill_1 FILLER_53_1270 ();
 sg13g2_decap_8 FILLER_53_1297 ();
 sg13g2_decap_8 FILLER_53_1304 ();
 sg13g2_fill_1 FILLER_53_1311 ();
 sg13g2_decap_8 FILLER_53_1322 ();
 sg13g2_decap_8 FILLER_53_1355 ();
 sg13g2_decap_8 FILLER_53_1362 ();
 sg13g2_fill_1 FILLER_53_1369 ();
 sg13g2_fill_2 FILLER_53_1374 ();
 sg13g2_fill_1 FILLER_53_1376 ();
 sg13g2_fill_1 FILLER_53_1417 ();
 sg13g2_decap_8 FILLER_53_1422 ();
 sg13g2_fill_2 FILLER_53_1429 ();
 sg13g2_decap_8 FILLER_53_1467 ();
 sg13g2_fill_1 FILLER_53_1474 ();
 sg13g2_fill_2 FILLER_53_1478 ();
 sg13g2_decap_8 FILLER_53_1484 ();
 sg13g2_decap_8 FILLER_53_1491 ();
 sg13g2_decap_8 FILLER_53_1498 ();
 sg13g2_decap_8 FILLER_53_1505 ();
 sg13g2_fill_1 FILLER_53_1512 ();
 sg13g2_decap_8 FILLER_53_1575 ();
 sg13g2_decap_8 FILLER_53_1582 ();
 sg13g2_fill_1 FILLER_53_1589 ();
 sg13g2_decap_8 FILLER_53_1598 ();
 sg13g2_decap_8 FILLER_53_1605 ();
 sg13g2_fill_1 FILLER_53_1612 ();
 sg13g2_decap_8 FILLER_53_1617 ();
 sg13g2_decap_8 FILLER_53_1624 ();
 sg13g2_decap_8 FILLER_53_1631 ();
 sg13g2_decap_8 FILLER_53_1638 ();
 sg13g2_decap_8 FILLER_53_1645 ();
 sg13g2_decap_8 FILLER_53_1652 ();
 sg13g2_decap_8 FILLER_53_1659 ();
 sg13g2_decap_8 FILLER_53_1666 ();
 sg13g2_fill_1 FILLER_53_1673 ();
 sg13g2_decap_8 FILLER_53_1678 ();
 sg13g2_decap_8 FILLER_53_1685 ();
 sg13g2_fill_2 FILLER_53_1692 ();
 sg13g2_fill_1 FILLER_53_1694 ();
 sg13g2_decap_4 FILLER_53_1705 ();
 sg13g2_decap_8 FILLER_53_1713 ();
 sg13g2_decap_8 FILLER_53_1720 ();
 sg13g2_fill_2 FILLER_53_1727 ();
 sg13g2_fill_1 FILLER_53_1729 ();
 sg13g2_decap_8 FILLER_53_1760 ();
 sg13g2_decap_8 FILLER_53_1767 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_16 ();
 sg13g2_fill_1 FILLER_54_43 ();
 sg13g2_fill_2 FILLER_54_54 ();
 sg13g2_fill_2 FILLER_54_60 ();
 sg13g2_decap_4 FILLER_54_88 ();
 sg13g2_decap_8 FILLER_54_102 ();
 sg13g2_fill_2 FILLER_54_109 ();
 sg13g2_fill_1 FILLER_54_111 ();
 sg13g2_fill_2 FILLER_54_134 ();
 sg13g2_fill_1 FILLER_54_136 ();
 sg13g2_fill_1 FILLER_54_141 ();
 sg13g2_fill_1 FILLER_54_146 ();
 sg13g2_decap_8 FILLER_54_155 ();
 sg13g2_fill_2 FILLER_54_162 ();
 sg13g2_fill_2 FILLER_54_184 ();
 sg13g2_fill_1 FILLER_54_186 ();
 sg13g2_fill_2 FILLER_54_195 ();
 sg13g2_fill_2 FILLER_54_207 ();
 sg13g2_fill_2 FILLER_54_238 ();
 sg13g2_fill_2 FILLER_54_250 ();
 sg13g2_fill_1 FILLER_54_282 ();
 sg13g2_fill_1 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_320 ();
 sg13g2_fill_1 FILLER_54_347 ();
 sg13g2_fill_2 FILLER_54_374 ();
 sg13g2_decap_4 FILLER_54_386 ();
 sg13g2_fill_1 FILLER_54_390 ();
 sg13g2_fill_2 FILLER_54_405 ();
 sg13g2_decap_8 FILLER_54_432 ();
 sg13g2_decap_8 FILLER_54_439 ();
 sg13g2_decap_8 FILLER_54_446 ();
 sg13g2_decap_8 FILLER_54_453 ();
 sg13g2_decap_4 FILLER_54_460 ();
 sg13g2_decap_8 FILLER_54_490 ();
 sg13g2_decap_8 FILLER_54_497 ();
 sg13g2_decap_8 FILLER_54_504 ();
 sg13g2_fill_1 FILLER_54_511 ();
 sg13g2_decap_8 FILLER_54_538 ();
 sg13g2_decap_4 FILLER_54_545 ();
 sg13g2_decap_4 FILLER_54_553 ();
 sg13g2_fill_1 FILLER_54_557 ();
 sg13g2_fill_2 FILLER_54_594 ();
 sg13g2_fill_2 FILLER_54_600 ();
 sg13g2_fill_1 FILLER_54_602 ();
 sg13g2_fill_1 FILLER_54_609 ();
 sg13g2_fill_2 FILLER_54_620 ();
 sg13g2_fill_2 FILLER_54_626 ();
 sg13g2_fill_1 FILLER_54_628 ();
 sg13g2_fill_1 FILLER_54_633 ();
 sg13g2_fill_2 FILLER_54_644 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_decap_4 FILLER_54_677 ();
 sg13g2_fill_2 FILLER_54_681 ();
 sg13g2_decap_8 FILLER_54_727 ();
 sg13g2_decap_8 FILLER_54_734 ();
 sg13g2_decap_8 FILLER_54_741 ();
 sg13g2_decap_8 FILLER_54_748 ();
 sg13g2_decap_4 FILLER_54_755 ();
 sg13g2_fill_1 FILLER_54_759 ();
 sg13g2_decap_4 FILLER_54_770 ();
 sg13g2_fill_1 FILLER_54_774 ();
 sg13g2_fill_2 FILLER_54_785 ();
 sg13g2_fill_1 FILLER_54_787 ();
 sg13g2_fill_1 FILLER_54_792 ();
 sg13g2_decap_8 FILLER_54_825 ();
 sg13g2_fill_2 FILLER_54_842 ();
 sg13g2_fill_2 FILLER_54_848 ();
 sg13g2_decap_4 FILLER_54_876 ();
 sg13g2_decap_8 FILLER_54_905 ();
 sg13g2_fill_1 FILLER_54_912 ();
 sg13g2_decap_8 FILLER_54_1082 ();
 sg13g2_fill_2 FILLER_54_1089 ();
 sg13g2_fill_1 FILLER_54_1095 ();
 sg13g2_decap_4 FILLER_54_1100 ();
 sg13g2_fill_2 FILLER_54_1116 ();
 sg13g2_fill_1 FILLER_54_1118 ();
 sg13g2_fill_1 FILLER_54_1158 ();
 sg13g2_fill_1 FILLER_54_1195 ();
 sg13g2_fill_1 FILLER_54_1200 ();
 sg13g2_fill_1 FILLER_54_1209 ();
 sg13g2_fill_1 FILLER_54_1220 ();
 sg13g2_fill_2 FILLER_54_1247 ();
 sg13g2_decap_4 FILLER_54_1289 ();
 sg13g2_fill_2 FILLER_54_1293 ();
 sg13g2_fill_2 FILLER_54_1324 ();
 sg13g2_fill_1 FILLER_54_1326 ();
 sg13g2_fill_2 FILLER_54_1367 ();
 sg13g2_decap_8 FILLER_54_1373 ();
 sg13g2_decap_8 FILLER_54_1380 ();
 sg13g2_decap_8 FILLER_54_1387 ();
 sg13g2_decap_4 FILLER_54_1394 ();
 sg13g2_decap_8 FILLER_54_1402 ();
 sg13g2_fill_2 FILLER_54_1409 ();
 sg13g2_decap_8 FILLER_54_1437 ();
 sg13g2_decap_4 FILLER_54_1444 ();
 sg13g2_decap_8 FILLER_54_1452 ();
 sg13g2_decap_8 FILLER_54_1459 ();
 sg13g2_fill_2 FILLER_54_1466 ();
 sg13g2_fill_2 FILLER_54_1485 ();
 sg13g2_decap_8 FILLER_54_1491 ();
 sg13g2_decap_8 FILLER_54_1498 ();
 sg13g2_decap_8 FILLER_54_1505 ();
 sg13g2_decap_4 FILLER_54_1512 ();
 sg13g2_fill_1 FILLER_54_1516 ();
 sg13g2_decap_8 FILLER_54_1545 ();
 sg13g2_fill_2 FILLER_54_1552 ();
 sg13g2_fill_1 FILLER_54_1554 ();
 sg13g2_decap_8 FILLER_54_1670 ();
 sg13g2_fill_1 FILLER_54_1677 ();
 sg13g2_decap_8 FILLER_54_1683 ();
 sg13g2_decap_8 FILLER_54_1690 ();
 sg13g2_decap_8 FILLER_54_1697 ();
 sg13g2_decap_8 FILLER_54_1704 ();
 sg13g2_decap_8 FILLER_54_1711 ();
 sg13g2_decap_8 FILLER_54_1718 ();
 sg13g2_decap_8 FILLER_54_1725 ();
 sg13g2_fill_1 FILLER_54_1732 ();
 sg13g2_decap_8 FILLER_54_1759 ();
 sg13g2_decap_8 FILLER_54_1766 ();
 sg13g2_fill_1 FILLER_54_1773 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_46 ();
 sg13g2_decap_8 FILLER_55_53 ();
 sg13g2_decap_4 FILLER_55_60 ();
 sg13g2_fill_1 FILLER_55_64 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_4 FILLER_55_77 ();
 sg13g2_fill_2 FILLER_55_81 ();
 sg13g2_decap_8 FILLER_55_103 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_decap_8 FILLER_55_135 ();
 sg13g2_decap_8 FILLER_55_172 ();
 sg13g2_decap_4 FILLER_55_179 ();
 sg13g2_fill_1 FILLER_55_183 ();
 sg13g2_decap_8 FILLER_55_188 ();
 sg13g2_decap_4 FILLER_55_195 ();
 sg13g2_fill_1 FILLER_55_199 ();
 sg13g2_fill_1 FILLER_55_208 ();
 sg13g2_fill_2 FILLER_55_238 ();
 sg13g2_fill_2 FILLER_55_244 ();
 sg13g2_decap_8 FILLER_55_252 ();
 sg13g2_decap_8 FILLER_55_259 ();
 sg13g2_decap_4 FILLER_55_266 ();
 sg13g2_fill_2 FILLER_55_284 ();
 sg13g2_fill_2 FILLER_55_300 ();
 sg13g2_fill_2 FILLER_55_306 ();
 sg13g2_fill_1 FILLER_55_308 ();
 sg13g2_fill_2 FILLER_55_313 ();
 sg13g2_fill_1 FILLER_55_315 ();
 sg13g2_fill_2 FILLER_55_326 ();
 sg13g2_fill_1 FILLER_55_328 ();
 sg13g2_decap_4 FILLER_55_333 ();
 sg13g2_fill_1 FILLER_55_337 ();
 sg13g2_fill_2 FILLER_55_404 ();
 sg13g2_fill_1 FILLER_55_416 ();
 sg13g2_fill_2 FILLER_55_447 ();
 sg13g2_decap_8 FILLER_55_495 ();
 sg13g2_decap_8 FILLER_55_502 ();
 sg13g2_decap_8 FILLER_55_509 ();
 sg13g2_decap_4 FILLER_55_516 ();
 sg13g2_fill_2 FILLER_55_520 ();
 sg13g2_decap_8 FILLER_55_530 ();
 sg13g2_decap_4 FILLER_55_537 ();
 sg13g2_fill_1 FILLER_55_541 ();
 sg13g2_decap_8 FILLER_55_588 ();
 sg13g2_fill_1 FILLER_55_595 ();
 sg13g2_decap_8 FILLER_55_606 ();
 sg13g2_fill_1 FILLER_55_613 ();
 sg13g2_fill_2 FILLER_55_632 ();
 sg13g2_decap_8 FILLER_55_644 ();
 sg13g2_fill_1 FILLER_55_651 ();
 sg13g2_fill_1 FILLER_55_656 ();
 sg13g2_fill_2 FILLER_55_674 ();
 sg13g2_decap_8 FILLER_55_686 ();
 sg13g2_fill_1 FILLER_55_693 ();
 sg13g2_decap_4 FILLER_55_698 ();
 sg13g2_fill_1 FILLER_55_702 ();
 sg13g2_fill_2 FILLER_55_724 ();
 sg13g2_fill_1 FILLER_55_726 ();
 sg13g2_fill_2 FILLER_55_747 ();
 sg13g2_decap_8 FILLER_55_759 ();
 sg13g2_decap_4 FILLER_55_766 ();
 sg13g2_fill_1 FILLER_55_816 ();
 sg13g2_fill_1 FILLER_55_823 ();
 sg13g2_fill_1 FILLER_55_828 ();
 sg13g2_fill_1 FILLER_55_855 ();
 sg13g2_decap_8 FILLER_55_882 ();
 sg13g2_decap_4 FILLER_55_889 ();
 sg13g2_fill_1 FILLER_55_893 ();
 sg13g2_decap_8 FILLER_55_898 ();
 sg13g2_decap_8 FILLER_55_905 ();
 sg13g2_decap_8 FILLER_55_912 ();
 sg13g2_fill_1 FILLER_55_924 ();
 sg13g2_fill_1 FILLER_55_936 ();
 sg13g2_fill_1 FILLER_55_951 ();
 sg13g2_decap_8 FILLER_55_981 ();
 sg13g2_fill_2 FILLER_55_998 ();
 sg13g2_fill_2 FILLER_55_1004 ();
 sg13g2_fill_2 FILLER_55_1010 ();
 sg13g2_fill_1 FILLER_55_1012 ();
 sg13g2_fill_1 FILLER_55_1023 ();
 sg13g2_fill_2 FILLER_55_1034 ();
 sg13g2_fill_1 FILLER_55_1036 ();
 sg13g2_fill_2 FILLER_55_1047 ();
 sg13g2_fill_1 FILLER_55_1049 ();
 sg13g2_fill_1 FILLER_55_1054 ();
 sg13g2_decap_8 FILLER_55_1127 ();
 sg13g2_decap_4 FILLER_55_1134 ();
 sg13g2_fill_1 FILLER_55_1138 ();
 sg13g2_fill_2 FILLER_55_1143 ();
 sg13g2_fill_1 FILLER_55_1145 ();
 sg13g2_fill_1 FILLER_55_1176 ();
 sg13g2_decap_8 FILLER_55_1187 ();
 sg13g2_decap_8 FILLER_55_1194 ();
 sg13g2_decap_4 FILLER_55_1201 ();
 sg13g2_fill_1 FILLER_55_1205 ();
 sg13g2_fill_1 FILLER_55_1227 ();
 sg13g2_fill_1 FILLER_55_1232 ();
 sg13g2_fill_1 FILLER_55_1243 ();
 sg13g2_fill_2 FILLER_55_1248 ();
 sg13g2_decap_8 FILLER_55_1281 ();
 sg13g2_decap_4 FILLER_55_1288 ();
 sg13g2_fill_2 FILLER_55_1292 ();
 sg13g2_fill_1 FILLER_55_1304 ();
 sg13g2_fill_1 FILLER_55_1309 ();
 sg13g2_fill_1 FILLER_55_1320 ();
 sg13g2_fill_1 FILLER_55_1342 ();
 sg13g2_fill_2 FILLER_55_1347 ();
 sg13g2_decap_8 FILLER_55_1385 ();
 sg13g2_decap_8 FILLER_55_1392 ();
 sg13g2_fill_2 FILLER_55_1399 ();
 sg13g2_decap_8 FILLER_55_1411 ();
 sg13g2_decap_4 FILLER_55_1418 ();
 sg13g2_fill_2 FILLER_55_1422 ();
 sg13g2_decap_8 FILLER_55_1427 ();
 sg13g2_decap_8 FILLER_55_1434 ();
 sg13g2_decap_8 FILLER_55_1504 ();
 sg13g2_decap_8 FILLER_55_1511 ();
 sg13g2_decap_8 FILLER_55_1518 ();
 sg13g2_fill_1 FILLER_55_1525 ();
 sg13g2_fill_1 FILLER_55_1538 ();
 sg13g2_fill_2 FILLER_55_1573 ();
 sg13g2_fill_2 FILLER_55_1589 ();
 sg13g2_fill_1 FILLER_55_1591 ();
 sg13g2_decap_8 FILLER_55_1606 ();
 sg13g2_decap_8 FILLER_55_1613 ();
 sg13g2_fill_1 FILLER_55_1620 ();
 sg13g2_fill_1 FILLER_55_1631 ();
 sg13g2_fill_2 FILLER_55_1658 ();
 sg13g2_fill_2 FILLER_55_1664 ();
 sg13g2_fill_2 FILLER_55_1671 ();
 sg13g2_decap_8 FILLER_55_1761 ();
 sg13g2_decap_4 FILLER_55_1768 ();
 sg13g2_fill_2 FILLER_55_1772 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_11 ();
 sg13g2_decap_8 FILLER_56_48 ();
 sg13g2_decap_8 FILLER_56_55 ();
 sg13g2_decap_8 FILLER_56_67 ();
 sg13g2_decap_8 FILLER_56_95 ();
 sg13g2_decap_8 FILLER_56_102 ();
 sg13g2_decap_8 FILLER_56_109 ();
 sg13g2_decap_4 FILLER_56_116 ();
 sg13g2_fill_2 FILLER_56_120 ();
 sg13g2_decap_8 FILLER_56_136 ();
 sg13g2_decap_8 FILLER_56_143 ();
 sg13g2_decap_8 FILLER_56_150 ();
 sg13g2_decap_8 FILLER_56_157 ();
 sg13g2_decap_8 FILLER_56_164 ();
 sg13g2_decap_4 FILLER_56_171 ();
 sg13g2_fill_2 FILLER_56_175 ();
 sg13g2_fill_1 FILLER_56_203 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_fill_2 FILLER_56_216 ();
 sg13g2_fill_2 FILLER_56_222 ();
 sg13g2_decap_4 FILLER_56_259 ();
 sg13g2_fill_2 FILLER_56_263 ();
 sg13g2_fill_2 FILLER_56_269 ();
 sg13g2_decap_8 FILLER_56_337 ();
 sg13g2_fill_1 FILLER_56_344 ();
 sg13g2_fill_2 FILLER_56_419 ();
 sg13g2_fill_1 FILLER_56_421 ();
 sg13g2_decap_4 FILLER_56_457 ();
 sg13g2_fill_2 FILLER_56_471 ();
 sg13g2_fill_2 FILLER_56_477 ();
 sg13g2_fill_1 FILLER_56_479 ();
 sg13g2_fill_2 FILLER_56_484 ();
 sg13g2_fill_1 FILLER_56_486 ();
 sg13g2_decap_4 FILLER_56_491 ();
 sg13g2_fill_2 FILLER_56_495 ();
 sg13g2_fill_2 FILLER_56_507 ();
 sg13g2_fill_1 FILLER_56_509 ();
 sg13g2_fill_2 FILLER_56_540 ();
 sg13g2_decap_8 FILLER_56_556 ();
 sg13g2_decap_8 FILLER_56_563 ();
 sg13g2_decap_4 FILLER_56_583 ();
 sg13g2_fill_2 FILLER_56_587 ();
 sg13g2_decap_8 FILLER_56_595 ();
 sg13g2_decap_8 FILLER_56_602 ();
 sg13g2_fill_1 FILLER_56_620 ();
 sg13g2_fill_1 FILLER_56_631 ();
 sg13g2_decap_8 FILLER_56_642 ();
 sg13g2_fill_1 FILLER_56_654 ();
 sg13g2_fill_2 FILLER_56_684 ();
 sg13g2_fill_2 FILLER_56_706 ();
 sg13g2_fill_1 FILLER_56_758 ();
 sg13g2_fill_2 FILLER_56_785 ();
 sg13g2_fill_1 FILLER_56_787 ();
 sg13g2_decap_8 FILLER_56_814 ();
 sg13g2_fill_2 FILLER_56_821 ();
 sg13g2_fill_1 FILLER_56_847 ();
 sg13g2_decap_4 FILLER_56_858 ();
 sg13g2_fill_2 FILLER_56_862 ();
 sg13g2_decap_4 FILLER_56_868 ();
 sg13g2_fill_2 FILLER_56_872 ();
 sg13g2_fill_2 FILLER_56_884 ();
 sg13g2_fill_1 FILLER_56_886 ();
 sg13g2_fill_2 FILLER_56_924 ();
 sg13g2_fill_1 FILLER_56_931 ();
 sg13g2_fill_2 FILLER_56_976 ();
 sg13g2_decap_8 FILLER_56_989 ();
 sg13g2_decap_8 FILLER_56_996 ();
 sg13g2_decap_8 FILLER_56_1003 ();
 sg13g2_decap_8 FILLER_56_1010 ();
 sg13g2_decap_4 FILLER_56_1017 ();
 sg13g2_fill_1 FILLER_56_1021 ();
 sg13g2_decap_8 FILLER_56_1034 ();
 sg13g2_fill_2 FILLER_56_1041 ();
 sg13g2_fill_1 FILLER_56_1043 ();
 sg13g2_fill_2 FILLER_56_1079 ();
 sg13g2_decap_4 FILLER_56_1120 ();
 sg13g2_fill_1 FILLER_56_1124 ();
 sg13g2_decap_4 FILLER_56_1151 ();
 sg13g2_fill_2 FILLER_56_1155 ();
 sg13g2_decap_4 FILLER_56_1167 ();
 sg13g2_decap_4 FILLER_56_1220 ();
 sg13g2_fill_1 FILLER_56_1228 ();
 sg13g2_fill_2 FILLER_56_1264 ();
 sg13g2_fill_1 FILLER_56_1266 ();
 sg13g2_decap_4 FILLER_56_1271 ();
 sg13g2_fill_1 FILLER_56_1275 ();
 sg13g2_fill_2 FILLER_56_1286 ();
 sg13g2_decap_4 FILLER_56_1314 ();
 sg13g2_fill_1 FILLER_56_1318 ();
 sg13g2_decap_8 FILLER_56_1401 ();
 sg13g2_decap_8 FILLER_56_1408 ();
 sg13g2_decap_8 FILLER_56_1415 ();
 sg13g2_fill_2 FILLER_56_1422 ();
 sg13g2_fill_1 FILLER_56_1428 ();
 sg13g2_decap_4 FILLER_56_1433 ();
 sg13g2_fill_1 FILLER_56_1437 ();
 sg13g2_decap_8 FILLER_56_1453 ();
 sg13g2_decap_4 FILLER_56_1460 ();
 sg13g2_fill_2 FILLER_56_1471 ();
 sg13g2_decap_4 FILLER_56_1517 ();
 sg13g2_fill_2 FILLER_56_1521 ();
 sg13g2_decap_4 FILLER_56_1527 ();
 sg13g2_fill_2 FILLER_56_1531 ();
 sg13g2_fill_1 FILLER_56_1537 ();
 sg13g2_fill_2 FILLER_56_1548 ();
 sg13g2_fill_1 FILLER_56_1652 ();
 sg13g2_fill_1 FILLER_56_1679 ();
 sg13g2_fill_1 FILLER_56_1706 ();
 sg13g2_fill_1 FILLER_56_1743 ();
 sg13g2_decap_4 FILLER_56_1770 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_11 ();
 sg13g2_fill_1 FILLER_57_49 ();
 sg13g2_fill_1 FILLER_57_76 ();
 sg13g2_fill_1 FILLER_57_87 ();
 sg13g2_fill_1 FILLER_57_114 ();
 sg13g2_fill_2 FILLER_57_151 ();
 sg13g2_fill_2 FILLER_57_163 ();
 sg13g2_fill_1 FILLER_57_165 ();
 sg13g2_fill_1 FILLER_57_170 ();
 sg13g2_fill_2 FILLER_57_181 ();
 sg13g2_fill_1 FILLER_57_183 ();
 sg13g2_fill_2 FILLER_57_204 ();
 sg13g2_decap_4 FILLER_57_241 ();
 sg13g2_decap_4 FILLER_57_249 ();
 sg13g2_fill_1 FILLER_57_263 ();
 sg13g2_decap_4 FILLER_57_270 ();
 sg13g2_fill_2 FILLER_57_274 ();
 sg13g2_decap_4 FILLER_57_302 ();
 sg13g2_fill_1 FILLER_57_327 ();
 sg13g2_fill_2 FILLER_57_354 ();
 sg13g2_fill_2 FILLER_57_360 ();
 sg13g2_fill_1 FILLER_57_372 ();
 sg13g2_decap_8 FILLER_57_412 ();
 sg13g2_decap_4 FILLER_57_419 ();
 sg13g2_fill_1 FILLER_57_423 ();
 sg13g2_fill_1 FILLER_57_428 ();
 sg13g2_fill_1 FILLER_57_474 ();
 sg13g2_decap_4 FILLER_57_501 ();
 sg13g2_decap_4 FILLER_57_508 ();
 sg13g2_fill_1 FILLER_57_512 ();
 sg13g2_decap_4 FILLER_57_530 ();
 sg13g2_fill_1 FILLER_57_534 ();
 sg13g2_fill_2 FILLER_57_567 ();
 sg13g2_decap_8 FILLER_57_575 ();
 sg13g2_fill_1 FILLER_57_582 ();
 sg13g2_fill_2 FILLER_57_588 ();
 sg13g2_fill_1 FILLER_57_590 ();
 sg13g2_decap_4 FILLER_57_599 ();
 sg13g2_fill_1 FILLER_57_603 ();
 sg13g2_decap_4 FILLER_57_645 ();
 sg13g2_fill_1 FILLER_57_666 ();
 sg13g2_fill_1 FILLER_57_693 ();
 sg13g2_fill_1 FILLER_57_726 ();
 sg13g2_decap_4 FILLER_57_763 ();
 sg13g2_fill_2 FILLER_57_771 ();
 sg13g2_fill_1 FILLER_57_777 ();
 sg13g2_decap_8 FILLER_57_798 ();
 sg13g2_fill_1 FILLER_57_851 ();
 sg13g2_decap_8 FILLER_57_864 ();
 sg13g2_decap_8 FILLER_57_871 ();
 sg13g2_decap_8 FILLER_57_878 ();
 sg13g2_fill_1 FILLER_57_885 ();
 sg13g2_decap_8 FILLER_57_895 ();
 sg13g2_fill_2 FILLER_57_902 ();
 sg13g2_fill_1 FILLER_57_909 ();
 sg13g2_fill_1 FILLER_57_927 ();
 sg13g2_fill_1 FILLER_57_984 ();
 sg13g2_decap_4 FILLER_57_1011 ();
 sg13g2_fill_1 FILLER_57_1015 ();
 sg13g2_decap_8 FILLER_57_1047 ();
 sg13g2_fill_1 FILLER_57_1054 ();
 sg13g2_decap_8 FILLER_57_1091 ();
 sg13g2_decap_8 FILLER_57_1098 ();
 sg13g2_decap_8 FILLER_57_1125 ();
 sg13g2_decap_4 FILLER_57_1132 ();
 sg13g2_decap_8 FILLER_57_1162 ();
 sg13g2_decap_8 FILLER_57_1169 ();
 sg13g2_fill_2 FILLER_57_1176 ();
 sg13g2_fill_1 FILLER_57_1182 ();
 sg13g2_decap_8 FILLER_57_1193 ();
 sg13g2_fill_1 FILLER_57_1200 ();
 sg13g2_decap_8 FILLER_57_1209 ();
 sg13g2_decap_8 FILLER_57_1216 ();
 sg13g2_decap_8 FILLER_57_1223 ();
 sg13g2_decap_8 FILLER_57_1230 ();
 sg13g2_decap_8 FILLER_57_1237 ();
 sg13g2_decap_8 FILLER_57_1254 ();
 sg13g2_decap_4 FILLER_57_1261 ();
 sg13g2_fill_1 FILLER_57_1265 ();
 sg13g2_fill_2 FILLER_57_1292 ();
 sg13g2_fill_1 FILLER_57_1294 ();
 sg13g2_decap_8 FILLER_57_1299 ();
 sg13g2_decap_8 FILLER_57_1306 ();
 sg13g2_fill_2 FILLER_57_1313 ();
 sg13g2_decap_4 FILLER_57_1408 ();
 sg13g2_decap_8 FILLER_57_1448 ();
 sg13g2_decap_8 FILLER_57_1455 ();
 sg13g2_decap_8 FILLER_57_1462 ();
 sg13g2_decap_4 FILLER_57_1469 ();
 sg13g2_fill_2 FILLER_57_1473 ();
 sg13g2_fill_2 FILLER_57_1478 ();
 sg13g2_decap_4 FILLER_57_1484 ();
 sg13g2_fill_2 FILLER_57_1488 ();
 sg13g2_decap_8 FILLER_57_1499 ();
 sg13g2_fill_2 FILLER_57_1552 ();
 sg13g2_fill_1 FILLER_57_1592 ();
 sg13g2_fill_2 FILLER_57_1603 ();
 sg13g2_fill_1 FILLER_57_1605 ();
 sg13g2_fill_2 FILLER_57_1616 ();
 sg13g2_fill_1 FILLER_57_1618 ();
 sg13g2_decap_8 FILLER_57_1623 ();
 sg13g2_decap_4 FILLER_57_1634 ();
 sg13g2_fill_1 FILLER_57_1638 ();
 sg13g2_decap_4 FILLER_57_1657 ();
 sg13g2_fill_2 FILLER_57_1661 ();
 sg13g2_fill_1 FILLER_57_1691 ();
 sg13g2_fill_2 FILLER_57_1715 ();
 sg13g2_fill_1 FILLER_57_1721 ();
 sg13g2_decap_8 FILLER_57_1758 ();
 sg13g2_decap_8 FILLER_57_1765 ();
 sg13g2_fill_2 FILLER_57_1772 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_9 ();
 sg13g2_fill_1 FILLER_58_20 ();
 sg13g2_fill_1 FILLER_58_25 ();
 sg13g2_fill_2 FILLER_58_30 ();
 sg13g2_fill_2 FILLER_58_58 ();
 sg13g2_fill_2 FILLER_58_64 ();
 sg13g2_fill_1 FILLER_58_66 ();
 sg13g2_fill_1 FILLER_58_159 ();
 sg13g2_fill_1 FILLER_58_186 ();
 sg13g2_fill_1 FILLER_58_201 ();
 sg13g2_decap_4 FILLER_58_208 ();
 sg13g2_fill_1 FILLER_58_212 ();
 sg13g2_fill_2 FILLER_58_236 ();
 sg13g2_decap_4 FILLER_58_276 ();
 sg13g2_fill_1 FILLER_58_280 ();
 sg13g2_decap_4 FILLER_58_285 ();
 sg13g2_fill_1 FILLER_58_289 ();
 sg13g2_decap_8 FILLER_58_305 ();
 sg13g2_fill_1 FILLER_58_373 ();
 sg13g2_decap_4 FILLER_58_400 ();
 sg13g2_decap_8 FILLER_58_414 ();
 sg13g2_decap_4 FILLER_58_421 ();
 sg13g2_fill_2 FILLER_58_425 ();
 sg13g2_fill_2 FILLER_58_447 ();
 sg13g2_fill_2 FILLER_58_505 ();
 sg13g2_fill_1 FILLER_58_557 ();
 sg13g2_fill_1 FILLER_58_592 ();
 sg13g2_fill_2 FILLER_58_603 ();
 sg13g2_fill_1 FILLER_58_619 ();
 sg13g2_fill_2 FILLER_58_655 ();
 sg13g2_fill_2 FILLER_58_737 ();
 sg13g2_fill_1 FILLER_58_743 ();
 sg13g2_fill_1 FILLER_58_748 ();
 sg13g2_fill_2 FILLER_58_755 ();
 sg13g2_fill_2 FILLER_58_763 ();
 sg13g2_fill_2 FILLER_58_775 ();
 sg13g2_fill_1 FILLER_58_777 ();
 sg13g2_decap_8 FILLER_58_781 ();
 sg13g2_decap_8 FILLER_58_788 ();
 sg13g2_decap_4 FILLER_58_795 ();
 sg13g2_fill_1 FILLER_58_824 ();
 sg13g2_fill_2 FILLER_58_833 ();
 sg13g2_fill_1 FILLER_58_840 ();
 sg13g2_fill_1 FILLER_58_886 ();
 sg13g2_fill_2 FILLER_58_900 ();
 sg13g2_fill_1 FILLER_58_956 ();
 sg13g2_fill_2 FILLER_58_968 ();
 sg13g2_fill_2 FILLER_58_1006 ();
 sg13g2_decap_8 FILLER_58_1018 ();
 sg13g2_decap_8 FILLER_58_1025 ();
 sg13g2_decap_4 FILLER_58_1061 ();
 sg13g2_fill_1 FILLER_58_1065 ();
 sg13g2_fill_2 FILLER_58_1102 ();
 sg13g2_fill_1 FILLER_58_1104 ();
 sg13g2_fill_1 FILLER_58_1126 ();
 sg13g2_decap_4 FILLER_58_1157 ();
 sg13g2_decap_4 FILLER_58_1166 ();
 sg13g2_fill_1 FILLER_58_1200 ();
 sg13g2_fill_1 FILLER_58_1211 ();
 sg13g2_fill_1 FILLER_58_1220 ();
 sg13g2_fill_1 FILLER_58_1231 ();
 sg13g2_fill_2 FILLER_58_1247 ();
 sg13g2_decap_4 FILLER_58_1278 ();
 sg13g2_fill_2 FILLER_58_1282 ();
 sg13g2_decap_8 FILLER_58_1289 ();
 sg13g2_decap_8 FILLER_58_1296 ();
 sg13g2_decap_8 FILLER_58_1303 ();
 sg13g2_decap_8 FILLER_58_1310 ();
 sg13g2_fill_2 FILLER_58_1317 ();
 sg13g2_fill_2 FILLER_58_1339 ();
 sg13g2_fill_1 FILLER_58_1377 ();
 sg13g2_fill_2 FILLER_58_1422 ();
 sg13g2_fill_2 FILLER_58_1429 ();
 sg13g2_decap_8 FILLER_58_1467 ();
 sg13g2_fill_2 FILLER_58_1474 ();
 sg13g2_fill_1 FILLER_58_1476 ();
 sg13g2_fill_1 FILLER_58_1539 ();
 sg13g2_fill_1 FILLER_58_1550 ();
 sg13g2_fill_2 FILLER_58_1557 ();
 sg13g2_decap_8 FILLER_58_1569 ();
 sg13g2_decap_8 FILLER_58_1576 ();
 sg13g2_fill_2 FILLER_58_1583 ();
 sg13g2_fill_1 FILLER_58_1585 ();
 sg13g2_decap_8 FILLER_58_1669 ();
 sg13g2_fill_1 FILLER_58_1676 ();
 sg13g2_decap_8 FILLER_58_1685 ();
 sg13g2_fill_2 FILLER_58_1692 ();
 sg13g2_fill_1 FILLER_58_1694 ();
 sg13g2_fill_1 FILLER_58_1705 ();
 sg13g2_decap_8 FILLER_58_1732 ();
 sg13g2_fill_2 FILLER_58_1739 ();
 sg13g2_decap_8 FILLER_58_1767 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_47 ();
 sg13g2_fill_2 FILLER_59_51 ();
 sg13g2_decap_4 FILLER_59_63 ();
 sg13g2_fill_1 FILLER_59_67 ();
 sg13g2_fill_2 FILLER_59_102 ();
 sg13g2_fill_1 FILLER_59_114 ();
 sg13g2_fill_1 FILLER_59_125 ();
 sg13g2_fill_1 FILLER_59_132 ();
 sg13g2_decap_4 FILLER_59_137 ();
 sg13g2_fill_1 FILLER_59_177 ();
 sg13g2_fill_2 FILLER_59_218 ();
 sg13g2_decap_8 FILLER_59_244 ();
 sg13g2_decap_8 FILLER_59_251 ();
 sg13g2_fill_2 FILLER_59_258 ();
 sg13g2_fill_1 FILLER_59_260 ();
 sg13g2_decap_8 FILLER_59_269 ();
 sg13g2_decap_8 FILLER_59_276 ();
 sg13g2_decap_8 FILLER_59_283 ();
 sg13g2_fill_2 FILLER_59_290 ();
 sg13g2_fill_2 FILLER_59_302 ();
 sg13g2_fill_1 FILLER_59_304 ();
 sg13g2_fill_1 FILLER_59_310 ();
 sg13g2_decap_4 FILLER_59_319 ();
 sg13g2_fill_1 FILLER_59_323 ();
 sg13g2_fill_1 FILLER_59_342 ();
 sg13g2_decap_8 FILLER_59_378 ();
 sg13g2_decap_4 FILLER_59_385 ();
 sg13g2_decap_4 FILLER_59_411 ();
 sg13g2_fill_1 FILLER_59_415 ();
 sg13g2_decap_4 FILLER_59_421 ();
 sg13g2_fill_1 FILLER_59_425 ();
 sg13g2_fill_2 FILLER_59_462 ();
 sg13g2_fill_1 FILLER_59_464 ();
 sg13g2_fill_2 FILLER_59_491 ();
 sg13g2_fill_2 FILLER_59_508 ();
 sg13g2_fill_1 FILLER_59_568 ();
 sg13g2_fill_2 FILLER_59_574 ();
 sg13g2_fill_1 FILLER_59_576 ();
 sg13g2_fill_1 FILLER_59_589 ();
 sg13g2_fill_1 FILLER_59_629 ();
 sg13g2_fill_1 FILLER_59_674 ();
 sg13g2_fill_1 FILLER_59_703 ();
 sg13g2_fill_2 FILLER_59_736 ();
 sg13g2_fill_1 FILLER_59_746 ();
 sg13g2_decap_4 FILLER_59_777 ();
 sg13g2_fill_2 FILLER_59_781 ();
 sg13g2_decap_8 FILLER_59_796 ();
 sg13g2_decap_4 FILLER_59_803 ();
 sg13g2_fill_1 FILLER_59_811 ();
 sg13g2_fill_2 FILLER_59_845 ();
 sg13g2_fill_2 FILLER_59_902 ();
 sg13g2_fill_1 FILLER_59_904 ();
 sg13g2_fill_1 FILLER_59_939 ();
 sg13g2_fill_2 FILLER_59_966 ();
 sg13g2_decap_8 FILLER_59_980 ();
 sg13g2_decap_4 FILLER_59_987 ();
 sg13g2_decap_4 FILLER_59_995 ();
 sg13g2_fill_1 FILLER_59_999 ();
 sg13g2_decap_8 FILLER_59_1008 ();
 sg13g2_decap_4 FILLER_59_1015 ();
 sg13g2_fill_1 FILLER_59_1019 ();
 sg13g2_decap_8 FILLER_59_1024 ();
 sg13g2_fill_1 FILLER_59_1031 ();
 sg13g2_fill_1 FILLER_59_1083 ();
 sg13g2_fill_2 FILLER_59_1088 ();
 sg13g2_decap_8 FILLER_59_1094 ();
 sg13g2_decap_4 FILLER_59_1101 ();
 sg13g2_fill_2 FILLER_59_1105 ();
 sg13g2_fill_2 FILLER_59_1156 ();
 sg13g2_fill_2 FILLER_59_1162 ();
 sg13g2_fill_1 FILLER_59_1164 ();
 sg13g2_fill_1 FILLER_59_1169 ();
 sg13g2_fill_2 FILLER_59_1196 ();
 sg13g2_fill_1 FILLER_59_1198 ();
 sg13g2_fill_2 FILLER_59_1208 ();
 sg13g2_fill_2 FILLER_59_1236 ();
 sg13g2_fill_1 FILLER_59_1238 ();
 sg13g2_decap_4 FILLER_59_1275 ();
 sg13g2_decap_4 FILLER_59_1319 ();
 sg13g2_fill_1 FILLER_59_1323 ();
 sg13g2_fill_2 FILLER_59_1355 ();
 sg13g2_fill_1 FILLER_59_1377 ();
 sg13g2_fill_1 FILLER_59_1382 ();
 sg13g2_fill_1 FILLER_59_1407 ();
 sg13g2_fill_2 FILLER_59_1424 ();
 sg13g2_fill_2 FILLER_59_1444 ();
 sg13g2_fill_1 FILLER_59_1446 ();
 sg13g2_decap_8 FILLER_59_1473 ();
 sg13g2_fill_1 FILLER_59_1480 ();
 sg13g2_decap_4 FILLER_59_1485 ();
 sg13g2_fill_1 FILLER_59_1489 ();
 sg13g2_fill_1 FILLER_59_1494 ();
 sg13g2_fill_2 FILLER_59_1516 ();
 sg13g2_fill_2 FILLER_59_1562 ();
 sg13g2_decap_8 FILLER_59_1572 ();
 sg13g2_decap_4 FILLER_59_1579 ();
 sg13g2_fill_1 FILLER_59_1587 ();
 sg13g2_decap_4 FILLER_59_1602 ();
 sg13g2_fill_2 FILLER_59_1606 ();
 sg13g2_decap_8 FILLER_59_1644 ();
 sg13g2_decap_8 FILLER_59_1651 ();
 sg13g2_decap_8 FILLER_59_1658 ();
 sg13g2_decap_8 FILLER_59_1665 ();
 sg13g2_fill_2 FILLER_59_1672 ();
 sg13g2_fill_1 FILLER_59_1674 ();
 sg13g2_decap_8 FILLER_59_1685 ();
 sg13g2_fill_2 FILLER_59_1692 ();
 sg13g2_decap_8 FILLER_59_1715 ();
 sg13g2_fill_2 FILLER_59_1722 ();
 sg13g2_fill_1 FILLER_59_1724 ();
 sg13g2_decap_8 FILLER_59_1761 ();
 sg13g2_decap_4 FILLER_59_1768 ();
 sg13g2_fill_2 FILLER_59_1772 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_2 FILLER_60_39 ();
 sg13g2_fill_1 FILLER_60_41 ();
 sg13g2_decap_8 FILLER_60_82 ();
 sg13g2_fill_1 FILLER_60_99 ();
 sg13g2_fill_2 FILLER_60_104 ();
 sg13g2_fill_1 FILLER_60_116 ();
 sg13g2_fill_1 FILLER_60_127 ();
 sg13g2_decap_4 FILLER_60_134 ();
 sg13g2_fill_1 FILLER_60_138 ();
 sg13g2_fill_1 FILLER_60_145 ();
 sg13g2_fill_1 FILLER_60_156 ();
 sg13g2_fill_2 FILLER_60_206 ();
 sg13g2_decap_8 FILLER_60_267 ();
 sg13g2_decap_8 FILLER_60_274 ();
 sg13g2_decap_4 FILLER_60_281 ();
 sg13g2_decap_8 FILLER_60_311 ();
 sg13g2_decap_4 FILLER_60_318 ();
 sg13g2_decap_8 FILLER_60_326 ();
 sg13g2_decap_4 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_337 ();
 sg13g2_fill_1 FILLER_60_364 ();
 sg13g2_fill_1 FILLER_60_446 ();
 sg13g2_fill_2 FILLER_60_491 ();
 sg13g2_fill_1 FILLER_60_592 ();
 sg13g2_fill_1 FILLER_60_665 ();
 sg13g2_decap_4 FILLER_60_675 ();
 sg13g2_decap_4 FILLER_60_686 ();
 sg13g2_fill_1 FILLER_60_716 ();
 sg13g2_fill_1 FILLER_60_750 ();
 sg13g2_fill_2 FILLER_60_787 ();
 sg13g2_fill_1 FILLER_60_789 ();
 sg13g2_fill_1 FILLER_60_799 ();
 sg13g2_fill_2 FILLER_60_860 ();
 sg13g2_fill_1 FILLER_60_862 ();
 sg13g2_decap_4 FILLER_60_901 ();
 sg13g2_fill_1 FILLER_60_905 ();
 sg13g2_fill_2 FILLER_60_927 ();
 sg13g2_fill_1 FILLER_60_959 ();
 sg13g2_fill_2 FILLER_60_996 ();
 sg13g2_fill_1 FILLER_60_998 ();
 sg13g2_fill_2 FILLER_60_1035 ();
 sg13g2_decap_4 FILLER_60_1047 ();
 sg13g2_fill_1 FILLER_60_1051 ();
 sg13g2_decap_8 FILLER_60_1056 ();
 sg13g2_fill_1 FILLER_60_1063 ();
 sg13g2_decap_8 FILLER_60_1068 ();
 sg13g2_fill_2 FILLER_60_1075 ();
 sg13g2_fill_1 FILLER_60_1077 ();
 sg13g2_fill_2 FILLER_60_1083 ();
 sg13g2_fill_1 FILLER_60_1085 ();
 sg13g2_decap_8 FILLER_60_1110 ();
 sg13g2_decap_4 FILLER_60_1117 ();
 sg13g2_fill_2 FILLER_60_1145 ();
 sg13g2_decap_8 FILLER_60_1151 ();
 sg13g2_decap_8 FILLER_60_1158 ();
 sg13g2_decap_4 FILLER_60_1165 ();
 sg13g2_fill_2 FILLER_60_1169 ();
 sg13g2_fill_2 FILLER_60_1224 ();
 sg13g2_fill_2 FILLER_60_1234 ();
 sg13g2_fill_1 FILLER_60_1236 ();
 sg13g2_fill_2 FILLER_60_1273 ();
 sg13g2_decap_4 FILLER_60_1311 ();
 sg13g2_decap_8 FILLER_60_1388 ();
 sg13g2_fill_1 FILLER_60_1405 ();
 sg13g2_fill_2 FILLER_60_1471 ();
 sg13g2_fill_1 FILLER_60_1473 ();
 sg13g2_decap_4 FILLER_60_1550 ();
 sg13g2_decap_4 FILLER_60_1619 ();
 sg13g2_fill_2 FILLER_60_1623 ();
 sg13g2_decap_4 FILLER_60_1656 ();
 sg13g2_fill_1 FILLER_60_1660 ();
 sg13g2_decap_4 FILLER_60_1708 ();
 sg13g2_fill_2 FILLER_60_1712 ();
 sg13g2_fill_2 FILLER_60_1738 ();
 sg13g2_fill_1 FILLER_60_1740 ();
 sg13g2_decap_8 FILLER_60_1767 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_fill_1 FILLER_61_49 ();
 sg13g2_fill_2 FILLER_61_76 ();
 sg13g2_fill_2 FILLER_61_104 ();
 sg13g2_fill_2 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_124 ();
 sg13g2_fill_2 FILLER_61_141 ();
 sg13g2_fill_2 FILLER_61_153 ();
 sg13g2_fill_1 FILLER_61_155 ();
 sg13g2_decap_8 FILLER_61_160 ();
 sg13g2_decap_4 FILLER_61_267 ();
 sg13g2_decap_8 FILLER_61_281 ();
 sg13g2_fill_1 FILLER_61_288 ();
 sg13g2_decap_8 FILLER_61_329 ();
 sg13g2_decap_4 FILLER_61_336 ();
 sg13g2_fill_1 FILLER_61_340 ();
 sg13g2_decap_4 FILLER_61_377 ();
 sg13g2_decap_4 FILLER_61_395 ();
 sg13g2_fill_2 FILLER_61_399 ();
 sg13g2_decap_8 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_61_422 ();
 sg13g2_decap_4 FILLER_61_433 ();
 sg13g2_fill_1 FILLER_61_437 ();
 sg13g2_decap_8 FILLER_61_442 ();
 sg13g2_decap_8 FILLER_61_449 ();
 sg13g2_fill_1 FILLER_61_456 ();
 sg13g2_fill_2 FILLER_61_488 ();
 sg13g2_fill_2 FILLER_61_500 ();
 sg13g2_fill_1 FILLER_61_516 ();
 sg13g2_fill_1 FILLER_61_520 ();
 sg13g2_fill_2 FILLER_61_526 ();
 sg13g2_fill_1 FILLER_61_632 ();
 sg13g2_fill_1 FILLER_61_662 ();
 sg13g2_fill_1 FILLER_61_699 ();
 sg13g2_fill_2 FILLER_61_710 ();
 sg13g2_fill_1 FILLER_61_730 ();
 sg13g2_decap_4 FILLER_61_787 ();
 sg13g2_fill_1 FILLER_61_886 ();
 sg13g2_fill_1 FILLER_61_911 ();
 sg13g2_fill_1 FILLER_61_916 ();
 sg13g2_fill_1 FILLER_61_921 ();
 sg13g2_fill_1 FILLER_61_932 ();
 sg13g2_fill_1 FILLER_61_943 ();
 sg13g2_decap_8 FILLER_61_948 ();
 sg13g2_decap_4 FILLER_61_955 ();
 sg13g2_fill_2 FILLER_61_959 ();
 sg13g2_decap_4 FILLER_61_996 ();
 sg13g2_fill_1 FILLER_61_1000 ();
 sg13g2_decap_8 FILLER_61_1026 ();
 sg13g2_decap_8 FILLER_61_1033 ();
 sg13g2_decap_4 FILLER_61_1040 ();
 sg13g2_fill_2 FILLER_61_1044 ();
 sg13g2_decap_4 FILLER_61_1072 ();
 sg13g2_fill_1 FILLER_61_1076 ();
 sg13g2_decap_8 FILLER_61_1081 ();
 sg13g2_decap_8 FILLER_61_1088 ();
 sg13g2_decap_8 FILLER_61_1095 ();
 sg13g2_decap_4 FILLER_61_1102 ();
 sg13g2_fill_1 FILLER_61_1106 ();
 sg13g2_decap_4 FILLER_61_1112 ();
 sg13g2_fill_1 FILLER_61_1116 ();
 sg13g2_decap_8 FILLER_61_1143 ();
 sg13g2_fill_2 FILLER_61_1150 ();
 sg13g2_fill_2 FILLER_61_1165 ();
 sg13g2_fill_1 FILLER_61_1167 ();
 sg13g2_fill_2 FILLER_61_1188 ();
 sg13g2_fill_1 FILLER_61_1190 ();
 sg13g2_fill_1 FILLER_61_1227 ();
 sg13g2_fill_1 FILLER_61_1299 ();
 sg13g2_decap_8 FILLER_61_1304 ();
 sg13g2_decap_4 FILLER_61_1311 ();
 sg13g2_fill_1 FILLER_61_1315 ();
 sg13g2_fill_2 FILLER_61_1347 ();
 sg13g2_fill_1 FILLER_61_1349 ();
 sg13g2_decap_4 FILLER_61_1354 ();
 sg13g2_fill_1 FILLER_61_1358 ();
 sg13g2_decap_8 FILLER_61_1363 ();
 sg13g2_decap_8 FILLER_61_1379 ();
 sg13g2_fill_1 FILLER_61_1386 ();
 sg13g2_fill_1 FILLER_61_1397 ();
 sg13g2_fill_2 FILLER_61_1408 ();
 sg13g2_decap_8 FILLER_61_1439 ();
 sg13g2_decap_8 FILLER_61_1446 ();
 sg13g2_fill_2 FILLER_61_1453 ();
 sg13g2_decap_8 FILLER_61_1463 ();
 sg13g2_decap_4 FILLER_61_1470 ();
 sg13g2_decap_8 FILLER_61_1486 ();
 sg13g2_fill_2 FILLER_61_1493 ();
 sg13g2_fill_1 FILLER_61_1495 ();
 sg13g2_fill_1 FILLER_61_1506 ();
 sg13g2_fill_2 FILLER_61_1517 ();
 sg13g2_fill_1 FILLER_61_1529 ();
 sg13g2_decap_4 FILLER_61_1540 ();
 sg13g2_decap_4 FILLER_61_1549 ();
 sg13g2_fill_2 FILLER_61_1614 ();
 sg13g2_decap_8 FILLER_61_1624 ();
 sg13g2_decap_8 FILLER_61_1631 ();
 sg13g2_fill_1 FILLER_61_1638 ();
 sg13g2_fill_2 FILLER_61_1649 ();
 sg13g2_fill_1 FILLER_61_1651 ();
 sg13g2_fill_2 FILLER_61_1656 ();
 sg13g2_fill_1 FILLER_61_1658 ();
 sg13g2_fill_2 FILLER_61_1689 ();
 sg13g2_decap_8 FILLER_61_1767 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_65 ();
 sg13g2_fill_2 FILLER_62_72 ();
 sg13g2_fill_1 FILLER_62_84 ();
 sg13g2_fill_2 FILLER_62_89 ();
 sg13g2_decap_8 FILLER_62_117 ();
 sg13g2_decap_4 FILLER_62_124 ();
 sg13g2_fill_2 FILLER_62_128 ();
 sg13g2_decap_8 FILLER_62_134 ();
 sg13g2_decap_8 FILLER_62_141 ();
 sg13g2_fill_1 FILLER_62_148 ();
 sg13g2_fill_2 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_207 ();
 sg13g2_decap_8 FILLER_62_214 ();
 sg13g2_decap_4 FILLER_62_221 ();
 sg13g2_decap_8 FILLER_62_262 ();
 sg13g2_decap_4 FILLER_62_269 ();
 sg13g2_fill_2 FILLER_62_273 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_fill_2 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_314 ();
 sg13g2_decap_8 FILLER_62_321 ();
 sg13g2_decap_8 FILLER_62_328 ();
 sg13g2_decap_8 FILLER_62_335 ();
 sg13g2_fill_2 FILLER_62_342 ();
 sg13g2_fill_1 FILLER_62_344 ();
 sg13g2_decap_8 FILLER_62_353 ();
 sg13g2_decap_4 FILLER_62_360 ();
 sg13g2_fill_1 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_417 ();
 sg13g2_decap_8 FILLER_62_424 ();
 sg13g2_decap_4 FILLER_62_431 ();
 sg13g2_fill_1 FILLER_62_435 ();
 sg13g2_decap_4 FILLER_62_469 ();
 sg13g2_fill_2 FILLER_62_473 ();
 sg13g2_fill_2 FILLER_62_479 ();
 sg13g2_fill_1 FILLER_62_498 ();
 sg13g2_fill_1 FILLER_62_511 ();
 sg13g2_fill_1 FILLER_62_524 ();
 sg13g2_decap_4 FILLER_62_574 ();
 sg13g2_fill_2 FILLER_62_578 ();
 sg13g2_fill_1 FILLER_62_599 ();
 sg13g2_fill_2 FILLER_62_622 ();
 sg13g2_fill_1 FILLER_62_688 ();
 sg13g2_fill_2 FILLER_62_693 ();
 sg13g2_fill_1 FILLER_62_705 ();
 sg13g2_fill_1 FILLER_62_735 ();
 sg13g2_fill_2 FILLER_62_754 ();
 sg13g2_fill_2 FILLER_62_773 ();
 sg13g2_fill_1 FILLER_62_784 ();
 sg13g2_fill_1 FILLER_62_815 ();
 sg13g2_fill_2 FILLER_62_836 ();
 sg13g2_fill_1 FILLER_62_846 ();
 sg13g2_fill_1 FILLER_62_851 ();
 sg13g2_fill_1 FILLER_62_888 ();
 sg13g2_fill_1 FILLER_62_915 ();
 sg13g2_decap_8 FILLER_62_942 ();
 sg13g2_decap_8 FILLER_62_949 ();
 sg13g2_decap_8 FILLER_62_956 ();
 sg13g2_fill_2 FILLER_62_963 ();
 sg13g2_fill_1 FILLER_62_965 ();
 sg13g2_fill_1 FILLER_62_987 ();
 sg13g2_fill_1 FILLER_62_997 ();
 sg13g2_decap_8 FILLER_62_1008 ();
 sg13g2_fill_2 FILLER_62_1041 ();
 sg13g2_fill_1 FILLER_62_1043 ();
 sg13g2_decap_8 FILLER_62_1054 ();
 sg13g2_decap_8 FILLER_62_1140 ();
 sg13g2_decap_8 FILLER_62_1147 ();
 sg13g2_decap_8 FILLER_62_1154 ();
 sg13g2_fill_2 FILLER_62_1161 ();
 sg13g2_decap_8 FILLER_62_1189 ();
 sg13g2_fill_2 FILLER_62_1196 ();
 sg13g2_fill_1 FILLER_62_1198 ();
 sg13g2_decap_8 FILLER_62_1225 ();
 sg13g2_decap_8 FILLER_62_1232 ();
 sg13g2_decap_4 FILLER_62_1239 ();
 sg13g2_fill_1 FILLER_62_1243 ();
 sg13g2_decap_8 FILLER_62_1270 ();
 sg13g2_fill_2 FILLER_62_1277 ();
 sg13g2_fill_1 FILLER_62_1279 ();
 sg13g2_fill_2 FILLER_62_1316 ();
 sg13g2_fill_2 FILLER_62_1321 ();
 sg13g2_fill_1 FILLER_62_1323 ();
 sg13g2_fill_1 FILLER_62_1328 ();
 sg13g2_fill_2 FILLER_62_1332 ();
 sg13g2_decap_8 FILLER_62_1347 ();
 sg13g2_decap_4 FILLER_62_1354 ();
 sg13g2_fill_1 FILLER_62_1358 ();
 sg13g2_fill_1 FILLER_62_1425 ();
 sg13g2_decap_4 FILLER_62_1430 ();
 sg13g2_fill_2 FILLER_62_1434 ();
 sg13g2_decap_4 FILLER_62_1441 ();
 sg13g2_fill_2 FILLER_62_1445 ();
 sg13g2_fill_2 FILLER_62_1450 ();
 sg13g2_fill_1 FILLER_62_1452 ();
 sg13g2_fill_2 FILLER_62_1468 ();
 sg13g2_decap_8 FILLER_62_1518 ();
 sg13g2_decap_4 FILLER_62_1525 ();
 sg13g2_fill_2 FILLER_62_1529 ();
 sg13g2_fill_2 FILLER_62_1543 ();
 sg13g2_fill_1 FILLER_62_1545 ();
 sg13g2_decap_4 FILLER_62_1568 ();
 sg13g2_decap_8 FILLER_62_1576 ();
 sg13g2_decap_8 FILLER_62_1583 ();
 sg13g2_decap_8 FILLER_62_1590 ();
 sg13g2_fill_2 FILLER_62_1597 ();
 sg13g2_fill_1 FILLER_62_1599 ();
 sg13g2_fill_2 FILLER_62_1640 ();
 sg13g2_fill_1 FILLER_62_1642 ();
 sg13g2_decap_4 FILLER_62_1709 ();
 sg13g2_fill_1 FILLER_62_1713 ();
 sg13g2_decap_4 FILLER_62_1769 ();
 sg13g2_fill_1 FILLER_62_1773 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_4 ();
 sg13g2_decap_4 FILLER_63_15 ();
 sg13g2_decap_8 FILLER_63_53 ();
 sg13g2_decap_8 FILLER_63_64 ();
 sg13g2_decap_8 FILLER_63_71 ();
 sg13g2_decap_8 FILLER_63_78 ();
 sg13g2_decap_8 FILLER_63_85 ();
 sg13g2_decap_4 FILLER_63_106 ();
 sg13g2_fill_1 FILLER_63_110 ();
 sg13g2_fill_2 FILLER_63_125 ();
 sg13g2_decap_4 FILLER_63_153 ();
 sg13g2_fill_1 FILLER_63_157 ();
 sg13g2_decap_8 FILLER_63_162 ();
 sg13g2_decap_8 FILLER_63_169 ();
 sg13g2_fill_2 FILLER_63_186 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_4 FILLER_63_210 ();
 sg13g2_fill_2 FILLER_63_214 ();
 sg13g2_decap_8 FILLER_63_244 ();
 sg13g2_decap_8 FILLER_63_251 ();
 sg13g2_decap_8 FILLER_63_258 ();
 sg13g2_decap_8 FILLER_63_265 ();
 sg13g2_decap_8 FILLER_63_272 ();
 sg13g2_fill_1 FILLER_63_279 ();
 sg13g2_decap_8 FILLER_63_284 ();
 sg13g2_decap_8 FILLER_63_291 ();
 sg13g2_decap_8 FILLER_63_298 ();
 sg13g2_decap_8 FILLER_63_305 ();
 sg13g2_fill_2 FILLER_63_312 ();
 sg13g2_decap_8 FILLER_63_324 ();
 sg13g2_fill_1 FILLER_63_345 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_fill_1 FILLER_63_387 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_fill_1 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_63_408 ();
 sg13g2_decap_4 FILLER_63_415 ();
 sg13g2_fill_1 FILLER_63_419 ();
 sg13g2_fill_2 FILLER_63_424 ();
 sg13g2_decap_8 FILLER_63_434 ();
 sg13g2_fill_1 FILLER_63_441 ();
 sg13g2_fill_2 FILLER_63_453 ();
 sg13g2_fill_1 FILLER_63_455 ();
 sg13g2_fill_1 FILLER_63_460 ();
 sg13g2_decap_4 FILLER_63_466 ();
 sg13g2_fill_1 FILLER_63_470 ();
 sg13g2_fill_2 FILLER_63_487 ();
 sg13g2_fill_1 FILLER_63_506 ();
 sg13g2_fill_1 FILLER_63_526 ();
 sg13g2_decap_4 FILLER_63_544 ();
 sg13g2_fill_2 FILLER_63_548 ();
 sg13g2_fill_1 FILLER_63_600 ();
 sg13g2_fill_2 FILLER_63_605 ();
 sg13g2_fill_2 FILLER_63_633 ();
 sg13g2_fill_1 FILLER_63_639 ();
 sg13g2_decap_8 FILLER_63_686 ();
 sg13g2_decap_8 FILLER_63_693 ();
 sg13g2_decap_4 FILLER_63_700 ();
 sg13g2_fill_2 FILLER_63_721 ();
 sg13g2_fill_2 FILLER_63_735 ();
 sg13g2_decap_8 FILLER_63_768 ();
 sg13g2_decap_8 FILLER_63_775 ();
 sg13g2_decap_8 FILLER_63_782 ();
 sg13g2_decap_4 FILLER_63_789 ();
 sg13g2_decap_8 FILLER_63_852 ();
 sg13g2_fill_2 FILLER_63_867 ();
 sg13g2_fill_1 FILLER_63_869 ();
 sg13g2_decap_4 FILLER_63_878 ();
 sg13g2_fill_2 FILLER_63_882 ();
 sg13g2_decap_4 FILLER_63_894 ();
 sg13g2_fill_2 FILLER_63_902 ();
 sg13g2_fill_1 FILLER_63_904 ();
 sg13g2_fill_1 FILLER_63_926 ();
 sg13g2_fill_1 FILLER_63_931 ();
 sg13g2_fill_1 FILLER_63_942 ();
 sg13g2_fill_1 FILLER_63_953 ();
 sg13g2_decap_8 FILLER_63_958 ();
 sg13g2_decap_8 FILLER_63_965 ();
 sg13g2_fill_2 FILLER_63_985 ();
 sg13g2_decap_4 FILLER_63_1016 ();
 sg13g2_fill_1 FILLER_63_1020 ();
 sg13g2_fill_2 FILLER_63_1051 ();
 sg13g2_decap_4 FILLER_63_1133 ();
 sg13g2_decap_8 FILLER_63_1145 ();
 sg13g2_decap_8 FILLER_63_1152 ();
 sg13g2_decap_8 FILLER_63_1159 ();
 sg13g2_fill_2 FILLER_63_1166 ();
 sg13g2_fill_1 FILLER_63_1168 ();
 sg13g2_decap_8 FILLER_63_1199 ();
 sg13g2_decap_8 FILLER_63_1215 ();
 sg13g2_fill_2 FILLER_63_1222 ();
 sg13g2_fill_1 FILLER_63_1224 ();
 sg13g2_decap_8 FILLER_63_1229 ();
 sg13g2_decap_8 FILLER_63_1236 ();
 sg13g2_decap_4 FILLER_63_1243 ();
 sg13g2_fill_1 FILLER_63_1247 ();
 sg13g2_fill_2 FILLER_63_1262 ();
 sg13g2_fill_1 FILLER_63_1264 ();
 sg13g2_decap_4 FILLER_63_1303 ();
 sg13g2_fill_2 FILLER_63_1307 ();
 sg13g2_fill_2 FILLER_63_1340 ();
 sg13g2_decap_8 FILLER_63_1355 ();
 sg13g2_decap_8 FILLER_63_1362 ();
 sg13g2_decap_4 FILLER_63_1369 ();
 sg13g2_fill_2 FILLER_63_1373 ();
 sg13g2_decap_4 FILLER_63_1379 ();
 sg13g2_decap_4 FILLER_63_1408 ();
 sg13g2_fill_1 FILLER_63_1412 ();
 sg13g2_fill_2 FILLER_63_1445 ();
 sg13g2_decap_4 FILLER_63_1485 ();
 sg13g2_fill_1 FILLER_63_1489 ();
 sg13g2_fill_1 FILLER_63_1500 ();
 sg13g2_fill_2 FILLER_63_1537 ();
 sg13g2_decap_8 FILLER_63_1591 ();
 sg13g2_decap_4 FILLER_63_1598 ();
 sg13g2_fill_2 FILLER_63_1602 ();
 sg13g2_decap_4 FILLER_63_1612 ();
 sg13g2_decap_8 FILLER_63_1646 ();
 sg13g2_decap_8 FILLER_63_1653 ();
 sg13g2_fill_2 FILLER_63_1660 ();
 sg13g2_decap_8 FILLER_63_1672 ();
 sg13g2_fill_2 FILLER_63_1679 ();
 sg13g2_fill_1 FILLER_63_1681 ();
 sg13g2_fill_1 FILLER_63_1686 ();
 sg13g2_fill_1 FILLER_63_1721 ();
 sg13g2_decap_4 FILLER_63_1742 ();
 sg13g2_fill_2 FILLER_63_1746 ();
 sg13g2_decap_8 FILLER_63_1752 ();
 sg13g2_decap_8 FILLER_63_1759 ();
 sg13g2_decap_8 FILLER_63_1766 ();
 sg13g2_fill_1 FILLER_63_1773 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_fill_1 FILLER_64_35 ();
 sg13g2_decap_4 FILLER_64_46 ();
 sg13g2_fill_2 FILLER_64_50 ();
 sg13g2_decap_8 FILLER_64_78 ();
 sg13g2_fill_2 FILLER_64_85 ();
 sg13g2_fill_1 FILLER_64_87 ();
 sg13g2_decap_8 FILLER_64_96 ();
 sg13g2_decap_8 FILLER_64_103 ();
 sg13g2_decap_8 FILLER_64_110 ();
 sg13g2_decap_4 FILLER_64_121 ();
 sg13g2_fill_1 FILLER_64_125 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_198 ();
 sg13g2_decap_8 FILLER_64_205 ();
 sg13g2_decap_4 FILLER_64_212 ();
 sg13g2_decap_4 FILLER_64_252 ();
 sg13g2_fill_2 FILLER_64_256 ();
 sg13g2_decap_8 FILLER_64_261 ();
 sg13g2_decap_8 FILLER_64_268 ();
 sg13g2_fill_2 FILLER_64_275 ();
 sg13g2_fill_1 FILLER_64_315 ();
 sg13g2_decap_4 FILLER_64_326 ();
 sg13g2_fill_2 FILLER_64_330 ();
 sg13g2_fill_1 FILLER_64_338 ();
 sg13g2_decap_4 FILLER_64_343 ();
 sg13g2_fill_1 FILLER_64_347 ();
 sg13g2_decap_4 FILLER_64_353 ();
 sg13g2_decap_8 FILLER_64_363 ();
 sg13g2_decap_8 FILLER_64_370 ();
 sg13g2_decap_8 FILLER_64_377 ();
 sg13g2_decap_8 FILLER_64_384 ();
 sg13g2_decap_8 FILLER_64_391 ();
 sg13g2_decap_8 FILLER_64_398 ();
 sg13g2_fill_2 FILLER_64_405 ();
 sg13g2_fill_1 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_64_414 ();
 sg13g2_decap_8 FILLER_64_421 ();
 sg13g2_decap_8 FILLER_64_428 ();
 sg13g2_decap_4 FILLER_64_435 ();
 sg13g2_fill_2 FILLER_64_439 ();
 sg13g2_fill_2 FILLER_64_518 ();
 sg13g2_fill_1 FILLER_64_570 ();
 sg13g2_decap_8 FILLER_64_628 ();
 sg13g2_fill_2 FILLER_64_635 ();
 sg13g2_fill_1 FILLER_64_637 ();
 sg13g2_decap_4 FILLER_64_646 ();
 sg13g2_fill_1 FILLER_64_650 ();
 sg13g2_fill_1 FILLER_64_665 ();
 sg13g2_fill_1 FILLER_64_725 ();
 sg13g2_decap_8 FILLER_64_780 ();
 sg13g2_decap_8 FILLER_64_787 ();
 sg13g2_decap_4 FILLER_64_794 ();
 sg13g2_fill_2 FILLER_64_798 ();
 sg13g2_decap_8 FILLER_64_862 ();
 sg13g2_fill_1 FILLER_64_869 ();
 sg13g2_fill_2 FILLER_64_945 ();
 sg13g2_fill_2 FILLER_64_973 ();
 sg13g2_fill_1 FILLER_64_1078 ();
 sg13g2_fill_2 FILLER_64_1122 ();
 sg13g2_decap_8 FILLER_64_1146 ();
 sg13g2_decap_8 FILLER_64_1153 ();
 sg13g2_decap_8 FILLER_64_1160 ();
 sg13g2_decap_8 FILLER_64_1167 ();
 sg13g2_fill_2 FILLER_64_1174 ();
 sg13g2_decap_8 FILLER_64_1235 ();
 sg13g2_decap_4 FILLER_64_1242 ();
 sg13g2_decap_8 FILLER_64_1292 ();
 sg13g2_fill_1 FILLER_64_1299 ();
 sg13g2_decap_4 FILLER_64_1304 ();
 sg13g2_fill_1 FILLER_64_1308 ();
 sg13g2_decap_8 FILLER_64_1362 ();
 sg13g2_fill_2 FILLER_64_1369 ();
 sg13g2_decap_4 FILLER_64_1397 ();
 sg13g2_fill_2 FILLER_64_1437 ();
 sg13g2_fill_1 FILLER_64_1455 ();
 sg13g2_fill_1 FILLER_64_1469 ();
 sg13g2_decap_8 FILLER_64_1493 ();
 sg13g2_fill_2 FILLER_64_1500 ();
 sg13g2_fill_1 FILLER_64_1502 ();
 sg13g2_fill_2 FILLER_64_1529 ();
 sg13g2_decap_4 FILLER_64_1557 ();
 sg13g2_fill_1 FILLER_64_1561 ();
 sg13g2_fill_1 FILLER_64_1608 ();
 sg13g2_decap_8 FILLER_64_1644 ();
 sg13g2_decap_4 FILLER_64_1651 ();
 sg13g2_fill_1 FILLER_64_1655 ();
 sg13g2_decap_8 FILLER_64_1692 ();
 sg13g2_decap_4 FILLER_64_1699 ();
 sg13g2_decap_8 FILLER_64_1729 ();
 sg13g2_fill_1 FILLER_64_1736 ();
 sg13g2_decap_8 FILLER_64_1767 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_fill_2 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_37 ();
 sg13g2_fill_2 FILLER_65_48 ();
 sg13g2_fill_1 FILLER_65_50 ();
 sg13g2_decap_8 FILLER_65_61 ();
 sg13g2_decap_8 FILLER_65_68 ();
 sg13g2_fill_1 FILLER_65_85 ();
 sg13g2_fill_2 FILLER_65_96 ();
 sg13g2_decap_8 FILLER_65_160 ();
 sg13g2_decap_4 FILLER_65_203 ();
 sg13g2_fill_1 FILLER_65_207 ();
 sg13g2_decap_8 FILLER_65_267 ();
 sg13g2_decap_8 FILLER_65_274 ();
 sg13g2_decap_8 FILLER_65_281 ();
 sg13g2_fill_1 FILLER_65_288 ();
 sg13g2_fill_1 FILLER_65_329 ();
 sg13g2_fill_1 FILLER_65_336 ();
 sg13g2_fill_2 FILLER_65_347 ();
 sg13g2_decap_4 FILLER_65_359 ();
 sg13g2_decap_4 FILLER_65_373 ();
 sg13g2_fill_1 FILLER_65_383 ();
 sg13g2_fill_1 FILLER_65_394 ();
 sg13g2_fill_2 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_413 ();
 sg13g2_fill_2 FILLER_65_440 ();
 sg13g2_decap_4 FILLER_65_446 ();
 sg13g2_fill_2 FILLER_65_455 ();
 sg13g2_fill_1 FILLER_65_462 ();
 sg13g2_decap_8 FILLER_65_469 ();
 sg13g2_decap_4 FILLER_65_476 ();
 sg13g2_fill_2 FILLER_65_480 ();
 sg13g2_fill_1 FILLER_65_509 ();
 sg13g2_fill_1 FILLER_65_541 ();
 sg13g2_decap_4 FILLER_65_547 ();
 sg13g2_fill_2 FILLER_65_551 ();
 sg13g2_fill_1 FILLER_65_579 ();
 sg13g2_fill_1 FILLER_65_618 ();
 sg13g2_decap_8 FILLER_65_637 ();
 sg13g2_decap_8 FILLER_65_644 ();
 sg13g2_decap_8 FILLER_65_656 ();
 sg13g2_decap_8 FILLER_65_663 ();
 sg13g2_decap_8 FILLER_65_670 ();
 sg13g2_decap_8 FILLER_65_677 ();
 sg13g2_fill_2 FILLER_65_684 ();
 sg13g2_fill_1 FILLER_65_686 ();
 sg13g2_decap_4 FILLER_65_691 ();
 sg13g2_fill_2 FILLER_65_695 ();
 sg13g2_fill_1 FILLER_65_721 ();
 sg13g2_fill_1 FILLER_65_748 ();
 sg13g2_fill_1 FILLER_65_753 ();
 sg13g2_decap_8 FILLER_65_768 ();
 sg13g2_decap_8 FILLER_65_775 ();
 sg13g2_decap_8 FILLER_65_782 ();
 sg13g2_decap_4 FILLER_65_789 ();
 sg13g2_fill_1 FILLER_65_803 ();
 sg13g2_decap_8 FILLER_65_858 ();
 sg13g2_decap_8 FILLER_65_865 ();
 sg13g2_fill_1 FILLER_65_872 ();
 sg13g2_decap_8 FILLER_65_908 ();
 sg13g2_decap_4 FILLER_65_915 ();
 sg13g2_fill_1 FILLER_65_919 ();
 sg13g2_fill_2 FILLER_65_925 ();
 sg13g2_fill_1 FILLER_65_927 ();
 sg13g2_fill_2 FILLER_65_932 ();
 sg13g2_fill_1 FILLER_65_934 ();
 sg13g2_fill_2 FILLER_65_990 ();
 sg13g2_fill_2 FILLER_65_1061 ();
 sg13g2_fill_2 FILLER_65_1067 ();
 sg13g2_fill_2 FILLER_65_1073 ();
 sg13g2_fill_1 FILLER_65_1096 ();
 sg13g2_fill_2 FILLER_65_1103 ();
 sg13g2_fill_1 FILLER_65_1115 ();
 sg13g2_fill_1 FILLER_65_1142 ();
 sg13g2_decap_8 FILLER_65_1148 ();
 sg13g2_decap_8 FILLER_65_1155 ();
 sg13g2_decap_4 FILLER_65_1162 ();
 sg13g2_fill_2 FILLER_65_1166 ();
 sg13g2_fill_1 FILLER_65_1194 ();
 sg13g2_fill_2 FILLER_65_1199 ();
 sg13g2_fill_2 FILLER_65_1211 ();
 sg13g2_fill_1 FILLER_65_1213 ();
 sg13g2_fill_1 FILLER_65_1224 ();
 sg13g2_fill_2 FILLER_65_1251 ();
 sg13g2_fill_2 FILLER_65_1263 ();
 sg13g2_fill_2 FILLER_65_1269 ();
 sg13g2_decap_8 FILLER_65_1275 ();
 sg13g2_fill_1 FILLER_65_1360 ();
 sg13g2_fill_2 FILLER_65_1391 ();
 sg13g2_fill_1 FILLER_65_1482 ();
 sg13g2_decap_8 FILLER_65_1513 ();
 sg13g2_decap_4 FILLER_65_1520 ();
 sg13g2_fill_1 FILLER_65_1524 ();
 sg13g2_fill_2 FILLER_65_1543 ();
 sg13g2_decap_4 FILLER_65_1549 ();
 sg13g2_fill_1 FILLER_65_1553 ();
 sg13g2_decap_4 FILLER_65_1564 ();
 sg13g2_decap_8 FILLER_65_1614 ();
 sg13g2_fill_2 FILLER_65_1621 ();
 sg13g2_decap_8 FILLER_65_1649 ();
 sg13g2_decap_8 FILLER_65_1656 ();
 sg13g2_decap_8 FILLER_65_1663 ();
 sg13g2_decap_8 FILLER_65_1670 ();
 sg13g2_decap_8 FILLER_65_1677 ();
 sg13g2_decap_8 FILLER_65_1684 ();
 sg13g2_decap_8 FILLER_65_1691 ();
 sg13g2_decap_8 FILLER_65_1744 ();
 sg13g2_decap_8 FILLER_65_1751 ();
 sg13g2_decap_8 FILLER_65_1758 ();
 sg13g2_decap_8 FILLER_65_1765 ();
 sg13g2_fill_2 FILLER_65_1772 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_33 ();
 sg13g2_fill_1 FILLER_66_39 ();
 sg13g2_fill_1 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_81 ();
 sg13g2_fill_2 FILLER_66_143 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_189 ();
 sg13g2_fill_2 FILLER_66_196 ();
 sg13g2_fill_1 FILLER_66_198 ();
 sg13g2_decap_8 FILLER_66_218 ();
 sg13g2_fill_2 FILLER_66_225 ();
 sg13g2_fill_2 FILLER_66_230 ();
 sg13g2_decap_8 FILLER_66_274 ();
 sg13g2_fill_1 FILLER_66_281 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_fill_1 FILLER_66_333 ();
 sg13g2_fill_2 FILLER_66_415 ();
 sg13g2_fill_1 FILLER_66_453 ();
 sg13g2_fill_1 FILLER_66_463 ();
 sg13g2_fill_2 FILLER_66_474 ();
 sg13g2_fill_1 FILLER_66_476 ();
 sg13g2_decap_4 FILLER_66_610 ();
 sg13g2_fill_1 FILLER_66_614 ();
 sg13g2_fill_1 FILLER_66_624 ();
 sg13g2_decap_8 FILLER_66_666 ();
 sg13g2_decap_8 FILLER_66_673 ();
 sg13g2_decap_8 FILLER_66_680 ();
 sg13g2_decap_4 FILLER_66_687 ();
 sg13g2_fill_1 FILLER_66_691 ();
 sg13g2_fill_2 FILLER_66_732 ();
 sg13g2_decap_8 FILLER_66_768 ();
 sg13g2_decap_8 FILLER_66_775 ();
 sg13g2_decap_8 FILLER_66_782 ();
 sg13g2_fill_2 FILLER_66_789 ();
 sg13g2_decap_4 FILLER_66_838 ();
 sg13g2_fill_1 FILLER_66_842 ();
 sg13g2_decap_4 FILLER_66_852 ();
 sg13g2_fill_2 FILLER_66_856 ();
 sg13g2_fill_1 FILLER_66_868 ();
 sg13g2_decap_4 FILLER_66_915 ();
 sg13g2_fill_1 FILLER_66_919 ();
 sg13g2_fill_2 FILLER_66_930 ();
 sg13g2_fill_1 FILLER_66_932 ();
 sg13g2_decap_8 FILLER_66_959 ();
 sg13g2_decap_4 FILLER_66_966 ();
 sg13g2_fill_2 FILLER_66_984 ();
 sg13g2_decap_4 FILLER_66_997 ();
 sg13g2_decap_8 FILLER_66_1010 ();
 sg13g2_decap_4 FILLER_66_1017 ();
 sg13g2_fill_2 FILLER_66_1021 ();
 sg13g2_fill_2 FILLER_66_1062 ();
 sg13g2_decap_8 FILLER_66_1130 ();
 sg13g2_decap_8 FILLER_66_1137 ();
 sg13g2_decap_8 FILLER_66_1144 ();
 sg13g2_decap_4 FILLER_66_1151 ();
 sg13g2_fill_2 FILLER_66_1155 ();
 sg13g2_decap_8 FILLER_66_1161 ();
 sg13g2_decap_4 FILLER_66_1168 ();
 sg13g2_fill_2 FILLER_66_1172 ();
 sg13g2_decap_4 FILLER_66_1198 ();
 sg13g2_fill_1 FILLER_66_1202 ();
 sg13g2_decap_4 FILLER_66_1229 ();
 sg13g2_fill_1 FILLER_66_1233 ();
 sg13g2_decap_8 FILLER_66_1238 ();
 sg13g2_fill_2 FILLER_66_1245 ();
 sg13g2_fill_1 FILLER_66_1247 ();
 sg13g2_fill_1 FILLER_66_1282 ();
 sg13g2_fill_1 FILLER_66_1319 ();
 sg13g2_fill_1 FILLER_66_1330 ();
 sg13g2_fill_2 FILLER_66_1387 ();
 sg13g2_fill_1 FILLER_66_1389 ();
 sg13g2_fill_1 FILLER_66_1404 ();
 sg13g2_fill_2 FILLER_66_1457 ();
 sg13g2_fill_1 FILLER_66_1466 ();
 sg13g2_fill_2 FILLER_66_1475 ();
 sg13g2_fill_2 FILLER_66_1481 ();
 sg13g2_decap_8 FILLER_66_1497 ();
 sg13g2_decap_8 FILLER_66_1504 ();
 sg13g2_decap_4 FILLER_66_1511 ();
 sg13g2_fill_1 FILLER_66_1515 ();
 sg13g2_fill_1 FILLER_66_1589 ();
 sg13g2_fill_1 FILLER_66_1594 ();
 sg13g2_fill_2 FILLER_66_1615 ();
 sg13g2_fill_2 FILLER_66_1643 ();
 sg13g2_fill_2 FILLER_66_1671 ();
 sg13g2_fill_2 FILLER_66_1699 ();
 sg13g2_fill_1 FILLER_66_1701 ();
 sg13g2_fill_1 FILLER_66_1706 ();
 sg13g2_fill_2 FILLER_66_1733 ();
 sg13g2_fill_1 FILLER_66_1735 ();
 sg13g2_decap_8 FILLER_66_1766 ();
 sg13g2_fill_1 FILLER_66_1773 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_15 ();
 sg13g2_fill_1 FILLER_67_26 ();
 sg13g2_fill_1 FILLER_67_53 ();
 sg13g2_fill_1 FILLER_67_59 ();
 sg13g2_decap_8 FILLER_67_86 ();
 sg13g2_fill_2 FILLER_67_93 ();
 sg13g2_fill_2 FILLER_67_150 ();
 sg13g2_decap_8 FILLER_67_156 ();
 sg13g2_fill_2 FILLER_67_163 ();
 sg13g2_fill_1 FILLER_67_226 ();
 sg13g2_decap_8 FILLER_67_272 ();
 sg13g2_decap_4 FILLER_67_279 ();
 sg13g2_fill_2 FILLER_67_283 ();
 sg13g2_fill_2 FILLER_67_289 ();
 sg13g2_fill_1 FILLER_67_291 ();
 sg13g2_fill_2 FILLER_67_395 ();
 sg13g2_fill_2 FILLER_67_446 ();
 sg13g2_fill_1 FILLER_67_458 ();
 sg13g2_decap_8 FILLER_67_465 ();
 sg13g2_decap_4 FILLER_67_472 ();
 sg13g2_fill_1 FILLER_67_496 ();
 sg13g2_decap_8 FILLER_67_567 ();
 sg13g2_fill_1 FILLER_67_596 ();
 sg13g2_fill_2 FILLER_67_602 ();
 sg13g2_fill_2 FILLER_67_614 ();
 sg13g2_fill_2 FILLER_67_642 ();
 sg13g2_fill_2 FILLER_67_684 ();
 sg13g2_fill_1 FILLER_67_705 ();
 sg13g2_fill_1 FILLER_67_714 ();
 sg13g2_decap_8 FILLER_67_760 ();
 sg13g2_decap_4 FILLER_67_767 ();
 sg13g2_fill_1 FILLER_67_771 ();
 sg13g2_decap_4 FILLER_67_778 ();
 sg13g2_fill_2 FILLER_67_782 ();
 sg13g2_fill_1 FILLER_67_813 ();
 sg13g2_decap_4 FILLER_67_850 ();
 sg13g2_fill_2 FILLER_67_854 ();
 sg13g2_fill_2 FILLER_67_895 ();
 sg13g2_fill_1 FILLER_67_897 ();
 sg13g2_fill_2 FILLER_67_924 ();
 sg13g2_fill_1 FILLER_67_926 ();
 sg13g2_fill_2 FILLER_67_941 ();
 sg13g2_fill_1 FILLER_67_943 ();
 sg13g2_decap_8 FILLER_67_948 ();
 sg13g2_decap_8 FILLER_67_959 ();
 sg13g2_decap_8 FILLER_67_966 ();
 sg13g2_decap_8 FILLER_67_973 ();
 sg13g2_decap_4 FILLER_67_980 ();
 sg13g2_fill_2 FILLER_67_984 ();
 sg13g2_fill_1 FILLER_67_989 ();
 sg13g2_fill_2 FILLER_67_1000 ();
 sg13g2_decap_8 FILLER_67_1007 ();
 sg13g2_decap_8 FILLER_67_1014 ();
 sg13g2_decap_8 FILLER_67_1021 ();
 sg13g2_decap_4 FILLER_67_1028 ();
 sg13g2_fill_1 FILLER_67_1032 ();
 sg13g2_decap_8 FILLER_67_1059 ();
 sg13g2_decap_8 FILLER_67_1066 ();
 sg13g2_decap_4 FILLER_67_1133 ();
 sg13g2_decap_4 FILLER_67_1145 ();
 sg13g2_fill_1 FILLER_67_1149 ();
 sg13g2_fill_1 FILLER_67_1176 ();
 sg13g2_fill_1 FILLER_67_1183 ();
 sg13g2_fill_1 FILLER_67_1228 ();
 sg13g2_decap_4 FILLER_67_1255 ();
 sg13g2_decap_4 FILLER_67_1295 ();
 sg13g2_fill_1 FILLER_67_1299 ();
 sg13g2_fill_1 FILLER_67_1304 ();
 sg13g2_fill_1 FILLER_67_1330 ();
 sg13g2_fill_1 FILLER_67_1365 ();
 sg13g2_decap_8 FILLER_67_1422 ();
 sg13g2_fill_1 FILLER_67_1429 ();
 sg13g2_decap_8 FILLER_67_1438 ();
 sg13g2_fill_2 FILLER_67_1445 ();
 sg13g2_fill_1 FILLER_67_1447 ();
 sg13g2_decap_8 FILLER_67_1487 ();
 sg13g2_decap_8 FILLER_67_1494 ();
 sg13g2_decap_8 FILLER_67_1501 ();
 sg13g2_decap_8 FILLER_67_1508 ();
 sg13g2_decap_4 FILLER_67_1515 ();
 sg13g2_fill_1 FILLER_67_1519 ();
 sg13g2_decap_8 FILLER_67_1530 ();
 sg13g2_fill_2 FILLER_67_1537 ();
 sg13g2_decap_8 FILLER_67_1553 ();
 sg13g2_decap_8 FILLER_67_1560 ();
 sg13g2_decap_4 FILLER_67_1567 ();
 sg13g2_decap_8 FILLER_67_1575 ();
 sg13g2_fill_2 FILLER_67_1582 ();
 sg13g2_decap_8 FILLER_67_1588 ();
 sg13g2_decap_4 FILLER_67_1595 ();
 sg13g2_decap_4 FILLER_67_1633 ();
 sg13g2_fill_1 FILLER_67_1637 ();
 sg13g2_fill_1 FILLER_67_1664 ();
 sg13g2_fill_1 FILLER_67_1679 ();
 sg13g2_decap_8 FILLER_67_1684 ();
 sg13g2_decap_4 FILLER_67_1691 ();
 sg13g2_decap_8 FILLER_67_1718 ();
 sg13g2_decap_4 FILLER_67_1725 ();
 sg13g2_decap_4 FILLER_67_1769 ();
 sg13g2_fill_1 FILLER_67_1773 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_4 ();
 sg13g2_fill_1 FILLER_68_31 ();
 sg13g2_fill_2 FILLER_68_46 ();
 sg13g2_fill_2 FILLER_68_60 ();
 sg13g2_fill_1 FILLER_68_98 ();
 sg13g2_fill_2 FILLER_68_131 ();
 sg13g2_decap_8 FILLER_68_143 ();
 sg13g2_decap_8 FILLER_68_150 ();
 sg13g2_fill_2 FILLER_68_169 ();
 sg13g2_fill_1 FILLER_68_171 ();
 sg13g2_fill_1 FILLER_68_208 ();
 sg13g2_fill_2 FILLER_68_240 ();
 sg13g2_decap_4 FILLER_68_250 ();
 sg13g2_fill_1 FILLER_68_258 ();
 sg13g2_fill_2 FILLER_68_288 ();
 sg13g2_fill_1 FILLER_68_295 ();
 sg13g2_fill_1 FILLER_68_300 ();
 sg13g2_fill_2 FILLER_68_309 ();
 sg13g2_fill_1 FILLER_68_331 ();
 sg13g2_fill_1 FILLER_68_342 ();
 sg13g2_fill_1 FILLER_68_357 ();
 sg13g2_fill_1 FILLER_68_410 ();
 sg13g2_fill_1 FILLER_68_463 ();
 sg13g2_decap_8 FILLER_68_469 ();
 sg13g2_decap_8 FILLER_68_476 ();
 sg13g2_fill_2 FILLER_68_483 ();
 sg13g2_fill_2 FILLER_68_525 ();
 sg13g2_fill_1 FILLER_68_537 ();
 sg13g2_decap_8 FILLER_68_542 ();
 sg13g2_decap_4 FILLER_68_549 ();
 sg13g2_decap_8 FILLER_68_563 ();
 sg13g2_decap_4 FILLER_68_570 ();
 sg13g2_fill_2 FILLER_68_574 ();
 sg13g2_decap_4 FILLER_68_617 ();
 sg13g2_fill_2 FILLER_68_621 ();
 sg13g2_fill_1 FILLER_68_627 ();
 sg13g2_decap_4 FILLER_68_638 ();
 sg13g2_decap_4 FILLER_68_652 ();
 sg13g2_fill_1 FILLER_68_656 ();
 sg13g2_fill_2 FILLER_68_687 ();
 sg13g2_fill_2 FILLER_68_710 ();
 sg13g2_fill_1 FILLER_68_742 ();
 sg13g2_decap_4 FILLER_68_779 ();
 sg13g2_fill_2 FILLER_68_783 ();
 sg13g2_fill_2 FILLER_68_811 ();
 sg13g2_fill_1 FILLER_68_817 ();
 sg13g2_fill_1 FILLER_68_822 ();
 sg13g2_fill_1 FILLER_68_833 ();
 sg13g2_fill_2 FILLER_68_860 ();
 sg13g2_decap_8 FILLER_68_866 ();
 sg13g2_fill_2 FILLER_68_873 ();
 sg13g2_fill_1 FILLER_68_875 ();
 sg13g2_fill_1 FILLER_68_887 ();
 sg13g2_decap_8 FILLER_68_892 ();
 sg13g2_decap_4 FILLER_68_899 ();
 sg13g2_fill_1 FILLER_68_903 ();
 sg13g2_decap_4 FILLER_68_913 ();
 sg13g2_fill_2 FILLER_68_926 ();
 sg13g2_fill_1 FILLER_68_928 ();
 sg13g2_fill_1 FILLER_68_933 ();
 sg13g2_fill_1 FILLER_68_955 ();
 sg13g2_fill_1 FILLER_68_982 ();
 sg13g2_fill_2 FILLER_68_993 ();
 sg13g2_decap_4 FILLER_68_1021 ();
 sg13g2_decap_8 FILLER_68_1073 ();
 sg13g2_decap_4 FILLER_68_1080 ();
 sg13g2_fill_1 FILLER_68_1084 ();
 sg13g2_fill_2 FILLER_68_1089 ();
 sg13g2_decap_4 FILLER_68_1141 ();
 sg13g2_fill_2 FILLER_68_1145 ();
 sg13g2_fill_1 FILLER_68_1173 ();
 sg13g2_fill_1 FILLER_68_1184 ();
 sg13g2_fill_2 FILLER_68_1224 ();
 sg13g2_decap_4 FILLER_68_1230 ();
 sg13g2_fill_2 FILLER_68_1234 ();
 sg13g2_decap_8 FILLER_68_1240 ();
 sg13g2_decap_4 FILLER_68_1247 ();
 sg13g2_fill_2 FILLER_68_1251 ();
 sg13g2_decap_4 FILLER_68_1258 ();
 sg13g2_fill_1 FILLER_68_1262 ();
 sg13g2_decap_4 FILLER_68_1267 ();
 sg13g2_fill_1 FILLER_68_1271 ();
 sg13g2_fill_1 FILLER_68_1308 ();
 sg13g2_fill_1 FILLER_68_1364 ();
 sg13g2_decap_8 FILLER_68_1417 ();
 sg13g2_fill_2 FILLER_68_1424 ();
 sg13g2_decap_8 FILLER_68_1439 ();
 sg13g2_decap_4 FILLER_68_1446 ();
 sg13g2_fill_1 FILLER_68_1450 ();
 sg13g2_fill_2 FILLER_68_1455 ();
 sg13g2_fill_1 FILLER_68_1457 ();
 sg13g2_fill_1 FILLER_68_1462 ();
 sg13g2_fill_1 FILLER_68_1473 ();
 sg13g2_fill_2 FILLER_68_1479 ();
 sg13g2_fill_2 FILLER_68_1507 ();
 sg13g2_fill_2 FILLER_68_1513 ();
 sg13g2_decap_8 FILLER_68_1567 ();
 sg13g2_fill_1 FILLER_68_1574 ();
 sg13g2_decap_8 FILLER_68_1585 ();
 sg13g2_decap_8 FILLER_68_1592 ();
 sg13g2_decap_4 FILLER_68_1599 ();
 sg13g2_decap_8 FILLER_68_1615 ();
 sg13g2_decap_8 FILLER_68_1622 ();
 sg13g2_fill_2 FILLER_68_1629 ();
 sg13g2_fill_1 FILLER_68_1655 ();
 sg13g2_fill_2 FILLER_68_1697 ();
 sg13g2_fill_2 FILLER_68_1703 ();
 sg13g2_decap_8 FILLER_68_1709 ();
 sg13g2_decap_8 FILLER_68_1716 ();
 sg13g2_decap_8 FILLER_68_1723 ();
 sg13g2_fill_1 FILLER_68_1730 ();
 sg13g2_decap_8 FILLER_68_1767 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_43 ();
 sg13g2_decap_8 FILLER_69_50 ();
 sg13g2_decap_4 FILLER_69_57 ();
 sg13g2_fill_1 FILLER_69_71 ();
 sg13g2_fill_2 FILLER_69_86 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_fill_1 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_110 ();
 sg13g2_fill_1 FILLER_69_117 ();
 sg13g2_fill_2 FILLER_69_121 ();
 sg13g2_fill_1 FILLER_69_123 ();
 sg13g2_decap_8 FILLER_69_150 ();
 sg13g2_decap_8 FILLER_69_157 ();
 sg13g2_decap_4 FILLER_69_164 ();
 sg13g2_decap_4 FILLER_69_178 ();
 sg13g2_fill_2 FILLER_69_182 ();
 sg13g2_decap_8 FILLER_69_233 ();
 sg13g2_decap_8 FILLER_69_240 ();
 sg13g2_decap_8 FILLER_69_247 ();
 sg13g2_fill_2 FILLER_69_254 ();
 sg13g2_fill_2 FILLER_69_265 ();
 sg13g2_decap_8 FILLER_69_271 ();
 sg13g2_fill_2 FILLER_69_290 ();
 sg13g2_decap_8 FILLER_69_338 ();
 sg13g2_decap_8 FILLER_69_345 ();
 sg13g2_fill_2 FILLER_69_352 ();
 sg13g2_fill_1 FILLER_69_363 ();
 sg13g2_fill_1 FILLER_69_372 ();
 sg13g2_decap_4 FILLER_69_401 ();
 sg13g2_fill_2 FILLER_69_405 ();
 sg13g2_fill_2 FILLER_69_411 ();
 sg13g2_decap_4 FILLER_69_427 ();
 sg13g2_fill_2 FILLER_69_431 ();
 sg13g2_decap_8 FILLER_69_443 ();
 sg13g2_decap_8 FILLER_69_464 ();
 sg13g2_decap_4 FILLER_69_471 ();
 sg13g2_fill_1 FILLER_69_475 ();
 sg13g2_decap_4 FILLER_69_484 ();
 sg13g2_fill_1 FILLER_69_488 ();
 sg13g2_fill_1 FILLER_69_503 ();
 sg13g2_fill_2 FILLER_69_525 ();
 sg13g2_fill_1 FILLER_69_527 ();
 sg13g2_decap_8 FILLER_69_554 ();
 sg13g2_decap_4 FILLER_69_561 ();
 sg13g2_decap_8 FILLER_69_569 ();
 sg13g2_decap_8 FILLER_69_576 ();
 sg13g2_fill_1 FILLER_69_583 ();
 sg13g2_fill_2 FILLER_69_644 ();
 sg13g2_decap_8 FILLER_69_650 ();
 sg13g2_decap_4 FILLER_69_657 ();
 sg13g2_fill_2 FILLER_69_661 ();
 sg13g2_fill_1 FILLER_69_668 ();
 sg13g2_decap_8 FILLER_69_673 ();
 sg13g2_decap_4 FILLER_69_680 ();
 sg13g2_fill_1 FILLER_69_721 ();
 sg13g2_fill_1 FILLER_69_729 ();
 sg13g2_fill_2 FILLER_69_740 ();
 sg13g2_decap_8 FILLER_69_777 ();
 sg13g2_decap_4 FILLER_69_784 ();
 sg13g2_fill_2 FILLER_69_788 ();
 sg13g2_decap_8 FILLER_69_794 ();
 sg13g2_decap_8 FILLER_69_801 ();
 sg13g2_decap_8 FILLER_69_808 ();
 sg13g2_decap_4 FILLER_69_815 ();
 sg13g2_decap_8 FILLER_69_849 ();
 sg13g2_decap_8 FILLER_69_856 ();
 sg13g2_decap_8 FILLER_69_863 ();
 sg13g2_decap_8 FILLER_69_870 ();
 sg13g2_decap_4 FILLER_69_877 ();
 sg13g2_fill_2 FILLER_69_881 ();
 sg13g2_decap_4 FILLER_69_887 ();
 sg13g2_fill_2 FILLER_69_891 ();
 sg13g2_decap_4 FILLER_69_936 ();
 sg13g2_fill_2 FILLER_69_940 ();
 sg13g2_fill_1 FILLER_69_952 ();
 sg13g2_fill_1 FILLER_69_979 ();
 sg13g2_fill_1 FILLER_69_990 ();
 sg13g2_fill_2 FILLER_69_1017 ();
 sg13g2_decap_4 FILLER_69_1024 ();
 sg13g2_decap_4 FILLER_69_1041 ();
 sg13g2_fill_1 FILLER_69_1045 ();
 sg13g2_fill_2 FILLER_69_1128 ();
 sg13g2_fill_1 FILLER_69_1130 ();
 sg13g2_decap_4 FILLER_69_1161 ();
 sg13g2_fill_2 FILLER_69_1165 ();
 sg13g2_fill_1 FILLER_69_1177 ();
 sg13g2_decap_8 FILLER_69_1245 ();
 sg13g2_decap_8 FILLER_69_1252 ();
 sg13g2_decap_8 FILLER_69_1259 ();
 sg13g2_decap_8 FILLER_69_1266 ();
 sg13g2_decap_8 FILLER_69_1273 ();
 sg13g2_decap_8 FILLER_69_1280 ();
 sg13g2_fill_2 FILLER_69_1287 ();
 sg13g2_decap_8 FILLER_69_1293 ();
 sg13g2_fill_2 FILLER_69_1332 ();
 sg13g2_fill_2 FILLER_69_1367 ();
 sg13g2_fill_2 FILLER_69_1374 ();
 sg13g2_fill_1 FILLER_69_1376 ();
 sg13g2_fill_1 FILLER_69_1381 ();
 sg13g2_decap_4 FILLER_69_1395 ();
 sg13g2_fill_1 FILLER_69_1399 ();
 sg13g2_decap_8 FILLER_69_1404 ();
 sg13g2_decap_8 FILLER_69_1411 ();
 sg13g2_decap_4 FILLER_69_1418 ();
 sg13g2_fill_1 FILLER_69_1422 ();
 sg13g2_fill_1 FILLER_69_1439 ();
 sg13g2_fill_1 FILLER_69_1484 ();
 sg13g2_fill_1 FILLER_69_1525 ();
 sg13g2_fill_1 FILLER_69_1533 ();
 sg13g2_fill_1 FILLER_69_1552 ();
 sg13g2_fill_2 FILLER_69_1589 ();
 sg13g2_decap_8 FILLER_69_1601 ();
 sg13g2_decap_8 FILLER_69_1608 ();
 sg13g2_decap_8 FILLER_69_1615 ();
 sg13g2_decap_8 FILLER_69_1622 ();
 sg13g2_fill_2 FILLER_69_1629 ();
 sg13g2_fill_1 FILLER_69_1631 ();
 sg13g2_decap_8 FILLER_69_1658 ();
 sg13g2_decap_8 FILLER_69_1665 ();
 sg13g2_decap_4 FILLER_69_1672 ();
 sg13g2_fill_2 FILLER_69_1676 ();
 sg13g2_decap_8 FILLER_69_1682 ();
 sg13g2_fill_1 FILLER_69_1725 ();
 sg13g2_decap_8 FILLER_69_1740 ();
 sg13g2_fill_1 FILLER_69_1747 ();
 sg13g2_decap_8 FILLER_69_1752 ();
 sg13g2_decap_8 FILLER_69_1759 ();
 sg13g2_decap_8 FILLER_69_1766 ();
 sg13g2_fill_1 FILLER_69_1773 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_26 ();
 sg13g2_decap_4 FILLER_70_54 ();
 sg13g2_decap_8 FILLER_70_78 ();
 sg13g2_decap_8 FILLER_70_85 ();
 sg13g2_decap_4 FILLER_70_124 ();
 sg13g2_decap_8 FILLER_70_142 ();
 sg13g2_decap_8 FILLER_70_149 ();
 sg13g2_decap_8 FILLER_70_156 ();
 sg13g2_decap_8 FILLER_70_163 ();
 sg13g2_fill_2 FILLER_70_170 ();
 sg13g2_decap_4 FILLER_70_198 ();
 sg13g2_fill_1 FILLER_70_202 ();
 sg13g2_decap_8 FILLER_70_239 ();
 sg13g2_decap_8 FILLER_70_246 ();
 sg13g2_fill_2 FILLER_70_253 ();
 sg13g2_fill_1 FILLER_70_255 ();
 sg13g2_decap_8 FILLER_70_260 ();
 sg13g2_decap_8 FILLER_70_267 ();
 sg13g2_decap_4 FILLER_70_274 ();
 sg13g2_decap_8 FILLER_70_283 ();
 sg13g2_fill_2 FILLER_70_290 ();
 sg13g2_decap_8 FILLER_70_332 ();
 sg13g2_decap_8 FILLER_70_339 ();
 sg13g2_decap_4 FILLER_70_356 ();
 sg13g2_fill_2 FILLER_70_360 ();
 sg13g2_decap_8 FILLER_70_380 ();
 sg13g2_decap_8 FILLER_70_387 ();
 sg13g2_fill_1 FILLER_70_394 ();
 sg13g2_fill_1 FILLER_70_425 ();
 sg13g2_fill_2 FILLER_70_434 ();
 sg13g2_decap_8 FILLER_70_446 ();
 sg13g2_fill_1 FILLER_70_453 ();
 sg13g2_fill_2 FILLER_70_464 ();
 sg13g2_fill_1 FILLER_70_466 ();
 sg13g2_fill_2 FILLER_70_473 ();
 sg13g2_decap_4 FILLER_70_483 ();
 sg13g2_fill_1 FILLER_70_487 ();
 sg13g2_decap_4 FILLER_70_548 ();
 sg13g2_fill_1 FILLER_70_552 ();
 sg13g2_decap_4 FILLER_70_556 ();
 sg13g2_fill_1 FILLER_70_560 ();
 sg13g2_fill_2 FILLER_70_597 ();
 sg13g2_fill_1 FILLER_70_599 ();
 sg13g2_decap_8 FILLER_70_604 ();
 sg13g2_decap_8 FILLER_70_611 ();
 sg13g2_fill_1 FILLER_70_618 ();
 sg13g2_decap_4 FILLER_70_623 ();
 sg13g2_fill_1 FILLER_70_627 ();
 sg13g2_decap_4 FILLER_70_677 ();
 sg13g2_decap_8 FILLER_70_699 ();
 sg13g2_decap_8 FILLER_70_706 ();
 sg13g2_fill_2 FILLER_70_713 ();
 sg13g2_decap_4 FILLER_70_721 ();
 sg13g2_fill_2 FILLER_70_782 ();
 sg13g2_fill_1 FILLER_70_784 ();
 sg13g2_fill_2 FILLER_70_799 ();
 sg13g2_fill_1 FILLER_70_801 ();
 sg13g2_decap_4 FILLER_70_810 ();
 sg13g2_fill_2 FILLER_70_814 ();
 sg13g2_fill_2 FILLER_70_830 ();
 sg13g2_fill_1 FILLER_70_832 ();
 sg13g2_decap_8 FILLER_70_837 ();
 sg13g2_decap_8 FILLER_70_844 ();
 sg13g2_decap_8 FILLER_70_851 ();
 sg13g2_decap_8 FILLER_70_858 ();
 sg13g2_decap_8 FILLER_70_865 ();
 sg13g2_decap_8 FILLER_70_872 ();
 sg13g2_fill_1 FILLER_70_879 ();
 sg13g2_decap_4 FILLER_70_907 ();
 sg13g2_decap_4 FILLER_70_921 ();
 sg13g2_decap_8 FILLER_70_933 ();
 sg13g2_fill_1 FILLER_70_940 ();
 sg13g2_decap_8 FILLER_70_951 ();
 sg13g2_fill_1 FILLER_70_958 ();
 sg13g2_fill_2 FILLER_70_973 ();
 sg13g2_decap_8 FILLER_70_996 ();
 sg13g2_decap_8 FILLER_70_1011 ();
 sg13g2_decap_8 FILLER_70_1018 ();
 sg13g2_decap_8 FILLER_70_1025 ();
 sg13g2_decap_8 FILLER_70_1032 ();
 sg13g2_decap_8 FILLER_70_1039 ();
 sg13g2_fill_2 FILLER_70_1046 ();
 sg13g2_fill_1 FILLER_70_1048 ();
 sg13g2_decap_4 FILLER_70_1054 ();
 sg13g2_fill_1 FILLER_70_1058 ();
 sg13g2_decap_8 FILLER_70_1073 ();
 sg13g2_decap_8 FILLER_70_1080 ();
 sg13g2_fill_2 FILLER_70_1087 ();
 sg13g2_fill_1 FILLER_70_1089 ();
 sg13g2_fill_2 FILLER_70_1112 ();
 sg13g2_fill_1 FILLER_70_1124 ();
 sg13g2_fill_1 FILLER_70_1138 ();
 sg13g2_decap_8 FILLER_70_1149 ();
 sg13g2_fill_1 FILLER_70_1166 ();
 sg13g2_fill_2 FILLER_70_1175 ();
 sg13g2_fill_2 FILLER_70_1181 ();
 sg13g2_fill_1 FILLER_70_1183 ();
 sg13g2_decap_8 FILLER_70_1188 ();
 sg13g2_fill_2 FILLER_70_1195 ();
 sg13g2_fill_1 FILLER_70_1197 ();
 sg13g2_fill_2 FILLER_70_1210 ();
 sg13g2_fill_1 FILLER_70_1225 ();
 sg13g2_decap_4 FILLER_70_1230 ();
 sg13g2_decap_4 FILLER_70_1244 ();
 sg13g2_fill_1 FILLER_70_1303 ();
 sg13g2_fill_1 FILLER_70_1333 ();
 sg13g2_decap_8 FILLER_70_1366 ();
 sg13g2_fill_1 FILLER_70_1373 ();
 sg13g2_fill_1 FILLER_70_1378 ();
 sg13g2_fill_2 FILLER_70_1395 ();
 sg13g2_decap_4 FILLER_70_1413 ();
 sg13g2_fill_2 FILLER_70_1417 ();
 sg13g2_fill_1 FILLER_70_1422 ();
 sg13g2_fill_2 FILLER_70_1428 ();
 sg13g2_fill_2 FILLER_70_1460 ();
 sg13g2_decap_4 FILLER_70_1488 ();
 sg13g2_decap_4 FILLER_70_1538 ();
 sg13g2_decap_8 FILLER_70_1628 ();
 sg13g2_fill_2 FILLER_70_1635 ();
 sg13g2_decap_8 FILLER_70_1691 ();
 sg13g2_decap_8 FILLER_70_1698 ();
 sg13g2_decap_8 FILLER_70_1759 ();
 sg13g2_decap_8 FILLER_70_1766 ();
 sg13g2_fill_1 FILLER_70_1773 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_34 ();
 sg13g2_decap_8 FILLER_71_75 ();
 sg13g2_fill_2 FILLER_71_82 ();
 sg13g2_decap_8 FILLER_71_94 ();
 sg13g2_decap_8 FILLER_71_101 ();
 sg13g2_decap_4 FILLER_71_108 ();
 sg13g2_decap_8 FILLER_71_122 ();
 sg13g2_fill_2 FILLER_71_129 ();
 sg13g2_decap_8 FILLER_71_141 ();
 sg13g2_decap_8 FILLER_71_148 ();
 sg13g2_decap_4 FILLER_71_155 ();
 sg13g2_decap_8 FILLER_71_183 ();
 sg13g2_decap_8 FILLER_71_194 ();
 sg13g2_decap_4 FILLER_71_201 ();
 sg13g2_fill_2 FILLER_71_205 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_4 FILLER_71_224 ();
 sg13g2_fill_1 FILLER_71_228 ();
 sg13g2_decap_4 FILLER_71_275 ();
 sg13g2_fill_2 FILLER_71_279 ();
 sg13g2_decap_8 FILLER_71_286 ();
 sg13g2_decap_8 FILLER_71_293 ();
 sg13g2_decap_4 FILLER_71_300 ();
 sg13g2_fill_2 FILLER_71_304 ();
 sg13g2_fill_2 FILLER_71_346 ();
 sg13g2_fill_1 FILLER_71_358 ();
 sg13g2_fill_1 FILLER_71_369 ();
 sg13g2_fill_1 FILLER_71_380 ();
 sg13g2_decap_4 FILLER_71_391 ();
 sg13g2_fill_1 FILLER_71_395 ();
 sg13g2_fill_1 FILLER_71_406 ();
 sg13g2_decap_4 FILLER_71_417 ();
 sg13g2_fill_2 FILLER_71_447 ();
 sg13g2_fill_1 FILLER_71_449 ();
 sg13g2_decap_4 FILLER_71_507 ();
 sg13g2_fill_1 FILLER_71_537 ();
 sg13g2_fill_2 FILLER_71_548 ();
 sg13g2_fill_1 FILLER_71_571 ();
 sg13g2_decap_8 FILLER_71_611 ();
 sg13g2_decap_8 FILLER_71_618 ();
 sg13g2_decap_8 FILLER_71_661 ();
 sg13g2_fill_2 FILLER_71_668 ();
 sg13g2_fill_2 FILLER_71_675 ();
 sg13g2_fill_2 FILLER_71_685 ();
 sg13g2_fill_2 FILLER_71_705 ();
 sg13g2_fill_1 FILLER_71_759 ();
 sg13g2_fill_1 FILLER_71_764 ();
 sg13g2_fill_1 FILLER_71_770 ();
 sg13g2_fill_1 FILLER_71_797 ();
 sg13g2_fill_1 FILLER_71_824 ();
 sg13g2_fill_1 FILLER_71_851 ();
 sg13g2_decap_8 FILLER_71_856 ();
 sg13g2_decap_4 FILLER_71_863 ();
 sg13g2_decap_4 FILLER_71_875 ();
 sg13g2_fill_1 FILLER_71_879 ();
 sg13g2_decap_4 FILLER_71_920 ();
 sg13g2_fill_2 FILLER_71_924 ();
 sg13g2_fill_2 FILLER_71_962 ();
 sg13g2_fill_2 FILLER_71_990 ();
 sg13g2_decap_8 FILLER_71_1038 ();
 sg13g2_decap_8 FILLER_71_1045 ();
 sg13g2_fill_2 FILLER_71_1052 ();
 sg13g2_decap_4 FILLER_71_1074 ();
 sg13g2_fill_1 FILLER_71_1108 ();
 sg13g2_decap_8 FILLER_71_1122 ();
 sg13g2_decap_8 FILLER_71_1129 ();
 sg13g2_fill_2 FILLER_71_1136 ();
 sg13g2_decap_8 FILLER_71_1142 ();
 sg13g2_decap_8 FILLER_71_1149 ();
 sg13g2_fill_1 FILLER_71_1156 ();
 sg13g2_fill_1 FILLER_71_1175 ();
 sg13g2_fill_1 FILLER_71_1218 ();
 sg13g2_fill_2 FILLER_71_1224 ();
 sg13g2_fill_2 FILLER_71_1237 ();
 sg13g2_fill_2 FILLER_71_1251 ();
 sg13g2_fill_1 FILLER_71_1263 ();
 sg13g2_fill_2 FILLER_71_1375 ();
 sg13g2_fill_1 FILLER_71_1377 ();
 sg13g2_decap_4 FILLER_71_1382 ();
 sg13g2_fill_1 FILLER_71_1402 ();
 sg13g2_fill_1 FILLER_71_1435 ();
 sg13g2_fill_1 FILLER_71_1449 ();
 sg13g2_decap_8 FILLER_71_1460 ();
 sg13g2_decap_4 FILLER_71_1467 ();
 sg13g2_fill_2 FILLER_71_1513 ();
 sg13g2_decap_8 FILLER_71_1520 ();
 sg13g2_decap_4 FILLER_71_1527 ();
 sg13g2_fill_1 FILLER_71_1531 ();
 sg13g2_fill_2 FILLER_71_1549 ();
 sg13g2_fill_1 FILLER_71_1569 ();
 sg13g2_fill_2 FILLER_71_1587 ();
 sg13g2_decap_4 FILLER_71_1599 ();
 sg13g2_decap_4 FILLER_71_1606 ();
 sg13g2_fill_2 FILLER_71_1610 ();
 sg13g2_decap_8 FILLER_71_1620 ();
 sg13g2_decap_8 FILLER_71_1627 ();
 sg13g2_decap_8 FILLER_71_1634 ();
 sg13g2_fill_2 FILLER_71_1641 ();
 sg13g2_fill_1 FILLER_71_1643 ();
 sg13g2_decap_4 FILLER_71_1674 ();
 sg13g2_decap_8 FILLER_71_1766 ();
 sg13g2_fill_1 FILLER_71_1773 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_45 ();
 sg13g2_fill_1 FILLER_72_72 ();
 sg13g2_fill_1 FILLER_72_99 ();
 sg13g2_fill_1 FILLER_72_110 ();
 sg13g2_fill_2 FILLER_72_121 ();
 sg13g2_fill_1 FILLER_72_123 ();
 sg13g2_fill_1 FILLER_72_170 ();
 sg13g2_fill_2 FILLER_72_211 ();
 sg13g2_decap_8 FILLER_72_223 ();
 sg13g2_fill_1 FILLER_72_230 ();
 sg13g2_decap_4 FILLER_72_277 ();
 sg13g2_decap_4 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_fill_1 FILLER_72_336 ();
 sg13g2_fill_2 FILLER_72_367 ();
 sg13g2_fill_1 FILLER_72_369 ();
 sg13g2_fill_2 FILLER_72_396 ();
 sg13g2_fill_2 FILLER_72_465 ();
 sg13g2_fill_2 FILLER_72_471 ();
 sg13g2_fill_1 FILLER_72_473 ();
 sg13g2_fill_2 FILLER_72_480 ();
 sg13g2_fill_1 FILLER_72_482 ();
 sg13g2_fill_2 FILLER_72_487 ();
 sg13g2_fill_1 FILLER_72_493 ();
 sg13g2_fill_2 FILLER_72_504 ();
 sg13g2_fill_1 FILLER_72_506 ();
 sg13g2_fill_2 FILLER_72_511 ();
 sg13g2_fill_1 FILLER_72_513 ();
 sg13g2_fill_1 FILLER_72_558 ();
 sg13g2_fill_1 FILLER_72_577 ();
 sg13g2_fill_2 FILLER_72_595 ();
 sg13g2_fill_1 FILLER_72_597 ();
 sg13g2_fill_2 FILLER_72_603 ();
 sg13g2_decap_8 FILLER_72_609 ();
 sg13g2_decap_4 FILLER_72_620 ();
 sg13g2_fill_2 FILLER_72_624 ();
 sg13g2_decap_8 FILLER_72_678 ();
 sg13g2_fill_1 FILLER_72_685 ();
 sg13g2_decap_8 FILLER_72_690 ();
 sg13g2_fill_2 FILLER_72_697 ();
 sg13g2_fill_2 FILLER_72_704 ();
 sg13g2_decap_8 FILLER_72_710 ();
 sg13g2_fill_1 FILLER_72_729 ();
 sg13g2_fill_2 FILLER_72_789 ();
 sg13g2_fill_1 FILLER_72_791 ();
 sg13g2_decap_4 FILLER_72_797 ();
 sg13g2_fill_2 FILLER_72_815 ();
 sg13g2_decap_4 FILLER_72_821 ();
 sg13g2_fill_2 FILLER_72_825 ();
 sg13g2_fill_1 FILLER_72_857 ();
 sg13g2_fill_1 FILLER_72_863 ();
 sg13g2_decap_8 FILLER_72_870 ();
 sg13g2_fill_1 FILLER_72_877 ();
 sg13g2_fill_2 FILLER_72_918 ();
 sg13g2_fill_1 FILLER_72_950 ();
 sg13g2_decap_8 FILLER_72_955 ();
 sg13g2_decap_8 FILLER_72_966 ();
 sg13g2_decap_4 FILLER_72_998 ();
 sg13g2_decap_8 FILLER_72_1032 ();
 sg13g2_decap_8 FILLER_72_1039 ();
 sg13g2_decap_4 FILLER_72_1113 ();
 sg13g2_fill_2 FILLER_72_1170 ();
 sg13g2_fill_1 FILLER_72_1172 ();
 sg13g2_fill_2 FILLER_72_1183 ();
 sg13g2_fill_1 FILLER_72_1224 ();
 sg13g2_fill_2 FILLER_72_1255 ();
 sg13g2_fill_2 FILLER_72_1275 ();
 sg13g2_fill_1 FILLER_72_1281 ();
 sg13g2_fill_2 FILLER_72_1308 ();
 sg13g2_fill_2 FILLER_72_1376 ();
 sg13g2_fill_1 FILLER_72_1378 ();
 sg13g2_fill_2 FILLER_72_1388 ();
 sg13g2_decap_4 FILLER_72_1395 ();
 sg13g2_fill_2 FILLER_72_1413 ();
 sg13g2_fill_1 FILLER_72_1418 ();
 sg13g2_fill_2 FILLER_72_1434 ();
 sg13g2_decap_4 FILLER_72_1482 ();
 sg13g2_fill_1 FILLER_72_1486 ();
 sg13g2_fill_2 FILLER_72_1541 ();
 sg13g2_fill_1 FILLER_72_1550 ();
 sg13g2_fill_1 FILLER_72_1598 ();
 sg13g2_fill_2 FILLER_72_1635 ();
 sg13g2_decap_8 FILLER_72_1683 ();
 sg13g2_decap_4 FILLER_72_1690 ();
 sg13g2_fill_1 FILLER_72_1694 ();
 sg13g2_decap_8 FILLER_72_1699 ();
 sg13g2_fill_1 FILLER_72_1706 ();
 sg13g2_decap_4 FILLER_72_1742 ();
 sg13g2_fill_2 FILLER_72_1746 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_7 ();
 sg13g2_fill_1 FILLER_73_9 ();
 sg13g2_fill_2 FILLER_73_72 ();
 sg13g2_decap_8 FILLER_73_82 ();
 sg13g2_decap_8 FILLER_73_89 ();
 sg13g2_decap_4 FILLER_73_96 ();
 sg13g2_fill_1 FILLER_73_146 ();
 sg13g2_fill_2 FILLER_73_161 ();
 sg13g2_fill_1 FILLER_73_163 ();
 sg13g2_decap_8 FILLER_73_190 ();
 sg13g2_fill_2 FILLER_73_243 ();
 sg13g2_fill_1 FILLER_73_245 ();
 sg13g2_fill_2 FILLER_73_279 ();
 sg13g2_decap_8 FILLER_73_286 ();
 sg13g2_decap_4 FILLER_73_293 ();
 sg13g2_fill_1 FILLER_73_297 ();
 sg13g2_fill_1 FILLER_73_302 ();
 sg13g2_fill_1 FILLER_73_313 ();
 sg13g2_fill_1 FILLER_73_340 ();
 sg13g2_decap_4 FILLER_73_351 ();
 sg13g2_fill_1 FILLER_73_355 ();
 sg13g2_fill_1 FILLER_73_360 ();
 sg13g2_fill_2 FILLER_73_453 ();
 sg13g2_decap_4 FILLER_73_464 ();
 sg13g2_fill_2 FILLER_73_478 ();
 sg13g2_decap_8 FILLER_73_484 ();
 sg13g2_fill_1 FILLER_73_491 ();
 sg13g2_fill_1 FILLER_73_512 ();
 sg13g2_decap_8 FILLER_73_521 ();
 sg13g2_fill_1 FILLER_73_528 ();
 sg13g2_decap_8 FILLER_73_575 ();
 sg13g2_decap_8 FILLER_73_582 ();
 sg13g2_decap_8 FILLER_73_589 ();
 sg13g2_decap_4 FILLER_73_596 ();
 sg13g2_fill_2 FILLER_73_604 ();
 sg13g2_fill_2 FILLER_73_616 ();
 sg13g2_fill_1 FILLER_73_618 ();
 sg13g2_fill_1 FILLER_73_669 ();
 sg13g2_decap_8 FILLER_73_675 ();
 sg13g2_decap_8 FILLER_73_682 ();
 sg13g2_decap_8 FILLER_73_689 ();
 sg13g2_decap_8 FILLER_73_696 ();
 sg13g2_decap_8 FILLER_73_703 ();
 sg13g2_decap_4 FILLER_73_710 ();
 sg13g2_fill_1 FILLER_73_759 ();
 sg13g2_decap_4 FILLER_73_806 ();
 sg13g2_fill_1 FILLER_73_862 ();
 sg13g2_fill_2 FILLER_73_868 ();
 sg13g2_fill_2 FILLER_73_874 ();
 sg13g2_decap_8 FILLER_73_944 ();
 sg13g2_fill_2 FILLER_73_951 ();
 sg13g2_fill_1 FILLER_73_953 ();
 sg13g2_fill_2 FILLER_73_975 ();
 sg13g2_decap_8 FILLER_73_1039 ();
 sg13g2_fill_2 FILLER_73_1046 ();
 sg13g2_decap_4 FILLER_73_1062 ();
 sg13g2_fill_2 FILLER_73_1150 ();
 sg13g2_fill_2 FILLER_73_1178 ();
 sg13g2_fill_1 FILLER_73_1206 ();
 sg13g2_decap_4 FILLER_73_1241 ();
 sg13g2_fill_2 FILLER_73_1245 ();
 sg13g2_fill_1 FILLER_73_1262 ();
 sg13g2_decap_4 FILLER_73_1279 ();
 sg13g2_fill_2 FILLER_73_1283 ();
 sg13g2_decap_8 FILLER_73_1290 ();
 sg13g2_fill_2 FILLER_73_1297 ();
 sg13g2_fill_1 FILLER_73_1299 ();
 sg13g2_fill_2 FILLER_73_1310 ();
 sg13g2_fill_1 FILLER_73_1312 ();
 sg13g2_fill_1 FILLER_73_1327 ();
 sg13g2_fill_1 FILLER_73_1341 ();
 sg13g2_fill_2 FILLER_73_1346 ();
 sg13g2_fill_2 FILLER_73_1384 ();
 sg13g2_fill_1 FILLER_73_1386 ();
 sg13g2_decap_4 FILLER_73_1403 ();
 sg13g2_fill_2 FILLER_73_1413 ();
 sg13g2_fill_2 FILLER_73_1444 ();
 sg13g2_fill_1 FILLER_73_1458 ();
 sg13g2_fill_1 FILLER_73_1485 ();
 sg13g2_fill_2 FILLER_73_1553 ();
 sg13g2_fill_1 FILLER_73_1562 ();
 sg13g2_fill_1 FILLER_73_1570 ();
 sg13g2_fill_1 FILLER_73_1612 ();
 sg13g2_fill_2 FILLER_73_1629 ();
 sg13g2_fill_1 FILLER_73_1631 ();
 sg13g2_fill_2 FILLER_73_1636 ();
 sg13g2_fill_1 FILLER_73_1638 ();
 sg13g2_fill_2 FILLER_73_1649 ();
 sg13g2_decap_8 FILLER_73_1676 ();
 sg13g2_decap_8 FILLER_73_1683 ();
 sg13g2_decap_8 FILLER_73_1690 ();
 sg13g2_decap_8 FILLER_73_1697 ();
 sg13g2_decap_4 FILLER_73_1704 ();
 sg13g2_fill_2 FILLER_73_1708 ();
 sg13g2_fill_2 FILLER_73_1771 ();
 sg13g2_fill_1 FILLER_73_1773 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_14 ();
 sg13g2_decap_4 FILLER_74_20 ();
 sg13g2_decap_4 FILLER_74_58 ();
 sg13g2_decap_8 FILLER_74_66 ();
 sg13g2_fill_1 FILLER_74_73 ();
 sg13g2_decap_4 FILLER_74_78 ();
 sg13g2_fill_2 FILLER_74_82 ();
 sg13g2_decap_4 FILLER_74_150 ();
 sg13g2_fill_1 FILLER_74_154 ();
 sg13g2_decap_4 FILLER_74_185 ();
 sg13g2_fill_1 FILLER_74_189 ();
 sg13g2_fill_2 FILLER_74_239 ();
 sg13g2_fill_1 FILLER_74_241 ();
 sg13g2_decap_4 FILLER_74_279 ();
 sg13g2_fill_1 FILLER_74_283 ();
 sg13g2_fill_1 FILLER_74_287 ();
 sg13g2_decap_4 FILLER_74_298 ();
 sg13g2_fill_2 FILLER_74_328 ();
 sg13g2_fill_1 FILLER_74_330 ();
 sg13g2_decap_8 FILLER_74_335 ();
 sg13g2_decap_8 FILLER_74_342 ();
 sg13g2_decap_4 FILLER_74_383 ();
 sg13g2_fill_2 FILLER_74_391 ();
 sg13g2_decap_8 FILLER_74_439 ();
 sg13g2_decap_8 FILLER_74_446 ();
 sg13g2_decap_8 FILLER_74_453 ();
 sg13g2_fill_2 FILLER_74_460 ();
 sg13g2_fill_1 FILLER_74_462 ();
 sg13g2_decap_8 FILLER_74_499 ();
 sg13g2_decap_8 FILLER_74_506 ();
 sg13g2_decap_8 FILLER_74_513 ();
 sg13g2_fill_2 FILLER_74_520 ();
 sg13g2_fill_1 FILLER_74_522 ();
 sg13g2_fill_1 FILLER_74_528 ();
 sg13g2_decap_8 FILLER_74_532 ();
 sg13g2_decap_8 FILLER_74_539 ();
 sg13g2_decap_8 FILLER_74_546 ();
 sg13g2_fill_1 FILLER_74_553 ();
 sg13g2_decap_4 FILLER_74_580 ();
 sg13g2_fill_1 FILLER_74_584 ();
 sg13g2_decap_4 FILLER_74_591 ();
 sg13g2_fill_2 FILLER_74_660 ();
 sg13g2_decap_8 FILLER_74_672 ();
 sg13g2_decap_8 FILLER_74_679 ();
 sg13g2_decap_8 FILLER_74_686 ();
 sg13g2_decap_4 FILLER_74_706 ();
 sg13g2_fill_1 FILLER_74_710 ();
 sg13g2_fill_2 FILLER_74_737 ();
 sg13g2_fill_1 FILLER_74_753 ();
 sg13g2_decap_4 FILLER_74_764 ();
 sg13g2_decap_4 FILLER_74_773 ();
 sg13g2_decap_8 FILLER_74_781 ();
 sg13g2_decap_8 FILLER_74_828 ();
 sg13g2_fill_2 FILLER_74_835 ();
 sg13g2_fill_1 FILLER_74_837 ();
 sg13g2_decap_8 FILLER_74_864 ();
 sg13g2_decap_4 FILLER_74_871 ();
 sg13g2_decap_8 FILLER_74_879 ();
 sg13g2_fill_1 FILLER_74_886 ();
 sg13g2_fill_2 FILLER_74_891 ();
 sg13g2_decap_4 FILLER_74_903 ();
 sg13g2_decap_4 FILLER_74_917 ();
 sg13g2_decap_4 FILLER_74_957 ();
 sg13g2_fill_1 FILLER_74_961 ();
 sg13g2_decap_8 FILLER_74_966 ();
 sg13g2_decap_4 FILLER_74_973 ();
 sg13g2_fill_2 FILLER_74_1026 ();
 sg13g2_decap_8 FILLER_74_1032 ();
 sg13g2_decap_8 FILLER_74_1039 ();
 sg13g2_fill_2 FILLER_74_1046 ();
 sg13g2_decap_4 FILLER_74_1053 ();
 sg13g2_fill_1 FILLER_74_1057 ();
 sg13g2_fill_1 FILLER_74_1063 ();
 sg13g2_fill_2 FILLER_74_1078 ();
 sg13g2_fill_1 FILLER_74_1084 ();
 sg13g2_fill_2 FILLER_74_1089 ();
 sg13g2_fill_2 FILLER_74_1101 ();
 sg13g2_fill_2 FILLER_74_1124 ();
 sg13g2_fill_1 FILLER_74_1201 ();
 sg13g2_fill_2 FILLER_74_1227 ();
 sg13g2_decap_8 FILLER_74_1233 ();
 sg13g2_fill_2 FILLER_74_1240 ();
 sg13g2_fill_1 FILLER_74_1242 ();
 sg13g2_decap_8 FILLER_74_1279 ();
 sg13g2_decap_4 FILLER_74_1286 ();
 sg13g2_fill_2 FILLER_74_1290 ();
 sg13g2_fill_1 FILLER_74_1358 ();
 sg13g2_fill_2 FILLER_74_1369 ();
 sg13g2_decap_8 FILLER_74_1410 ();
 sg13g2_decap_4 FILLER_74_1417 ();
 sg13g2_fill_2 FILLER_74_1427 ();
 sg13g2_decap_8 FILLER_74_1478 ();
 sg13g2_decap_8 FILLER_74_1485 ();
 sg13g2_decap_8 FILLER_74_1496 ();
 sg13g2_decap_8 FILLER_74_1503 ();
 sg13g2_fill_1 FILLER_74_1561 ();
 sg13g2_fill_2 FILLER_74_1570 ();
 sg13g2_fill_2 FILLER_74_1585 ();
 sg13g2_fill_1 FILLER_74_1675 ();
 sg13g2_decap_4 FILLER_74_1686 ();
 sg13g2_decap_4 FILLER_74_1726 ();
 sg13g2_fill_1 FILLER_74_1740 ();
 sg13g2_decap_8 FILLER_74_1767 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_4 FILLER_75_21 ();
 sg13g2_fill_1 FILLER_75_25 ();
 sg13g2_decap_8 FILLER_75_66 ();
 sg13g2_decap_4 FILLER_75_73 ();
 sg13g2_fill_2 FILLER_75_77 ();
 sg13g2_fill_2 FILLER_75_89 ();
 sg13g2_decap_8 FILLER_75_101 ();
 sg13g2_decap_8 FILLER_75_142 ();
 sg13g2_decap_8 FILLER_75_149 ();
 sg13g2_fill_2 FILLER_75_156 ();
 sg13g2_fill_1 FILLER_75_158 ();
 sg13g2_fill_1 FILLER_75_163 ();
 sg13g2_decap_8 FILLER_75_172 ();
 sg13g2_decap_8 FILLER_75_179 ();
 sg13g2_fill_2 FILLER_75_195 ();
 sg13g2_fill_1 FILLER_75_201 ();
 sg13g2_fill_1 FILLER_75_206 ();
 sg13g2_fill_2 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_226 ();
 sg13g2_decap_4 FILLER_75_233 ();
 sg13g2_fill_2 FILLER_75_237 ();
 sg13g2_decap_4 FILLER_75_243 ();
 sg13g2_fill_1 FILLER_75_284 ();
 sg13g2_fill_2 FILLER_75_320 ();
 sg13g2_fill_1 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_327 ();
 sg13g2_decap_8 FILLER_75_334 ();
 sg13g2_fill_2 FILLER_75_341 ();
 sg13g2_decap_4 FILLER_75_348 ();
 sg13g2_fill_2 FILLER_75_352 ();
 sg13g2_decap_8 FILLER_75_358 ();
 sg13g2_decap_8 FILLER_75_365 ();
 sg13g2_decap_8 FILLER_75_372 ();
 sg13g2_decap_8 FILLER_75_379 ();
 sg13g2_decap_8 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_decap_8 FILLER_75_407 ();
 sg13g2_decap_4 FILLER_75_414 ();
 sg13g2_fill_2 FILLER_75_418 ();
 sg13g2_fill_2 FILLER_75_424 ();
 sg13g2_decap_8 FILLER_75_430 ();
 sg13g2_fill_2 FILLER_75_437 ();
 sg13g2_fill_1 FILLER_75_439 ();
 sg13g2_decap_8 FILLER_75_445 ();
 sg13g2_decap_8 FILLER_75_452 ();
 sg13g2_decap_8 FILLER_75_489 ();
 sg13g2_decap_8 FILLER_75_496 ();
 sg13g2_fill_2 FILLER_75_503 ();
 sg13g2_fill_1 FILLER_75_528 ();
 sg13g2_fill_2 FILLER_75_560 ();
 sg13g2_fill_2 FILLER_75_566 ();
 sg13g2_fill_1 FILLER_75_568 ();
 sg13g2_fill_1 FILLER_75_574 ();
 sg13g2_fill_2 FILLER_75_585 ();
 sg13g2_fill_1 FILLER_75_587 ();
 sg13g2_fill_1 FILLER_75_592 ();
 sg13g2_fill_1 FILLER_75_598 ();
 sg13g2_fill_2 FILLER_75_604 ();
 sg13g2_fill_2 FILLER_75_611 ();
 sg13g2_decap_8 FILLER_75_617 ();
 sg13g2_decap_8 FILLER_75_648 ();
 sg13g2_decap_4 FILLER_75_655 ();
 sg13g2_fill_2 FILLER_75_679 ();
 sg13g2_decap_8 FILLER_75_686 ();
 sg13g2_decap_4 FILLER_75_693 ();
 sg13g2_decap_8 FILLER_75_738 ();
 sg13g2_decap_4 FILLER_75_745 ();
 sg13g2_fill_2 FILLER_75_749 ();
 sg13g2_decap_8 FILLER_75_761 ();
 sg13g2_decap_8 FILLER_75_768 ();
 sg13g2_decap_8 FILLER_75_775 ();
 sg13g2_decap_4 FILLER_75_782 ();
 sg13g2_decap_4 FILLER_75_822 ();
 sg13g2_fill_1 FILLER_75_826 ();
 sg13g2_decap_4 FILLER_75_858 ();
 sg13g2_decap_8 FILLER_75_867 ();
 sg13g2_decap_8 FILLER_75_874 ();
 sg13g2_decap_8 FILLER_75_881 ();
 sg13g2_decap_8 FILLER_75_888 ();
 sg13g2_fill_1 FILLER_75_895 ();
 sg13g2_decap_8 FILLER_75_917 ();
 sg13g2_decap_8 FILLER_75_928 ();
 sg13g2_fill_2 FILLER_75_935 ();
 sg13g2_fill_1 FILLER_75_937 ();
 sg13g2_decap_4 FILLER_75_948 ();
 sg13g2_fill_1 FILLER_75_952 ();
 sg13g2_decap_8 FILLER_75_979 ();
 sg13g2_fill_2 FILLER_75_986 ();
 sg13g2_fill_1 FILLER_75_988 ();
 sg13g2_decap_8 FILLER_75_1029 ();
 sg13g2_decap_8 FILLER_75_1036 ();
 sg13g2_fill_2 FILLER_75_1053 ();
 sg13g2_fill_1 FILLER_75_1055 ();
 sg13g2_decap_8 FILLER_75_1066 ();
 sg13g2_decap_8 FILLER_75_1073 ();
 sg13g2_decap_4 FILLER_75_1080 ();
 sg13g2_fill_1 FILLER_75_1084 ();
 sg13g2_fill_1 FILLER_75_1126 ();
 sg13g2_decap_8 FILLER_75_1132 ();
 sg13g2_fill_1 FILLER_75_1169 ();
 sg13g2_fill_1 FILLER_75_1191 ();
 sg13g2_fill_1 FILLER_75_1196 ();
 sg13g2_fill_1 FILLER_75_1207 ();
 sg13g2_decap_4 FILLER_75_1234 ();
 sg13g2_decap_8 FILLER_75_1243 ();
 sg13g2_fill_2 FILLER_75_1250 ();
 sg13g2_fill_1 FILLER_75_1252 ();
 sg13g2_decap_8 FILLER_75_1267 ();
 sg13g2_fill_2 FILLER_75_1278 ();
 sg13g2_fill_1 FILLER_75_1280 ();
 sg13g2_decap_8 FILLER_75_1312 ();
 sg13g2_decap_8 FILLER_75_1319 ();
 sg13g2_fill_2 FILLER_75_1326 ();
 sg13g2_fill_1 FILLER_75_1375 ();
 sg13g2_decap_8 FILLER_75_1420 ();
 sg13g2_fill_2 FILLER_75_1427 ();
 sg13g2_decap_8 FILLER_75_1434 ();
 sg13g2_decap_4 FILLER_75_1441 ();
 sg13g2_fill_2 FILLER_75_1445 ();
 sg13g2_decap_8 FILLER_75_1461 ();
 sg13g2_fill_2 FILLER_75_1468 ();
 sg13g2_decap_4 FILLER_75_1474 ();
 sg13g2_decap_4 FILLER_75_1488 ();
 sg13g2_decap_8 FILLER_75_1502 ();
 sg13g2_decap_4 FILLER_75_1509 ();
 sg13g2_fill_1 FILLER_75_1513 ();
 sg13g2_decap_4 FILLER_75_1524 ();
 sg13g2_fill_2 FILLER_75_1528 ();
 sg13g2_fill_1 FILLER_75_1534 ();
 sg13g2_fill_1 FILLER_75_1539 ();
 sg13g2_fill_1 FILLER_75_1550 ();
 sg13g2_fill_1 FILLER_75_1605 ();
 sg13g2_fill_2 FILLER_75_1610 ();
 sg13g2_decap_4 FILLER_75_1650 ();
 sg13g2_decap_4 FILLER_75_1658 ();
 sg13g2_fill_2 FILLER_75_1662 ();
 sg13g2_fill_2 FILLER_75_1698 ();
 sg13g2_fill_2 FILLER_75_1710 ();
 sg13g2_fill_2 FILLER_75_1716 ();
 sg13g2_fill_1 FILLER_75_1718 ();
 sg13g2_fill_2 FILLER_75_1729 ();
 sg13g2_fill_1 FILLER_75_1731 ();
 sg13g2_decap_8 FILLER_75_1762 ();
 sg13g2_decap_4 FILLER_75_1769 ();
 sg13g2_fill_1 FILLER_75_1773 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_4 FILLER_76_14 ();
 sg13g2_fill_1 FILLER_76_18 ();
 sg13g2_decap_8 FILLER_76_55 ();
 sg13g2_decap_4 FILLER_76_62 ();
 sg13g2_fill_2 FILLER_76_66 ();
 sg13g2_fill_1 FILLER_76_78 ();
 sg13g2_fill_2 FILLER_76_89 ();
 sg13g2_fill_1 FILLER_76_117 ();
 sg13g2_fill_1 FILLER_76_128 ();
 sg13g2_fill_1 FILLER_76_139 ();
 sg13g2_fill_2 FILLER_76_150 ();
 sg13g2_fill_2 FILLER_76_156 ();
 sg13g2_decap_4 FILLER_76_171 ();
 sg13g2_fill_1 FILLER_76_175 ();
 sg13g2_fill_1 FILLER_76_224 ();
 sg13g2_fill_2 FILLER_76_250 ();
 sg13g2_fill_2 FILLER_76_256 ();
 sg13g2_decap_8 FILLER_76_325 ();
 sg13g2_decap_8 FILLER_76_332 ();
 sg13g2_decap_4 FILLER_76_354 ();
 sg13g2_fill_1 FILLER_76_358 ();
 sg13g2_fill_1 FILLER_76_366 ();
 sg13g2_decap_8 FILLER_76_372 ();
 sg13g2_decap_8 FILLER_76_379 ();
 sg13g2_decap_8 FILLER_76_386 ();
 sg13g2_fill_1 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_decap_8 FILLER_76_429 ();
 sg13g2_decap_8 FILLER_76_436 ();
 sg13g2_decap_8 FILLER_76_443 ();
 sg13g2_fill_1 FILLER_76_455 ();
 sg13g2_decap_4 FILLER_76_466 ();
 sg13g2_fill_2 FILLER_76_470 ();
 sg13g2_fill_1 FILLER_76_476 ();
 sg13g2_decap_4 FILLER_76_503 ();
 sg13g2_decap_4 FILLER_76_573 ();
 sg13g2_fill_2 FILLER_76_608 ();
 sg13g2_decap_8 FILLER_76_614 ();
 sg13g2_fill_2 FILLER_76_621 ();
 sg13g2_fill_1 FILLER_76_623 ();
 sg13g2_decap_4 FILLER_76_695 ();
 sg13g2_fill_2 FILLER_76_699 ();
 sg13g2_fill_1 FILLER_76_741 ();
 sg13g2_decap_4 FILLER_76_752 ();
 sg13g2_fill_2 FILLER_76_756 ();
 sg13g2_decap_8 FILLER_76_768 ();
 sg13g2_decap_8 FILLER_76_775 ();
 sg13g2_decap_4 FILLER_76_782 ();
 sg13g2_fill_1 FILLER_76_786 ();
 sg13g2_decap_8 FILLER_76_797 ();
 sg13g2_fill_1 FILLER_76_804 ();
 sg13g2_fill_2 FILLER_76_809 ();
 sg13g2_decap_8 FILLER_76_858 ();
 sg13g2_decap_8 FILLER_76_865 ();
 sg13g2_decap_4 FILLER_76_872 ();
 sg13g2_decap_4 FILLER_76_902 ();
 sg13g2_fill_1 FILLER_76_906 ();
 sg13g2_decap_8 FILLER_76_917 ();
 sg13g2_decap_8 FILLER_76_924 ();
 sg13g2_fill_1 FILLER_76_931 ();
 sg13g2_decap_8 FILLER_76_936 ();
 sg13g2_decap_8 FILLER_76_943 ();
 sg13g2_fill_1 FILLER_76_950 ();
 sg13g2_decap_8 FILLER_76_971 ();
 sg13g2_decap_8 FILLER_76_978 ();
 sg13g2_fill_1 FILLER_76_985 ();
 sg13g2_decap_8 FILLER_76_1022 ();
 sg13g2_decap_8 FILLER_76_1029 ();
 sg13g2_decap_8 FILLER_76_1036 ();
 sg13g2_decap_8 FILLER_76_1043 ();
 sg13g2_decap_8 FILLER_76_1050 ();
 sg13g2_decap_8 FILLER_76_1067 ();
 sg13g2_fill_2 FILLER_76_1074 ();
 sg13g2_decap_4 FILLER_76_1086 ();
 sg13g2_fill_1 FILLER_76_1090 ();
 sg13g2_decap_4 FILLER_76_1096 ();
 sg13g2_fill_1 FILLER_76_1100 ();
 sg13g2_fill_2 FILLER_76_1118 ();
 sg13g2_fill_2 FILLER_76_1135 ();
 sg13g2_fill_1 FILLER_76_1137 ();
 sg13g2_fill_2 FILLER_76_1148 ();
 sg13g2_decap_8 FILLER_76_1160 ();
 sg13g2_decap_8 FILLER_76_1167 ();
 sg13g2_decap_8 FILLER_76_1174 ();
 sg13g2_decap_8 FILLER_76_1185 ();
 sg13g2_decap_8 FILLER_76_1202 ();
 sg13g2_fill_2 FILLER_76_1209 ();
 sg13g2_fill_1 FILLER_76_1211 ();
 sg13g2_fill_1 FILLER_76_1216 ();
 sg13g2_decap_8 FILLER_76_1221 ();
 sg13g2_decap_8 FILLER_76_1228 ();
 sg13g2_decap_8 FILLER_76_1235 ();
 sg13g2_decap_8 FILLER_76_1242 ();
 sg13g2_decap_8 FILLER_76_1249 ();
 sg13g2_decap_8 FILLER_76_1256 ();
 sg13g2_decap_4 FILLER_76_1263 ();
 sg13g2_fill_1 FILLER_76_1297 ();
 sg13g2_fill_1 FILLER_76_1308 ();
 sg13g2_fill_2 FILLER_76_1335 ();
 sg13g2_fill_1 FILLER_76_1347 ();
 sg13g2_decap_8 FILLER_76_1358 ();
 sg13g2_decap_4 FILLER_76_1365 ();
 sg13g2_fill_1 FILLER_76_1395 ();
 sg13g2_fill_2 FILLER_76_1422 ();
 sg13g2_fill_1 FILLER_76_1424 ();
 sg13g2_decap_8 FILLER_76_1429 ();
 sg13g2_decap_8 FILLER_76_1436 ();
 sg13g2_decap_8 FILLER_76_1443 ();
 sg13g2_fill_1 FILLER_76_1450 ();
 sg13g2_decap_8 FILLER_76_1507 ();
 sg13g2_decap_8 FILLER_76_1514 ();
 sg13g2_fill_2 FILLER_76_1521 ();
 sg13g2_fill_1 FILLER_76_1559 ();
 sg13g2_fill_1 FILLER_76_1570 ();
 sg13g2_fill_1 FILLER_76_1581 ();
 sg13g2_fill_1 FILLER_76_1619 ();
 sg13g2_fill_1 FILLER_76_1646 ();
 sg13g2_decap_8 FILLER_76_1683 ();
 sg13g2_decap_8 FILLER_76_1690 ();
 sg13g2_decap_8 FILLER_76_1697 ();
 sg13g2_decap_4 FILLER_76_1704 ();
 sg13g2_decap_8 FILLER_76_1764 ();
 sg13g2_fill_2 FILLER_76_1771 ();
 sg13g2_fill_1 FILLER_76_1773 ();
 sg13g2_decap_4 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_4 ();
 sg13g2_fill_2 FILLER_77_19 ();
 sg13g2_fill_2 FILLER_77_57 ();
 sg13g2_fill_1 FILLER_77_59 ();
 sg13g2_fill_2 FILLER_77_86 ();
 sg13g2_fill_2 FILLER_77_114 ();
 sg13g2_decap_4 FILLER_77_126 ();
 sg13g2_decap_4 FILLER_77_140 ();
 sg13g2_fill_1 FILLER_77_191 ();
 sg13g2_fill_1 FILLER_77_205 ();
 sg13g2_fill_1 FILLER_77_287 ();
 sg13g2_fill_1 FILLER_77_298 ();
 sg13g2_fill_2 FILLER_77_315 ();
 sg13g2_fill_1 FILLER_77_321 ();
 sg13g2_fill_1 FILLER_77_350 ();
 sg13g2_decap_4 FILLER_77_365 ();
 sg13g2_fill_2 FILLER_77_369 ();
 sg13g2_decap_4 FILLER_77_412 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_448 ();
 sg13g2_fill_1 FILLER_77_455 ();
 sg13g2_fill_2 FILLER_77_492 ();
 sg13g2_fill_1 FILLER_77_494 ();
 sg13g2_decap_8 FILLER_77_550 ();
 sg13g2_decap_8 FILLER_77_577 ();
 sg13g2_decap_4 FILLER_77_584 ();
 sg13g2_fill_1 FILLER_77_588 ();
 sg13g2_decap_8 FILLER_77_625 ();
 sg13g2_decap_4 FILLER_77_632 ();
 sg13g2_fill_1 FILLER_77_636 ();
 sg13g2_fill_2 FILLER_77_693 ();
 sg13g2_fill_1 FILLER_77_695 ();
 sg13g2_decap_8 FILLER_77_700 ();
 sg13g2_decap_4 FILLER_77_707 ();
 sg13g2_decap_4 FILLER_77_715 ();
 sg13g2_fill_2 FILLER_77_750 ();
 sg13g2_fill_2 FILLER_77_778 ();
 sg13g2_fill_1 FILLER_77_805 ();
 sg13g2_fill_2 FILLER_77_816 ();
 sg13g2_fill_1 FILLER_77_818 ();
 sg13g2_decap_8 FILLER_77_865 ();
 sg13g2_fill_1 FILLER_77_872 ();
 sg13g2_fill_1 FILLER_77_887 ();
 sg13g2_decap_8 FILLER_77_940 ();
 sg13g2_fill_1 FILLER_77_947 ();
 sg13g2_decap_8 FILLER_77_974 ();
 sg13g2_fill_1 FILLER_77_995 ();
 sg13g2_decap_8 FILLER_77_1026 ();
 sg13g2_decap_4 FILLER_77_1033 ();
 sg13g2_fill_2 FILLER_77_1077 ();
 sg13g2_decap_4 FILLER_77_1084 ();
 sg13g2_fill_2 FILLER_77_1098 ();
 sg13g2_fill_2 FILLER_77_1120 ();
 sg13g2_fill_2 FILLER_77_1148 ();
 sg13g2_fill_2 FILLER_77_1154 ();
 sg13g2_fill_2 FILLER_77_1202 ();
 sg13g2_fill_1 FILLER_77_1204 ();
 sg13g2_decap_8 FILLER_77_1231 ();
 sg13g2_decap_4 FILLER_77_1238 ();
 sg13g2_fill_1 FILLER_77_1242 ();
 sg13g2_decap_4 FILLER_77_1269 ();
 sg13g2_fill_1 FILLER_77_1273 ();
 sg13g2_fill_2 FILLER_77_1284 ();
 sg13g2_decap_4 FILLER_77_1333 ();
 sg13g2_fill_1 FILLER_77_1337 ();
 sg13g2_decap_8 FILLER_77_1359 ();
 sg13g2_decap_8 FILLER_77_1366 ();
 sg13g2_fill_2 FILLER_77_1373 ();
 sg13g2_fill_1 FILLER_77_1375 ();
 sg13g2_decap_8 FILLER_77_1468 ();
 sg13g2_decap_8 FILLER_77_1475 ();
 sg13g2_fill_1 FILLER_77_1482 ();
 sg13g2_decap_4 FILLER_77_1517 ();
 sg13g2_fill_2 FILLER_77_1521 ();
 sg13g2_fill_1 FILLER_77_1533 ();
 sg13g2_fill_2 FILLER_77_1577 ();
 sg13g2_fill_2 FILLER_77_1622 ();
 sg13g2_fill_2 FILLER_77_1637 ();
 sg13g2_decap_4 FILLER_77_1698 ();
 sg13g2_fill_2 FILLER_77_1702 ();
 sg13g2_decap_8 FILLER_77_1748 ();
 sg13g2_decap_8 FILLER_77_1755 ();
 sg13g2_decap_8 FILLER_77_1762 ();
 sg13g2_decap_4 FILLER_77_1769 ();
 sg13g2_fill_1 FILLER_77_1773 ();
 sg13g2_decap_4 FILLER_78_0 ();
 sg13g2_decap_4 FILLER_78_34 ();
 sg13g2_fill_1 FILLER_78_106 ();
 sg13g2_fill_1 FILLER_78_141 ();
 sg13g2_fill_1 FILLER_78_168 ();
 sg13g2_fill_1 FILLER_78_179 ();
 sg13g2_fill_1 FILLER_78_206 ();
 sg13g2_fill_1 FILLER_78_211 ();
 sg13g2_fill_1 FILLER_78_231 ();
 sg13g2_fill_1 FILLER_78_245 ();
 sg13g2_fill_2 FILLER_78_275 ();
 sg13g2_decap_8 FILLER_78_432 ();
 sg13g2_decap_4 FILLER_78_439 ();
 sg13g2_fill_1 FILLER_78_443 ();
 sg13g2_decap_8 FILLER_78_495 ();
 sg13g2_fill_2 FILLER_78_502 ();
 sg13g2_fill_1 FILLER_78_530 ();
 sg13g2_fill_2 FILLER_78_567 ();
 sg13g2_fill_1 FILLER_78_595 ();
 sg13g2_fill_2 FILLER_78_606 ();
 sg13g2_fill_1 FILLER_78_634 ();
 sg13g2_fill_2 FILLER_78_661 ();
 sg13g2_decap_8 FILLER_78_699 ();
 sg13g2_decap_8 FILLER_78_706 ();
 sg13g2_decap_4 FILLER_78_713 ();
 sg13g2_fill_2 FILLER_78_789 ();
 sg13g2_fill_1 FILLER_78_817 ();
 sg13g2_fill_1 FILLER_78_828 ();
 sg13g2_fill_1 FILLER_78_855 ();
 sg13g2_fill_2 FILLER_78_882 ();
 sg13g2_fill_2 FILLER_78_924 ();
 sg13g2_fill_1 FILLER_78_952 ();
 sg13g2_fill_1 FILLER_78_979 ();
 sg13g2_fill_1 FILLER_78_990 ();
 sg13g2_decap_8 FILLER_78_1017 ();
 sg13g2_decap_8 FILLER_78_1024 ();
 sg13g2_decap_4 FILLER_78_1031 ();
 sg13g2_fill_2 FILLER_78_1035 ();
 sg13g2_fill_1 FILLER_78_1063 ();
 sg13g2_fill_1 FILLER_78_1068 ();
 sg13g2_fill_1 FILLER_78_1099 ();
 sg13g2_decap_4 FILLER_78_1105 ();
 sg13g2_fill_1 FILLER_78_1109 ();
 sg13g2_fill_2 FILLER_78_1170 ();
 sg13g2_fill_1 FILLER_78_1216 ();
 sg13g2_fill_2 FILLER_78_1227 ();
 sg13g2_fill_2 FILLER_78_1255 ();
 sg13g2_decap_8 FILLER_78_1283 ();
 sg13g2_fill_1 FILLER_78_1320 ();
 sg13g2_fill_2 FILLER_78_1397 ();
 sg13g2_decap_8 FILLER_78_1409 ();
 sg13g2_fill_1 FILLER_78_1416 ();
 sg13g2_decap_4 FILLER_78_1443 ();
 sg13g2_decap_8 FILLER_78_1473 ();
 sg13g2_fill_1 FILLER_78_1490 ();
 sg13g2_fill_1 FILLER_78_1495 ();
 sg13g2_fill_1 FILLER_78_1522 ();
 sg13g2_fill_1 FILLER_78_1559 ();
 sg13g2_fill_1 FILLER_78_1570 ();
 sg13g2_fill_2 FILLER_78_1645 ();
 sg13g2_fill_2 FILLER_78_1673 ();
 sg13g2_fill_2 FILLER_78_1679 ();
 sg13g2_fill_1 FILLER_78_1681 ();
 sg13g2_decap_4 FILLER_78_1692 ();
 sg13g2_fill_1 FILLER_78_1696 ();
 sg13g2_decap_4 FILLER_78_1701 ();
 sg13g2_fill_1 FILLER_78_1705 ();
 sg13g2_fill_2 FILLER_78_1716 ();
 sg13g2_fill_1 FILLER_78_1718 ();
 sg13g2_fill_1 FILLER_78_1723 ();
 sg13g2_decap_8 FILLER_78_1738 ();
 sg13g2_decap_8 FILLER_78_1745 ();
 sg13g2_decap_8 FILLER_78_1752 ();
 sg13g2_decap_8 FILLER_78_1759 ();
 sg13g2_decap_8 FILLER_78_1766 ();
 sg13g2_fill_1 FILLER_78_1773 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_9 ();
 sg13g2_fill_2 FILLER_79_40 ();
 sg13g2_fill_2 FILLER_79_94 ();
 sg13g2_fill_1 FILLER_79_96 ();
 sg13g2_fill_1 FILLER_79_101 ();
 sg13g2_fill_2 FILLER_79_131 ();
 sg13g2_fill_1 FILLER_79_133 ();
 sg13g2_fill_1 FILLER_79_211 ();
 sg13g2_fill_2 FILLER_79_219 ();
 sg13g2_fill_2 FILLER_79_230 ();
 sg13g2_fill_1 FILLER_79_238 ();
 sg13g2_fill_1 FILLER_79_304 ();
 sg13g2_fill_2 FILLER_79_324 ();
 sg13g2_fill_1 FILLER_79_330 ();
 sg13g2_fill_1 FILLER_79_336 ();
 sg13g2_fill_1 FILLER_79_376 ();
 sg13g2_decap_8 FILLER_79_449 ();
 sg13g2_decap_8 FILLER_79_456 ();
 sg13g2_fill_1 FILLER_79_463 ();
 sg13g2_fill_2 FILLER_79_469 ();
 sg13g2_fill_1 FILLER_79_471 ();
 sg13g2_fill_2 FILLER_79_545 ();
 sg13g2_fill_1 FILLER_79_547 ();
 sg13g2_decap_4 FILLER_79_560 ();
 sg13g2_fill_2 FILLER_79_590 ();
 sg13g2_fill_1 FILLER_79_592 ();
 sg13g2_fill_2 FILLER_79_629 ();
 sg13g2_fill_1 FILLER_79_641 ();
 sg13g2_fill_2 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_705 ();
 sg13g2_decap_8 FILLER_79_712 ();
 sg13g2_fill_2 FILLER_79_719 ();
 sg13g2_fill_2 FILLER_79_781 ();
 sg13g2_fill_1 FILLER_79_866 ();
 sg13g2_fill_1 FILLER_79_875 ();
 sg13g2_fill_1 FILLER_79_902 ();
 sg13g2_fill_1 FILLER_79_913 ();
 sg13g2_fill_1 FILLER_79_938 ();
 sg13g2_fill_1 FILLER_79_965 ();
 sg13g2_fill_1 FILLER_79_970 ();
 sg13g2_fill_1 FILLER_79_1023 ();
 sg13g2_fill_1 FILLER_79_1028 ();
 sg13g2_fill_2 FILLER_79_1033 ();
 sg13g2_fill_1 FILLER_79_1035 ();
 sg13g2_decap_4 FILLER_79_1086 ();
 sg13g2_fill_2 FILLER_79_1090 ();
 sg13g2_fill_1 FILLER_79_1118 ();
 sg13g2_decap_8 FILLER_79_1145 ();
 sg13g2_fill_2 FILLER_79_1152 ();
 sg13g2_fill_1 FILLER_79_1195 ();
 sg13g2_decap_4 FILLER_79_1226 ();
 sg13g2_fill_2 FILLER_79_1230 ();
 sg13g2_fill_1 FILLER_79_1236 ();
 sg13g2_fill_1 FILLER_79_1255 ();
 sg13g2_fill_2 FILLER_79_1266 ();
 sg13g2_fill_2 FILLER_79_1272 ();
 sg13g2_fill_2 FILLER_79_1279 ();
 sg13g2_fill_1 FILLER_79_1281 ();
 sg13g2_decap_8 FILLER_79_1300 ();
 sg13g2_decap_8 FILLER_79_1307 ();
 sg13g2_fill_2 FILLER_79_1314 ();
 sg13g2_fill_1 FILLER_79_1316 ();
 sg13g2_fill_2 FILLER_79_1353 ();
 sg13g2_fill_1 FILLER_79_1381 ();
 sg13g2_fill_2 FILLER_79_1386 ();
 sg13g2_fill_2 FILLER_79_1414 ();
 sg13g2_fill_2 FILLER_79_1442 ();
 sg13g2_fill_1 FILLER_79_1453 ();
 sg13g2_decap_4 FILLER_79_1458 ();
 sg13g2_decap_4 FILLER_79_1518 ();
 sg13g2_fill_1 FILLER_79_1522 ();
 sg13g2_fill_2 FILLER_79_1572 ();
 sg13g2_fill_1 FILLER_79_1578 ();
 sg13g2_fill_2 FILLER_79_1589 ();
 sg13g2_fill_2 FILLER_79_1595 ();
 sg13g2_fill_2 FILLER_79_1602 ();
 sg13g2_decap_4 FILLER_79_1634 ();
 sg13g2_decap_8 FILLER_79_1742 ();
 sg13g2_decap_8 FILLER_79_1749 ();
 sg13g2_decap_8 FILLER_79_1756 ();
 sg13g2_decap_8 FILLER_79_1763 ();
 sg13g2_decap_4 FILLER_79_1770 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_4 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_22 ();
 sg13g2_decap_8 FILLER_80_29 ();
 sg13g2_decap_8 FILLER_80_36 ();
 sg13g2_decap_8 FILLER_80_43 ();
 sg13g2_decap_8 FILLER_80_50 ();
 sg13g2_fill_1 FILLER_80_57 ();
 sg13g2_fill_1 FILLER_80_92 ();
 sg13g2_fill_1 FILLER_80_215 ();
 sg13g2_fill_1 FILLER_80_279 ();
 sg13g2_decap_4 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_369 ();
 sg13g2_fill_1 FILLER_80_411 ();
 sg13g2_fill_1 FILLER_80_416 ();
 sg13g2_decap_8 FILLER_80_434 ();
 sg13g2_decap_8 FILLER_80_441 ();
 sg13g2_decap_8 FILLER_80_448 ();
 sg13g2_decap_8 FILLER_80_455 ();
 sg13g2_fill_2 FILLER_80_462 ();
 sg13g2_decap_4 FILLER_80_474 ();
 sg13g2_fill_2 FILLER_80_478 ();
 sg13g2_fill_2 FILLER_80_484 ();
 sg13g2_decap_8 FILLER_80_496 ();
 sg13g2_decap_8 FILLER_80_507 ();
 sg13g2_fill_1 FILLER_80_514 ();
 sg13g2_decap_8 FILLER_80_523 ();
 sg13g2_fill_1 FILLER_80_530 ();
 sg13g2_decap_4 FILLER_80_561 ();
 sg13g2_fill_1 FILLER_80_565 ();
 sg13g2_fill_2 FILLER_80_570 ();
 sg13g2_fill_1 FILLER_80_572 ();
 sg13g2_fill_1 FILLER_80_581 ();
 sg13g2_decap_8 FILLER_80_587 ();
 sg13g2_decap_8 FILLER_80_594 ();
 sg13g2_decap_8 FILLER_80_601 ();
 sg13g2_decap_4 FILLER_80_608 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_632 ();
 sg13g2_decap_8 FILLER_80_639 ();
 sg13g2_decap_4 FILLER_80_646 ();
 sg13g2_fill_2 FILLER_80_650 ();
 sg13g2_decap_4 FILLER_80_656 ();
 sg13g2_fill_2 FILLER_80_660 ();
 sg13g2_fill_2 FILLER_80_672 ();
 sg13g2_fill_2 FILLER_80_678 ();
 sg13g2_fill_1 FILLER_80_680 ();
 sg13g2_fill_2 FILLER_80_685 ();
 sg13g2_fill_1 FILLER_80_687 ();
 sg13g2_fill_2 FILLER_80_692 ();
 sg13g2_fill_1 FILLER_80_694 ();
 sg13g2_decap_8 FILLER_80_699 ();
 sg13g2_decap_8 FILLER_80_706 ();
 sg13g2_decap_8 FILLER_80_713 ();
 sg13g2_decap_8 FILLER_80_720 ();
 sg13g2_fill_2 FILLER_80_727 ();
 sg13g2_decap_4 FILLER_80_743 ();
 sg13g2_fill_1 FILLER_80_747 ();
 sg13g2_fill_2 FILLER_80_758 ();
 sg13g2_fill_1 FILLER_80_760 ();
 sg13g2_fill_2 FILLER_80_765 ();
 sg13g2_fill_2 FILLER_80_771 ();
 sg13g2_fill_1 FILLER_80_773 ();
 sg13g2_fill_2 FILLER_80_778 ();
 sg13g2_decap_4 FILLER_80_784 ();
 sg13g2_fill_2 FILLER_80_788 ();
 sg13g2_fill_2 FILLER_80_794 ();
 sg13g2_fill_1 FILLER_80_796 ();
 sg13g2_decap_8 FILLER_80_801 ();
 sg13g2_decap_8 FILLER_80_808 ();
 sg13g2_decap_8 FILLER_80_815 ();
 sg13g2_decap_4 FILLER_80_822 ();
 sg13g2_fill_2 FILLER_80_834 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_fill_1 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_852 ();
 sg13g2_decap_4 FILLER_80_859 ();
 sg13g2_fill_1 FILLER_80_863 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_decap_4 FILLER_80_875 ();
 sg13g2_fill_1 FILLER_80_879 ();
 sg13g2_decap_4 FILLER_80_889 ();
 sg13g2_fill_1 FILLER_80_893 ();
 sg13g2_fill_2 FILLER_80_898 ();
 sg13g2_decap_4 FILLER_80_909 ();
 sg13g2_decap_8 FILLER_80_921 ();
 sg13g2_decap_4 FILLER_80_928 ();
 sg13g2_decap_4 FILLER_80_942 ();
 sg13g2_fill_2 FILLER_80_950 ();
 sg13g2_decap_8 FILLER_80_966 ();
 sg13g2_decap_4 FILLER_80_973 ();
 sg13g2_fill_1 FILLER_80_977 ();
 sg13g2_decap_8 FILLER_80_982 ();
 sg13g2_decap_8 FILLER_80_989 ();
 sg13g2_fill_2 FILLER_80_996 ();
 sg13g2_decap_4 FILLER_80_1002 ();
 sg13g2_decap_4 FILLER_80_1010 ();
 sg13g2_fill_1 FILLER_80_1014 ();
 sg13g2_decap_8 FILLER_80_1020 ();
 sg13g2_decap_8 FILLER_80_1027 ();
 sg13g2_decap_8 FILLER_80_1034 ();
 sg13g2_fill_2 FILLER_80_1041 ();
 sg13g2_fill_1 FILLER_80_1043 ();
 sg13g2_decap_4 FILLER_80_1048 ();
 sg13g2_decap_8 FILLER_80_1057 ();
 sg13g2_decap_4 FILLER_80_1064 ();
 sg13g2_decap_8 FILLER_80_1094 ();
 sg13g2_decap_8 FILLER_80_1105 ();
 sg13g2_decap_4 FILLER_80_1112 ();
 sg13g2_fill_2 FILLER_80_1116 ();
 sg13g2_decap_8 FILLER_80_1130 ();
 sg13g2_decap_8 FILLER_80_1137 ();
 sg13g2_decap_8 FILLER_80_1144 ();
 sg13g2_decap_8 FILLER_80_1151 ();
 sg13g2_decap_4 FILLER_80_1158 ();
 sg13g2_decap_8 FILLER_80_1170 ();
 sg13g2_decap_8 FILLER_80_1177 ();
 sg13g2_decap_8 FILLER_80_1184 ();
 sg13g2_fill_2 FILLER_80_1191 ();
 sg13g2_fill_1 FILLER_80_1193 ();
 sg13g2_decap_8 FILLER_80_1228 ();
 sg13g2_decap_8 FILLER_80_1235 ();
 sg13g2_decap_8 FILLER_80_1242 ();
 sg13g2_decap_8 FILLER_80_1249 ();
 sg13g2_decap_8 FILLER_80_1256 ();
 sg13g2_decap_8 FILLER_80_1263 ();
 sg13g2_decap_8 FILLER_80_1270 ();
 sg13g2_decap_8 FILLER_80_1277 ();
 sg13g2_fill_1 FILLER_80_1284 ();
 sg13g2_decap_8 FILLER_80_1311 ();
 sg13g2_decap_8 FILLER_80_1318 ();
 sg13g2_decap_4 FILLER_80_1325 ();
 sg13g2_fill_1 FILLER_80_1329 ();
 sg13g2_decap_4 FILLER_80_1342 ();
 sg13g2_fill_1 FILLER_80_1346 ();
 sg13g2_decap_4 FILLER_80_1352 ();
 sg13g2_fill_2 FILLER_80_1356 ();
 sg13g2_fill_2 FILLER_80_1366 ();
 sg13g2_decap_8 FILLER_80_1377 ();
 sg13g2_fill_2 FILLER_80_1384 ();
 sg13g2_decap_8 FILLER_80_1400 ();
 sg13g2_decap_4 FILLER_80_1407 ();
 sg13g2_fill_1 FILLER_80_1411 ();
 sg13g2_fill_1 FILLER_80_1422 ();
 sg13g2_fill_2 FILLER_80_1427 ();
 sg13g2_fill_2 FILLER_80_1433 ();
 sg13g2_decap_8 FILLER_80_1439 ();
 sg13g2_decap_8 FILLER_80_1446 ();
 sg13g2_decap_8 FILLER_80_1453 ();
 sg13g2_decap_8 FILLER_80_1460 ();
 sg13g2_fill_1 FILLER_80_1467 ();
 sg13g2_decap_8 FILLER_80_1472 ();
 sg13g2_decap_4 FILLER_80_1479 ();
 sg13g2_fill_2 FILLER_80_1483 ();
 sg13g2_decap_4 FILLER_80_1490 ();
 sg13g2_fill_1 FILLER_80_1494 ();
 sg13g2_decap_4 FILLER_80_1499 ();
 sg13g2_decap_4 FILLER_80_1529 ();
 sg13g2_fill_2 FILLER_80_1533 ();
 sg13g2_fill_1 FILLER_80_1558 ();
 sg13g2_decap_8 FILLER_80_1600 ();
 sg13g2_decap_4 FILLER_80_1607 ();
 sg13g2_fill_2 FILLER_80_1611 ();
 sg13g2_decap_8 FILLER_80_1626 ();
 sg13g2_decap_8 FILLER_80_1633 ();
 sg13g2_decap_4 FILLER_80_1640 ();
 sg13g2_decap_4 FILLER_80_1648 ();
 sg13g2_fill_1 FILLER_80_1656 ();
 sg13g2_decap_8 FILLER_80_1661 ();
 sg13g2_fill_2 FILLER_80_1668 ();
 sg13g2_fill_1 FILLER_80_1670 ();
 sg13g2_fill_2 FILLER_80_1675 ();
 sg13g2_fill_1 FILLER_80_1677 ();
 sg13g2_decap_8 FILLER_80_1683 ();
 sg13g2_decap_8 FILLER_80_1690 ();
 sg13g2_fill_2 FILLER_80_1697 ();
 sg13g2_fill_1 FILLER_80_1699 ();
 sg13g2_decap_8 FILLER_80_1705 ();
 sg13g2_decap_8 FILLER_80_1712 ();
 sg13g2_decap_4 FILLER_80_1719 ();
 sg13g2_fill_1 FILLER_80_1723 ();
 sg13g2_decap_8 FILLER_80_1728 ();
 sg13g2_decap_8 FILLER_80_1735 ();
 sg13g2_decap_8 FILLER_80_1742 ();
 sg13g2_decap_8 FILLER_80_1749 ();
 sg13g2_decap_8 FILLER_80_1756 ();
 sg13g2_decap_8 FILLER_80_1763 ();
 sg13g2_decap_4 FILLER_80_1770 ();
endmodule
