module tt_um_simon_cipher (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire clknet_leaf_0_clk;
 wire net100;
 wire \bitserial_cipher.bit_counter[0] ;
 wire \bitserial_cipher.bit_counter[1] ;
 wire \bitserial_cipher.bit_counter[2] ;
 wire \bitserial_cipher.bit_counter[3] ;
 wire \bitserial_cipher.bit_counter[4] ;
 wire \bitserial_cipher.bit_counter[5] ;
 wire \bitserial_cipher.cipher_out ;
 wire \bitserial_cipher.datapath.fifo_ff56 ;
 wire \bitserial_cipher.datapath.fifo_ff57 ;
 wire \bitserial_cipher.datapath.fifo_ff58 ;
 wire \bitserial_cipher.datapath.fifo_ff59 ;
 wire \bitserial_cipher.datapath.fifo_ff60 ;
 wire \bitserial_cipher.datapath.fifo_ff61 ;
 wire \bitserial_cipher.datapath.fifo_ff62 ;
 wire \bitserial_cipher.datapath.fifo_ff63 ;
 wire \bitserial_cipher.datapath.key_in ;
 wire \bitserial_cipher.datapath.lut_ff56 ;
 wire \bitserial_cipher.datapath.lut_ff57 ;
 wire \bitserial_cipher.datapath.lut_ff58 ;
 wire \bitserial_cipher.datapath.lut_ff59 ;
 wire \bitserial_cipher.datapath.lut_ff60 ;
 wire \bitserial_cipher.datapath.lut_ff61 ;
 wire \bitserial_cipher.datapath.lut_ff62 ;
 wire \bitserial_cipher.datapath.lut_ff63 ;
 wire \bitserial_cipher.datapath.round_counter[0] ;
 wire \bitserial_cipher.datapath.round_counter[1] ;
 wire \bitserial_cipher.datapath.round_counter[2] ;
 wire \bitserial_cipher.datapath.round_counter[3] ;
 wire \bitserial_cipher.datapath.round_counter[4] ;
 wire \bitserial_cipher.datapath.round_counter[5] ;
 wire \bitserial_cipher.datapath.round_counter[6] ;
 wire \bitserial_cipher.datapath.shift_in2 ;
 wire \bitserial_cipher.datapath.shifter1[10] ;
 wire \bitserial_cipher.datapath.shifter1[11] ;
 wire \bitserial_cipher.datapath.shifter1[12] ;
 wire \bitserial_cipher.datapath.shifter1[13] ;
 wire \bitserial_cipher.datapath.shifter1[14] ;
 wire \bitserial_cipher.datapath.shifter1[15] ;
 wire \bitserial_cipher.datapath.shifter1[16] ;
 wire \bitserial_cipher.datapath.shifter1[17] ;
 wire \bitserial_cipher.datapath.shifter1[18] ;
 wire \bitserial_cipher.datapath.shifter1[19] ;
 wire \bitserial_cipher.datapath.shifter1[1] ;
 wire \bitserial_cipher.datapath.shifter1[20] ;
 wire \bitserial_cipher.datapath.shifter1[21] ;
 wire \bitserial_cipher.datapath.shifter1[22] ;
 wire \bitserial_cipher.datapath.shifter1[23] ;
 wire \bitserial_cipher.datapath.shifter1[24] ;
 wire \bitserial_cipher.datapath.shifter1[25] ;
 wire \bitserial_cipher.datapath.shifter1[26] ;
 wire \bitserial_cipher.datapath.shifter1[27] ;
 wire \bitserial_cipher.datapath.shifter1[28] ;
 wire \bitserial_cipher.datapath.shifter1[29] ;
 wire \bitserial_cipher.datapath.shifter1[2] ;
 wire \bitserial_cipher.datapath.shifter1[30] ;
 wire \bitserial_cipher.datapath.shifter1[31] ;
 wire \bitserial_cipher.datapath.shifter1[32] ;
 wire \bitserial_cipher.datapath.shifter1[33] ;
 wire \bitserial_cipher.datapath.shifter1[34] ;
 wire \bitserial_cipher.datapath.shifter1[35] ;
 wire \bitserial_cipher.datapath.shifter1[36] ;
 wire \bitserial_cipher.datapath.shifter1[37] ;
 wire \bitserial_cipher.datapath.shifter1[38] ;
 wire \bitserial_cipher.datapath.shifter1[39] ;
 wire \bitserial_cipher.datapath.shifter1[3] ;
 wire \bitserial_cipher.datapath.shifter1[40] ;
 wire \bitserial_cipher.datapath.shifter1[41] ;
 wire \bitserial_cipher.datapath.shifter1[42] ;
 wire \bitserial_cipher.datapath.shifter1[43] ;
 wire \bitserial_cipher.datapath.shifter1[44] ;
 wire \bitserial_cipher.datapath.shifter1[45] ;
 wire \bitserial_cipher.datapath.shifter1[46] ;
 wire \bitserial_cipher.datapath.shifter1[47] ;
 wire \bitserial_cipher.datapath.shifter1[48] ;
 wire \bitserial_cipher.datapath.shifter1[49] ;
 wire \bitserial_cipher.datapath.shifter1[4] ;
 wire \bitserial_cipher.datapath.shifter1[50] ;
 wire \bitserial_cipher.datapath.shifter1[51] ;
 wire \bitserial_cipher.datapath.shifter1[52] ;
 wire \bitserial_cipher.datapath.shifter1[53] ;
 wire \bitserial_cipher.datapath.shifter1[54] ;
 wire \bitserial_cipher.datapath.shifter1[55] ;
 wire \bitserial_cipher.datapath.shifter1[5] ;
 wire \bitserial_cipher.datapath.shifter1[6] ;
 wire \bitserial_cipher.datapath.shifter1[7] ;
 wire \bitserial_cipher.datapath.shifter1[8] ;
 wire \bitserial_cipher.datapath.shifter1[9] ;
 wire \bitserial_cipher.datapath.shifter2[10] ;
 wire \bitserial_cipher.datapath.shifter2[11] ;
 wire \bitserial_cipher.datapath.shifter2[12] ;
 wire \bitserial_cipher.datapath.shifter2[13] ;
 wire \bitserial_cipher.datapath.shifter2[14] ;
 wire \bitserial_cipher.datapath.shifter2[15] ;
 wire \bitserial_cipher.datapath.shifter2[16] ;
 wire \bitserial_cipher.datapath.shifter2[17] ;
 wire \bitserial_cipher.datapath.shifter2[18] ;
 wire \bitserial_cipher.datapath.shifter2[19] ;
 wire \bitserial_cipher.datapath.shifter2[1] ;
 wire \bitserial_cipher.datapath.shifter2[20] ;
 wire \bitserial_cipher.datapath.shifter2[21] ;
 wire \bitserial_cipher.datapath.shifter2[22] ;
 wire \bitserial_cipher.datapath.shifter2[23] ;
 wire \bitserial_cipher.datapath.shifter2[24] ;
 wire \bitserial_cipher.datapath.shifter2[25] ;
 wire \bitserial_cipher.datapath.shifter2[26] ;
 wire \bitserial_cipher.datapath.shifter2[27] ;
 wire \bitserial_cipher.datapath.shifter2[28] ;
 wire \bitserial_cipher.datapath.shifter2[29] ;
 wire \bitserial_cipher.datapath.shifter2[2] ;
 wire \bitserial_cipher.datapath.shifter2[30] ;
 wire \bitserial_cipher.datapath.shifter2[31] ;
 wire \bitserial_cipher.datapath.shifter2[32] ;
 wire \bitserial_cipher.datapath.shifter2[33] ;
 wire \bitserial_cipher.datapath.shifter2[34] ;
 wire \bitserial_cipher.datapath.shifter2[35] ;
 wire \bitserial_cipher.datapath.shifter2[36] ;
 wire \bitserial_cipher.datapath.shifter2[37] ;
 wire \bitserial_cipher.datapath.shifter2[38] ;
 wire \bitserial_cipher.datapath.shifter2[39] ;
 wire \bitserial_cipher.datapath.shifter2[3] ;
 wire \bitserial_cipher.datapath.shifter2[40] ;
 wire \bitserial_cipher.datapath.shifter2[41] ;
 wire \bitserial_cipher.datapath.shifter2[42] ;
 wire \bitserial_cipher.datapath.shifter2[43] ;
 wire \bitserial_cipher.datapath.shifter2[44] ;
 wire \bitserial_cipher.datapath.shifter2[45] ;
 wire \bitserial_cipher.datapath.shifter2[46] ;
 wire \bitserial_cipher.datapath.shifter2[47] ;
 wire \bitserial_cipher.datapath.shifter2[48] ;
 wire \bitserial_cipher.datapath.shifter2[49] ;
 wire \bitserial_cipher.datapath.shifter2[4] ;
 wire \bitserial_cipher.datapath.shifter2[50] ;
 wire \bitserial_cipher.datapath.shifter2[51] ;
 wire \bitserial_cipher.datapath.shifter2[52] ;
 wire \bitserial_cipher.datapath.shifter2[53] ;
 wire \bitserial_cipher.datapath.shifter2[54] ;
 wire \bitserial_cipher.datapath.shifter2[55] ;
 wire \bitserial_cipher.datapath.shifter2[56] ;
 wire \bitserial_cipher.datapath.shifter2[57] ;
 wire \bitserial_cipher.datapath.shifter2[58] ;
 wire \bitserial_cipher.datapath.shifter2[59] ;
 wire \bitserial_cipher.datapath.shifter2[5] ;
 wire \bitserial_cipher.datapath.shifter2[60] ;
 wire \bitserial_cipher.datapath.shifter2[61] ;
 wire \bitserial_cipher.datapath.shifter2[62] ;
 wire \bitserial_cipher.datapath.shifter2[63] ;
 wire \bitserial_cipher.datapath.shifter2[6] ;
 wire \bitserial_cipher.datapath.shifter2[7] ;
 wire \bitserial_cipher.datapath.shifter2[8] ;
 wire \bitserial_cipher.datapath.shifter2[9] ;
 wire \bitserial_cipher.datapath.valid ;
 wire \bitserial_cipher.key_exp.fifo_ff0 ;
 wire \bitserial_cipher.key_exp.fifo_ff1 ;
 wire \bitserial_cipher.key_exp.fifo_ff2 ;
 wire \bitserial_cipher.key_exp.fifo_ff3 ;
 wire \bitserial_cipher.key_exp.lut_ff0 ;
 wire \bitserial_cipher.key_exp.lut_ff1 ;
 wire \bitserial_cipher.key_exp.lut_ff2 ;
 wire \bitserial_cipher.key_exp.lut_ff3 ;
 wire \bitserial_cipher.key_exp.shift_out1 ;
 wire \bitserial_cipher.key_exp.shifter1[10] ;
 wire \bitserial_cipher.key_exp.shifter1[11] ;
 wire \bitserial_cipher.key_exp.shifter1[12] ;
 wire \bitserial_cipher.key_exp.shifter1[13] ;
 wire \bitserial_cipher.key_exp.shifter1[14] ;
 wire \bitserial_cipher.key_exp.shifter1[15] ;
 wire \bitserial_cipher.key_exp.shifter1[16] ;
 wire \bitserial_cipher.key_exp.shifter1[17] ;
 wire \bitserial_cipher.key_exp.shifter1[18] ;
 wire \bitserial_cipher.key_exp.shifter1[19] ;
 wire \bitserial_cipher.key_exp.shifter1[1] ;
 wire \bitserial_cipher.key_exp.shifter1[20] ;
 wire \bitserial_cipher.key_exp.shifter1[21] ;
 wire \bitserial_cipher.key_exp.shifter1[22] ;
 wire \bitserial_cipher.key_exp.shifter1[23] ;
 wire \bitserial_cipher.key_exp.shifter1[24] ;
 wire \bitserial_cipher.key_exp.shifter1[25] ;
 wire \bitserial_cipher.key_exp.shifter1[26] ;
 wire \bitserial_cipher.key_exp.shifter1[27] ;
 wire \bitserial_cipher.key_exp.shifter1[28] ;
 wire \bitserial_cipher.key_exp.shifter1[29] ;
 wire \bitserial_cipher.key_exp.shifter1[2] ;
 wire \bitserial_cipher.key_exp.shifter1[30] ;
 wire \bitserial_cipher.key_exp.shifter1[31] ;
 wire \bitserial_cipher.key_exp.shifter1[32] ;
 wire \bitserial_cipher.key_exp.shifter1[33] ;
 wire \bitserial_cipher.key_exp.shifter1[34] ;
 wire \bitserial_cipher.key_exp.shifter1[35] ;
 wire \bitserial_cipher.key_exp.shifter1[36] ;
 wire \bitserial_cipher.key_exp.shifter1[37] ;
 wire \bitserial_cipher.key_exp.shifter1[38] ;
 wire \bitserial_cipher.key_exp.shifter1[39] ;
 wire \bitserial_cipher.key_exp.shifter1[3] ;
 wire \bitserial_cipher.key_exp.shifter1[40] ;
 wire \bitserial_cipher.key_exp.shifter1[41] ;
 wire \bitserial_cipher.key_exp.shifter1[42] ;
 wire \bitserial_cipher.key_exp.shifter1[43] ;
 wire \bitserial_cipher.key_exp.shifter1[44] ;
 wire \bitserial_cipher.key_exp.shifter1[45] ;
 wire \bitserial_cipher.key_exp.shifter1[46] ;
 wire \bitserial_cipher.key_exp.shifter1[47] ;
 wire \bitserial_cipher.key_exp.shifter1[48] ;
 wire \bitserial_cipher.key_exp.shifter1[49] ;
 wire \bitserial_cipher.key_exp.shifter1[4] ;
 wire \bitserial_cipher.key_exp.shifter1[50] ;
 wire \bitserial_cipher.key_exp.shifter1[51] ;
 wire \bitserial_cipher.key_exp.shifter1[52] ;
 wire \bitserial_cipher.key_exp.shifter1[53] ;
 wire \bitserial_cipher.key_exp.shifter1[54] ;
 wire \bitserial_cipher.key_exp.shifter1[55] ;
 wire \bitserial_cipher.key_exp.shifter1[56] ;
 wire \bitserial_cipher.key_exp.shifter1[57] ;
 wire \bitserial_cipher.key_exp.shifter1[58] ;
 wire \bitserial_cipher.key_exp.shifter1[59] ;
 wire \bitserial_cipher.key_exp.shifter1[5] ;
 wire \bitserial_cipher.key_exp.shifter1[6] ;
 wire \bitserial_cipher.key_exp.shifter1[7] ;
 wire \bitserial_cipher.key_exp.shifter1[8] ;
 wire \bitserial_cipher.key_exp.shifter1[9] ;
 wire \bitserial_cipher.key_exp.shifter2[10] ;
 wire \bitserial_cipher.key_exp.shifter2[11] ;
 wire \bitserial_cipher.key_exp.shifter2[12] ;
 wire \bitserial_cipher.key_exp.shifter2[13] ;
 wire \bitserial_cipher.key_exp.shifter2[14] ;
 wire \bitserial_cipher.key_exp.shifter2[15] ;
 wire \bitserial_cipher.key_exp.shifter2[16] ;
 wire \bitserial_cipher.key_exp.shifter2[17] ;
 wire \bitserial_cipher.key_exp.shifter2[18] ;
 wire \bitserial_cipher.key_exp.shifter2[19] ;
 wire \bitserial_cipher.key_exp.shifter2[1] ;
 wire \bitserial_cipher.key_exp.shifter2[20] ;
 wire \bitserial_cipher.key_exp.shifter2[21] ;
 wire \bitserial_cipher.key_exp.shifter2[22] ;
 wire \bitserial_cipher.key_exp.shifter2[23] ;
 wire \bitserial_cipher.key_exp.shifter2[24] ;
 wire \bitserial_cipher.key_exp.shifter2[25] ;
 wire \bitserial_cipher.key_exp.shifter2[26] ;
 wire \bitserial_cipher.key_exp.shifter2[27] ;
 wire \bitserial_cipher.key_exp.shifter2[28] ;
 wire \bitserial_cipher.key_exp.shifter2[29] ;
 wire \bitserial_cipher.key_exp.shifter2[2] ;
 wire \bitserial_cipher.key_exp.shifter2[30] ;
 wire \bitserial_cipher.key_exp.shifter2[31] ;
 wire \bitserial_cipher.key_exp.shifter2[32] ;
 wire \bitserial_cipher.key_exp.shifter2[33] ;
 wire \bitserial_cipher.key_exp.shifter2[34] ;
 wire \bitserial_cipher.key_exp.shifter2[35] ;
 wire \bitserial_cipher.key_exp.shifter2[36] ;
 wire \bitserial_cipher.key_exp.shifter2[37] ;
 wire \bitserial_cipher.key_exp.shifter2[38] ;
 wire \bitserial_cipher.key_exp.shifter2[39] ;
 wire \bitserial_cipher.key_exp.shifter2[3] ;
 wire \bitserial_cipher.key_exp.shifter2[40] ;
 wire \bitserial_cipher.key_exp.shifter2[41] ;
 wire \bitserial_cipher.key_exp.shifter2[42] ;
 wire \bitserial_cipher.key_exp.shifter2[43] ;
 wire \bitserial_cipher.key_exp.shifter2[44] ;
 wire \bitserial_cipher.key_exp.shifter2[45] ;
 wire \bitserial_cipher.key_exp.shifter2[46] ;
 wire \bitserial_cipher.key_exp.shifter2[47] ;
 wire \bitserial_cipher.key_exp.shifter2[48] ;
 wire \bitserial_cipher.key_exp.shifter2[49] ;
 wire \bitserial_cipher.key_exp.shifter2[4] ;
 wire \bitserial_cipher.key_exp.shifter2[50] ;
 wire \bitserial_cipher.key_exp.shifter2[51] ;
 wire \bitserial_cipher.key_exp.shifter2[52] ;
 wire \bitserial_cipher.key_exp.shifter2[53] ;
 wire \bitserial_cipher.key_exp.shifter2[54] ;
 wire \bitserial_cipher.key_exp.shifter2[55] ;
 wire \bitserial_cipher.key_exp.shifter2[56] ;
 wire \bitserial_cipher.key_exp.shifter2[57] ;
 wire \bitserial_cipher.key_exp.shifter2[58] ;
 wire \bitserial_cipher.key_exp.shifter2[59] ;
 wire \bitserial_cipher.key_exp.shifter2[5] ;
 wire \bitserial_cipher.key_exp.shifter2[60] ;
 wire \bitserial_cipher.key_exp.shifter2[61] ;
 wire \bitserial_cipher.key_exp.shifter2[62] ;
 wire \bitserial_cipher.key_exp.shifter2[63] ;
 wire \bitserial_cipher.key_exp.shifter2[6] ;
 wire \bitserial_cipher.key_exp.shifter2[7] ;
 wire \bitserial_cipher.key_exp.shifter2[8] ;
 wire \bitserial_cipher.key_exp.shifter2[9] ;
 wire \bitserial_cipher.zero ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_1 _1099_ (.A(ui_in[6]),
    .X(_0543_));
 sg13g2_buf_1 _1100_ (.A(_0543_),
    .X(_0544_));
 sg13g2_buf_1 _1101_ (.A(_0544_),
    .X(_0545_));
 sg13g2_buf_2 _1102_ (.A(ui_in[7]),
    .X(_0546_));
 sg13g2_buf_1 _1103_ (.A(_0546_),
    .X(_0547_));
 sg13g2_inv_1 _1104_ (.Y(_0548_),
    .A(\bitserial_cipher.bit_counter[0] ));
 sg13g2_nand2_1 _1105_ (.Y(_0549_),
    .A(net73),
    .B(_0004_));
 sg13g2_o21ai_1 _1106_ (.B1(_0549_),
    .Y(_0550_),
    .A1(net73),
    .A2(_0548_));
 sg13g2_nand2_1 _1107_ (.Y(_0551_),
    .A(net73),
    .B(\bitserial_cipher.bit_counter[0] ));
 sg13g2_nor2_1 _1108_ (.A(_0545_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_a21oi_1 _1109_ (.A1(_0545_),
    .A2(_0550_),
    .Y(_0553_),
    .B1(_0552_));
 sg13g2_buf_1 _1110_ (.A(net1),
    .X(_0554_));
 sg13g2_buf_1 _1111_ (.A(net75),
    .X(_0555_));
 sg13g2_buf_1 _1112_ (.A(net72),
    .X(_0556_));
 sg13g2_nor2b_1 _1113_ (.A(_0553_),
    .B_N(net47),
    .Y(_0005_));
 sg13g2_buf_1 _1114_ (.A(_0546_),
    .X(_0557_));
 sg13g2_buf_1 _1115_ (.A(_0557_),
    .X(_0558_));
 sg13g2_buf_1 _1116_ (.A(net76),
    .X(_0559_));
 sg13g2_inv_2 _1117_ (.Y(_0560_),
    .A(\bitserial_cipher.bit_counter[1] ));
 sg13g2_nand3_1 _1118_ (.B(\bitserial_cipher.bit_counter[0] ),
    .C(_0560_),
    .A(net70),
    .Y(_0561_));
 sg13g2_o21ai_1 _1119_ (.B1(_0561_),
    .Y(_0562_),
    .A1(net70),
    .A2(_0560_));
 sg13g2_and2_1 _1120_ (.A(_0559_),
    .B(\bitserial_cipher.bit_counter[1] ),
    .X(_0563_));
 sg13g2_a22oi_1 _1121_ (.Y(_0564_),
    .B1(_0563_),
    .B2(_0551_),
    .A2(_0562_),
    .A1(net46));
 sg13g2_nor2b_1 _1122_ (.A(_0564_),
    .B_N(net47),
    .Y(_0006_));
 sg13g2_inv_1 _1123_ (.Y(_0565_),
    .A(\bitserial_cipher.bit_counter[2] ));
 sg13g2_nor2_1 _1124_ (.A(_0548_),
    .B(_0560_),
    .Y(_0566_));
 sg13g2_nand3_1 _1125_ (.B(_0565_),
    .C(_0566_),
    .A(net70),
    .Y(_0567_));
 sg13g2_o21ai_1 _1126_ (.B1(_0567_),
    .Y(_0568_),
    .A1(net70),
    .A2(_0565_));
 sg13g2_nand3_1 _1127_ (.B(\bitserial_cipher.bit_counter[0] ),
    .C(\bitserial_cipher.bit_counter[1] ),
    .A(_0546_),
    .Y(_0569_));
 sg13g2_and2_1 _1128_ (.A(net48),
    .B(\bitserial_cipher.bit_counter[2] ),
    .X(_0570_));
 sg13g2_a22oi_1 _1129_ (.Y(_0571_),
    .B1(_0569_),
    .B2(_0570_),
    .A2(_0568_),
    .A1(net46));
 sg13g2_nor2b_1 _1130_ (.A(_0571_),
    .B_N(net47),
    .Y(_0007_));
 sg13g2_inv_1 _1131_ (.Y(_0572_),
    .A(\bitserial_cipher.bit_counter[3] ));
 sg13g2_nand4_1 _1132_ (.B(_0572_),
    .C(\bitserial_cipher.bit_counter[2] ),
    .A(_0544_),
    .Y(_0573_),
    .D(_0566_));
 sg13g2_o21ai_1 _1133_ (.B1(_0573_),
    .Y(_0574_),
    .A1(net70),
    .A2(_0572_));
 sg13g2_and2_1 _1134_ (.A(net70),
    .B(\bitserial_cipher.bit_counter[3] ),
    .X(_0575_));
 sg13g2_or2_1 _1135_ (.X(_0576_),
    .B(_0569_),
    .A(_0565_));
 sg13g2_a22oi_1 _1136_ (.Y(_0577_),
    .B1(_0575_),
    .B2(_0576_),
    .A2(_0574_),
    .A1(net46));
 sg13g2_nor2b_1 _1137_ (.A(_0577_),
    .B_N(net47),
    .Y(_0008_));
 sg13g2_buf_1 _1138_ (.A(net75),
    .X(_0578_));
 sg13g2_or2_1 _1139_ (.X(_0579_),
    .B(_0546_),
    .A(net76));
 sg13g2_buf_2 _1140_ (.A(_0579_),
    .X(_0580_));
 sg13g2_nand2_1 _1141_ (.Y(_0581_),
    .A(net69),
    .B(_0580_));
 sg13g2_nand3_1 _1142_ (.B(\bitserial_cipher.bit_counter[3] ),
    .C(\bitserial_cipher.bit_counter[2] ),
    .A(net76),
    .Y(_0582_));
 sg13g2_nor2_1 _1143_ (.A(_0569_),
    .B(_0582_),
    .Y(_0583_));
 sg13g2_xnor2_1 _1144_ (.Y(_0584_),
    .A(\bitserial_cipher.bit_counter[4] ),
    .B(_0583_));
 sg13g2_nor2_1 _1145_ (.A(_0581_),
    .B(_0584_),
    .Y(_0009_));
 sg13g2_nand2_1 _1146_ (.Y(_0585_),
    .A(\bitserial_cipher.bit_counter[4] ),
    .B(_0583_));
 sg13g2_xor2_1 _1147_ (.B(_0585_),
    .A(\bitserial_cipher.bit_counter[5] ),
    .X(_0586_));
 sg13g2_nor2_1 _1148_ (.A(_0581_),
    .B(_0586_),
    .Y(_0010_));
 sg13g2_mux2_1 _1149_ (.A0(\bitserial_cipher.datapath.fifo_ff56 ),
    .A1(\bitserial_cipher.datapath.fifo_ff57 ),
    .S(net48),
    .X(_0587_));
 sg13g2_and2_1 _1150_ (.A(net47),
    .B(_0587_),
    .X(_0011_));
 sg13g2_mux2_1 _1151_ (.A0(\bitserial_cipher.datapath.fifo_ff57 ),
    .A1(\bitserial_cipher.datapath.fifo_ff58 ),
    .S(net48),
    .X(_0588_));
 sg13g2_and2_1 _1152_ (.A(net47),
    .B(_0588_),
    .X(_0012_));
 sg13g2_mux2_1 _1153_ (.A0(\bitserial_cipher.datapath.fifo_ff58 ),
    .A1(\bitserial_cipher.datapath.fifo_ff59 ),
    .S(net48),
    .X(_0589_));
 sg13g2_and2_1 _1154_ (.A(net47),
    .B(_0589_),
    .X(_0013_));
 sg13g2_mux2_1 _1155_ (.A0(\bitserial_cipher.datapath.fifo_ff59 ),
    .A1(\bitserial_cipher.datapath.fifo_ff60 ),
    .S(net48),
    .X(_0590_));
 sg13g2_and2_1 _1156_ (.A(net47),
    .B(_0590_),
    .X(_0014_));
 sg13g2_buf_1 _1157_ (.A(net72),
    .X(_0591_));
 sg13g2_mux2_1 _1158_ (.A0(\bitserial_cipher.datapath.fifo_ff60 ),
    .A1(\bitserial_cipher.datapath.fifo_ff61 ),
    .S(net48),
    .X(_0592_));
 sg13g2_and2_1 _1159_ (.A(net45),
    .B(_0592_),
    .X(_0015_));
 sg13g2_buf_1 _1160_ (.A(net74),
    .X(_0593_));
 sg13g2_mux2_1 _1161_ (.A0(\bitserial_cipher.datapath.fifo_ff61 ),
    .A1(\bitserial_cipher.datapath.fifo_ff62 ),
    .S(_0593_),
    .X(_0594_));
 sg13g2_and2_1 _1162_ (.A(net45),
    .B(_0594_),
    .X(_0016_));
 sg13g2_mux2_1 _1163_ (.A0(\bitserial_cipher.datapath.fifo_ff62 ),
    .A1(\bitserial_cipher.datapath.fifo_ff63 ),
    .S(_0593_),
    .X(_0595_));
 sg13g2_and2_1 _1164_ (.A(net45),
    .B(_0595_),
    .X(_0017_));
 sg13g2_buf_2 _1165_ (.A(_0000_),
    .X(_0596_));
 sg13g2_xnor2_1 _1166_ (.Y(_0597_),
    .A(\bitserial_cipher.cipher_out ),
    .B(\bitserial_cipher.datapath.key_in ));
 sg13g2_buf_2 _1167_ (.A(\bitserial_cipher.datapath.round_counter[0] ),
    .X(_0598_));
 sg13g2_mux2_1 _1168_ (.A0(\bitserial_cipher.datapath.fifo_ff62 ),
    .A1(\bitserial_cipher.datapath.lut_ff62 ),
    .S(_0598_),
    .X(_0599_));
 sg13g2_xnor2_1 _1169_ (.Y(_0600_),
    .A(_0597_),
    .B(_0599_));
 sg13g2_buf_1 _1170_ (.A(_0598_),
    .X(_0601_));
 sg13g2_nand2_1 _1171_ (.Y(_0602_),
    .A(\bitserial_cipher.datapath.fifo_ff63 ),
    .B(\bitserial_cipher.datapath.fifo_ff56 ));
 sg13g2_nand3_1 _1172_ (.B(\bitserial_cipher.datapath.lut_ff63 ),
    .C(\bitserial_cipher.datapath.lut_ff56 ),
    .A(net43),
    .Y(_0603_));
 sg13g2_o21ai_1 _1173_ (.B1(_0603_),
    .Y(_0604_),
    .A1(net43),
    .A2(_0602_));
 sg13g2_xnor2_1 _1174_ (.Y(_0605_),
    .A(_0600_),
    .B(_0604_));
 sg13g2_nand2_1 _1175_ (.Y(_0606_),
    .A(_0596_),
    .B(\bitserial_cipher.datapath.shift_in2 ));
 sg13g2_o21ai_1 _1176_ (.B1(_0606_),
    .Y(_0607_),
    .A1(_0596_),
    .A2(_0605_));
 sg13g2_nor2b_1 _1177_ (.A(_0547_),
    .B_N(net2),
    .Y(_0608_));
 sg13g2_a21oi_1 _1178_ (.A1(net73),
    .A2(_0607_),
    .Y(_0609_),
    .B1(_0608_));
 sg13g2_nor2_1 _1179_ (.A(net48),
    .B(\bitserial_cipher.datapath.fifo_ff63 ),
    .Y(_0610_));
 sg13g2_a21oi_1 _1180_ (.A1(net48),
    .A2(_0609_),
    .Y(_0611_),
    .B1(_0610_));
 sg13g2_and2_1 _1181_ (.A(net45),
    .B(_0611_),
    .X(_0018_));
 sg13g2_and2_1 _1182_ (.A(net45),
    .B(\bitserial_cipher.datapath.lut_ff57 ),
    .X(_0019_));
 sg13g2_and2_1 _1183_ (.A(net45),
    .B(\bitserial_cipher.datapath.lut_ff58 ),
    .X(_0020_));
 sg13g2_and2_1 _1184_ (.A(net45),
    .B(\bitserial_cipher.datapath.lut_ff59 ),
    .X(_0021_));
 sg13g2_and2_1 _1185_ (.A(_0591_),
    .B(\bitserial_cipher.datapath.lut_ff60 ),
    .X(_0022_));
 sg13g2_and2_1 _1186_ (.A(_0591_),
    .B(\bitserial_cipher.datapath.lut_ff61 ),
    .X(_0023_));
 sg13g2_and2_1 _1187_ (.A(net45),
    .B(\bitserial_cipher.datapath.lut_ff62 ),
    .X(_0024_));
 sg13g2_buf_1 _1188_ (.A(net72),
    .X(_0612_));
 sg13g2_and2_1 _1189_ (.A(net42),
    .B(\bitserial_cipher.datapath.lut_ff63 ),
    .X(_0025_));
 sg13g2_nand2_1 _1190_ (.Y(_0613_),
    .A(net43),
    .B(\bitserial_cipher.datapath.shift_in2 ));
 sg13g2_o21ai_1 _1191_ (.B1(_0613_),
    .Y(_0614_),
    .A1(net43),
    .A2(_0605_));
 sg13g2_and2_1 _1192_ (.A(net42),
    .B(_0614_),
    .X(_0026_));
 sg13g2_mux2_1 _1193_ (.A0(\bitserial_cipher.datapath.shift_in2 ),
    .A1(\bitserial_cipher.datapath.shifter1[1] ),
    .S(net44),
    .X(_0615_));
 sg13g2_and2_1 _1194_ (.A(net42),
    .B(_0615_),
    .X(_0027_));
 sg13g2_mux2_1 _1195_ (.A0(\bitserial_cipher.datapath.shifter1[10] ),
    .A1(\bitserial_cipher.datapath.shifter1[11] ),
    .S(net44),
    .X(_0616_));
 sg13g2_and2_1 _1196_ (.A(net42),
    .B(_0616_),
    .X(_0028_));
 sg13g2_mux2_1 _1197_ (.A0(\bitserial_cipher.datapath.shifter1[11] ),
    .A1(\bitserial_cipher.datapath.shifter1[12] ),
    .S(net44),
    .X(_0617_));
 sg13g2_and2_1 _1198_ (.A(net42),
    .B(_0617_),
    .X(_0029_));
 sg13g2_mux2_1 _1199_ (.A0(\bitserial_cipher.datapath.shifter1[12] ),
    .A1(\bitserial_cipher.datapath.shifter1[13] ),
    .S(net44),
    .X(_0618_));
 sg13g2_and2_1 _1200_ (.A(net42),
    .B(_0618_),
    .X(_0030_));
 sg13g2_mux2_1 _1201_ (.A0(\bitserial_cipher.datapath.shifter1[13] ),
    .A1(\bitserial_cipher.datapath.shifter1[14] ),
    .S(net44),
    .X(_0619_));
 sg13g2_and2_1 _1202_ (.A(net42),
    .B(_0619_),
    .X(_0031_));
 sg13g2_mux2_1 _1203_ (.A0(\bitserial_cipher.datapath.shifter1[14] ),
    .A1(\bitserial_cipher.datapath.shifter1[15] ),
    .S(net44),
    .X(_0620_));
 sg13g2_and2_1 _1204_ (.A(net42),
    .B(_0620_),
    .X(_0032_));
 sg13g2_mux2_1 _1205_ (.A0(\bitserial_cipher.datapath.shifter1[15] ),
    .A1(\bitserial_cipher.datapath.shifter1[16] ),
    .S(net44),
    .X(_0621_));
 sg13g2_and2_1 _1206_ (.A(_0612_),
    .B(_0621_),
    .X(_0033_));
 sg13g2_mux2_1 _1207_ (.A0(\bitserial_cipher.datapath.shifter1[16] ),
    .A1(\bitserial_cipher.datapath.shifter1[17] ),
    .S(net44),
    .X(_0622_));
 sg13g2_and2_1 _1208_ (.A(_0612_),
    .B(_0622_),
    .X(_0034_));
 sg13g2_buf_1 _1209_ (.A(_0555_),
    .X(_0623_));
 sg13g2_buf_1 _1210_ (.A(net74),
    .X(_0624_));
 sg13g2_mux2_1 _1211_ (.A0(\bitserial_cipher.datapath.shifter1[17] ),
    .A1(\bitserial_cipher.datapath.shifter1[18] ),
    .S(net40),
    .X(_0625_));
 sg13g2_and2_1 _1212_ (.A(net41),
    .B(_0625_),
    .X(_0035_));
 sg13g2_mux2_1 _1213_ (.A0(\bitserial_cipher.datapath.shifter1[18] ),
    .A1(\bitserial_cipher.datapath.shifter1[19] ),
    .S(net40),
    .X(_0626_));
 sg13g2_and2_1 _1214_ (.A(net41),
    .B(_0626_),
    .X(_0036_));
 sg13g2_mux2_1 _1215_ (.A0(\bitserial_cipher.datapath.shifter1[19] ),
    .A1(\bitserial_cipher.datapath.shifter1[20] ),
    .S(net40),
    .X(_0627_));
 sg13g2_and2_1 _1216_ (.A(net41),
    .B(_0627_),
    .X(_0037_));
 sg13g2_mux2_1 _1217_ (.A0(\bitserial_cipher.datapath.shifter1[1] ),
    .A1(\bitserial_cipher.datapath.shifter1[2] ),
    .S(net40),
    .X(_0628_));
 sg13g2_and2_1 _1218_ (.A(net41),
    .B(_0628_),
    .X(_0038_));
 sg13g2_mux2_1 _1219_ (.A0(\bitserial_cipher.datapath.shifter1[20] ),
    .A1(\bitserial_cipher.datapath.shifter1[21] ),
    .S(_0624_),
    .X(_0629_));
 sg13g2_and2_1 _1220_ (.A(_0623_),
    .B(_0629_),
    .X(_0039_));
 sg13g2_mux2_1 _1221_ (.A0(\bitserial_cipher.datapath.shifter1[21] ),
    .A1(\bitserial_cipher.datapath.shifter1[22] ),
    .S(net40),
    .X(_0630_));
 sg13g2_and2_1 _1222_ (.A(net41),
    .B(_0630_),
    .X(_0040_));
 sg13g2_mux2_1 _1223_ (.A0(\bitserial_cipher.datapath.shifter1[22] ),
    .A1(\bitserial_cipher.datapath.shifter1[23] ),
    .S(net40),
    .X(_0631_));
 sg13g2_and2_1 _1224_ (.A(net41),
    .B(_0631_),
    .X(_0041_));
 sg13g2_mux2_1 _1225_ (.A0(\bitserial_cipher.datapath.shifter1[23] ),
    .A1(\bitserial_cipher.datapath.shifter1[24] ),
    .S(_0624_),
    .X(_0632_));
 sg13g2_and2_1 _1226_ (.A(_0623_),
    .B(_0632_),
    .X(_0042_));
 sg13g2_mux2_1 _1227_ (.A0(\bitserial_cipher.datapath.shifter1[24] ),
    .A1(\bitserial_cipher.datapath.shifter1[25] ),
    .S(net40),
    .X(_0633_));
 sg13g2_and2_1 _1228_ (.A(net41),
    .B(_0633_),
    .X(_0043_));
 sg13g2_mux2_1 _1229_ (.A0(\bitserial_cipher.datapath.shifter1[25] ),
    .A1(\bitserial_cipher.datapath.shifter1[26] ),
    .S(net40),
    .X(_0634_));
 sg13g2_and2_1 _1230_ (.A(net41),
    .B(_0634_),
    .X(_0044_));
 sg13g2_buf_1 _1231_ (.A(net72),
    .X(_0635_));
 sg13g2_buf_1 _1232_ (.A(net74),
    .X(_0636_));
 sg13g2_mux2_1 _1233_ (.A0(\bitserial_cipher.datapath.shifter1[26] ),
    .A1(\bitserial_cipher.datapath.shifter1[27] ),
    .S(_0636_),
    .X(_0637_));
 sg13g2_and2_1 _1234_ (.A(net39),
    .B(_0637_),
    .X(_0045_));
 sg13g2_mux2_1 _1235_ (.A0(\bitserial_cipher.datapath.shifter1[27] ),
    .A1(\bitserial_cipher.datapath.shifter1[28] ),
    .S(_0636_),
    .X(_0638_));
 sg13g2_and2_1 _1236_ (.A(_0635_),
    .B(_0638_),
    .X(_0046_));
 sg13g2_mux2_1 _1237_ (.A0(\bitserial_cipher.datapath.shifter1[28] ),
    .A1(\bitserial_cipher.datapath.shifter1[29] ),
    .S(net38),
    .X(_0639_));
 sg13g2_and2_1 _1238_ (.A(net39),
    .B(_0639_),
    .X(_0047_));
 sg13g2_mux2_1 _1239_ (.A0(\bitserial_cipher.datapath.shifter1[29] ),
    .A1(\bitserial_cipher.datapath.shifter1[30] ),
    .S(net38),
    .X(_0640_));
 sg13g2_and2_1 _1240_ (.A(net39),
    .B(_0640_),
    .X(_0048_));
 sg13g2_mux2_1 _1241_ (.A0(\bitserial_cipher.datapath.shifter1[2] ),
    .A1(\bitserial_cipher.datapath.shifter1[3] ),
    .S(net38),
    .X(_0641_));
 sg13g2_and2_1 _1242_ (.A(net39),
    .B(_0641_),
    .X(_0049_));
 sg13g2_mux2_1 _1243_ (.A0(\bitserial_cipher.datapath.shifter1[30] ),
    .A1(\bitserial_cipher.datapath.shifter1[31] ),
    .S(net38),
    .X(_0642_));
 sg13g2_and2_1 _1244_ (.A(_0635_),
    .B(_0642_),
    .X(_0050_));
 sg13g2_mux2_1 _1245_ (.A0(\bitserial_cipher.datapath.shifter1[31] ),
    .A1(\bitserial_cipher.datapath.shifter1[32] ),
    .S(net38),
    .X(_0643_));
 sg13g2_and2_1 _1246_ (.A(net39),
    .B(_0643_),
    .X(_0051_));
 sg13g2_mux2_1 _1247_ (.A0(\bitserial_cipher.datapath.shifter1[32] ),
    .A1(\bitserial_cipher.datapath.shifter1[33] ),
    .S(net38),
    .X(_0644_));
 sg13g2_and2_1 _1248_ (.A(net39),
    .B(_0644_),
    .X(_0052_));
 sg13g2_mux2_1 _1249_ (.A0(\bitserial_cipher.datapath.shifter1[33] ),
    .A1(\bitserial_cipher.datapath.shifter1[34] ),
    .S(net38),
    .X(_0645_));
 sg13g2_and2_1 _1250_ (.A(net39),
    .B(_0645_),
    .X(_0053_));
 sg13g2_mux2_1 _1251_ (.A0(\bitserial_cipher.datapath.shifter1[34] ),
    .A1(\bitserial_cipher.datapath.shifter1[35] ),
    .S(net38),
    .X(_0646_));
 sg13g2_and2_1 _1252_ (.A(net39),
    .B(_0646_),
    .X(_0054_));
 sg13g2_buf_1 _1253_ (.A(_0555_),
    .X(_0647_));
 sg13g2_buf_1 _1254_ (.A(net74),
    .X(_0648_));
 sg13g2_mux2_1 _1255_ (.A0(\bitserial_cipher.datapath.shifter1[35] ),
    .A1(\bitserial_cipher.datapath.shifter1[36] ),
    .S(net36),
    .X(_0649_));
 sg13g2_and2_1 _1256_ (.A(net37),
    .B(_0649_),
    .X(_0055_));
 sg13g2_mux2_1 _1257_ (.A0(\bitserial_cipher.datapath.shifter1[36] ),
    .A1(\bitserial_cipher.datapath.shifter1[37] ),
    .S(net36),
    .X(_0650_));
 sg13g2_and2_1 _1258_ (.A(_0647_),
    .B(_0650_),
    .X(_0056_));
 sg13g2_mux2_1 _1259_ (.A0(\bitserial_cipher.datapath.shifter1[37] ),
    .A1(\bitserial_cipher.datapath.shifter1[38] ),
    .S(_0648_),
    .X(_0651_));
 sg13g2_and2_1 _1260_ (.A(_0647_),
    .B(_0651_),
    .X(_0057_));
 sg13g2_mux2_1 _1261_ (.A0(\bitserial_cipher.datapath.shifter1[38] ),
    .A1(\bitserial_cipher.datapath.shifter1[39] ),
    .S(_0648_),
    .X(_0652_));
 sg13g2_and2_1 _1262_ (.A(net37),
    .B(_0652_),
    .X(_0058_));
 sg13g2_mux2_1 _1263_ (.A0(\bitserial_cipher.datapath.shifter1[39] ),
    .A1(\bitserial_cipher.datapath.shifter1[40] ),
    .S(net36),
    .X(_0653_));
 sg13g2_and2_1 _1264_ (.A(net37),
    .B(_0653_),
    .X(_0059_));
 sg13g2_mux2_1 _1265_ (.A0(\bitserial_cipher.datapath.shifter1[3] ),
    .A1(\bitserial_cipher.datapath.shifter1[4] ),
    .S(net36),
    .X(_0654_));
 sg13g2_and2_1 _1266_ (.A(net37),
    .B(_0654_),
    .X(_0060_));
 sg13g2_mux2_1 _1267_ (.A0(\bitserial_cipher.datapath.shifter1[40] ),
    .A1(\bitserial_cipher.datapath.shifter1[41] ),
    .S(net36),
    .X(_0655_));
 sg13g2_and2_1 _1268_ (.A(net37),
    .B(_0655_),
    .X(_0061_));
 sg13g2_mux2_1 _1269_ (.A0(\bitserial_cipher.datapath.shifter1[41] ),
    .A1(\bitserial_cipher.datapath.shifter1[42] ),
    .S(net36),
    .X(_0656_));
 sg13g2_and2_1 _1270_ (.A(net37),
    .B(_0656_),
    .X(_0062_));
 sg13g2_mux2_1 _1271_ (.A0(\bitserial_cipher.datapath.shifter1[42] ),
    .A1(\bitserial_cipher.datapath.shifter1[43] ),
    .S(net36),
    .X(_0657_));
 sg13g2_and2_1 _1272_ (.A(net37),
    .B(_0657_),
    .X(_0063_));
 sg13g2_mux2_1 _1273_ (.A0(\bitserial_cipher.datapath.shifter1[43] ),
    .A1(\bitserial_cipher.datapath.shifter1[44] ),
    .S(net36),
    .X(_0658_));
 sg13g2_and2_1 _1274_ (.A(net37),
    .B(_0658_),
    .X(_0064_));
 sg13g2_buf_1 _1275_ (.A(net72),
    .X(_0659_));
 sg13g2_buf_1 _1276_ (.A(net74),
    .X(_0660_));
 sg13g2_mux2_1 _1277_ (.A0(\bitserial_cipher.datapath.shifter1[44] ),
    .A1(\bitserial_cipher.datapath.shifter1[45] ),
    .S(net34),
    .X(_0661_));
 sg13g2_and2_1 _1278_ (.A(net35),
    .B(_0661_),
    .X(_0065_));
 sg13g2_mux2_1 _1279_ (.A0(\bitserial_cipher.datapath.shifter1[45] ),
    .A1(\bitserial_cipher.datapath.shifter1[46] ),
    .S(net34),
    .X(_0662_));
 sg13g2_and2_1 _1280_ (.A(net35),
    .B(_0662_),
    .X(_0066_));
 sg13g2_mux2_1 _1281_ (.A0(\bitserial_cipher.datapath.shifter1[46] ),
    .A1(\bitserial_cipher.datapath.shifter1[47] ),
    .S(net34),
    .X(_0663_));
 sg13g2_and2_1 _1282_ (.A(net35),
    .B(_0663_),
    .X(_0067_));
 sg13g2_mux2_1 _1283_ (.A0(\bitserial_cipher.datapath.shifter1[47] ),
    .A1(\bitserial_cipher.datapath.shifter1[48] ),
    .S(net34),
    .X(_0664_));
 sg13g2_and2_1 _1284_ (.A(net35),
    .B(_0664_),
    .X(_0068_));
 sg13g2_mux2_1 _1285_ (.A0(\bitserial_cipher.datapath.shifter1[48] ),
    .A1(\bitserial_cipher.datapath.shifter1[49] ),
    .S(net34),
    .X(_0665_));
 sg13g2_and2_1 _1286_ (.A(net35),
    .B(_0665_),
    .X(_0069_));
 sg13g2_mux2_1 _1287_ (.A0(\bitserial_cipher.datapath.shifter1[49] ),
    .A1(\bitserial_cipher.datapath.shifter1[50] ),
    .S(net34),
    .X(_0666_));
 sg13g2_and2_1 _1288_ (.A(net35),
    .B(_0666_),
    .X(_0070_));
 sg13g2_mux2_1 _1289_ (.A0(\bitserial_cipher.datapath.shifter1[4] ),
    .A1(\bitserial_cipher.datapath.shifter1[5] ),
    .S(net34),
    .X(_0667_));
 sg13g2_and2_1 _1290_ (.A(net35),
    .B(_0667_),
    .X(_0071_));
 sg13g2_mux2_1 _1291_ (.A0(\bitserial_cipher.datapath.shifter1[50] ),
    .A1(\bitserial_cipher.datapath.shifter1[51] ),
    .S(net34),
    .X(_0668_));
 sg13g2_and2_1 _1292_ (.A(net35),
    .B(_0668_),
    .X(_0072_));
 sg13g2_mux2_1 _1293_ (.A0(\bitserial_cipher.datapath.shifter1[51] ),
    .A1(\bitserial_cipher.datapath.shifter1[52] ),
    .S(_0660_),
    .X(_0669_));
 sg13g2_and2_1 _1294_ (.A(_0659_),
    .B(_0669_),
    .X(_0073_));
 sg13g2_mux2_1 _1295_ (.A0(\bitserial_cipher.datapath.shifter1[52] ),
    .A1(\bitserial_cipher.datapath.shifter1[53] ),
    .S(_0660_),
    .X(_0670_));
 sg13g2_and2_1 _1296_ (.A(_0659_),
    .B(_0670_),
    .X(_0074_));
 sg13g2_buf_1 _1297_ (.A(net72),
    .X(_0671_));
 sg13g2_buf_1 _1298_ (.A(net74),
    .X(_0672_));
 sg13g2_mux2_1 _1299_ (.A0(\bitserial_cipher.datapath.shifter1[53] ),
    .A1(\bitserial_cipher.datapath.shifter1[54] ),
    .S(_0672_),
    .X(_0673_));
 sg13g2_and2_1 _1300_ (.A(_0671_),
    .B(_0673_),
    .X(_0075_));
 sg13g2_mux2_1 _1301_ (.A0(\bitserial_cipher.datapath.shifter1[54] ),
    .A1(\bitserial_cipher.datapath.shifter1[55] ),
    .S(net32),
    .X(_0674_));
 sg13g2_and2_1 _1302_ (.A(net33),
    .B(_0674_),
    .X(_0076_));
 sg13g2_inv_1 _1303_ (.Y(_0675_),
    .A(_0546_));
 sg13g2_inv_1 _1304_ (.Y(_0676_),
    .A(_0598_));
 sg13g2_nor3_1 _1305_ (.A(\bitserial_cipher.bit_counter[3] ),
    .B(\bitserial_cipher.bit_counter[4] ),
    .C(\bitserial_cipher.bit_counter[5] ),
    .Y(_0677_));
 sg13g2_xnor2_1 _1306_ (.Y(_0678_),
    .A(_0676_),
    .B(_0677_));
 sg13g2_nor2_1 _1307_ (.A(_0675_),
    .B(_0678_),
    .Y(_0679_));
 sg13g2_mux2_1 _1308_ (.A0(\bitserial_cipher.datapath.fifo_ff56 ),
    .A1(\bitserial_cipher.datapath.lut_ff56 ),
    .S(_0679_),
    .X(_0680_));
 sg13g2_mux2_1 _1309_ (.A0(\bitserial_cipher.datapath.shifter1[55] ),
    .A1(_0680_),
    .S(net32),
    .X(_0681_));
 sg13g2_and2_1 _1310_ (.A(net33),
    .B(_0681_),
    .X(_0077_));
 sg13g2_mux2_1 _1311_ (.A0(\bitserial_cipher.datapath.shifter1[5] ),
    .A1(\bitserial_cipher.datapath.shifter1[6] ),
    .S(net32),
    .X(_0682_));
 sg13g2_and2_1 _1312_ (.A(net33),
    .B(_0682_),
    .X(_0078_));
 sg13g2_mux2_1 _1313_ (.A0(\bitserial_cipher.datapath.shifter1[6] ),
    .A1(\bitserial_cipher.datapath.shifter1[7] ),
    .S(net32),
    .X(_0683_));
 sg13g2_and2_1 _1314_ (.A(net33),
    .B(_0683_),
    .X(_0079_));
 sg13g2_mux2_1 _1315_ (.A0(\bitserial_cipher.datapath.shifter1[7] ),
    .A1(\bitserial_cipher.datapath.shifter1[8] ),
    .S(net32),
    .X(_0684_));
 sg13g2_and2_1 _1316_ (.A(net33),
    .B(_0684_),
    .X(_0080_));
 sg13g2_mux2_1 _1317_ (.A0(\bitserial_cipher.datapath.shifter1[8] ),
    .A1(\bitserial_cipher.datapath.shifter1[9] ),
    .S(net32),
    .X(_0685_));
 sg13g2_and2_1 _1318_ (.A(net33),
    .B(_0685_),
    .X(_0081_));
 sg13g2_mux2_1 _1319_ (.A0(\bitserial_cipher.datapath.shifter1[9] ),
    .A1(\bitserial_cipher.datapath.shifter1[10] ),
    .S(net32),
    .X(_0686_));
 sg13g2_and2_1 _1320_ (.A(net33),
    .B(_0686_),
    .X(_0082_));
 sg13g2_mux2_1 _1321_ (.A0(\bitserial_cipher.cipher_out ),
    .A1(\bitserial_cipher.datapath.shifter2[1] ),
    .S(_0672_),
    .X(_0687_));
 sg13g2_and2_1 _1322_ (.A(_0671_),
    .B(_0687_),
    .X(_0083_));
 sg13g2_mux2_1 _1323_ (.A0(\bitserial_cipher.datapath.shifter2[10] ),
    .A1(\bitserial_cipher.datapath.shifter2[11] ),
    .S(net32),
    .X(_0688_));
 sg13g2_and2_1 _1324_ (.A(net33),
    .B(_0688_),
    .X(_0084_));
 sg13g2_buf_1 _1325_ (.A(net72),
    .X(_0689_));
 sg13g2_buf_1 _1326_ (.A(net74),
    .X(_0690_));
 sg13g2_mux2_1 _1327_ (.A0(\bitserial_cipher.datapath.shifter2[11] ),
    .A1(\bitserial_cipher.datapath.shifter2[12] ),
    .S(net30),
    .X(_0691_));
 sg13g2_and2_1 _1328_ (.A(_0689_),
    .B(_0691_),
    .X(_0085_));
 sg13g2_mux2_1 _1329_ (.A0(\bitserial_cipher.datapath.shifter2[12] ),
    .A1(\bitserial_cipher.datapath.shifter2[13] ),
    .S(net30),
    .X(_0692_));
 sg13g2_and2_1 _1330_ (.A(_0689_),
    .B(_0692_),
    .X(_0086_));
 sg13g2_mux2_1 _1331_ (.A0(\bitserial_cipher.datapath.shifter2[13] ),
    .A1(\bitserial_cipher.datapath.shifter2[14] ),
    .S(_0690_),
    .X(_0693_));
 sg13g2_and2_1 _1332_ (.A(net31),
    .B(_0693_),
    .X(_0087_));
 sg13g2_mux2_1 _1333_ (.A0(\bitserial_cipher.datapath.shifter2[14] ),
    .A1(\bitserial_cipher.datapath.shifter2[15] ),
    .S(_0690_),
    .X(_0694_));
 sg13g2_and2_1 _1334_ (.A(net31),
    .B(_0694_),
    .X(_0088_));
 sg13g2_mux2_1 _1335_ (.A0(\bitserial_cipher.datapath.shifter2[15] ),
    .A1(\bitserial_cipher.datapath.shifter2[16] ),
    .S(net30),
    .X(_0695_));
 sg13g2_and2_1 _1336_ (.A(net31),
    .B(_0695_),
    .X(_0089_));
 sg13g2_mux2_1 _1337_ (.A0(\bitserial_cipher.datapath.shifter2[16] ),
    .A1(\bitserial_cipher.datapath.shifter2[17] ),
    .S(net30),
    .X(_0696_));
 sg13g2_and2_1 _1338_ (.A(net31),
    .B(_0696_),
    .X(_0090_));
 sg13g2_mux2_1 _1339_ (.A0(\bitserial_cipher.datapath.shifter2[17] ),
    .A1(\bitserial_cipher.datapath.shifter2[18] ),
    .S(net30),
    .X(_0697_));
 sg13g2_and2_1 _1340_ (.A(net31),
    .B(_0697_),
    .X(_0091_));
 sg13g2_mux2_1 _1341_ (.A0(\bitserial_cipher.datapath.shifter2[18] ),
    .A1(\bitserial_cipher.datapath.shifter2[19] ),
    .S(net30),
    .X(_0698_));
 sg13g2_and2_1 _1342_ (.A(net31),
    .B(_0698_),
    .X(_0092_));
 sg13g2_mux2_1 _1343_ (.A0(\bitserial_cipher.datapath.shifter2[19] ),
    .A1(\bitserial_cipher.datapath.shifter2[20] ),
    .S(net30),
    .X(_0699_));
 sg13g2_and2_1 _1344_ (.A(net31),
    .B(_0699_),
    .X(_0093_));
 sg13g2_mux2_1 _1345_ (.A0(\bitserial_cipher.datapath.shifter2[1] ),
    .A1(\bitserial_cipher.datapath.shifter2[2] ),
    .S(net30),
    .X(_0700_));
 sg13g2_and2_1 _1346_ (.A(net31),
    .B(_0700_),
    .X(_0094_));
 sg13g2_buf_1 _1347_ (.A(net72),
    .X(_0701_));
 sg13g2_buf_1 _1348_ (.A(net74),
    .X(_0702_));
 sg13g2_mux2_1 _1349_ (.A0(\bitserial_cipher.datapath.shifter2[20] ),
    .A1(\bitserial_cipher.datapath.shifter2[21] ),
    .S(net28),
    .X(_0703_));
 sg13g2_and2_1 _1350_ (.A(net29),
    .B(_0703_),
    .X(_0095_));
 sg13g2_mux2_1 _1351_ (.A0(\bitserial_cipher.datapath.shifter2[21] ),
    .A1(\bitserial_cipher.datapath.shifter2[22] ),
    .S(net28),
    .X(_0704_));
 sg13g2_and2_1 _1352_ (.A(net29),
    .B(_0704_),
    .X(_0096_));
 sg13g2_mux2_1 _1353_ (.A0(\bitserial_cipher.datapath.shifter2[22] ),
    .A1(\bitserial_cipher.datapath.shifter2[23] ),
    .S(net28),
    .X(_0705_));
 sg13g2_and2_1 _1354_ (.A(net29),
    .B(_0705_),
    .X(_0097_));
 sg13g2_mux2_1 _1355_ (.A0(\bitserial_cipher.datapath.shifter2[23] ),
    .A1(\bitserial_cipher.datapath.shifter2[24] ),
    .S(net28),
    .X(_0706_));
 sg13g2_and2_1 _1356_ (.A(net29),
    .B(_0706_),
    .X(_0098_));
 sg13g2_mux2_1 _1357_ (.A0(\bitserial_cipher.datapath.shifter2[24] ),
    .A1(\bitserial_cipher.datapath.shifter2[25] ),
    .S(_0702_),
    .X(_0707_));
 sg13g2_and2_1 _1358_ (.A(_0701_),
    .B(_0707_),
    .X(_0099_));
 sg13g2_mux2_1 _1359_ (.A0(\bitserial_cipher.datapath.shifter2[25] ),
    .A1(\bitserial_cipher.datapath.shifter2[26] ),
    .S(net28),
    .X(_0708_));
 sg13g2_and2_1 _1360_ (.A(net29),
    .B(_0708_),
    .X(_0100_));
 sg13g2_mux2_1 _1361_ (.A0(\bitserial_cipher.datapath.shifter2[26] ),
    .A1(\bitserial_cipher.datapath.shifter2[27] ),
    .S(_0702_),
    .X(_0709_));
 sg13g2_and2_1 _1362_ (.A(_0701_),
    .B(_0709_),
    .X(_0101_));
 sg13g2_mux2_1 _1363_ (.A0(\bitserial_cipher.datapath.shifter2[27] ),
    .A1(\bitserial_cipher.datapath.shifter2[28] ),
    .S(net28),
    .X(_0710_));
 sg13g2_and2_1 _1364_ (.A(net29),
    .B(_0710_),
    .X(_0102_));
 sg13g2_mux2_1 _1365_ (.A0(\bitserial_cipher.datapath.shifter2[28] ),
    .A1(\bitserial_cipher.datapath.shifter2[29] ),
    .S(net28),
    .X(_0711_));
 sg13g2_and2_1 _1366_ (.A(net29),
    .B(_0711_),
    .X(_0103_));
 sg13g2_mux2_1 _1367_ (.A0(\bitserial_cipher.datapath.shifter2[29] ),
    .A1(\bitserial_cipher.datapath.shifter2[30] ),
    .S(net28),
    .X(_0712_));
 sg13g2_and2_1 _1368_ (.A(net29),
    .B(_0712_),
    .X(_0104_));
 sg13g2_buf_1 _1369_ (.A(net75),
    .X(_0713_));
 sg13g2_buf_1 _1370_ (.A(net68),
    .X(_0714_));
 sg13g2_buf_1 _1371_ (.A(net76),
    .X(_0715_));
 sg13g2_mux2_1 _1372_ (.A0(\bitserial_cipher.datapath.shifter2[2] ),
    .A1(\bitserial_cipher.datapath.shifter2[3] ),
    .S(net67),
    .X(_0716_));
 sg13g2_and2_1 _1373_ (.A(net27),
    .B(_0716_),
    .X(_0105_));
 sg13g2_mux2_1 _1374_ (.A0(\bitserial_cipher.datapath.shifter2[30] ),
    .A1(\bitserial_cipher.datapath.shifter2[31] ),
    .S(net67),
    .X(_0717_));
 sg13g2_and2_1 _1375_ (.A(net27),
    .B(_0717_),
    .X(_0106_));
 sg13g2_mux2_1 _1376_ (.A0(\bitserial_cipher.datapath.shifter2[31] ),
    .A1(\bitserial_cipher.datapath.shifter2[32] ),
    .S(net67),
    .X(_0718_));
 sg13g2_and2_1 _1377_ (.A(net27),
    .B(_0718_),
    .X(_0107_));
 sg13g2_mux2_1 _1378_ (.A0(\bitserial_cipher.datapath.shifter2[32] ),
    .A1(\bitserial_cipher.datapath.shifter2[33] ),
    .S(net67),
    .X(_0719_));
 sg13g2_and2_1 _1379_ (.A(net27),
    .B(_0719_),
    .X(_0108_));
 sg13g2_mux2_1 _1380_ (.A0(\bitserial_cipher.datapath.shifter2[33] ),
    .A1(\bitserial_cipher.datapath.shifter2[34] ),
    .S(net67),
    .X(_0720_));
 sg13g2_and2_1 _1381_ (.A(net27),
    .B(_0720_),
    .X(_0109_));
 sg13g2_mux2_1 _1382_ (.A0(\bitserial_cipher.datapath.shifter2[34] ),
    .A1(\bitserial_cipher.datapath.shifter2[35] ),
    .S(net67),
    .X(_0721_));
 sg13g2_and2_1 _1383_ (.A(net27),
    .B(_0721_),
    .X(_0110_));
 sg13g2_mux2_1 _1384_ (.A0(\bitserial_cipher.datapath.shifter2[35] ),
    .A1(\bitserial_cipher.datapath.shifter2[36] ),
    .S(net67),
    .X(_0722_));
 sg13g2_and2_1 _1385_ (.A(net27),
    .B(_0722_),
    .X(_0111_));
 sg13g2_mux2_1 _1386_ (.A0(\bitserial_cipher.datapath.shifter2[36] ),
    .A1(\bitserial_cipher.datapath.shifter2[37] ),
    .S(net67),
    .X(_0723_));
 sg13g2_and2_1 _1387_ (.A(net27),
    .B(_0723_),
    .X(_0112_));
 sg13g2_mux2_1 _1388_ (.A0(\bitserial_cipher.datapath.shifter2[37] ),
    .A1(\bitserial_cipher.datapath.shifter2[38] ),
    .S(_0715_),
    .X(_0724_));
 sg13g2_and2_1 _1389_ (.A(_0714_),
    .B(_0724_),
    .X(_0113_));
 sg13g2_mux2_1 _1390_ (.A0(\bitserial_cipher.datapath.shifter2[38] ),
    .A1(\bitserial_cipher.datapath.shifter2[39] ),
    .S(_0715_),
    .X(_0725_));
 sg13g2_and2_1 _1391_ (.A(_0714_),
    .B(_0725_),
    .X(_0114_));
 sg13g2_buf_1 _1392_ (.A(net68),
    .X(_0726_));
 sg13g2_buf_1 _1393_ (.A(net76),
    .X(_0727_));
 sg13g2_mux2_1 _1394_ (.A0(\bitserial_cipher.datapath.shifter2[39] ),
    .A1(\bitserial_cipher.datapath.shifter2[40] ),
    .S(_0727_),
    .X(_0728_));
 sg13g2_and2_1 _1395_ (.A(net26),
    .B(_0728_),
    .X(_0115_));
 sg13g2_mux2_1 _1396_ (.A0(\bitserial_cipher.datapath.shifter2[3] ),
    .A1(\bitserial_cipher.datapath.shifter2[4] ),
    .S(_0727_),
    .X(_0729_));
 sg13g2_and2_1 _1397_ (.A(_0726_),
    .B(_0729_),
    .X(_0116_));
 sg13g2_mux2_1 _1398_ (.A0(\bitserial_cipher.datapath.shifter2[40] ),
    .A1(\bitserial_cipher.datapath.shifter2[41] ),
    .S(net66),
    .X(_0730_));
 sg13g2_and2_1 _1399_ (.A(net26),
    .B(_0730_),
    .X(_0117_));
 sg13g2_mux2_1 _1400_ (.A0(\bitserial_cipher.datapath.shifter2[41] ),
    .A1(\bitserial_cipher.datapath.shifter2[42] ),
    .S(net66),
    .X(_0731_));
 sg13g2_and2_1 _1401_ (.A(_0726_),
    .B(_0731_),
    .X(_0118_));
 sg13g2_mux2_1 _1402_ (.A0(\bitserial_cipher.datapath.shifter2[42] ),
    .A1(\bitserial_cipher.datapath.shifter2[43] ),
    .S(net66),
    .X(_0732_));
 sg13g2_and2_1 _1403_ (.A(net26),
    .B(_0732_),
    .X(_0119_));
 sg13g2_mux2_1 _1404_ (.A0(\bitserial_cipher.datapath.shifter2[43] ),
    .A1(\bitserial_cipher.datapath.shifter2[44] ),
    .S(net66),
    .X(_0733_));
 sg13g2_and2_1 _1405_ (.A(net26),
    .B(_0733_),
    .X(_0120_));
 sg13g2_mux2_1 _1406_ (.A0(\bitserial_cipher.datapath.shifter2[44] ),
    .A1(\bitserial_cipher.datapath.shifter2[45] ),
    .S(net66),
    .X(_0734_));
 sg13g2_and2_1 _1407_ (.A(net26),
    .B(_0734_),
    .X(_0121_));
 sg13g2_mux2_1 _1408_ (.A0(\bitserial_cipher.datapath.shifter2[45] ),
    .A1(\bitserial_cipher.datapath.shifter2[46] ),
    .S(net66),
    .X(_0735_));
 sg13g2_and2_1 _1409_ (.A(net26),
    .B(_0735_),
    .X(_0122_));
 sg13g2_mux2_1 _1410_ (.A0(\bitserial_cipher.datapath.shifter2[46] ),
    .A1(\bitserial_cipher.datapath.shifter2[47] ),
    .S(net66),
    .X(_0736_));
 sg13g2_and2_1 _1411_ (.A(net26),
    .B(_0736_),
    .X(_0123_));
 sg13g2_mux2_1 _1412_ (.A0(\bitserial_cipher.datapath.shifter2[47] ),
    .A1(\bitserial_cipher.datapath.shifter2[48] ),
    .S(net66),
    .X(_0737_));
 sg13g2_and2_1 _1413_ (.A(net26),
    .B(_0737_),
    .X(_0124_));
 sg13g2_buf_1 _1414_ (.A(net68),
    .X(_0738_));
 sg13g2_buf_1 _1415_ (.A(net76),
    .X(_0739_));
 sg13g2_mux2_1 _1416_ (.A0(\bitserial_cipher.datapath.shifter2[48] ),
    .A1(\bitserial_cipher.datapath.shifter2[49] ),
    .S(net65),
    .X(_0740_));
 sg13g2_and2_1 _1417_ (.A(net25),
    .B(_0740_),
    .X(_0125_));
 sg13g2_mux2_1 _1418_ (.A0(\bitserial_cipher.datapath.shifter2[49] ),
    .A1(\bitserial_cipher.datapath.shifter2[50] ),
    .S(net65),
    .X(_0741_));
 sg13g2_and2_1 _1419_ (.A(net25),
    .B(_0741_),
    .X(_0126_));
 sg13g2_mux2_1 _1420_ (.A0(\bitserial_cipher.datapath.shifter2[4] ),
    .A1(\bitserial_cipher.datapath.shifter2[5] ),
    .S(net65),
    .X(_0742_));
 sg13g2_and2_1 _1421_ (.A(net25),
    .B(_0742_),
    .X(_0127_));
 sg13g2_mux2_1 _1422_ (.A0(\bitserial_cipher.datapath.shifter2[50] ),
    .A1(\bitserial_cipher.datapath.shifter2[51] ),
    .S(net65),
    .X(_0743_));
 sg13g2_and2_1 _1423_ (.A(net25),
    .B(_0743_),
    .X(_0128_));
 sg13g2_mux2_1 _1424_ (.A0(\bitserial_cipher.datapath.shifter2[51] ),
    .A1(\bitserial_cipher.datapath.shifter2[52] ),
    .S(net65),
    .X(_0744_));
 sg13g2_and2_1 _1425_ (.A(net25),
    .B(_0744_),
    .X(_0129_));
 sg13g2_mux2_1 _1426_ (.A0(\bitserial_cipher.datapath.shifter2[52] ),
    .A1(\bitserial_cipher.datapath.shifter2[53] ),
    .S(net65),
    .X(_0745_));
 sg13g2_and2_1 _1427_ (.A(net25),
    .B(_0745_),
    .X(_0130_));
 sg13g2_mux2_1 _1428_ (.A0(\bitserial_cipher.datapath.shifter2[53] ),
    .A1(\bitserial_cipher.datapath.shifter2[54] ),
    .S(net65),
    .X(_0746_));
 sg13g2_and2_1 _1429_ (.A(net25),
    .B(_0746_),
    .X(_0131_));
 sg13g2_mux2_1 _1430_ (.A0(\bitserial_cipher.datapath.shifter2[54] ),
    .A1(\bitserial_cipher.datapath.shifter2[55] ),
    .S(net65),
    .X(_0747_));
 sg13g2_and2_1 _1431_ (.A(net25),
    .B(_0747_),
    .X(_0132_));
 sg13g2_mux2_1 _1432_ (.A0(\bitserial_cipher.datapath.shifter2[55] ),
    .A1(\bitserial_cipher.datapath.shifter2[56] ),
    .S(_0739_),
    .X(_0748_));
 sg13g2_and2_1 _1433_ (.A(_0738_),
    .B(_0748_),
    .X(_0133_));
 sg13g2_mux2_1 _1434_ (.A0(\bitserial_cipher.datapath.shifter2[56] ),
    .A1(\bitserial_cipher.datapath.shifter2[57] ),
    .S(_0739_),
    .X(_0749_));
 sg13g2_and2_1 _1435_ (.A(_0738_),
    .B(_0749_),
    .X(_0134_));
 sg13g2_buf_1 _1436_ (.A(net68),
    .X(_0750_));
 sg13g2_buf_1 _1437_ (.A(net76),
    .X(_0751_));
 sg13g2_mux2_1 _1438_ (.A0(\bitserial_cipher.datapath.shifter2[57] ),
    .A1(\bitserial_cipher.datapath.shifter2[58] ),
    .S(net64),
    .X(_0752_));
 sg13g2_and2_1 _1439_ (.A(net24),
    .B(_0752_),
    .X(_0135_));
 sg13g2_mux2_1 _1440_ (.A0(\bitserial_cipher.datapath.shifter2[58] ),
    .A1(\bitserial_cipher.datapath.shifter2[59] ),
    .S(net64),
    .X(_0753_));
 sg13g2_and2_1 _1441_ (.A(net24),
    .B(_0753_),
    .X(_0136_));
 sg13g2_mux2_1 _1442_ (.A0(\bitserial_cipher.datapath.shifter2[59] ),
    .A1(\bitserial_cipher.datapath.shifter2[60] ),
    .S(net64),
    .X(_0754_));
 sg13g2_and2_1 _1443_ (.A(net24),
    .B(_0754_),
    .X(_0137_));
 sg13g2_mux2_1 _1444_ (.A0(\bitserial_cipher.datapath.shifter2[5] ),
    .A1(\bitserial_cipher.datapath.shifter2[6] ),
    .S(net64),
    .X(_0755_));
 sg13g2_and2_1 _1445_ (.A(net24),
    .B(_0755_),
    .X(_0138_));
 sg13g2_mux2_1 _1446_ (.A0(\bitserial_cipher.datapath.shifter2[60] ),
    .A1(\bitserial_cipher.datapath.shifter2[61] ),
    .S(net64),
    .X(_0756_));
 sg13g2_and2_1 _1447_ (.A(net24),
    .B(_0756_),
    .X(_0139_));
 sg13g2_mux2_1 _1448_ (.A0(\bitserial_cipher.datapath.shifter2[61] ),
    .A1(\bitserial_cipher.datapath.shifter2[62] ),
    .S(net64),
    .X(_0757_));
 sg13g2_and2_1 _1449_ (.A(_0750_),
    .B(_0757_),
    .X(_0140_));
 sg13g2_mux2_1 _1450_ (.A0(\bitserial_cipher.datapath.shifter2[62] ),
    .A1(\bitserial_cipher.datapath.shifter2[63] ),
    .S(_0751_),
    .X(_0758_));
 sg13g2_and2_1 _1451_ (.A(net24),
    .B(_0758_),
    .X(_0141_));
 sg13g2_mux2_1 _1452_ (.A0(\bitserial_cipher.datapath.shifter2[63] ),
    .A1(\bitserial_cipher.datapath.shift_in2 ),
    .S(_0751_),
    .X(_0759_));
 sg13g2_and2_1 _1453_ (.A(_0750_),
    .B(_0759_),
    .X(_0142_));
 sg13g2_mux2_1 _1454_ (.A0(\bitserial_cipher.datapath.shifter2[6] ),
    .A1(\bitserial_cipher.datapath.shifter2[7] ),
    .S(net64),
    .X(_0760_));
 sg13g2_and2_1 _1455_ (.A(net24),
    .B(_0760_),
    .X(_0143_));
 sg13g2_mux2_1 _1456_ (.A0(\bitserial_cipher.datapath.shifter2[7] ),
    .A1(\bitserial_cipher.datapath.shifter2[8] ),
    .S(net64),
    .X(_0761_));
 sg13g2_and2_1 _1457_ (.A(net24),
    .B(_0761_),
    .X(_0144_));
 sg13g2_buf_1 _1458_ (.A(net68),
    .X(_0762_));
 sg13g2_mux2_1 _1459_ (.A0(\bitserial_cipher.datapath.shifter2[8] ),
    .A1(\bitserial_cipher.datapath.shifter2[9] ),
    .S(net70),
    .X(_0763_));
 sg13g2_and2_1 _1460_ (.A(net23),
    .B(_0763_),
    .X(_0145_));
 sg13g2_mux2_1 _1461_ (.A0(\bitserial_cipher.datapath.shifter2[9] ),
    .A1(\bitserial_cipher.datapath.shifter2[10] ),
    .S(net70),
    .X(_0764_));
 sg13g2_and2_1 _1462_ (.A(net23),
    .B(_0764_),
    .X(_0146_));
 sg13g2_mux2_1 _1463_ (.A0(\bitserial_cipher.key_exp.fifo_ff0 ),
    .A1(\bitserial_cipher.key_exp.fifo_ff1 ),
    .S(net46),
    .X(_0765_));
 sg13g2_and2_1 _1464_ (.A(net23),
    .B(_0765_),
    .X(_0147_));
 sg13g2_mux2_1 _1465_ (.A0(\bitserial_cipher.key_exp.fifo_ff1 ),
    .A1(\bitserial_cipher.key_exp.fifo_ff2 ),
    .S(net46),
    .X(_0766_));
 sg13g2_and2_1 _1466_ (.A(net23),
    .B(_0766_),
    .X(_0148_));
 sg13g2_mux2_1 _1467_ (.A0(\bitserial_cipher.key_exp.fifo_ff2 ),
    .A1(\bitserial_cipher.key_exp.fifo_ff3 ),
    .S(_0558_),
    .X(_0767_));
 sg13g2_and2_1 _1468_ (.A(net23),
    .B(_0767_),
    .X(_0149_));
 sg13g2_inv_1 _1469_ (.Y(_0768_),
    .A(\bitserial_cipher.key_exp.fifo_ff3 ));
 sg13g2_nand2_1 _1470_ (.Y(_0769_),
    .A(net46),
    .B(\bitserial_cipher.key_exp.shift_out1 ));
 sg13g2_o21ai_1 _1471_ (.B1(_0769_),
    .Y(_0770_),
    .A1(_0558_),
    .A2(_0768_));
 sg13g2_and2_1 _1472_ (.A(net23),
    .B(_0770_),
    .X(_0150_));
 sg13g2_nor4_2 _1473_ (.A(\bitserial_cipher.bit_counter[3] ),
    .B(\bitserial_cipher.bit_counter[2] ),
    .C(\bitserial_cipher.bit_counter[4] ),
    .Y(_0771_),
    .D(\bitserial_cipher.bit_counter[5] ));
 sg13g2_and2_1 _1474_ (.A(net76),
    .B(_0771_),
    .X(_0772_));
 sg13g2_buf_1 _1475_ (.A(_0772_),
    .X(_0773_));
 sg13g2_nand2_2 _1476_ (.Y(_0774_),
    .A(net73),
    .B(_0773_));
 sg13g2_mux2_1 _1477_ (.A0(\bitserial_cipher.key_exp.lut_ff1 ),
    .A1(\bitserial_cipher.key_exp.lut_ff0 ),
    .S(_0774_),
    .X(_0775_));
 sg13g2_and2_1 _1478_ (.A(net23),
    .B(_0775_),
    .X(_0151_));
 sg13g2_mux2_1 _1479_ (.A0(\bitserial_cipher.key_exp.lut_ff2 ),
    .A1(\bitserial_cipher.key_exp.lut_ff1 ),
    .S(_0774_),
    .X(_0776_));
 sg13g2_and2_1 _1480_ (.A(_0762_),
    .B(_0776_),
    .X(_0152_));
 sg13g2_mux2_1 _1481_ (.A0(\bitserial_cipher.key_exp.lut_ff3 ),
    .A1(\bitserial_cipher.key_exp.lut_ff2 ),
    .S(_0774_),
    .X(_0777_));
 sg13g2_and2_1 _1482_ (.A(_0762_),
    .B(_0777_),
    .X(_0153_));
 sg13g2_buf_1 _1483_ (.A(\bitserial_cipher.datapath.round_counter[3] ),
    .X(_0778_));
 sg13g2_buf_1 _1484_ (.A(\bitserial_cipher.datapath.round_counter[2] ),
    .X(_0779_));
 sg13g2_nor2_1 _1485_ (.A(_0778_),
    .B(net62),
    .Y(_0780_));
 sg13g2_buf_8 _1486_ (.A(\bitserial_cipher.datapath.round_counter[4] ),
    .X(_0781_));
 sg13g2_nor2b_1 _1487_ (.A(_0780_),
    .B_N(net61),
    .Y(_0782_));
 sg13g2_buf_8 _1488_ (.A(net63),
    .X(_0783_));
 sg13g2_buf_8 _1489_ (.A(net62),
    .X(_0784_));
 sg13g2_inv_1 _1490_ (.Y(_0785_),
    .A(\bitserial_cipher.datapath.round_counter[6] ));
 sg13g2_buf_1 _1491_ (.A(\bitserial_cipher.datapath.round_counter[1] ),
    .X(_0786_));
 sg13g2_nor2_1 _1492_ (.A(_0786_),
    .B(_0598_),
    .Y(_0787_));
 sg13g2_nand4_1 _1493_ (.B(net21),
    .C(_0785_),
    .A(net22),
    .Y(_0788_),
    .D(_0787_));
 sg13g2_buf_1 _1494_ (.A(\bitserial_cipher.datapath.round_counter[5] ),
    .X(_0789_));
 sg13g2_nor2_1 _1495_ (.A(_0778_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_buf_8 _1496_ (.A(_0001_),
    .X(_0791_));
 sg13g2_nor2b_1 _1497_ (.A(_0598_),
    .B_N(_0791_),
    .Y(_0792_));
 sg13g2_or3_1 _1498_ (.A(net63),
    .B(net62),
    .C(net61),
    .X(_0793_));
 sg13g2_a221oi_1 _1499_ (.B2(_0792_),
    .C1(_0793_),
    .B1(_0790_),
    .A1(_0676_),
    .Y(_0794_),
    .A2(_0785_));
 sg13g2_a21o_1 _1500_ (.A2(_0788_),
    .A1(_0782_),
    .B1(_0794_),
    .X(_0795_));
 sg13g2_nor2b_1 _1501_ (.A(net62),
    .B_N(net63),
    .Y(_0796_));
 sg13g2_nor2b_2 _1502_ (.A(_0596_),
    .B_N(\bitserial_cipher.datapath.round_counter[1] ),
    .Y(_0797_));
 sg13g2_nor2b_1 _1503_ (.A(_0598_),
    .B_N(net63),
    .Y(_0798_));
 sg13g2_nor2_1 _1504_ (.A(net60),
    .B(net21),
    .Y(_0799_));
 sg13g2_a22oi_1 _1505_ (.Y(_0800_),
    .B1(_0798_),
    .B2(_0799_),
    .A2(_0797_),
    .A1(_0796_));
 sg13g2_nand2b_1 _1506_ (.Y(_0801_),
    .B(net62),
    .A_N(_0596_));
 sg13g2_or3_1 _1507_ (.A(net60),
    .B(net63),
    .C(_0801_),
    .X(_0802_));
 sg13g2_nor2b_1 _1508_ (.A(_0789_),
    .B_N(_0791_),
    .Y(_0803_));
 sg13g2_nor2_2 _1509_ (.A(net63),
    .B(\bitserial_cipher.datapath.round_counter[4] ),
    .Y(_0804_));
 sg13g2_a21oi_2 _1510_ (.B1(_0785_),
    .Y(_0805_),
    .A2(_0804_),
    .A1(_0803_));
 sg13g2_a21o_1 _1511_ (.A2(_0802_),
    .A1(_0800_),
    .B1(_0805_),
    .X(_0806_));
 sg13g2_nor3_2 _1512_ (.A(net63),
    .B(net62),
    .C(\bitserial_cipher.datapath.round_counter[4] ),
    .Y(_0807_));
 sg13g2_nor2_1 _1513_ (.A(_0807_),
    .B(_0782_),
    .Y(_0808_));
 sg13g2_and2_1 _1514_ (.A(_0598_),
    .B(_0596_),
    .X(_0809_));
 sg13g2_nand2_1 _1515_ (.Y(_0810_),
    .A(net60),
    .B(_0002_));
 sg13g2_nor2b_1 _1516_ (.A(net63),
    .B_N(net62),
    .Y(_0811_));
 sg13g2_nand2b_1 _1517_ (.Y(_0812_),
    .B(_0596_),
    .A_N(\bitserial_cipher.datapath.round_counter[1] ));
 sg13g2_nor2b_1 _1518_ (.A(_0002_),
    .B_N(_0781_),
    .Y(_0813_));
 sg13g2_a221oi_1 _1519_ (.B2(_0796_),
    .C1(_0813_),
    .B1(_0812_),
    .A1(_0810_),
    .Y(_0814_),
    .A2(_0811_));
 sg13g2_or3_1 _1520_ (.A(_0805_),
    .B(_0809_),
    .C(_0814_),
    .X(_0815_));
 sg13g2_nand2b_1 _1521_ (.Y(_0816_),
    .B(net21),
    .A_N(_0791_));
 sg13g2_buf_1 _1522_ (.A(_0789_),
    .X(_0817_));
 sg13g2_buf_8 _1523_ (.A(_0003_),
    .X(_0818_));
 sg13g2_nand2b_1 _1524_ (.Y(_0819_),
    .B(net59),
    .A_N(net20));
 sg13g2_a21oi_1 _1525_ (.A1(_0804_),
    .A2(_0816_),
    .Y(_0820_),
    .B1(_0819_));
 sg13g2_or4_1 _1526_ (.A(_0779_),
    .B(_0789_),
    .C(_0003_),
    .D(_0791_),
    .X(_0286_));
 sg13g2_nand3_1 _1527_ (.B(net59),
    .C(_0791_),
    .A(net20),
    .Y(_0287_));
 sg13g2_or2_1 _1528_ (.X(_0288_),
    .B(net61),
    .A(net22));
 sg13g2_a21oi_1 _1529_ (.A1(_0286_),
    .A2(_0287_),
    .Y(_0289_),
    .B1(_0288_));
 sg13g2_and3_1 _1530_ (.X(_0290_),
    .A(_0548_),
    .B(_0560_),
    .C(_0771_));
 sg13g2_o21ai_1 _1531_ (.B1(_0290_),
    .Y(_0291_),
    .A1(_0820_),
    .A2(_0289_));
 sg13g2_a221oi_1 _1532_ (.B2(_0815_),
    .C1(_0291_),
    .B1(_0808_),
    .A1(_0795_),
    .Y(_0292_),
    .A2(_0806_));
 sg13g2_xnor2_1 _1533_ (.Y(_0293_),
    .A(net21),
    .B(net59));
 sg13g2_nor2_1 _1534_ (.A(net20),
    .B(_0293_),
    .Y(_0294_));
 sg13g2_inv_1 _1535_ (.Y(_0295_),
    .A(net20));
 sg13g2_nor2_1 _1536_ (.A(_0295_),
    .B(_0818_),
    .Y(_0296_));
 sg13g2_nand2_1 _1537_ (.Y(_0297_),
    .A(_0791_),
    .B(_0804_));
 sg13g2_mux2_1 _1538_ (.A0(_0294_),
    .A1(_0296_),
    .S(_0297_),
    .X(_0298_));
 sg13g2_nor3_1 _1539_ (.A(_0601_),
    .B(_0793_),
    .C(_0805_),
    .Y(_0299_));
 sg13g2_nand3_1 _1540_ (.B(_0298_),
    .C(_0299_),
    .A(_0290_),
    .Y(_0300_));
 sg13g2_nand2b_1 _1541_ (.Y(_0301_),
    .B(_0300_),
    .A_N(_0292_));
 sg13g2_and2_1 _1542_ (.A(_0786_),
    .B(_0002_),
    .X(_0302_));
 sg13g2_nor2b_1 _1543_ (.A(net62),
    .B_N(_0596_),
    .Y(_0303_));
 sg13g2_nor2b_1 _1544_ (.A(_0784_),
    .B_N(_0002_),
    .Y(_0304_));
 sg13g2_nor4_1 _1545_ (.A(_0809_),
    .B(_0302_),
    .C(_0303_),
    .D(_0304_),
    .Y(_0305_));
 sg13g2_or2_1 _1546_ (.X(_0306_),
    .B(_0797_),
    .A(_0787_));
 sg13g2_nor2_1 _1547_ (.A(_0002_),
    .B(_0801_),
    .Y(_0307_));
 sg13g2_a221oi_1 _1548_ (.B2(_0780_),
    .C1(_0307_),
    .B1(_0306_),
    .A1(net22),
    .Y(_0308_),
    .A2(_0305_));
 sg13g2_o21ai_1 _1549_ (.B1(_0808_),
    .Y(_0309_),
    .A1(_0805_),
    .A2(_0308_));
 sg13g2_a21o_1 _1550_ (.A2(_0804_),
    .A1(_0803_),
    .B1(_0785_),
    .X(_0310_));
 sg13g2_nand3_1 _1551_ (.B(_0784_),
    .C(_0310_),
    .A(_0676_),
    .Y(_0311_));
 sg13g2_nand3_1 _1552_ (.B(_0782_),
    .C(_0311_),
    .A(net60),
    .Y(_0312_));
 sg13g2_nand3_1 _1553_ (.B(_0818_),
    .C(_0297_),
    .A(_0817_),
    .Y(_0313_));
 sg13g2_nand4_1 _1554_ (.B(_0791_),
    .C(_0804_),
    .A(_0295_),
    .Y(_0314_),
    .D(_0293_));
 sg13g2_nand2_1 _1555_ (.Y(_0315_),
    .A(_0310_),
    .B(_0797_));
 sg13g2_nor2b_1 _1556_ (.A(net60),
    .B_N(_0779_),
    .Y(_0316_));
 sg13g2_o21ai_1 _1557_ (.B1(_0781_),
    .Y(_0317_),
    .A1(_0783_),
    .A2(_0316_));
 sg13g2_nand2b_1 _1558_ (.Y(_0318_),
    .B(_0783_),
    .A_N(_0601_));
 sg13g2_a21oi_1 _1559_ (.A1(_0596_),
    .A2(_0318_),
    .Y(_0319_),
    .B1(\bitserial_cipher.datapath.round_counter[6] ));
 sg13g2_o21ai_1 _1560_ (.B1(_0290_),
    .Y(_0320_),
    .A1(_0317_),
    .A2(_0319_));
 sg13g2_a221oi_1 _1561_ (.B2(_0794_),
    .C1(_0320_),
    .B1(_0315_),
    .A1(_0313_),
    .Y(_0321_),
    .A2(_0314_));
 sg13g2_and3_1 _1562_ (.X(_0322_),
    .A(_0309_),
    .B(_0312_),
    .C(_0321_));
 sg13g2_nor3_1 _1563_ (.A(\bitserial_cipher.datapath.round_counter[1] ),
    .B(_0598_),
    .C(_0789_),
    .Y(_0323_));
 sg13g2_nand3_1 _1564_ (.B(_0807_),
    .C(_0323_),
    .A(net59),
    .Y(_0324_));
 sg13g2_nor2b_1 _1565_ (.A(\bitserial_cipher.bit_counter[0] ),
    .B_N(\bitserial_cipher.key_exp.lut_ff3 ),
    .Y(_0325_));
 sg13g2_xor2_1 _1566_ (.B(\bitserial_cipher.key_exp.shift_out1 ),
    .A(\bitserial_cipher.datapath.key_in ),
    .X(_0326_));
 sg13g2_nand3_1 _1567_ (.B(_0771_),
    .C(_0326_),
    .A(_0560_),
    .Y(_0327_));
 sg13g2_a21oi_1 _1568_ (.A1(_0324_),
    .A2(_0325_),
    .Y(_0328_),
    .B1(_0327_));
 sg13g2_nand2_1 _1569_ (.Y(_0329_),
    .A(_0560_),
    .B(_0771_));
 sg13g2_nor2_1 _1570_ (.A(_0329_),
    .B(_0326_),
    .Y(_0330_));
 sg13g2_a21oi_1 _1571_ (.A1(_0548_),
    .A2(_0324_),
    .Y(_0331_),
    .B1(_0768_));
 sg13g2_mux2_1 _1572_ (.A0(_0328_),
    .A1(_0330_),
    .S(_0331_),
    .X(_0332_));
 sg13g2_and2_1 _1573_ (.A(_0324_),
    .B(_0325_),
    .X(_0333_));
 sg13g2_nand2_1 _1574_ (.Y(_0334_),
    .A(\bitserial_cipher.key_exp.fifo_ff3 ),
    .B(_0326_));
 sg13g2_nand2b_1 _1575_ (.Y(_0335_),
    .B(_0768_),
    .A_N(_0326_));
 sg13g2_a22oi_1 _1576_ (.Y(_0336_),
    .B1(_0334_),
    .B2(_0335_),
    .A2(_0771_),
    .A1(_0560_));
 sg13g2_a21o_1 _1577_ (.A2(_0330_),
    .A1(_0333_),
    .B1(_0336_),
    .X(_0337_));
 sg13g2_nand3_1 _1578_ (.B(net1),
    .C(_0773_),
    .A(_0547_),
    .Y(_0338_));
 sg13g2_nor3_1 _1579_ (.A(_0332_),
    .B(_0337_),
    .C(_0338_),
    .Y(_0339_));
 sg13g2_o21ai_1 _1580_ (.B1(_0339_),
    .Y(_0340_),
    .A1(_0301_),
    .A2(_0322_));
 sg13g2_nor2_1 _1581_ (.A(_0332_),
    .B(_0337_),
    .Y(_0341_));
 sg13g2_or4_1 _1582_ (.A(_0301_),
    .B(_0322_),
    .C(_0341_),
    .D(_0338_),
    .X(_0342_));
 sg13g2_nand3_1 _1583_ (.B(\bitserial_cipher.key_exp.lut_ff3 ),
    .C(_0774_),
    .A(net69),
    .Y(_0343_));
 sg13g2_nand3_1 _1584_ (.B(_0342_),
    .C(_0343_),
    .A(_0340_),
    .Y(_0154_));
 sg13g2_nand3_1 _1585_ (.B(\bitserial_cipher.bit_counter[5] ),
    .C(_0583_),
    .A(\bitserial_cipher.bit_counter[4] ),
    .Y(_0344_));
 sg13g2_buf_2 _1586_ (.A(_0344_),
    .X(_0345_));
 sg13g2_buf_1 _1587_ (.A(_0345_),
    .X(_0346_));
 sg13g2_nand3_1 _1588_ (.B(_0580_),
    .C(net5),
    .A(net43),
    .Y(_0347_));
 sg13g2_o21ai_1 _1589_ (.B1(_0347_),
    .Y(_0348_),
    .A1(net43),
    .A2(net5));
 sg13g2_and2_1 _1590_ (.A(net23),
    .B(_0348_),
    .X(_0155_));
 sg13g2_buf_1 _1591_ (.A(net68),
    .X(_0349_));
 sg13g2_xnor2_1 _1592_ (.Y(_0350_),
    .A(net60),
    .B(net43));
 sg13g2_nand3_1 _1593_ (.B(_0580_),
    .C(net5),
    .A(net60),
    .Y(_0351_));
 sg13g2_o21ai_1 _1594_ (.B1(_0351_),
    .Y(_0352_),
    .A1(net5),
    .A2(_0350_));
 sg13g2_and2_1 _1595_ (.A(net19),
    .B(_0352_),
    .X(_0156_));
 sg13g2_nand2_1 _1596_ (.Y(_0353_),
    .A(net60),
    .B(net43));
 sg13g2_xnor2_1 _1597_ (.Y(_0354_),
    .A(_0791_),
    .B(_0353_));
 sg13g2_nand3_1 _1598_ (.B(_0580_),
    .C(_0345_),
    .A(net21),
    .Y(_0355_));
 sg13g2_o21ai_1 _1599_ (.B1(_0355_),
    .Y(_0356_),
    .A1(net5),
    .A2(_0354_));
 sg13g2_and2_1 _1600_ (.A(net19),
    .B(_0356_),
    .X(_0157_));
 sg13g2_nand2_1 _1601_ (.Y(_0357_),
    .A(net21),
    .B(_0797_));
 sg13g2_xor2_1 _1602_ (.B(_0357_),
    .A(net22),
    .X(_0358_));
 sg13g2_nand3_1 _1603_ (.B(_0580_),
    .C(_0345_),
    .A(net22),
    .Y(_0359_));
 sg13g2_o21ai_1 _1604_ (.B1(_0359_),
    .Y(_0360_),
    .A1(net5),
    .A2(_0358_));
 sg13g2_and2_1 _1605_ (.A(_0349_),
    .B(_0360_),
    .X(_0158_));
 sg13g2_nand2_1 _1606_ (.Y(_0361_),
    .A(net22),
    .B(net21));
 sg13g2_nor2_1 _1607_ (.A(_0361_),
    .B(_0353_),
    .Y(_0362_));
 sg13g2_nand2_1 _1608_ (.Y(_0363_),
    .A(_0580_),
    .B(_0345_));
 sg13g2_o21ai_1 _1609_ (.B1(_0363_),
    .Y(_0364_),
    .A1(_0346_),
    .A2(_0362_));
 sg13g2_nor4_1 _1610_ (.A(net61),
    .B(_0361_),
    .C(net5),
    .D(_0353_),
    .Y(_0365_));
 sg13g2_a21oi_1 _1611_ (.A1(net61),
    .A2(_0364_),
    .Y(_0366_),
    .B1(_0365_));
 sg13g2_nor2b_1 _1612_ (.A(_0366_),
    .B_N(_0556_),
    .Y(_0159_));
 sg13g2_nand4_1 _1613_ (.B(net21),
    .C(net61),
    .A(net22),
    .Y(_0367_),
    .D(_0797_));
 sg13g2_nand2b_1 _1614_ (.Y(_0368_),
    .B(_0367_),
    .A_N(_0345_));
 sg13g2_nand2_1 _1615_ (.Y(_0369_),
    .A(_0363_),
    .B(_0368_));
 sg13g2_nor3_1 _1616_ (.A(net20),
    .B(_0346_),
    .C(_0367_),
    .Y(_0370_));
 sg13g2_a21oi_1 _1617_ (.A1(net20),
    .A2(_0369_),
    .Y(_0371_),
    .B1(_0370_));
 sg13g2_nor2b_1 _1618_ (.A(_0371_),
    .B_N(_0556_),
    .Y(_0160_));
 sg13g2_nand3_1 _1619_ (.B(net61),
    .C(_0362_),
    .A(net20),
    .Y(_0372_));
 sg13g2_xnor2_1 _1620_ (.Y(_0373_),
    .A(net59),
    .B(_0372_));
 sg13g2_nand3_1 _1621_ (.B(_0580_),
    .C(_0345_),
    .A(\bitserial_cipher.datapath.round_counter[6] ),
    .Y(_0374_));
 sg13g2_o21ai_1 _1622_ (.B1(_0374_),
    .Y(_0375_),
    .A1(net5),
    .A2(_0373_));
 sg13g2_and2_1 _1623_ (.A(_0349_),
    .B(_0375_),
    .X(_0161_));
 sg13g2_mux2_1 _1624_ (.A0(\bitserial_cipher.key_exp.shift_out1 ),
    .A1(\bitserial_cipher.key_exp.shifter1[1] ),
    .S(net46),
    .X(_0376_));
 sg13g2_and2_1 _1625_ (.A(net19),
    .B(_0376_),
    .X(_0162_));
 sg13g2_mux2_1 _1626_ (.A0(\bitserial_cipher.key_exp.shifter1[10] ),
    .A1(\bitserial_cipher.key_exp.shifter1[11] ),
    .S(net46),
    .X(_0377_));
 sg13g2_and2_1 _1627_ (.A(net19),
    .B(_0377_),
    .X(_0163_));
 sg13g2_buf_1 _1628_ (.A(net71),
    .X(_0378_));
 sg13g2_mux2_1 _1629_ (.A0(\bitserial_cipher.key_exp.shifter1[11] ),
    .A1(\bitserial_cipher.key_exp.shifter1[12] ),
    .S(net18),
    .X(_0379_));
 sg13g2_and2_1 _1630_ (.A(net19),
    .B(_0379_),
    .X(_0164_));
 sg13g2_mux2_1 _1631_ (.A0(\bitserial_cipher.key_exp.shifter1[12] ),
    .A1(\bitserial_cipher.key_exp.shifter1[13] ),
    .S(net18),
    .X(_0380_));
 sg13g2_and2_1 _1632_ (.A(net19),
    .B(_0380_),
    .X(_0165_));
 sg13g2_mux2_1 _1633_ (.A0(\bitserial_cipher.key_exp.shifter1[13] ),
    .A1(\bitserial_cipher.key_exp.shifter1[14] ),
    .S(_0378_),
    .X(_0381_));
 sg13g2_and2_1 _1634_ (.A(net19),
    .B(_0381_),
    .X(_0166_));
 sg13g2_mux2_1 _1635_ (.A0(\bitserial_cipher.key_exp.shifter1[14] ),
    .A1(\bitserial_cipher.key_exp.shifter1[15] ),
    .S(_0378_),
    .X(_0382_));
 sg13g2_and2_1 _1636_ (.A(net19),
    .B(_0382_),
    .X(_0167_));
 sg13g2_buf_1 _1637_ (.A(net68),
    .X(_0383_));
 sg13g2_mux2_1 _1638_ (.A0(\bitserial_cipher.key_exp.shifter1[15] ),
    .A1(\bitserial_cipher.key_exp.shifter1[16] ),
    .S(net18),
    .X(_0384_));
 sg13g2_and2_1 _1639_ (.A(net17),
    .B(_0384_),
    .X(_0168_));
 sg13g2_mux2_1 _1640_ (.A0(\bitserial_cipher.key_exp.shifter1[16] ),
    .A1(\bitserial_cipher.key_exp.shifter1[17] ),
    .S(net18),
    .X(_0385_));
 sg13g2_and2_1 _1641_ (.A(net17),
    .B(_0385_),
    .X(_0169_));
 sg13g2_mux2_1 _1642_ (.A0(\bitserial_cipher.key_exp.shifter1[17] ),
    .A1(\bitserial_cipher.key_exp.shifter1[18] ),
    .S(net18),
    .X(_0386_));
 sg13g2_and2_1 _1643_ (.A(_0383_),
    .B(_0386_),
    .X(_0170_));
 sg13g2_mux2_1 _1644_ (.A0(\bitserial_cipher.key_exp.shifter1[18] ),
    .A1(\bitserial_cipher.key_exp.shifter1[19] ),
    .S(net18),
    .X(_0387_));
 sg13g2_and2_1 _1645_ (.A(net17),
    .B(_0387_),
    .X(_0171_));
 sg13g2_mux2_1 _1646_ (.A0(\bitserial_cipher.key_exp.shifter1[19] ),
    .A1(\bitserial_cipher.key_exp.shifter1[20] ),
    .S(net18),
    .X(_0388_));
 sg13g2_and2_1 _1647_ (.A(net17),
    .B(_0388_),
    .X(_0172_));
 sg13g2_mux2_1 _1648_ (.A0(\bitserial_cipher.key_exp.shifter1[1] ),
    .A1(\bitserial_cipher.key_exp.shifter1[2] ),
    .S(net18),
    .X(_0389_));
 sg13g2_and2_1 _1649_ (.A(_0383_),
    .B(_0389_),
    .X(_0173_));
 sg13g2_buf_1 _1650_ (.A(net71),
    .X(_0390_));
 sg13g2_mux2_1 _1651_ (.A0(\bitserial_cipher.key_exp.shifter1[20] ),
    .A1(\bitserial_cipher.key_exp.shifter1[21] ),
    .S(net16),
    .X(_0391_));
 sg13g2_and2_1 _1652_ (.A(net17),
    .B(_0391_),
    .X(_0174_));
 sg13g2_mux2_1 _1653_ (.A0(\bitserial_cipher.key_exp.shifter1[21] ),
    .A1(\bitserial_cipher.key_exp.shifter1[22] ),
    .S(net16),
    .X(_0392_));
 sg13g2_and2_1 _1654_ (.A(net17),
    .B(_0392_),
    .X(_0175_));
 sg13g2_mux2_1 _1655_ (.A0(\bitserial_cipher.key_exp.shifter1[22] ),
    .A1(\bitserial_cipher.key_exp.shifter1[23] ),
    .S(net16),
    .X(_0393_));
 sg13g2_and2_1 _1656_ (.A(net17),
    .B(_0393_),
    .X(_0176_));
 sg13g2_mux2_1 _1657_ (.A0(\bitserial_cipher.key_exp.shifter1[23] ),
    .A1(\bitserial_cipher.key_exp.shifter1[24] ),
    .S(_0390_),
    .X(_0394_));
 sg13g2_and2_1 _1658_ (.A(net17),
    .B(_0394_),
    .X(_0177_));
 sg13g2_buf_1 _1659_ (.A(net68),
    .X(_0395_));
 sg13g2_mux2_1 _1660_ (.A0(\bitserial_cipher.key_exp.shifter1[24] ),
    .A1(\bitserial_cipher.key_exp.shifter1[25] ),
    .S(_0390_),
    .X(_0396_));
 sg13g2_and2_1 _1661_ (.A(net15),
    .B(_0396_),
    .X(_0178_));
 sg13g2_mux2_1 _1662_ (.A0(\bitserial_cipher.key_exp.shifter1[25] ),
    .A1(\bitserial_cipher.key_exp.shifter1[26] ),
    .S(net16),
    .X(_0397_));
 sg13g2_and2_1 _1663_ (.A(net15),
    .B(_0397_),
    .X(_0179_));
 sg13g2_mux2_1 _1664_ (.A0(\bitserial_cipher.key_exp.shifter1[26] ),
    .A1(\bitserial_cipher.key_exp.shifter1[27] ),
    .S(net16),
    .X(_0398_));
 sg13g2_and2_1 _1665_ (.A(net15),
    .B(_0398_),
    .X(_0180_));
 sg13g2_mux2_1 _1666_ (.A0(\bitserial_cipher.key_exp.shifter1[27] ),
    .A1(\bitserial_cipher.key_exp.shifter1[28] ),
    .S(net16),
    .X(_0399_));
 sg13g2_and2_1 _1667_ (.A(net15),
    .B(_0399_),
    .X(_0181_));
 sg13g2_mux2_1 _1668_ (.A0(\bitserial_cipher.key_exp.shifter1[28] ),
    .A1(\bitserial_cipher.key_exp.shifter1[29] ),
    .S(net16),
    .X(_0400_));
 sg13g2_and2_1 _1669_ (.A(net15),
    .B(_0400_),
    .X(_0182_));
 sg13g2_mux2_1 _1670_ (.A0(\bitserial_cipher.key_exp.shifter1[29] ),
    .A1(\bitserial_cipher.key_exp.shifter1[30] ),
    .S(net16),
    .X(_0401_));
 sg13g2_and2_1 _1671_ (.A(_0395_),
    .B(_0401_),
    .X(_0183_));
 sg13g2_buf_1 _1672_ (.A(net71),
    .X(_0402_));
 sg13g2_mux2_1 _1673_ (.A0(\bitserial_cipher.key_exp.shifter1[2] ),
    .A1(\bitserial_cipher.key_exp.shifter1[3] ),
    .S(net14),
    .X(_0403_));
 sg13g2_and2_1 _1674_ (.A(net15),
    .B(_0403_),
    .X(_0184_));
 sg13g2_mux2_1 _1675_ (.A0(\bitserial_cipher.key_exp.shifter1[30] ),
    .A1(\bitserial_cipher.key_exp.shifter1[31] ),
    .S(net14),
    .X(_0404_));
 sg13g2_and2_1 _1676_ (.A(net15),
    .B(_0404_),
    .X(_0185_));
 sg13g2_mux2_1 _1677_ (.A0(\bitserial_cipher.key_exp.shifter1[31] ),
    .A1(\bitserial_cipher.key_exp.shifter1[32] ),
    .S(net14),
    .X(_0405_));
 sg13g2_and2_1 _1678_ (.A(_0395_),
    .B(_0405_),
    .X(_0186_));
 sg13g2_mux2_1 _1679_ (.A0(\bitserial_cipher.key_exp.shifter1[32] ),
    .A1(\bitserial_cipher.key_exp.shifter1[33] ),
    .S(net14),
    .X(_0406_));
 sg13g2_and2_1 _1680_ (.A(net15),
    .B(_0406_),
    .X(_0187_));
 sg13g2_buf_1 _1681_ (.A(_0713_),
    .X(_0407_));
 sg13g2_mux2_1 _1682_ (.A0(\bitserial_cipher.key_exp.shifter1[33] ),
    .A1(\bitserial_cipher.key_exp.shifter1[34] ),
    .S(net14),
    .X(_0408_));
 sg13g2_and2_1 _1683_ (.A(net13),
    .B(_0408_),
    .X(_0188_));
 sg13g2_mux2_1 _1684_ (.A0(\bitserial_cipher.key_exp.shifter1[34] ),
    .A1(\bitserial_cipher.key_exp.shifter1[35] ),
    .S(net14),
    .X(_0409_));
 sg13g2_and2_1 _1685_ (.A(net13),
    .B(_0409_),
    .X(_0189_));
 sg13g2_mux2_1 _1686_ (.A0(\bitserial_cipher.key_exp.shifter1[35] ),
    .A1(\bitserial_cipher.key_exp.shifter1[36] ),
    .S(net14),
    .X(_0410_));
 sg13g2_and2_1 _1687_ (.A(net13),
    .B(_0410_),
    .X(_0190_));
 sg13g2_mux2_1 _1688_ (.A0(\bitserial_cipher.key_exp.shifter1[36] ),
    .A1(\bitserial_cipher.key_exp.shifter1[37] ),
    .S(net14),
    .X(_0411_));
 sg13g2_and2_1 _1689_ (.A(net13),
    .B(_0411_),
    .X(_0191_));
 sg13g2_mux2_1 _1690_ (.A0(\bitserial_cipher.key_exp.shifter1[37] ),
    .A1(\bitserial_cipher.key_exp.shifter1[38] ),
    .S(_0402_),
    .X(_0412_));
 sg13g2_and2_1 _1691_ (.A(net13),
    .B(_0412_),
    .X(_0192_));
 sg13g2_mux2_1 _1692_ (.A0(\bitserial_cipher.key_exp.shifter1[38] ),
    .A1(\bitserial_cipher.key_exp.shifter1[39] ),
    .S(_0402_),
    .X(_0413_));
 sg13g2_and2_1 _1693_ (.A(net13),
    .B(_0413_),
    .X(_0193_));
 sg13g2_buf_1 _1694_ (.A(net71),
    .X(_0414_));
 sg13g2_mux2_1 _1695_ (.A0(\bitserial_cipher.key_exp.shifter1[39] ),
    .A1(\bitserial_cipher.key_exp.shifter1[40] ),
    .S(net12),
    .X(_0415_));
 sg13g2_and2_1 _1696_ (.A(net13),
    .B(_0415_),
    .X(_0194_));
 sg13g2_mux2_1 _1697_ (.A0(\bitserial_cipher.key_exp.shifter1[3] ),
    .A1(\bitserial_cipher.key_exp.shifter1[4] ),
    .S(_0414_),
    .X(_0416_));
 sg13g2_and2_1 _1698_ (.A(net13),
    .B(_0416_),
    .X(_0195_));
 sg13g2_mux2_1 _1699_ (.A0(\bitserial_cipher.key_exp.shifter1[40] ),
    .A1(\bitserial_cipher.key_exp.shifter1[41] ),
    .S(net12),
    .X(_0417_));
 sg13g2_and2_1 _1700_ (.A(_0407_),
    .B(_0417_),
    .X(_0196_));
 sg13g2_mux2_1 _1701_ (.A0(\bitserial_cipher.key_exp.shifter1[41] ),
    .A1(\bitserial_cipher.key_exp.shifter1[42] ),
    .S(net12),
    .X(_0418_));
 sg13g2_and2_1 _1702_ (.A(_0407_),
    .B(_0418_),
    .X(_0197_));
 sg13g2_buf_1 _1703_ (.A(_0713_),
    .X(_0419_));
 sg13g2_mux2_1 _1704_ (.A0(\bitserial_cipher.key_exp.shifter1[42] ),
    .A1(\bitserial_cipher.key_exp.shifter1[43] ),
    .S(net12),
    .X(_0420_));
 sg13g2_and2_1 _1705_ (.A(net11),
    .B(_0420_),
    .X(_0198_));
 sg13g2_mux2_1 _1706_ (.A0(\bitserial_cipher.key_exp.shifter1[43] ),
    .A1(\bitserial_cipher.key_exp.shifter1[44] ),
    .S(_0414_),
    .X(_0421_));
 sg13g2_and2_1 _1707_ (.A(net11),
    .B(_0421_),
    .X(_0199_));
 sg13g2_mux2_1 _1708_ (.A0(\bitserial_cipher.key_exp.shifter1[44] ),
    .A1(\bitserial_cipher.key_exp.shifter1[45] ),
    .S(net12),
    .X(_0422_));
 sg13g2_and2_1 _1709_ (.A(net11),
    .B(_0422_),
    .X(_0200_));
 sg13g2_mux2_1 _1710_ (.A0(\bitserial_cipher.key_exp.shifter1[45] ),
    .A1(\bitserial_cipher.key_exp.shifter1[46] ),
    .S(net12),
    .X(_0423_));
 sg13g2_and2_1 _1711_ (.A(net11),
    .B(_0423_),
    .X(_0201_));
 sg13g2_mux2_1 _1712_ (.A0(\bitserial_cipher.key_exp.shifter1[46] ),
    .A1(\bitserial_cipher.key_exp.shifter1[47] ),
    .S(net12),
    .X(_0424_));
 sg13g2_and2_1 _1713_ (.A(net11),
    .B(_0424_),
    .X(_0202_));
 sg13g2_mux2_1 _1714_ (.A0(\bitserial_cipher.key_exp.shifter1[47] ),
    .A1(\bitserial_cipher.key_exp.shifter1[48] ),
    .S(net12),
    .X(_0425_));
 sg13g2_and2_1 _1715_ (.A(_0419_),
    .B(_0425_),
    .X(_0203_));
 sg13g2_buf_1 _1716_ (.A(net71),
    .X(_0426_));
 sg13g2_mux2_1 _1717_ (.A0(\bitserial_cipher.key_exp.shifter1[48] ),
    .A1(\bitserial_cipher.key_exp.shifter1[49] ),
    .S(net10),
    .X(_0427_));
 sg13g2_and2_1 _1718_ (.A(_0419_),
    .B(_0427_),
    .X(_0204_));
 sg13g2_mux2_1 _1719_ (.A0(\bitserial_cipher.key_exp.shifter1[49] ),
    .A1(\bitserial_cipher.key_exp.shifter1[50] ),
    .S(net10),
    .X(_0428_));
 sg13g2_and2_1 _1720_ (.A(net11),
    .B(_0428_),
    .X(_0205_));
 sg13g2_mux2_1 _1721_ (.A0(\bitserial_cipher.key_exp.shifter1[4] ),
    .A1(\bitserial_cipher.key_exp.shifter1[5] ),
    .S(net10),
    .X(_0429_));
 sg13g2_and2_1 _1722_ (.A(net11),
    .B(_0429_),
    .X(_0206_));
 sg13g2_mux2_1 _1723_ (.A0(\bitserial_cipher.key_exp.shifter1[50] ),
    .A1(\bitserial_cipher.key_exp.shifter1[51] ),
    .S(_0426_),
    .X(_0430_));
 sg13g2_and2_1 _1724_ (.A(net11),
    .B(_0430_),
    .X(_0207_));
 sg13g2_buf_1 _1725_ (.A(net75),
    .X(_0431_));
 sg13g2_mux2_1 _1726_ (.A0(\bitserial_cipher.key_exp.shifter1[51] ),
    .A1(\bitserial_cipher.key_exp.shifter1[52] ),
    .S(_0426_),
    .X(_0432_));
 sg13g2_and2_1 _1727_ (.A(net58),
    .B(_0432_),
    .X(_0208_));
 sg13g2_mux2_1 _1728_ (.A0(\bitserial_cipher.key_exp.shifter1[52] ),
    .A1(\bitserial_cipher.key_exp.shifter1[53] ),
    .S(net10),
    .X(_0433_));
 sg13g2_and2_1 _1729_ (.A(net58),
    .B(_0433_),
    .X(_0209_));
 sg13g2_mux2_1 _1730_ (.A0(\bitserial_cipher.key_exp.shifter1[53] ),
    .A1(\bitserial_cipher.key_exp.shifter1[54] ),
    .S(net10),
    .X(_0434_));
 sg13g2_and2_1 _1731_ (.A(net58),
    .B(_0434_),
    .X(_0210_));
 sg13g2_mux2_1 _1732_ (.A0(\bitserial_cipher.key_exp.shifter1[54] ),
    .A1(\bitserial_cipher.key_exp.shifter1[55] ),
    .S(net10),
    .X(_0435_));
 sg13g2_and2_1 _1733_ (.A(net58),
    .B(_0435_),
    .X(_0211_));
 sg13g2_mux2_1 _1734_ (.A0(\bitserial_cipher.key_exp.shifter1[55] ),
    .A1(\bitserial_cipher.key_exp.shifter1[56] ),
    .S(net10),
    .X(_0436_));
 sg13g2_and2_1 _1735_ (.A(net58),
    .B(_0436_),
    .X(_0212_));
 sg13g2_mux2_1 _1736_ (.A0(\bitserial_cipher.key_exp.shifter1[56] ),
    .A1(\bitserial_cipher.key_exp.shifter1[57] ),
    .S(net10),
    .X(_0437_));
 sg13g2_and2_1 _1737_ (.A(net58),
    .B(_0437_),
    .X(_0213_));
 sg13g2_buf_1 _1738_ (.A(_0557_),
    .X(_0438_));
 sg13g2_mux2_1 _1739_ (.A0(\bitserial_cipher.key_exp.shifter1[57] ),
    .A1(\bitserial_cipher.key_exp.shifter1[58] ),
    .S(net9),
    .X(_0439_));
 sg13g2_and2_1 _1740_ (.A(net58),
    .B(_0439_),
    .X(_0214_));
 sg13g2_mux2_1 _1741_ (.A0(\bitserial_cipher.key_exp.shifter1[58] ),
    .A1(\bitserial_cipher.key_exp.shifter1[59] ),
    .S(net9),
    .X(_0440_));
 sg13g2_and2_1 _1742_ (.A(_0431_),
    .B(_0440_),
    .X(_0215_));
 sg13g2_nor2_1 _1743_ (.A(\bitserial_cipher.key_exp.fifo_ff0 ),
    .B(_0324_),
    .Y(_0441_));
 sg13g2_nand2b_1 _1744_ (.Y(_0442_),
    .B(\bitserial_cipher.datapath.round_counter[6] ),
    .A_N(net59));
 sg13g2_and3_1 _1745_ (.X(_0443_),
    .A(_0807_),
    .B(_0323_),
    .C(_0442_));
 sg13g2_nor2_1 _1746_ (.A(\bitserial_cipher.key_exp.lut_ff0 ),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_o21ai_1 _1747_ (.B1(_0771_),
    .Y(_0445_),
    .A1(_0441_),
    .A2(_0444_));
 sg13g2_and3_1 _1748_ (.X(_0446_),
    .A(_0559_),
    .B(net73),
    .C(_0445_));
 sg13g2_nor2b_1 _1749_ (.A(net73),
    .B_N(\bitserial_cipher.key_exp.shifter1[59] ),
    .Y(_0447_));
 sg13g2_o21ai_1 _1750_ (.B1(net69),
    .Y(_0448_),
    .A1(_0446_),
    .A2(_0447_));
 sg13g2_nor2b_1 _1751_ (.A(_0292_),
    .B_N(_0300_),
    .Y(_0449_));
 sg13g2_nand3_1 _1752_ (.B(_0312_),
    .C(_0321_),
    .A(_0309_),
    .Y(_0450_));
 sg13g2_nand2_1 _1753_ (.Y(_0451_),
    .A(_0543_),
    .B(\bitserial_cipher.key_exp.lut_ff0 ));
 sg13g2_nand4_1 _1754_ (.B(\bitserial_cipher.key_exp.fifo_ff0 ),
    .C(_0807_),
    .A(net59),
    .Y(_0452_),
    .D(_0323_));
 sg13g2_o21ai_1 _1755_ (.B1(_0452_),
    .Y(_0453_),
    .A1(_0443_),
    .A2(_0451_));
 sg13g2_a21oi_1 _1756_ (.A1(_0773_),
    .A2(_0453_),
    .Y(_0454_),
    .B1(_0675_));
 sg13g2_and4_1 _1757_ (.A(_0449_),
    .B(_0450_),
    .C(_0341_),
    .D(_0454_),
    .X(_0455_));
 sg13g2_o21ai_1 _1758_ (.B1(_0454_),
    .Y(_0456_),
    .A1(_0332_),
    .A2(_0337_));
 sg13g2_a21oi_1 _1759_ (.A1(_0449_),
    .A2(_0450_),
    .Y(_0457_),
    .B1(_0456_));
 sg13g2_nor3_1 _1760_ (.A(_0448_),
    .B(_0455_),
    .C(_0457_),
    .Y(_0216_));
 sg13g2_mux2_1 _1761_ (.A0(\bitserial_cipher.key_exp.shifter1[5] ),
    .A1(\bitserial_cipher.key_exp.shifter1[6] ),
    .S(net9),
    .X(_0458_));
 sg13g2_and2_1 _1762_ (.A(_0431_),
    .B(_0458_),
    .X(_0217_));
 sg13g2_mux2_1 _1763_ (.A0(\bitserial_cipher.key_exp.shifter1[6] ),
    .A1(\bitserial_cipher.key_exp.shifter1[7] ),
    .S(net9),
    .X(_0459_));
 sg13g2_and2_1 _1764_ (.A(net58),
    .B(_0459_),
    .X(_0218_));
 sg13g2_buf_1 _1765_ (.A(net75),
    .X(_0460_));
 sg13g2_mux2_1 _1766_ (.A0(\bitserial_cipher.key_exp.shifter1[7] ),
    .A1(\bitserial_cipher.key_exp.shifter1[8] ),
    .S(net9),
    .X(_0461_));
 sg13g2_and2_1 _1767_ (.A(net57),
    .B(_0461_),
    .X(_0219_));
 sg13g2_mux2_1 _1768_ (.A0(\bitserial_cipher.key_exp.shifter1[8] ),
    .A1(\bitserial_cipher.key_exp.shifter1[9] ),
    .S(net9),
    .X(_0462_));
 sg13g2_and2_1 _1769_ (.A(net57),
    .B(_0462_),
    .X(_0220_));
 sg13g2_mux2_1 _1770_ (.A0(\bitserial_cipher.key_exp.shifter1[9] ),
    .A1(\bitserial_cipher.key_exp.shifter1[10] ),
    .S(net9),
    .X(_0463_));
 sg13g2_and2_1 _1771_ (.A(net57),
    .B(_0463_),
    .X(_0221_));
 sg13g2_mux2_1 _1772_ (.A0(\bitserial_cipher.datapath.key_in ),
    .A1(\bitserial_cipher.key_exp.shifter2[1] ),
    .S(net9),
    .X(_0464_));
 sg13g2_and2_1 _1773_ (.A(net57),
    .B(_0464_),
    .X(_0222_));
 sg13g2_mux2_1 _1774_ (.A0(\bitserial_cipher.key_exp.shifter2[10] ),
    .A1(\bitserial_cipher.key_exp.shifter2[11] ),
    .S(_0438_),
    .X(_0465_));
 sg13g2_and2_1 _1775_ (.A(net57),
    .B(_0465_),
    .X(_0223_));
 sg13g2_mux2_1 _1776_ (.A0(\bitserial_cipher.key_exp.shifter2[11] ),
    .A1(\bitserial_cipher.key_exp.shifter2[12] ),
    .S(_0438_),
    .X(_0466_));
 sg13g2_and2_1 _1777_ (.A(net57),
    .B(_0466_),
    .X(_0224_));
 sg13g2_buf_1 _1778_ (.A(net71),
    .X(_0467_));
 sg13g2_mux2_1 _1779_ (.A0(\bitserial_cipher.key_exp.shifter2[12] ),
    .A1(\bitserial_cipher.key_exp.shifter2[13] ),
    .S(net8),
    .X(_0468_));
 sg13g2_and2_1 _1780_ (.A(net57),
    .B(_0468_),
    .X(_0225_));
 sg13g2_mux2_1 _1781_ (.A0(\bitserial_cipher.key_exp.shifter2[13] ),
    .A1(\bitserial_cipher.key_exp.shifter2[14] ),
    .S(_0467_),
    .X(_0469_));
 sg13g2_and2_1 _1782_ (.A(net57),
    .B(_0469_),
    .X(_0226_));
 sg13g2_mux2_1 _1783_ (.A0(\bitserial_cipher.key_exp.shifter2[14] ),
    .A1(\bitserial_cipher.key_exp.shifter2[15] ),
    .S(net8),
    .X(_0470_));
 sg13g2_and2_1 _1784_ (.A(_0460_),
    .B(_0470_),
    .X(_0227_));
 sg13g2_mux2_1 _1785_ (.A0(\bitserial_cipher.key_exp.shifter2[15] ),
    .A1(\bitserial_cipher.key_exp.shifter2[16] ),
    .S(net8),
    .X(_0471_));
 sg13g2_and2_1 _1786_ (.A(_0460_),
    .B(_0471_),
    .X(_0228_));
 sg13g2_buf_1 _1787_ (.A(net75),
    .X(_0472_));
 sg13g2_mux2_1 _1788_ (.A0(\bitserial_cipher.key_exp.shifter2[16] ),
    .A1(\bitserial_cipher.key_exp.shifter2[17] ),
    .S(_0467_),
    .X(_0473_));
 sg13g2_and2_1 _1789_ (.A(net56),
    .B(_0473_),
    .X(_0229_));
 sg13g2_mux2_1 _1790_ (.A0(\bitserial_cipher.key_exp.shifter2[17] ),
    .A1(\bitserial_cipher.key_exp.shifter2[18] ),
    .S(net8),
    .X(_0474_));
 sg13g2_and2_1 _1791_ (.A(net56),
    .B(_0474_),
    .X(_0230_));
 sg13g2_mux2_1 _1792_ (.A0(\bitserial_cipher.key_exp.shifter2[18] ),
    .A1(\bitserial_cipher.key_exp.shifter2[19] ),
    .S(net8),
    .X(_0475_));
 sg13g2_and2_1 _1793_ (.A(net56),
    .B(_0475_),
    .X(_0231_));
 sg13g2_mux2_1 _1794_ (.A0(\bitserial_cipher.key_exp.shifter2[19] ),
    .A1(\bitserial_cipher.key_exp.shifter2[20] ),
    .S(net8),
    .X(_0476_));
 sg13g2_and2_1 _1795_ (.A(net56),
    .B(_0476_),
    .X(_0232_));
 sg13g2_mux2_1 _1796_ (.A0(\bitserial_cipher.key_exp.shifter2[1] ),
    .A1(\bitserial_cipher.key_exp.shifter2[2] ),
    .S(net8),
    .X(_0477_));
 sg13g2_and2_1 _1797_ (.A(net56),
    .B(_0477_),
    .X(_0233_));
 sg13g2_mux2_1 _1798_ (.A0(\bitserial_cipher.key_exp.shifter2[20] ),
    .A1(\bitserial_cipher.key_exp.shifter2[21] ),
    .S(net8),
    .X(_0478_));
 sg13g2_and2_1 _1799_ (.A(net56),
    .B(_0478_),
    .X(_0234_));
 sg13g2_buf_1 _1800_ (.A(net71),
    .X(_0479_));
 sg13g2_mux2_1 _1801_ (.A0(\bitserial_cipher.key_exp.shifter2[21] ),
    .A1(\bitserial_cipher.key_exp.shifter2[22] ),
    .S(net7),
    .X(_0480_));
 sg13g2_and2_1 _1802_ (.A(net56),
    .B(_0480_),
    .X(_0235_));
 sg13g2_mux2_1 _1803_ (.A0(\bitserial_cipher.key_exp.shifter2[22] ),
    .A1(\bitserial_cipher.key_exp.shifter2[23] ),
    .S(net7),
    .X(_0481_));
 sg13g2_and2_1 _1804_ (.A(net56),
    .B(_0481_),
    .X(_0236_));
 sg13g2_mux2_1 _1805_ (.A0(\bitserial_cipher.key_exp.shifter2[23] ),
    .A1(\bitserial_cipher.key_exp.shifter2[24] ),
    .S(net7),
    .X(_0482_));
 sg13g2_and2_1 _1806_ (.A(_0472_),
    .B(_0482_),
    .X(_0237_));
 sg13g2_mux2_1 _1807_ (.A0(\bitserial_cipher.key_exp.shifter2[24] ),
    .A1(\bitserial_cipher.key_exp.shifter2[25] ),
    .S(net7),
    .X(_0483_));
 sg13g2_and2_1 _1808_ (.A(_0472_),
    .B(_0483_),
    .X(_0238_));
 sg13g2_buf_1 _1809_ (.A(net75),
    .X(_0484_));
 sg13g2_mux2_1 _1810_ (.A0(\bitserial_cipher.key_exp.shifter2[25] ),
    .A1(\bitserial_cipher.key_exp.shifter2[26] ),
    .S(net7),
    .X(_0485_));
 sg13g2_and2_1 _1811_ (.A(net55),
    .B(_0485_),
    .X(_0239_));
 sg13g2_mux2_1 _1812_ (.A0(\bitserial_cipher.key_exp.shifter2[26] ),
    .A1(\bitserial_cipher.key_exp.shifter2[27] ),
    .S(_0479_),
    .X(_0486_));
 sg13g2_and2_1 _1813_ (.A(net55),
    .B(_0486_),
    .X(_0240_));
 sg13g2_mux2_1 _1814_ (.A0(\bitserial_cipher.key_exp.shifter2[27] ),
    .A1(\bitserial_cipher.key_exp.shifter2[28] ),
    .S(net7),
    .X(_0487_));
 sg13g2_and2_1 _1815_ (.A(net55),
    .B(_0487_),
    .X(_0241_));
 sg13g2_mux2_1 _1816_ (.A0(\bitserial_cipher.key_exp.shifter2[28] ),
    .A1(\bitserial_cipher.key_exp.shifter2[29] ),
    .S(net7),
    .X(_0488_));
 sg13g2_and2_1 _1817_ (.A(net55),
    .B(_0488_),
    .X(_0242_));
 sg13g2_mux2_1 _1818_ (.A0(\bitserial_cipher.key_exp.shifter2[29] ),
    .A1(\bitserial_cipher.key_exp.shifter2[30] ),
    .S(net7),
    .X(_0489_));
 sg13g2_and2_1 _1819_ (.A(net55),
    .B(_0489_),
    .X(_0243_));
 sg13g2_mux2_1 _1820_ (.A0(\bitserial_cipher.key_exp.shifter2[2] ),
    .A1(\bitserial_cipher.key_exp.shifter2[3] ),
    .S(_0479_),
    .X(_0490_));
 sg13g2_and2_1 _1821_ (.A(net55),
    .B(_0490_),
    .X(_0244_));
 sg13g2_buf_1 _1822_ (.A(net71),
    .X(_0491_));
 sg13g2_mux2_1 _1823_ (.A0(\bitserial_cipher.key_exp.shifter2[30] ),
    .A1(\bitserial_cipher.key_exp.shifter2[31] ),
    .S(net6),
    .X(_0492_));
 sg13g2_and2_1 _1824_ (.A(_0484_),
    .B(_0492_),
    .X(_0245_));
 sg13g2_mux2_1 _1825_ (.A0(\bitserial_cipher.key_exp.shifter2[31] ),
    .A1(\bitserial_cipher.key_exp.shifter2[32] ),
    .S(net6),
    .X(_0493_));
 sg13g2_and2_1 _1826_ (.A(_0484_),
    .B(_0493_),
    .X(_0246_));
 sg13g2_mux2_1 _1827_ (.A0(\bitserial_cipher.key_exp.shifter2[32] ),
    .A1(\bitserial_cipher.key_exp.shifter2[33] ),
    .S(_0491_),
    .X(_0494_));
 sg13g2_and2_1 _1828_ (.A(net55),
    .B(_0494_),
    .X(_0247_));
 sg13g2_mux2_1 _1829_ (.A0(\bitserial_cipher.key_exp.shifter2[33] ),
    .A1(\bitserial_cipher.key_exp.shifter2[34] ),
    .S(net6),
    .X(_0495_));
 sg13g2_and2_1 _1830_ (.A(net55),
    .B(_0495_),
    .X(_0248_));
 sg13g2_buf_1 _1831_ (.A(net75),
    .X(_0496_));
 sg13g2_mux2_1 _1832_ (.A0(\bitserial_cipher.key_exp.shifter2[34] ),
    .A1(\bitserial_cipher.key_exp.shifter2[35] ),
    .S(net6),
    .X(_0497_));
 sg13g2_and2_1 _1833_ (.A(_0496_),
    .B(_0497_),
    .X(_0249_));
 sg13g2_mux2_1 _1834_ (.A0(\bitserial_cipher.key_exp.shifter2[35] ),
    .A1(\bitserial_cipher.key_exp.shifter2[36] ),
    .S(net6),
    .X(_0498_));
 sg13g2_and2_1 _1835_ (.A(net54),
    .B(_0498_),
    .X(_0250_));
 sg13g2_mux2_1 _1836_ (.A0(\bitserial_cipher.key_exp.shifter2[36] ),
    .A1(\bitserial_cipher.key_exp.shifter2[37] ),
    .S(net6),
    .X(_0499_));
 sg13g2_and2_1 _1837_ (.A(net54),
    .B(_0499_),
    .X(_0251_));
 sg13g2_mux2_1 _1838_ (.A0(\bitserial_cipher.key_exp.shifter2[37] ),
    .A1(\bitserial_cipher.key_exp.shifter2[38] ),
    .S(net6),
    .X(_0500_));
 sg13g2_and2_1 _1839_ (.A(net54),
    .B(_0500_),
    .X(_0252_));
 sg13g2_mux2_1 _1840_ (.A0(\bitserial_cipher.key_exp.shifter2[38] ),
    .A1(\bitserial_cipher.key_exp.shifter2[39] ),
    .S(_0491_),
    .X(_0501_));
 sg13g2_and2_1 _1841_ (.A(net54),
    .B(_0501_),
    .X(_0253_));
 sg13g2_mux2_1 _1842_ (.A0(\bitserial_cipher.key_exp.shifter2[39] ),
    .A1(\bitserial_cipher.key_exp.shifter2[40] ),
    .S(net6),
    .X(_0502_));
 sg13g2_and2_1 _1843_ (.A(_0496_),
    .B(_0502_),
    .X(_0254_));
 sg13g2_buf_1 _1844_ (.A(_0546_),
    .X(_0503_));
 sg13g2_mux2_1 _1845_ (.A0(\bitserial_cipher.key_exp.shifter2[3] ),
    .A1(\bitserial_cipher.key_exp.shifter2[4] ),
    .S(net53),
    .X(_0504_));
 sg13g2_and2_1 _1846_ (.A(net54),
    .B(_0504_),
    .X(_0255_));
 sg13g2_mux2_1 _1847_ (.A0(\bitserial_cipher.key_exp.shifter2[40] ),
    .A1(\bitserial_cipher.key_exp.shifter2[41] ),
    .S(net53),
    .X(_0505_));
 sg13g2_and2_1 _1848_ (.A(net54),
    .B(_0505_),
    .X(_0256_));
 sg13g2_mux2_1 _1849_ (.A0(\bitserial_cipher.key_exp.shifter2[41] ),
    .A1(\bitserial_cipher.key_exp.shifter2[42] ),
    .S(net53),
    .X(_0506_));
 sg13g2_and2_1 _1850_ (.A(net54),
    .B(_0506_),
    .X(_0257_));
 sg13g2_mux2_1 _1851_ (.A0(\bitserial_cipher.key_exp.shifter2[42] ),
    .A1(\bitserial_cipher.key_exp.shifter2[43] ),
    .S(net53),
    .X(_0507_));
 sg13g2_and2_1 _1852_ (.A(net54),
    .B(_0507_),
    .X(_0258_));
 sg13g2_buf_1 _1853_ (.A(_0554_),
    .X(_0508_));
 sg13g2_mux2_1 _1854_ (.A0(\bitserial_cipher.key_exp.shifter2[43] ),
    .A1(\bitserial_cipher.key_exp.shifter2[44] ),
    .S(net53),
    .X(_0509_));
 sg13g2_and2_1 _1855_ (.A(net52),
    .B(_0509_),
    .X(_0259_));
 sg13g2_mux2_1 _1856_ (.A0(\bitserial_cipher.key_exp.shifter2[44] ),
    .A1(\bitserial_cipher.key_exp.shifter2[45] ),
    .S(net53),
    .X(_0510_));
 sg13g2_and2_1 _1857_ (.A(net52),
    .B(_0510_),
    .X(_0260_));
 sg13g2_mux2_1 _1858_ (.A0(\bitserial_cipher.key_exp.shifter2[45] ),
    .A1(\bitserial_cipher.key_exp.shifter2[46] ),
    .S(net53),
    .X(_0511_));
 sg13g2_and2_1 _1859_ (.A(net52),
    .B(_0511_),
    .X(_0261_));
 sg13g2_mux2_1 _1860_ (.A0(\bitserial_cipher.key_exp.shifter2[46] ),
    .A1(\bitserial_cipher.key_exp.shifter2[47] ),
    .S(net53),
    .X(_0512_));
 sg13g2_and2_1 _1861_ (.A(net52),
    .B(_0512_),
    .X(_0262_));
 sg13g2_mux2_1 _1862_ (.A0(\bitserial_cipher.key_exp.shifter2[47] ),
    .A1(\bitserial_cipher.key_exp.shifter2[48] ),
    .S(_0503_),
    .X(_0513_));
 sg13g2_and2_1 _1863_ (.A(net52),
    .B(_0513_),
    .X(_0263_));
 sg13g2_mux2_1 _1864_ (.A0(\bitserial_cipher.key_exp.shifter2[48] ),
    .A1(\bitserial_cipher.key_exp.shifter2[49] ),
    .S(_0503_),
    .X(_0514_));
 sg13g2_and2_1 _1865_ (.A(net52),
    .B(_0514_),
    .X(_0264_));
 sg13g2_buf_1 _1866_ (.A(_0546_),
    .X(_0515_));
 sg13g2_mux2_1 _1867_ (.A0(\bitserial_cipher.key_exp.shifter2[49] ),
    .A1(\bitserial_cipher.key_exp.shifter2[50] ),
    .S(net51),
    .X(_0516_));
 sg13g2_and2_1 _1868_ (.A(_0508_),
    .B(_0516_),
    .X(_0265_));
 sg13g2_mux2_1 _1869_ (.A0(\bitserial_cipher.key_exp.shifter2[4] ),
    .A1(\bitserial_cipher.key_exp.shifter2[5] ),
    .S(net51),
    .X(_0517_));
 sg13g2_and2_1 _1870_ (.A(net52),
    .B(_0517_),
    .X(_0266_));
 sg13g2_mux2_1 _1871_ (.A0(\bitserial_cipher.key_exp.shifter2[50] ),
    .A1(\bitserial_cipher.key_exp.shifter2[51] ),
    .S(net51),
    .X(_0518_));
 sg13g2_and2_1 _1872_ (.A(_0508_),
    .B(_0518_),
    .X(_0267_));
 sg13g2_mux2_1 _1873_ (.A0(\bitserial_cipher.key_exp.shifter2[51] ),
    .A1(\bitserial_cipher.key_exp.shifter2[52] ),
    .S(net51),
    .X(_0519_));
 sg13g2_and2_1 _1874_ (.A(net52),
    .B(_0519_),
    .X(_0268_));
 sg13g2_buf_1 _1875_ (.A(_0554_),
    .X(_0520_));
 sg13g2_mux2_1 _1876_ (.A0(\bitserial_cipher.key_exp.shifter2[52] ),
    .A1(\bitserial_cipher.key_exp.shifter2[53] ),
    .S(net51),
    .X(_0521_));
 sg13g2_and2_1 _1877_ (.A(net50),
    .B(_0521_),
    .X(_0269_));
 sg13g2_mux2_1 _1878_ (.A0(\bitserial_cipher.key_exp.shifter2[53] ),
    .A1(\bitserial_cipher.key_exp.shifter2[54] ),
    .S(_0515_),
    .X(_0522_));
 sg13g2_and2_1 _1879_ (.A(net50),
    .B(_0522_),
    .X(_0270_));
 sg13g2_mux2_1 _1880_ (.A0(\bitserial_cipher.key_exp.shifter2[54] ),
    .A1(\bitserial_cipher.key_exp.shifter2[55] ),
    .S(net51),
    .X(_0523_));
 sg13g2_and2_1 _1881_ (.A(_0520_),
    .B(_0523_),
    .X(_0271_));
 sg13g2_mux2_1 _1882_ (.A0(\bitserial_cipher.key_exp.shifter2[55] ),
    .A1(\bitserial_cipher.key_exp.shifter2[56] ),
    .S(_0515_),
    .X(_0524_));
 sg13g2_and2_1 _1883_ (.A(_0520_),
    .B(_0524_),
    .X(_0272_));
 sg13g2_mux2_1 _1884_ (.A0(\bitserial_cipher.key_exp.shifter2[56] ),
    .A1(\bitserial_cipher.key_exp.shifter2[57] ),
    .S(net51),
    .X(_0525_));
 sg13g2_and2_1 _1885_ (.A(net50),
    .B(_0525_),
    .X(_0273_));
 sg13g2_mux2_1 _1886_ (.A0(\bitserial_cipher.key_exp.shifter2[57] ),
    .A1(\bitserial_cipher.key_exp.shifter2[58] ),
    .S(net51),
    .X(_0526_));
 sg13g2_and2_1 _1887_ (.A(net50),
    .B(_0526_),
    .X(_0274_));
 sg13g2_buf_1 _1888_ (.A(_0546_),
    .X(_0527_));
 sg13g2_mux2_1 _1889_ (.A0(\bitserial_cipher.key_exp.shifter2[58] ),
    .A1(\bitserial_cipher.key_exp.shifter2[59] ),
    .S(net49),
    .X(_0528_));
 sg13g2_and2_1 _1890_ (.A(net50),
    .B(_0528_),
    .X(_0275_));
 sg13g2_mux2_1 _1891_ (.A0(\bitserial_cipher.key_exp.shifter2[59] ),
    .A1(\bitserial_cipher.key_exp.shifter2[60] ),
    .S(_0527_),
    .X(_0529_));
 sg13g2_and2_1 _1892_ (.A(net50),
    .B(_0529_),
    .X(_0276_));
 sg13g2_mux2_1 _1893_ (.A0(\bitserial_cipher.key_exp.shifter2[5] ),
    .A1(\bitserial_cipher.key_exp.shifter2[6] ),
    .S(net49),
    .X(_0530_));
 sg13g2_and2_1 _1894_ (.A(net50),
    .B(_0530_),
    .X(_0277_));
 sg13g2_mux2_1 _1895_ (.A0(\bitserial_cipher.key_exp.shifter2[60] ),
    .A1(\bitserial_cipher.key_exp.shifter2[61] ),
    .S(_0527_),
    .X(_0531_));
 sg13g2_and2_1 _1896_ (.A(net50),
    .B(_0531_),
    .X(_0278_));
 sg13g2_mux2_1 _1897_ (.A0(\bitserial_cipher.key_exp.shifter2[61] ),
    .A1(\bitserial_cipher.key_exp.shifter2[62] ),
    .S(net49),
    .X(_0532_));
 sg13g2_and2_1 _1898_ (.A(net69),
    .B(_0532_),
    .X(_0279_));
 sg13g2_mux2_1 _1899_ (.A0(\bitserial_cipher.key_exp.shifter2[62] ),
    .A1(\bitserial_cipher.key_exp.shifter2[63] ),
    .S(net49),
    .X(_0533_));
 sg13g2_and2_1 _1900_ (.A(net69),
    .B(_0533_),
    .X(_0280_));
 sg13g2_nor4_1 _1901_ (.A(_0817_),
    .B(\bitserial_cipher.datapath.round_counter[6] ),
    .C(_0793_),
    .D(_0812_),
    .Y(_0534_));
 sg13g2_nor2b_1 _1902_ (.A(_0534_),
    .B_N(_0773_),
    .Y(_0535_));
 sg13g2_mux2_1 _1903_ (.A0(\bitserial_cipher.key_exp.fifo_ff0 ),
    .A1(\bitserial_cipher.key_exp.lut_ff0 ),
    .S(_0535_),
    .X(_0536_));
 sg13g2_mux2_1 _1904_ (.A0(\bitserial_cipher.key_exp.shifter2[63] ),
    .A1(_0536_),
    .S(net49),
    .X(_0537_));
 sg13g2_and2_1 _1905_ (.A(net69),
    .B(_0537_),
    .X(_0281_));
 sg13g2_mux2_1 _1906_ (.A0(\bitserial_cipher.key_exp.shifter2[6] ),
    .A1(\bitserial_cipher.key_exp.shifter2[7] ),
    .S(net49),
    .X(_0538_));
 sg13g2_and2_1 _1907_ (.A(net69),
    .B(_0538_),
    .X(_0282_));
 sg13g2_mux2_1 _1908_ (.A0(\bitserial_cipher.key_exp.shifter2[7] ),
    .A1(\bitserial_cipher.key_exp.shifter2[8] ),
    .S(net49),
    .X(_0539_));
 sg13g2_and2_1 _1909_ (.A(net69),
    .B(_0539_),
    .X(_0283_));
 sg13g2_mux2_1 _1910_ (.A0(\bitserial_cipher.key_exp.shifter2[8] ),
    .A1(\bitserial_cipher.key_exp.shifter2[9] ),
    .S(net49),
    .X(_0540_));
 sg13g2_and2_1 _1911_ (.A(_0578_),
    .B(_0540_),
    .X(_0284_));
 sg13g2_mux2_1 _1912_ (.A0(\bitserial_cipher.key_exp.shifter2[9] ),
    .A1(\bitserial_cipher.key_exp.shifter2[10] ),
    .S(net73),
    .X(_0541_));
 sg13g2_and2_1 _1913_ (.A(_0578_),
    .B(_0541_),
    .X(_0285_));
 sg13g2_nor4_1 _1914_ (.A(net22),
    .B(net20),
    .C(net61),
    .D(net59),
    .Y(_0542_));
 sg13g2_and2_1 _1915_ (.A(_0316_),
    .B(_0542_),
    .X(\bitserial_cipher.datapath.valid ));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi \bitserial_cipher.datapath.bit_counter[0]$_SDFFE_PP0P__100  (.L_HI(net100));
 sg13g2_buf_1 _1918_ (.A(net77),
    .X(\bitserial_cipher.zero ));
 sg13g2_buf_1 _1919_ (.A(net78),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1920_ (.A(net79),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1921_ (.A(net80),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1922_ (.A(net81),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1923_ (.A(net82),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1924_ (.A(net83),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1925_ (.A(net84),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1926_ (.A(net85),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1927_ (.A(net86),
    .X(uio_out[0]));
 sg13g2_buf_1 _1928_ (.A(net87),
    .X(uio_out[1]));
 sg13g2_buf_1 _1929_ (.A(net88),
    .X(uio_out[2]));
 sg13g2_buf_1 _1930_ (.A(net89),
    .X(uio_out[3]));
 sg13g2_buf_1 _1931_ (.A(net90),
    .X(uio_out[4]));
 sg13g2_buf_1 _1932_ (.A(net91),
    .X(uio_out[5]));
 sg13g2_buf_1 _1933_ (.A(net92),
    .X(uio_out[6]));
 sg13g2_buf_1 _1934_ (.A(net93),
    .X(uio_out[7]));
 sg13g2_buf_1 _1935_ (.A(\bitserial_cipher.cipher_out ),
    .X(net3));
 sg13g2_buf_1 _1936_ (.A(net94),
    .X(uo_out[1]));
 sg13g2_buf_1 _1937_ (.A(net95),
    .X(uo_out[2]));
 sg13g2_buf_1 _1938_ (.A(net96),
    .X(uo_out[3]));
 sg13g2_buf_1 _1939_ (.A(net97),
    .X(uo_out[4]));
 sg13g2_buf_1 _1940_ (.A(net98),
    .X(uo_out[5]));
 sg13g2_buf_1 _1941_ (.A(net99),
    .X(uo_out[6]));
 sg13g2_buf_1 _1942_ (.A(\bitserial_cipher.datapath.valid ),
    .X(net4));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.bit_counter[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net100),
    .D(_0005_),
    .Q_N(_0004_),
    .Q(\bitserial_cipher.bit_counter[0] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.bit_counter[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net101),
    .D(_0006_),
    .Q_N(_1096_),
    .Q(\bitserial_cipher.bit_counter[1] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.bit_counter[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net102),
    .D(_0007_),
    .Q_N(_1095_),
    .Q(\bitserial_cipher.bit_counter[2] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.bit_counter[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net103),
    .D(_0008_),
    .Q_N(_1094_),
    .Q(\bitserial_cipher.bit_counter[3] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.bit_counter[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net104),
    .D(_0009_),
    .Q_N(_1093_),
    .Q(\bitserial_cipher.bit_counter[4] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.bit_counter[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net105),
    .D(_0010_),
    .Q_N(_1092_),
    .Q(\bitserial_cipher.bit_counter[5] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.fifo_ff56$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net106),
    .D(_0011_),
    .Q_N(_1091_),
    .Q(\bitserial_cipher.datapath.fifo_ff56 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.fifo_ff57$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net107),
    .D(_0012_),
    .Q_N(_1090_),
    .Q(\bitserial_cipher.datapath.fifo_ff57 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.fifo_ff58$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net108),
    .D(_0013_),
    .Q_N(_1089_),
    .Q(\bitserial_cipher.datapath.fifo_ff58 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.fifo_ff59$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net109),
    .D(_0014_),
    .Q_N(_1088_),
    .Q(\bitserial_cipher.datapath.fifo_ff59 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.fifo_ff60$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net110),
    .D(_0015_),
    .Q_N(_1087_),
    .Q(\bitserial_cipher.datapath.fifo_ff60 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.fifo_ff61$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net111),
    .D(_0016_),
    .Q_N(_1086_),
    .Q(\bitserial_cipher.datapath.fifo_ff61 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.fifo_ff62$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net112),
    .D(_0017_),
    .Q_N(_1085_),
    .Q(\bitserial_cipher.datapath.fifo_ff62 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.fifo_ff63$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net113),
    .D(_0018_),
    .Q_N(_1084_),
    .Q(\bitserial_cipher.datapath.fifo_ff63 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.lut_ff56$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net114),
    .D(_0019_),
    .Q_N(_1083_),
    .Q(\bitserial_cipher.datapath.lut_ff56 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.lut_ff57$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net115),
    .D(_0020_),
    .Q_N(_1082_),
    .Q(\bitserial_cipher.datapath.lut_ff57 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.lut_ff58$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net116),
    .D(_0021_),
    .Q_N(_1081_),
    .Q(\bitserial_cipher.datapath.lut_ff58 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.lut_ff59$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net117),
    .D(_0022_),
    .Q_N(_1080_),
    .Q(\bitserial_cipher.datapath.lut_ff59 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.lut_ff60$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net118),
    .D(_0023_),
    .Q_N(_1079_),
    .Q(\bitserial_cipher.datapath.lut_ff60 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.lut_ff61$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net119),
    .D(_0024_),
    .Q_N(_1078_),
    .Q(\bitserial_cipher.datapath.lut_ff61 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.lut_ff62$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net120),
    .D(_0025_),
    .Q_N(_1077_),
    .Q(\bitserial_cipher.datapath.lut_ff62 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.lut_ff63$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net121),
    .D(_0026_),
    .Q_N(_1076_),
    .Q(\bitserial_cipher.datapath.lut_ff63 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net122),
    .D(_0027_),
    .Q_N(_1075_),
    .Q(\bitserial_cipher.datapath.shift_in2 ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net123),
    .D(_0028_),
    .Q_N(_1074_),
    .Q(\bitserial_cipher.datapath.shifter1[10] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net124),
    .D(_0029_),
    .Q_N(_1073_),
    .Q(\bitserial_cipher.datapath.shifter1[11] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net125),
    .D(_0030_),
    .Q_N(_1072_),
    .Q(\bitserial_cipher.datapath.shifter1[12] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net126),
    .D(_0031_),
    .Q_N(_1071_),
    .Q(\bitserial_cipher.datapath.shifter1[13] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net127),
    .D(_0032_),
    .Q_N(_1070_),
    .Q(\bitserial_cipher.datapath.shifter1[14] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net128),
    .D(_0033_),
    .Q_N(_1069_),
    .Q(\bitserial_cipher.datapath.shifter1[15] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net129),
    .D(_0034_),
    .Q_N(_1068_),
    .Q(\bitserial_cipher.datapath.shifter1[16] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net130),
    .D(_0035_),
    .Q_N(_1067_),
    .Q(\bitserial_cipher.datapath.shifter1[17] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net131),
    .D(_0036_),
    .Q_N(_1066_),
    .Q(\bitserial_cipher.datapath.shifter1[18] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net132),
    .D(_0037_),
    .Q_N(_1065_),
    .Q(\bitserial_cipher.datapath.shifter1[19] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net133),
    .D(_0038_),
    .Q_N(_1064_),
    .Q(\bitserial_cipher.datapath.shifter1[1] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net134),
    .D(_0039_),
    .Q_N(_1063_),
    .Q(\bitserial_cipher.datapath.shifter1[20] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net135),
    .D(_0040_),
    .Q_N(_1062_),
    .Q(\bitserial_cipher.datapath.shifter1[21] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net136),
    .D(_0041_),
    .Q_N(_1061_),
    .Q(\bitserial_cipher.datapath.shifter1[22] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net137),
    .D(_0042_),
    .Q_N(_1060_),
    .Q(\bitserial_cipher.datapath.shifter1[23] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net138),
    .D(_0043_),
    .Q_N(_1059_),
    .Q(\bitserial_cipher.datapath.shifter1[24] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net139),
    .D(_0044_),
    .Q_N(_1058_),
    .Q(\bitserial_cipher.datapath.shifter1[25] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net140),
    .D(_0045_),
    .Q_N(_1057_),
    .Q(\bitserial_cipher.datapath.shifter1[26] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net141),
    .D(_0046_),
    .Q_N(_1056_),
    .Q(\bitserial_cipher.datapath.shifter1[27] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net142),
    .D(_0047_),
    .Q_N(_1055_),
    .Q(\bitserial_cipher.datapath.shifter1[28] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net143),
    .D(_0048_),
    .Q_N(_1054_),
    .Q(\bitserial_cipher.datapath.shifter1[29] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net144),
    .D(_0049_),
    .Q_N(_1053_),
    .Q(\bitserial_cipher.datapath.shifter1[2] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net145),
    .D(_0050_),
    .Q_N(_1052_),
    .Q(\bitserial_cipher.datapath.shifter1[30] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net146),
    .D(_0051_),
    .Q_N(_1051_),
    .Q(\bitserial_cipher.datapath.shifter1[31] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net147),
    .D(_0052_),
    .Q_N(_1050_),
    .Q(\bitserial_cipher.datapath.shifter1[32] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net148),
    .D(_0053_),
    .Q_N(_1049_),
    .Q(\bitserial_cipher.datapath.shifter1[33] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net149),
    .D(_0054_),
    .Q_N(_1048_),
    .Q(\bitserial_cipher.datapath.shifter1[34] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net150),
    .D(_0055_),
    .Q_N(_1047_),
    .Q(\bitserial_cipher.datapath.shifter1[35] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net151),
    .D(_0056_),
    .Q_N(_1046_),
    .Q(\bitserial_cipher.datapath.shifter1[36] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net152),
    .D(_0057_),
    .Q_N(_1045_),
    .Q(\bitserial_cipher.datapath.shifter1[37] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net153),
    .D(_0058_),
    .Q_N(_1044_),
    .Q(\bitserial_cipher.datapath.shifter1[38] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net154),
    .D(_0059_),
    .Q_N(_1043_),
    .Q(\bitserial_cipher.datapath.shifter1[39] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net155),
    .D(_0060_),
    .Q_N(_1042_),
    .Q(\bitserial_cipher.datapath.shifter1[3] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net156),
    .D(_0061_),
    .Q_N(_1041_),
    .Q(\bitserial_cipher.datapath.shifter1[40] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net157),
    .D(_0062_),
    .Q_N(_1040_),
    .Q(\bitserial_cipher.datapath.shifter1[41] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net158),
    .D(_0063_),
    .Q_N(_1039_),
    .Q(\bitserial_cipher.datapath.shifter1[42] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net159),
    .D(_0064_),
    .Q_N(_1038_),
    .Q(\bitserial_cipher.datapath.shifter1[43] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net160),
    .D(_0065_),
    .Q_N(_1037_),
    .Q(\bitserial_cipher.datapath.shifter1[44] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net161),
    .D(_0066_),
    .Q_N(_1036_),
    .Q(\bitserial_cipher.datapath.shifter1[45] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net162),
    .D(_0067_),
    .Q_N(_1035_),
    .Q(\bitserial_cipher.datapath.shifter1[46] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net163),
    .D(_0068_),
    .Q_N(_1034_),
    .Q(\bitserial_cipher.datapath.shifter1[47] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net164),
    .D(_0069_),
    .Q_N(_1033_),
    .Q(\bitserial_cipher.datapath.shifter1[48] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net165),
    .D(_0070_),
    .Q_N(_1032_),
    .Q(\bitserial_cipher.datapath.shifter1[49] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net166),
    .D(_0071_),
    .Q_N(_1031_),
    .Q(\bitserial_cipher.datapath.shifter1[4] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net167),
    .D(_0072_),
    .Q_N(_1030_),
    .Q(\bitserial_cipher.datapath.shifter1[50] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net168),
    .D(_0073_),
    .Q_N(_1029_),
    .Q(\bitserial_cipher.datapath.shifter1[51] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net169),
    .D(_0074_),
    .Q_N(_1028_),
    .Q(\bitserial_cipher.datapath.shifter1[52] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net170),
    .D(_0075_),
    .Q_N(_1027_),
    .Q(\bitserial_cipher.datapath.shifter1[53] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net171),
    .D(_0076_),
    .Q_N(_1026_),
    .Q(\bitserial_cipher.datapath.shifter1[54] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net172),
    .D(_0077_),
    .Q_N(_1025_),
    .Q(\bitserial_cipher.datapath.shifter1[55] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net173),
    .D(_0078_),
    .Q_N(_1024_),
    .Q(\bitserial_cipher.datapath.shifter1[5] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net174),
    .D(_0079_),
    .Q_N(_1023_),
    .Q(\bitserial_cipher.datapath.shifter1[6] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net175),
    .D(_0080_),
    .Q_N(_1022_),
    .Q(\bitserial_cipher.datapath.shifter1[7] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net176),
    .D(_0081_),
    .Q_N(_1021_),
    .Q(\bitserial_cipher.datapath.shifter1[8] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net177),
    .D(_0082_),
    .Q_N(_1020_),
    .Q(\bitserial_cipher.datapath.shifter1[9] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net178),
    .D(_0083_),
    .Q_N(_1019_),
    .Q(\bitserial_cipher.cipher_out ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net179),
    .D(_0084_),
    .Q_N(_1018_),
    .Q(\bitserial_cipher.datapath.shifter2[10] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net180),
    .D(_0085_),
    .Q_N(_1017_),
    .Q(\bitserial_cipher.datapath.shifter2[11] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net181),
    .D(_0086_),
    .Q_N(_1016_),
    .Q(\bitserial_cipher.datapath.shifter2[12] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net182),
    .D(_0087_),
    .Q_N(_1015_),
    .Q(\bitserial_cipher.datapath.shifter2[13] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net183),
    .D(_0088_),
    .Q_N(_1014_),
    .Q(\bitserial_cipher.datapath.shifter2[14] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net184),
    .D(_0089_),
    .Q_N(_1013_),
    .Q(\bitserial_cipher.datapath.shifter2[15] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net185),
    .D(_0090_),
    .Q_N(_1012_),
    .Q(\bitserial_cipher.datapath.shifter2[16] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net186),
    .D(_0091_),
    .Q_N(_1011_),
    .Q(\bitserial_cipher.datapath.shifter2[17] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net187),
    .D(_0092_),
    .Q_N(_1010_),
    .Q(\bitserial_cipher.datapath.shifter2[18] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net188),
    .D(_0093_),
    .Q_N(_1009_),
    .Q(\bitserial_cipher.datapath.shifter2[19] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net189),
    .D(_0094_),
    .Q_N(_1008_),
    .Q(\bitserial_cipher.datapath.shifter2[1] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net190),
    .D(_0095_),
    .Q_N(_1007_),
    .Q(\bitserial_cipher.datapath.shifter2[20] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net191),
    .D(_0096_),
    .Q_N(_1006_),
    .Q(\bitserial_cipher.datapath.shifter2[21] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net192),
    .D(_0097_),
    .Q_N(_1005_),
    .Q(\bitserial_cipher.datapath.shifter2[22] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net193),
    .D(_0098_),
    .Q_N(_1004_),
    .Q(\bitserial_cipher.datapath.shifter2[23] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net194),
    .D(_0099_),
    .Q_N(_1003_),
    .Q(\bitserial_cipher.datapath.shifter2[24] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net195),
    .D(_0100_),
    .Q_N(_1002_),
    .Q(\bitserial_cipher.datapath.shifter2[25] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net196),
    .D(_0101_),
    .Q_N(_1001_),
    .Q(\bitserial_cipher.datapath.shifter2[26] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net197),
    .D(_0102_),
    .Q_N(_1000_),
    .Q(\bitserial_cipher.datapath.shifter2[27] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net198),
    .D(_0103_),
    .Q_N(_0999_),
    .Q(\bitserial_cipher.datapath.shifter2[28] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net199),
    .D(_0104_),
    .Q_N(_0998_),
    .Q(\bitserial_cipher.datapath.shifter2[29] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net200),
    .D(_0105_),
    .Q_N(_0997_),
    .Q(\bitserial_cipher.datapath.shifter2[2] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net201),
    .D(_0106_),
    .Q_N(_0996_),
    .Q(\bitserial_cipher.datapath.shifter2[30] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net202),
    .D(_0107_),
    .Q_N(_0995_),
    .Q(\bitserial_cipher.datapath.shifter2[31] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net203),
    .D(_0108_),
    .Q_N(_0994_),
    .Q(\bitserial_cipher.datapath.shifter2[32] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net204),
    .D(_0109_),
    .Q_N(_0993_),
    .Q(\bitserial_cipher.datapath.shifter2[33] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net205),
    .D(_0110_),
    .Q_N(_0992_),
    .Q(\bitserial_cipher.datapath.shifter2[34] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net206),
    .D(_0111_),
    .Q_N(_0991_),
    .Q(\bitserial_cipher.datapath.shifter2[35] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net207),
    .D(_0112_),
    .Q_N(_0990_),
    .Q(\bitserial_cipher.datapath.shifter2[36] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net208),
    .D(_0113_),
    .Q_N(_0989_),
    .Q(\bitserial_cipher.datapath.shifter2[37] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net209),
    .D(_0114_),
    .Q_N(_0988_),
    .Q(\bitserial_cipher.datapath.shifter2[38] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net210),
    .D(_0115_),
    .Q_N(_0987_),
    .Q(\bitserial_cipher.datapath.shifter2[39] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net211),
    .D(_0116_),
    .Q_N(_0986_),
    .Q(\bitserial_cipher.datapath.shifter2[3] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net212),
    .D(_0117_),
    .Q_N(_0985_),
    .Q(\bitserial_cipher.datapath.shifter2[40] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net213),
    .D(_0118_),
    .Q_N(_0984_),
    .Q(\bitserial_cipher.datapath.shifter2[41] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net214),
    .D(_0119_),
    .Q_N(_0983_),
    .Q(\bitserial_cipher.datapath.shifter2[42] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net215),
    .D(_0120_),
    .Q_N(_0982_),
    .Q(\bitserial_cipher.datapath.shifter2[43] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net216),
    .D(_0121_),
    .Q_N(_0981_),
    .Q(\bitserial_cipher.datapath.shifter2[44] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net217),
    .D(_0122_),
    .Q_N(_0980_),
    .Q(\bitserial_cipher.datapath.shifter2[45] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net218),
    .D(_0123_),
    .Q_N(_0979_),
    .Q(\bitserial_cipher.datapath.shifter2[46] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net219),
    .D(_0124_),
    .Q_N(_0978_),
    .Q(\bitserial_cipher.datapath.shifter2[47] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net220),
    .D(_0125_),
    .Q_N(_0977_),
    .Q(\bitserial_cipher.datapath.shifter2[48] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net221),
    .D(_0126_),
    .Q_N(_0976_),
    .Q(\bitserial_cipher.datapath.shifter2[49] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net222),
    .D(_0127_),
    .Q_N(_0975_),
    .Q(\bitserial_cipher.datapath.shifter2[4] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net223),
    .D(_0128_),
    .Q_N(_0974_),
    .Q(\bitserial_cipher.datapath.shifter2[50] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net224),
    .D(_0129_),
    .Q_N(_0973_),
    .Q(\bitserial_cipher.datapath.shifter2[51] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net225),
    .D(_0130_),
    .Q_N(_0972_),
    .Q(\bitserial_cipher.datapath.shifter2[52] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net226),
    .D(_0131_),
    .Q_N(_0971_),
    .Q(\bitserial_cipher.datapath.shifter2[53] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net227),
    .D(_0132_),
    .Q_N(_0970_),
    .Q(\bitserial_cipher.datapath.shifter2[54] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net228),
    .D(_0133_),
    .Q_N(_0969_),
    .Q(\bitserial_cipher.datapath.shifter2[55] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net229),
    .D(_0134_),
    .Q_N(_0968_),
    .Q(\bitserial_cipher.datapath.shifter2[56] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net230),
    .D(_0135_),
    .Q_N(_0967_),
    .Q(\bitserial_cipher.datapath.shifter2[57] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net231),
    .D(_0136_),
    .Q_N(_0966_),
    .Q(\bitserial_cipher.datapath.shifter2[58] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net232),
    .D(_0137_),
    .Q_N(_0965_),
    .Q(\bitserial_cipher.datapath.shifter2[59] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net233),
    .D(_0138_),
    .Q_N(_0964_),
    .Q(\bitserial_cipher.datapath.shifter2[5] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net234),
    .D(_0139_),
    .Q_N(_0963_),
    .Q(\bitserial_cipher.datapath.shifter2[60] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net235),
    .D(_0140_),
    .Q_N(_0962_),
    .Q(\bitserial_cipher.datapath.shifter2[61] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net236),
    .D(_0141_),
    .Q_N(_0961_),
    .Q(\bitserial_cipher.datapath.shifter2[62] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net237),
    .D(_0142_),
    .Q_N(_0960_),
    .Q(\bitserial_cipher.datapath.shifter2[63] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net238),
    .D(_0143_),
    .Q_N(_0959_),
    .Q(\bitserial_cipher.datapath.shifter2[6] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net239),
    .D(_0144_),
    .Q_N(_0958_),
    .Q(\bitserial_cipher.datapath.shifter2[7] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net240),
    .D(_0145_),
    .Q_N(_0957_),
    .Q(\bitserial_cipher.datapath.shifter2[8] ));
 sg13g2_dfrbp_1 \bitserial_cipher.datapath.shifter2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net241),
    .D(_0146_),
    .Q_N(_0956_),
    .Q(\bitserial_cipher.datapath.shifter2[9] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.fifo_ff0$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net242),
    .D(_0147_),
    .Q_N(_0955_),
    .Q(\bitserial_cipher.key_exp.fifo_ff0 ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.fifo_ff1$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net243),
    .D(_0148_),
    .Q_N(_0954_),
    .Q(\bitserial_cipher.key_exp.fifo_ff1 ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.fifo_ff2$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net244),
    .D(_0149_),
    .Q_N(_0953_),
    .Q(\bitserial_cipher.key_exp.fifo_ff2 ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.fifo_ff3$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net245),
    .D(_0150_),
    .Q_N(_0952_),
    .Q(\bitserial_cipher.key_exp.fifo_ff3 ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.lut_ff0$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net246),
    .D(_0151_),
    .Q_N(_0951_),
    .Q(\bitserial_cipher.key_exp.lut_ff0 ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.lut_ff1$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net247),
    .D(_0152_),
    .Q_N(_0950_),
    .Q(\bitserial_cipher.key_exp.lut_ff1 ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.lut_ff2$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net248),
    .D(_0153_),
    .Q_N(_0949_),
    .Q(\bitserial_cipher.key_exp.lut_ff2 ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.lut_ff3$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net249),
    .D(_0154_),
    .Q_N(_0948_),
    .Q(\bitserial_cipher.key_exp.lut_ff3 ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.round_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net250),
    .D(_0155_),
    .Q_N(_0000_),
    .Q(\bitserial_cipher.datapath.round_counter[0] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.round_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net251),
    .D(_0156_),
    .Q_N(_0002_),
    .Q(\bitserial_cipher.datapath.round_counter[1] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.round_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net252),
    .D(_0157_),
    .Q_N(_0001_),
    .Q(\bitserial_cipher.datapath.round_counter[2] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.round_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net253),
    .D(_0158_),
    .Q_N(_0947_),
    .Q(\bitserial_cipher.datapath.round_counter[3] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.round_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net254),
    .D(_0159_),
    .Q_N(_0946_),
    .Q(\bitserial_cipher.datapath.round_counter[4] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.round_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net255),
    .D(_0160_),
    .Q_N(_0945_),
    .Q(\bitserial_cipher.datapath.round_counter[5] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.round_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net256),
    .D(_0161_),
    .Q_N(_0003_),
    .Q(\bitserial_cipher.datapath.round_counter[6] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net257),
    .D(_0162_),
    .Q_N(_0944_),
    .Q(\bitserial_cipher.key_exp.shift_out1 ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net258),
    .D(_0163_),
    .Q_N(_0943_),
    .Q(\bitserial_cipher.key_exp.shifter1[10] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net259),
    .D(_0164_),
    .Q_N(_0942_),
    .Q(\bitserial_cipher.key_exp.shifter1[11] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net260),
    .D(_0165_),
    .Q_N(_0941_),
    .Q(\bitserial_cipher.key_exp.shifter1[12] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net261),
    .D(_0166_),
    .Q_N(_0940_),
    .Q(\bitserial_cipher.key_exp.shifter1[13] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net262),
    .D(_0167_),
    .Q_N(_0939_),
    .Q(\bitserial_cipher.key_exp.shifter1[14] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net263),
    .D(_0168_),
    .Q_N(_0938_),
    .Q(\bitserial_cipher.key_exp.shifter1[15] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net264),
    .D(_0169_),
    .Q_N(_0937_),
    .Q(\bitserial_cipher.key_exp.shifter1[16] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net265),
    .D(_0170_),
    .Q_N(_0936_),
    .Q(\bitserial_cipher.key_exp.shifter1[17] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net266),
    .D(_0171_),
    .Q_N(_0935_),
    .Q(\bitserial_cipher.key_exp.shifter1[18] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net267),
    .D(_0172_),
    .Q_N(_0934_),
    .Q(\bitserial_cipher.key_exp.shifter1[19] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net268),
    .D(_0173_),
    .Q_N(_0933_),
    .Q(\bitserial_cipher.key_exp.shifter1[1] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net269),
    .D(_0174_),
    .Q_N(_0932_),
    .Q(\bitserial_cipher.key_exp.shifter1[20] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net270),
    .D(_0175_),
    .Q_N(_0931_),
    .Q(\bitserial_cipher.key_exp.shifter1[21] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net271),
    .D(_0176_),
    .Q_N(_0930_),
    .Q(\bitserial_cipher.key_exp.shifter1[22] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net272),
    .D(_0177_),
    .Q_N(_0929_),
    .Q(\bitserial_cipher.key_exp.shifter1[23] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net273),
    .D(_0178_),
    .Q_N(_0928_),
    .Q(\bitserial_cipher.key_exp.shifter1[24] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net274),
    .D(_0179_),
    .Q_N(_0927_),
    .Q(\bitserial_cipher.key_exp.shifter1[25] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net275),
    .D(_0180_),
    .Q_N(_0926_),
    .Q(\bitserial_cipher.key_exp.shifter1[26] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net276),
    .D(_0181_),
    .Q_N(_0925_),
    .Q(\bitserial_cipher.key_exp.shifter1[27] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net277),
    .D(_0182_),
    .Q_N(_0924_),
    .Q(\bitserial_cipher.key_exp.shifter1[28] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net278),
    .D(_0183_),
    .Q_N(_0923_),
    .Q(\bitserial_cipher.key_exp.shifter1[29] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net279),
    .D(_0184_),
    .Q_N(_0922_),
    .Q(\bitserial_cipher.key_exp.shifter1[2] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net280),
    .D(_0185_),
    .Q_N(_0921_),
    .Q(\bitserial_cipher.key_exp.shifter1[30] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net281),
    .D(_0186_),
    .Q_N(_0920_),
    .Q(\bitserial_cipher.key_exp.shifter1[31] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net282),
    .D(_0187_),
    .Q_N(_0919_),
    .Q(\bitserial_cipher.key_exp.shifter1[32] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net283),
    .D(_0188_),
    .Q_N(_0918_),
    .Q(\bitserial_cipher.key_exp.shifter1[33] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net284),
    .D(_0189_),
    .Q_N(_0917_),
    .Q(\bitserial_cipher.key_exp.shifter1[34] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net285),
    .D(_0190_),
    .Q_N(_0916_),
    .Q(\bitserial_cipher.key_exp.shifter1[35] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net286),
    .D(_0191_),
    .Q_N(_0915_),
    .Q(\bitserial_cipher.key_exp.shifter1[36] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net287),
    .D(_0192_),
    .Q_N(_0914_),
    .Q(\bitserial_cipher.key_exp.shifter1[37] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net288),
    .D(_0193_),
    .Q_N(_0913_),
    .Q(\bitserial_cipher.key_exp.shifter1[38] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net289),
    .D(_0194_),
    .Q_N(_0912_),
    .Q(\bitserial_cipher.key_exp.shifter1[39] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net290),
    .D(_0195_),
    .Q_N(_0911_),
    .Q(\bitserial_cipher.key_exp.shifter1[3] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net291),
    .D(_0196_),
    .Q_N(_0910_),
    .Q(\bitserial_cipher.key_exp.shifter1[40] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net292),
    .D(_0197_),
    .Q_N(_0909_),
    .Q(\bitserial_cipher.key_exp.shifter1[41] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net293),
    .D(_0198_),
    .Q_N(_0908_),
    .Q(\bitserial_cipher.key_exp.shifter1[42] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net294),
    .D(_0199_),
    .Q_N(_0907_),
    .Q(\bitserial_cipher.key_exp.shifter1[43] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net295),
    .D(_0200_),
    .Q_N(_0906_),
    .Q(\bitserial_cipher.key_exp.shifter1[44] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net296),
    .D(_0201_),
    .Q_N(_0905_),
    .Q(\bitserial_cipher.key_exp.shifter1[45] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net297),
    .D(_0202_),
    .Q_N(_0904_),
    .Q(\bitserial_cipher.key_exp.shifter1[46] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net298),
    .D(_0203_),
    .Q_N(_0903_),
    .Q(\bitserial_cipher.key_exp.shifter1[47] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net299),
    .D(_0204_),
    .Q_N(_0902_),
    .Q(\bitserial_cipher.key_exp.shifter1[48] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net300),
    .D(_0205_),
    .Q_N(_0901_),
    .Q(\bitserial_cipher.key_exp.shifter1[49] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net301),
    .D(_0206_),
    .Q_N(_0900_),
    .Q(\bitserial_cipher.key_exp.shifter1[4] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net302),
    .D(_0207_),
    .Q_N(_0899_),
    .Q(\bitserial_cipher.key_exp.shifter1[50] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net303),
    .D(_0208_),
    .Q_N(_0898_),
    .Q(\bitserial_cipher.key_exp.shifter1[51] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net304),
    .D(_0209_),
    .Q_N(_0897_),
    .Q(\bitserial_cipher.key_exp.shifter1[52] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net305),
    .D(_0210_),
    .Q_N(_0896_),
    .Q(\bitserial_cipher.key_exp.shifter1[53] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net306),
    .D(_0211_),
    .Q_N(_0895_),
    .Q(\bitserial_cipher.key_exp.shifter1[54] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net307),
    .D(_0212_),
    .Q_N(_0894_),
    .Q(\bitserial_cipher.key_exp.shifter1[55] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net308),
    .D(_0213_),
    .Q_N(_0893_),
    .Q(\bitserial_cipher.key_exp.shifter1[56] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net309),
    .D(_0214_),
    .Q_N(_0892_),
    .Q(\bitserial_cipher.key_exp.shifter1[57] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net310),
    .D(_0215_),
    .Q_N(_0891_),
    .Q(\bitserial_cipher.key_exp.shifter1[58] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net311),
    .D(_0216_),
    .Q_N(_0890_),
    .Q(\bitserial_cipher.key_exp.shifter1[59] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net312),
    .D(_0217_),
    .Q_N(_0889_),
    .Q(\bitserial_cipher.key_exp.shifter1[5] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net313),
    .D(_0218_),
    .Q_N(_0888_),
    .Q(\bitserial_cipher.key_exp.shifter1[6] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net314),
    .D(_0219_),
    .Q_N(_0887_),
    .Q(\bitserial_cipher.key_exp.shifter1[7] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net315),
    .D(_0220_),
    .Q_N(_0886_),
    .Q(\bitserial_cipher.key_exp.shifter1[8] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net316),
    .D(_0221_),
    .Q_N(_0885_),
    .Q(\bitserial_cipher.key_exp.shifter1[9] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net317),
    .D(_0222_),
    .Q_N(_0884_),
    .Q(\bitserial_cipher.datapath.key_in ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net318),
    .D(_0223_),
    .Q_N(_0883_),
    .Q(\bitserial_cipher.key_exp.shifter2[10] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net319),
    .D(_0224_),
    .Q_N(_0882_),
    .Q(\bitserial_cipher.key_exp.shifter2[11] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net320),
    .D(_0225_),
    .Q_N(_0881_),
    .Q(\bitserial_cipher.key_exp.shifter2[12] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net321),
    .D(_0226_),
    .Q_N(_0880_),
    .Q(\bitserial_cipher.key_exp.shifter2[13] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net322),
    .D(_0227_),
    .Q_N(_0879_),
    .Q(\bitserial_cipher.key_exp.shifter2[14] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net323),
    .D(_0228_),
    .Q_N(_0878_),
    .Q(\bitserial_cipher.key_exp.shifter2[15] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net324),
    .D(_0229_),
    .Q_N(_0877_),
    .Q(\bitserial_cipher.key_exp.shifter2[16] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net325),
    .D(_0230_),
    .Q_N(_0876_),
    .Q(\bitserial_cipher.key_exp.shifter2[17] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net326),
    .D(_0231_),
    .Q_N(_0875_),
    .Q(\bitserial_cipher.key_exp.shifter2[18] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net327),
    .D(_0232_),
    .Q_N(_0874_),
    .Q(\bitserial_cipher.key_exp.shifter2[19] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net328),
    .D(_0233_),
    .Q_N(_0873_),
    .Q(\bitserial_cipher.key_exp.shifter2[1] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net329),
    .D(_0234_),
    .Q_N(_0872_),
    .Q(\bitserial_cipher.key_exp.shifter2[20] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net330),
    .D(_0235_),
    .Q_N(_0871_),
    .Q(\bitserial_cipher.key_exp.shifter2[21] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net331),
    .D(_0236_),
    .Q_N(_0870_),
    .Q(\bitserial_cipher.key_exp.shifter2[22] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net332),
    .D(_0237_),
    .Q_N(_0869_),
    .Q(\bitserial_cipher.key_exp.shifter2[23] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net333),
    .D(_0238_),
    .Q_N(_0868_),
    .Q(\bitserial_cipher.key_exp.shifter2[24] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net334),
    .D(_0239_),
    .Q_N(_0867_),
    .Q(\bitserial_cipher.key_exp.shifter2[25] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net335),
    .D(_0240_),
    .Q_N(_0866_),
    .Q(\bitserial_cipher.key_exp.shifter2[26] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net336),
    .D(_0241_),
    .Q_N(_0865_),
    .Q(\bitserial_cipher.key_exp.shifter2[27] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net337),
    .D(_0242_),
    .Q_N(_0864_),
    .Q(\bitserial_cipher.key_exp.shifter2[28] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net338),
    .D(_0243_),
    .Q_N(_0863_),
    .Q(\bitserial_cipher.key_exp.shifter2[29] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net339),
    .D(_0244_),
    .Q_N(_0862_),
    .Q(\bitserial_cipher.key_exp.shifter2[2] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net340),
    .D(_0245_),
    .Q_N(_0861_),
    .Q(\bitserial_cipher.key_exp.shifter2[30] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net341),
    .D(_0246_),
    .Q_N(_0860_),
    .Q(\bitserial_cipher.key_exp.shifter2[31] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net342),
    .D(_0247_),
    .Q_N(_0859_),
    .Q(\bitserial_cipher.key_exp.shifter2[32] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net343),
    .D(_0248_),
    .Q_N(_0858_),
    .Q(\bitserial_cipher.key_exp.shifter2[33] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net344),
    .D(_0249_),
    .Q_N(_0857_),
    .Q(\bitserial_cipher.key_exp.shifter2[34] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net345),
    .D(_0250_),
    .Q_N(_0856_),
    .Q(\bitserial_cipher.key_exp.shifter2[35] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net346),
    .D(_0251_),
    .Q_N(_0855_),
    .Q(\bitserial_cipher.key_exp.shifter2[36] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net347),
    .D(_0252_),
    .Q_N(_0854_),
    .Q(\bitserial_cipher.key_exp.shifter2[37] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net348),
    .D(_0253_),
    .Q_N(_0853_),
    .Q(\bitserial_cipher.key_exp.shifter2[38] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net349),
    .D(_0254_),
    .Q_N(_0852_),
    .Q(\bitserial_cipher.key_exp.shifter2[39] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net350),
    .D(_0255_),
    .Q_N(_0851_),
    .Q(\bitserial_cipher.key_exp.shifter2[3] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net351),
    .D(_0256_),
    .Q_N(_0850_),
    .Q(\bitserial_cipher.key_exp.shifter2[40] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net352),
    .D(_0257_),
    .Q_N(_0849_),
    .Q(\bitserial_cipher.key_exp.shifter2[41] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net353),
    .D(_0258_),
    .Q_N(_0848_),
    .Q(\bitserial_cipher.key_exp.shifter2[42] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net354),
    .D(_0259_),
    .Q_N(_0847_),
    .Q(\bitserial_cipher.key_exp.shifter2[43] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net355),
    .D(_0260_),
    .Q_N(_0846_),
    .Q(\bitserial_cipher.key_exp.shifter2[44] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net356),
    .D(_0261_),
    .Q_N(_0845_),
    .Q(\bitserial_cipher.key_exp.shifter2[45] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net357),
    .D(_0262_),
    .Q_N(_0844_),
    .Q(\bitserial_cipher.key_exp.shifter2[46] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net358),
    .D(_0263_),
    .Q_N(_0843_),
    .Q(\bitserial_cipher.key_exp.shifter2[47] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net359),
    .D(_0264_),
    .Q_N(_0842_),
    .Q(\bitserial_cipher.key_exp.shifter2[48] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net360),
    .D(_0265_),
    .Q_N(_0841_),
    .Q(\bitserial_cipher.key_exp.shifter2[49] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net361),
    .D(_0266_),
    .Q_N(_0840_),
    .Q(\bitserial_cipher.key_exp.shifter2[4] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net362),
    .D(_0267_),
    .Q_N(_0839_),
    .Q(\bitserial_cipher.key_exp.shifter2[50] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net363),
    .D(_0268_),
    .Q_N(_0838_),
    .Q(\bitserial_cipher.key_exp.shifter2[51] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net364),
    .D(_0269_),
    .Q_N(_0837_),
    .Q(\bitserial_cipher.key_exp.shifter2[52] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net365),
    .D(_0270_),
    .Q_N(_0836_),
    .Q(\bitserial_cipher.key_exp.shifter2[53] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net366),
    .D(_0271_),
    .Q_N(_0835_),
    .Q(\bitserial_cipher.key_exp.shifter2[54] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net367),
    .D(_0272_),
    .Q_N(_0834_),
    .Q(\bitserial_cipher.key_exp.shifter2[55] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net368),
    .D(_0273_),
    .Q_N(_0833_),
    .Q(\bitserial_cipher.key_exp.shifter2[56] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net369),
    .D(_0274_),
    .Q_N(_0832_),
    .Q(\bitserial_cipher.key_exp.shifter2[57] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net370),
    .D(_0275_),
    .Q_N(_0831_),
    .Q(\bitserial_cipher.key_exp.shifter2[58] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net371),
    .D(_0276_),
    .Q_N(_0830_),
    .Q(\bitserial_cipher.key_exp.shifter2[59] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net372),
    .D(_0277_),
    .Q_N(_0829_),
    .Q(\bitserial_cipher.key_exp.shifter2[5] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net373),
    .D(_0278_),
    .Q_N(_0828_),
    .Q(\bitserial_cipher.key_exp.shifter2[60] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net374),
    .D(_0279_),
    .Q_N(_0827_),
    .Q(\bitserial_cipher.key_exp.shifter2[61] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net375),
    .D(_0280_),
    .Q_N(_0826_),
    .Q(\bitserial_cipher.key_exp.shifter2[62] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net376),
    .D(_0281_),
    .Q_N(_0825_),
    .Q(\bitserial_cipher.key_exp.shifter2[63] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net377),
    .D(_0282_),
    .Q_N(_0824_),
    .Q(\bitserial_cipher.key_exp.shifter2[6] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net378),
    .D(_0283_),
    .Q_N(_0823_),
    .Q(\bitserial_cipher.key_exp.shifter2[7] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net379),
    .D(_0284_),
    .Q_N(_0822_),
    .Q(\bitserial_cipher.key_exp.shifter2[8] ));
 sg13g2_dfrbp_1 \bitserial_cipher.key_exp.shifter2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net380),
    .D(_0285_),
    .Q_N(_0821_),
    .Q(\bitserial_cipher.key_exp.shifter2[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout5 (.A(_0346_),
    .X(net5));
 sg13g2_buf_4 fanout6 (.X(net6),
    .A(_0491_));
 sg13g2_buf_4 fanout7 (.X(net7),
    .A(_0479_));
 sg13g2_buf_4 fanout8 (.X(net8),
    .A(_0467_));
 sg13g2_buf_4 fanout9 (.X(net9),
    .A(_0438_));
 sg13g2_buf_4 fanout10 (.X(net10),
    .A(_0426_));
 sg13g2_buf_1 fanout11 (.A(_0419_),
    .X(net11));
 sg13g2_buf_4 fanout12 (.X(net12),
    .A(_0414_));
 sg13g2_buf_1 fanout13 (.A(_0407_),
    .X(net13));
 sg13g2_buf_4 fanout14 (.X(net14),
    .A(_0402_));
 sg13g2_buf_1 fanout15 (.A(_0395_),
    .X(net15));
 sg13g2_buf_4 fanout16 (.X(net16),
    .A(_0390_));
 sg13g2_buf_1 fanout17 (.A(_0383_),
    .X(net17));
 sg13g2_buf_4 fanout18 (.X(net18),
    .A(_0378_));
 sg13g2_buf_2 fanout19 (.A(_0349_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0817_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0784_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0783_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0762_),
    .X(net23));
 sg13g2_buf_1 fanout24 (.A(_0750_),
    .X(net24));
 sg13g2_buf_1 fanout25 (.A(_0738_),
    .X(net25));
 sg13g2_buf_1 fanout26 (.A(_0726_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0714_),
    .X(net27));
 sg13g2_buf_4 fanout28 (.X(net28),
    .A(_0702_));
 sg13g2_buf_1 fanout29 (.A(_0701_),
    .X(net29));
 sg13g2_buf_4 fanout30 (.X(net30),
    .A(_0690_));
 sg13g2_buf_1 fanout31 (.A(_0689_),
    .X(net31));
 sg13g2_buf_4 fanout32 (.X(net32),
    .A(_0672_));
 sg13g2_buf_2 fanout33 (.A(_0671_),
    .X(net33));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(_0660_));
 sg13g2_buf_1 fanout35 (.A(_0659_),
    .X(net35));
 sg13g2_buf_4 fanout36 (.X(net36),
    .A(_0648_));
 sg13g2_buf_1 fanout37 (.A(_0647_),
    .X(net37));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(_0636_));
 sg13g2_buf_1 fanout39 (.A(_0635_),
    .X(net39));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(_0624_));
 sg13g2_buf_1 fanout41 (.A(_0623_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0612_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0601_),
    .X(net43));
 sg13g2_buf_4 fanout44 (.X(net44),
    .A(_0593_));
 sg13g2_buf_1 fanout45 (.A(_0591_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0558_),
    .X(net46));
 sg13g2_buf_1 fanout47 (.A(_0556_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0545_),
    .X(net48));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(_0527_));
 sg13g2_buf_2 fanout50 (.A(_0520_),
    .X(net50));
 sg13g2_buf_4 fanout51 (.X(net51),
    .A(_0515_));
 sg13g2_buf_1 fanout52 (.A(_0508_),
    .X(net52));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(_0503_));
 sg13g2_buf_1 fanout54 (.A(_0496_),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(_0484_),
    .X(net55));
 sg13g2_buf_1 fanout56 (.A(_0472_),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(_0460_),
    .X(net57));
 sg13g2_buf_1 fanout58 (.A(_0431_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0818_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0786_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0781_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0779_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0778_),
    .X(net63));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(_0751_));
 sg13g2_buf_4 fanout65 (.X(net65),
    .A(_0739_));
 sg13g2_buf_4 fanout66 (.X(net66),
    .A(_0727_));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(_0715_));
 sg13g2_buf_2 fanout68 (.A(_0713_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0578_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0559_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0557_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0555_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0547_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0544_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0554_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0543_),
    .X(net76));
 sg13g2_tielo _1918__77 (.L_LO(net77));
 sg13g2_tielo _1919__78 (.L_LO(net78));
 sg13g2_tielo _1920__79 (.L_LO(net79));
 sg13g2_tielo _1921__80 (.L_LO(net80));
 sg13g2_tielo _1922__81 (.L_LO(net81));
 sg13g2_tielo _1923__82 (.L_LO(net82));
 sg13g2_tielo _1924__83 (.L_LO(net83));
 sg13g2_tielo _1925__84 (.L_LO(net84));
 sg13g2_tielo _1926__85 (.L_LO(net85));
 sg13g2_tielo _1927__86 (.L_LO(net86));
 sg13g2_tielo _1928__87 (.L_LO(net87));
 sg13g2_tielo _1929__88 (.L_LO(net88));
 sg13g2_tielo _1930__89 (.L_LO(net89));
 sg13g2_tielo _1931__90 (.L_LO(net90));
 sg13g2_tielo _1932__91 (.L_LO(net91));
 sg13g2_tielo _1933__92 (.L_LO(net92));
 sg13g2_tielo _1934__93 (.L_LO(net93));
 sg13g2_tielo _1936__94 (.L_LO(net94));
 sg13g2_tielo _1937__95 (.L_LO(net95));
 sg13g2_tielo _1938__96 (.L_LO(net96));
 sg13g2_tielo _1939__97 (.L_LO(net97));
 sg13g2_tielo _1940__98 (.L_LO(net98));
 sg13g2_tielo _1941__99 (.L_LO(net99));
 sg13g2_tiehi \bitserial_cipher.datapath.bit_counter[1]$_SDFFE_PP0P__101  (.L_HI(net101));
 sg13g2_tiehi \bitserial_cipher.datapath.bit_counter[2]$_SDFFE_PP0P__102  (.L_HI(net102));
 sg13g2_tiehi \bitserial_cipher.datapath.bit_counter[3]$_SDFFE_PP0P__103  (.L_HI(net103));
 sg13g2_tiehi \bitserial_cipher.datapath.bit_counter[4]$_SDFFE_PP0P__104  (.L_HI(net104));
 sg13g2_tiehi \bitserial_cipher.datapath.bit_counter[5]$_SDFFE_PP0P__105  (.L_HI(net105));
 sg13g2_tiehi \bitserial_cipher.datapath.fifo_ff56$_SDFFE_PN0P__106  (.L_HI(net106));
 sg13g2_tiehi \bitserial_cipher.datapath.fifo_ff57$_SDFFE_PN0P__107  (.L_HI(net107));
 sg13g2_tiehi \bitserial_cipher.datapath.fifo_ff58$_SDFFE_PN0P__108  (.L_HI(net108));
 sg13g2_tiehi \bitserial_cipher.datapath.fifo_ff59$_SDFFE_PN0P__109  (.L_HI(net109));
 sg13g2_tiehi \bitserial_cipher.datapath.fifo_ff60$_SDFFE_PN0P__110  (.L_HI(net110));
 sg13g2_tiehi \bitserial_cipher.datapath.fifo_ff61$_SDFFE_PN0P__111  (.L_HI(net111));
 sg13g2_tiehi \bitserial_cipher.datapath.fifo_ff62$_SDFFE_PN0P__112  (.L_HI(net112));
 sg13g2_tiehi \bitserial_cipher.datapath.fifo_ff63$_SDFFE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \bitserial_cipher.datapath.lut_ff56$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_tiehi \bitserial_cipher.datapath.lut_ff57$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \bitserial_cipher.datapath.lut_ff58$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \bitserial_cipher.datapath.lut_ff59$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_tiehi \bitserial_cipher.datapath.lut_ff60$_SDFF_PN0__118  (.L_HI(net118));
 sg13g2_tiehi \bitserial_cipher.datapath.lut_ff61$_SDFF_PN0__119  (.L_HI(net119));
 sg13g2_tiehi \bitserial_cipher.datapath.lut_ff62$_SDFF_PN0__120  (.L_HI(net120));
 sg13g2_tiehi \bitserial_cipher.datapath.lut_ff63$_SDFF_PN0__121  (.L_HI(net121));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[0]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[10]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[11]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[12]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[13]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[14]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[15]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[16]$_SDFFE_PN0P__129  (.L_HI(net129));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[17]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[18]$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[19]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[1]$_SDFFE_PN0P__133  (.L_HI(net133));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[20]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[21]$_SDFFE_PN0P__135  (.L_HI(net135));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[22]$_SDFFE_PN0P__136  (.L_HI(net136));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[23]$_SDFFE_PN0P__137  (.L_HI(net137));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[24]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[25]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[26]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[27]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[28]$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[29]$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[2]$_SDFFE_PN0P__144  (.L_HI(net144));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[30]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[31]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[32]$_SDFFE_PN0P__147  (.L_HI(net147));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[33]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[34]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[35]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[36]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[37]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[38]$_SDFFE_PN0P__153  (.L_HI(net153));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[39]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[3]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[40]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[41]$_SDFFE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[42]$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[43]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[44]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[45]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[46]$_SDFFE_PN0P__162  (.L_HI(net162));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[47]$_SDFFE_PN0P__163  (.L_HI(net163));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[48]$_SDFFE_PN0P__164  (.L_HI(net164));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[49]$_SDFFE_PN0P__165  (.L_HI(net165));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[4]$_SDFFE_PN0P__166  (.L_HI(net166));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[50]$_SDFFE_PN0P__167  (.L_HI(net167));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[51]$_SDFFE_PN0P__168  (.L_HI(net168));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[52]$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[53]$_SDFFE_PN0P__170  (.L_HI(net170));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[54]$_SDFFE_PN0P__171  (.L_HI(net171));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[55]$_SDFFE_PN0P__172  (.L_HI(net172));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[5]$_SDFFE_PN0P__173  (.L_HI(net173));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[6]$_SDFFE_PN0P__174  (.L_HI(net174));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[7]$_SDFFE_PN0P__175  (.L_HI(net175));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[8]$_SDFFE_PN0P__176  (.L_HI(net176));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter1[9]$_SDFFE_PN0P__177  (.L_HI(net177));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[0]$_SDFFE_PN0P__178  (.L_HI(net178));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[10]$_SDFFE_PN0P__179  (.L_HI(net179));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[11]$_SDFFE_PN0P__180  (.L_HI(net180));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[12]$_SDFFE_PN0P__181  (.L_HI(net181));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[13]$_SDFFE_PN0P__182  (.L_HI(net182));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[14]$_SDFFE_PN0P__183  (.L_HI(net183));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[15]$_SDFFE_PN0P__184  (.L_HI(net184));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[16]$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[17]$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[18]$_SDFFE_PN0P__187  (.L_HI(net187));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[19]$_SDFFE_PN0P__188  (.L_HI(net188));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[1]$_SDFFE_PN0P__189  (.L_HI(net189));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[20]$_SDFFE_PN0P__190  (.L_HI(net190));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[21]$_SDFFE_PN0P__191  (.L_HI(net191));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[22]$_SDFFE_PN0P__192  (.L_HI(net192));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[23]$_SDFFE_PN0P__193  (.L_HI(net193));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[24]$_SDFFE_PN0P__194  (.L_HI(net194));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[25]$_SDFFE_PN0P__195  (.L_HI(net195));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[26]$_SDFFE_PN0P__196  (.L_HI(net196));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[27]$_SDFFE_PN0P__197  (.L_HI(net197));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[28]$_SDFFE_PN0P__198  (.L_HI(net198));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[29]$_SDFFE_PN0P__199  (.L_HI(net199));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[2]$_SDFFE_PN0P__200  (.L_HI(net200));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[30]$_SDFFE_PN0P__201  (.L_HI(net201));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[31]$_SDFFE_PN0P__202  (.L_HI(net202));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[32]$_SDFFE_PN0P__203  (.L_HI(net203));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[33]$_SDFFE_PN0P__204  (.L_HI(net204));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[34]$_SDFFE_PN0P__205  (.L_HI(net205));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[35]$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[36]$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[37]$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[38]$_SDFFE_PN0P__209  (.L_HI(net209));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[39]$_SDFFE_PN0P__210  (.L_HI(net210));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[3]$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[40]$_SDFFE_PN0P__212  (.L_HI(net212));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[41]$_SDFFE_PN0P__213  (.L_HI(net213));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[42]$_SDFFE_PN0P__214  (.L_HI(net214));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[43]$_SDFFE_PN0P__215  (.L_HI(net215));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[44]$_SDFFE_PN0P__216  (.L_HI(net216));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[45]$_SDFFE_PN0P__217  (.L_HI(net217));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[46]$_SDFFE_PN0P__218  (.L_HI(net218));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[47]$_SDFFE_PN0P__219  (.L_HI(net219));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[48]$_SDFFE_PN0P__220  (.L_HI(net220));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[49]$_SDFFE_PN0P__221  (.L_HI(net221));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[4]$_SDFFE_PN0P__222  (.L_HI(net222));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[50]$_SDFFE_PN0P__223  (.L_HI(net223));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[51]$_SDFFE_PN0P__224  (.L_HI(net224));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[52]$_SDFFE_PN0P__225  (.L_HI(net225));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[53]$_SDFFE_PN0P__226  (.L_HI(net226));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[54]$_SDFFE_PN0P__227  (.L_HI(net227));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[55]$_SDFFE_PN0P__228  (.L_HI(net228));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[56]$_SDFFE_PN0P__229  (.L_HI(net229));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[57]$_SDFFE_PN0P__230  (.L_HI(net230));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[58]$_SDFFE_PN0P__231  (.L_HI(net231));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[59]$_SDFFE_PN0P__232  (.L_HI(net232));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[5]$_SDFFE_PN0P__233  (.L_HI(net233));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[60]$_SDFFE_PN0P__234  (.L_HI(net234));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[61]$_SDFFE_PN0P__235  (.L_HI(net235));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[62]$_SDFFE_PN0P__236  (.L_HI(net236));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[63]$_SDFFE_PN0P__237  (.L_HI(net237));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[6]$_SDFFE_PN0P__238  (.L_HI(net238));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[7]$_SDFFE_PN0P__239  (.L_HI(net239));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[8]$_SDFFE_PN0P__240  (.L_HI(net240));
 sg13g2_tiehi \bitserial_cipher.datapath.shifter2[9]$_SDFFE_PN0P__241  (.L_HI(net241));
 sg13g2_tiehi \bitserial_cipher.key_exp.fifo_ff0$_SDFFE_PN0P__242  (.L_HI(net242));
 sg13g2_tiehi \bitserial_cipher.key_exp.fifo_ff1$_SDFFE_PN0P__243  (.L_HI(net243));
 sg13g2_tiehi \bitserial_cipher.key_exp.fifo_ff2$_SDFFE_PN0P__244  (.L_HI(net244));
 sg13g2_tiehi \bitserial_cipher.key_exp.fifo_ff3$_SDFFE_PN0P__245  (.L_HI(net245));
 sg13g2_tiehi \bitserial_cipher.key_exp.lut_ff0$_SDFFE_PN0P__246  (.L_HI(net246));
 sg13g2_tiehi \bitserial_cipher.key_exp.lut_ff1$_SDFFE_PN0P__247  (.L_HI(net247));
 sg13g2_tiehi \bitserial_cipher.key_exp.lut_ff2$_SDFFE_PN0P__248  (.L_HI(net248));
 sg13g2_tiehi \bitserial_cipher.key_exp.lut_ff3$_SDFFE_PN0P__249  (.L_HI(net249));
 sg13g2_tiehi \bitserial_cipher.key_exp.round_counter[0]$_SDFFE_PN0P__250  (.L_HI(net250));
 sg13g2_tiehi \bitserial_cipher.key_exp.round_counter[1]$_SDFFE_PN0P__251  (.L_HI(net251));
 sg13g2_tiehi \bitserial_cipher.key_exp.round_counter[2]$_SDFFE_PN0P__252  (.L_HI(net252));
 sg13g2_tiehi \bitserial_cipher.key_exp.round_counter[3]$_SDFFE_PN0P__253  (.L_HI(net253));
 sg13g2_tiehi \bitserial_cipher.key_exp.round_counter[4]$_SDFFE_PN0P__254  (.L_HI(net254));
 sg13g2_tiehi \bitserial_cipher.key_exp.round_counter[5]$_SDFFE_PN0P__255  (.L_HI(net255));
 sg13g2_tiehi \bitserial_cipher.key_exp.round_counter[6]$_SDFFE_PN0P__256  (.L_HI(net256));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[0]$_SDFFE_PN0P__257  (.L_HI(net257));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[10]$_SDFFE_PN0P__258  (.L_HI(net258));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[11]$_SDFFE_PN0P__259  (.L_HI(net259));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[12]$_SDFFE_PN0P__260  (.L_HI(net260));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[13]$_SDFFE_PN0P__261  (.L_HI(net261));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[14]$_SDFFE_PN0P__262  (.L_HI(net262));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[15]$_SDFFE_PN0P__263  (.L_HI(net263));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[16]$_SDFFE_PN0P__264  (.L_HI(net264));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[17]$_SDFFE_PN0P__265  (.L_HI(net265));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[18]$_SDFFE_PN0P__266  (.L_HI(net266));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[19]$_SDFFE_PN0P__267  (.L_HI(net267));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[1]$_SDFFE_PN0P__268  (.L_HI(net268));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[20]$_SDFFE_PN0P__269  (.L_HI(net269));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[21]$_SDFFE_PN0P__270  (.L_HI(net270));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[22]$_SDFFE_PN0P__271  (.L_HI(net271));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[23]$_SDFFE_PN0P__272  (.L_HI(net272));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[24]$_SDFFE_PN0P__273  (.L_HI(net273));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[25]$_SDFFE_PN0P__274  (.L_HI(net274));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[26]$_SDFFE_PN0P__275  (.L_HI(net275));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[27]$_SDFFE_PN0P__276  (.L_HI(net276));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[28]$_SDFFE_PN0P__277  (.L_HI(net277));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[29]$_SDFFE_PN0P__278  (.L_HI(net278));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[2]$_SDFFE_PN0P__279  (.L_HI(net279));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[30]$_SDFFE_PN0P__280  (.L_HI(net280));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[31]$_SDFFE_PN0P__281  (.L_HI(net281));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[32]$_SDFFE_PN0P__282  (.L_HI(net282));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[33]$_SDFFE_PN0P__283  (.L_HI(net283));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[34]$_SDFFE_PN0P__284  (.L_HI(net284));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[35]$_SDFFE_PN0P__285  (.L_HI(net285));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[36]$_SDFFE_PN0P__286  (.L_HI(net286));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[37]$_SDFFE_PN0P__287  (.L_HI(net287));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[38]$_SDFFE_PN0P__288  (.L_HI(net288));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[39]$_SDFFE_PN0P__289  (.L_HI(net289));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[3]$_SDFFE_PN0P__290  (.L_HI(net290));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[40]$_SDFFE_PN0P__291  (.L_HI(net291));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[41]$_SDFFE_PN0P__292  (.L_HI(net292));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[42]$_SDFFE_PN0P__293  (.L_HI(net293));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[43]$_SDFFE_PN0P__294  (.L_HI(net294));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[44]$_SDFFE_PN0P__295  (.L_HI(net295));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[45]$_SDFFE_PN0P__296  (.L_HI(net296));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[46]$_SDFFE_PN0P__297  (.L_HI(net297));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[47]$_SDFFE_PN0P__298  (.L_HI(net298));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[48]$_SDFFE_PN0P__299  (.L_HI(net299));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[49]$_SDFFE_PN0P__300  (.L_HI(net300));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[4]$_SDFFE_PN0P__301  (.L_HI(net301));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[50]$_SDFFE_PN0P__302  (.L_HI(net302));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[51]$_SDFFE_PN0P__303  (.L_HI(net303));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[52]$_SDFFE_PN0P__304  (.L_HI(net304));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[53]$_SDFFE_PN0P__305  (.L_HI(net305));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[54]$_SDFFE_PN0P__306  (.L_HI(net306));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[55]$_SDFFE_PN0P__307  (.L_HI(net307));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[56]$_SDFFE_PN0P__308  (.L_HI(net308));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[57]$_SDFFE_PN0P__309  (.L_HI(net309));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[58]$_SDFFE_PN0P__310  (.L_HI(net310));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[59]$_SDFFE_PN0P__311  (.L_HI(net311));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[5]$_SDFFE_PN0P__312  (.L_HI(net312));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[6]$_SDFFE_PN0P__313  (.L_HI(net313));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[7]$_SDFFE_PN0P__314  (.L_HI(net314));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[8]$_SDFFE_PN0P__315  (.L_HI(net315));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter1[9]$_SDFFE_PN0P__316  (.L_HI(net316));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[0]$_SDFFE_PN0P__317  (.L_HI(net317));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[10]$_SDFFE_PN0P__318  (.L_HI(net318));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[11]$_SDFFE_PN0P__319  (.L_HI(net319));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[12]$_SDFFE_PN0P__320  (.L_HI(net320));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[13]$_SDFFE_PN0P__321  (.L_HI(net321));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[14]$_SDFFE_PN0P__322  (.L_HI(net322));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[15]$_SDFFE_PN0P__323  (.L_HI(net323));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[16]$_SDFFE_PN0P__324  (.L_HI(net324));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[17]$_SDFFE_PN0P__325  (.L_HI(net325));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[18]$_SDFFE_PN0P__326  (.L_HI(net326));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[19]$_SDFFE_PN0P__327  (.L_HI(net327));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[1]$_SDFFE_PN0P__328  (.L_HI(net328));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[20]$_SDFFE_PN0P__329  (.L_HI(net329));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[21]$_SDFFE_PN0P__330  (.L_HI(net330));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[22]$_SDFFE_PN0P__331  (.L_HI(net331));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[23]$_SDFFE_PN0P__332  (.L_HI(net332));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[24]$_SDFFE_PN0P__333  (.L_HI(net333));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[25]$_SDFFE_PN0P__334  (.L_HI(net334));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[26]$_SDFFE_PN0P__335  (.L_HI(net335));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[27]$_SDFFE_PN0P__336  (.L_HI(net336));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[28]$_SDFFE_PN0P__337  (.L_HI(net337));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[29]$_SDFFE_PN0P__338  (.L_HI(net338));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[2]$_SDFFE_PN0P__339  (.L_HI(net339));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[30]$_SDFFE_PN0P__340  (.L_HI(net340));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[31]$_SDFFE_PN0P__341  (.L_HI(net341));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[32]$_SDFFE_PN0P__342  (.L_HI(net342));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[33]$_SDFFE_PN0P__343  (.L_HI(net343));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[34]$_SDFFE_PN0P__344  (.L_HI(net344));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[35]$_SDFFE_PN0P__345  (.L_HI(net345));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[36]$_SDFFE_PN0P__346  (.L_HI(net346));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[37]$_SDFFE_PN0P__347  (.L_HI(net347));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[38]$_SDFFE_PN0P__348  (.L_HI(net348));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[39]$_SDFFE_PN0P__349  (.L_HI(net349));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[3]$_SDFFE_PN0P__350  (.L_HI(net350));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[40]$_SDFFE_PN0P__351  (.L_HI(net351));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[41]$_SDFFE_PN0P__352  (.L_HI(net352));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[42]$_SDFFE_PN0P__353  (.L_HI(net353));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[43]$_SDFFE_PN0P__354  (.L_HI(net354));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[44]$_SDFFE_PN0P__355  (.L_HI(net355));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[45]$_SDFFE_PN0P__356  (.L_HI(net356));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[46]$_SDFFE_PN0P__357  (.L_HI(net357));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[47]$_SDFFE_PN0P__358  (.L_HI(net358));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[48]$_SDFFE_PN0P__359  (.L_HI(net359));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[49]$_SDFFE_PN0P__360  (.L_HI(net360));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[4]$_SDFFE_PN0P__361  (.L_HI(net361));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[50]$_SDFFE_PN0P__362  (.L_HI(net362));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[51]$_SDFFE_PN0P__363  (.L_HI(net363));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[52]$_SDFFE_PN0P__364  (.L_HI(net364));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[53]$_SDFFE_PN0P__365  (.L_HI(net365));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[54]$_SDFFE_PN0P__366  (.L_HI(net366));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[55]$_SDFFE_PN0P__367  (.L_HI(net367));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[56]$_SDFFE_PN0P__368  (.L_HI(net368));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[57]$_SDFFE_PN0P__369  (.L_HI(net369));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[58]$_SDFFE_PN0P__370  (.L_HI(net370));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[59]$_SDFFE_PN0P__371  (.L_HI(net371));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[5]$_SDFFE_PN0P__372  (.L_HI(net372));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[60]$_SDFFE_PN0P__373  (.L_HI(net373));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[61]$_SDFFE_PN0P__374  (.L_HI(net374));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[62]$_SDFFE_PN0P__375  (.L_HI(net375));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[63]$_SDFFE_PN0P__376  (.L_HI(net376));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[6]$_SDFFE_PN0P__377  (.L_HI(net377));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[7]$_SDFFE_PN0P__378  (.L_HI(net378));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[8]$_SDFFE_PN0P__379  (.L_HI(net379));
 sg13g2_tiehi \bitserial_cipher.key_exp.shifter2[9]$_SDFFE_PN0P__380  (.L_HI(net380));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_35_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_leaf_13_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_14_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_fill_2 FILLER_0_84 ();
 sg13g2_fill_2 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_150 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_decap_8 FILLER_0_171 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_fill_2 FILLER_0_206 ();
 sg13g2_decap_4 FILLER_0_234 ();
 sg13g2_fill_1 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_272 ();
 sg13g2_fill_1 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_fill_2 FILLER_0_313 ();
 sg13g2_fill_1 FILLER_0_315 ();
 sg13g2_fill_2 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_8 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_0_414 ();
 sg13g2_decap_8 FILLER_0_421 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_fill_2 FILLER_1_63 ();
 sg13g2_decap_4 FILLER_1_109 ();
 sg13g2_fill_2 FILLER_1_128 ();
 sg13g2_fill_1 FILLER_1_130 ();
 sg13g2_decap_4 FILLER_1_145 ();
 sg13g2_fill_2 FILLER_1_149 ();
 sg13g2_decap_8 FILLER_1_181 ();
 sg13g2_fill_2 FILLER_1_188 ();
 sg13g2_decap_8 FILLER_1_194 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_decap_4 FILLER_1_208 ();
 sg13g2_fill_2 FILLER_1_212 ();
 sg13g2_decap_4 FILLER_1_218 ();
 sg13g2_fill_1 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_4 FILLER_2_70 ();
 sg13g2_fill_1 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_79 ();
 sg13g2_fill_1 FILLER_2_86 ();
 sg13g2_decap_4 FILLER_2_92 ();
 sg13g2_fill_2 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_169 ();
 sg13g2_fill_2 FILLER_2_176 ();
 sg13g2_fill_2 FILLER_2_209 ();
 sg13g2_fill_2 FILLER_2_277 ();
 sg13g2_fill_2 FILLER_2_284 ();
 sg13g2_fill_1 FILLER_2_286 ();
 sg13g2_fill_1 FILLER_2_310 ();
 sg13g2_fill_1 FILLER_2_342 ();
 sg13g2_fill_2 FILLER_2_374 ();
 sg13g2_fill_1 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_4 FILLER_3_63 ();
 sg13g2_fill_1 FILLER_3_67 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_fill_1 FILLER_3_182 ();
 sg13g2_fill_1 FILLER_3_188 ();
 sg13g2_decap_4 FILLER_3_215 ();
 sg13g2_decap_4 FILLER_3_238 ();
 sg13g2_fill_2 FILLER_3_255 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_fill_1 FILLER_3_266 ();
 sg13g2_fill_1 FILLER_3_271 ();
 sg13g2_fill_1 FILLER_3_328 ();
 sg13g2_fill_2 FILLER_3_352 ();
 sg13g2_fill_1 FILLER_3_354 ();
 sg13g2_decap_4 FILLER_3_359 ();
 sg13g2_fill_1 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_63 ();
 sg13g2_fill_2 FILLER_4_100 ();
 sg13g2_fill_1 FILLER_4_102 ();
 sg13g2_fill_1 FILLER_4_149 ();
 sg13g2_fill_1 FILLER_4_193 ();
 sg13g2_fill_1 FILLER_4_198 ();
 sg13g2_decap_4 FILLER_4_203 ();
 sg13g2_fill_1 FILLER_4_207 ();
 sg13g2_fill_1 FILLER_4_234 ();
 sg13g2_fill_2 FILLER_4_281 ();
 sg13g2_fill_1 FILLER_4_283 ();
 sg13g2_fill_1 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_9 ();
 sg13g2_fill_2 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_62 ();
 sg13g2_decap_4 FILLER_5_69 ();
 sg13g2_fill_1 FILLER_5_99 ();
 sg13g2_fill_2 FILLER_5_110 ();
 sg13g2_fill_1 FILLER_5_122 ();
 sg13g2_fill_2 FILLER_5_149 ();
 sg13g2_fill_2 FILLER_5_177 ();
 sg13g2_fill_1 FILLER_5_215 ();
 sg13g2_decap_4 FILLER_5_220 ();
 sg13g2_fill_2 FILLER_5_224 ();
 sg13g2_fill_1 FILLER_5_251 ();
 sg13g2_fill_2 FILLER_5_267 ();
 sg13g2_fill_1 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_311 ();
 sg13g2_fill_1 FILLER_5_348 ();
 sg13g2_fill_2 FILLER_5_357 ();
 sg13g2_fill_1 FILLER_5_359 ();
 sg13g2_fill_2 FILLER_5_364 ();
 sg13g2_fill_1 FILLER_5_366 ();
 sg13g2_fill_1 FILLER_5_381 ();
 sg13g2_fill_1 FILLER_5_387 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_27 ();
 sg13g2_fill_1 FILLER_6_33 ();
 sg13g2_fill_1 FILLER_6_44 ();
 sg13g2_fill_1 FILLER_6_49 ();
 sg13g2_fill_1 FILLER_6_175 ();
 sg13g2_decap_4 FILLER_6_191 ();
 sg13g2_fill_2 FILLER_6_199 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_fill_2 FILLER_6_262 ();
 sg13g2_fill_2 FILLER_6_294 ();
 sg13g2_fill_2 FILLER_6_322 ();
 sg13g2_fill_1 FILLER_6_338 ();
 sg13g2_decap_4 FILLER_6_398 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_fill_1 FILLER_7_36 ();
 sg13g2_fill_2 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_54 ();
 sg13g2_fill_2 FILLER_7_65 ();
 sg13g2_fill_2 FILLER_7_71 ();
 sg13g2_fill_1 FILLER_7_83 ();
 sg13g2_fill_2 FILLER_7_115 ();
 sg13g2_fill_2 FILLER_7_143 ();
 sg13g2_fill_1 FILLER_7_145 ();
 sg13g2_fill_2 FILLER_7_155 ();
 sg13g2_fill_1 FILLER_7_157 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_fill_1 FILLER_7_224 ();
 sg13g2_fill_2 FILLER_7_244 ();
 sg13g2_fill_2 FILLER_7_285 ();
 sg13g2_fill_2 FILLER_7_297 ();
 sg13g2_fill_2 FILLER_7_309 ();
 sg13g2_fill_1 FILLER_7_316 ();
 sg13g2_fill_2 FILLER_7_387 ();
 sg13g2_fill_2 FILLER_7_399 ();
 sg13g2_fill_1 FILLER_7_401 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_82 ();
 sg13g2_fill_1 FILLER_8_103 ();
 sg13g2_fill_1 FILLER_8_112 ();
 sg13g2_fill_1 FILLER_8_123 ();
 sg13g2_fill_2 FILLER_8_128 ();
 sg13g2_fill_1 FILLER_8_135 ();
 sg13g2_fill_1 FILLER_8_140 ();
 sg13g2_fill_1 FILLER_8_276 ();
 sg13g2_fill_1 FILLER_8_307 ();
 sg13g2_fill_2 FILLER_8_326 ();
 sg13g2_fill_1 FILLER_8_351 ();
 sg13g2_fill_2 FILLER_8_367 ();
 sg13g2_fill_2 FILLER_8_405 ();
 sg13g2_fill_1 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_52 ();
 sg13g2_fill_2 FILLER_9_59 ();
 sg13g2_fill_1 FILLER_9_61 ();
 sg13g2_decap_8 FILLER_9_66 ();
 sg13g2_fill_2 FILLER_9_73 ();
 sg13g2_fill_1 FILLER_9_75 ();
 sg13g2_decap_4 FILLER_9_137 ();
 sg13g2_fill_2 FILLER_9_194 ();
 sg13g2_fill_2 FILLER_9_201 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_4 FILLER_9_214 ();
 sg13g2_fill_2 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_4 FILLER_9_424 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_11 ();
 sg13g2_fill_1 FILLER_10_86 ();
 sg13g2_fill_1 FILLER_10_111 ();
 sg13g2_fill_2 FILLER_10_116 ();
 sg13g2_decap_4 FILLER_10_132 ();
 sg13g2_fill_1 FILLER_10_243 ();
 sg13g2_fill_2 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_274 ();
 sg13g2_fill_1 FILLER_10_280 ();
 sg13g2_fill_2 FILLER_10_290 ();
 sg13g2_fill_1 FILLER_10_302 ();
 sg13g2_fill_2 FILLER_10_313 ();
 sg13g2_fill_1 FILLER_10_332 ();
 sg13g2_fill_2 FILLER_10_338 ();
 sg13g2_fill_1 FILLER_10_340 ();
 sg13g2_fill_1 FILLER_10_350 ();
 sg13g2_fill_1 FILLER_10_361 ();
 sg13g2_fill_1 FILLER_10_366 ();
 sg13g2_fill_1 FILLER_10_382 ();
 sg13g2_fill_1 FILLER_10_393 ();
 sg13g2_fill_1 FILLER_10_398 ();
 sg13g2_fill_1 FILLER_11_46 ();
 sg13g2_fill_1 FILLER_11_51 ();
 sg13g2_fill_1 FILLER_11_67 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_fill_1 FILLER_11_99 ();
 sg13g2_fill_1 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_153 ();
 sg13g2_fill_2 FILLER_11_206 ();
 sg13g2_decap_8 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_223 ();
 sg13g2_fill_2 FILLER_11_230 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_27 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_fill_2 FILLER_12_118 ();
 sg13g2_fill_1 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_130 ();
 sg13g2_fill_1 FILLER_12_140 ();
 sg13g2_fill_1 FILLER_12_297 ();
 sg13g2_fill_2 FILLER_12_317 ();
 sg13g2_fill_1 FILLER_12_319 ();
 sg13g2_fill_2 FILLER_12_365 ();
 sg13g2_fill_2 FILLER_12_372 ();
 sg13g2_fill_1 FILLER_12_374 ();
 sg13g2_fill_2 FILLER_12_383 ();
 sg13g2_fill_1 FILLER_12_385 ();
 sg13g2_fill_2 FILLER_12_391 ();
 sg13g2_fill_1 FILLER_12_393 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_140 ();
 sg13g2_fill_2 FILLER_13_154 ();
 sg13g2_fill_1 FILLER_13_210 ();
 sg13g2_fill_1 FILLER_13_215 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_fill_1 FILLER_13_230 ();
 sg13g2_decap_4 FILLER_13_241 ();
 sg13g2_fill_2 FILLER_13_245 ();
 sg13g2_fill_1 FILLER_13_252 ();
 sg13g2_fill_1 FILLER_13_279 ();
 sg13g2_fill_1 FILLER_13_306 ();
 sg13g2_fill_2 FILLER_13_338 ();
 sg13g2_fill_2 FILLER_13_345 ();
 sg13g2_fill_2 FILLER_13_357 ();
 sg13g2_fill_1 FILLER_13_385 ();
 sg13g2_fill_1 FILLER_13_390 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_422 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_fill_2 FILLER_14_65 ();
 sg13g2_decap_8 FILLER_14_71 ();
 sg13g2_fill_2 FILLER_14_78 ();
 sg13g2_fill_1 FILLER_14_175 ();
 sg13g2_fill_1 FILLER_14_181 ();
 sg13g2_fill_1 FILLER_14_208 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_242 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_291 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_decap_4 FILLER_14_361 ();
 sg13g2_fill_2 FILLER_14_365 ();
 sg13g2_fill_2 FILLER_14_371 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_111 ();
 sg13g2_fill_1 FILLER_15_144 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_fill_1 FILLER_15_184 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_decap_4 FILLER_15_201 ();
 sg13g2_fill_2 FILLER_15_219 ();
 sg13g2_fill_1 FILLER_15_262 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_fill_1 FILLER_15_283 ();
 sg13g2_fill_1 FILLER_15_315 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_fill_1 FILLER_15_348 ();
 sg13g2_fill_2 FILLER_15_375 ();
 sg13g2_fill_1 FILLER_15_381 ();
 sg13g2_fill_2 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_53 ();
 sg13g2_fill_2 FILLER_16_64 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_decap_4 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_144 ();
 sg13g2_fill_2 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_210 ();
 sg13g2_decap_4 FILLER_16_248 ();
 sg13g2_fill_1 FILLER_16_278 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_299 ();
 sg13g2_fill_2 FILLER_16_304 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_fill_2 FILLER_17_31 ();
 sg13g2_fill_2 FILLER_17_59 ();
 sg13g2_fill_1 FILLER_17_61 ();
 sg13g2_fill_1 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_247 ();
 sg13g2_fill_1 FILLER_17_341 ();
 sg13g2_fill_1 FILLER_17_352 ();
 sg13g2_fill_1 FILLER_17_361 ();
 sg13g2_fill_2 FILLER_17_381 ();
 sg13g2_fill_1 FILLER_17_403 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_15 ();
 sg13g2_fill_1 FILLER_18_116 ();
 sg13g2_fill_2 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_fill_2 FILLER_18_212 ();
 sg13g2_fill_2 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_fill_1 FILLER_18_391 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_fill_1 FILLER_19_45 ();
 sg13g2_fill_2 FILLER_19_50 ();
 sg13g2_fill_2 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_decap_4 FILLER_19_100 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_fill_2 FILLER_19_184 ();
 sg13g2_fill_2 FILLER_19_190 ();
 sg13g2_decap_4 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_272 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_299 ();
 sg13g2_fill_2 FILLER_19_304 ();
 sg13g2_fill_2 FILLER_19_310 ();
 sg13g2_decap_4 FILLER_19_341 ();
 sg13g2_fill_1 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_4 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_decap_4 FILLER_19_377 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_fill_1 FILLER_19_387 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_15 ();
 sg13g2_decap_4 FILLER_20_114 ();
 sg13g2_fill_2 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_151 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_decap_4 FILLER_20_205 ();
 sg13g2_fill_1 FILLER_20_209 ();
 sg13g2_decap_4 FILLER_20_214 ();
 sg13g2_decap_4 FILLER_20_257 ();
 sg13g2_decap_4 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_fill_2 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_361 ();
 sg13g2_fill_2 FILLER_20_393 ();
 sg13g2_decap_4 FILLER_20_400 ();
 sg13g2_fill_1 FILLER_20_404 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_decap_4 FILLER_20_425 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_2 FILLER_21_52 ();
 sg13g2_fill_2 FILLER_21_58 ();
 sg13g2_fill_2 FILLER_21_64 ();
 sg13g2_fill_2 FILLER_21_71 ();
 sg13g2_fill_1 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_decap_4 FILLER_21_116 ();
 sg13g2_fill_1 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_decap_4 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_198 ();
 sg13g2_fill_2 FILLER_21_204 ();
 sg13g2_fill_1 FILLER_21_206 ();
 sg13g2_decap_4 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_decap_4 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_226 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_fill_2 FILLER_21_282 ();
 sg13g2_fill_1 FILLER_21_284 ();
 sg13g2_fill_2 FILLER_21_293 ();
 sg13g2_decap_4 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_fill_1 FILLER_21_369 ();
 sg13g2_fill_2 FILLER_21_402 ();
 sg13g2_fill_1 FILLER_22_77 ();
 sg13g2_fill_2 FILLER_22_82 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_decap_4 FILLER_22_107 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_decap_4 FILLER_22_148 ();
 sg13g2_decap_8 FILLER_22_156 ();
 sg13g2_fill_1 FILLER_22_163 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_fill_1 FILLER_22_183 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_268 ();
 sg13g2_fill_2 FILLER_22_310 ();
 sg13g2_decap_4 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_fill_2 FILLER_22_326 ();
 sg13g2_fill_1 FILLER_22_328 ();
 sg13g2_fill_1 FILLER_22_333 ();
 sg13g2_fill_2 FILLER_22_360 ();
 sg13g2_fill_2 FILLER_22_393 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_27 ();
 sg13g2_fill_1 FILLER_23_62 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_fill_2 FILLER_23_151 ();
 sg13g2_fill_2 FILLER_23_184 ();
 sg13g2_fill_1 FILLER_23_186 ();
 sg13g2_decap_4 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_208 ();
 sg13g2_decap_4 FILLER_23_221 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_1 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_fill_2 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_304 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_fill_2 FILLER_23_397 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_36 ();
 sg13g2_decap_4 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_125 ();
 sg13g2_fill_2 FILLER_24_173 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_230 ();
 sg13g2_decap_4 FILLER_24_282 ();
 sg13g2_decap_4 FILLER_24_290 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_fill_2 FILLER_24_410 ();
 sg13g2_decap_4 FILLER_24_425 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_fill_2 FILLER_25_55 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_decap_4 FILLER_25_62 ();
 sg13g2_decap_4 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_146 ();
 sg13g2_fill_1 FILLER_25_152 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_fill_1 FILLER_25_173 ();
 sg13g2_fill_1 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_fill_2 FILLER_25_216 ();
 sg13g2_fill_2 FILLER_25_253 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_fill_2 FILLER_25_344 ();
 sg13g2_fill_2 FILLER_25_351 ();
 sg13g2_fill_2 FILLER_25_379 ();
 sg13g2_fill_2 FILLER_25_391 ();
 sg13g2_fill_1 FILLER_25_393 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_41 ();
 sg13g2_fill_2 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_fill_2 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_4 FILLER_26_192 ();
 sg13g2_fill_2 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_fill_1 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_236 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_257 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_2 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_298 ();
 sg13g2_fill_2 FILLER_26_305 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_27 ();
 sg13g2_fill_1 FILLER_27_59 ();
 sg13g2_fill_1 FILLER_27_64 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_97 ();
 sg13g2_fill_2 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_273 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_decap_4 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_fill_1 FILLER_27_364 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_fill_1 FILLER_27_383 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_146 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_decap_4 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_fill_2 FILLER_28_171 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_fill_2 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_393 ();
 sg13g2_fill_1 FILLER_28_398 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_decap_4 FILLER_29_242 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_333 ();
 sg13g2_fill_1 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_356 ();
 sg13g2_fill_2 FILLER_29_377 ();
 sg13g2_fill_1 FILLER_29_379 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_1 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_31 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_68 ();
 sg13g2_fill_1 FILLER_30_74 ();
 sg13g2_fill_2 FILLER_30_79 ();
 sg13g2_fill_1 FILLER_30_86 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_decap_4 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_148 ();
 sg13g2_decap_4 FILLER_30_158 ();
 sg13g2_fill_2 FILLER_30_162 ();
 sg13g2_fill_2 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_184 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_232 ();
 sg13g2_fill_1 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_272 ();
 sg13g2_fill_1 FILLER_30_283 ();
 sg13g2_fill_1 FILLER_30_291 ();
 sg13g2_fill_2 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_395 ();
 sg13g2_fill_1 FILLER_30_397 ();
 sg13g2_fill_1 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_105 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_fill_2 FILLER_31_112 ();
 sg13g2_fill_1 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_129 ();
 sg13g2_decap_4 FILLER_31_175 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_fill_1 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_247 ();
 sg13g2_decap_4 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_302 ();
 sg13g2_fill_1 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_fill_1 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_380 ();
 sg13g2_fill_2 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_fill_1 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_decap_4 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_216 ();
 sg13g2_fill_1 FILLER_32_227 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_fill_2 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_303 ();
 sg13g2_decap_4 FILLER_32_335 ();
 sg13g2_fill_2 FILLER_32_375 ();
 sg13g2_fill_1 FILLER_32_381 ();
 sg13g2_fill_2 FILLER_32_386 ();
 sg13g2_fill_2 FILLER_33_26 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_59 ();
 sg13g2_fill_2 FILLER_33_102 ();
 sg13g2_fill_1 FILLER_33_104 ();
 sg13g2_fill_1 FILLER_33_143 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_204 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_2 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_1 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_44 ();
 sg13g2_fill_1 FILLER_34_89 ();
 sg13g2_fill_1 FILLER_34_126 ();
 sg13g2_fill_2 FILLER_34_157 ();
 sg13g2_decap_4 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_168 ();
 sg13g2_decap_4 FILLER_34_174 ();
 sg13g2_fill_2 FILLER_34_189 ();
 sg13g2_fill_1 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_210 ();
 sg13g2_fill_1 FILLER_34_219 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_242 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_2 FILLER_34_269 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_decap_4 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_303 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_368 ();
 sg13g2_fill_2 FILLER_34_378 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_fill_1 FILLER_34_401 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_fill_2 FILLER_35_81 ();
 sg13g2_fill_2 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_138 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_fill_1 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_277 ();
 sg13g2_fill_2 FILLER_35_301 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_31 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_fill_2 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_180 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_204 ();
 sg13g2_fill_2 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_309 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_1 FILLER_37_31 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_1 FILLER_37_204 ();
 sg13g2_fill_1 FILLER_37_283 ();
 sg13g2_fill_2 FILLER_37_310 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_fill_2 FILLER_37_369 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_fill_2 FILLER_38_79 ();
 sg13g2_fill_2 FILLER_38_104 ();
 sg13g2_fill_1 FILLER_38_106 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_166 ();
 sg13g2_decap_4 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_263 ();
 sg13g2_fill_2 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_351 ();
 sg13g2_fill_1 FILLER_38_358 ();
 sg13g2_fill_1 FILLER_38_369 ();
 sg13g2_fill_2 FILLER_38_380 ();
 sg13g2_fill_2 FILLER_38_402 ();
endmodule
