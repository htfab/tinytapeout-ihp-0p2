VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA tt_um_ccattuto_conway_via1_2_2200_440_1_5_410_410
  VIARULE via1Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal1 Via1 Metal2 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.01 0.125 0.05 0.005 ;
  ROWCOL 1 5 ;
END tt_um_ccattuto_conway_via1_2_2200_440_1_5_410_410

VIA tt_um_ccattuto_conway_via2_3_2200_440_1_5_410_410
  VIARULE via2Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal2 Via2 Metal3 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 1 5 ;
END tt_um_ccattuto_conway_via2_3_2200_440_1_5_410_410

VIA tt_um_ccattuto_conway_via3_4_2200_440_1_5_410_410
  VIARULE via3Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.005 0.05 0.05 0.005 ;
  ROWCOL 1 5 ;
END tt_um_ccattuto_conway_via3_4_2200_440_1_5_410_410

VIA tt_um_ccattuto_conway_via4_5_2200_440_1_5_410_410
  VIARULE via4Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal4 Via4 Metal5 ;
  CUTSPACING 0.22 0.22 ;
  ENCLOSURE 0.05 0.005 0.185 0.05 ;
  ROWCOL 1 5 ;
END tt_um_ccattuto_conway_via4_5_2200_440_1_5_410_410

MACRO tt_um_ccattuto_conway
  FOREIGN tt_um_ccattuto_conway 0 0 ;
  CLASS BLOCK ;
  SIZE 642.24 BY 313.74 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  198.57 312.74 198.87 313.74 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  202.41 312.74 202.71 313.74 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  194.73 312.74 195.03 313.74 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  190.89 312.74 191.19 313.74 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  187.05 312.74 187.35 313.74 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  183.21 312.74 183.51 313.74 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  179.37 312.74 179.67 313.74 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  175.53 312.74 175.83 313.74 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  171.69 312.74 171.99 313.74 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  167.85 312.74 168.15 313.74 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  164.01 312.74 164.31 313.74 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  160.17 312.74 160.47 313.74 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  156.33 312.74 156.63 313.74 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  152.49 312.74 152.79 313.74 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  148.65 312.74 148.95 313.74 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  144.81 312.74 145.11 313.74 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  140.97 312.74 141.27 313.74 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  137.13 312.74 137.43 313.74 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  133.29 312.74 133.59 313.74 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  68.01 312.74 68.31 313.74 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  64.17 312.74 64.47 313.74 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  60.33 312.74 60.63 313.74 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  56.49 312.74 56.79 313.74 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  52.65 312.74 52.95 313.74 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  48.81 312.74 49.11 313.74 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  44.97 312.74 45.27 313.74 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  41.13 312.74 41.43 313.74 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  98.73 312.74 99.03 313.74 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  94.89 312.74 95.19 313.74 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  91.05 312.74 91.35 313.74 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  87.21 312.74 87.51 313.74 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  83.37 312.74 83.67 313.74 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  79.53 312.74 79.83 313.74 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  75.69 312.74 75.99 313.74 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  71.85 312.74 72.15 313.74 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  129.45 312.74 129.75 313.74 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  125.61 312.74 125.91 313.74 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  121.77 312.74 122.07 313.74 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  117.93 312.74 118.23 313.74 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  114.09 312.74 114.39 313.74 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  110.25 312.74 110.55 313.74 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  106.41 312.74 106.71 313.74 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT  102.57 312.74 102.87 313.74 ;
    END
  END uo_out[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT  620.18 3.56 622.38 310.18 ;
        RECT  544.58 3.56 546.78 310.18 ;
        RECT  468.98 3.56 471.18 310.18 ;
        RECT  393.38 3.56 395.58 310.18 ;
        RECT  317.78 3.56 319.98 310.18 ;
        RECT  242.18 3.56 244.38 310.18 ;
        RECT  166.58 3.56 168.78 310.18 ;
        RECT  90.98 3.56 93.18 310.18 ;
        RECT  15.38 3.56 17.58 310.18 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT  582.38 3.56 584.58 310.18 ;
        RECT  506.78 3.56 508.98 310.18 ;
        RECT  431.18 3.56 433.38 310.18 ;
        RECT  355.58 3.56 357.78 310.18 ;
        RECT  279.98 3.56 282.18 310.18 ;
        RECT  204.38 3.56 206.58 310.18 ;
        RECT  128.78 3.56 130.98 310.18 ;
        RECT  53.18 3.56 55.38 310.18 ;
    END
  END VPWR
  OBS
    LAYER Metal1 ;
     RECT  1.775 3.56 639.36 313.74 ;
    LAYER Metal2 ;
     RECT  1.775 3.56 639.36 313.74 ;
    LAYER Metal3 ;
     RECT  1.775 3.56 639.36 313.74 ;
    LAYER Metal4 ;
     RECT  1.775 3.56 639.36 313.74 ;
    LAYER Metal5 ;
     RECT  1.775 3.56 639.36 313.74 ;
  END
END tt_um_ccattuto_conway
END LIBRARY
