module tt_um_MichaelBell_tinyQV (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire clknet_leaf_0_clk;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire net1396;
 wire \addr[0] ;
 wire \addr[10] ;
 wire \addr[11] ;
 wire \addr[12] ;
 wire \addr[13] ;
 wire \addr[14] ;
 wire \addr[15] ;
 wire \addr[16] ;
 wire \addr[17] ;
 wire \addr[18] ;
 wire \addr[19] ;
 wire \addr[1] ;
 wire \addr[20] ;
 wire \addr[21] ;
 wire \addr[22] ;
 wire \addr[23] ;
 wire \addr[24] ;
 wire \addr[25] ;
 wire \addr[26] ;
 wire \addr[27] ;
 wire \addr[2] ;
 wire \addr[3] ;
 wire \addr[4] ;
 wire \addr[5] ;
 wire \addr[6] ;
 wire \addr[7] ;
 wire \addr[8] ;
 wire \addr[9] ;
 wire \data_to_write[0] ;
 wire \data_to_write[10] ;
 wire \data_to_write[11] ;
 wire \data_to_write[12] ;
 wire \data_to_write[13] ;
 wire \data_to_write[14] ;
 wire \data_to_write[15] ;
 wire \data_to_write[16] ;
 wire \data_to_write[17] ;
 wire \data_to_write[18] ;
 wire \data_to_write[19] ;
 wire \data_to_write[1] ;
 wire \data_to_write[20] ;
 wire \data_to_write[21] ;
 wire \data_to_write[22] ;
 wire \data_to_write[23] ;
 wire \data_to_write[24] ;
 wire \data_to_write[25] ;
 wire \data_to_write[26] ;
 wire \data_to_write[27] ;
 wire \data_to_write[28] ;
 wire \data_to_write[29] ;
 wire \data_to_write[2] ;
 wire \data_to_write[30] ;
 wire \data_to_write[31] ;
 wire \data_to_write[3] ;
 wire \data_to_write[4] ;
 wire \data_to_write[5] ;
 wire \data_to_write[6] ;
 wire \data_to_write[7] ;
 wire \data_to_write[8] ;
 wire \data_to_write[9] ;
 wire debug_data_continue;
 wire debug_instr_valid;
 wire \debug_rd[0] ;
 wire \debug_rd[1] ;
 wire \debug_rd[2] ;
 wire \debug_rd[3] ;
 wire \debug_rd_r[0] ;
 wire \debug_rd_r[1] ;
 wire \debug_rd_r[2] ;
 wire \debug_rd_r[3] ;
 wire debug_register_data;
 wire debug_uart_txd;
 wire \gpio_out[0] ;
 wire \gpio_out[1] ;
 wire \gpio_out[2] ;
 wire \gpio_out[3] ;
 wire \gpio_out[4] ;
 wire \gpio_out[5] ;
 wire \gpio_out[6] ;
 wire \gpio_out[7] ;
 wire \gpio_out_sel[0] ;
 wire \gpio_out_sel[1] ;
 wire \gpio_out_sel[2] ;
 wire \gpio_out_sel[3] ;
 wire \gpio_out_sel[4] ;
 wire \gpio_out_sel[5] ;
 wire \gpio_out_sel[6] ;
 wire \gpio_out_sel[7] ;
 wire \gpio_out_sel[8] ;
 wire \gpio_out_sel[9] ;
 wire \i_debug_uart_tx.cycle_counter[0] ;
 wire \i_debug_uart_tx.cycle_counter[1] ;
 wire \i_debug_uart_tx.cycle_counter[2] ;
 wire \i_debug_uart_tx.cycle_counter[3] ;
 wire \i_debug_uart_tx.cycle_counter[4] ;
 wire \i_debug_uart_tx.data_to_send[0] ;
 wire \i_debug_uart_tx.data_to_send[1] ;
 wire \i_debug_uart_tx.data_to_send[2] ;
 wire \i_debug_uart_tx.data_to_send[3] ;
 wire \i_debug_uart_tx.data_to_send[4] ;
 wire \i_debug_uart_tx.data_to_send[5] ;
 wire \i_debug_uart_tx.data_to_send[6] ;
 wire \i_debug_uart_tx.data_to_send[7] ;
 wire \i_debug_uart_tx.fsm_state[0] ;
 wire \i_debug_uart_tx.fsm_state[1] ;
 wire \i_debug_uart_tx.fsm_state[2] ;
 wire \i_debug_uart_tx.fsm_state[3] ;
 wire \i_debug_uart_tx.resetn ;
 wire \i_pwm.pwm_count[0] ;
 wire \i_pwm.pwm_count[1] ;
 wire \i_pwm.pwm_count[2] ;
 wire \i_pwm.pwm_count[3] ;
 wire \i_pwm.pwm_count[4] ;
 wire \i_pwm.pwm_count[5] ;
 wire \i_pwm.pwm_count[6] ;
 wire \i_pwm.pwm_count[7] ;
 wire \i_pwm.pwm_level[0] ;
 wire \i_pwm.pwm_level[1] ;
 wire \i_pwm.pwm_level[2] ;
 wire \i_pwm.pwm_level[3] ;
 wire \i_pwm.pwm_level[4] ;
 wire \i_pwm.pwm_level[5] ;
 wire \i_pwm.pwm_level[6] ;
 wire \i_pwm.pwm_level[7] ;
 wire \i_spi.bits_remaining[0] ;
 wire \i_spi.bits_remaining[1] ;
 wire \i_spi.bits_remaining[2] ;
 wire \i_spi.bits_remaining[3] ;
 wire \i_spi.busy ;
 wire \i_spi.clock_count[0] ;
 wire \i_spi.clock_count[1] ;
 wire \i_spi.clock_divider[0] ;
 wire \i_spi.clock_divider[1] ;
 wire \i_spi.data[0] ;
 wire \i_spi.data[1] ;
 wire \i_spi.data[2] ;
 wire \i_spi.data[3] ;
 wire \i_spi.data[4] ;
 wire \i_spi.data[5] ;
 wire \i_spi.data[6] ;
 wire \i_spi.data[7] ;
 wire \i_spi.end_txn_reg ;
 wire \i_spi.read_latency ;
 wire \i_spi.spi_clk_out ;
 wire \i_spi.spi_dc ;
 wire \i_spi.spi_select ;
 wire \i_tinyqv.cpu.additional_mem_ops[0] ;
 wire \i_tinyqv.cpu.additional_mem_ops[1] ;
 wire \i_tinyqv.cpu.additional_mem_ops[2] ;
 wire \i_tinyqv.cpu.alu_op[0] ;
 wire \i_tinyqv.cpu.alu_op[1] ;
 wire \i_tinyqv.cpu.alu_op[2] ;
 wire \i_tinyqv.cpu.alu_op[3] ;
 wire \i_tinyqv.cpu.counter[2] ;
 wire \i_tinyqv.cpu.counter[3] ;
 wire \i_tinyqv.cpu.counter[4] ;
 wire \i_tinyqv.cpu.data_read_n[0] ;
 wire \i_tinyqv.cpu.data_read_n[1] ;
 wire \i_tinyqv.cpu.data_ready_core ;
 wire \i_tinyqv.cpu.data_ready_latch ;
 wire \i_tinyqv.cpu.data_write_n[0] ;
 wire \i_tinyqv.cpu.data_write_n[1] ;
 wire \i_tinyqv.cpu.i_core.cmp ;
 wire \i_tinyqv.cpu.i_core.cmp_out ;
 wire \i_tinyqv.cpu.i_core.cy ;
 wire \i_tinyqv.cpu.i_core.cy_out ;
 wire \i_tinyqv.cpu.i_core.cycle[0] ;
 wire \i_tinyqv.cpu.i_core.cycle[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[0] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[2] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[3] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[4] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[5] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[6] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.cy ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.rstn ;
 wire \i_tinyqv.cpu.i_core.i_instrret.add ;
 wire \i_tinyqv.cpu.i_core.i_instrret.cy ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[0] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[1] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[2] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[3] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[10] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[11] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[12] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[13] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[14] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[15] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[16] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[17] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[18] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[19] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[20] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[21] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[22] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[23] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[24] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[25] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[26] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[27] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[28] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[29] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[30] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[31] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[4] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[5] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[6] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[7] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[8] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[9] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[0] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[10] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[11] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[1] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[2] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[3] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[5] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[6] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[7] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[8] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[9] ;
 wire \i_tinyqv.cpu.i_core.interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.is_double_fault_r ;
 wire \i_tinyqv.cpu.i_core.is_interrupt ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.load_done ;
 wire \i_tinyqv.cpu.i_core.load_top_bit ;
 wire \i_tinyqv.cpu.i_core.mcause[0] ;
 wire \i_tinyqv.cpu.i_core.mcause[1] ;
 wire \i_tinyqv.cpu.i_core.mcause[3] ;
 wire \i_tinyqv.cpu.i_core.mcause[4] ;
 wire \i_tinyqv.cpu.i_core.mem_op[0] ;
 wire \i_tinyqv.cpu.i_core.mem_op[1] ;
 wire \i_tinyqv.cpu.i_core.mem_op[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[0] ;
 wire \i_tinyqv.cpu.i_core.mepc[10] ;
 wire \i_tinyqv.cpu.i_core.mepc[11] ;
 wire \i_tinyqv.cpu.i_core.mepc[12] ;
 wire \i_tinyqv.cpu.i_core.mepc[13] ;
 wire \i_tinyqv.cpu.i_core.mepc[14] ;
 wire \i_tinyqv.cpu.i_core.mepc[15] ;
 wire \i_tinyqv.cpu.i_core.mepc[16] ;
 wire \i_tinyqv.cpu.i_core.mepc[17] ;
 wire \i_tinyqv.cpu.i_core.mepc[18] ;
 wire \i_tinyqv.cpu.i_core.mepc[19] ;
 wire \i_tinyqv.cpu.i_core.mepc[1] ;
 wire \i_tinyqv.cpu.i_core.mepc[20] ;
 wire \i_tinyqv.cpu.i_core.mepc[21] ;
 wire \i_tinyqv.cpu.i_core.mepc[22] ;
 wire \i_tinyqv.cpu.i_core.mepc[23] ;
 wire \i_tinyqv.cpu.i_core.mepc[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[3] ;
 wire \i_tinyqv.cpu.i_core.mepc[4] ;
 wire \i_tinyqv.cpu.i_core.mepc[5] ;
 wire \i_tinyqv.cpu.i_core.mepc[6] ;
 wire \i_tinyqv.cpu.i_core.mepc[7] ;
 wire \i_tinyqv.cpu.i_core.mepc[8] ;
 wire \i_tinyqv.cpu.i_core.mepc[9] ;
 wire \i_tinyqv.cpu.i_core.mie[16] ;
 wire \i_tinyqv.cpu.i_core.mie[17] ;
 wire \i_tinyqv.cpu.i_core.mie[18] ;
 wire \i_tinyqv.cpu.i_core.mie[19] ;
 wire \i_tinyqv.cpu.i_core.mip[16] ;
 wire \i_tinyqv.cpu.i_core.mip[17] ;
 wire \i_tinyqv.cpu.i_core.mstatus_mie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mpie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mte ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[0] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[10] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[11] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[12] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[13] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[14] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[15] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[1] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[2] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[3] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[4] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[5] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[6] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[7] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[8] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[9] ;
 wire \i_tinyqv.cpu.i_core.time_hi[0] ;
 wire \i_tinyqv.cpu.i_core.time_hi[1] ;
 wire \i_tinyqv.cpu.i_core.time_hi[2] ;
 wire \i_tinyqv.cpu.imm[12] ;
 wire \i_tinyqv.cpu.imm[13] ;
 wire \i_tinyqv.cpu.imm[14] ;
 wire \i_tinyqv.cpu.imm[15] ;
 wire \i_tinyqv.cpu.imm[16] ;
 wire \i_tinyqv.cpu.imm[17] ;
 wire \i_tinyqv.cpu.imm[18] ;
 wire \i_tinyqv.cpu.imm[19] ;
 wire \i_tinyqv.cpu.imm[20] ;
 wire \i_tinyqv.cpu.imm[21] ;
 wire \i_tinyqv.cpu.imm[22] ;
 wire \i_tinyqv.cpu.imm[23] ;
 wire \i_tinyqv.cpu.imm[24] ;
 wire \i_tinyqv.cpu.imm[25] ;
 wire \i_tinyqv.cpu.imm[26] ;
 wire \i_tinyqv.cpu.imm[27] ;
 wire \i_tinyqv.cpu.imm[28] ;
 wire \i_tinyqv.cpu.imm[29] ;
 wire \i_tinyqv.cpu.imm[30] ;
 wire \i_tinyqv.cpu.imm[31] ;
 wire \i_tinyqv.cpu.instr_data[0][0] ;
 wire \i_tinyqv.cpu.instr_data[0][10] ;
 wire \i_tinyqv.cpu.instr_data[0][11] ;
 wire \i_tinyqv.cpu.instr_data[0][12] ;
 wire \i_tinyqv.cpu.instr_data[0][13] ;
 wire \i_tinyqv.cpu.instr_data[0][14] ;
 wire \i_tinyqv.cpu.instr_data[0][15] ;
 wire \i_tinyqv.cpu.instr_data[0][1] ;
 wire \i_tinyqv.cpu.instr_data[0][2] ;
 wire \i_tinyqv.cpu.instr_data[0][3] ;
 wire \i_tinyqv.cpu.instr_data[0][4] ;
 wire \i_tinyqv.cpu.instr_data[0][5] ;
 wire \i_tinyqv.cpu.instr_data[0][6] ;
 wire \i_tinyqv.cpu.instr_data[0][7] ;
 wire \i_tinyqv.cpu.instr_data[0][8] ;
 wire \i_tinyqv.cpu.instr_data[0][9] ;
 wire \i_tinyqv.cpu.instr_data[1][0] ;
 wire \i_tinyqv.cpu.instr_data[1][10] ;
 wire \i_tinyqv.cpu.instr_data[1][11] ;
 wire \i_tinyqv.cpu.instr_data[1][12] ;
 wire \i_tinyqv.cpu.instr_data[1][13] ;
 wire \i_tinyqv.cpu.instr_data[1][14] ;
 wire \i_tinyqv.cpu.instr_data[1][15] ;
 wire \i_tinyqv.cpu.instr_data[1][1] ;
 wire \i_tinyqv.cpu.instr_data[1][2] ;
 wire \i_tinyqv.cpu.instr_data[1][3] ;
 wire \i_tinyqv.cpu.instr_data[1][4] ;
 wire \i_tinyqv.cpu.instr_data[1][5] ;
 wire \i_tinyqv.cpu.instr_data[1][6] ;
 wire \i_tinyqv.cpu.instr_data[1][7] ;
 wire \i_tinyqv.cpu.instr_data[1][8] ;
 wire \i_tinyqv.cpu.instr_data[1][9] ;
 wire \i_tinyqv.cpu.instr_data[2][0] ;
 wire \i_tinyqv.cpu.instr_data[2][10] ;
 wire \i_tinyqv.cpu.instr_data[2][11] ;
 wire \i_tinyqv.cpu.instr_data[2][12] ;
 wire \i_tinyqv.cpu.instr_data[2][13] ;
 wire \i_tinyqv.cpu.instr_data[2][14] ;
 wire \i_tinyqv.cpu.instr_data[2][15] ;
 wire \i_tinyqv.cpu.instr_data[2][1] ;
 wire \i_tinyqv.cpu.instr_data[2][2] ;
 wire \i_tinyqv.cpu.instr_data[2][3] ;
 wire \i_tinyqv.cpu.instr_data[2][4] ;
 wire \i_tinyqv.cpu.instr_data[2][5] ;
 wire \i_tinyqv.cpu.instr_data[2][6] ;
 wire \i_tinyqv.cpu.instr_data[2][7] ;
 wire \i_tinyqv.cpu.instr_data[2][8] ;
 wire \i_tinyqv.cpu.instr_data[2][9] ;
 wire \i_tinyqv.cpu.instr_data[3][0] ;
 wire \i_tinyqv.cpu.instr_data[3][10] ;
 wire \i_tinyqv.cpu.instr_data[3][11] ;
 wire \i_tinyqv.cpu.instr_data[3][12] ;
 wire \i_tinyqv.cpu.instr_data[3][13] ;
 wire \i_tinyqv.cpu.instr_data[3][14] ;
 wire \i_tinyqv.cpu.instr_data[3][15] ;
 wire \i_tinyqv.cpu.instr_data[3][1] ;
 wire \i_tinyqv.cpu.instr_data[3][2] ;
 wire \i_tinyqv.cpu.instr_data[3][3] ;
 wire \i_tinyqv.cpu.instr_data[3][4] ;
 wire \i_tinyqv.cpu.instr_data[3][5] ;
 wire \i_tinyqv.cpu.instr_data[3][6] ;
 wire \i_tinyqv.cpu.instr_data[3][7] ;
 wire \i_tinyqv.cpu.instr_data[3][8] ;
 wire \i_tinyqv.cpu.instr_data[3][9] ;
 wire \i_tinyqv.cpu.instr_data_in[0] ;
 wire \i_tinyqv.cpu.instr_data_in[10] ;
 wire \i_tinyqv.cpu.instr_data_in[11] ;
 wire \i_tinyqv.cpu.instr_data_in[12] ;
 wire \i_tinyqv.cpu.instr_data_in[13] ;
 wire \i_tinyqv.cpu.instr_data_in[14] ;
 wire \i_tinyqv.cpu.instr_data_in[15] ;
 wire \i_tinyqv.cpu.instr_data_in[1] ;
 wire \i_tinyqv.cpu.instr_data_in[2] ;
 wire \i_tinyqv.cpu.instr_data_in[3] ;
 wire \i_tinyqv.cpu.instr_data_in[4] ;
 wire \i_tinyqv.cpu.instr_data_in[5] ;
 wire \i_tinyqv.cpu.instr_data_in[6] ;
 wire \i_tinyqv.cpu.instr_data_in[7] ;
 wire \i_tinyqv.cpu.instr_data_in[8] ;
 wire \i_tinyqv.cpu.instr_data_in[9] ;
 wire \i_tinyqv.cpu.instr_data_start[10] ;
 wire \i_tinyqv.cpu.instr_data_start[11] ;
 wire \i_tinyqv.cpu.instr_data_start[12] ;
 wire \i_tinyqv.cpu.instr_data_start[13] ;
 wire \i_tinyqv.cpu.instr_data_start[14] ;
 wire \i_tinyqv.cpu.instr_data_start[15] ;
 wire \i_tinyqv.cpu.instr_data_start[16] ;
 wire \i_tinyqv.cpu.instr_data_start[17] ;
 wire \i_tinyqv.cpu.instr_data_start[18] ;
 wire \i_tinyqv.cpu.instr_data_start[19] ;
 wire \i_tinyqv.cpu.instr_data_start[20] ;
 wire \i_tinyqv.cpu.instr_data_start[21] ;
 wire \i_tinyqv.cpu.instr_data_start[22] ;
 wire \i_tinyqv.cpu.instr_data_start[23] ;
 wire \i_tinyqv.cpu.instr_data_start[3] ;
 wire \i_tinyqv.cpu.instr_data_start[4] ;
 wire \i_tinyqv.cpu.instr_data_start[5] ;
 wire \i_tinyqv.cpu.instr_data_start[6] ;
 wire \i_tinyqv.cpu.instr_data_start[7] ;
 wire \i_tinyqv.cpu.instr_data_start[8] ;
 wire \i_tinyqv.cpu.instr_data_start[9] ;
 wire \i_tinyqv.cpu.instr_fetch_running ;
 wire \i_tinyqv.cpu.instr_fetch_started ;
 wire \i_tinyqv.cpu.instr_fetch_stopped ;
 wire \i_tinyqv.cpu.instr_len[1] ;
 wire \i_tinyqv.cpu.instr_len[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[1] ;
 wire \i_tinyqv.cpu.instr_write_offset[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[3] ;
 wire \i_tinyqv.cpu.is_alu_imm ;
 wire \i_tinyqv.cpu.is_alu_reg ;
 wire \i_tinyqv.cpu.is_auipc ;
 wire \i_tinyqv.cpu.is_branch ;
 wire \i_tinyqv.cpu.is_jal ;
 wire \i_tinyqv.cpu.is_jalr ;
 wire \i_tinyqv.cpu.is_load ;
 wire \i_tinyqv.cpu.is_lui ;
 wire \i_tinyqv.cpu.is_store ;
 wire \i_tinyqv.cpu.is_system ;
 wire \i_tinyqv.cpu.load_started ;
 wire \i_tinyqv.cpu.mem_op_increment_reg ;
 wire \i_tinyqv.cpu.no_write_in_progress ;
 wire \i_tinyqv.cpu.pc[1] ;
 wire \i_tinyqv.cpu.pc[2] ;
 wire \i_tinyqv.cpu.was_early_branch ;
 wire \i_tinyqv.mem.data_from_read[16] ;
 wire \i_tinyqv.mem.data_from_read[17] ;
 wire \i_tinyqv.mem.data_from_read[18] ;
 wire \i_tinyqv.mem.data_from_read[19] ;
 wire \i_tinyqv.mem.data_from_read[20] ;
 wire \i_tinyqv.mem.data_from_read[21] ;
 wire \i_tinyqv.mem.data_from_read[22] ;
 wire \i_tinyqv.mem.data_from_read[23] ;
 wire \i_tinyqv.mem.data_stall ;
 wire \i_tinyqv.mem.instr_active ;
 wire \i_tinyqv.mem.q_ctrl.addr[0] ;
 wire \i_tinyqv.mem.q_ctrl.addr[10] ;
 wire \i_tinyqv.mem.q_ctrl.addr[11] ;
 wire \i_tinyqv.mem.q_ctrl.addr[12] ;
 wire \i_tinyqv.mem.q_ctrl.addr[13] ;
 wire \i_tinyqv.mem.q_ctrl.addr[14] ;
 wire \i_tinyqv.mem.q_ctrl.addr[15] ;
 wire \i_tinyqv.mem.q_ctrl.addr[16] ;
 wire \i_tinyqv.mem.q_ctrl.addr[17] ;
 wire \i_tinyqv.mem.q_ctrl.addr[18] ;
 wire \i_tinyqv.mem.q_ctrl.addr[19] ;
 wire \i_tinyqv.mem.q_ctrl.addr[1] ;
 wire \i_tinyqv.mem.q_ctrl.addr[20] ;
 wire \i_tinyqv.mem.q_ctrl.addr[21] ;
 wire \i_tinyqv.mem.q_ctrl.addr[22] ;
 wire \i_tinyqv.mem.q_ctrl.addr[23] ;
 wire \i_tinyqv.mem.q_ctrl.addr[2] ;
 wire \i_tinyqv.mem.q_ctrl.addr[3] ;
 wire \i_tinyqv.mem.q_ctrl.addr[4] ;
 wire \i_tinyqv.mem.q_ctrl.addr[5] ;
 wire \i_tinyqv.mem.q_ctrl.addr[6] ;
 wire \i_tinyqv.mem.q_ctrl.addr[7] ;
 wire \i_tinyqv.mem.q_ctrl.addr[8] ;
 wire \i_tinyqv.mem.q_ctrl.addr[9] ;
 wire \i_tinyqv.mem.q_ctrl.data_ready ;
 wire \i_tinyqv.mem.q_ctrl.data_req ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[0] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[1] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[2] ;
 wire \i_tinyqv.mem.q_ctrl.is_writing ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_a_sel ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_b_sel ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[0] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[1] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[2] ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_out ;
 wire \i_tinyqv.mem.q_ctrl.spi_data_oe[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_flash_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_a_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_b_select ;
 wire \i_tinyqv.mem.q_ctrl.stop_txn_reg ;
 wire \i_tinyqv.mem.qspi_data_buf[10] ;
 wire \i_tinyqv.mem.qspi_data_buf[11] ;
 wire \i_tinyqv.mem.qspi_data_buf[12] ;
 wire \i_tinyqv.mem.qspi_data_buf[13] ;
 wire \i_tinyqv.mem.qspi_data_buf[14] ;
 wire \i_tinyqv.mem.qspi_data_buf[15] ;
 wire \i_tinyqv.mem.qspi_data_buf[24] ;
 wire \i_tinyqv.mem.qspi_data_buf[25] ;
 wire \i_tinyqv.mem.qspi_data_buf[26] ;
 wire \i_tinyqv.mem.qspi_data_buf[27] ;
 wire \i_tinyqv.mem.qspi_data_buf[28] ;
 wire \i_tinyqv.mem.qspi_data_buf[29] ;
 wire \i_tinyqv.mem.qspi_data_buf[30] ;
 wire \i_tinyqv.mem.qspi_data_buf[31] ;
 wire \i_tinyqv.mem.qspi_data_buf[8] ;
 wire \i_tinyqv.mem.qspi_data_buf[9] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[0] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[1] ;
 wire \i_tinyqv.mem.qspi_write_done ;
 wire \i_uart_rx.bit_sample ;
 wire \i_uart_rx.cycle_counter[0] ;
 wire \i_uart_rx.cycle_counter[10] ;
 wire \i_uart_rx.cycle_counter[1] ;
 wire \i_uart_rx.cycle_counter[2] ;
 wire \i_uart_rx.cycle_counter[3] ;
 wire \i_uart_rx.cycle_counter[4] ;
 wire \i_uart_rx.cycle_counter[5] ;
 wire \i_uart_rx.cycle_counter[6] ;
 wire \i_uart_rx.cycle_counter[7] ;
 wire \i_uart_rx.cycle_counter[8] ;
 wire \i_uart_rx.cycle_counter[9] ;
 wire \i_uart_rx.fsm_state[0] ;
 wire \i_uart_rx.fsm_state[1] ;
 wire \i_uart_rx.fsm_state[2] ;
 wire \i_uart_rx.fsm_state[3] ;
 wire \i_uart_rx.recieved_data[0] ;
 wire \i_uart_rx.recieved_data[1] ;
 wire \i_uart_rx.recieved_data[2] ;
 wire \i_uart_rx.recieved_data[3] ;
 wire \i_uart_rx.recieved_data[4] ;
 wire \i_uart_rx.recieved_data[5] ;
 wire \i_uart_rx.recieved_data[6] ;
 wire \i_uart_rx.recieved_data[7] ;
 wire \i_uart_rx.rxd_reg[0] ;
 wire \i_uart_rx.rxd_reg[1] ;
 wire \i_uart_rx.uart_rts ;
 wire \i_uart_tx.cycle_counter[0] ;
 wire \i_uart_tx.cycle_counter[10] ;
 wire \i_uart_tx.cycle_counter[1] ;
 wire \i_uart_tx.cycle_counter[2] ;
 wire \i_uart_tx.cycle_counter[3] ;
 wire \i_uart_tx.cycle_counter[4] ;
 wire \i_uart_tx.cycle_counter[5] ;
 wire \i_uart_tx.cycle_counter[6] ;
 wire \i_uart_tx.cycle_counter[7] ;
 wire \i_uart_tx.cycle_counter[8] ;
 wire \i_uart_tx.cycle_counter[9] ;
 wire \i_uart_tx.data_to_send[0] ;
 wire \i_uart_tx.data_to_send[1] ;
 wire \i_uart_tx.data_to_send[2] ;
 wire \i_uart_tx.data_to_send[3] ;
 wire \i_uart_tx.data_to_send[4] ;
 wire \i_uart_tx.data_to_send[5] ;
 wire \i_uart_tx.data_to_send[6] ;
 wire \i_uart_tx.data_to_send[7] ;
 wire \i_uart_tx.fsm_state[0] ;
 wire \i_uart_tx.fsm_state[1] ;
 wire \i_uart_tx.fsm_state[2] ;
 wire \i_uart_tx.fsm_state[3] ;
 wire \i_uart_tx.txd_reg ;
 wire uio_out7;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_8 _06226_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .X(_00766_));
 sg13g2_buf_1 _06227_ (.A(net339),
    .X(_00767_));
 sg13g2_buf_8 _06228_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .X(_00768_));
 sg13g2_buf_8 _06229_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .X(_00769_));
 sg13g2_and2_1 _06230_ (.A(_00768_),
    .B(net338),
    .X(_00770_));
 sg13g2_nor2b_1 _06231_ (.A(net293),
    .B_N(_00770_),
    .Y(_00771_));
 sg13g2_buf_8 _06232_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .X(_00772_));
 sg13g2_buf_8 _06233_ (.A(_00772_),
    .X(_00773_));
 sg13g2_mux2_1 _06234_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .S(net292),
    .X(_00774_));
 sg13g2_buf_8 _06235_ (.A(net338),
    .X(_00775_));
 sg13g2_nand2b_1 _06236_ (.Y(_00776_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .A_N(net291));
 sg13g2_nand3_1 _06237_ (.B(net291),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .A(net293),
    .Y(_00777_));
 sg13g2_o21ai_1 _06238_ (.B1(_00777_),
    .Y(_00778_),
    .A1(net293),
    .A2(_00776_));
 sg13g2_buf_8 _06239_ (.A(net292),
    .X(_00779_));
 sg13g2_buf_8 _06240_ (.A(_00768_),
    .X(_00780_));
 sg13g2_inv_1 _06241_ (.Y(_00781_),
    .A(_00780_));
 sg13g2_nor2_1 _06242_ (.A(net242),
    .B(_00781_),
    .Y(_00782_));
 sg13g2_buf_1 _06243_ (.A(net339),
    .X(_00783_));
 sg13g2_mux2_1 _06244_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .S(net292),
    .X(_00784_));
 sg13g2_nor2b_1 _06245_ (.A(net338),
    .B_N(_00768_),
    .Y(_00785_));
 sg13g2_and3_1 _06246_ (.X(_00786_),
    .A(_00783_),
    .B(_00784_),
    .C(_00785_));
 sg13g2_a221oi_1 _06247_ (.B2(_00782_),
    .C1(_00786_),
    .B1(_00778_),
    .A1(_00771_),
    .Y(_00787_),
    .A2(_00774_));
 sg13g2_inv_1 _06248_ (.Y(_00788_),
    .A(net292));
 sg13g2_buf_8 _06249_ (.A(\i_tinyqv.cpu.counter[2] ),
    .X(_00789_));
 sg13g2_buf_8 _06250_ (.A(_00789_),
    .X(_00790_));
 sg13g2_buf_8 _06251_ (.A(\i_tinyqv.cpu.counter[3] ),
    .X(_00791_));
 sg13g2_buf_2 _06252_ (.A(\i_tinyqv.cpu.counter[4] ),
    .X(_00792_));
 sg13g2_nand3b_1 _06253_ (.B(net337),
    .C(net336),
    .Y(_00793_),
    .A_N(net288));
 sg13g2_buf_2 _06254_ (.A(_00793_),
    .X(_00794_));
 sg13g2_nand2_1 _06255_ (.Y(_00795_),
    .A(net293),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ));
 sg13g2_o21ai_1 _06256_ (.B1(_00795_),
    .Y(_00796_),
    .A1(net289),
    .A2(_00794_));
 sg13g2_nor2b_1 _06257_ (.A(_00768_),
    .B_N(net338),
    .Y(_00797_));
 sg13g2_nand3_1 _06258_ (.B(_00796_),
    .C(_00797_),
    .A(_00788_),
    .Y(_00798_));
 sg13g2_nand2_1 _06259_ (.Y(_00799_),
    .A(_00787_),
    .B(_00798_));
 sg13g2_nand2b_1 _06260_ (.Y(_00800_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .A_N(net291));
 sg13g2_buf_1 _06261_ (.A(net338),
    .X(_00801_));
 sg13g2_nand3_1 _06262_ (.B(net287),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .A(net293),
    .Y(_00802_));
 sg13g2_o21ai_1 _06263_ (.B1(_00802_),
    .Y(_00803_),
    .A1(net289),
    .A2(_00800_));
 sg13g2_buf_1 _06264_ (.A(_00768_),
    .X(_00804_));
 sg13g2_nand2b_1 _06265_ (.Y(_00805_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .A_N(net286));
 sg13g2_nand3b_1 _06266_ (.B(net286),
    .C(net293),
    .Y(_00806_),
    .A_N(_00092_));
 sg13g2_o21ai_1 _06267_ (.B1(_00806_),
    .Y(_00807_),
    .A1(net289),
    .A2(_00805_));
 sg13g2_a22oi_1 _06268_ (.Y(_00808_),
    .B1(_00807_),
    .B2(net287),
    .A2(_00803_),
    .A1(_00781_));
 sg13g2_nor2b_1 _06269_ (.A(_00772_),
    .B_N(net339),
    .Y(_00809_));
 sg13g2_buf_2 _06270_ (.A(_00809_),
    .X(_00810_));
 sg13g2_nand3_1 _06271_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .C(_00810_),
    .A(_00781_),
    .Y(_00811_));
 sg13g2_nor2b_1 _06272_ (.A(net339),
    .B_N(_00772_),
    .Y(_00812_));
 sg13g2_buf_2 _06273_ (.A(_00812_),
    .X(_00813_));
 sg13g2_nand3_1 _06274_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .C(_00813_),
    .A(net286),
    .Y(_00814_));
 sg13g2_a21o_1 _06275_ (.A2(_00814_),
    .A1(_00811_),
    .B1(net287),
    .X(_00815_));
 sg13g2_o21ai_1 _06276_ (.B1(_00815_),
    .Y(_00816_),
    .A1(_00788_),
    .A2(_00808_));
 sg13g2_buf_2 _06277_ (.A(\i_tinyqv.cpu.alu_op[1] ),
    .X(_00817_));
 sg13g2_buf_1 _06278_ (.A(\i_tinyqv.cpu.alu_op[2] ),
    .X(_00818_));
 sg13g2_and2_1 _06279_ (.A(_00817_),
    .B(_00818_),
    .X(_00819_));
 sg13g2_buf_2 _06280_ (.A(_00819_),
    .X(_00820_));
 sg13g2_nor2b_1 _06281_ (.A(_00091_),
    .B_N(_00820_),
    .Y(_00821_));
 sg13g2_buf_1 _06282_ (.A(_00821_),
    .X(_00822_));
 sg13g2_buf_2 _06283_ (.A(debug_instr_valid),
    .X(_00823_));
 sg13g2_o21ai_1 _06284_ (.B1(_00823_),
    .Y(_00824_),
    .A1(\i_tinyqv.cpu.is_jal ),
    .A2(\i_tinyqv.cpu.is_auipc ));
 sg13g2_inv_1 _06285_ (.Y(_00825_),
    .A(_00824_));
 sg13g2_nor2_2 _06286_ (.A(net203),
    .B(_00825_),
    .Y(_00826_));
 sg13g2_o21ai_1 _06287_ (.B1(_00826_),
    .Y(_00827_),
    .A1(_00799_),
    .A2(_00816_));
 sg13g2_nor2_2 _06288_ (.A(_00822_),
    .B(_00824_),
    .Y(_00828_));
 sg13g2_buf_1 _06289_ (.A(\i_tinyqv.cpu.instr_data_start[15] ),
    .X(_00829_));
 sg13g2_nand2_1 _06290_ (.Y(_00830_),
    .A(net337),
    .B(_00829_));
 sg13g2_buf_1 _06291_ (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .X(_00831_));
 sg13g2_nand2b_1 _06292_ (.Y(_00832_),
    .B(_00831_),
    .A_N(_00791_));
 sg13g2_buf_1 _06293_ (.A(net336),
    .X(_00833_));
 sg13g2_a21oi_1 _06294_ (.A1(_00830_),
    .A2(_00832_),
    .Y(_00834_),
    .B1(net285));
 sg13g2_buf_8 _06295_ (.A(net337),
    .X(_00835_));
 sg13g2_buf_1 _06296_ (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .X(_00836_));
 sg13g2_nand2b_1 _06297_ (.Y(_00837_),
    .B(net334),
    .A_N(_00835_));
 sg13g2_a21oi_1 _06298_ (.A1(net285),
    .A2(_00837_),
    .Y(_00838_),
    .B1(net288));
 sg13g2_buf_8 _06299_ (.A(net284),
    .X(_00839_));
 sg13g2_buf_1 _06300_ (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .X(_00840_));
 sg13g2_inv_1 _06301_ (.Y(_00841_),
    .A(_00840_));
 sg13g2_nor2_1 _06302_ (.A(net337),
    .B(net336),
    .Y(_00842_));
 sg13g2_buf_1 _06303_ (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .X(_00843_));
 sg13g2_inv_1 _06304_ (.Y(_00844_),
    .A(net333));
 sg13g2_a22oi_1 _06305_ (.Y(_00845_),
    .B1(_00842_),
    .B2(_00844_),
    .A2(_00841_),
    .A1(net241));
 sg13g2_o21ai_1 _06306_ (.B1(_00845_),
    .Y(_00846_),
    .A1(_00834_),
    .A2(_00838_));
 sg13g2_buf_1 _06307_ (.A(net288),
    .X(_00847_));
 sg13g2_nor2b_1 _06308_ (.A(net284),
    .B_N(net336),
    .Y(_00848_));
 sg13g2_nand3_1 _06309_ (.B(\i_tinyqv.cpu.instr_data_start[23] ),
    .C(_00848_),
    .A(net240),
    .Y(_00849_));
 sg13g2_nand2_1 _06310_ (.Y(_00850_),
    .A(net240),
    .B(_00834_));
 sg13g2_nand3_1 _06311_ (.B(_00849_),
    .C(_00850_),
    .A(_00846_),
    .Y(_00851_));
 sg13g2_buf_1 _06312_ (.A(_00851_),
    .X(_00852_));
 sg13g2_nand2_1 _06313_ (.Y(_00853_),
    .A(_00828_),
    .B(_00852_));
 sg13g2_nand2_1 _06314_ (.Y(_00854_),
    .A(_00827_),
    .B(_00853_));
 sg13g2_buf_1 _06315_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .X(_00855_));
 sg13g2_inv_1 _06316_ (.Y(_00856_),
    .A(net332));
 sg13g2_buf_8 _06317_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .X(_00857_));
 sg13g2_buf_1 _06318_ (.A(net331),
    .X(_00858_));
 sg13g2_buf_1 _06319_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .X(_00859_));
 sg13g2_buf_8 _06320_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .X(_00860_));
 sg13g2_and2_1 _06321_ (.A(_00859_),
    .B(_00860_),
    .X(_00861_));
 sg13g2_buf_1 _06322_ (.A(_00861_),
    .X(_00862_));
 sg13g2_buf_8 _06323_ (.A(_00859_),
    .X(_00863_));
 sg13g2_nor2_1 _06324_ (.A(net282),
    .B(_00860_),
    .Y(_00864_));
 sg13g2_a22oi_1 _06325_ (.Y(_00865_),
    .B1(_00864_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .A2(_00862_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ));
 sg13g2_nor3_1 _06326_ (.A(_00856_),
    .B(_00858_),
    .C(_00865_),
    .Y(_00866_));
 sg13g2_nor2_1 _06327_ (.A(_00860_),
    .B(_00857_),
    .Y(_00867_));
 sg13g2_and2_1 _06328_ (.A(_00860_),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .X(_00868_));
 sg13g2_buf_1 _06329_ (.A(_00868_),
    .X(_00869_));
 sg13g2_a22oi_1 _06330_ (.Y(_00870_),
    .B1(_00869_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .A2(_00867_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ));
 sg13g2_nor2b_1 _06331_ (.A(net332),
    .B_N(_00859_),
    .Y(_00871_));
 sg13g2_buf_2 _06332_ (.A(_00871_),
    .X(_00872_));
 sg13g2_nor2b_1 _06333_ (.A(_00870_),
    .B_N(_00872_),
    .Y(_00873_));
 sg13g2_buf_8 _06334_ (.A(net282),
    .X(_00874_));
 sg13g2_nor2b_1 _06335_ (.A(net331),
    .B_N(_00860_),
    .Y(_00875_));
 sg13g2_and2_1 _06336_ (.A(net332),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .X(_00876_));
 sg13g2_buf_8 _06337_ (.A(net332),
    .X(_00877_));
 sg13g2_nor2b_1 _06338_ (.A(net281),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .Y(_00878_));
 sg13g2_buf_8 _06339_ (.A(_00860_),
    .X(_00879_));
 sg13g2_nor2b_1 _06340_ (.A(net280),
    .B_N(net331),
    .Y(_00880_));
 sg13g2_a22oi_1 _06341_ (.Y(_00881_),
    .B1(_00878_),
    .B2(_00880_),
    .A2(_00876_),
    .A1(_00875_));
 sg13g2_nand3b_1 _06342_ (.B(net331),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .Y(_00882_),
    .A_N(net282));
 sg13g2_nand3b_1 _06343_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .C(_00863_),
    .Y(_00883_),
    .A_N(_00857_));
 sg13g2_nand2b_1 _06344_ (.Y(_00884_),
    .B(net280),
    .A_N(net332));
 sg13g2_a21o_1 _06345_ (.A2(_00883_),
    .A1(_00882_),
    .B1(_00884_),
    .X(_00885_));
 sg13g2_o21ai_1 _06346_ (.B1(_00885_),
    .Y(_00886_),
    .A1(net239),
    .A2(_00881_));
 sg13g2_nor3_1 _06347_ (.A(_00866_),
    .B(_00873_),
    .C(_00886_),
    .Y(_00887_));
 sg13g2_buf_2 _06348_ (.A(\i_tinyqv.cpu.alu_op[3] ),
    .X(_00888_));
 sg13g2_buf_1 _06349_ (.A(_00094_),
    .X(_00889_));
 sg13g2_nor2b_1 _06350_ (.A(_00888_),
    .B_N(_00889_),
    .Y(_00890_));
 sg13g2_a21o_1 _06351_ (.A2(_00820_),
    .A1(_00888_),
    .B1(_00890_),
    .X(_00891_));
 sg13g2_buf_1 _06352_ (.A(_00891_),
    .X(_00892_));
 sg13g2_buf_2 _06353_ (.A(\i_tinyqv.cpu.is_branch ),
    .X(_00893_));
 sg13g2_buf_1 _06354_ (.A(\i_tinyqv.cpu.is_alu_reg ),
    .X(_00894_));
 sg13g2_o21ai_1 _06355_ (.B1(_00823_),
    .Y(_00895_),
    .A1(_00893_),
    .A2(_00894_));
 sg13g2_buf_2 _06356_ (.A(_00895_),
    .X(_00896_));
 sg13g2_buf_1 _06357_ (.A(_00896_),
    .X(_00897_));
 sg13g2_inv_1 _06358_ (.Y(_00898_),
    .A(net336));
 sg13g2_nor2b_1 _06359_ (.A(_00789_),
    .B_N(net337),
    .Y(_00899_));
 sg13g2_buf_2 _06360_ (.A(_00899_),
    .X(_00900_));
 sg13g2_and2_1 _06361_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .B(net282),
    .X(_00901_));
 sg13g2_buf_2 _06362_ (.A(_00901_),
    .X(_00902_));
 sg13g2_nand4_1 _06363_ (.B(_00900_),
    .C(_00902_),
    .A(_00898_),
    .Y(_00903_),
    .D(_00867_));
 sg13g2_nor2b_1 _06364_ (.A(net280),
    .B_N(net332),
    .Y(_00904_));
 sg13g2_mux2_1 _06365_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .S(_00863_),
    .X(_00905_));
 sg13g2_nand3_1 _06366_ (.B(_00904_),
    .C(_00905_),
    .A(net283),
    .Y(_00906_));
 sg13g2_nor2b_1 _06367_ (.A(_00095_),
    .B_N(net282),
    .Y(_00907_));
 sg13g2_nor2b_1 _06368_ (.A(net239),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .Y(_00908_));
 sg13g2_and3_1 _06369_ (.X(_00909_),
    .A(_00855_),
    .B(net280),
    .C(net331));
 sg13g2_o21ai_1 _06370_ (.B1(_00909_),
    .Y(_00910_),
    .A1(_00907_),
    .A2(_00908_));
 sg13g2_nand3_1 _06371_ (.B(_00872_),
    .C(_00880_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .Y(_00911_));
 sg13g2_nand4_1 _06372_ (.B(_00906_),
    .C(_00910_),
    .A(_00903_),
    .Y(_00912_),
    .D(_00911_));
 sg13g2_nor3_1 _06373_ (.A(_00892_),
    .B(net224),
    .C(_00912_),
    .Y(_00913_));
 sg13g2_inv_1 _06374_ (.Y(_00914_),
    .A(net224));
 sg13g2_buf_1 _06375_ (.A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .X(_00915_));
 sg13g2_buf_2 _06376_ (.A(\i_tinyqv.cpu.imm[14] ),
    .X(_00916_));
 sg13g2_buf_1 _06377_ (.A(\i_tinyqv.cpu.imm[22] ),
    .X(_00917_));
 sg13g2_mux4_1 _06378_ (.S0(net284),
    .A0(_00915_),
    .A1(_00916_),
    .A2(_00917_),
    .A3(\i_tinyqv.cpu.imm[30] ),
    .S1(net285),
    .X(_00918_));
 sg13g2_buf_1 _06379_ (.A(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .X(_00919_));
 sg13g2_buf_1 _06380_ (.A(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .X(_00920_));
 sg13g2_buf_2 _06381_ (.A(\i_tinyqv.cpu.imm[18] ),
    .X(_00921_));
 sg13g2_mux4_1 _06382_ (.S0(net284),
    .A0(net330),
    .A1(_00920_),
    .A2(_00921_),
    .A3(\i_tinyqv.cpu.imm[26] ),
    .S1(net285),
    .X(_00922_));
 sg13g2_inv_1 _06383_ (.Y(_00923_),
    .A(_00790_));
 sg13g2_buf_1 _06384_ (.A(_00923_),
    .X(_00924_));
 sg13g2_mux2_1 _06385_ (.A0(_00918_),
    .A1(_00922_),
    .S(net223),
    .X(_00925_));
 sg13g2_buf_1 _06386_ (.A(_00925_),
    .X(_00926_));
 sg13g2_nor3_1 _06387_ (.A(_00892_),
    .B(_00914_),
    .C(_00926_),
    .Y(_00927_));
 sg13g2_a21oi_1 _06388_ (.A1(_00887_),
    .A2(_00913_),
    .Y(_00928_),
    .B1(_00927_));
 sg13g2_or4_1 _06389_ (.A(_00866_),
    .B(_00873_),
    .C(_00886_),
    .D(_00912_),
    .X(_00929_));
 sg13g2_buf_2 _06390_ (.A(_00929_),
    .X(_00930_));
 sg13g2_nand2b_1 _06391_ (.Y(_00931_),
    .B(net224),
    .A_N(_00926_));
 sg13g2_and2_1 _06392_ (.A(_00892_),
    .B(_00931_),
    .X(_00932_));
 sg13g2_o21ai_1 _06393_ (.B1(_00932_),
    .Y(_00933_),
    .A1(net224),
    .A2(_00930_));
 sg13g2_nand2_1 _06394_ (.Y(_00934_),
    .A(_00928_),
    .B(_00933_));
 sg13g2_o21ai_1 _06395_ (.B1(_00931_),
    .Y(_00935_),
    .A1(net224),
    .A2(_00930_));
 sg13g2_buf_1 _06396_ (.A(_00935_),
    .X(_00936_));
 sg13g2_mux2_1 _06397_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .S(_00860_),
    .X(_00937_));
 sg13g2_inv_2 _06398_ (.Y(_00938_),
    .A(net331));
 sg13g2_a221oi_1 _06399_ (.B2(_00938_),
    .C1(_00856_),
    .B1(_00937_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .Y(_00939_),
    .A2(_00869_));
 sg13g2_a21oi_1 _06400_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .A2(_00880_),
    .Y(_00940_),
    .B1(net281));
 sg13g2_or3_1 _06401_ (.A(_00874_),
    .B(_00939_),
    .C(_00940_),
    .X(_00941_));
 sg13g2_nor2b_1 _06402_ (.A(net281),
    .B_N(net280),
    .Y(_00942_));
 sg13g2_a22oi_1 _06403_ (.Y(_00943_),
    .B1(_00942_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .A2(_00904_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ));
 sg13g2_nand3b_1 _06404_ (.B(net283),
    .C(net239),
    .Y(_00944_),
    .A_N(_00943_));
 sg13g2_nor2b_1 _06405_ (.A(net239),
    .B_N(_00855_),
    .Y(_00945_));
 sg13g2_a22oi_1 _06406_ (.Y(_00946_),
    .B1(_00945_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .A2(_00872_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ));
 sg13g2_nand2b_1 _06407_ (.Y(_00947_),
    .B(_00880_),
    .A_N(_00946_));
 sg13g2_nor2b_1 _06408_ (.A(_00092_),
    .B_N(net331),
    .Y(_00948_));
 sg13g2_nor2b_1 _06409_ (.A(net331),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .Y(_00949_));
 sg13g2_and3_1 _06410_ (.X(_00950_),
    .A(net332),
    .B(net282),
    .C(net280));
 sg13g2_o21ai_1 _06411_ (.B1(_00950_),
    .Y(_00951_),
    .A1(_00948_),
    .A2(_00949_));
 sg13g2_nor2_1 _06412_ (.A(net332),
    .B(net282),
    .Y(_00952_));
 sg13g2_nand4_1 _06413_ (.B(_00900_),
    .C(_00875_),
    .A(net336),
    .Y(_00953_),
    .D(_00952_));
 sg13g2_mux2_1 _06414_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .S(_00860_),
    .X(_00954_));
 sg13g2_nand3_1 _06415_ (.B(_00872_),
    .C(_00954_),
    .A(_00938_),
    .Y(_00955_));
 sg13g2_nand3_1 _06416_ (.B(_00869_),
    .C(_00952_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .Y(_00956_));
 sg13g2_and4_1 _06417_ (.A(_00951_),
    .B(_00953_),
    .C(_00955_),
    .D(_00956_),
    .X(_00957_));
 sg13g2_nand4_1 _06418_ (.B(_00944_),
    .C(_00947_),
    .A(_00941_),
    .Y(_00958_),
    .D(_00957_));
 sg13g2_buf_2 _06419_ (.A(_00958_),
    .X(_00959_));
 sg13g2_buf_2 _06420_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .X(_00960_));
 sg13g2_buf_2 _06421_ (.A(\i_tinyqv.cpu.imm[15] ),
    .X(_00961_));
 sg13g2_mux4_1 _06422_ (.S0(net284),
    .A0(_00960_),
    .A1(_00961_),
    .A2(\i_tinyqv.cpu.imm[23] ),
    .A3(\i_tinyqv.cpu.imm[31] ),
    .S1(net285),
    .X(_00962_));
 sg13g2_buf_1 _06423_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .X(_00963_));
 sg13g2_buf_1 _06424_ (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .X(_00964_));
 sg13g2_buf_2 _06425_ (.A(\i_tinyqv.cpu.imm[19] ),
    .X(_00965_));
 sg13g2_mux4_1 _06426_ (.S0(net284),
    .A0(net329),
    .A1(net328),
    .A2(_00965_),
    .A3(\i_tinyqv.cpu.imm[27] ),
    .S1(net336),
    .X(_00966_));
 sg13g2_mux2_1 _06427_ (.A0(_00962_),
    .A1(_00966_),
    .S(_00923_),
    .X(_00967_));
 sg13g2_buf_1 _06428_ (.A(_00967_),
    .X(_00968_));
 sg13g2_nand2b_1 _06429_ (.Y(_00969_),
    .B(_00896_),
    .A_N(_00968_));
 sg13g2_o21ai_1 _06430_ (.B1(_00969_),
    .Y(_00970_),
    .A1(_00897_),
    .A2(_00959_));
 sg13g2_buf_2 _06431_ (.A(_00970_),
    .X(_00971_));
 sg13g2_a21oi_1 _06432_ (.A1(_00888_),
    .A2(_00820_),
    .Y(_00972_),
    .B1(_00890_));
 sg13g2_buf_2 _06433_ (.A(_00972_),
    .X(_00973_));
 sg13g2_o21ai_1 _06434_ (.B1(_00973_),
    .Y(_00974_),
    .A1(_00936_),
    .A2(_00971_));
 sg13g2_mux2_1 _06435_ (.A0(_00930_),
    .A1(_00926_),
    .S(net224),
    .X(_00975_));
 sg13g2_buf_2 _06436_ (.A(_00975_),
    .X(_00976_));
 sg13g2_mux2_1 _06437_ (.A0(_00959_),
    .A1(_00968_),
    .S(net224),
    .X(_00977_));
 sg13g2_buf_2 _06438_ (.A(_00977_),
    .X(_00978_));
 sg13g2_buf_1 _06439_ (.A(_00892_),
    .X(_00979_));
 sg13g2_o21ai_1 _06440_ (.B1(net187),
    .Y(_00980_),
    .A1(_00976_),
    .A2(_00978_));
 sg13g2_nand2_1 _06441_ (.Y(_00981_),
    .A(_00974_),
    .B(_00980_));
 sg13g2_o21ai_1 _06442_ (.B1(_00981_),
    .Y(_00982_),
    .A1(_00854_),
    .A2(_00934_));
 sg13g2_inv_1 _06443_ (.Y(_00983_),
    .A(_00826_));
 sg13g2_nand3b_1 _06444_ (.B(net291),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .Y(_00984_),
    .A_N(net290));
 sg13g2_nand3b_1 _06445_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .C(net290),
    .Y(_00985_),
    .A_N(net291));
 sg13g2_a21o_1 _06446_ (.A2(_00985_),
    .A1(_00984_),
    .B1(_00788_),
    .X(_00986_));
 sg13g2_nor2b_1 _06447_ (.A(net291),
    .B_N(net292),
    .Y(_00987_));
 sg13g2_nor2b_1 _06448_ (.A(net290),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .Y(_00988_));
 sg13g2_nor2b_1 _06449_ (.A(net242),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .Y(_00989_));
 sg13g2_a221oi_1 _06450_ (.B2(_00770_),
    .C1(net289),
    .B1(_00989_),
    .A1(_00987_),
    .Y(_00990_),
    .A2(_00988_));
 sg13g2_a21o_1 _06451_ (.A2(_00986_),
    .A1(net289),
    .B1(_00990_),
    .X(_00991_));
 sg13g2_nand2_1 _06452_ (.Y(_00992_),
    .A(_00779_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ));
 sg13g2_nand3b_1 _06453_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .C(_00766_),
    .Y(_00993_),
    .A_N(net292));
 sg13g2_o21ai_1 _06454_ (.B1(_00993_),
    .Y(_00994_),
    .A1(net289),
    .A2(_00992_));
 sg13g2_nor2_1 _06455_ (.A(_00779_),
    .B(net291),
    .Y(_00995_));
 sg13g2_inv_1 _06456_ (.Y(_00996_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ));
 sg13g2_nand2b_1 _06457_ (.Y(_00997_),
    .B(net339),
    .A_N(_00768_));
 sg13g2_nand3b_1 _06458_ (.B(net290),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .Y(_00998_),
    .A_N(net339));
 sg13g2_o21ai_1 _06459_ (.B1(_00998_),
    .Y(_00999_),
    .A1(_00996_),
    .A2(_00997_));
 sg13g2_a22oi_1 _06460_ (.Y(_01000_),
    .B1(_00995_),
    .B2(_00999_),
    .A2(_00994_),
    .A1(_00797_));
 sg13g2_and3_1 _06461_ (.X(_01001_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .B(_00785_),
    .C(_00813_));
 sg13g2_mux2_1 _06462_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .S(net338),
    .X(_01002_));
 sg13g2_and3_1 _06463_ (.X(_01003_),
    .A(_00780_),
    .B(_00810_),
    .C(_01002_));
 sg13g2_nand2b_1 _06464_ (.Y(_01004_),
    .B(net339),
    .A_N(_00095_));
 sg13g2_nand2b_1 _06465_ (.Y(_01005_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .A_N(_00766_));
 sg13g2_nand3_1 _06466_ (.B(_00768_),
    .C(net291),
    .A(_00773_),
    .Y(_01006_));
 sg13g2_a21oi_1 _06467_ (.A1(_01004_),
    .A2(_01005_),
    .Y(_01007_),
    .B1(_01006_));
 sg13g2_nand2b_1 _06468_ (.Y(_01008_),
    .B(net337),
    .A_N(_00789_));
 sg13g2_buf_1 _06469_ (.A(_01008_),
    .X(_01009_));
 sg13g2_nand2b_1 _06470_ (.Y(_01010_),
    .B(net292),
    .A_N(net338));
 sg13g2_nor4_1 _06471_ (.A(net336),
    .B(_01009_),
    .C(_01010_),
    .D(_00997_),
    .Y(_01011_));
 sg13g2_nor4_2 _06472_ (.A(_01001_),
    .B(_01003_),
    .C(_01007_),
    .Y(_01012_),
    .D(_01011_));
 sg13g2_and3_1 _06473_ (.X(_01013_),
    .A(_00991_),
    .B(_01000_),
    .C(_01012_));
 sg13g2_buf_1 _06474_ (.A(_01013_),
    .X(_01014_));
 sg13g2_inv_1 _06475_ (.Y(_01015_),
    .A(net337));
 sg13g2_buf_1 _06476_ (.A(_01015_),
    .X(_01016_));
 sg13g2_buf_1 _06477_ (.A(\i_tinyqv.cpu.instr_data_start[18] ),
    .X(_01017_));
 sg13g2_a21o_1 _06478_ (.A2(net327),
    .A1(net238),
    .B1(_00898_),
    .X(_01018_));
 sg13g2_buf_1 _06479_ (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .X(_01019_));
 sg13g2_nand2_1 _06480_ (.Y(_01020_),
    .A(net284),
    .B(net326));
 sg13g2_buf_1 _06481_ (.A(\i_tinyqv.cpu.instr_data_start[6] ),
    .X(_01021_));
 sg13g2_nand2b_1 _06482_ (.Y(_01022_),
    .B(_01021_),
    .A_N(_00835_));
 sg13g2_a21oi_1 _06483_ (.A1(_01020_),
    .A2(_01022_),
    .Y(_01023_),
    .B1(net285));
 sg13g2_a21oi_1 _06484_ (.A1(_00923_),
    .A2(_01018_),
    .Y(_01024_),
    .B1(_01023_));
 sg13g2_buf_1 _06485_ (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .X(_01025_));
 sg13g2_buf_2 _06486_ (.A(\i_tinyqv.cpu.pc[2] ),
    .X(_01026_));
 sg13g2_inv_1 _06487_ (.Y(_01027_),
    .A(_01026_));
 sg13g2_nand2_1 _06488_ (.Y(_01028_),
    .A(_01027_),
    .B(_00842_));
 sg13g2_o21ai_1 _06489_ (.B1(_01028_),
    .Y(_01029_),
    .A1(net238),
    .A2(net325));
 sg13g2_buf_2 _06490_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .X(_01030_));
 sg13g2_and2_1 _06491_ (.A(_01030_),
    .B(_00848_),
    .X(_01031_));
 sg13g2_o21ai_1 _06492_ (.B1(net240),
    .Y(_01032_),
    .A1(_01023_),
    .A2(_01031_));
 sg13g2_o21ai_1 _06493_ (.B1(_01032_),
    .Y(_01033_),
    .A1(_01024_),
    .A2(_01029_));
 sg13g2_nand2_1 _06494_ (.Y(_01034_),
    .A(_00828_),
    .B(_01033_));
 sg13g2_o21ai_1 _06495_ (.B1(_01034_),
    .Y(_01035_),
    .A1(_00983_),
    .A2(net163));
 sg13g2_buf_2 _06496_ (.A(_01035_),
    .X(_01036_));
 sg13g2_and2_1 _06497_ (.A(net293),
    .B(net287),
    .X(_01037_));
 sg13g2_nand2b_1 _06498_ (.Y(_01038_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .A_N(_00768_));
 sg13g2_nand3b_1 _06499_ (.B(net290),
    .C(_00773_),
    .Y(_01039_),
    .A_N(_00096_));
 sg13g2_o21ai_1 _06500_ (.B1(_01039_),
    .Y(_01040_),
    .A1(net242),
    .A2(_01038_));
 sg13g2_nand2b_1 _06501_ (.Y(_01041_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .A_N(net290));
 sg13g2_nand3_1 _06502_ (.B(net290),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A(net293),
    .Y(_01042_));
 sg13g2_o21ai_1 _06503_ (.B1(_01042_),
    .Y(_01043_),
    .A1(_00767_),
    .A2(_01041_));
 sg13g2_a22oi_1 _06504_ (.Y(_01044_),
    .B1(_01043_),
    .B2(_00987_),
    .A2(_01040_),
    .A1(_01037_));
 sg13g2_buf_2 _06505_ (.A(_01044_),
    .X(_01045_));
 sg13g2_mux4_1 _06506_ (.S0(net292),
    .A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .A2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .A3(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .S1(net338),
    .X(_01046_));
 sg13g2_nand3b_1 _06507_ (.B(_00804_),
    .C(_01046_),
    .Y(_01047_),
    .A_N(_00767_));
 sg13g2_nor2_1 _06508_ (.A(net290),
    .B(_00775_),
    .Y(_01048_));
 sg13g2_nand3_1 _06509_ (.B(_00810_),
    .C(_01048_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .Y(_01049_));
 sg13g2_mux2_1 _06510_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .S(net339),
    .X(_01050_));
 sg13g2_nand3_1 _06511_ (.B(_00797_),
    .C(_01050_),
    .A(net242),
    .Y(_01051_));
 sg13g2_mux2_1 _06512_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .S(_00769_),
    .X(_01052_));
 sg13g2_nand3_1 _06513_ (.B(_00810_),
    .C(_01052_),
    .A(net286),
    .Y(_01053_));
 sg13g2_and4_1 _06514_ (.A(_01047_),
    .B(_01049_),
    .C(_01051_),
    .D(_01053_),
    .X(_01054_));
 sg13g2_buf_8 _06515_ (.A(_01054_),
    .X(_01055_));
 sg13g2_nand2_1 _06516_ (.Y(_01056_),
    .A(_01045_),
    .B(_01055_));
 sg13g2_buf_2 _06517_ (.A(_01056_),
    .X(_01057_));
 sg13g2_buf_2 _06518_ (.A(\i_tinyqv.cpu.instr_data_start[13] ),
    .X(_01058_));
 sg13g2_nand2_1 _06519_ (.Y(_01059_),
    .A(net241),
    .B(_01058_));
 sg13g2_nand2b_1 _06520_ (.Y(_01060_),
    .B(\i_tinyqv.cpu.instr_data_start[5] ),
    .A_N(net241));
 sg13g2_a21oi_1 _06521_ (.A1(_01059_),
    .A2(_01060_),
    .Y(_01061_),
    .B1(net285));
 sg13g2_buf_1 _06522_ (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .X(_01062_));
 sg13g2_nand2b_1 _06523_ (.Y(_01063_),
    .B(net324),
    .A_N(net241));
 sg13g2_a21oi_1 _06524_ (.A1(_00833_),
    .A2(_01063_),
    .Y(_01064_),
    .B1(net240));
 sg13g2_buf_2 _06525_ (.A(\i_tinyqv.cpu.instr_data_start[9] ),
    .X(_01065_));
 sg13g2_inv_2 _06526_ (.Y(_01066_),
    .A(_01065_));
 sg13g2_buf_2 _06527_ (.A(\i_tinyqv.cpu.pc[1] ),
    .X(_01067_));
 sg13g2_inv_1 _06528_ (.Y(_01068_),
    .A(_01067_));
 sg13g2_a22oi_1 _06529_ (.Y(_01069_),
    .B1(_00842_),
    .B2(_01068_),
    .A2(_01066_),
    .A1(net241));
 sg13g2_o21ai_1 _06530_ (.B1(_01069_),
    .Y(_01070_),
    .A1(_01061_),
    .A2(_01064_));
 sg13g2_buf_1 _06531_ (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .X(_01071_));
 sg13g2_and2_1 _06532_ (.A(net323),
    .B(_00848_),
    .X(_01072_));
 sg13g2_o21ai_1 _06533_ (.B1(net240),
    .Y(_01073_),
    .A1(_01061_),
    .A2(_01072_));
 sg13g2_nand2_1 _06534_ (.Y(_01074_),
    .A(_01070_),
    .B(_01073_));
 sg13g2_a22oi_1 _06535_ (.Y(_01075_),
    .B1(_01074_),
    .B2(_00828_),
    .A2(_01057_),
    .A1(_00826_));
 sg13g2_buf_2 _06536_ (.A(_01075_),
    .X(_01076_));
 sg13g2_mux2_1 _06537_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .S(net283),
    .X(_01077_));
 sg13g2_nand2_1 _06538_ (.Y(_01078_),
    .A(_00872_),
    .B(_01077_));
 sg13g2_nor2b_1 _06539_ (.A(net283),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .Y(_01079_));
 sg13g2_and2_1 _06540_ (.A(net283),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .X(_01080_));
 sg13g2_a22oi_1 _06541_ (.Y(_01081_),
    .B1(_01080_),
    .B2(_00952_),
    .A2(_01079_),
    .A1(_00902_));
 sg13g2_buf_8 _06542_ (.A(net280),
    .X(_01082_));
 sg13g2_mux2_1 _06543_ (.A0(_01078_),
    .A1(_01081_),
    .S(net237),
    .X(_01083_));
 sg13g2_a221oi_1 _06544_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .C1(net281),
    .B1(_00864_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .Y(_01084_),
    .A2(_00862_));
 sg13g2_inv_1 _06545_ (.Y(_01085_),
    .A(_00096_));
 sg13g2_a221oi_1 _06546_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .C1(_00856_),
    .B1(_00864_),
    .A1(_01085_),
    .Y(_01086_),
    .A2(_00862_));
 sg13g2_or3_1 _06547_ (.A(_00938_),
    .B(_01084_),
    .C(_01086_),
    .X(_01087_));
 sg13g2_and3_1 _06548_ (.X(_01088_),
    .A(net283),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .C(_00904_));
 sg13g2_and3_1 _06549_ (.X(_01089_),
    .A(_00938_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .C(_00942_));
 sg13g2_o21ai_1 _06550_ (.B1(net239),
    .Y(_01090_),
    .A1(_01088_),
    .A2(_01089_));
 sg13g2_mux2_1 _06551_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .S(net283),
    .X(_01091_));
 sg13g2_a22oi_1 _06552_ (.Y(_01092_),
    .B1(_01091_),
    .B2(_01082_),
    .A2(_00867_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ));
 sg13g2_nand2b_1 _06553_ (.Y(_01093_),
    .B(_00945_),
    .A_N(_01092_));
 sg13g2_and4_1 _06554_ (.A(_01083_),
    .B(_01087_),
    .C(_01090_),
    .D(_01093_),
    .X(_01094_));
 sg13g2_buf_2 _06555_ (.A(_01094_),
    .X(_01095_));
 sg13g2_buf_2 _06556_ (.A(\i_tinyqv.cpu.imm[17] ),
    .X(_01096_));
 sg13g2_buf_1 _06557_ (.A(\i_tinyqv.cpu.imm[21] ),
    .X(_01097_));
 sg13g2_mux4_1 _06558_ (.S0(net288),
    .A0(_01096_),
    .A1(_01097_),
    .A2(\i_tinyqv.cpu.imm[25] ),
    .A3(\i_tinyqv.cpu.imm[29] ),
    .S1(net241),
    .X(_01098_));
 sg13g2_buf_1 _06559_ (.A(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .X(_01099_));
 sg13g2_buf_2 _06560_ (.A(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .X(_01100_));
 sg13g2_buf_2 _06561_ (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .X(_01101_));
 sg13g2_buf_1 _06562_ (.A(\i_tinyqv.cpu.imm[13] ),
    .X(_01102_));
 sg13g2_mux4_1 _06563_ (.S0(net288),
    .A0(_01099_),
    .A1(_01100_),
    .A2(_01101_),
    .A3(_01102_),
    .S1(net241),
    .X(_01103_));
 sg13g2_buf_1 _06564_ (.A(_00898_),
    .X(_01104_));
 sg13g2_mux2_1 _06565_ (.A0(_01098_),
    .A1(_01103_),
    .S(net236),
    .X(_01105_));
 sg13g2_buf_1 _06566_ (.A(_01105_),
    .X(_01106_));
 sg13g2_nor2_1 _06567_ (.A(_00914_),
    .B(_01106_),
    .Y(_01107_));
 sg13g2_a21oi_2 _06568_ (.B1(_01107_),
    .Y(_01108_),
    .A2(_01095_),
    .A1(_00914_));
 sg13g2_buf_2 _06569_ (.A(\i_tinyqv.cpu.imm[16] ),
    .X(_01109_));
 sg13g2_buf_2 _06570_ (.A(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .X(_01110_));
 sg13g2_mux4_1 _06571_ (.S0(_00792_),
    .A0(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .A1(_01109_),
    .A2(_01110_),
    .A3(\i_tinyqv.cpu.imm[24] ),
    .S1(net284),
    .X(_01111_));
 sg13g2_buf_2 _06572_ (.A(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .X(_01112_));
 sg13g2_buf_2 _06573_ (.A(\i_tinyqv.cpu.imm[12] ),
    .X(_01113_));
 sg13g2_buf_2 _06574_ (.A(\i_tinyqv.cpu.imm[20] ),
    .X(_01114_));
 sg13g2_mux4_1 _06575_ (.S0(net337),
    .A0(_01112_),
    .A1(_01113_),
    .A2(_01114_),
    .A3(\i_tinyqv.cpu.imm[28] ),
    .S1(_00792_),
    .X(_01115_));
 sg13g2_and2_1 _06576_ (.A(net288),
    .B(_01115_),
    .X(_01116_));
 sg13g2_a21oi_2 _06577_ (.B1(_01116_),
    .Y(_01117_),
    .A2(_01111_),
    .A1(_00923_));
 sg13g2_mux2_1 _06578_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .S(net237),
    .X(_01118_));
 sg13g2_nand2_1 _06579_ (.Y(_01119_),
    .A(_01082_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_o21ai_1 _06580_ (.B1(_01119_),
    .Y(_01120_),
    .A1(net237),
    .A2(_00794_));
 sg13g2_mux2_1 _06581_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .S(_00879_),
    .X(_01121_));
 sg13g2_and2_1 _06582_ (.A(_00872_),
    .B(_01121_),
    .X(_01122_));
 sg13g2_a221oi_1 _06583_ (.B2(_00902_),
    .C1(_01122_),
    .B1(_01120_),
    .A1(_00945_),
    .Y(_01123_),
    .A2(_01118_));
 sg13g2_nor2_1 _06584_ (.A(net283),
    .B(_00896_),
    .Y(_01124_));
 sg13g2_nand3b_1 _06585_ (.B(net237),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .Y(_01125_),
    .A_N(net239));
 sg13g2_nand3b_1 _06586_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .C(net239),
    .Y(_01126_),
    .A_N(net280));
 sg13g2_a21o_1 _06587_ (.A2(_01126_),
    .A1(_01125_),
    .B1(_00856_),
    .X(_01127_));
 sg13g2_nand3b_1 _06588_ (.B(net237),
    .C(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .Y(_01128_),
    .A_N(_00877_));
 sg13g2_nand3b_1 _06589_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .C(_00877_),
    .Y(_01129_),
    .A_N(_00879_));
 sg13g2_a21o_1 _06590_ (.A2(_01129_),
    .A1(_01128_),
    .B1(net239),
    .X(_01130_));
 sg13g2_nor2_1 _06591_ (.A(net281),
    .B(net237),
    .Y(_01131_));
 sg13g2_mux2_1 _06592_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .S(net282),
    .X(_01132_));
 sg13g2_mux2_1 _06593_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .S(net281),
    .X(_01133_));
 sg13g2_a22oi_1 _06594_ (.Y(_01134_),
    .B1(_01133_),
    .B2(_00862_),
    .A2(_01132_),
    .A1(_01131_));
 sg13g2_nor2_1 _06595_ (.A(_00938_),
    .B(_00896_),
    .Y(_01135_));
 sg13g2_and4_1 _06596_ (.A(_01127_),
    .B(_01130_),
    .C(_01134_),
    .D(_01135_),
    .X(_01136_));
 sg13g2_a221oi_1 _06597_ (.B2(_01124_),
    .C1(_01136_),
    .B1(_01123_),
    .A1(_00896_),
    .Y(_01137_),
    .A2(_01117_));
 sg13g2_buf_1 _06598_ (.A(_01137_),
    .X(_01138_));
 sg13g2_nand2b_1 _06599_ (.Y(_01139_),
    .B(_00973_),
    .A_N(_01138_));
 sg13g2_a21oi_1 _06600_ (.A1(_01076_),
    .A2(_01108_),
    .Y(_01140_),
    .B1(_01139_));
 sg13g2_a21o_1 _06601_ (.A2(_01095_),
    .A1(_00914_),
    .B1(_01107_),
    .X(_01141_));
 sg13g2_nand2_1 _06602_ (.Y(_01142_),
    .A(_00892_),
    .B(_01138_));
 sg13g2_a21oi_1 _06603_ (.A1(_01076_),
    .A2(_01141_),
    .Y(_01143_),
    .B1(_01142_));
 sg13g2_nor2_1 _06604_ (.A(net288),
    .B(net241),
    .Y(_01144_));
 sg13g2_nand2_1 _06605_ (.Y(_01145_),
    .A(net236),
    .B(_01144_));
 sg13g2_buf_2 _06606_ (.A(_01145_),
    .X(_01146_));
 sg13g2_nand2_1 _06607_ (.Y(_01147_),
    .A(_00097_),
    .B(_01146_));
 sg13g2_o21ai_1 _06608_ (.B1(_01147_),
    .Y(_01148_),
    .A1(_00973_),
    .A2(_01146_));
 sg13g2_buf_2 _06609_ (.A(_01148_),
    .X(_01149_));
 sg13g2_nor2b_1 _06610_ (.A(net286),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .Y(_01150_));
 sg13g2_and2_1 _06611_ (.A(net286),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .X(_01151_));
 sg13g2_a22oi_1 _06612_ (.Y(_01152_),
    .B1(_01151_),
    .B2(_00810_),
    .A2(_01150_),
    .A1(_00813_));
 sg13g2_nor2b_1 _06613_ (.A(net286),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .Y(_01153_));
 sg13g2_and2_1 _06614_ (.A(_00804_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .X(_01154_));
 sg13g2_a221oi_1 _06615_ (.B2(_00810_),
    .C1(net287),
    .B1(_01154_),
    .A1(_00813_),
    .Y(_01155_),
    .A2(_01153_));
 sg13g2_a21o_1 _06616_ (.A2(_01152_),
    .A1(net287),
    .B1(_01155_),
    .X(_01156_));
 sg13g2_mux2_1 _06617_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .S(_00775_),
    .X(_01157_));
 sg13g2_nand3_1 _06618_ (.B(net242),
    .C(_01157_),
    .A(_00783_),
    .Y(_01158_));
 sg13g2_nand3b_1 _06619_ (.B(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .C(_00995_),
    .Y(_01159_),
    .A_N(net289));
 sg13g2_a21o_1 _06620_ (.A2(_01159_),
    .A1(_01158_),
    .B1(_00781_),
    .X(_01160_));
 sg13g2_and2_1 _06621_ (.A(_00785_),
    .B(_00813_),
    .X(_01161_));
 sg13g2_mux2_1 _06622_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .S(net242),
    .X(_01162_));
 sg13g2_nor3_1 _06623_ (.A(_00794_),
    .B(_01010_),
    .C(_00997_),
    .Y(_01163_));
 sg13g2_a221oi_1 _06624_ (.B2(_00771_),
    .C1(_01163_),
    .B1(_01162_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .Y(_01164_),
    .A2(_01161_));
 sg13g2_nand2_1 _06625_ (.Y(_01165_),
    .A(_00801_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ));
 sg13g2_nand2b_1 _06626_ (.Y(_01166_),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .A_N(_00801_));
 sg13g2_nand3_1 _06627_ (.B(_01165_),
    .C(_01166_),
    .A(_00788_),
    .Y(_01167_));
 sg13g2_nand2_1 _06628_ (.Y(_01168_),
    .A(net287),
    .B(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_a21oi_1 _06629_ (.A1(net242),
    .A2(_01168_),
    .Y(_01169_),
    .B1(_00997_));
 sg13g2_a21oi_1 _06630_ (.A1(_01167_),
    .A2(_01169_),
    .Y(_01170_),
    .B1(_00825_));
 sg13g2_nand4_1 _06631_ (.B(_01160_),
    .C(_01164_),
    .A(_01156_),
    .Y(_01171_),
    .D(_01170_));
 sg13g2_buf_1 _06632_ (.A(_01171_),
    .X(_01172_));
 sg13g2_nand2b_1 _06633_ (.Y(_01173_),
    .B(_00820_),
    .A_N(_00091_));
 sg13g2_buf_2 _06634_ (.A(_01173_),
    .X(_01174_));
 sg13g2_buf_2 _06635_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .X(_01175_));
 sg13g2_mux2_1 _06636_ (.A0(\i_tinyqv.cpu.instr_data_start[16] ),
    .A1(_01175_),
    .S(_00790_),
    .X(_01176_));
 sg13g2_a21oi_1 _06637_ (.A1(_01016_),
    .A2(_01176_),
    .Y(_01177_),
    .B1(_00898_));
 sg13g2_buf_1 _06638_ (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .X(_01178_));
 sg13g2_buf_2 _06639_ (.A(\i_tinyqv.cpu.instr_data_start[4] ),
    .X(_01179_));
 sg13g2_mux2_1 _06640_ (.A0(_01179_),
    .A1(\i_tinyqv.cpu.instr_data_start[12] ),
    .S(_00791_),
    .X(_01180_));
 sg13g2_a221oi_1 _06641_ (.B2(net288),
    .C1(_00833_),
    .B1(_01180_),
    .A1(_01178_),
    .Y(_01181_),
    .A2(_00900_));
 sg13g2_o21ai_1 _06642_ (.B1(_00825_),
    .Y(_01182_),
    .A1(_01177_),
    .A2(_01181_));
 sg13g2_and2_1 _06643_ (.A(_01174_),
    .B(_01182_),
    .X(_01183_));
 sg13g2_buf_1 _06644_ (.A(_01183_),
    .X(_01184_));
 sg13g2_nand2_2 _06645_ (.Y(_01185_),
    .A(_01172_),
    .B(_01184_));
 sg13g2_nand2_1 _06646_ (.Y(_01186_),
    .A(_01149_),
    .B(_01185_));
 sg13g2_o21ai_1 _06647_ (.B1(_01186_),
    .Y(_01187_),
    .A1(_01140_),
    .A2(_01143_));
 sg13g2_nor3_1 _06648_ (.A(_01149_),
    .B(_01185_),
    .C(_01076_),
    .Y(_01188_));
 sg13g2_xnor2_1 _06649_ (.Y(_01189_),
    .A(net187),
    .B(_01108_));
 sg13g2_o21ai_1 _06650_ (.B1(_01076_),
    .Y(_01190_),
    .A1(_01149_),
    .A2(_01185_));
 sg13g2_o21ai_1 _06651_ (.B1(_01190_),
    .Y(_01191_),
    .A1(_01188_),
    .A2(_01189_));
 sg13g2_nand2_2 _06652_ (.Y(_01192_),
    .A(_01187_),
    .B(_01191_));
 sg13g2_nand2_1 _06653_ (.Y(_01193_),
    .A(_01036_),
    .B(_01192_));
 sg13g2_xnor2_1 _06654_ (.Y(_01194_),
    .A(_00892_),
    .B(_00978_));
 sg13g2_nand3_1 _06655_ (.B(_01000_),
    .C(_01012_),
    .A(_00991_),
    .Y(_01195_));
 sg13g2_buf_2 _06656_ (.A(_01195_),
    .X(_01196_));
 sg13g2_a22oi_1 _06657_ (.Y(_01197_),
    .B1(_01196_),
    .B2(_00826_),
    .A2(_01033_),
    .A1(_00828_));
 sg13g2_buf_2 _06658_ (.A(_01197_),
    .X(_01198_));
 sg13g2_nand3_1 _06659_ (.B(_01187_),
    .C(_01191_),
    .A(_01198_),
    .Y(_01199_));
 sg13g2_o21ai_1 _06660_ (.B1(_01199_),
    .Y(_01200_),
    .A1(_00854_),
    .A2(_01194_));
 sg13g2_nand2_1 _06661_ (.Y(_01201_),
    .A(_00854_),
    .B(_01194_));
 sg13g2_a22oi_1 _06662_ (.Y(\i_tinyqv.cpu.i_core.cy_out ),
    .B1(_01200_),
    .B2(_01201_),
    .A2(_01193_),
    .A1(_00982_));
 sg13g2_buf_1 _06663_ (.A(_00823_),
    .X(_01202_));
 sg13g2_buf_1 _06664_ (.A(\i_tinyqv.cpu.is_load ),
    .X(_01203_));
 sg13g2_buf_1 _06665_ (.A(\i_tinyqv.cpu.is_store ),
    .X(_01204_));
 sg13g2_o21ai_1 _06666_ (.B1(_00098_),
    .Y(_01205_),
    .A1(_01203_),
    .A2(_01204_));
 sg13g2_and2_1 _06667_ (.A(net279),
    .B(_01205_),
    .X(_01206_));
 sg13g2_buf_1 _06668_ (.A(_01206_),
    .X(_01207_));
 sg13g2_inv_1 _06669_ (.Y(_01208_),
    .A(_01207_));
 sg13g2_buf_1 _06670_ (.A(_00088_),
    .X(_01209_));
 sg13g2_nand2_1 _06671_ (.Y(_01210_),
    .A(net240),
    .B(_00839_));
 sg13g2_buf_2 _06672_ (.A(_01210_),
    .X(_01211_));
 sg13g2_nor2_1 _06673_ (.A(_01209_),
    .B(_01211_),
    .Y(_01212_));
 sg13g2_buf_1 _06674_ (.A(_01212_),
    .X(_01213_));
 sg13g2_buf_1 _06675_ (.A(_00099_),
    .X(_01214_));
 sg13g2_inv_1 _06676_ (.Y(_01215_),
    .A(_01214_));
 sg13g2_buf_1 _06677_ (.A(_01215_),
    .X(_01216_));
 sg13g2_buf_1 _06678_ (.A(net235),
    .X(_01217_));
 sg13g2_buf_1 _06679_ (.A(_00090_),
    .X(_01218_));
 sg13g2_buf_1 _06680_ (.A(\i_tinyqv.cpu.is_system ),
    .X(_01219_));
 sg13g2_and2_1 _06681_ (.A(_00823_),
    .B(_01219_),
    .X(_01220_));
 sg13g2_buf_1 _06682_ (.A(\i_tinyqv.cpu.alu_op[0] ),
    .X(_01221_));
 sg13g2_nor2_1 _06683_ (.A(_01221_),
    .B(_00817_),
    .Y(_01222_));
 sg13g2_nor2_1 _06684_ (.A(_01110_),
    .B(_01101_),
    .Y(_01223_));
 sg13g2_nand4_1 _06685_ (.B(_01220_),
    .C(_01222_),
    .A(_01218_),
    .Y(_01224_),
    .D(_01223_));
 sg13g2_buf_1 _06686_ (.A(_01224_),
    .X(_01225_));
 sg13g2_nand2_1 _06687_ (.Y(_01226_),
    .A(_00089_),
    .B(_01225_));
 sg13g2_buf_1 _06688_ (.A(_01226_),
    .X(_01227_));
 sg13g2_and2_1 _06689_ (.A(_01204_),
    .B(\i_tinyqv.cpu.no_write_in_progress ),
    .X(_01228_));
 sg13g2_buf_1 _06690_ (.A(_01228_),
    .X(_01229_));
 sg13g2_nor4_1 _06691_ (.A(_01219_),
    .B(_00893_),
    .C(\i_tinyqv.cpu.is_auipc ),
    .D(_01229_),
    .Y(_01230_));
 sg13g2_nor2_1 _06692_ (.A(\i_tinyqv.cpu.is_jal ),
    .B(\i_tinyqv.cpu.is_jalr ),
    .Y(_01231_));
 sg13g2_inv_1 _06693_ (.Y(_01232_),
    .A(_01231_));
 sg13g2_o21ai_1 _06694_ (.B1(_01202_),
    .Y(_01233_),
    .A1(\i_tinyqv.cpu.is_lui ),
    .A2(_01232_));
 sg13g2_nand4_1 _06695_ (.B(_01230_),
    .C(_01205_),
    .A(net279),
    .Y(_01234_),
    .D(_01233_));
 sg13g2_nor4_2 _06696_ (.A(net222),
    .B(_01174_),
    .C(net186),
    .Y(_01235_),
    .D(_01234_));
 sg13g2_buf_1 _06697_ (.A(_01221_),
    .X(_01236_));
 sg13g2_nand2b_1 _06698_ (.Y(_01237_),
    .B(net242),
    .A_N(_00808_));
 sg13g2_buf_2 _06699_ (.A(_01237_),
    .X(_01238_));
 sg13g2_and3_1 _06700_ (.X(_01239_),
    .A(_00787_),
    .B(_00798_),
    .C(_00815_));
 sg13g2_buf_2 _06701_ (.A(_01239_),
    .X(_01240_));
 sg13g2_a21oi_2 _06702_ (.B1(_00983_),
    .Y(_01241_),
    .A2(_01240_),
    .A1(_01238_));
 sg13g2_and2_1 _06703_ (.A(_00828_),
    .B(_00852_),
    .X(_01242_));
 sg13g2_buf_1 _06704_ (.A(_01242_),
    .X(_01243_));
 sg13g2_nor4_1 _06705_ (.A(_01241_),
    .B(_01243_),
    .C(_00976_),
    .D(_01198_),
    .Y(_01244_));
 sg13g2_nor3_1 _06706_ (.A(_00976_),
    .B(_00971_),
    .C(_01198_),
    .Y(_01245_));
 sg13g2_nor3_1 _06707_ (.A(_01241_),
    .B(_01243_),
    .C(_00971_),
    .Y(_01246_));
 sg13g2_nor4_1 _06708_ (.A(net187),
    .B(_01244_),
    .C(_01245_),
    .D(_01246_),
    .Y(_01247_));
 sg13g2_nor3_1 _06709_ (.A(_01241_),
    .B(_01243_),
    .C(_00978_),
    .Y(_01248_));
 sg13g2_nor4_1 _06710_ (.A(_01241_),
    .B(_01243_),
    .C(_00936_),
    .D(_01198_),
    .Y(_01249_));
 sg13g2_nor3_1 _06711_ (.A(_00936_),
    .B(_00978_),
    .C(_01198_),
    .Y(_01250_));
 sg13g2_nor4_1 _06712_ (.A(_00973_),
    .B(_01248_),
    .C(_01249_),
    .D(_01250_),
    .Y(_01251_));
 sg13g2_nor3_1 _06713_ (.A(_01236_),
    .B(_00889_),
    .C(_00822_),
    .Y(_01252_));
 sg13g2_o21ai_1 _06714_ (.B1(_01252_),
    .Y(_01253_),
    .A1(_01247_),
    .A2(_01251_));
 sg13g2_xnor2_1 _06715_ (.Y(_01254_),
    .A(_01076_),
    .B(_01141_));
 sg13g2_nand3_1 _06716_ (.B(_01184_),
    .C(_01138_),
    .A(_01172_),
    .Y(_01255_));
 sg13g2_buf_1 _06717_ (.A(_01255_),
    .X(_01256_));
 sg13g2_a21o_1 _06718_ (.A2(_01184_),
    .A1(_01172_),
    .B1(_01138_),
    .X(_01257_));
 sg13g2_nand2b_1 _06719_ (.Y(_01258_),
    .B(_00889_),
    .A_N(_01221_));
 sg13g2_buf_1 _06720_ (.A(net285),
    .X(_01259_));
 sg13g2_nand2_2 _06721_ (.Y(_01260_),
    .A(_00924_),
    .B(net238));
 sg13g2_nor2_1 _06722_ (.A(net234),
    .B(_01260_),
    .Y(_01261_));
 sg13g2_nor2_1 _06723_ (.A(\i_tinyqv.cpu.i_core.cmp ),
    .B(_01261_),
    .Y(_01262_));
 sg13g2_a221oi_1 _06724_ (.B2(_01174_),
    .C1(_01262_),
    .B1(_01258_),
    .A1(_01256_),
    .Y(_01263_),
    .A2(_01257_));
 sg13g2_and2_1 _06725_ (.A(_01254_),
    .B(_01263_),
    .X(_01264_));
 sg13g2_nand3_1 _06726_ (.B(_00853_),
    .C(_00971_),
    .A(_00827_),
    .Y(_01265_));
 sg13g2_buf_1 _06727_ (.A(_01265_),
    .X(_01266_));
 sg13g2_o21ai_1 _06728_ (.B1(_00978_),
    .Y(_01267_),
    .A1(_01241_),
    .A2(_01243_));
 sg13g2_buf_1 _06729_ (.A(_01267_),
    .X(_01268_));
 sg13g2_xnor2_1 _06730_ (.Y(_01269_),
    .A(_00976_),
    .B(_01198_));
 sg13g2_a21oi_1 _06731_ (.A1(_01266_),
    .A2(_01268_),
    .Y(_01270_),
    .B1(_01269_));
 sg13g2_nor3_1 _06732_ (.A(net187),
    .B(_00976_),
    .C(_00978_),
    .Y(_01271_));
 sg13g2_nor3_1 _06733_ (.A(_00973_),
    .B(_00936_),
    .C(_00971_),
    .Y(_01272_));
 sg13g2_o21ai_1 _06734_ (.B1(_01036_),
    .Y(_01273_),
    .A1(_01271_),
    .A2(_01272_));
 sg13g2_a22oi_1 _06735_ (.Y(_01274_),
    .B1(_00928_),
    .B2(_00933_),
    .A2(_00853_),
    .A1(_00827_));
 sg13g2_nand2_1 _06736_ (.Y(_01275_),
    .A(_01236_),
    .B(_01174_));
 sg13g2_a221oi_1 _06737_ (.B2(_01036_),
    .C1(_01275_),
    .B1(_01274_),
    .A1(_00854_),
    .Y(_01276_),
    .A2(_01194_));
 sg13g2_a22oi_1 _06738_ (.Y(_01277_),
    .B1(_01273_),
    .B2(_01276_),
    .A2(_01270_),
    .A1(_01264_));
 sg13g2_a21oi_1 _06739_ (.A1(_01254_),
    .A2(_01263_),
    .Y(_01278_),
    .B1(net187));
 sg13g2_and4_1 _06740_ (.A(net187),
    .B(_01266_),
    .C(_01268_),
    .D(_01269_),
    .X(_01279_));
 sg13g2_a21o_1 _06741_ (.A2(_01278_),
    .A1(_01270_),
    .B1(_01279_),
    .X(_01280_));
 sg13g2_a22oi_1 _06742_ (.Y(_01281_),
    .B1(_01280_),
    .B2(_01192_),
    .A2(_01277_),
    .A1(_01253_));
 sg13g2_buf_1 _06743_ (.A(_01281_),
    .X(\i_tinyqv.cpu.i_core.cmp_out ));
 sg13g2_xnor2_1 _06744_ (.Y(_01282_),
    .A(net278),
    .B(\i_tinyqv.cpu.i_core.cmp_out ));
 sg13g2_nor2_1 _06745_ (.A(net186),
    .B(_01234_),
    .Y(_01283_));
 sg13g2_inv_1 _06746_ (.Y(_01284_),
    .A(_01283_));
 sg13g2_nor2_1 _06747_ (.A(_00894_),
    .B(\i_tinyqv.cpu.is_alu_imm ),
    .Y(_01285_));
 sg13g2_buf_1 _06748_ (.A(_01214_),
    .X(_01286_));
 sg13g2_nor2_1 _06749_ (.A(_00820_),
    .B(_01222_),
    .Y(_01287_));
 sg13g2_xnor2_1 _06750_ (.Y(_01288_),
    .A(net277),
    .B(_01287_));
 sg13g2_nor2b_1 _06751_ (.A(_00098_),
    .B_N(_01203_),
    .Y(_01289_));
 sg13g2_nand3_1 _06752_ (.B(_01285_),
    .C(_01289_),
    .A(\i_tinyqv.cpu.i_core.load_done ),
    .Y(_01290_));
 sg13g2_o21ai_1 _06753_ (.B1(_01290_),
    .Y(_01291_),
    .A1(_01285_),
    .A2(_01288_));
 sg13g2_and2_1 _06754_ (.A(net279),
    .B(_01291_),
    .X(_01292_));
 sg13g2_nor3_1 _06755_ (.A(net203),
    .B(_01284_),
    .C(_01292_),
    .Y(_01293_));
 sg13g2_a21oi_1 _06756_ (.A1(_01235_),
    .A2(_01282_),
    .Y(_01294_),
    .B1(_01293_));
 sg13g2_nand2_1 _06757_ (.Y(_01295_),
    .A(net174),
    .B(_01294_));
 sg13g2_a21oi_1 _06758_ (.A1(_00089_),
    .A2(_01208_),
    .Y(_00031_),
    .B1(_01295_));
 sg13g2_buf_1 _06759_ (.A(\i_tinyqv.mem.q_ctrl.data_req ),
    .X(_01296_));
 sg13g2_inv_1 _06760_ (.Y(_01297_),
    .A(_01296_));
 sg13g2_buf_1 _06761_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .X(_01298_));
 sg13g2_nor3_1 _06762_ (.A(\addr[26] ),
    .B(\addr[25] ),
    .C(\addr[27] ),
    .Y(_01299_));
 sg13g2_buf_1 _06763_ (.A(_01299_),
    .X(_01300_));
 sg13g2_buf_1 _06764_ (.A(\i_tinyqv.cpu.data_write_n[1] ),
    .X(_01301_));
 sg13g2_nand2_1 _06765_ (.Y(_01302_),
    .A(_01301_),
    .B(\i_tinyqv.cpu.data_read_n[1] ));
 sg13g2_buf_1 _06766_ (.A(_00159_),
    .X(_01303_));
 sg13g2_a21oi_1 _06767_ (.A1(net276),
    .A2(_01302_),
    .Y(_01304_),
    .B1(_01303_));
 sg13g2_nand2_2 _06768_ (.Y(_01305_),
    .A(net276),
    .B(_01302_));
 sg13g2_buf_1 _06769_ (.A(\i_tinyqv.cpu.data_write_n[0] ),
    .X(_01306_));
 sg13g2_nand2_1 _06770_ (.Y(_01307_),
    .A(_01306_),
    .B(\i_tinyqv.cpu.data_read_n[0] ));
 sg13g2_xor2_1 _06771_ (.B(_01307_),
    .A(_01303_),
    .X(_01308_));
 sg13g2_nor3_1 _06772_ (.A(net322),
    .B(_01305_),
    .C(_01308_),
    .Y(_01309_));
 sg13g2_a21oi_1 _06773_ (.A1(net322),
    .A2(_01304_),
    .Y(_01310_),
    .B1(_01309_));
 sg13g2_nor2_1 _06774_ (.A(_01297_),
    .B(_01310_),
    .Y(_00084_));
 sg13g2_mux2_1 _06775_ (.A0(\i_uart_tx.txd_reg ),
    .A1(\gpio_out[0] ),
    .S(\gpio_out_sel[0] ),
    .X(net28));
 sg13g2_buf_1 _06776_ (.A(debug_register_data),
    .X(_01311_));
 sg13g2_nor2b_1 _06777_ (.A(net321),
    .B_N(\i_spi.spi_select ),
    .Y(_01312_));
 sg13g2_a21oi_1 _06778_ (.A1(\debug_rd_r[2] ),
    .A2(net321),
    .Y(_01313_),
    .B1(_01312_));
 sg13g2_nand2_1 _06779_ (.Y(_01314_),
    .A(\gpio_out_sel[4] ),
    .B(\gpio_out[4] ));
 sg13g2_o21ai_1 _06780_ (.B1(_01314_),
    .Y(net32),
    .A1(\gpio_out_sel[4] ),
    .A2(_01313_));
 sg13g2_mux2_1 _06781_ (.A0(\i_uart_rx.uart_rts ),
    .A1(\gpio_out[1] ),
    .S(\gpio_out_sel[1] ),
    .X(net29));
 sg13g2_inv_1 _06782_ (.Y(_01315_),
    .A(\i_spi.spi_clk_out ));
 sg13g2_nor2_1 _06783_ (.A(_01315_),
    .B(net321),
    .Y(_01316_));
 sg13g2_a21oi_1 _06784_ (.A1(net321),
    .A2(\debug_rd_r[3] ),
    .Y(_01317_),
    .B1(_01316_));
 sg13g2_nand2_1 _06785_ (.Y(_01318_),
    .A(\gpio_out_sel[5] ),
    .B(\gpio_out[5] ));
 sg13g2_o21ai_1 _06786_ (.B1(_01318_),
    .Y(net33),
    .A1(\gpio_out_sel[5] ),
    .A2(_01317_));
 sg13g2_nor2b_1 _06787_ (.A(net321),
    .B_N(\i_spi.spi_dc ),
    .Y(_01319_));
 sg13g2_a21oi_1 _06788_ (.A1(net321),
    .A2(\debug_rd_r[0] ),
    .Y(_01320_),
    .B1(_01319_));
 sg13g2_nand2_1 _06789_ (.Y(_01321_),
    .A(\gpio_out_sel[2] ),
    .B(\gpio_out[2] ));
 sg13g2_o21ai_1 _06790_ (.B1(_01321_),
    .Y(net30),
    .A1(\gpio_out_sel[2] ),
    .A2(_01320_));
 sg13g2_mux2_1 _06791_ (.A0(debug_uart_txd),
    .A1(\gpio_out[6] ),
    .S(\gpio_out_sel[6] ),
    .X(net34));
 sg13g2_nor2b_1 _06792_ (.A(_01311_),
    .B_N(\i_spi.data[7] ),
    .Y(_01322_));
 sg13g2_a21oi_1 _06793_ (.A1(net321),
    .A2(\debug_rd_r[1] ),
    .Y(_01323_),
    .B1(_01322_));
 sg13g2_nand2_1 _06794_ (.Y(_01324_),
    .A(\gpio_out_sel[3] ),
    .B(\gpio_out[3] ));
 sg13g2_o21ai_1 _06795_ (.B1(_01324_),
    .Y(net31),
    .A1(\gpio_out_sel[3] ),
    .A2(_01323_));
 sg13g2_a21o_1 _06796_ (.A2(_01282_),
    .A1(_01235_),
    .B1(_01293_),
    .X(_01325_));
 sg13g2_buf_2 _06797_ (.A(_01325_),
    .X(_01326_));
 sg13g2_buf_1 _06798_ (.A(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .X(_01327_));
 sg13g2_nor3_2 _06799_ (.A(_01327_),
    .B(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .C(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .Y(_01328_));
 sg13g2_and3_1 _06800_ (.X(_01329_),
    .A(_01212_),
    .B(_01207_),
    .C(_01328_));
 sg13g2_buf_1 _06801_ (.A(_01329_),
    .X(_01330_));
 sg13g2_inv_1 _06802_ (.Y(_01331_),
    .A(_01330_));
 sg13g2_buf_1 _06803_ (.A(ui_in[3]),
    .X(_01332_));
 sg13g2_o21ai_1 _06804_ (.B1(net341),
    .Y(_01333_),
    .A1(_01326_),
    .A2(_01331_));
 sg13g2_inv_1 _06805_ (.Y(_01334_),
    .A(_01332_));
 sg13g2_buf_1 _06806_ (.A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .X(_01335_));
 sg13g2_buf_1 _06807_ (.A(\i_tinyqv.mem.instr_active ),
    .X(_01336_));
 sg13g2_buf_1 _06808_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .X(_01337_));
 sg13g2_nor2b_1 _06809_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B_N(net318),
    .Y(_01338_));
 sg13g2_buf_1 _06810_ (.A(_01338_),
    .X(_01339_));
 sg13g2_nand3_1 _06811_ (.B(_01336_),
    .C(_01339_),
    .A(net319),
    .Y(_01340_));
 sg13g2_buf_1 _06812_ (.A(_01340_),
    .X(_01341_));
 sg13g2_nand2_1 _06813_ (.Y(_01342_),
    .A(net320),
    .B(_01341_));
 sg13g2_buf_1 _06814_ (.A(net5),
    .X(_01343_));
 sg13g2_buf_1 _06815_ (.A(ui_in[5]),
    .X(_01344_));
 sg13g2_nand2_1 _06816_ (.Y(_01345_),
    .A(net340),
    .B(_01344_));
 sg13g2_a21oi_1 _06817_ (.A1(_01333_),
    .A2(_01342_),
    .Y(_01346_),
    .B1(_01345_));
 sg13g2_a21o_1 _06818_ (.A2(_01301_),
    .A1(_01306_),
    .B1(net276),
    .X(_01347_));
 sg13g2_buf_1 _06819_ (.A(_01347_),
    .X(_01348_));
 sg13g2_or3_1 _06820_ (.A(\addr[26] ),
    .B(\addr[25] ),
    .C(\addr[27] ),
    .X(_01349_));
 sg13g2_buf_2 _06821_ (.A(_01349_),
    .X(_01350_));
 sg13g2_nand2_1 _06822_ (.Y(_01351_),
    .A(\i_tinyqv.cpu.data_read_n[0] ),
    .B(\i_tinyqv.cpu.data_read_n[1] ));
 sg13g2_a21oi_1 _06823_ (.A1(_01350_),
    .A2(_01351_),
    .Y(_01352_),
    .B1(_01334_));
 sg13g2_a21oi_1 _06824_ (.A1(_01334_),
    .A2(_01348_),
    .Y(_01353_),
    .B1(_01352_));
 sg13g2_nand2b_1 _06825_ (.Y(_01354_),
    .B(net319),
    .A_N(_01310_));
 sg13g2_buf_2 _06826_ (.A(_00085_),
    .X(_01355_));
 sg13g2_inv_1 _06827_ (.Y(_01356_),
    .A(_01355_));
 sg13g2_a21oi_1 _06828_ (.A1(_00156_),
    .A2(_01354_),
    .Y(_01357_),
    .B1(_01356_));
 sg13g2_buf_1 _06829_ (.A(_01357_),
    .X(_01358_));
 sg13g2_nand2b_1 _06830_ (.Y(_01359_),
    .B(net276),
    .A_N(net162));
 sg13g2_buf_1 _06831_ (.A(_01359_),
    .X(_01360_));
 sg13g2_buf_1 _06832_ (.A(\i_tinyqv.cpu.i_core.mip[17] ),
    .X(_01361_));
 sg13g2_nand2_1 _06833_ (.Y(_01362_),
    .A(\i_tinyqv.cpu.i_core.mie[17] ),
    .B(_01361_));
 sg13g2_buf_1 _06834_ (.A(\i_tinyqv.cpu.i_core.mip[16] ),
    .X(_01363_));
 sg13g2_nand2_1 _06835_ (.Y(_01364_),
    .A(\i_tinyqv.cpu.i_core.mie[16] ),
    .B(_01363_));
 sg13g2_nand2_1 _06836_ (.Y(_01365_),
    .A(_01362_),
    .B(_01364_));
 sg13g2_buf_1 _06837_ (.A(\i_uart_rx.fsm_state[0] ),
    .X(_01366_));
 sg13g2_inv_1 _06838_ (.Y(_01367_),
    .A(net317));
 sg13g2_buf_2 _06839_ (.A(\i_uart_rx.fsm_state[2] ),
    .X(_01368_));
 sg13g2_buf_1 _06840_ (.A(\i_uart_rx.fsm_state[1] ),
    .X(_01369_));
 sg13g2_buf_1 _06841_ (.A(\i_uart_rx.fsm_state[3] ),
    .X(_01370_));
 sg13g2_nand2_1 _06842_ (.Y(_01371_),
    .A(net316),
    .B(net315));
 sg13g2_nor2_1 _06843_ (.A(_01368_),
    .B(_01371_),
    .Y(_01372_));
 sg13g2_inv_1 _06844_ (.Y(_01373_),
    .A(_01372_));
 sg13g2_nor2_2 _06845_ (.A(_01367_),
    .B(_01373_),
    .Y(_01374_));
 sg13g2_buf_2 _06846_ (.A(\i_uart_tx.fsm_state[1] ),
    .X(_01375_));
 sg13g2_buf_2 _06847_ (.A(\i_uart_tx.fsm_state[2] ),
    .X(_01376_));
 sg13g2_nor2_2 _06848_ (.A(_01375_),
    .B(_01376_),
    .Y(_01377_));
 sg13g2_buf_2 _06849_ (.A(\i_uart_tx.fsm_state[0] ),
    .X(_01378_));
 sg13g2_buf_2 _06850_ (.A(\i_uart_tx.fsm_state[3] ),
    .X(_01379_));
 sg13g2_nor2_1 _06851_ (.A(_01378_),
    .B(_01379_),
    .Y(_01380_));
 sg13g2_and2_1 _06852_ (.A(_01377_),
    .B(_01380_),
    .X(_01381_));
 sg13g2_buf_2 _06853_ (.A(_01381_),
    .X(_01382_));
 sg13g2_a22oi_1 _06854_ (.Y(_01383_),
    .B1(_01382_),
    .B2(\i_tinyqv.cpu.i_core.mie[19] ),
    .A2(_01374_),
    .A1(\i_tinyqv.cpu.i_core.mie[18] ));
 sg13g2_inv_1 _06855_ (.Y(_01384_),
    .A(_01383_));
 sg13g2_buf_1 _06856_ (.A(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .X(_01385_));
 sg13g2_o21ai_1 _06857_ (.B1(_01385_),
    .Y(_01386_),
    .A1(_01365_),
    .A2(_01384_));
 sg13g2_nor2_1 _06858_ (.A(net341),
    .B(_01386_),
    .Y(_01387_));
 sg13g2_a21oi_1 _06859_ (.A1(net341),
    .A2(_01360_),
    .Y(_01388_),
    .B1(_01387_));
 sg13g2_nor2_1 _06860_ (.A(net340),
    .B(_01388_),
    .Y(_01389_));
 sg13g2_a21oi_1 _06861_ (.A1(_01343_),
    .A2(_01353_),
    .Y(_01390_),
    .B1(_01389_));
 sg13g2_nand2b_1 _06862_ (.Y(_01391_),
    .B(_01390_),
    .A_N(_01344_));
 sg13g2_buf_1 _06863_ (.A(\gpio_out_sel[7] ),
    .X(_01392_));
 sg13g2_buf_1 _06864_ (.A(\gpio_out_sel[8] ),
    .X(_01393_));
 sg13g2_nor2_1 _06865_ (.A(_01392_),
    .B(_01393_),
    .Y(_01394_));
 sg13g2_nand3_1 _06866_ (.B(_01391_),
    .C(_01394_),
    .A(net6),
    .Y(_01395_));
 sg13g2_inv_1 _06867_ (.Y(_01396_),
    .A(\i_pwm.pwm_count[7] ));
 sg13g2_inv_1 _06868_ (.Y(_01397_),
    .A(\i_pwm.pwm_level[7] ));
 sg13g2_buf_1 _06869_ (.A(\i_pwm.pwm_count[6] ),
    .X(_01398_));
 sg13g2_nand2b_1 _06870_ (.Y(_01399_),
    .B(_01398_),
    .A_N(\i_pwm.pwm_level[6] ));
 sg13g2_buf_1 _06871_ (.A(\i_pwm.pwm_count[5] ),
    .X(_01400_));
 sg13g2_buf_1 _06872_ (.A(\i_pwm.pwm_count[4] ),
    .X(_01401_));
 sg13g2_inv_1 _06873_ (.Y(_01402_),
    .A(\i_pwm.pwm_level[4] ));
 sg13g2_nor2_1 _06874_ (.A(_01401_),
    .B(_01402_),
    .Y(_01403_));
 sg13g2_buf_1 _06875_ (.A(\i_pwm.pwm_count[2] ),
    .X(_01404_));
 sg13g2_inv_1 _06876_ (.Y(_01405_),
    .A(\i_pwm.pwm_level[2] ));
 sg13g2_inv_1 _06877_ (.Y(_01406_),
    .A(_01404_));
 sg13g2_buf_2 _06878_ (.A(\i_pwm.pwm_count[1] ),
    .X(_01407_));
 sg13g2_nand2b_1 _06879_ (.Y(_01408_),
    .B(_01407_),
    .A_N(\i_pwm.pwm_level[1] ));
 sg13g2_buf_1 _06880_ (.A(\i_pwm.pwm_count[0] ),
    .X(_01409_));
 sg13g2_nor2b_1 _06881_ (.A(net314),
    .B_N(\i_pwm.pwm_level[0] ),
    .Y(_01410_));
 sg13g2_nor2b_1 _06882_ (.A(_01407_),
    .B_N(\i_pwm.pwm_level[1] ),
    .Y(_01411_));
 sg13g2_a221oi_1 _06883_ (.B2(_01410_),
    .C1(_01411_),
    .B1(_01408_),
    .A1(_01406_),
    .Y(_01412_),
    .A2(\i_pwm.pwm_level[2] ));
 sg13g2_a21oi_1 _06884_ (.A1(_01404_),
    .A2(_01405_),
    .Y(_01413_),
    .B1(_01412_));
 sg13g2_nand2_1 _06885_ (.Y(_01414_),
    .A(\i_pwm.pwm_level[3] ),
    .B(_01413_));
 sg13g2_buf_1 _06886_ (.A(\i_pwm.pwm_count[3] ),
    .X(_01415_));
 sg13g2_nor2_1 _06887_ (.A(\i_pwm.pwm_level[3] ),
    .B(_01413_),
    .Y(_01416_));
 sg13g2_a221oi_1 _06888_ (.B2(_01415_),
    .C1(_01416_),
    .B1(_01414_),
    .A1(_01401_),
    .Y(_01417_),
    .A2(_01402_));
 sg13g2_or2_1 _06889_ (.X(_01418_),
    .B(_01417_),
    .A(_01403_));
 sg13g2_nor2_1 _06890_ (.A(\i_pwm.pwm_level[5] ),
    .B(_01418_),
    .Y(_01419_));
 sg13g2_nand2_1 _06891_ (.Y(_01420_),
    .A(\i_pwm.pwm_level[5] ),
    .B(_01418_));
 sg13g2_o21ai_1 _06892_ (.B1(_01420_),
    .Y(_01421_),
    .A1(_01400_),
    .A2(_01419_));
 sg13g2_nor2b_1 _06893_ (.A(_01398_),
    .B_N(\i_pwm.pwm_level[6] ),
    .Y(_01422_));
 sg13g2_a21oi_1 _06894_ (.A1(_01399_),
    .A2(_01421_),
    .Y(_01423_),
    .B1(_01422_));
 sg13g2_o21ai_1 _06895_ (.B1(_01423_),
    .Y(_01424_),
    .A1(\i_pwm.pwm_count[7] ),
    .A2(_01397_));
 sg13g2_o21ai_1 _06896_ (.B1(_01424_),
    .Y(_01425_),
    .A1(_01396_),
    .A2(\i_pwm.pwm_level[7] ));
 sg13g2_a21oi_1 _06897_ (.A1(_01392_),
    .A2(\gpio_out[7] ),
    .Y(_01426_),
    .B1(_01393_));
 sg13g2_a21o_1 _06898_ (.A2(_01425_),
    .A1(_01393_),
    .B1(_01426_),
    .X(_01427_));
 sg13g2_o21ai_1 _06899_ (.B1(_01427_),
    .Y(_01428_),
    .A1(_01346_),
    .A2(_01395_));
 sg13g2_buf_2 _06900_ (.A(\i_tinyqv.cpu.instr_len[1] ),
    .X(_01429_));
 sg13g2_nand2_1 _06901_ (.Y(_01430_),
    .A(_01067_),
    .B(_01429_));
 sg13g2_buf_2 _06902_ (.A(\i_tinyqv.cpu.instr_len[2] ),
    .X(_01431_));
 sg13g2_xor2_1 _06903_ (.B(_01431_),
    .A(_01026_),
    .X(_01432_));
 sg13g2_xnor2_1 _06904_ (.Y(_01433_),
    .A(_01430_),
    .B(_01432_));
 sg13g2_nor2_1 _06905_ (.A(_00823_),
    .B(_00102_),
    .Y(_01434_));
 sg13g2_a21oi_1 _06906_ (.A1(_00823_),
    .A2(_01433_),
    .Y(_01435_),
    .B1(_01434_));
 sg13g2_buf_1 _06907_ (.A(_01435_),
    .X(_01436_));
 sg13g2_buf_1 _06908_ (.A(net202),
    .X(_01437_));
 sg13g2_xnor2_1 _06909_ (.Y(_01438_),
    .A(_01067_),
    .B(_01429_));
 sg13g2_mux2_1 _06910_ (.A0(_00101_),
    .A1(_01438_),
    .S(_00823_),
    .X(_01439_));
 sg13g2_buf_1 _06911_ (.A(_01439_),
    .X(_01440_));
 sg13g2_buf_1 _06912_ (.A(net221),
    .X(_01441_));
 sg13g2_mux2_1 _06913_ (.A0(_00124_),
    .A1(_00125_),
    .S(net201),
    .X(_01442_));
 sg13g2_inv_1 _06914_ (.Y(_01443_),
    .A(net221));
 sg13g2_buf_1 _06915_ (.A(_01443_),
    .X(_01444_));
 sg13g2_nand2_1 _06916_ (.Y(_01445_),
    .A(_00127_),
    .B(net184));
 sg13g2_nand2_1 _06917_ (.Y(_01446_),
    .A(_00126_),
    .B(net201));
 sg13g2_a21oi_1 _06918_ (.A1(_01445_),
    .A2(_01446_),
    .Y(_01447_),
    .B1(_01436_));
 sg13g2_a21oi_1 _06919_ (.A1(net185),
    .A2(_01442_),
    .Y(_01448_),
    .B1(_01447_));
 sg13g2_buf_1 _06920_ (.A(_01448_),
    .X(_01449_));
 sg13g2_mux2_1 _06921_ (.A0(_00128_),
    .A1(_00129_),
    .S(net201),
    .X(_01450_));
 sg13g2_nand2_1 _06922_ (.Y(_01451_),
    .A(_00131_),
    .B(net184));
 sg13g2_nand2_1 _06923_ (.Y(_01452_),
    .A(_00130_),
    .B(net201));
 sg13g2_a21oi_1 _06924_ (.A1(_01451_),
    .A2(_01452_),
    .Y(_01453_),
    .B1(net185));
 sg13g2_a21o_1 _06925_ (.A2(_01450_),
    .A1(net185),
    .B1(_01453_),
    .X(_01454_));
 sg13g2_buf_1 _06926_ (.A(_01454_),
    .X(_01455_));
 sg13g2_mux2_1 _06927_ (.A0(_00120_),
    .A1(_00121_),
    .S(net201),
    .X(_01456_));
 sg13g2_nand2_1 _06928_ (.Y(_01457_),
    .A(_00123_),
    .B(net184));
 sg13g2_nand2_1 _06929_ (.Y(_01458_),
    .A(_00122_),
    .B(net201));
 sg13g2_a21oi_1 _06930_ (.A1(_01457_),
    .A2(_01458_),
    .Y(_01459_),
    .B1(net185));
 sg13g2_a21oi_1 _06931_ (.A1(net185),
    .A2(_01456_),
    .Y(_01460_),
    .B1(_01459_));
 sg13g2_buf_2 _06932_ (.A(_01460_),
    .X(_01461_));
 sg13g2_nor3_2 _06933_ (.A(net137),
    .B(_01455_),
    .C(_01461_),
    .Y(_01462_));
 sg13g2_mux2_1 _06934_ (.A0(_00116_),
    .A1(_00117_),
    .S(net221),
    .X(_01463_));
 sg13g2_nand2_1 _06935_ (.Y(_01464_),
    .A(_00119_),
    .B(_01443_));
 sg13g2_nand2_1 _06936_ (.Y(_01465_),
    .A(_00118_),
    .B(_01440_));
 sg13g2_a21oi_1 _06937_ (.A1(_01464_),
    .A2(_01465_),
    .Y(_01466_),
    .B1(net202));
 sg13g2_a21o_1 _06938_ (.A2(_01463_),
    .A1(net202),
    .B1(_01466_),
    .X(_01467_));
 sg13g2_buf_2 _06939_ (.A(_01467_),
    .X(_01468_));
 sg13g2_mux4_1 _06940_ (.S0(net201),
    .A0(_00115_),
    .A1(_00114_),
    .A2(_00112_),
    .A3(_00113_),
    .S1(net202),
    .X(_01469_));
 sg13g2_buf_2 _06941_ (.A(_01469_),
    .X(_01470_));
 sg13g2_nand2_1 _06942_ (.Y(_01471_),
    .A(_01468_),
    .B(_01470_));
 sg13g2_mux4_1 _06943_ (.S0(net221),
    .A0(\i_tinyqv.cpu.instr_data[3][3] ),
    .A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .A2(\i_tinyqv.cpu.instr_data[1][3] ),
    .A3(\i_tinyqv.cpu.instr_data[0][3] ),
    .S1(net202),
    .X(_01472_));
 sg13g2_mux2_1 _06944_ (.A0(_00108_),
    .A1(_00109_),
    .S(net221),
    .X(_01473_));
 sg13g2_mux2_1 _06945_ (.A0(_00111_),
    .A1(_00110_),
    .S(net221),
    .X(_01474_));
 sg13g2_nor2b_1 _06946_ (.A(net202),
    .B_N(_01474_),
    .Y(_01475_));
 sg13g2_a21oi_1 _06947_ (.A1(net202),
    .A2(_01473_),
    .Y(_01476_),
    .B1(_01475_));
 sg13g2_buf_1 _06948_ (.A(_01476_),
    .X(_01477_));
 sg13g2_mux4_1 _06949_ (.S0(net221),
    .A0(\i_tinyqv.cpu.instr_data[3][2] ),
    .A1(\i_tinyqv.cpu.instr_data[2][2] ),
    .A2(\i_tinyqv.cpu.instr_data[1][2] ),
    .A3(\i_tinyqv.cpu.instr_data[0][2] ),
    .S1(net202),
    .X(_01478_));
 sg13g2_buf_1 _06950_ (.A(_01478_),
    .X(_01479_));
 sg13g2_inv_2 _06951_ (.Y(_01480_),
    .A(net173));
 sg13g2_nand2b_1 _06952_ (.Y(_01481_),
    .B(_01480_),
    .A_N(net161));
 sg13g2_or2_1 _06953_ (.X(_01482_),
    .B(_01481_),
    .A(_01472_));
 sg13g2_buf_1 _06954_ (.A(_01482_),
    .X(_01483_));
 sg13g2_nor2_1 _06955_ (.A(_01471_),
    .B(_01483_),
    .Y(_01484_));
 sg13g2_mux2_1 _06956_ (.A0(_00103_),
    .A1(_00104_),
    .S(net201),
    .X(_01485_));
 sg13g2_nand2_1 _06957_ (.Y(_01486_),
    .A(_00106_),
    .B(net184));
 sg13g2_nand2_1 _06958_ (.Y(_01487_),
    .A(_00105_),
    .B(_01441_));
 sg13g2_a21oi_1 _06959_ (.A1(_01486_),
    .A2(_01487_),
    .Y(_01488_),
    .B1(_01437_));
 sg13g2_a21o_1 _06960_ (.A2(_01485_),
    .A1(net185),
    .B1(_01488_),
    .X(_01489_));
 sg13g2_buf_2 _06961_ (.A(_01489_),
    .X(_01490_));
 sg13g2_buf_1 _06962_ (.A(net221),
    .X(_01491_));
 sg13g2_mux2_1 _06963_ (.A0(\i_tinyqv.cpu.instr_data[1][0] ),
    .A1(\i_tinyqv.cpu.instr_data[0][0] ),
    .S(net200),
    .X(_01492_));
 sg13g2_nand2_1 _06964_ (.Y(_01493_),
    .A(\i_tinyqv.cpu.instr_data[3][0] ),
    .B(net184));
 sg13g2_nand2_1 _06965_ (.Y(_01494_),
    .A(\i_tinyqv.cpu.instr_data[2][0] ),
    .B(_01441_));
 sg13g2_a21oi_1 _06966_ (.A1(_01493_),
    .A2(_01494_),
    .Y(_01495_),
    .B1(_01437_));
 sg13g2_a21o_1 _06967_ (.A2(_01492_),
    .A1(net185),
    .B1(_01495_),
    .X(_01496_));
 sg13g2_buf_1 _06968_ (.A(_01496_),
    .X(_01497_));
 sg13g2_nor2_2 _06969_ (.A(_01490_),
    .B(_01497_),
    .Y(_01498_));
 sg13g2_nand3_1 _06970_ (.B(_01484_),
    .C(_01498_),
    .A(_01462_),
    .Y(_01499_));
 sg13g2_buf_1 _06971_ (.A(_01499_),
    .X(_01500_));
 sg13g2_buf_1 _06972_ (.A(net185),
    .X(_01501_));
 sg13g2_mux4_1 _06973_ (.S0(net200),
    .A0(_00147_),
    .A1(_00146_),
    .A2(_00144_),
    .A3(_00145_),
    .S1(net172),
    .X(_01502_));
 sg13g2_buf_1 _06974_ (.A(_01502_),
    .X(_01503_));
 sg13g2_mux4_1 _06975_ (.S0(_01491_),
    .A0(_00143_),
    .A1(_00142_),
    .A2(_00140_),
    .A3(_00141_),
    .S1(net172),
    .X(_01504_));
 sg13g2_buf_1 _06976_ (.A(_01504_),
    .X(_01505_));
 sg13g2_nand2_1 _06977_ (.Y(_01506_),
    .A(net147),
    .B(_01505_));
 sg13g2_buf_1 _06978_ (.A(net172),
    .X(_01507_));
 sg13g2_mux2_1 _06979_ (.A0(_00148_),
    .A1(_00149_),
    .S(net200),
    .X(_01508_));
 sg13g2_nand2_1 _06980_ (.Y(_01509_),
    .A(_00151_),
    .B(net184));
 sg13g2_nand2_1 _06981_ (.Y(_01510_),
    .A(_00150_),
    .B(net200));
 sg13g2_a21oi_1 _06982_ (.A1(_01509_),
    .A2(_01510_),
    .Y(_01511_),
    .B1(net172));
 sg13g2_a21o_1 _06983_ (.A2(_01508_),
    .A1(net160),
    .B1(_01511_),
    .X(_01512_));
 sg13g2_buf_1 _06984_ (.A(_01512_),
    .X(_01513_));
 sg13g2_mux2_1 _06985_ (.A0(_00136_),
    .A1(_00137_),
    .S(net200),
    .X(_01514_));
 sg13g2_nand2_1 _06986_ (.Y(_01515_),
    .A(_00139_),
    .B(_01444_));
 sg13g2_nand2_1 _06987_ (.Y(_01516_),
    .A(_00138_),
    .B(_01491_));
 sg13g2_a21oi_1 _06988_ (.A1(_01515_),
    .A2(_01516_),
    .Y(_01517_),
    .B1(net172));
 sg13g2_a21o_1 _06989_ (.A2(_01514_),
    .A1(net160),
    .B1(_01517_),
    .X(_01518_));
 sg13g2_buf_1 _06990_ (.A(_01518_),
    .X(_01519_));
 sg13g2_mux2_1 _06991_ (.A0(_00132_),
    .A1(_00133_),
    .S(net200),
    .X(_01520_));
 sg13g2_nand2_1 _06992_ (.Y(_01521_),
    .A(_00135_),
    .B(net184));
 sg13g2_nand2_1 _06993_ (.Y(_01522_),
    .A(_00134_),
    .B(net200));
 sg13g2_a21oi_1 _06994_ (.A1(_01521_),
    .A2(_01522_),
    .Y(_01523_),
    .B1(net172));
 sg13g2_a21oi_1 _06995_ (.A1(net160),
    .A2(_01520_),
    .Y(_01524_),
    .B1(_01523_));
 sg13g2_buf_1 _06996_ (.A(_01524_),
    .X(_01525_));
 sg13g2_nand3_1 _06997_ (.B(_01519_),
    .C(net136),
    .A(_01513_),
    .Y(_01526_));
 sg13g2_nor3_2 _06998_ (.A(_01500_),
    .B(_01506_),
    .C(_01526_),
    .Y(_01527_));
 sg13g2_a21oi_1 _06999_ (.A1(_01507_),
    .A2(_01492_),
    .Y(_01528_),
    .B1(_01495_));
 sg13g2_buf_2 _07000_ (.A(_01528_),
    .X(_01529_));
 sg13g2_a21o_1 _07001_ (.A2(_01456_),
    .A1(net172),
    .B1(_01459_),
    .X(_01530_));
 sg13g2_buf_1 _07002_ (.A(_01530_),
    .X(_01531_));
 sg13g2_nor2_2 _07003_ (.A(net137),
    .B(net135),
    .Y(_01532_));
 sg13g2_buf_1 _07004_ (.A(_01472_),
    .X(_01533_));
 sg13g2_nor4_2 _07005_ (.A(_01468_),
    .B(_01470_),
    .C(_01480_),
    .Y(_01534_),
    .D(net161));
 sg13g2_nand2_1 _07006_ (.Y(_01535_),
    .A(_01533_),
    .B(_01534_));
 sg13g2_buf_1 _07007_ (.A(_01535_),
    .X(_01536_));
 sg13g2_nor2_1 _07008_ (.A(_01490_),
    .B(_01536_),
    .Y(_01537_));
 sg13g2_a21oi_1 _07009_ (.A1(_01490_),
    .A2(_01532_),
    .Y(_01538_),
    .B1(_01537_));
 sg13g2_nor2_2 _07010_ (.A(_01529_),
    .B(_01538_),
    .Y(_01539_));
 sg13g2_or2_1 _07011_ (.X(_01540_),
    .B(_01539_),
    .A(_01527_));
 sg13g2_buf_1 _07012_ (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .X(_01541_));
 sg13g2_inv_1 _07013_ (.Y(_01542_),
    .A(_01541_));
 sg13g2_and2_1 _07014_ (.A(_00089_),
    .B(_01225_),
    .X(_01543_));
 sg13g2_buf_1 _07015_ (.A(_01543_),
    .X(_01544_));
 sg13g2_nor2b_2 _07016_ (.A(_01231_),
    .B_N(_01202_),
    .Y(_01545_));
 sg13g2_inv_1 _07017_ (.Y(_01546_),
    .A(_01110_));
 sg13g2_inv_1 _07018_ (.Y(_01547_),
    .A(_01101_));
 sg13g2_nor2_1 _07019_ (.A(_01546_),
    .B(_01547_),
    .Y(_01548_));
 sg13g2_nand4_1 _07020_ (.B(_01220_),
    .C(_01222_),
    .A(_01218_),
    .Y(_01549_),
    .D(_01548_));
 sg13g2_buf_1 _07021_ (.A(_01549_),
    .X(_01550_));
 sg13g2_nor2b_1 _07022_ (.A(_01545_),
    .B_N(_01550_),
    .Y(_01551_));
 sg13g2_or2_1 _07023_ (.X(_01552_),
    .B(_01211_),
    .A(_01209_));
 sg13g2_buf_1 _07024_ (.A(_01552_),
    .X(_01553_));
 sg13g2_a21oi_1 _07025_ (.A1(net183),
    .A2(_01551_),
    .Y(_01554_),
    .B1(_01553_));
 sg13g2_buf_1 _07026_ (.A(_01554_),
    .X(_01555_));
 sg13g2_buf_1 _07027_ (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .X(_01556_));
 sg13g2_inv_1 _07028_ (.Y(_01557_),
    .A(_01556_));
 sg13g2_nand2_1 _07029_ (.Y(_01558_),
    .A(net279),
    .B(_00893_));
 sg13g2_buf_1 _07030_ (.A(_01558_),
    .X(_01559_));
 sg13g2_nor3_1 _07031_ (.A(_01557_),
    .B(_01553_),
    .C(_01559_),
    .Y(_01560_));
 sg13g2_nor3_1 _07032_ (.A(_01556_),
    .B(_01553_),
    .C(_01559_),
    .Y(_01561_));
 sg13g2_mux2_1 _07033_ (.A0(_01560_),
    .A1(_01561_),
    .S(\i_tinyqv.cpu.i_core.cmp_out ),
    .X(_01562_));
 sg13g2_buf_1 _07034_ (.A(_01562_),
    .X(_01563_));
 sg13g2_nor3_1 _07035_ (.A(_01542_),
    .B(net146),
    .C(net86),
    .Y(_01564_));
 sg13g2_buf_1 _07036_ (.A(net279),
    .X(_01565_));
 sg13g2_nand2b_1 _07037_ (.Y(_01566_),
    .B(_01212_),
    .A_N(_01565_));
 sg13g2_o21ai_1 _07038_ (.B1(_01566_),
    .Y(_01567_),
    .A1(_01326_),
    .A2(_01331_));
 sg13g2_buf_2 _07039_ (.A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .X(_01568_));
 sg13g2_a21oi_1 _07040_ (.A1(_01067_),
    .A2(_01429_),
    .Y(_01569_),
    .B1(_01431_));
 sg13g2_nand3_1 _07041_ (.B(_01429_),
    .C(_01431_),
    .A(_01067_),
    .Y(_01570_));
 sg13g2_o21ai_1 _07042_ (.B1(_01570_),
    .Y(_01571_),
    .A1(_01027_),
    .A2(_01569_));
 sg13g2_buf_1 _07043_ (.A(_01571_),
    .X(_01572_));
 sg13g2_nor2b_1 _07044_ (.A(_00100_),
    .B_N(_01572_),
    .Y(_01573_));
 sg13g2_xnor2_1 _07045_ (.Y(_01574_),
    .A(_01568_),
    .B(_01573_));
 sg13g2_buf_1 _07046_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .X(_01575_));
 sg13g2_nand2_1 _07047_ (.Y(_01576_),
    .A(_00107_),
    .B(_01444_));
 sg13g2_nand2_1 _07048_ (.Y(_01577_),
    .A(_01501_),
    .B(_01576_));
 sg13g2_or2_1 _07049_ (.X(_01578_),
    .B(_01576_),
    .A(_01501_));
 sg13g2_nand3_1 _07050_ (.B(_01578_),
    .C(_01577_),
    .A(net313),
    .Y(_01579_));
 sg13g2_o21ai_1 _07051_ (.B1(_01579_),
    .Y(_01580_),
    .A1(net313),
    .A2(_01577_));
 sg13g2_nor4_1 _07052_ (.A(net313),
    .B(_01507_),
    .C(_01574_),
    .D(_01576_),
    .Y(_01581_));
 sg13g2_a21o_1 _07053_ (.A2(_01580_),
    .A1(_01574_),
    .B1(_01581_),
    .X(_01582_));
 sg13g2_a21oi_1 _07054_ (.A1(net172),
    .A2(_01485_),
    .Y(_01583_),
    .B1(_01488_));
 sg13g2_buf_1 _07055_ (.A(_01583_),
    .X(_01584_));
 sg13g2_nand2_1 _07056_ (.Y(_01585_),
    .A(_01584_),
    .B(_01497_));
 sg13g2_buf_2 _07057_ (.A(\i_tinyqv.cpu.instr_write_offset[1] ),
    .X(_01586_));
 sg13g2_buf_1 _07058_ (.A(net200),
    .X(_01587_));
 sg13g2_xnor2_1 _07059_ (.Y(_01588_),
    .A(_01586_),
    .B(_01587_));
 sg13g2_nand2_1 _07060_ (.Y(_01589_),
    .A(_01585_),
    .B(_01588_));
 sg13g2_buf_1 _07061_ (.A(_01553_),
    .X(_01590_));
 sg13g2_nor2_1 _07062_ (.A(net159),
    .B(_01386_),
    .Y(_01591_));
 sg13g2_inv_1 _07063_ (.Y(_01592_),
    .A(_00087_));
 sg13g2_a221oi_1 _07064_ (.B2(_01294_),
    .C1(_01592_),
    .B1(_01591_),
    .A1(_01582_),
    .Y(_01593_),
    .A2(_01589_));
 sg13g2_buf_2 _07065_ (.A(_01593_),
    .X(_01594_));
 sg13g2_nand4_1 _07066_ (.B(_01564_),
    .C(_01567_),
    .A(_01540_),
    .Y(_01595_),
    .D(_01594_));
 sg13g2_buf_2 _07067_ (.A(_01595_),
    .X(_01596_));
 sg13g2_inv_1 _07068_ (.Y(_01597_),
    .A(_00086_));
 sg13g2_nor2_1 _07069_ (.A(net146),
    .B(net86),
    .Y(_01598_));
 sg13g2_nor2_1 _07070_ (.A(_01592_),
    .B(_01598_),
    .Y(_01599_));
 sg13g2_nor3_1 _07071_ (.A(_01597_),
    .B(net341),
    .C(_01599_),
    .Y(_01600_));
 sg13g2_nand2b_1 _07072_ (.Y(_01601_),
    .B(_01344_),
    .A_N(net340));
 sg13g2_a21oi_1 _07073_ (.A1(_01565_),
    .A2(net341),
    .Y(_01602_),
    .B1(_01601_));
 sg13g2_nand2_1 _07074_ (.Y(_01603_),
    .A(_01427_),
    .B(_01602_));
 sg13g2_a21o_1 _07075_ (.A2(_01600_),
    .A1(_01596_),
    .B1(_01603_),
    .X(_01604_));
 sg13g2_nand2_1 _07076_ (.Y(_01605_),
    .A(debug_data_continue),
    .B(net320));
 sg13g2_o21ai_1 _07077_ (.B1(_01605_),
    .Y(_01606_),
    .A1(net320),
    .A2(_01146_));
 sg13g2_nand2_1 _07078_ (.Y(_01607_),
    .A(net319),
    .B(_01336_));
 sg13g2_nand3_1 _07079_ (.B(_01339_),
    .C(_01607_),
    .A(_01356_),
    .Y(_01608_));
 sg13g2_nor2_1 _07080_ (.A(_00086_),
    .B(_01341_),
    .Y(_01609_));
 sg13g2_nor2b_1 _07081_ (.A(_01609_),
    .B_N(_00107_),
    .Y(_01610_));
 sg13g2_nor3_2 _07082_ (.A(_00086_),
    .B(_00107_),
    .C(_01341_),
    .Y(_01611_));
 sg13g2_xor2_1 _07083_ (.B(_00160_),
    .A(_00102_),
    .X(_01612_));
 sg13g2_mux2_1 _07084_ (.A0(_01610_),
    .A1(_01611_),
    .S(_01612_),
    .X(_01613_));
 sg13g2_nor2_1 _07085_ (.A(_01610_),
    .B(_01611_),
    .Y(_01614_));
 sg13g2_nor2_1 _07086_ (.A(_00101_),
    .B(_01612_),
    .Y(_01615_));
 sg13g2_a22oi_1 _07087_ (.Y(_01616_),
    .B1(_01614_),
    .B2(_01615_),
    .A2(_01613_),
    .A1(_00101_));
 sg13g2_buf_1 _07088_ (.A(_01616_),
    .X(_01617_));
 sg13g2_nand2_1 _07089_ (.Y(_01618_),
    .A(_01575_),
    .B(_01611_));
 sg13g2_xor2_1 _07090_ (.B(_01618_),
    .A(_01568_),
    .X(_01619_));
 sg13g2_nor3_1 _07091_ (.A(_01608_),
    .B(_01617_),
    .C(_01619_),
    .Y(_01620_));
 sg13g2_xnor2_1 _07092_ (.Y(_01621_),
    .A(_01568_),
    .B(_01618_));
 sg13g2_nor3_1 _07093_ (.A(_01608_),
    .B(_01617_),
    .C(_01621_),
    .Y(_01622_));
 sg13g2_nand2_1 _07094_ (.Y(_01623_),
    .A(_01253_),
    .B(_01277_));
 sg13g2_a21oi_1 _07095_ (.A1(_01270_),
    .A2(_01278_),
    .Y(_01624_),
    .B1(_01279_));
 sg13g2_and4_1 _07096_ (.A(net278),
    .B(_01235_),
    .C(_01623_),
    .D(_01624_),
    .X(_01625_));
 sg13g2_nand2b_1 _07097_ (.Y(_01626_),
    .B(_01235_),
    .A_N(net278));
 sg13g2_a21oi_1 _07098_ (.A1(_01187_),
    .A2(_01191_),
    .Y(_01627_),
    .B1(_01626_));
 sg13g2_nor3_1 _07099_ (.A(net203),
    .B(_01284_),
    .C(_01292_),
    .Y(_01628_));
 sg13g2_a21oi_1 _07100_ (.A1(_01280_),
    .A2(_01627_),
    .Y(_01629_),
    .B1(_01628_));
 sg13g2_o21ai_1 _07101_ (.B1(_01629_),
    .Y(_01630_),
    .A1(_01623_),
    .A2(_01626_));
 sg13g2_nand2_1 _07102_ (.Y(_01631_),
    .A(_01330_),
    .B(_01572_));
 sg13g2_nor3_2 _07103_ (.A(_01625_),
    .B(_01630_),
    .C(_01631_),
    .Y(_01632_));
 sg13g2_mux2_1 _07104_ (.A0(_01620_),
    .A1(_01622_),
    .S(_01632_),
    .X(_01633_));
 sg13g2_buf_1 _07105_ (.A(_01633_),
    .X(_01634_));
 sg13g2_nor2_1 _07106_ (.A(net340),
    .B(net320),
    .Y(_01635_));
 sg13g2_a221oi_1 _07107_ (.B2(_01635_),
    .C1(_01344_),
    .B1(_01634_),
    .A1(net340),
    .Y(_01636_),
    .A2(_01606_));
 sg13g2_or2_1 _07108_ (.X(_01637_),
    .B(_01307_),
    .A(_01302_));
 sg13g2_nand2_2 _07109_ (.Y(_01638_),
    .A(net276),
    .B(_01637_));
 sg13g2_nor3_1 _07110_ (.A(_01617_),
    .B(_01619_),
    .C(_01638_),
    .Y(_01639_));
 sg13g2_nor3_1 _07111_ (.A(_01617_),
    .B(_01621_),
    .C(_01638_),
    .Y(_01640_));
 sg13g2_mux2_1 _07112_ (.A0(_01639_),
    .A1(_01640_),
    .S(_01632_),
    .X(_01641_));
 sg13g2_nand2_1 _07113_ (.Y(_01642_),
    .A(_01335_),
    .B(_01339_));
 sg13g2_buf_1 _07114_ (.A(_01642_),
    .X(_01643_));
 sg13g2_o21ai_1 _07115_ (.B1(_01336_),
    .Y(_01644_),
    .A1(_01643_),
    .A2(_01638_));
 sg13g2_nor2_1 _07116_ (.A(net319),
    .B(_01296_),
    .Y(_01645_));
 sg13g2_nor3_1 _07117_ (.A(debug_data_continue),
    .B(_01310_),
    .C(_01645_),
    .Y(_01646_));
 sg13g2_buf_1 _07118_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .X(_01647_));
 sg13g2_buf_1 _07119_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .X(_01648_));
 sg13g2_inv_1 _07120_ (.Y(_01649_),
    .A(_01648_));
 sg13g2_buf_1 _07121_ (.A(_00157_),
    .X(_01650_));
 sg13g2_nand2_1 _07122_ (.Y(_01651_),
    .A(net275),
    .B(net311));
 sg13g2_nor2_1 _07123_ (.A(net312),
    .B(_01651_),
    .Y(_01652_));
 sg13g2_buf_1 _07124_ (.A(_01652_),
    .X(_01653_));
 sg13g2_nand2_1 _07125_ (.Y(_01654_),
    .A(_00156_),
    .B(_01653_));
 sg13g2_o21ai_1 _07126_ (.B1(_01654_),
    .Y(_01655_),
    .A1(_01336_),
    .A2(_01646_));
 sg13g2_nor3_1 _07127_ (.A(net340),
    .B(net341),
    .C(_01655_),
    .Y(_01656_));
 sg13g2_o21ai_1 _07128_ (.B1(_01656_),
    .Y(_01657_),
    .A1(_01641_),
    .A2(_01644_));
 sg13g2_and2_1 _07129_ (.A(_01636_),
    .B(_01657_),
    .X(_01658_));
 sg13g2_nor2_2 _07130_ (.A(_01597_),
    .B(_01599_),
    .Y(_01659_));
 sg13g2_nand2b_1 _07131_ (.Y(_01660_),
    .B(\i_tinyqv.cpu.instr_fetch_started ),
    .A_N(_01634_));
 sg13g2_nand4_1 _07132_ (.B(_01596_),
    .C(_01656_),
    .A(_01659_),
    .Y(_01661_),
    .D(_01660_));
 sg13g2_and3_1 _07133_ (.X(_01662_),
    .A(_01564_),
    .B(_01567_),
    .C(_01594_));
 sg13g2_buf_1 _07134_ (.A(_01662_),
    .X(_01663_));
 sg13g2_nor2_1 _07135_ (.A(net320),
    .B(_01598_),
    .Y(_01664_));
 sg13g2_o21ai_1 _07136_ (.B1(_01344_),
    .Y(_01665_),
    .A1(net340),
    .A2(net341));
 sg13g2_a21o_1 _07137_ (.A2(_01664_),
    .A1(net340),
    .B1(_01665_),
    .X(_01666_));
 sg13g2_o21ai_1 _07138_ (.B1(net341),
    .Y(_01667_),
    .A1(net146),
    .A2(net86));
 sg13g2_a21oi_1 _07139_ (.A1(net320),
    .A2(_01539_),
    .Y(_01668_),
    .B1(_01345_));
 sg13g2_nor3_1 _07140_ (.A(\i_tinyqv.cpu.is_auipc ),
    .B(_00894_),
    .C(\i_tinyqv.cpu.is_alu_imm ),
    .Y(_01669_));
 sg13g2_nand2b_1 _07141_ (.Y(_01670_),
    .B(net279),
    .A_N(_01669_));
 sg13g2_buf_2 _07142_ (.A(_01670_),
    .X(_01671_));
 sg13g2_buf_2 _07143_ (.A(_00818_),
    .X(_01672_));
 sg13g2_nor2b_1 _07144_ (.A(net274),
    .B_N(_00817_),
    .Y(_01673_));
 sg13g2_nand2_1 _07145_ (.Y(_01674_),
    .A(_00888_),
    .B(_01673_));
 sg13g2_buf_1 _07146_ (.A(_01674_),
    .X(_01675_));
 sg13g2_nor3_1 _07147_ (.A(net222),
    .B(_01671_),
    .C(net198),
    .Y(_01676_));
 sg13g2_nand2_1 _07148_ (.Y(_01677_),
    .A(net279),
    .B(_01219_));
 sg13g2_nor2_1 _07149_ (.A(_01677_),
    .B(_01222_),
    .Y(_01678_));
 sg13g2_inv_1 _07150_ (.Y(_01679_),
    .A(_01678_));
 sg13g2_nand3_1 _07151_ (.B(\i_tinyqv.cpu.data_ready_core ),
    .C(_01289_),
    .A(net279),
    .Y(_01680_));
 sg13g2_buf_1 _07152_ (.A(_01680_),
    .X(_01681_));
 sg13g2_nand4_1 _07153_ (.B(_01671_),
    .C(_01679_),
    .A(_01233_),
    .Y(_01682_),
    .D(_01681_));
 sg13g2_nor2b_1 _07154_ (.A(_01676_),
    .B_N(_01682_),
    .Y(_01683_));
 sg13g2_buf_1 _07155_ (.A(_01683_),
    .X(_01684_));
 sg13g2_mux2_1 _07156_ (.A0(_01527_),
    .A1(_01684_),
    .S(net320),
    .X(_01685_));
 sg13g2_nor3_1 _07157_ (.A(net6),
    .B(_01392_),
    .C(_01393_),
    .Y(_01686_));
 sg13g2_o21ai_1 _07158_ (.B1(_01686_),
    .Y(_01687_),
    .A1(_01601_),
    .A2(_01685_));
 sg13g2_a21oi_1 _07159_ (.A1(_01667_),
    .A2(_01668_),
    .Y(_01688_),
    .B1(_01687_));
 sg13g2_o21ai_1 _07160_ (.B1(_01688_),
    .Y(_01689_),
    .A1(_01663_),
    .A2(_01666_));
 sg13g2_a21oi_1 _07161_ (.A1(_01658_),
    .A2(_01661_),
    .Y(_01690_),
    .B1(_01689_));
 sg13g2_a21o_1 _07162_ (.A2(_01604_),
    .A1(_01428_),
    .B1(_01690_),
    .X(net35));
 sg13g2_buf_1 _07163_ (.A(\i_debug_uart_tx.resetn ),
    .X(_01691_));
 sg13g2_buf_1 _07164_ (.A(_01691_),
    .X(_01692_));
 sg13g2_nand2_1 _07165_ (.Y(_01693_),
    .A(_01692_),
    .B(\gpio_out[0] ));
 sg13g2_buf_1 _07166_ (.A(\addr[2] ),
    .X(_01694_));
 sg13g2_buf_1 _07167_ (.A(\addr[3] ),
    .X(_01695_));
 sg13g2_nor2_2 _07168_ (.A(_01694_),
    .B(_01695_),
    .Y(_01696_));
 sg13g2_buf_1 _07169_ (.A(\addr[4] ),
    .X(_01697_));
 sg13g2_buf_2 _07170_ (.A(\addr[5] ),
    .X(_01698_));
 sg13g2_nor4_1 _07171_ (.A(\addr[16] ),
    .B(\addr[19] ),
    .C(\addr[18] ),
    .D(\addr[21] ),
    .Y(_01699_));
 sg13g2_nor4_1 _07172_ (.A(\addr[20] ),
    .B(\addr[23] ),
    .C(\addr[22] ),
    .D(\addr[24] ),
    .Y(_01700_));
 sg13g2_nor4_1 _07173_ (.A(\addr[0] ),
    .B(\addr[7] ),
    .C(\addr[6] ),
    .D(\addr[9] ),
    .Y(_01701_));
 sg13g2_inv_1 _07174_ (.Y(_01702_),
    .A(\addr[27] ));
 sg13g2_nor4_1 _07175_ (.A(_01702_),
    .B(\addr[1] ),
    .C(\addr[14] ),
    .D(\addr[17] ),
    .Y(_01703_));
 sg13g2_and4_1 _07176_ (.A(_01699_),
    .B(_01700_),
    .C(_01701_),
    .D(_01703_),
    .X(_01704_));
 sg13g2_nor4_1 _07177_ (.A(\addr[11] ),
    .B(\addr[10] ),
    .C(\addr[13] ),
    .D(\addr[15] ),
    .Y(_01705_));
 sg13g2_nor4_1 _07178_ (.A(\addr[26] ),
    .B(\addr[25] ),
    .C(\addr[8] ),
    .D(\addr[12] ),
    .Y(_01706_));
 sg13g2_nand3_1 _07179_ (.B(_01705_),
    .C(_01706_),
    .A(_01704_),
    .Y(_01707_));
 sg13g2_buf_1 _07180_ (.A(_01707_),
    .X(_01708_));
 sg13g2_nor3_1 _07181_ (.A(net310),
    .B(_01698_),
    .C(_01708_),
    .Y(_01709_));
 sg13g2_nand2_1 _07182_ (.Y(_01710_),
    .A(_01696_),
    .B(_01709_));
 sg13g2_nor2_1 _07183_ (.A(_01348_),
    .B(_01710_),
    .Y(_01711_));
 sg13g2_buf_2 _07184_ (.A(_01711_),
    .X(_01712_));
 sg13g2_buf_1 _07185_ (.A(_01712_),
    .X(_01713_));
 sg13g2_buf_1 _07186_ (.A(\data_to_write[0] ),
    .X(_01714_));
 sg13g2_nand2_1 _07187_ (.Y(_01715_),
    .A(net309),
    .B(net134));
 sg13g2_o21ai_1 _07188_ (.B1(_01715_),
    .Y(_00000_),
    .A1(_01693_),
    .A2(net134));
 sg13g2_buf_1 _07189_ (.A(_01691_),
    .X(_01716_));
 sg13g2_nand2_1 _07190_ (.Y(_01717_),
    .A(_01716_),
    .B(\gpio_out[1] ));
 sg13g2_buf_1 _07191_ (.A(\data_to_write[1] ),
    .X(_01718_));
 sg13g2_nand2_1 _07192_ (.Y(_01719_),
    .A(net308),
    .B(_01713_));
 sg13g2_o21ai_1 _07193_ (.B1(_01719_),
    .Y(_00001_),
    .A1(net134),
    .A2(_01717_));
 sg13g2_nand2_1 _07194_ (.Y(_01720_),
    .A(net231),
    .B(\gpio_out[2] ));
 sg13g2_buf_1 _07195_ (.A(\data_to_write[2] ),
    .X(_01721_));
 sg13g2_nand2_1 _07196_ (.Y(_01722_),
    .A(net307),
    .B(_01712_));
 sg13g2_o21ai_1 _07197_ (.B1(_01722_),
    .Y(_00002_),
    .A1(net134),
    .A2(_01720_));
 sg13g2_nand2_1 _07198_ (.Y(_01723_),
    .A(net231),
    .B(\gpio_out[3] ));
 sg13g2_buf_2 _07199_ (.A(\data_to_write[3] ),
    .X(_01724_));
 sg13g2_nand2_1 _07200_ (.Y(_01725_),
    .A(_01724_),
    .B(_01712_));
 sg13g2_o21ai_1 _07201_ (.B1(_01725_),
    .Y(_00003_),
    .A1(net134),
    .A2(_01723_));
 sg13g2_nand2_1 _07202_ (.Y(_01726_),
    .A(net231),
    .B(\gpio_out[4] ));
 sg13g2_buf_1 _07203_ (.A(\data_to_write[4] ),
    .X(_01727_));
 sg13g2_nand2_1 _07204_ (.Y(_01728_),
    .A(net306),
    .B(_01712_));
 sg13g2_o21ai_1 _07205_ (.B1(_01728_),
    .Y(_00004_),
    .A1(net134),
    .A2(_01726_));
 sg13g2_nand2_1 _07206_ (.Y(_01729_),
    .A(net231),
    .B(\gpio_out[5] ));
 sg13g2_buf_1 _07207_ (.A(\data_to_write[5] ),
    .X(_01730_));
 sg13g2_nand2_1 _07208_ (.Y(_01731_),
    .A(net305),
    .B(_01712_));
 sg13g2_o21ai_1 _07209_ (.B1(_01731_),
    .Y(_00005_),
    .A1(net134),
    .A2(_01729_));
 sg13g2_buf_1 _07210_ (.A(net232),
    .X(_01732_));
 sg13g2_nand2_1 _07211_ (.Y(_01733_),
    .A(net220),
    .B(\gpio_out[6] ));
 sg13g2_buf_1 _07212_ (.A(\data_to_write[6] ),
    .X(_01734_));
 sg13g2_nand2_1 _07213_ (.Y(_01735_),
    .A(net304),
    .B(_01712_));
 sg13g2_o21ai_1 _07214_ (.B1(_01735_),
    .Y(_00006_),
    .A1(_01713_),
    .A2(_01733_));
 sg13g2_nand2_1 _07215_ (.Y(_01736_),
    .A(net220),
    .B(\gpio_out[7] ));
 sg13g2_buf_2 _07216_ (.A(\data_to_write[7] ),
    .X(_01737_));
 sg13g2_nand2_1 _07217_ (.Y(_01738_),
    .A(_01737_),
    .B(_01712_));
 sg13g2_o21ai_1 _07218_ (.B1(_01738_),
    .Y(_00007_),
    .A1(net134),
    .A2(_01736_));
 sg13g2_nand2_1 _07219_ (.Y(_01739_),
    .A(_01692_),
    .B(\gpio_out_sel[0] ));
 sg13g2_nor2_1 _07220_ (.A(_01698_),
    .B(_01708_),
    .Y(_01740_));
 sg13g2_nand2b_1 _07221_ (.Y(_01741_),
    .B(_01740_),
    .A_N(net310));
 sg13g2_buf_1 _07222_ (.A(_01694_),
    .X(_01742_));
 sg13g2_buf_1 _07223_ (.A(_01695_),
    .X(_01743_));
 sg13g2_nand2_1 _07224_ (.Y(_01744_),
    .A(net273),
    .B(net272));
 sg13g2_nor3_1 _07225_ (.A(_01348_),
    .B(_01741_),
    .C(_01744_),
    .Y(_01745_));
 sg13g2_buf_1 _07226_ (.A(_01745_),
    .X(_01746_));
 sg13g2_buf_1 _07227_ (.A(net145),
    .X(_01747_));
 sg13g2_nand2_1 _07228_ (.Y(_01748_),
    .A(net309),
    .B(net145));
 sg13g2_o21ai_1 _07229_ (.B1(_01748_),
    .Y(_00008_),
    .A1(_01739_),
    .A2(net133));
 sg13g2_nand2_1 _07230_ (.Y(_01749_),
    .A(_01732_),
    .B(\gpio_out_sel[1] ));
 sg13g2_nand2_1 _07231_ (.Y(_01750_),
    .A(net308),
    .B(net145));
 sg13g2_o21ai_1 _07232_ (.B1(_01750_),
    .Y(_00009_),
    .A1(net133),
    .A2(_01749_));
 sg13g2_nand2_1 _07233_ (.Y(_01751_),
    .A(_01732_),
    .B(\gpio_out_sel[2] ));
 sg13g2_nand2_1 _07234_ (.Y(_01752_),
    .A(net307),
    .B(net145));
 sg13g2_o21ai_1 _07235_ (.B1(_01752_),
    .Y(_00010_),
    .A1(net133),
    .A2(_01751_));
 sg13g2_nand2_1 _07236_ (.Y(_01753_),
    .A(net220),
    .B(\gpio_out_sel[3] ));
 sg13g2_nand2_1 _07237_ (.Y(_01754_),
    .A(_01724_),
    .B(net145));
 sg13g2_o21ai_1 _07238_ (.B1(_01754_),
    .Y(_00011_),
    .A1(_01747_),
    .A2(_01753_));
 sg13g2_nand2_1 _07239_ (.Y(_01755_),
    .A(net220),
    .B(\gpio_out_sel[4] ));
 sg13g2_nand2_1 _07240_ (.Y(_01756_),
    .A(net306),
    .B(net145));
 sg13g2_o21ai_1 _07241_ (.B1(_01756_),
    .Y(_00012_),
    .A1(net133),
    .A2(_01755_));
 sg13g2_nand2_1 _07242_ (.Y(_01757_),
    .A(net220),
    .B(\gpio_out_sel[5] ));
 sg13g2_nand2_1 _07243_ (.Y(_01758_),
    .A(net305),
    .B(_01746_));
 sg13g2_o21ai_1 _07244_ (.B1(_01758_),
    .Y(_00013_),
    .A1(_01747_),
    .A2(_01757_));
 sg13g2_nand2_1 _07245_ (.Y(_01759_),
    .A(net220),
    .B(\gpio_out_sel[6] ));
 sg13g2_nand2_1 _07246_ (.Y(_01760_),
    .A(net304),
    .B(net145));
 sg13g2_o21ai_1 _07247_ (.B1(_01760_),
    .Y(_00014_),
    .A1(net133),
    .A2(_01759_));
 sg13g2_nand2_1 _07248_ (.Y(_01761_),
    .A(net232),
    .B(_01392_));
 sg13g2_o21ai_1 _07249_ (.B1(_01761_),
    .Y(_01762_),
    .A1(net232),
    .A2(_01343_));
 sg13g2_mux2_1 _07250_ (.A0(_01762_),
    .A1(_01737_),
    .S(net133),
    .X(_00015_));
 sg13g2_nand2_1 _07251_ (.Y(_01763_),
    .A(net220),
    .B(_01393_));
 sg13g2_nand2_1 _07252_ (.Y(_01764_),
    .A(\data_to_write[8] ),
    .B(net145));
 sg13g2_o21ai_1 _07253_ (.B1(_01764_),
    .Y(_00016_),
    .A1(net133),
    .A2(_01763_));
 sg13g2_nand2_1 _07254_ (.Y(_01765_),
    .A(net220),
    .B(\gpio_out_sel[9] ));
 sg13g2_nand2_1 _07255_ (.Y(_01766_),
    .A(\data_to_write[9] ),
    .B(_01746_));
 sg13g2_o21ai_1 _07256_ (.B1(_01766_),
    .Y(_00017_),
    .A1(net133),
    .A2(_01765_));
 sg13g2_buf_1 _07257_ (.A(_00166_),
    .X(_01767_));
 sg13g2_buf_1 _07258_ (.A(_01767_),
    .X(_01768_));
 sg13g2_inv_1 _07259_ (.Y(_01769_),
    .A(_01204_));
 sg13g2_nand2_1 _07260_ (.Y(_01770_),
    .A(_01294_),
    .B(_01330_));
 sg13g2_nand2_1 _07261_ (.Y(_01771_),
    .A(_01203_),
    .B(_01770_));
 sg13g2_buf_1 _07262_ (.A(\i_tinyqv.cpu.i_core.cycle[0] ),
    .X(_01772_));
 sg13g2_buf_1 _07263_ (.A(_01772_),
    .X(_01773_));
 sg13g2_buf_1 _07264_ (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .X(_01774_));
 sg13g2_nor2_1 _07265_ (.A(net270),
    .B(_01774_),
    .Y(_01775_));
 sg13g2_or2_1 _07266_ (.X(_01776_),
    .B(_01289_),
    .A(_01229_));
 sg13g2_nand4_1 _07267_ (.B(net174),
    .C(_01775_),
    .A(net233),
    .Y(_01777_),
    .D(_01776_));
 sg13g2_buf_1 _07268_ (.A(_01777_),
    .X(_01778_));
 sg13g2_a21o_1 _07269_ (.A2(_01771_),
    .A1(_01769_),
    .B1(_01778_),
    .X(_01779_));
 sg13g2_nor2_1 _07270_ (.A(_01328_),
    .B(_01778_),
    .Y(_01780_));
 sg13g2_a22oi_1 _07271_ (.Y(_01781_),
    .B1(_01780_),
    .B2(_01204_),
    .A2(_01779_),
    .A1(debug_data_continue));
 sg13g2_nand2_1 _07272_ (.Y(_01782_),
    .A(_01203_),
    .B(_01780_));
 sg13g2_o21ai_1 _07273_ (.B1(_01782_),
    .Y(_00030_),
    .A1(net271),
    .A2(_01781_));
 sg13g2_buf_1 _07274_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .X(_01783_));
 sg13g2_buf_1 _07275_ (.A(_01783_),
    .X(_01784_));
 sg13g2_a21oi_1 _07276_ (.A1(_01238_),
    .A2(_01240_),
    .Y(_01785_),
    .B1(net277));
 sg13g2_buf_1 _07277_ (.A(_01785_),
    .X(_01786_));
 sg13g2_nand2_1 _07278_ (.Y(_01787_),
    .A(net269),
    .B(net132));
 sg13g2_inv_1 _07279_ (.Y(_01788_),
    .A(_01787_));
 sg13g2_nand2_1 _07280_ (.Y(_01789_),
    .A(_01167_),
    .B(_01169_));
 sg13g2_nand4_1 _07281_ (.B(_01160_),
    .C(_01164_),
    .A(_01156_),
    .Y(_01790_),
    .D(_01789_));
 sg13g2_buf_2 _07282_ (.A(_01790_),
    .X(_01791_));
 sg13g2_nand3_1 _07283_ (.B(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .C(_01791_),
    .A(_01772_),
    .Y(_01792_));
 sg13g2_buf_1 _07284_ (.A(_01792_),
    .X(_01793_));
 sg13g2_buf_1 _07285_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .X(_01794_));
 sg13g2_nand2_1 _07286_ (.Y(_01795_),
    .A(_01216_),
    .B(net303));
 sg13g2_buf_2 _07287_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .X(_01796_));
 sg13g2_nand2_2 _07288_ (.Y(_01797_),
    .A(net235),
    .B(_01796_));
 sg13g2_a21oi_2 _07289_ (.B1(_01797_),
    .Y(_01798_),
    .A2(_01055_),
    .A1(_01045_));
 sg13g2_or3_1 _07290_ (.A(net163),
    .B(_01795_),
    .C(_01798_),
    .X(_01799_));
 sg13g2_o21ai_1 _07291_ (.B1(_01798_),
    .Y(_01800_),
    .A1(net163),
    .A2(_01795_));
 sg13g2_nand3_1 _07292_ (.B(_01799_),
    .C(_01800_),
    .A(_01793_),
    .Y(_01801_));
 sg13g2_a21o_1 _07293_ (.A2(_01800_),
    .A1(_01799_),
    .B1(_01793_),
    .X(_01802_));
 sg13g2_nand2_1 _07294_ (.Y(_01803_),
    .A(_01801_),
    .B(_01802_));
 sg13g2_inv_1 _07295_ (.Y(_01804_),
    .A(_01772_));
 sg13g2_inv_1 _07296_ (.Y(_01805_),
    .A(_01796_));
 sg13g2_and4_1 _07297_ (.A(_01156_),
    .B(_01160_),
    .C(_01164_),
    .D(_01789_),
    .X(_01806_));
 sg13g2_buf_1 _07298_ (.A(_01806_),
    .X(_01807_));
 sg13g2_nor3_2 _07299_ (.A(_01804_),
    .B(_01805_),
    .C(net158),
    .Y(_01808_));
 sg13g2_inv_2 _07300_ (.Y(_01809_),
    .A(_01783_));
 sg13g2_nor3_2 _07301_ (.A(net277),
    .B(_01809_),
    .C(net163),
    .Y(_01810_));
 sg13g2_a21oi_1 _07302_ (.A1(_01045_),
    .A2(_01055_),
    .Y(_01811_),
    .B1(_01795_));
 sg13g2_buf_2 _07303_ (.A(_01811_),
    .X(_01812_));
 sg13g2_o21ai_1 _07304_ (.B1(_01812_),
    .Y(_01813_),
    .A1(_01808_),
    .A2(_01810_));
 sg13g2_buf_1 _07305_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .X(_01814_));
 sg13g2_a21oi_1 _07306_ (.A1(_01808_),
    .A2(_01810_),
    .Y(_01815_),
    .B1(_01814_));
 sg13g2_and2_1 _07307_ (.A(_01814_),
    .B(_01812_),
    .X(_01816_));
 sg13g2_or2_1 _07308_ (.X(_01817_),
    .B(_01810_),
    .A(_01808_));
 sg13g2_and3_1 _07309_ (.X(_01818_),
    .A(_01814_),
    .B(_01808_),
    .C(_01810_));
 sg13g2_a221oi_1 _07310_ (.B2(_01817_),
    .C1(_01818_),
    .B1(_01816_),
    .A1(_01813_),
    .Y(_01819_),
    .A2(_01815_));
 sg13g2_xnor2_1 _07311_ (.Y(_01820_),
    .A(_01803_),
    .B(_01819_));
 sg13g2_nor2_1 _07312_ (.A(_01788_),
    .B(_01820_),
    .Y(_01821_));
 sg13g2_buf_1 _07313_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .X(_01822_));
 sg13g2_nor2_1 _07314_ (.A(_01804_),
    .B(net158),
    .Y(_01823_));
 sg13g2_buf_1 _07315_ (.A(_01823_),
    .X(_01824_));
 sg13g2_buf_1 _07316_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .X(_01825_));
 sg13g2_a21oi_1 _07317_ (.A1(_01822_),
    .A2(net131),
    .Y(_01826_),
    .B1(_01825_));
 sg13g2_a21oi_1 _07318_ (.A1(_01045_),
    .A2(_01055_),
    .Y(_01827_),
    .B1(net277));
 sg13g2_buf_8 _07319_ (.A(_01827_),
    .X(_01828_));
 sg13g2_buf_1 _07320_ (.A(net157),
    .X(_01829_));
 sg13g2_nand2b_1 _07321_ (.Y(_01830_),
    .B(net144),
    .A_N(net303));
 sg13g2_buf_1 _07322_ (.A(_01791_),
    .X(_01831_));
 sg13g2_nand2_1 _07323_ (.Y(_01832_),
    .A(net270),
    .B(_01831_));
 sg13g2_buf_2 _07324_ (.A(_01832_),
    .X(_01833_));
 sg13g2_nand3_1 _07325_ (.B(_01833_),
    .C(net144),
    .A(_01825_),
    .Y(_01834_));
 sg13g2_o21ai_1 _07326_ (.B1(_01834_),
    .Y(_01835_),
    .A1(_01826_),
    .A2(_01830_));
 sg13g2_nand2_1 _07327_ (.Y(_01836_),
    .A(net235),
    .B(_01057_));
 sg13g2_buf_1 _07328_ (.A(_01836_),
    .X(_01837_));
 sg13g2_a21oi_1 _07329_ (.A1(_01794_),
    .A2(net130),
    .Y(_01838_),
    .B1(_01825_));
 sg13g2_nand3_1 _07330_ (.B(_01822_),
    .C(net131),
    .A(net269),
    .Y(_01839_));
 sg13g2_nand2_1 _07331_ (.Y(_01840_),
    .A(net269),
    .B(net157));
 sg13g2_nand4_1 _07332_ (.B(_01825_),
    .C(net131),
    .A(net303),
    .Y(_01841_),
    .D(_01840_));
 sg13g2_o21ai_1 _07333_ (.B1(_01841_),
    .Y(_01842_),
    .A1(_01838_),
    .A2(_01839_));
 sg13g2_a21oi_1 _07334_ (.A1(net269),
    .A2(_01835_),
    .Y(_01843_),
    .B1(_01842_));
 sg13g2_nand2_1 _07335_ (.Y(_01844_),
    .A(net303),
    .B(net157));
 sg13g2_nand3_1 _07336_ (.B(_01796_),
    .C(_01791_),
    .A(net270),
    .Y(_01845_));
 sg13g2_buf_8 _07337_ (.A(_01196_),
    .X(_01846_));
 sg13g2_a22oi_1 _07338_ (.Y(_01847_),
    .B1(net143),
    .B2(net270),
    .A2(net142),
    .A1(net222));
 sg13g2_a21o_1 _07339_ (.A2(_01845_),
    .A1(_01809_),
    .B1(_01847_),
    .X(_01848_));
 sg13g2_nor2_1 _07340_ (.A(_01783_),
    .B(_01805_),
    .Y(_01849_));
 sg13g2_nand2_1 _07341_ (.Y(_01850_),
    .A(_01812_),
    .B(_01849_));
 sg13g2_nor2_1 _07342_ (.A(_01809_),
    .B(_01796_),
    .Y(_01851_));
 sg13g2_o21ai_1 _07343_ (.B1(_01851_),
    .Y(_01852_),
    .A1(net277),
    .A2(net163));
 sg13g2_nor2_1 _07344_ (.A(_01809_),
    .B(_01805_),
    .Y(_01853_));
 sg13g2_nand3_1 _07345_ (.B(net142),
    .C(_01853_),
    .A(net222),
    .Y(_01854_));
 sg13g2_nand3_1 _07346_ (.B(_01852_),
    .C(_01854_),
    .A(_01850_),
    .Y(_01855_));
 sg13g2_nand2_1 _07347_ (.Y(_01856_),
    .A(net235),
    .B(net142));
 sg13g2_buf_2 _07348_ (.A(_01856_),
    .X(_01857_));
 sg13g2_nand2_1 _07349_ (.Y(_01858_),
    .A(_01784_),
    .B(_01812_));
 sg13g2_nor3_1 _07350_ (.A(net131),
    .B(_01857_),
    .C(_01858_),
    .Y(_01859_));
 sg13g2_a221oi_1 _07351_ (.B2(net131),
    .C1(_01859_),
    .B1(_01855_),
    .A1(_01844_),
    .Y(_01860_),
    .A2(_01848_));
 sg13g2_xnor2_1 _07352_ (.Y(_01861_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .B(_01860_));
 sg13g2_or2_1 _07353_ (.X(_01862_),
    .B(_01861_),
    .A(_01843_));
 sg13g2_buf_2 _07354_ (.A(_01862_),
    .X(_01863_));
 sg13g2_nand2_1 _07355_ (.Y(_01864_),
    .A(_01788_),
    .B(_01820_));
 sg13g2_nand2_1 _07356_ (.Y(_01865_),
    .A(_01863_),
    .B(_01864_));
 sg13g2_nand2b_1 _07357_ (.Y(_01866_),
    .B(_01865_),
    .A_N(_01821_));
 sg13g2_nor2_1 _07358_ (.A(net277),
    .B(net163),
    .Y(_01867_));
 sg13g2_buf_1 _07359_ (.A(_01867_),
    .X(_01868_));
 sg13g2_xnor2_1 _07360_ (.Y(_01869_),
    .A(_01796_),
    .B(net129));
 sg13g2_nor2_1 _07361_ (.A(_01833_),
    .B(_01858_),
    .Y(_01870_));
 sg13g2_nand3_1 _07362_ (.B(_01812_),
    .C(_01845_),
    .A(_01809_),
    .Y(_01871_));
 sg13g2_nand4_1 _07363_ (.B(_01833_),
    .C(net129),
    .A(_01784_),
    .Y(_01872_),
    .D(_01844_));
 sg13g2_nand3_1 _07364_ (.B(_01857_),
    .C(_01812_),
    .A(net269),
    .Y(_01873_));
 sg13g2_nand3_1 _07365_ (.B(_01872_),
    .C(_01873_),
    .A(_01871_),
    .Y(_01874_));
 sg13g2_nand2b_1 _07366_ (.Y(_01875_),
    .B(_01849_),
    .A_N(_01812_));
 sg13g2_o21ai_1 _07367_ (.B1(_01853_),
    .Y(_01876_),
    .A1(net277),
    .A2(_01014_));
 sg13g2_buf_8 _07368_ (.A(net142),
    .X(_01877_));
 sg13g2_nand3_1 _07369_ (.B(net128),
    .C(_01851_),
    .A(net222),
    .Y(_01878_));
 sg13g2_nand3_1 _07370_ (.B(_01876_),
    .C(_01878_),
    .A(_01875_),
    .Y(_01879_));
 sg13g2_inv_1 _07371_ (.Y(_01880_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[2] ));
 sg13g2_nor2_1 _07372_ (.A(_01880_),
    .B(_01833_),
    .Y(_01881_));
 sg13g2_and2_1 _07373_ (.A(_01879_),
    .B(_01881_),
    .X(_01882_));
 sg13g2_a221oi_1 _07374_ (.B2(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .C1(_01882_),
    .B1(_01874_),
    .A1(_01869_),
    .Y(_01883_),
    .A2(_01870_));
 sg13g2_buf_1 _07375_ (.A(_01883_),
    .X(_01884_));
 sg13g2_nor3_1 _07376_ (.A(_01884_),
    .B(_01863_),
    .C(_01864_),
    .Y(_01885_));
 sg13g2_a221oi_1 _07377_ (.B2(_01884_),
    .C1(_01885_),
    .B1(_01866_),
    .A1(_01821_),
    .Y(_01886_),
    .A2(_01863_));
 sg13g2_a21oi_1 _07378_ (.A1(_01812_),
    .A2(_01808_),
    .Y(_01887_),
    .B1(_01810_));
 sg13g2_a21o_1 _07379_ (.A2(_01845_),
    .A1(_01844_),
    .B1(_01887_),
    .X(_01888_));
 sg13g2_nand3_1 _07380_ (.B(_01801_),
    .C(_01802_),
    .A(_01814_),
    .Y(_01889_));
 sg13g2_a21oi_1 _07381_ (.A1(_01801_),
    .A2(_01802_),
    .Y(_01890_),
    .B1(_01814_));
 sg13g2_a21o_1 _07382_ (.A2(_01889_),
    .A1(_01888_),
    .B1(_01890_),
    .X(_01891_));
 sg13g2_nor2_1 _07383_ (.A(_00799_),
    .B(_00816_),
    .Y(_01892_));
 sg13g2_buf_1 _07384_ (.A(_01892_),
    .X(_01893_));
 sg13g2_nor2_1 _07385_ (.A(_01893_),
    .B(_01795_),
    .Y(_01894_));
 sg13g2_nor2_1 _07386_ (.A(net277),
    .B(_01805_),
    .Y(_01895_));
 sg13g2_nand2_1 _07387_ (.Y(_01896_),
    .A(net142),
    .B(_01895_));
 sg13g2_buf_1 _07388_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .X(_01897_));
 sg13g2_and2_1 _07389_ (.A(_01772_),
    .B(net302),
    .X(_01898_));
 sg13g2_buf_1 _07390_ (.A(_01898_),
    .X(_01899_));
 sg13g2_nand2_1 _07391_ (.Y(_01900_),
    .A(net235),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[3] ));
 sg13g2_a21o_1 _07392_ (.A2(_01055_),
    .A1(_01045_),
    .B1(_01900_),
    .X(_01901_));
 sg13g2_buf_2 _07393_ (.A(_01901_),
    .X(_01902_));
 sg13g2_a21o_1 _07394_ (.A2(_01899_),
    .A1(_01791_),
    .B1(_01902_),
    .X(_01903_));
 sg13g2_buf_1 _07395_ (.A(_01903_),
    .X(_01904_));
 sg13g2_nand3_1 _07396_ (.B(_01899_),
    .C(_01902_),
    .A(_01791_),
    .Y(_01905_));
 sg13g2_buf_1 _07397_ (.A(_01905_),
    .X(_01906_));
 sg13g2_nand3_1 _07398_ (.B(_01904_),
    .C(_01906_),
    .A(_01896_),
    .Y(_01907_));
 sg13g2_a21oi_1 _07399_ (.A1(_01791_),
    .A2(_01899_),
    .Y(_01908_),
    .B1(_01902_));
 sg13g2_and3_1 _07400_ (.X(_01909_),
    .A(_01791_),
    .B(_01899_),
    .C(_01902_));
 sg13g2_buf_1 _07401_ (.A(_01909_),
    .X(_01910_));
 sg13g2_nor2_2 _07402_ (.A(net163),
    .B(_01797_),
    .Y(_01911_));
 sg13g2_o21ai_1 _07403_ (.B1(_01911_),
    .Y(_01912_),
    .A1(_01908_),
    .A2(_01910_));
 sg13g2_and2_1 _07404_ (.A(_01907_),
    .B(_01912_),
    .X(_01913_));
 sg13g2_buf_1 _07405_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .X(_01914_));
 sg13g2_nor2b_1 _07406_ (.A(_01286_),
    .B_N(net303),
    .Y(_01915_));
 sg13g2_nand3_1 _07407_ (.B(_01915_),
    .C(_01798_),
    .A(net142),
    .Y(_01916_));
 sg13g2_a21oi_1 _07408_ (.A1(net142),
    .A2(_01915_),
    .Y(_01917_),
    .B1(_01798_));
 sg13g2_a21oi_2 _07409_ (.B1(_01917_),
    .Y(_01918_),
    .A2(_01916_),
    .A1(_01793_));
 sg13g2_xnor2_1 _07410_ (.Y(_01919_),
    .A(_01914_),
    .B(_01918_));
 sg13g2_xnor2_1 _07411_ (.Y(_01920_),
    .A(_01913_),
    .B(_01919_));
 sg13g2_xor2_1 _07412_ (.B(_01920_),
    .A(_01894_),
    .X(_01921_));
 sg13g2_xnor2_1 _07413_ (.Y(_01922_),
    .A(_01891_),
    .B(_01921_));
 sg13g2_xor2_1 _07414_ (.B(_01922_),
    .A(_01886_),
    .X(_00018_));
 sg13g2_nand2b_1 _07415_ (.Y(_01923_),
    .B(_01891_),
    .A_N(_01921_));
 sg13g2_inv_1 _07416_ (.Y(_01924_),
    .A(_01820_));
 sg13g2_a21oi_1 _07417_ (.A1(_01888_),
    .A2(_01889_),
    .Y(_01925_),
    .B1(_01890_));
 sg13g2_a221oi_1 _07418_ (.B2(_01921_),
    .C1(_01863_),
    .B1(_01925_),
    .A1(_01787_),
    .Y(_01926_),
    .A2(_01924_));
 sg13g2_nand2_1 _07419_ (.Y(_01927_),
    .A(_01923_),
    .B(_01926_));
 sg13g2_or3_1 _07420_ (.A(_01884_),
    .B(_01843_),
    .C(_01861_),
    .X(_01928_));
 sg13g2_nor2_1 _07421_ (.A(_01864_),
    .B(_01928_),
    .Y(_01929_));
 sg13g2_and3_1 _07422_ (.X(_01930_),
    .A(_01871_),
    .B(_01872_),
    .C(_01873_));
 sg13g2_a22oi_1 _07423_ (.Y(_01931_),
    .B1(_01879_),
    .B2(_01881_),
    .A2(_01870_),
    .A1(_01869_));
 sg13g2_o21ai_1 _07424_ (.B1(_01931_),
    .Y(_01932_),
    .A1(_01880_),
    .A2(_01930_));
 sg13g2_o21ai_1 _07425_ (.B1(_01932_),
    .Y(_01933_),
    .A1(_01788_),
    .A2(_01820_));
 sg13g2_nand3_1 _07426_ (.B(_01928_),
    .C(_01933_),
    .A(_01864_),
    .Y(_01934_));
 sg13g2_o21ai_1 _07427_ (.B1(_01934_),
    .Y(_01935_),
    .A1(_01929_),
    .A2(_01922_));
 sg13g2_and2_1 _07428_ (.A(_01927_),
    .B(_01935_),
    .X(_01936_));
 sg13g2_buf_1 _07429_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .X(_01937_));
 sg13g2_and2_1 _07430_ (.A(_01772_),
    .B(_01937_),
    .X(_01938_));
 sg13g2_buf_1 _07431_ (.A(_01938_),
    .X(_01939_));
 sg13g2_nand2_1 _07432_ (.Y(_01940_),
    .A(net143),
    .B(_01939_));
 sg13g2_nor2b_1 _07433_ (.A(_01214_),
    .B_N(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .Y(_01941_));
 sg13g2_buf_2 _07434_ (.A(_01941_),
    .X(_01942_));
 sg13g2_nand2_1 _07435_ (.Y(_01943_),
    .A(net235),
    .B(net302));
 sg13g2_a21o_1 _07436_ (.A2(_01055_),
    .A1(_01045_),
    .B1(_01943_),
    .X(_01944_));
 sg13g2_buf_1 _07437_ (.A(_01944_),
    .X(_01945_));
 sg13g2_nand3_1 _07438_ (.B(_01942_),
    .C(_01945_),
    .A(_01196_),
    .Y(_01946_));
 sg13g2_buf_1 _07439_ (.A(_01946_),
    .X(_01947_));
 sg13g2_a21o_1 _07440_ (.A2(_01942_),
    .A1(_01196_),
    .B1(_01945_),
    .X(_01948_));
 sg13g2_buf_1 _07441_ (.A(_01948_),
    .X(_01949_));
 sg13g2_nand2_2 _07442_ (.Y(_01950_),
    .A(_01947_),
    .B(_01949_));
 sg13g2_xnor2_1 _07443_ (.Y(_01951_),
    .A(_01940_),
    .B(_01950_));
 sg13g2_inv_1 _07444_ (.Y(_01952_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ));
 sg13g2_nand2_1 _07445_ (.Y(_01953_),
    .A(_01772_),
    .B(net302));
 sg13g2_o21ai_1 _07446_ (.B1(_01902_),
    .Y(_01954_),
    .A1(net158),
    .A2(_01953_));
 sg13g2_nor3_1 _07447_ (.A(net158),
    .B(_01953_),
    .C(_01902_),
    .Y(_01955_));
 sg13g2_a21oi_2 _07448_ (.B1(_01955_),
    .Y(_01956_),
    .A2(_01954_),
    .A1(_01911_));
 sg13g2_xnor2_1 _07449_ (.Y(_01957_),
    .A(_01952_),
    .B(_01956_));
 sg13g2_xnor2_1 _07450_ (.Y(_01958_),
    .A(_01951_),
    .B(_01957_));
 sg13g2_a21oi_1 _07451_ (.A1(_01238_),
    .A2(_01240_),
    .Y(_01959_),
    .B1(_01797_));
 sg13g2_buf_1 _07452_ (.A(_01959_),
    .X(_01960_));
 sg13g2_nand4_1 _07453_ (.B(_01904_),
    .C(_01906_),
    .A(_01896_),
    .Y(_01961_),
    .D(net127));
 sg13g2_and2_1 _07454_ (.A(_01000_),
    .B(_01012_),
    .X(_01962_));
 sg13g2_a221oi_1 _07455_ (.B2(_01962_),
    .C1(_01797_),
    .B1(_00991_),
    .A1(_01238_),
    .Y(_01963_),
    .A2(_01240_));
 sg13g2_o21ai_1 _07456_ (.B1(_01963_),
    .Y(_01964_),
    .A1(_01908_),
    .A2(_01910_));
 sg13g2_a21oi_1 _07457_ (.A1(_01961_),
    .A2(_01964_),
    .Y(_01965_),
    .B1(_01918_));
 sg13g2_inv_1 _07458_ (.Y(_01966_),
    .A(_01914_));
 sg13g2_and2_1 _07459_ (.A(_01966_),
    .B(net127),
    .X(_01967_));
 sg13g2_nand2_2 _07460_ (.Y(_01968_),
    .A(_01238_),
    .B(_01240_));
 sg13g2_a221oi_1 _07461_ (.B2(_01906_),
    .C1(_01911_),
    .B1(_01904_),
    .A1(_01968_),
    .Y(_01969_),
    .A2(_01895_));
 sg13g2_mux2_1 _07462_ (.A0(_01967_),
    .A1(_01969_),
    .S(_01918_),
    .X(_01970_));
 sg13g2_or4_1 _07463_ (.A(_01896_),
    .B(_01908_),
    .C(_01910_),
    .D(net127),
    .X(_01971_));
 sg13g2_nand2b_1 _07464_ (.Y(_01972_),
    .B(_01914_),
    .A_N(_01960_));
 sg13g2_a21o_1 _07465_ (.A2(_01916_),
    .A1(_01793_),
    .B1(_01917_),
    .X(_01973_));
 sg13g2_a21oi_1 _07466_ (.A1(_01971_),
    .A2(_01972_),
    .Y(_01974_),
    .B1(_01973_));
 sg13g2_and2_1 _07467_ (.A(_01896_),
    .B(net127),
    .X(_01975_));
 sg13g2_nor2_1 _07468_ (.A(_01896_),
    .B(net127),
    .Y(_01976_));
 sg13g2_nor2_1 _07469_ (.A(_01911_),
    .B(net127),
    .Y(_01977_));
 sg13g2_nand2_1 _07470_ (.Y(_01978_),
    .A(_01904_),
    .B(_01906_));
 sg13g2_mux4_1 _07471_ (.S0(_01978_),
    .A0(_01975_),
    .A1(_01963_),
    .A2(_01976_),
    .A3(_01977_),
    .S1(_01914_),
    .X(_01979_));
 sg13g2_nor4_1 _07472_ (.A(_01965_),
    .B(_01970_),
    .C(_01974_),
    .D(_01979_),
    .Y(_01980_));
 sg13g2_xnor2_1 _07473_ (.Y(_01981_),
    .A(_01958_),
    .B(_01980_));
 sg13g2_o21ai_1 _07474_ (.B1(_01925_),
    .Y(_01982_),
    .A1(_01894_),
    .A2(_01920_));
 sg13g2_nand2_1 _07475_ (.Y(_01983_),
    .A(_01894_),
    .B(_01920_));
 sg13g2_nand2_1 _07476_ (.Y(_01984_),
    .A(_01982_),
    .B(_01983_));
 sg13g2_nand2_1 _07477_ (.Y(_01985_),
    .A(_01981_),
    .B(_01984_));
 sg13g2_nand3b_1 _07478_ (.B(_01982_),
    .C(_01983_),
    .Y(_01986_),
    .A_N(_01981_));
 sg13g2_and2_1 _07479_ (.A(_01985_),
    .B(_01986_),
    .X(_01987_));
 sg13g2_xnor2_1 _07480_ (.Y(_00021_),
    .A(_01936_),
    .B(_01987_));
 sg13g2_nor2_1 _07481_ (.A(_01981_),
    .B(_01984_),
    .Y(_01988_));
 sg13g2_o21ai_1 _07482_ (.B1(_01985_),
    .Y(_01989_),
    .A1(_01936_),
    .A2(_01988_));
 sg13g2_nand2_1 _07483_ (.Y(_01990_),
    .A(_01958_),
    .B(net127));
 sg13g2_nand3_1 _07484_ (.B(_01907_),
    .C(_01912_),
    .A(_01918_),
    .Y(_01991_));
 sg13g2_a21oi_1 _07485_ (.A1(_01907_),
    .A2(_01912_),
    .Y(_01992_),
    .B1(_01918_));
 sg13g2_a21oi_1 _07486_ (.A1(_01966_),
    .A2(_01991_),
    .Y(_01993_),
    .B1(_01992_));
 sg13g2_o21ai_1 _07487_ (.B1(_01993_),
    .Y(_01994_),
    .A1(_01958_),
    .A2(net127));
 sg13g2_and2_1 _07488_ (.A(_01990_),
    .B(_01994_),
    .X(_01995_));
 sg13g2_buf_2 _07489_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .X(_01996_));
 sg13g2_inv_1 _07490_ (.Y(_01997_),
    .A(_01996_));
 sg13g2_nor3_2 _07491_ (.A(_01804_),
    .B(_01997_),
    .C(_01807_),
    .Y(_01998_));
 sg13g2_nand3_1 _07492_ (.B(net302),
    .C(net128),
    .A(net222),
    .Y(_01999_));
 sg13g2_and2_1 _07493_ (.A(_01937_),
    .B(net157),
    .X(_02000_));
 sg13g2_buf_1 _07494_ (.A(_02000_),
    .X(_02001_));
 sg13g2_xnor2_1 _07495_ (.Y(_02002_),
    .A(_01999_),
    .B(_02001_));
 sg13g2_xnor2_1 _07496_ (.Y(_02003_),
    .A(_01998_),
    .B(_02002_));
 sg13g2_a22oi_1 _07497_ (.Y(_02004_),
    .B1(_01939_),
    .B2(net143),
    .A2(_01942_),
    .A1(net128));
 sg13g2_nand4_1 _07498_ (.B(net143),
    .C(_01942_),
    .A(net128),
    .Y(_02005_),
    .D(_01939_));
 sg13g2_o21ai_1 _07499_ (.B1(_02005_),
    .Y(_02006_),
    .A1(_01945_),
    .A2(_02004_));
 sg13g2_xor2_1 _07500_ (.B(_02006_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .X(_02007_));
 sg13g2_xor2_1 _07501_ (.B(_02007_),
    .A(_02003_),
    .X(_02008_));
 sg13g2_a221oi_1 _07502_ (.B2(_01949_),
    .C1(_01940_),
    .B1(_01947_),
    .A1(_01968_),
    .Y(_02009_),
    .A2(_01942_));
 sg13g2_and2_1 _07503_ (.A(net143),
    .B(_01939_),
    .X(_02010_));
 sg13g2_buf_1 _07504_ (.A(_02010_),
    .X(_02011_));
 sg13g2_and3_1 _07505_ (.X(_02012_),
    .A(net128),
    .B(_01942_),
    .C(_01945_));
 sg13g2_a21oi_1 _07506_ (.A1(net128),
    .A2(_01942_),
    .Y(_02013_),
    .B1(_01945_));
 sg13g2_a21oi_1 _07507_ (.A1(_01238_),
    .A2(_01240_),
    .Y(_02014_),
    .B1(_01900_));
 sg13g2_nor4_1 _07508_ (.A(_02011_),
    .B(_02012_),
    .C(_02013_),
    .D(_02014_),
    .Y(_02015_));
 sg13g2_o21ai_1 _07509_ (.B1(_01956_),
    .Y(_02016_),
    .A1(_02009_),
    .A2(_02015_));
 sg13g2_o21ai_1 _07510_ (.B1(_01942_),
    .Y(_02017_),
    .A1(_00799_),
    .A2(_00816_));
 sg13g2_buf_1 _07511_ (.A(_02017_),
    .X(_02018_));
 sg13g2_nand3_1 _07512_ (.B(_01956_),
    .C(_02018_),
    .A(_01952_),
    .Y(_02019_));
 sg13g2_nand4_1 _07513_ (.B(_02011_),
    .C(_01950_),
    .A(_01952_),
    .Y(_02020_),
    .D(_02018_));
 sg13g2_or4_1 _07514_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .B(_02011_),
    .C(_01950_),
    .D(_02014_),
    .X(_02021_));
 sg13g2_and4_1 _07515_ (.A(_02016_),
    .B(_02019_),
    .C(_02020_),
    .D(_02021_),
    .X(_02022_));
 sg13g2_buf_1 _07516_ (.A(_02022_),
    .X(_02023_));
 sg13g2_a221oi_1 _07517_ (.B2(_01939_),
    .C1(_01900_),
    .B1(net143),
    .A1(_01238_),
    .Y(_02024_),
    .A2(_01240_));
 sg13g2_o21ai_1 _07518_ (.B1(_02024_),
    .Y(_02025_),
    .A1(_02012_),
    .A2(_02013_));
 sg13g2_nand4_1 _07519_ (.B(_01947_),
    .C(_01949_),
    .A(_02011_),
    .Y(_02026_),
    .D(_02014_));
 sg13g2_a21oi_1 _07520_ (.A1(_02025_),
    .A2(_02026_),
    .Y(_02027_),
    .B1(_01956_));
 sg13g2_nor3_1 _07521_ (.A(_01952_),
    .B(_01956_),
    .C(_02018_),
    .Y(_02028_));
 sg13g2_nor3_1 _07522_ (.A(_01952_),
    .B(_01940_),
    .C(_02018_),
    .Y(_02029_));
 sg13g2_and2_1 _07523_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .B(_02024_),
    .X(_02030_));
 sg13g2_mux2_1 _07524_ (.A0(_02029_),
    .A1(_02030_),
    .S(_01950_),
    .X(_02031_));
 sg13g2_nor3_1 _07525_ (.A(_02027_),
    .B(_02028_),
    .C(_02031_),
    .Y(_02032_));
 sg13g2_nand3_1 _07526_ (.B(_02023_),
    .C(_02032_),
    .A(_02008_),
    .Y(_02033_));
 sg13g2_a21o_1 _07527_ (.A2(_02032_),
    .A1(_02023_),
    .B1(_02008_),
    .X(_02034_));
 sg13g2_nand2_1 _07528_ (.Y(_02035_),
    .A(_02033_),
    .B(_02034_));
 sg13g2_xnor2_1 _07529_ (.Y(_02036_),
    .A(_01995_),
    .B(_02035_));
 sg13g2_xor2_1 _07530_ (.B(_02036_),
    .A(_01989_),
    .X(_00022_));
 sg13g2_a22oi_1 _07531_ (.Y(_02037_),
    .B1(_02033_),
    .B2(_02034_),
    .A2(_01994_),
    .A1(_01990_));
 sg13g2_a221oi_1 _07532_ (.B2(_01984_),
    .C1(_02037_),
    .B1(_01981_),
    .A1(_01923_),
    .Y(_02038_),
    .A2(_01926_));
 sg13g2_nand4_1 _07533_ (.B(_01994_),
    .C(_02033_),
    .A(_01990_),
    .Y(_02039_),
    .D(_02034_));
 sg13g2_o21ai_1 _07534_ (.B1(_02039_),
    .Y(_02040_),
    .A1(_01986_),
    .A2(_02037_));
 sg13g2_a21oi_2 _07535_ (.B1(_02040_),
    .Y(_02041_),
    .A2(_02038_),
    .A1(_01935_));
 sg13g2_xnor2_1 _07536_ (.Y(_02042_),
    .A(_02003_),
    .B(_02007_));
 sg13g2_or3_1 _07537_ (.A(_02027_),
    .B(_02028_),
    .C(_02031_),
    .X(_02043_));
 sg13g2_a21oi_1 _07538_ (.A1(_02042_),
    .A2(_02023_),
    .Y(_02044_),
    .B1(_02043_));
 sg13g2_buf_2 _07539_ (.A(_02044_),
    .X(_02045_));
 sg13g2_a22oi_1 _07540_ (.Y(_02046_),
    .B1(_01998_),
    .B2(_02001_),
    .A2(net129),
    .A1(net302));
 sg13g2_nor2_1 _07541_ (.A(_01998_),
    .B(_02001_),
    .Y(_02047_));
 sg13g2_nor2_1 _07542_ (.A(_02046_),
    .B(_02047_),
    .Y(_02048_));
 sg13g2_buf_1 _07543_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[7] ),
    .X(_02049_));
 sg13g2_buf_1 _07544_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .X(_02050_));
 sg13g2_nand3_1 _07545_ (.B(net300),
    .C(_01791_),
    .A(_01772_),
    .Y(_02051_));
 sg13g2_buf_1 _07546_ (.A(_02051_),
    .X(_02052_));
 sg13g2_and2_1 _07547_ (.A(net301),
    .B(net126),
    .X(_02053_));
 sg13g2_nor2_1 _07548_ (.A(net301),
    .B(net126),
    .Y(_02054_));
 sg13g2_nand2_2 _07549_ (.Y(_02055_),
    .A(_01996_),
    .B(net157));
 sg13g2_nand3_1 _07550_ (.B(_01937_),
    .C(_01196_),
    .A(net235),
    .Y(_02056_));
 sg13g2_buf_1 _07551_ (.A(_02056_),
    .X(_02057_));
 sg13g2_xor2_1 _07552_ (.B(_02057_),
    .A(_02055_),
    .X(_02058_));
 sg13g2_buf_1 _07553_ (.A(_02058_),
    .X(_02059_));
 sg13g2_o21ai_1 _07554_ (.B1(_02059_),
    .Y(_02060_),
    .A1(_02053_),
    .A2(_02054_));
 sg13g2_inv_1 _07555_ (.Y(_02061_),
    .A(net301));
 sg13g2_and2_1 _07556_ (.A(_02061_),
    .B(net126),
    .X(_02062_));
 sg13g2_nor2_1 _07557_ (.A(_02061_),
    .B(net126),
    .Y(_02063_));
 sg13g2_xnor2_1 _07558_ (.Y(_02064_),
    .A(_02055_),
    .B(_02057_));
 sg13g2_o21ai_1 _07559_ (.B1(_02064_),
    .Y(_02065_),
    .A1(_02062_),
    .A2(_02063_));
 sg13g2_and3_1 _07560_ (.X(_02066_),
    .A(_02048_),
    .B(_02060_),
    .C(_02065_));
 sg13g2_buf_1 _07561_ (.A(_02066_),
    .X(_02067_));
 sg13g2_a21oi_1 _07562_ (.A1(_02060_),
    .A2(_02065_),
    .Y(_02068_),
    .B1(_02048_));
 sg13g2_or2_1 _07563_ (.X(_02069_),
    .B(_02068_),
    .A(_02067_));
 sg13g2_nand2_1 _07564_ (.Y(_02070_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .B(_02006_));
 sg13g2_nor2_1 _07565_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .B(_02006_),
    .Y(_02071_));
 sg13g2_a21oi_2 _07566_ (.B1(_02071_),
    .Y(_02072_),
    .A2(_02070_),
    .A1(_02003_));
 sg13g2_nand2_1 _07567_ (.Y(_02073_),
    .A(net302),
    .B(net132));
 sg13g2_xor2_1 _07568_ (.B(_02073_),
    .A(_02072_),
    .X(_02074_));
 sg13g2_xnor2_1 _07569_ (.Y(_02075_),
    .A(_02069_),
    .B(_02074_));
 sg13g2_xnor2_1 _07570_ (.Y(_02076_),
    .A(_02045_),
    .B(_02075_));
 sg13g2_xnor2_1 _07571_ (.Y(_00023_),
    .A(_02041_),
    .B(_02076_));
 sg13g2_nor2_1 _07572_ (.A(_02055_),
    .B(_02052_),
    .Y(_02077_));
 sg13g2_a21oi_1 _07573_ (.A1(_02055_),
    .A2(_02052_),
    .Y(_02078_),
    .B1(_02057_));
 sg13g2_nor2_1 _07574_ (.A(_02077_),
    .B(_02078_),
    .Y(_02079_));
 sg13g2_nand3_1 _07575_ (.B(_01996_),
    .C(net142),
    .A(net222),
    .Y(_02080_));
 sg13g2_nand2_1 _07576_ (.Y(_02081_),
    .A(net300),
    .B(_01828_));
 sg13g2_xnor2_1 _07577_ (.Y(_02082_),
    .A(_02080_),
    .B(_02081_));
 sg13g2_buf_2 _07578_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .X(_02083_));
 sg13g2_nand3_1 _07579_ (.B(_02083_),
    .C(net143),
    .A(_01773_),
    .Y(_02084_));
 sg13g2_buf_1 _07580_ (.A(_02084_),
    .X(_02085_));
 sg13g2_xnor2_1 _07581_ (.Y(_02086_),
    .A(_02082_),
    .B(_02085_));
 sg13g2_xnor2_1 _07582_ (.Y(_02087_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .B(_02086_));
 sg13g2_xnor2_1 _07583_ (.Y(_02088_),
    .A(_02079_),
    .B(_02087_));
 sg13g2_nand2_1 _07584_ (.Y(_02089_),
    .A(_01937_),
    .B(net132));
 sg13g2_buf_1 _07585_ (.A(_02089_),
    .X(_02090_));
 sg13g2_nand3_1 _07586_ (.B(net126),
    .C(net101),
    .A(_02059_),
    .Y(_02091_));
 sg13g2_and2_1 _07587_ (.A(net300),
    .B(net131),
    .X(_02092_));
 sg13g2_buf_1 _07588_ (.A(_02092_),
    .X(_02093_));
 sg13g2_nand3_1 _07589_ (.B(_02093_),
    .C(net101),
    .A(_02064_),
    .Y(_02094_));
 sg13g2_or2_1 _07590_ (.X(_02095_),
    .B(_02047_),
    .A(_02046_));
 sg13g2_buf_1 _07591_ (.A(_02095_),
    .X(_02096_));
 sg13g2_a21o_1 _07592_ (.A2(_02094_),
    .A1(_02091_),
    .B1(_02096_),
    .X(_02097_));
 sg13g2_and3_1 _07593_ (.X(_02098_),
    .A(net301),
    .B(net126),
    .C(_02089_));
 sg13g2_and2_1 _07594_ (.A(net301),
    .B(net101),
    .X(_02099_));
 sg13g2_and4_1 _07595_ (.A(net301),
    .B(_02064_),
    .C(_02093_),
    .D(_02090_),
    .X(_02100_));
 sg13g2_a221oi_1 _07596_ (.B2(_02048_),
    .C1(_02100_),
    .B1(_02099_),
    .A1(_02059_),
    .Y(_02101_),
    .A2(_02098_));
 sg13g2_nor3_1 _07597_ (.A(_02064_),
    .B(net126),
    .C(net101),
    .Y(_02102_));
 sg13g2_nor3_1 _07598_ (.A(_02059_),
    .B(_02093_),
    .C(net101),
    .Y(_02103_));
 sg13g2_o21ai_1 _07599_ (.B1(_02096_),
    .Y(_02104_),
    .A1(_02102_),
    .A2(_02103_));
 sg13g2_nor3_1 _07600_ (.A(net301),
    .B(net126),
    .C(net101),
    .Y(_02105_));
 sg13g2_nor2_1 _07601_ (.A(_02049_),
    .B(net101),
    .Y(_02106_));
 sg13g2_nor4_1 _07602_ (.A(net301),
    .B(_02059_),
    .C(_02093_),
    .D(net101),
    .Y(_02107_));
 sg13g2_a221oi_1 _07603_ (.B2(_02096_),
    .C1(_02107_),
    .B1(_02106_),
    .A1(_02059_),
    .Y(_02108_),
    .A2(_02105_));
 sg13g2_nand4_1 _07604_ (.B(_02101_),
    .C(_02104_),
    .A(_02097_),
    .Y(_02109_),
    .D(_02108_));
 sg13g2_xnor2_1 _07605_ (.Y(_02110_),
    .A(_02088_),
    .B(_02109_));
 sg13g2_o21ai_1 _07606_ (.B1(_02073_),
    .Y(_02111_),
    .A1(_02067_),
    .A2(_02068_));
 sg13g2_nor2_1 _07607_ (.A(_02072_),
    .B(_02111_),
    .Y(_02112_));
 sg13g2_nor3_2 _07608_ (.A(_02067_),
    .B(_02068_),
    .C(_02073_),
    .Y(_02113_));
 sg13g2_a21oi_2 _07609_ (.B1(_02113_),
    .Y(_02114_),
    .A2(_02111_),
    .A1(_02072_));
 sg13g2_a21oi_1 _07610_ (.A1(_02045_),
    .A2(_02114_),
    .Y(_02115_),
    .B1(_02112_));
 sg13g2_nand2b_1 _07611_ (.Y(_02116_),
    .B(_02115_),
    .A_N(_02041_));
 sg13g2_nand2_1 _07612_ (.Y(_02117_),
    .A(_02072_),
    .B(_02113_));
 sg13g2_o21ai_1 _07613_ (.B1(_02117_),
    .Y(_02118_),
    .A1(_02045_),
    .A2(_02114_));
 sg13g2_nand2b_1 _07614_ (.Y(_02119_),
    .B(_02041_),
    .A_N(_02118_));
 sg13g2_nor2_1 _07615_ (.A(_02045_),
    .B(_02117_),
    .Y(_02120_));
 sg13g2_a221oi_1 _07616_ (.B2(_02119_),
    .C1(_02120_),
    .B1(_02116_),
    .A1(_02045_),
    .Y(_02121_),
    .A2(_02112_));
 sg13g2_xnor2_1 _07617_ (.Y(_00024_),
    .A(_02110_),
    .B(_02121_));
 sg13g2_a22oi_1 _07618_ (.Y(_02122_),
    .B1(_02110_),
    .B2(_02114_),
    .A2(_02075_),
    .A1(_02045_));
 sg13g2_nand2b_1 _07619_ (.Y(_02123_),
    .B(_02111_),
    .A_N(_02045_));
 sg13g2_a21oi_1 _07620_ (.A1(_02114_),
    .A2(_02123_),
    .Y(_02124_),
    .B1(_02110_));
 sg13g2_xor2_1 _07621_ (.B(_02109_),
    .A(_02088_),
    .X(_02125_));
 sg13g2_nor2b_1 _07622_ (.A(_02045_),
    .B_N(_02072_),
    .Y(_02126_));
 sg13g2_o21ai_1 _07623_ (.B1(_02126_),
    .Y(_02127_),
    .A1(_02125_),
    .A2(_02113_));
 sg13g2_nand2b_1 _07624_ (.Y(_02128_),
    .B(_02127_),
    .A_N(_02124_));
 sg13g2_a21oi_1 _07625_ (.A1(_02041_),
    .A2(_02122_),
    .Y(_02129_),
    .B1(_02128_));
 sg13g2_nor2_1 _07626_ (.A(_02081_),
    .B(_02085_),
    .Y(_02130_));
 sg13g2_a21oi_2 _07627_ (.B1(_02080_),
    .Y(_02131_),
    .A2(_02085_),
    .A1(_02081_));
 sg13g2_or2_1 _07628_ (.X(_02132_),
    .B(_02131_),
    .A(_02130_));
 sg13g2_nand3_1 _07629_ (.B(net300),
    .C(_01846_),
    .A(net222),
    .Y(_02133_));
 sg13g2_and2_1 _07630_ (.A(_02083_),
    .B(_01827_),
    .X(_02134_));
 sg13g2_buf_1 _07631_ (.A(_02134_),
    .X(_02135_));
 sg13g2_xnor2_1 _07632_ (.Y(_02136_),
    .A(_02133_),
    .B(_02135_));
 sg13g2_buf_2 _07633_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .X(_02137_));
 sg13g2_inv_1 _07634_ (.Y(_02138_),
    .A(_02137_));
 sg13g2_nor3_2 _07635_ (.A(_01804_),
    .B(_02138_),
    .C(_01807_),
    .Y(_02139_));
 sg13g2_xnor2_1 _07636_ (.Y(_02140_),
    .A(_02136_),
    .B(_02139_));
 sg13g2_xor2_1 _07637_ (.B(_02140_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .X(_02141_));
 sg13g2_xnor2_1 _07638_ (.Y(_02142_),
    .A(_02132_),
    .B(_02141_));
 sg13g2_o21ai_1 _07639_ (.B1(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .Y(_02143_),
    .A1(_02077_),
    .A2(_02078_));
 sg13g2_nor3_1 _07640_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .B(_02077_),
    .C(_02078_),
    .Y(_02144_));
 sg13g2_a21oi_2 _07641_ (.B1(_02144_),
    .Y(_02145_),
    .A2(_02143_),
    .A1(_02086_));
 sg13g2_nand2_1 _07642_ (.Y(_02146_),
    .A(_01996_),
    .B(net132));
 sg13g2_xor2_1 _07643_ (.B(_02146_),
    .A(_02145_),
    .X(_02147_));
 sg13g2_xnor2_1 _07644_ (.Y(_02148_),
    .A(_02142_),
    .B(_02147_));
 sg13g2_inv_1 _07645_ (.Y(_02149_),
    .A(_02090_));
 sg13g2_nand2_1 _07646_ (.Y(_02150_),
    .A(_02088_),
    .B(_02149_));
 sg13g2_xnor2_1 _07647_ (.Y(_02151_),
    .A(_02064_),
    .B(_02093_));
 sg13g2_inv_1 _07648_ (.Y(_02152_),
    .A(_02151_));
 sg13g2_o21ai_1 _07649_ (.B1(_02049_),
    .Y(_02153_),
    .A1(_02048_),
    .A2(_02151_));
 sg13g2_o21ai_1 _07650_ (.B1(_02153_),
    .Y(_02154_),
    .A1(_02096_),
    .A2(_02152_));
 sg13g2_o21ai_1 _07651_ (.B1(_02154_),
    .Y(_02155_),
    .A1(_02088_),
    .A2(_02149_));
 sg13g2_nand3b_1 _07652_ (.B(_02150_),
    .C(_02155_),
    .Y(_02156_),
    .A_N(_02148_));
 sg13g2_nand2_1 _07653_ (.Y(_02157_),
    .A(_02150_),
    .B(_02155_));
 sg13g2_nand2_1 _07654_ (.Y(_02158_),
    .A(_02148_),
    .B(_02157_));
 sg13g2_and2_1 _07655_ (.A(_02156_),
    .B(_02158_),
    .X(_02159_));
 sg13g2_xnor2_1 _07656_ (.Y(_00025_),
    .A(_02129_),
    .B(_02159_));
 sg13g2_nor2_1 _07657_ (.A(_02148_),
    .B(_02157_),
    .Y(_02160_));
 sg13g2_a21oi_2 _07658_ (.B1(_02160_),
    .Y(_02161_),
    .A2(_02158_),
    .A1(_02129_));
 sg13g2_nor2_1 _07659_ (.A(_02135_),
    .B(_02139_),
    .Y(_02162_));
 sg13g2_a22oi_1 _07660_ (.Y(_02163_),
    .B1(_02135_),
    .B2(_02139_),
    .A2(net129),
    .A1(net300));
 sg13g2_or2_1 _07661_ (.X(_02164_),
    .B(_02163_),
    .A(_02162_));
 sg13g2_buf_1 _07662_ (.A(_02164_),
    .X(_02165_));
 sg13g2_buf_1 _07663_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .X(_02166_));
 sg13g2_inv_1 _07664_ (.Y(_02167_),
    .A(_02166_));
 sg13g2_buf_2 _07665_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .X(_02168_));
 sg13g2_nand3_1 _07666_ (.B(_02168_),
    .C(net143),
    .A(_01773_),
    .Y(_02169_));
 sg13g2_buf_2 _07667_ (.A(_02169_),
    .X(_02170_));
 sg13g2_nand2_2 _07668_ (.Y(_02171_),
    .A(_02137_),
    .B(net157));
 sg13g2_nand3_1 _07669_ (.B(_02083_),
    .C(_01196_),
    .A(net235),
    .Y(_02172_));
 sg13g2_buf_1 _07670_ (.A(_02172_),
    .X(_02173_));
 sg13g2_xnor2_1 _07671_ (.Y(_02174_),
    .A(_02171_),
    .B(_02173_));
 sg13g2_xnor2_1 _07672_ (.Y(_02175_),
    .A(_02170_),
    .B(_02174_));
 sg13g2_xnor2_1 _07673_ (.Y(_02176_),
    .A(_02167_),
    .B(_02175_));
 sg13g2_xnor2_1 _07674_ (.Y(_02177_),
    .A(_02165_),
    .B(_02176_));
 sg13g2_o21ai_1 _07675_ (.B1(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .Y(_02178_),
    .A1(_02130_),
    .A2(_02131_));
 sg13g2_nor3_1 _07676_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .B(_02130_),
    .C(_02131_),
    .Y(_02179_));
 sg13g2_a21oi_2 _07677_ (.B1(_02179_),
    .Y(_02180_),
    .A2(_02178_),
    .A1(_02140_));
 sg13g2_nand2_1 _07678_ (.Y(_02181_),
    .A(net300),
    .B(net132));
 sg13g2_xor2_1 _07679_ (.B(_02181_),
    .A(_02180_),
    .X(_02182_));
 sg13g2_xnor2_1 _07680_ (.Y(_02183_),
    .A(_02177_),
    .B(_02182_));
 sg13g2_nand3_1 _07681_ (.B(net132),
    .C(_02145_),
    .A(_01996_),
    .Y(_02184_));
 sg13g2_nor2_1 _07682_ (.A(_02130_),
    .B(_02131_),
    .Y(_02185_));
 sg13g2_nand3b_1 _07683_ (.B(_02145_),
    .C(_02185_),
    .Y(_02186_),
    .A_N(_02141_));
 sg13g2_nand3_1 _07684_ (.B(_02132_),
    .C(_02141_),
    .A(_02145_),
    .Y(_02187_));
 sg13g2_nand2b_1 _07685_ (.Y(_02188_),
    .B(_02185_),
    .A_N(_02146_));
 sg13g2_or2_1 _07686_ (.X(_02189_),
    .B(_02146_),
    .A(_02185_));
 sg13g2_mux2_1 _07687_ (.A0(_02188_),
    .A1(_02189_),
    .S(_02141_),
    .X(_02190_));
 sg13g2_and4_1 _07688_ (.A(_02184_),
    .B(_02186_),
    .C(_02187_),
    .D(_02190_),
    .X(_02191_));
 sg13g2_xnor2_1 _07689_ (.Y(_02192_),
    .A(_02183_),
    .B(_02191_));
 sg13g2_xnor2_1 _07690_ (.Y(_00026_),
    .A(_02161_),
    .B(_02192_));
 sg13g2_nand4_1 _07691_ (.B(_02186_),
    .C(_02187_),
    .A(_02184_),
    .Y(_02193_),
    .D(_02190_));
 sg13g2_nand2_1 _07692_ (.Y(_02194_),
    .A(_02161_),
    .B(_02193_));
 sg13g2_nor2_1 _07693_ (.A(_02161_),
    .B(_02193_),
    .Y(_02195_));
 sg13g2_a21oi_1 _07694_ (.A1(_02183_),
    .A2(_02194_),
    .Y(_02196_),
    .B1(_02195_));
 sg13g2_nand3_1 _07695_ (.B(net132),
    .C(_02180_),
    .A(net300),
    .Y(_02197_));
 sg13g2_nor2b_1 _07696_ (.A(_02180_),
    .B_N(_02181_),
    .Y(_02198_));
 sg13g2_a21o_1 _07697_ (.A2(_02197_),
    .A1(_02177_),
    .B1(_02198_),
    .X(_02199_));
 sg13g2_buf_1 _07698_ (.A(_02199_),
    .X(_02200_));
 sg13g2_nand2_1 _07699_ (.Y(_02201_),
    .A(_02170_),
    .B(_02171_));
 sg13g2_o21ai_1 _07700_ (.B1(_02173_),
    .Y(_02202_),
    .A1(_02170_),
    .A2(_02171_));
 sg13g2_nand2_1 _07701_ (.Y(_02203_),
    .A(_02201_),
    .B(_02202_));
 sg13g2_buf_1 _07702_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .X(_02204_));
 sg13g2_nand2_1 _07703_ (.Y(_02205_),
    .A(_02204_),
    .B(net131));
 sg13g2_nand2_1 _07704_ (.Y(_02206_),
    .A(_02168_),
    .B(net157));
 sg13g2_nand3_1 _07705_ (.B(_02137_),
    .C(_01846_),
    .A(_01216_),
    .Y(_02207_));
 sg13g2_xnor2_1 _07706_ (.Y(_02208_),
    .A(_02206_),
    .B(_02207_));
 sg13g2_xnor2_1 _07707_ (.Y(_02209_),
    .A(_02205_),
    .B(_02208_));
 sg13g2_xor2_1 _07708_ (.B(_02209_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .X(_02210_));
 sg13g2_xnor2_1 _07709_ (.Y(_02211_),
    .A(_02203_),
    .B(_02210_));
 sg13g2_and2_1 _07710_ (.A(_02083_),
    .B(_01785_),
    .X(_02212_));
 sg13g2_buf_1 _07711_ (.A(_02212_),
    .X(_02213_));
 sg13g2_nor3_1 _07712_ (.A(_02170_),
    .B(_02174_),
    .C(_02213_),
    .Y(_02214_));
 sg13g2_inv_1 _07713_ (.Y(_02215_),
    .A(_02168_));
 sg13g2_nor2_1 _07714_ (.A(_02215_),
    .B(_01833_),
    .Y(_02216_));
 sg13g2_xor2_1 _07715_ (.B(_02173_),
    .A(_02171_),
    .X(_02217_));
 sg13g2_nor3_1 _07716_ (.A(_02216_),
    .B(_02217_),
    .C(net116),
    .Y(_02218_));
 sg13g2_o21ai_1 _07717_ (.B1(_02165_),
    .Y(_02219_),
    .A1(_02214_),
    .A2(_02218_));
 sg13g2_nor3_1 _07718_ (.A(_02166_),
    .B(_02170_),
    .C(net116),
    .Y(_02220_));
 sg13g2_nor2_1 _07719_ (.A(_02166_),
    .B(net116),
    .Y(_02221_));
 sg13g2_nor4_1 _07720_ (.A(_02166_),
    .B(_02216_),
    .C(_02217_),
    .D(net116),
    .Y(_02222_));
 sg13g2_a221oi_1 _07721_ (.B2(_02165_),
    .C1(_02222_),
    .B1(_02221_),
    .A1(_02217_),
    .Y(_02223_),
    .A2(_02220_));
 sg13g2_nand3_1 _07722_ (.B(_02217_),
    .C(net116),
    .A(_02170_),
    .Y(_02224_));
 sg13g2_nand3_1 _07723_ (.B(_02174_),
    .C(net116),
    .A(_02216_),
    .Y(_02225_));
 sg13g2_a21o_1 _07724_ (.A2(_02225_),
    .A1(_02224_),
    .B1(_02165_),
    .X(_02226_));
 sg13g2_nand4_1 _07725_ (.B(_02170_),
    .C(_02217_),
    .A(_02166_),
    .Y(_02227_),
    .D(net116));
 sg13g2_nand4_1 _07726_ (.B(_02216_),
    .C(_02174_),
    .A(_02166_),
    .Y(_02228_),
    .D(net116));
 sg13g2_nand2_1 _07727_ (.Y(_02229_),
    .A(_02083_),
    .B(_01785_));
 sg13g2_or4_1 _07728_ (.A(_02167_),
    .B(_02162_),
    .C(_02163_),
    .D(_02229_),
    .X(_02230_));
 sg13g2_and3_1 _07729_ (.X(_02231_),
    .A(_02227_),
    .B(_02228_),
    .C(_02230_));
 sg13g2_nand4_1 _07730_ (.B(_02223_),
    .C(_02226_),
    .A(_02219_),
    .Y(_02232_),
    .D(_02231_));
 sg13g2_xnor2_1 _07731_ (.Y(_02233_),
    .A(_02211_),
    .B(_02232_));
 sg13g2_xnor2_1 _07732_ (.Y(_02234_),
    .A(_02200_),
    .B(_02233_));
 sg13g2_xnor2_1 _07733_ (.Y(_00027_),
    .A(_02196_),
    .B(_02234_));
 sg13g2_or2_1 _07734_ (.X(_02235_),
    .B(_02233_),
    .A(_02200_));
 sg13g2_inv_1 _07735_ (.Y(_02236_),
    .A(_02235_));
 sg13g2_nand2_1 _07736_ (.Y(_02237_),
    .A(_02200_),
    .B(_02233_));
 sg13g2_o21ai_1 _07737_ (.B1(_02237_),
    .Y(_02238_),
    .A1(_02196_),
    .A2(_02236_));
 sg13g2_nor2_1 _07738_ (.A(_02211_),
    .B(_02229_),
    .Y(_02239_));
 sg13g2_nor2_1 _07739_ (.A(_02165_),
    .B(_02175_),
    .Y(_02240_));
 sg13g2_nor2_1 _07740_ (.A(_02166_),
    .B(_02240_),
    .Y(_02241_));
 sg13g2_a221oi_1 _07741_ (.B2(_02229_),
    .C1(_02241_),
    .B1(_02211_),
    .A1(_02165_),
    .Y(_02242_),
    .A2(_02175_));
 sg13g2_nor2_2 _07742_ (.A(_02239_),
    .B(_02242_),
    .Y(_02243_));
 sg13g2_nand2_1 _07743_ (.Y(_02244_),
    .A(_02205_),
    .B(_02206_));
 sg13g2_o21ai_1 _07744_ (.B1(_02207_),
    .Y(_02245_),
    .A1(_02205_),
    .A2(_02206_));
 sg13g2_nand2_1 _07745_ (.Y(_02246_),
    .A(_02244_),
    .B(_02245_));
 sg13g2_inv_1 _07746_ (.Y(_02247_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[12] ));
 sg13g2_buf_2 _07747_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .X(_02248_));
 sg13g2_nand2_1 _07748_ (.Y(_02249_),
    .A(_02248_),
    .B(_01824_));
 sg13g2_nand2_1 _07749_ (.Y(_02250_),
    .A(_02204_),
    .B(_01828_));
 sg13g2_nand3_1 _07750_ (.B(_02168_),
    .C(_01877_),
    .A(_01217_),
    .Y(_02251_));
 sg13g2_xnor2_1 _07751_ (.Y(_02252_),
    .A(_02250_),
    .B(_02251_));
 sg13g2_xnor2_1 _07752_ (.Y(_02253_),
    .A(_02249_),
    .B(_02252_));
 sg13g2_xnor2_1 _07753_ (.Y(_02254_),
    .A(_02247_),
    .B(_02253_));
 sg13g2_xnor2_1 _07754_ (.Y(_02255_),
    .A(_02246_),
    .B(_02254_));
 sg13g2_nor2_1 _07755_ (.A(_02203_),
    .B(_02209_),
    .Y(_02256_));
 sg13g2_nand2_1 _07756_ (.Y(_02257_),
    .A(_02203_),
    .B(_02209_));
 sg13g2_o21ai_1 _07757_ (.B1(_02257_),
    .Y(_02258_),
    .A1(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .A2(_02256_));
 sg13g2_nand2_1 _07758_ (.Y(_02259_),
    .A(_02137_),
    .B(net132));
 sg13g2_xnor2_1 _07759_ (.Y(_02260_),
    .A(_02258_),
    .B(_02259_));
 sg13g2_xnor2_1 _07760_ (.Y(_02261_),
    .A(_02255_),
    .B(_02260_));
 sg13g2_xor2_1 _07761_ (.B(_02261_),
    .A(_02243_),
    .X(_02262_));
 sg13g2_xnor2_1 _07762_ (.Y(_00028_),
    .A(_02238_),
    .B(_02262_));
 sg13g2_a22oi_1 _07763_ (.Y(_02263_),
    .B1(_02200_),
    .B2(_02233_),
    .A2(_02191_),
    .A1(_02183_));
 sg13g2_and2_1 _07764_ (.A(_02156_),
    .B(_02263_),
    .X(_02264_));
 sg13g2_and3_1 _07765_ (.X(_02265_),
    .A(_02122_),
    .B(_02156_),
    .C(_02263_));
 sg13g2_and3_1 _07766_ (.X(_02266_),
    .A(_02148_),
    .B(_02157_),
    .C(_02263_));
 sg13g2_a221oi_1 _07767_ (.B2(_02041_),
    .C1(_02266_),
    .B1(_02265_),
    .A1(_02128_),
    .Y(_02267_),
    .A2(_02264_));
 sg13g2_nor2_1 _07768_ (.A(_02243_),
    .B(_02261_),
    .Y(_02268_));
 sg13g2_nand2b_1 _07769_ (.Y(_02269_),
    .B(_02193_),
    .A_N(_02183_));
 sg13g2_and2_1 _07770_ (.A(_02200_),
    .B(_02233_),
    .X(_02270_));
 sg13g2_a21oi_1 _07771_ (.A1(_02235_),
    .A2(_02269_),
    .Y(_02271_),
    .B1(_02270_));
 sg13g2_nor2_1 _07772_ (.A(_02268_),
    .B(_02271_),
    .Y(_02272_));
 sg13g2_a22oi_1 _07773_ (.Y(_02273_),
    .B1(_02267_),
    .B2(_02272_),
    .A2(_02261_),
    .A1(_02243_));
 sg13g2_a21oi_2 _07774_ (.B1(_02258_),
    .Y(_02274_),
    .A2(_02259_),
    .A1(_02255_));
 sg13g2_nor2_1 _07775_ (.A(_02255_),
    .B(_02259_),
    .Y(_02275_));
 sg13g2_nor2_2 _07776_ (.A(_02274_),
    .B(_02275_),
    .Y(_02276_));
 sg13g2_a21o_1 _07777_ (.A2(_02253_),
    .A1(_02246_),
    .B1(_02247_),
    .X(_02277_));
 sg13g2_o21ai_1 _07778_ (.B1(_02277_),
    .Y(_02278_),
    .A1(_02246_),
    .A2(_02253_));
 sg13g2_buf_2 _07779_ (.A(_02278_),
    .X(_02279_));
 sg13g2_nand2_1 _07780_ (.Y(_02280_),
    .A(_02249_),
    .B(_02250_));
 sg13g2_o21ai_1 _07781_ (.B1(_02251_),
    .Y(_02281_),
    .A1(_02249_),
    .A2(_02250_));
 sg13g2_nand2_1 _07782_ (.Y(_02282_),
    .A(_02280_),
    .B(_02281_));
 sg13g2_buf_1 _07783_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .X(_02283_));
 sg13g2_buf_1 _07784_ (.A(net131),
    .X(_02284_));
 sg13g2_nand2_1 _07785_ (.Y(_02285_),
    .A(net299),
    .B(net115));
 sg13g2_nand2_1 _07786_ (.Y(_02286_),
    .A(_02248_),
    .B(net144));
 sg13g2_nand2_1 _07787_ (.Y(_02287_),
    .A(_02204_),
    .B(net129));
 sg13g2_xnor2_1 _07788_ (.Y(_02288_),
    .A(_02286_),
    .B(_02287_));
 sg13g2_xnor2_1 _07789_ (.Y(_02289_),
    .A(_02285_),
    .B(_02288_));
 sg13g2_xor2_1 _07790_ (.B(_02289_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[13] ),
    .X(_02290_));
 sg13g2_xnor2_1 _07791_ (.Y(_02291_),
    .A(_02282_),
    .B(_02290_));
 sg13g2_buf_1 _07792_ (.A(_01786_),
    .X(_02292_));
 sg13g2_nand2_1 _07793_ (.Y(_02293_),
    .A(_02168_),
    .B(_02292_));
 sg13g2_xor2_1 _07794_ (.B(_02293_),
    .A(_02291_),
    .X(_02294_));
 sg13g2_xnor2_1 _07795_ (.Y(_02295_),
    .A(_02279_),
    .B(_02294_));
 sg13g2_xnor2_1 _07796_ (.Y(_02296_),
    .A(_02276_),
    .B(_02295_));
 sg13g2_xnor2_1 _07797_ (.Y(_00029_),
    .A(_02273_),
    .B(_02296_));
 sg13g2_nand2_1 _07798_ (.Y(_02297_),
    .A(_02282_),
    .B(_02289_));
 sg13g2_nor2_1 _07799_ (.A(_02282_),
    .B(_02289_),
    .Y(_02298_));
 sg13g2_a21oi_2 _07800_ (.B1(_02298_),
    .Y(_02299_),
    .A2(_02297_),
    .A1(\i_tinyqv.cpu.i_core.multiplier.accum[13] ));
 sg13g2_nand2_1 _07801_ (.Y(_02300_),
    .A(_02285_),
    .B(_02286_));
 sg13g2_o21ai_1 _07802_ (.B1(_02287_),
    .Y(_02301_),
    .A1(_02285_),
    .A2(_02286_));
 sg13g2_nand2_1 _07803_ (.Y(_02302_),
    .A(_02300_),
    .B(_02301_));
 sg13g2_buf_1 _07804_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .X(_02303_));
 sg13g2_nand2_1 _07805_ (.Y(_02304_),
    .A(_02303_),
    .B(_01824_));
 sg13g2_nand2_2 _07806_ (.Y(_02305_),
    .A(net299),
    .B(net157));
 sg13g2_nand3_1 _07807_ (.B(_02248_),
    .C(_01877_),
    .A(_01217_),
    .Y(_02306_));
 sg13g2_xnor2_1 _07808_ (.Y(_02307_),
    .A(_02305_),
    .B(_02306_));
 sg13g2_xnor2_1 _07809_ (.Y(_02308_),
    .A(_02304_),
    .B(_02307_));
 sg13g2_xor2_1 _07810_ (.B(_02308_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[14] ),
    .X(_02309_));
 sg13g2_xnor2_1 _07811_ (.Y(_02310_),
    .A(_02302_),
    .B(_02309_));
 sg13g2_nand2_1 _07812_ (.Y(_02311_),
    .A(_02204_),
    .B(_01786_));
 sg13g2_xor2_1 _07813_ (.B(_02311_),
    .A(_02310_),
    .X(_02312_));
 sg13g2_xnor2_1 _07814_ (.Y(_02313_),
    .A(_02299_),
    .B(_02312_));
 sg13g2_nor2_2 _07815_ (.A(_02291_),
    .B(_02293_),
    .Y(_02314_));
 sg13g2_nor2b_1 _07816_ (.A(_02276_),
    .B_N(_02279_),
    .Y(_02315_));
 sg13g2_nand2_1 _07817_ (.Y(_02316_),
    .A(_02291_),
    .B(_02293_));
 sg13g2_nor2_1 _07818_ (.A(_02279_),
    .B(_02316_),
    .Y(_02317_));
 sg13g2_a22oi_1 _07819_ (.Y(_02318_),
    .B1(_02317_),
    .B2(_02276_),
    .A2(_02315_),
    .A1(_02314_));
 sg13g2_a21oi_1 _07820_ (.A1(_02279_),
    .A2(_02316_),
    .Y(_02319_),
    .B1(_02314_));
 sg13g2_a21oi_1 _07821_ (.A1(_02276_),
    .A2(_02319_),
    .Y(_02320_),
    .B1(_02317_));
 sg13g2_nor2_1 _07822_ (.A(_02276_),
    .B(_02319_),
    .Y(_02321_));
 sg13g2_a21oi_1 _07823_ (.A1(_02279_),
    .A2(_02314_),
    .Y(_02322_),
    .B1(_02321_));
 sg13g2_mux2_1 _07824_ (.A0(_02320_),
    .A1(_02322_),
    .S(_02273_),
    .X(_02323_));
 sg13g2_nand2_1 _07825_ (.Y(_02324_),
    .A(_02318_),
    .B(_02323_));
 sg13g2_xnor2_1 _07826_ (.Y(_00019_),
    .A(_02313_),
    .B(_02324_));
 sg13g2_o21ai_1 _07827_ (.B1(_02279_),
    .Y(_02325_),
    .A1(_02274_),
    .A2(_02275_));
 sg13g2_nor2_1 _07828_ (.A(_02313_),
    .B(_02314_),
    .Y(_02326_));
 sg13g2_or3_1 _07829_ (.A(_02274_),
    .B(_02275_),
    .C(_02279_),
    .X(_02327_));
 sg13g2_and2_1 _07830_ (.A(_02313_),
    .B(_02327_),
    .X(_02328_));
 sg13g2_nor4_1 _07831_ (.A(_02268_),
    .B(_02271_),
    .C(_02314_),
    .D(_02328_),
    .Y(_02329_));
 sg13g2_nand2_1 _07832_ (.Y(_02330_),
    .A(_02243_),
    .B(_02261_));
 sg13g2_nor3_1 _07833_ (.A(_02330_),
    .B(_02314_),
    .C(_02328_),
    .Y(_02331_));
 sg13g2_a221oi_1 _07834_ (.B2(_02267_),
    .C1(_02331_),
    .B1(_02329_),
    .A1(_02325_),
    .Y(_02332_),
    .A2(_02326_));
 sg13g2_inv_1 _07835_ (.Y(_02333_),
    .A(_02313_));
 sg13g2_inv_1 _07836_ (.Y(_02334_),
    .A(_02316_));
 sg13g2_and2_1 _07837_ (.A(_02313_),
    .B(_02316_),
    .X(_02335_));
 sg13g2_nor4_1 _07838_ (.A(_02268_),
    .B(_02271_),
    .C(_02315_),
    .D(_02335_),
    .Y(_02336_));
 sg13g2_nand3_1 _07839_ (.B(_02261_),
    .C(_02325_),
    .A(_02243_),
    .Y(_02337_));
 sg13g2_a21oi_1 _07840_ (.A1(_02327_),
    .A2(_02337_),
    .Y(_02338_),
    .B1(_02335_));
 sg13g2_a221oi_1 _07841_ (.B2(_02267_),
    .C1(_02338_),
    .B1(_02336_),
    .A1(_02333_),
    .Y(_02339_),
    .A2(_02334_));
 sg13g2_and2_1 _07842_ (.A(_02332_),
    .B(_02339_),
    .X(_02340_));
 sg13g2_nand2_1 _07843_ (.Y(_02341_),
    .A(_02299_),
    .B(_02310_));
 sg13g2_o21ai_1 _07844_ (.B1(_02311_),
    .Y(_02342_),
    .A1(_02299_),
    .A2(_02310_));
 sg13g2_nand2_1 _07845_ (.Y(_02343_),
    .A(_02341_),
    .B(_02342_));
 sg13g2_nand2_1 _07846_ (.Y(_02344_),
    .A(_02304_),
    .B(_02305_));
 sg13g2_o21ai_1 _07847_ (.B1(_02306_),
    .Y(_02345_),
    .A1(_02304_),
    .A2(_02305_));
 sg13g2_nand2_1 _07848_ (.Y(_02346_),
    .A(_02344_),
    .B(_02345_));
 sg13g2_nand2_1 _07849_ (.Y(_02347_),
    .A(net299),
    .B(net129));
 sg13g2_nand2_1 _07850_ (.Y(_02348_),
    .A(_02303_),
    .B(net144));
 sg13g2_xnor2_1 _07851_ (.Y(_02349_),
    .A(_02347_),
    .B(_02348_));
 sg13g2_buf_1 _07852_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .X(_02350_));
 sg13g2_nand2_1 _07853_ (.Y(_02351_),
    .A(_02350_),
    .B(net115));
 sg13g2_xnor2_1 _07854_ (.Y(_02352_),
    .A(_02349_),
    .B(_02351_));
 sg13g2_xor2_1 _07855_ (.B(_02352_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .X(_02353_));
 sg13g2_xnor2_1 _07856_ (.Y(_02354_),
    .A(_02346_),
    .B(_02353_));
 sg13g2_nand2_1 _07857_ (.Y(_02355_),
    .A(_02302_),
    .B(_02308_));
 sg13g2_nor2_1 _07858_ (.A(_02302_),
    .B(_02308_),
    .Y(_02356_));
 sg13g2_a21oi_2 _07859_ (.B1(_02356_),
    .Y(_02357_),
    .A2(_02355_),
    .A1(\i_tinyqv.cpu.i_core.multiplier.accum[14] ));
 sg13g2_nand2_1 _07860_ (.Y(_02358_),
    .A(_02248_),
    .B(_02292_));
 sg13g2_xnor2_1 _07861_ (.Y(_02359_),
    .A(_02357_),
    .B(_02358_));
 sg13g2_xnor2_1 _07862_ (.Y(_02360_),
    .A(_02354_),
    .B(_02359_));
 sg13g2_nor2_1 _07863_ (.A(_02343_),
    .B(_02360_),
    .Y(_02361_));
 sg13g2_nand2_1 _07864_ (.Y(_02362_),
    .A(_02343_),
    .B(_02360_));
 sg13g2_nand2b_1 _07865_ (.Y(_02363_),
    .B(_02362_),
    .A_N(_02361_));
 sg13g2_xnor2_1 _07866_ (.Y(_00020_),
    .A(_02340_),
    .B(_02363_));
 sg13g2_nor2b_1 _07867_ (.A(_01669_),
    .B_N(net233),
    .Y(_02364_));
 sg13g2_buf_1 _07868_ (.A(_02364_),
    .X(_02365_));
 sg13g2_nand2b_1 _07869_ (.Y(_02366_),
    .B(net270),
    .A_N(_01774_));
 sg13g2_buf_1 _07870_ (.A(_02366_),
    .X(_02367_));
 sg13g2_nand2b_1 _07871_ (.Y(_02368_),
    .B(net278),
    .A_N(_00817_));
 sg13g2_buf_1 _07872_ (.A(_02368_),
    .X(_02369_));
 sg13g2_nor2_1 _07873_ (.A(_02367_),
    .B(_02369_),
    .Y(_02370_));
 sg13g2_buf_2 _07874_ (.A(_02370_),
    .X(_02371_));
 sg13g2_buf_2 _07875_ (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .X(_02372_));
 sg13g2_xor2_1 _07876_ (.B(_02372_),
    .A(net274),
    .X(_02373_));
 sg13g2_mux2_1 _07877_ (.A0(_00198_),
    .A1(_00197_),
    .S(_02373_),
    .X(_02374_));
 sg13g2_buf_2 _07878_ (.A(net335),
    .X(_02375_));
 sg13g2_buf_1 _07879_ (.A(_02372_),
    .X(_02376_));
 sg13g2_mux4_1 _07880_ (.S0(net268),
    .A0(_00190_),
    .A1(_00189_),
    .A2(_00192_),
    .A3(_00191_),
    .S1(net267),
    .X(_02377_));
 sg13g2_buf_1 _07881_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .X(_02378_));
 sg13g2_xnor2_1 _07882_ (.Y(_02379_),
    .A(net335),
    .B(_02378_));
 sg13g2_xnor2_1 _07883_ (.Y(_02380_),
    .A(_00847_),
    .B(_02379_));
 sg13g2_buf_2 _07884_ (.A(_02380_),
    .X(_02381_));
 sg13g2_buf_1 _07885_ (.A(_02381_),
    .X(_02382_));
 sg13g2_mux2_1 _07886_ (.A0(_02374_),
    .A1(_02377_),
    .S(net181),
    .X(_02383_));
 sg13g2_buf_1 _07887_ (.A(_02372_),
    .X(_02384_));
 sg13g2_mux4_1 _07888_ (.S0(net268),
    .A0(_00195_),
    .A1(_00196_),
    .A2(_00193_),
    .A3(_00194_),
    .S1(net266),
    .X(_02385_));
 sg13g2_mux4_1 _07889_ (.S0(net268),
    .A0(_00194_),
    .A1(_00193_),
    .A2(_00196_),
    .A3(_00195_),
    .S1(net267),
    .X(_02386_));
 sg13g2_mux2_1 _07890_ (.A0(_02385_),
    .A1(_02386_),
    .S(net181),
    .X(_02387_));
 sg13g2_buf_2 _07891_ (.A(net335),
    .X(_02388_));
 sg13g2_mux4_1 _07892_ (.S0(net265),
    .A0(_00182_),
    .A1(_00181_),
    .A2(_00184_),
    .A3(_00183_),
    .S1(net267),
    .X(_02389_));
 sg13g2_buf_1 _07893_ (.A(_00173_),
    .X(_02390_));
 sg13g2_buf_1 _07894_ (.A(_02372_),
    .X(_02391_));
 sg13g2_mux4_1 _07895_ (.S0(net265),
    .A0(_00174_),
    .A1(_02390_),
    .A2(_00176_),
    .A3(_00175_),
    .S1(net264),
    .X(_02392_));
 sg13g2_mux2_1 _07896_ (.A0(_02389_),
    .A1(_02392_),
    .S(_02381_),
    .X(_02393_));
 sg13g2_mux4_1 _07897_ (.S0(net265),
    .A0(_00186_),
    .A1(_00185_),
    .A2(_00188_),
    .A3(_00187_),
    .S1(net267),
    .X(_02394_));
 sg13g2_mux4_1 _07898_ (.S0(net265),
    .A0(_00178_),
    .A1(_00177_),
    .A2(_00180_),
    .A3(_00179_),
    .S1(net267),
    .X(_02395_));
 sg13g2_mux2_1 _07899_ (.A0(_02394_),
    .A1(_02395_),
    .S(net181),
    .X(_02396_));
 sg13g2_buf_1 _07900_ (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .X(_02397_));
 sg13g2_buf_1 _07901_ (.A(_00839_),
    .X(_02398_));
 sg13g2_buf_1 _07902_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .X(_02399_));
 sg13g2_xor2_1 _07903_ (.B(_02399_),
    .A(net219),
    .X(_02400_));
 sg13g2_nor2b_1 _07904_ (.A(_02378_),
    .B_N(net274),
    .Y(_02401_));
 sg13g2_a21oi_1 _07905_ (.A1(net223),
    .A2(_02378_),
    .Y(_02402_),
    .B1(_02401_));
 sg13g2_xnor2_1 _07906_ (.Y(_02403_),
    .A(_02400_),
    .B(_02402_));
 sg13g2_buf_4 _07907_ (.X(_02404_),
    .A(_02403_));
 sg13g2_mux4_1 _07908_ (.S0(net298),
    .A0(_02383_),
    .A1(_02387_),
    .A2(_02393_),
    .A3(_02396_),
    .S1(_02404_),
    .X(_02405_));
 sg13g2_buf_1 _07909_ (.A(_02381_),
    .X(_02406_));
 sg13g2_buf_1 _07910_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .X(_02407_));
 sg13g2_nand2_2 _07911_ (.Y(_02408_),
    .A(_00888_),
    .B(_02407_));
 sg13g2_nand2_1 _07912_ (.Y(_02409_),
    .A(net274),
    .B(_00203_));
 sg13g2_nand2b_1 _07913_ (.Y(_02410_),
    .B(_00172_),
    .A_N(net274));
 sg13g2_a21oi_1 _07914_ (.A1(_02409_),
    .A2(_02410_),
    .Y(_02411_),
    .B1(net264));
 sg13g2_a21oi_1 _07915_ (.A1(net266),
    .A2(_02408_),
    .Y(_02412_),
    .B1(_02411_));
 sg13g2_mux4_1 _07916_ (.S0(net274),
    .A0(_00175_),
    .A1(_00176_),
    .A2(_02390_),
    .A3(_00174_),
    .S1(_02372_),
    .X(_02413_));
 sg13g2_nand2_1 _07917_ (.Y(_02414_),
    .A(_02381_),
    .B(_02413_));
 sg13g2_o21ai_1 _07918_ (.B1(_02414_),
    .Y(_02415_),
    .A1(net180),
    .A2(_02412_));
 sg13g2_buf_1 _07919_ (.A(_00199_),
    .X(_02416_));
 sg13g2_buf_1 _07920_ (.A(_00201_),
    .X(_02417_));
 sg13g2_mux4_1 _07921_ (.S0(net274),
    .A0(_02416_),
    .A1(_00200_),
    .A2(_02417_),
    .A3(_00202_),
    .S1(net264),
    .X(_02418_));
 sg13g2_nor2b_1 _07922_ (.A(_02381_),
    .B_N(_02408_),
    .Y(_02419_));
 sg13g2_a21o_1 _07923_ (.A2(_02418_),
    .A1(net180),
    .B1(_02419_),
    .X(_02420_));
 sg13g2_mux4_1 _07924_ (.S0(net265),
    .A0(_00183_),
    .A1(_00184_),
    .A2(_00181_),
    .A3(_00182_),
    .S1(net264),
    .X(_02421_));
 sg13g2_mux4_1 _07925_ (.S0(net274),
    .A0(_00191_),
    .A1(_00192_),
    .A2(_00189_),
    .A3(_00190_),
    .S1(net264),
    .X(_02422_));
 sg13g2_mux2_1 _07926_ (.A0(_02421_),
    .A1(_02422_),
    .S(_02381_),
    .X(_02423_));
 sg13g2_mux4_1 _07927_ (.S0(_01672_),
    .A0(_00179_),
    .A1(_00180_),
    .A2(_00177_),
    .A3(_00178_),
    .S1(net264),
    .X(_02424_));
 sg13g2_mux4_1 _07928_ (.S0(_01672_),
    .A0(_00187_),
    .A1(_00188_),
    .A2(_00185_),
    .A3(_00186_),
    .S1(net264),
    .X(_02425_));
 sg13g2_mux2_1 _07929_ (.A0(_02424_),
    .A1(_02425_),
    .S(net181),
    .X(_02426_));
 sg13g2_mux4_1 _07930_ (.S0(net298),
    .A0(_02415_),
    .A1(_02420_),
    .A2(_02423_),
    .A3(_02426_),
    .S1(_02404_),
    .X(_02427_));
 sg13g2_buf_1 _07931_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .X(_02428_));
 sg13g2_xor2_1 _07932_ (.B(net234),
    .A(net335),
    .X(_02429_));
 sg13g2_xnor2_1 _07933_ (.Y(_02430_),
    .A(_02428_),
    .B(_02429_));
 sg13g2_nor2b_1 _07934_ (.A(net219),
    .B_N(_02399_),
    .Y(_02431_));
 sg13g2_a21oi_1 _07935_ (.A1(net219),
    .A2(net335),
    .Y(_02432_),
    .B1(_02431_));
 sg13g2_nand2_1 _07936_ (.Y(_02433_),
    .A(net219),
    .B(_02399_));
 sg13g2_o21ai_1 _07937_ (.B1(_02433_),
    .Y(_02434_),
    .A1(net219),
    .A2(net335));
 sg13g2_nor2_1 _07938_ (.A(_00847_),
    .B(_02434_),
    .Y(_02435_));
 sg13g2_a21oi_1 _07939_ (.A1(net240),
    .A2(_02432_),
    .Y(_02436_),
    .B1(_02435_));
 sg13g2_xnor2_1 _07940_ (.Y(_02437_),
    .A(net219),
    .B(net335));
 sg13g2_a22oi_1 _07941_ (.Y(_02438_),
    .B1(_02437_),
    .B2(_02399_),
    .A2(_02436_),
    .A1(_02378_));
 sg13g2_nand2b_1 _07942_ (.Y(_02439_),
    .B(_02438_),
    .A_N(_02430_));
 sg13g2_buf_4 _07943_ (.X(_02440_),
    .A(_02439_));
 sg13g2_mux2_1 _07944_ (.A0(_02405_),
    .A1(_02427_),
    .S(_02440_),
    .X(_02441_));
 sg13g2_nand2b_1 _07945_ (.Y(_02442_),
    .B(_02428_),
    .A_N(_02438_));
 sg13g2_nor2b_1 _07946_ (.A(_02428_),
    .B_N(_02438_),
    .Y(_02443_));
 sg13g2_a21oi_2 _07947_ (.B1(_02443_),
    .Y(_02444_),
    .A2(_02429_),
    .A1(_02442_));
 sg13g2_mux2_1 _07948_ (.A0(_02441_),
    .A1(_02408_),
    .S(_02444_),
    .X(_02445_));
 sg13g2_buf_1 _07949_ (.A(net335),
    .X(_02446_));
 sg13g2_mux4_1 _07950_ (.S0(net263),
    .A0(_00192_),
    .A1(_00191_),
    .A2(_00194_),
    .A3(_00193_),
    .S1(net266),
    .X(_02447_));
 sg13g2_mux4_1 _07951_ (.S0(_02375_),
    .A0(_00184_),
    .A1(_00183_),
    .A2(_00186_),
    .A3(_00185_),
    .S1(net266),
    .X(_02448_));
 sg13g2_mux2_1 _07952_ (.A0(_02447_),
    .A1(_02448_),
    .S(net180),
    .X(_02449_));
 sg13g2_mux4_1 _07953_ (.S0(_02446_),
    .A0(_00196_),
    .A1(_00195_),
    .A2(_00198_),
    .A3(_00197_),
    .S1(net266),
    .X(_02450_));
 sg13g2_mux4_1 _07954_ (.S0(net268),
    .A0(_00188_),
    .A1(_00187_),
    .A2(_00190_),
    .A3(_00189_),
    .S1(_02384_),
    .X(_02451_));
 sg13g2_mux2_1 _07955_ (.A0(_02450_),
    .A1(_02451_),
    .S(_02382_),
    .X(_02452_));
 sg13g2_mux4_1 _07956_ (.S0(_02372_),
    .A0(_02390_),
    .A1(_02416_),
    .A2(_00174_),
    .A3(_00200_),
    .S1(net263),
    .X(_02453_));
 sg13g2_mux4_1 _07957_ (.S0(net265),
    .A0(_00181_),
    .A1(_00182_),
    .A2(_00179_),
    .A3(_00180_),
    .S1(net267),
    .X(_02454_));
 sg13g2_mux2_1 _07958_ (.A0(_02453_),
    .A1(_02454_),
    .S(net181),
    .X(_02455_));
 sg13g2_mux4_1 _07959_ (.S0(net268),
    .A0(_02417_),
    .A1(_00202_),
    .A2(_00172_),
    .A3(_00203_),
    .S1(net267),
    .X(_02456_));
 sg13g2_mux4_1 _07960_ (.S0(net265),
    .A0(_00177_),
    .A1(_00178_),
    .A2(_00175_),
    .A3(_00176_),
    .S1(net264),
    .X(_02457_));
 sg13g2_mux2_1 _07961_ (.A0(_02456_),
    .A1(_02457_),
    .S(net181),
    .X(_02458_));
 sg13g2_mux4_1 _07962_ (.S0(net298),
    .A0(_02449_),
    .A1(_02452_),
    .A2(_02455_),
    .A3(_02458_),
    .S1(_02440_),
    .X(_02459_));
 sg13g2_mux4_1 _07963_ (.S0(net268),
    .A0(_00176_),
    .A1(_00175_),
    .A2(_00178_),
    .A3(_00177_),
    .S1(net266),
    .X(_02460_));
 sg13g2_mux4_1 _07964_ (.S0(_02372_),
    .A0(_00203_),
    .A1(_00202_),
    .A2(_00172_),
    .A3(_02417_),
    .S1(net263),
    .X(_02461_));
 sg13g2_mux2_1 _07965_ (.A0(_02460_),
    .A1(_02461_),
    .S(_02382_),
    .X(_02462_));
 sg13g2_mux4_1 _07966_ (.S0(net268),
    .A0(_00180_),
    .A1(_00179_),
    .A2(_00182_),
    .A3(_00181_),
    .S1(_02384_),
    .X(_02463_));
 sg13g2_mux4_1 _07967_ (.S0(net268),
    .A0(_00200_),
    .A1(_02416_),
    .A2(_00174_),
    .A3(_02390_),
    .S1(net267),
    .X(_02464_));
 sg13g2_mux2_1 _07968_ (.A0(_02463_),
    .A1(_02464_),
    .S(net181),
    .X(_02465_));
 sg13g2_mux4_1 _07969_ (.S0(_02388_),
    .A0(_00189_),
    .A1(_00190_),
    .A2(_00187_),
    .A3(_00188_),
    .S1(_02376_),
    .X(_02466_));
 sg13g2_mux4_1 _07970_ (.S0(_02388_),
    .A0(_00197_),
    .A1(_00198_),
    .A2(_00195_),
    .A3(_00196_),
    .S1(_02391_),
    .X(_02467_));
 sg13g2_mux2_1 _07971_ (.A0(_02466_),
    .A1(_02467_),
    .S(net181),
    .X(_02468_));
 sg13g2_mux4_1 _07972_ (.S0(_02375_),
    .A0(_00185_),
    .A1(_00186_),
    .A2(_00183_),
    .A3(_00184_),
    .S1(_02376_),
    .X(_02469_));
 sg13g2_mux4_1 _07973_ (.S0(net265),
    .A0(_00193_),
    .A1(_00194_),
    .A2(_00191_),
    .A3(_00192_),
    .S1(_02391_),
    .X(_02470_));
 sg13g2_mux2_1 _07974_ (.A0(_02469_),
    .A1(_02470_),
    .S(_02381_),
    .X(_02471_));
 sg13g2_mux4_1 _07975_ (.S0(net298),
    .A0(_02462_),
    .A1(_02465_),
    .A2(_02468_),
    .A3(_02471_),
    .S1(_02440_),
    .X(_02472_));
 sg13g2_mux2_1 _07976_ (.A0(_02459_),
    .A1(_02472_),
    .S(_02404_),
    .X(_02473_));
 sg13g2_mux2_1 _07977_ (.A0(_02473_),
    .A1(_02408_),
    .S(_02444_),
    .X(_02474_));
 sg13g2_mux2_1 _07978_ (.A0(_02445_),
    .A1(_02474_),
    .S(net263),
    .X(_02475_));
 sg13g2_and4_1 _07979_ (.A(_00858_),
    .B(_01127_),
    .C(_01130_),
    .D(_01134_),
    .X(_02476_));
 sg13g2_a21oi_2 _07980_ (.B1(_02476_),
    .Y(_02477_),
    .A2(_01123_),
    .A1(_00938_));
 sg13g2_nand2_1 _07981_ (.Y(_02478_),
    .A(net224),
    .B(_01117_));
 sg13g2_o21ai_1 _07982_ (.B1(_02478_),
    .Y(_02479_),
    .A1(_00897_),
    .A2(_02477_));
 sg13g2_nor2_1 _07983_ (.A(net278),
    .B(net203),
    .Y(_02480_));
 sg13g2_and3_1 _07984_ (.X(_02481_),
    .A(_01218_),
    .B(_00889_),
    .C(_02480_));
 sg13g2_buf_1 _07985_ (.A(_02481_),
    .X(_02482_));
 sg13g2_xnor2_1 _07986_ (.Y(_02483_),
    .A(_00973_),
    .B(_01149_));
 sg13g2_nand2_1 _07987_ (.Y(_02484_),
    .A(_02482_),
    .B(_02483_));
 sg13g2_nor2b_1 _07988_ (.A(_02484_),
    .B_N(_01185_),
    .Y(_02485_));
 sg13g2_nand3_1 _07989_ (.B(_00889_),
    .C(_02480_),
    .A(_01218_),
    .Y(_02486_));
 sg13g2_buf_1 _07990_ (.A(_02486_),
    .X(_02487_));
 sg13g2_nor2_1 _07991_ (.A(net278),
    .B(_01218_),
    .Y(_02488_));
 sg13g2_nor2_1 _07992_ (.A(net203),
    .B(_02488_),
    .Y(_02489_));
 sg13g2_o21ai_1 _07993_ (.B1(_02489_),
    .Y(_02490_),
    .A1(_02487_),
    .A2(_02483_));
 sg13g2_nand2_1 _07994_ (.Y(_02491_),
    .A(_01256_),
    .B(_01257_));
 sg13g2_inv_1 _07995_ (.Y(_02492_),
    .A(_02491_));
 sg13g2_or3_1 _07996_ (.A(_01218_),
    .B(_00889_),
    .C(net203),
    .X(_02493_));
 sg13g2_buf_1 _07997_ (.A(_02493_),
    .X(_02494_));
 sg13g2_a21oi_1 _07998_ (.A1(_02484_),
    .A2(_02494_),
    .Y(_02495_),
    .B1(_01256_));
 sg13g2_a221oi_1 _07999_ (.B2(_02492_),
    .C1(_02495_),
    .B1(_02490_),
    .A1(_02479_),
    .Y(_02496_),
    .A2(_02485_));
 sg13g2_a21o_1 _08000_ (.A2(net115),
    .A1(net269),
    .B1(_01822_),
    .X(_02497_));
 sg13g2_a21oi_1 _08001_ (.A1(_01839_),
    .A2(_02497_),
    .Y(_02498_),
    .B1(net198));
 sg13g2_a21oi_1 _08002_ (.A1(net198),
    .A2(_02496_),
    .Y(_02499_),
    .B1(_02498_));
 sg13g2_nor2_1 _08003_ (.A(_02499_),
    .B(_02371_),
    .Y(_02500_));
 sg13g2_a21oi_1 _08004_ (.A1(_02371_),
    .A2(_02475_),
    .Y(_02501_),
    .B1(_02500_));
 sg13g2_buf_1 _08005_ (.A(_01146_),
    .X(_02502_));
 sg13g2_nand2b_1 _08006_ (.Y(_02503_),
    .B(_01673_),
    .A_N(_00888_));
 sg13g2_nor3_1 _08007_ (.A(net170),
    .B(_02367_),
    .C(_02503_),
    .Y(_02504_));
 sg13g2_mux2_1 _08008_ (.A0(_02501_),
    .A1(\i_tinyqv.cpu.i_core.cmp ),
    .S(_02504_),
    .X(_02505_));
 sg13g2_nor3_1 _08009_ (.A(_00172_),
    .B(_01174_),
    .C(_02367_),
    .Y(_02506_));
 sg13g2_a21oi_1 _08010_ (.A1(_01174_),
    .A2(_02505_),
    .Y(_02507_),
    .B1(_02506_));
 sg13g2_buf_1 _08011_ (.A(_01681_),
    .X(_02508_));
 sg13g2_buf_1 _08012_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .X(_02509_));
 sg13g2_buf_1 _08013_ (.A(net219),
    .X(_02510_));
 sg13g2_a21oi_1 _08014_ (.A1(net196),
    .A2(_01557_),
    .Y(_02511_),
    .B1(net234));
 sg13g2_nor2_1 _08015_ (.A(_02509_),
    .B(_02511_),
    .Y(_02512_));
 sg13g2_buf_1 _08016_ (.A(_02512_),
    .X(_02513_));
 sg13g2_buf_1 _08017_ (.A(net234),
    .X(_02514_));
 sg13g2_inv_1 _08018_ (.Y(_02515_),
    .A(_01698_));
 sg13g2_nand2_1 _08019_ (.Y(_02516_),
    .A(net310),
    .B(_01698_));
 sg13g2_inv_1 _08020_ (.Y(_02517_),
    .A(_01695_));
 sg13g2_a22oi_1 _08021_ (.Y(_02518_),
    .B1(_02516_),
    .B2(_02517_),
    .A2(_02515_),
    .A1(_01694_));
 sg13g2_nor2_1 _08022_ (.A(_01708_),
    .B(_02518_),
    .Y(_02519_));
 sg13g2_buf_2 _08023_ (.A(_02519_),
    .X(_02520_));
 sg13g2_nor2_2 _08024_ (.A(_01741_),
    .B(_01744_),
    .Y(_02521_));
 sg13g2_nand2b_1 _08025_ (.Y(_02522_),
    .B(_02521_),
    .A_N(_00171_));
 sg13g2_buf_1 _08026_ (.A(\i_tinyqv.cpu.instr_data_in[8] ),
    .X(_02523_));
 sg13g2_nor2_1 _08027_ (.A(_01305_),
    .B(_01307_),
    .Y(_02524_));
 sg13g2_nand2_1 _08028_ (.Y(_02525_),
    .A(net162),
    .B(_02524_));
 sg13g2_buf_1 _08029_ (.A(_02525_),
    .X(_02526_));
 sg13g2_nand2b_1 _08030_ (.Y(_02527_),
    .B(net125),
    .A_N(\i_tinyqv.mem.qspi_data_buf[8] ));
 sg13g2_o21ai_1 _08031_ (.B1(_02527_),
    .Y(_02528_),
    .A1(_02523_),
    .A2(net125));
 sg13g2_a221oi_1 _08032_ (.B2(_01300_),
    .C1(_01009_),
    .B1(_02528_),
    .A1(_02520_),
    .Y(_02529_),
    .A2(_02522_));
 sg13g2_buf_1 _08033_ (.A(net276),
    .X(_02530_));
 sg13g2_nor2b_1 _08034_ (.A(_01305_),
    .B_N(_01307_),
    .Y(_02531_));
 sg13g2_nand2_1 _08035_ (.Y(_02532_),
    .A(net162),
    .B(_02531_));
 sg13g2_buf_1 _08036_ (.A(_02532_),
    .X(_02533_));
 sg13g2_inv_1 _08037_ (.Y(_02534_),
    .A(\i_tinyqv.cpu.instr_data_in[0] ));
 sg13g2_nand2_1 _08038_ (.Y(_02535_),
    .A(_02534_),
    .B(_02533_));
 sg13g2_o21ai_1 _08039_ (.B1(_02535_),
    .Y(_02536_),
    .A1(_02523_),
    .A2(net124));
 sg13g2_nor2_1 _08040_ (.A(net310),
    .B(_01708_),
    .Y(_02537_));
 sg13g2_nand2_1 _08041_ (.Y(_02538_),
    .A(_01698_),
    .B(_02537_));
 sg13g2_nor3_1 _08042_ (.A(_01694_),
    .B(_01743_),
    .C(_02538_),
    .Y(_02539_));
 sg13g2_buf_1 _08043_ (.A(_02539_),
    .X(_02540_));
 sg13g2_nand2_2 _08044_ (.Y(_02541_),
    .A(_02515_),
    .B(_02537_));
 sg13g2_nand2_1 _08045_ (.Y(_02542_),
    .A(_01694_),
    .B(_02517_));
 sg13g2_nor2_1 _08046_ (.A(_02541_),
    .B(_02542_),
    .Y(_02543_));
 sg13g2_nor3_2 _08047_ (.A(net273),
    .B(net272),
    .C(_02541_),
    .Y(_02544_));
 sg13g2_and2_1 _08048_ (.A(net28),
    .B(_02544_),
    .X(_02545_));
 sg13g2_a221oi_1 _08049_ (.B2(net2),
    .C1(_02545_),
    .B1(_02543_),
    .A1(\i_spi.data[0] ),
    .Y(_02546_),
    .A2(net141));
 sg13g2_nand2_1 _08050_ (.Y(_02547_),
    .A(_01377_),
    .B(_01380_));
 sg13g2_and2_1 _08051_ (.A(net310),
    .B(_01740_),
    .X(_02548_));
 sg13g2_buf_1 _08052_ (.A(_02548_),
    .X(_02549_));
 sg13g2_buf_1 _08053_ (.A(_00169_),
    .X(_02550_));
 sg13g2_nor2_1 _08054_ (.A(_02550_),
    .B(_02538_),
    .Y(_02551_));
 sg13g2_a21oi_1 _08055_ (.A1(_02547_),
    .A2(_02549_),
    .Y(_02552_),
    .B1(_02551_));
 sg13g2_nor2_1 _08056_ (.A(_02542_),
    .B(_02552_),
    .Y(_02553_));
 sg13g2_buf_2 _08057_ (.A(\i_debug_uart_tx.fsm_state[1] ),
    .X(_02554_));
 sg13g2_buf_2 _08058_ (.A(\i_debug_uart_tx.fsm_state[2] ),
    .X(_02555_));
 sg13g2_nor2_2 _08059_ (.A(_02554_),
    .B(_02555_),
    .Y(_02556_));
 sg13g2_buf_2 _08060_ (.A(\i_debug_uart_tx.fsm_state[0] ),
    .X(_02557_));
 sg13g2_buf_2 _08061_ (.A(\i_debug_uart_tx.fsm_state[3] ),
    .X(_02558_));
 sg13g2_nor2_1 _08062_ (.A(_02557_),
    .B(_02558_),
    .Y(_02559_));
 sg13g2_and2_1 _08063_ (.A(_02556_),
    .B(_02559_),
    .X(_02560_));
 sg13g2_buf_1 _08064_ (.A(_02560_),
    .X(_02561_));
 sg13g2_nand2_1 _08065_ (.Y(_02562_),
    .A(net310),
    .B(net217));
 sg13g2_o21ai_1 _08066_ (.B1(_02562_),
    .Y(_02563_),
    .A1(_01697_),
    .A2(\gpio_out_sel[0] ));
 sg13g2_a21oi_1 _08067_ (.A1(net273),
    .A2(_02563_),
    .Y(_02564_),
    .B1(_02517_));
 sg13g2_nor2_1 _08068_ (.A(_01698_),
    .B(_02564_),
    .Y(_02565_));
 sg13g2_nor2_1 _08069_ (.A(net272),
    .B(net310),
    .Y(_02566_));
 sg13g2_and2_1 _08070_ (.A(_01696_),
    .B(_02549_),
    .X(_02567_));
 sg13g2_buf_1 _08071_ (.A(_02567_),
    .X(_02568_));
 sg13g2_nand2_1 _08072_ (.Y(_02569_),
    .A(\i_uart_rx.recieved_data[0] ),
    .B(net123));
 sg13g2_o21ai_1 _08073_ (.B1(_02569_),
    .Y(_02570_),
    .A1(_02565_),
    .A2(_02566_));
 sg13g2_nor3_1 _08074_ (.A(_01708_),
    .B(_02553_),
    .C(_02570_),
    .Y(_02571_));
 sg13g2_a221oi_1 _08075_ (.B2(_02571_),
    .C1(_01260_),
    .B1(_02546_),
    .A1(_02530_),
    .Y(_02572_),
    .A2(_02536_));
 sg13g2_buf_1 _08076_ (.A(net240),
    .X(_02573_));
 sg13g2_buf_1 _08077_ (.A(net216),
    .X(_02574_));
 sg13g2_nand2_2 _08078_ (.Y(_02575_),
    .A(net195),
    .B(net238));
 sg13g2_buf_1 _08079_ (.A(\i_tinyqv.cpu.instr_data_in[12] ),
    .X(_02576_));
 sg13g2_buf_1 _08080_ (.A(\i_tinyqv.cpu.instr_data_in[4] ),
    .X(_02577_));
 sg13g2_mux2_1 _08081_ (.A0(_02576_),
    .A1(_02577_),
    .S(net124),
    .X(_02578_));
 sg13g2_nor2_1 _08082_ (.A(_02541_),
    .B(_01744_),
    .Y(_02579_));
 sg13g2_a22oi_1 _08083_ (.Y(_02580_),
    .B1(net141),
    .B2(\i_spi.data[4] ),
    .A2(_02579_),
    .A1(\gpio_out_sel[4] ));
 sg13g2_nand2_1 _08084_ (.Y(_02581_),
    .A(net5),
    .B(_02543_));
 sg13g2_inv_1 _08085_ (.Y(_02582_),
    .A(_02520_));
 sg13g2_a221oi_1 _08086_ (.B2(\i_uart_rx.recieved_data[4] ),
    .C1(_02582_),
    .B1(net123),
    .A1(net32),
    .Y(_02583_),
    .A2(_02544_));
 sg13g2_nand3_1 _08087_ (.B(_02581_),
    .C(_02583_),
    .A(_02580_),
    .Y(_02584_));
 sg13g2_o21ai_1 _08088_ (.B1(_02584_),
    .Y(_02585_),
    .A1(_01350_),
    .A2(_02578_));
 sg13g2_mux2_1 _08089_ (.A0(_02576_),
    .A1(\i_tinyqv.mem.qspi_data_buf[12] ),
    .S(net125),
    .X(_02586_));
 sg13g2_nor2_1 _08090_ (.A(_01211_),
    .B(_02520_),
    .Y(_02587_));
 sg13g2_o21ai_1 _08091_ (.B1(_02587_),
    .Y(_02588_),
    .A1(_01350_),
    .A2(_02586_));
 sg13g2_o21ai_1 _08092_ (.B1(_02588_),
    .Y(_02589_),
    .A1(_02575_),
    .A2(_02585_));
 sg13g2_nor4_1 _08093_ (.A(net218),
    .B(_02529_),
    .C(_02572_),
    .D(_02589_),
    .Y(_02590_));
 sg13g2_buf_1 _08094_ (.A(net196),
    .X(_02591_));
 sg13g2_buf_1 _08095_ (.A(net216),
    .X(_02592_));
 sg13g2_and2_1 _08096_ (.A(net194),
    .B(\i_tinyqv.mem.data_from_read[20] ),
    .X(_02593_));
 sg13g2_a21oi_1 _08097_ (.A1(net223),
    .A2(\i_tinyqv.mem.data_from_read[16] ),
    .Y(_02594_),
    .B1(_02593_));
 sg13g2_mux4_1 _08098_ (.S0(net216),
    .A0(\i_tinyqv.mem.qspi_data_buf[24] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[28] ),
    .A2(_02523_),
    .A3(_02576_),
    .S1(net162),
    .X(_02595_));
 sg13g2_nand2_1 _08099_ (.Y(_02596_),
    .A(net196),
    .B(_02595_));
 sg13g2_o21ai_1 _08100_ (.B1(_02596_),
    .Y(_02597_),
    .A1(net179),
    .A2(_02594_));
 sg13g2_o21ai_1 _08101_ (.B1(net234),
    .Y(_02598_),
    .A1(_01300_),
    .A2(_02520_));
 sg13g2_buf_1 _08102_ (.A(_02598_),
    .X(_02599_));
 sg13g2_a21oi_1 _08103_ (.A1(net230),
    .A2(_02597_),
    .Y(_02600_),
    .B1(_02599_));
 sg13g2_nor3_1 _08104_ (.A(_02513_),
    .B(_02590_),
    .C(_02600_),
    .Y(_02601_));
 sg13g2_a21oi_1 _08105_ (.A1(\i_tinyqv.cpu.i_core.load_top_bit ),
    .A2(net156),
    .Y(_02602_),
    .B1(_02601_));
 sg13g2_buf_2 _08106_ (.A(_00163_),
    .X(_02603_));
 sg13g2_nand2_1 _08107_ (.Y(_02604_),
    .A(net333),
    .B(_01572_));
 sg13g2_buf_2 _08108_ (.A(_02604_),
    .X(_02605_));
 sg13g2_xnor2_1 _08109_ (.Y(_02606_),
    .A(_02603_),
    .B(_02605_));
 sg13g2_buf_1 _08110_ (.A(\i_tinyqv.cpu.instr_data_start[12] ),
    .X(_02607_));
 sg13g2_buf_1 _08111_ (.A(_00840_),
    .X(_02608_));
 sg13g2_and3_1 _08112_ (.X(_02609_),
    .A(_01025_),
    .B(_01065_),
    .C(_01178_));
 sg13g2_buf_1 _08113_ (.A(_02609_),
    .X(_02610_));
 sg13g2_buf_1 _08114_ (.A(_00831_),
    .X(_02611_));
 sg13g2_buf_1 _08115_ (.A(_01021_),
    .X(_02612_));
 sg13g2_buf_1 _08116_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .X(_02613_));
 sg13g2_nand4_1 _08117_ (.B(net260),
    .C(net296),
    .A(_02611_),
    .Y(_02614_),
    .D(_01179_));
 sg13g2_buf_1 _08118_ (.A(_02614_),
    .X(_02615_));
 sg13g2_nor2_2 _08119_ (.A(_02605_),
    .B(_02615_),
    .Y(_02616_));
 sg13g2_nand3_1 _08120_ (.B(_02610_),
    .C(_02616_),
    .A(net262),
    .Y(_02617_));
 sg13g2_xnor2_1 _08121_ (.Y(_02618_),
    .A(_02607_),
    .B(_02617_));
 sg13g2_nand2_1 _08122_ (.Y(_02619_),
    .A(_02398_),
    .B(_02618_));
 sg13g2_o21ai_1 _08123_ (.B1(_02619_),
    .Y(_02620_),
    .A1(net219),
    .A2(_02606_));
 sg13g2_buf_1 _08124_ (.A(_01178_),
    .X(_02621_));
 sg13g2_inv_1 _08125_ (.Y(_02622_),
    .A(net259));
 sg13g2_xnor2_1 _08126_ (.Y(_02623_),
    .A(_02622_),
    .B(_02616_));
 sg13g2_a22oi_1 _08127_ (.Y(_02624_),
    .B1(_02623_),
    .B2(_00900_),
    .A2(_02620_),
    .A1(net194));
 sg13g2_buf_1 _08128_ (.A(\i_tinyqv.cpu.instr_data_start[16] ),
    .X(_02625_));
 sg13g2_buf_1 _08129_ (.A(_00829_),
    .X(_02626_));
 sg13g2_nand2_1 _08130_ (.Y(_02627_),
    .A(net258),
    .B(net326));
 sg13g2_and4_1 _08131_ (.A(_02608_),
    .B(_01058_),
    .C(net297),
    .D(_02610_),
    .X(_02628_));
 sg13g2_buf_1 _08132_ (.A(_02628_),
    .X(_02629_));
 sg13g2_nand2_1 _08133_ (.Y(_02630_),
    .A(_02629_),
    .B(_02616_));
 sg13g2_nor2_1 _08134_ (.A(_02627_),
    .B(_02630_),
    .Y(_02631_));
 sg13g2_xnor2_1 _08135_ (.Y(_02632_),
    .A(net295),
    .B(_02631_));
 sg13g2_nand2_1 _08136_ (.Y(_02633_),
    .A(net334),
    .B(net327));
 sg13g2_nand4_1 _08137_ (.B(net326),
    .C(net324),
    .A(_00829_),
    .Y(_02634_),
    .D(net295));
 sg13g2_nor3_1 _08138_ (.A(_02633_),
    .B(_02615_),
    .C(_02634_),
    .Y(_02635_));
 sg13g2_nand2_1 _08139_ (.Y(_02636_),
    .A(_02629_),
    .B(_02635_));
 sg13g2_nor2_1 _08140_ (.A(_02605_),
    .B(_02636_),
    .Y(_02637_));
 sg13g2_xor2_1 _08141_ (.B(_02637_),
    .A(_01175_),
    .X(_02638_));
 sg13g2_nand2_1 _08142_ (.Y(_02639_),
    .A(net216),
    .B(_02638_));
 sg13g2_o21ai_1 _08143_ (.B1(_02639_),
    .Y(_02640_),
    .A1(net216),
    .A2(_02632_));
 sg13g2_nand3_1 _08144_ (.B(_00093_),
    .C(_02640_),
    .A(net234),
    .Y(_02641_));
 sg13g2_o21ai_1 _08145_ (.B1(_02641_),
    .Y(_02642_),
    .A1(_01259_),
    .A2(_02624_));
 sg13g2_a21oi_1 _08146_ (.A1(_01232_),
    .A2(_02642_),
    .Y(_02643_),
    .B1(\i_tinyqv.cpu.is_lui ));
 sg13g2_nand2b_1 _08147_ (.Y(_02644_),
    .B(net233),
    .A_N(_02643_));
 sg13g2_nor3_1 _08148_ (.A(_00960_),
    .B(_01100_),
    .C(_01112_),
    .Y(_02645_));
 sg13g2_buf_1 _08149_ (.A(_00920_),
    .X(_02646_));
 sg13g2_nor2_1 _08150_ (.A(net328),
    .B(_02646_),
    .Y(_02647_));
 sg13g2_nand3_1 _08151_ (.B(_02645_),
    .C(_02647_),
    .A(_01548_),
    .Y(_02648_));
 sg13g2_buf_1 _08152_ (.A(_02648_),
    .X(_02649_));
 sg13g2_buf_1 _08153_ (.A(_00915_),
    .X(_02650_));
 sg13g2_inv_1 _08154_ (.Y(_02651_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[0] ));
 sg13g2_nor3_1 _08155_ (.A(_00919_),
    .B(_01099_),
    .C(_02651_),
    .Y(_02652_));
 sg13g2_buf_1 _08156_ (.A(_01099_),
    .X(_02653_));
 sg13g2_inv_1 _08157_ (.Y(_02654_),
    .A(net255));
 sg13g2_inv_1 _08158_ (.Y(_02655_),
    .A(net256));
 sg13g2_nor3_1 _08159_ (.A(net330),
    .B(_02655_),
    .C(_02654_),
    .Y(_02656_));
 sg13g2_a21o_1 _08160_ (.A2(_02654_),
    .A1(net330),
    .B1(_02656_),
    .X(_02657_));
 sg13g2_a22oi_1 _08161_ (.Y(_02658_),
    .B1(_02657_),
    .B2(_02651_),
    .A2(_02652_),
    .A1(net256));
 sg13g2_nor3_1 _08162_ (.A(net329),
    .B(_02649_),
    .C(_02658_),
    .Y(_02659_));
 sg13g2_nor2b_1 _08163_ (.A(net329),
    .B_N(_02652_),
    .Y(_02660_));
 sg13g2_nand4_1 _08164_ (.B(_02655_),
    .C(net257),
    .A(net328),
    .Y(_02661_),
    .D(_01223_));
 sg13g2_nor4_1 _08165_ (.A(_00960_),
    .B(_01100_),
    .C(_01112_),
    .D(_02661_),
    .Y(_02662_));
 sg13g2_and2_1 _08166_ (.A(_02660_),
    .B(_02662_),
    .X(_02663_));
 sg13g2_buf_1 _08167_ (.A(_02663_),
    .X(_02664_));
 sg13g2_nor2_1 _08168_ (.A(net256),
    .B(_02649_),
    .Y(_02665_));
 sg13g2_and2_1 _08169_ (.A(_02660_),
    .B(_02665_),
    .X(_02666_));
 sg13g2_buf_1 _08170_ (.A(_02666_),
    .X(_02667_));
 sg13g2_nor3_1 _08171_ (.A(net329),
    .B(net330),
    .C(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .Y(_02668_));
 sg13g2_and3_1 _08172_ (.X(_02669_),
    .A(_02654_),
    .B(_02665_),
    .C(_02668_));
 sg13g2_buf_1 _08173_ (.A(_02669_),
    .X(_02670_));
 sg13g2_and2_1 _08174_ (.A(_02662_),
    .B(_02668_),
    .X(_02671_));
 sg13g2_buf_1 _08175_ (.A(_02671_),
    .X(_02672_));
 sg13g2_nor4_1 _08176_ (.A(_02664_),
    .B(_02667_),
    .C(_02670_),
    .D(_02672_),
    .Y(_02673_));
 sg13g2_nor2b_1 _08177_ (.A(_02659_),
    .B_N(_02673_),
    .Y(_02674_));
 sg13g2_nor3_2 _08178_ (.A(_01232_),
    .B(_01679_),
    .C(_02674_),
    .Y(_02675_));
 sg13g2_inv_1 _08179_ (.Y(_02676_),
    .A(_02649_));
 sg13g2_nand2_2 _08180_ (.Y(_02677_),
    .A(net256),
    .B(_02676_));
 sg13g2_nand2_1 _08181_ (.Y(_02678_),
    .A(_02653_),
    .B(_02668_));
 sg13g2_nand2_1 _08182_ (.Y(_02679_),
    .A(\i_tinyqv.cpu.i_core.mcause[4] ),
    .B(_01146_));
 sg13g2_nor3_1 _08183_ (.A(_02677_),
    .B(_02678_),
    .C(_02679_),
    .Y(_02680_));
 sg13g2_nor2_2 _08184_ (.A(net223),
    .B(_02398_),
    .Y(_02681_));
 sg13g2_and2_1 _08185_ (.A(_01209_),
    .B(_02681_),
    .X(_02682_));
 sg13g2_buf_1 _08186_ (.A(_02682_),
    .X(_02683_));
 sg13g2_o21ai_1 _08187_ (.B1(_02683_),
    .Y(_02684_),
    .A1(_02667_),
    .A2(_02680_));
 sg13g2_nor2_2 _08188_ (.A(_01016_),
    .B(net236),
    .Y(_02685_));
 sg13g2_nand3_1 _08189_ (.B(_02660_),
    .C(_02676_),
    .A(net256),
    .Y(_02686_));
 sg13g2_nor2_1 _08190_ (.A(_02685_),
    .B(_02686_),
    .Y(_02687_));
 sg13g2_nor3_2 _08191_ (.A(_01146_),
    .B(_02677_),
    .C(_02678_),
    .Y(_02688_));
 sg13g2_a22oi_1 _08192_ (.Y(_02689_),
    .B1(_02688_),
    .B2(\i_tinyqv.cpu.i_core.mcause[0] ),
    .A2(_02687_),
    .A1(\i_tinyqv.cpu.i_core.mepc[0] ));
 sg13g2_nor2_1 _08193_ (.A(net255),
    .B(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .Y(_02690_));
 sg13g2_a21oi_1 _08194_ (.A1(net255),
    .A2(_00170_),
    .Y(_02691_),
    .B1(_02690_));
 sg13g2_nor2_1 _08195_ (.A(net329),
    .B(_01099_),
    .Y(_02692_));
 sg13g2_nor2_2 _08196_ (.A(_01209_),
    .B(_01260_),
    .Y(_02693_));
 sg13g2_nand4_1 _08197_ (.B(_02651_),
    .C(_02692_),
    .A(net330),
    .Y(_02694_),
    .D(_02693_));
 sg13g2_buf_1 _08198_ (.A(_02694_),
    .X(_02695_));
 sg13g2_nor3_2 _08199_ (.A(_02650_),
    .B(_02649_),
    .C(_02695_),
    .Y(_02696_));
 sg13g2_a22oi_1 _08200_ (.Y(_02697_),
    .B1(_02696_),
    .B2(\i_tinyqv.cpu.i_core.mie[16] ),
    .A2(_02691_),
    .A1(_02672_));
 sg13g2_buf_1 _08201_ (.A(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .X(_02698_));
 sg13g2_nor2_2 _08202_ (.A(_02677_),
    .B(_02695_),
    .Y(_02699_));
 sg13g2_a22oi_1 _08203_ (.Y(_02700_),
    .B1(_02699_),
    .B2(_01363_),
    .A2(_02664_),
    .A1(_02698_));
 sg13g2_nand4_1 _08204_ (.B(_02689_),
    .C(_02697_),
    .A(_02684_),
    .Y(_02701_),
    .D(_02700_));
 sg13g2_nand2_1 _08205_ (.Y(_02702_),
    .A(_02675_),
    .B(_02701_));
 sg13g2_nand2_1 _08206_ (.Y(_02703_),
    .A(net233),
    .B(\i_tinyqv.cpu.is_lui ));
 sg13g2_inv_2 _08207_ (.Y(_02704_),
    .A(_02703_));
 sg13g2_a22oi_1 _08208_ (.Y(_02705_),
    .B1(_02704_),
    .B2(_01117_),
    .A2(_02702_),
    .A1(_02644_));
 sg13g2_nand2_1 _08209_ (.Y(_02706_),
    .A(net197),
    .B(_02705_));
 sg13g2_o21ai_1 _08210_ (.B1(_02706_),
    .Y(_02707_),
    .A1(net197),
    .A2(_02602_));
 sg13g2_nor2_1 _08211_ (.A(_02365_),
    .B(_02707_),
    .Y(_02708_));
 sg13g2_a21oi_1 _08212_ (.A1(_02365_),
    .A2(_02507_),
    .Y(_02709_),
    .B1(_02708_));
 sg13g2_buf_1 _08213_ (.A(_02709_),
    .X(_02710_));
 sg13g2_buf_1 _08214_ (.A(_02710_),
    .X(\debug_rd[0] ));
 sg13g2_buf_2 _08215_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .X(_02711_));
 sg13g2_buf_2 _08216_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .X(_02712_));
 sg13g2_nand2_2 _08217_ (.Y(_02713_),
    .A(_02711_),
    .B(_02712_));
 sg13g2_buf_2 _08218_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .X(_02714_));
 sg13g2_buf_1 _08219_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .X(_02715_));
 sg13g2_nand3_1 _08220_ (.B(_02715_),
    .C(_01684_),
    .A(_02714_),
    .Y(_02716_));
 sg13g2_buf_2 _08221_ (.A(_02716_),
    .X(_02717_));
 sg13g2_nor2_2 _08222_ (.A(_02713_),
    .B(_02717_),
    .Y(_02718_));
 sg13g2_mux2_1 _08223_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .A1(net80),
    .S(_02718_),
    .X(_00052_));
 sg13g2_nor2_1 _08224_ (.A(net203),
    .B(_02504_),
    .Y(_02719_));
 sg13g2_mux2_1 _08225_ (.A0(_02467_),
    .A1(_02447_),
    .S(net180),
    .X(_02720_));
 sg13g2_mux2_1 _08226_ (.A0(_02448_),
    .A1(_02460_),
    .S(net180),
    .X(_02721_));
 sg13g2_mux4_1 _08227_ (.S0(_02404_),
    .A0(_02452_),
    .A1(_02465_),
    .A2(_02720_),
    .A3(_02721_),
    .S1(net298),
    .X(_02722_));
 sg13g2_a21o_1 _08228_ (.A2(_02453_),
    .A1(_02406_),
    .B1(_02419_),
    .X(_02723_));
 sg13g2_mux2_1 _08229_ (.A0(_02454_),
    .A1(_02466_),
    .S(_02406_),
    .X(_02724_));
 sg13g2_mux4_1 _08230_ (.S0(_02404_),
    .A0(_02458_),
    .A1(_02471_),
    .A2(_02723_),
    .A3(_02724_),
    .S1(net298),
    .X(_02725_));
 sg13g2_mux2_1 _08231_ (.A0(_02722_),
    .A1(_02725_),
    .S(_02440_),
    .X(_02726_));
 sg13g2_mux2_1 _08232_ (.A0(_02726_),
    .A1(_02408_),
    .S(_02444_),
    .X(_02727_));
 sg13g2_mux2_1 _08233_ (.A0(_02383_),
    .A1(_02415_),
    .S(_02440_),
    .X(_02728_));
 sg13g2_mux4_1 _08234_ (.S0(net180),
    .A0(_02386_),
    .A1(_02394_),
    .A2(_02418_),
    .A3(_02424_),
    .S1(_02440_),
    .X(_02729_));
 sg13g2_nor2b_1 _08235_ (.A(net298),
    .B_N(_02729_),
    .Y(_02730_));
 sg13g2_a21oi_1 _08236_ (.A1(net298),
    .A2(_02728_),
    .Y(_02731_),
    .B1(_02730_));
 sg13g2_mux4_1 _08237_ (.S0(net263),
    .A0(_00202_),
    .A1(_02417_),
    .A2(_00200_),
    .A3(_02416_),
    .S1(net266),
    .X(_02732_));
 sg13g2_mux2_1 _08238_ (.A0(_02395_),
    .A1(_02732_),
    .S(net180),
    .X(_02733_));
 sg13g2_mux2_1 _08239_ (.A0(_02425_),
    .A1(_02385_),
    .S(net180),
    .X(_02734_));
 sg13g2_mux4_1 _08240_ (.S0(_02440_),
    .A0(_02733_),
    .A1(_02734_),
    .A2(_02393_),
    .A3(_02423_),
    .S1(_02397_),
    .X(_02735_));
 sg13g2_nand2_1 _08241_ (.Y(_02736_),
    .A(_02404_),
    .B(_02735_));
 sg13g2_o21ai_1 _08242_ (.B1(_02736_),
    .Y(_02737_),
    .A1(_02404_),
    .A2(_02731_));
 sg13g2_mux2_1 _08243_ (.A0(_02737_),
    .A1(_02408_),
    .S(_02444_),
    .X(_02738_));
 sg13g2_mux2_1 _08244_ (.A0(_02727_),
    .A1(_02738_),
    .S(net263),
    .X(_02739_));
 sg13g2_nand2_1 _08245_ (.Y(_02740_),
    .A(_01186_),
    .B(_02479_));
 sg13g2_o21ai_1 _08246_ (.B1(_02740_),
    .Y(_02741_),
    .A1(_01149_),
    .A2(_01185_));
 sg13g2_nand2_1 _08247_ (.Y(_02742_),
    .A(_01149_),
    .B(_01256_));
 sg13g2_nand3_1 _08248_ (.B(_01257_),
    .C(_02742_),
    .A(net187),
    .Y(_02743_));
 sg13g2_o21ai_1 _08249_ (.B1(_02743_),
    .Y(_02744_),
    .A1(net187),
    .A2(_02741_));
 sg13g2_o21ai_1 _08250_ (.B1(_02489_),
    .Y(_02745_),
    .A1(_02487_),
    .A2(_02744_));
 sg13g2_nor2b_1 _08251_ (.A(_01254_),
    .B_N(_02745_),
    .Y(_02746_));
 sg13g2_inv_1 _08252_ (.Y(_02747_),
    .A(_01076_));
 sg13g2_nand2_1 _08253_ (.Y(_02748_),
    .A(_02482_),
    .B(_02744_));
 sg13g2_nor3_1 _08254_ (.A(_02747_),
    .B(_01108_),
    .C(_02748_),
    .Y(_02749_));
 sg13g2_nand2_1 _08255_ (.Y(_02750_),
    .A(_02747_),
    .B(_01108_));
 sg13g2_a21oi_1 _08256_ (.A1(_02494_),
    .A2(_02748_),
    .Y(_02751_),
    .B1(_02750_));
 sg13g2_nor3_1 _08257_ (.A(_02746_),
    .B(_02749_),
    .C(_02751_),
    .Y(_02752_));
 sg13g2_o21ai_1 _08258_ (.B1(net115),
    .Y(_02753_),
    .A1(_01822_),
    .A2(net303));
 sg13g2_nand2_1 _08259_ (.Y(_02754_),
    .A(net115),
    .B(net130));
 sg13g2_o21ai_1 _08260_ (.B1(_01844_),
    .Y(_02755_),
    .A1(net303),
    .A2(_02754_));
 sg13g2_a22oi_1 _08261_ (.Y(_02756_),
    .B1(_02755_),
    .B2(_01822_),
    .A2(_02753_),
    .A1(net144));
 sg13g2_o21ai_1 _08262_ (.B1(net269),
    .Y(_02757_),
    .A1(_01822_),
    .A2(net144));
 sg13g2_nand3_1 _08263_ (.B(net115),
    .C(_02757_),
    .A(net303),
    .Y(_02758_));
 sg13g2_o21ai_1 _08264_ (.B1(_02758_),
    .Y(_02759_),
    .A1(_01809_),
    .A2(_02756_));
 sg13g2_xor2_1 _08265_ (.B(_02759_),
    .A(_01825_),
    .X(_02760_));
 sg13g2_nor2_1 _08266_ (.A(net198),
    .B(_02760_),
    .Y(_02761_));
 sg13g2_a21oi_1 _08267_ (.A1(net198),
    .A2(_02752_),
    .Y(_02762_),
    .B1(_02761_));
 sg13g2_nor2_1 _08268_ (.A(_02371_),
    .B(_02762_),
    .Y(_02763_));
 sg13g2_a21oi_1 _08269_ (.A1(_02371_),
    .A2(_02739_),
    .Y(_02764_),
    .B1(_02763_));
 sg13g2_or2_1 _08270_ (.X(_02765_),
    .B(_02367_),
    .A(_01174_));
 sg13g2_buf_1 _08271_ (.A(_02765_),
    .X(_02766_));
 sg13g2_nor2_1 _08272_ (.A(_02417_),
    .B(_02766_),
    .Y(_02767_));
 sg13g2_a21oi_1 _08273_ (.A1(_02719_),
    .A2(_02764_),
    .Y(_02768_),
    .B1(_02767_));
 sg13g2_buf_1 _08274_ (.A(\i_tinyqv.cpu.instr_data_in[13] ),
    .X(_02769_));
 sg13g2_mux2_1 _08275_ (.A0(_02769_),
    .A1(\i_tinyqv.mem.qspi_data_buf[13] ),
    .S(net125),
    .X(_02770_));
 sg13g2_o21ai_1 _08276_ (.B1(_02587_),
    .Y(_02771_),
    .A1(_01350_),
    .A2(_02770_));
 sg13g2_nand2_1 _08277_ (.Y(_02772_),
    .A(net236),
    .B(_02771_));
 sg13g2_buf_1 _08278_ (.A(\i_tinyqv.cpu.instr_data_in[5] ),
    .X(_02773_));
 sg13g2_mux2_1 _08279_ (.A0(_02769_),
    .A1(_02773_),
    .S(net124),
    .X(_02774_));
 sg13g2_a22oi_1 _08280_ (.Y(_02775_),
    .B1(net141),
    .B2(\i_spi.data[5] ),
    .A2(_02579_),
    .A1(\gpio_out_sel[5] ));
 sg13g2_nand2_1 _08281_ (.Y(_02776_),
    .A(_01344_),
    .B(_02543_));
 sg13g2_a221oi_1 _08282_ (.B2(\i_uart_rx.recieved_data[5] ),
    .C1(_02582_),
    .B1(net123),
    .A1(net33),
    .Y(_02777_),
    .A2(_02544_));
 sg13g2_nand3_1 _08283_ (.B(_02776_),
    .C(_02777_),
    .A(_02775_),
    .Y(_02778_));
 sg13g2_o21ai_1 _08284_ (.B1(_02778_),
    .Y(_02779_),
    .A1(_01350_),
    .A2(_02774_));
 sg13g2_nor2b_1 _08285_ (.A(_01742_),
    .B_N(\i_uart_rx.recieved_data[1] ),
    .Y(_02780_));
 sg13g2_a21oi_1 _08286_ (.A1(_01742_),
    .A2(_01374_),
    .Y(_02781_),
    .B1(_02780_));
 sg13g2_nor2_1 _08287_ (.A(_01743_),
    .B(_02781_),
    .Y(_02782_));
 sg13g2_a22oi_1 _08288_ (.Y(_02783_),
    .B1(_02549_),
    .B2(_02782_),
    .A2(_02540_),
    .A1(\i_spi.data[1] ));
 sg13g2_nor2_1 _08289_ (.A(_01741_),
    .B(_02542_),
    .Y(_02784_));
 sg13g2_a22oi_1 _08290_ (.Y(_02785_),
    .B1(_02784_),
    .B2(net3),
    .A2(_02521_),
    .A1(\gpio_out_sel[1] ));
 sg13g2_nand3_1 _08291_ (.B(_01696_),
    .C(_01709_),
    .A(net29),
    .Y(_02786_));
 sg13g2_nand4_1 _08292_ (.B(_02783_),
    .C(_02785_),
    .A(_02520_),
    .Y(_02787_),
    .D(_02786_));
 sg13g2_buf_1 _08293_ (.A(\i_tinyqv.cpu.instr_data_in[9] ),
    .X(_02788_));
 sg13g2_nor2_1 _08294_ (.A(_02788_),
    .B(_02533_),
    .Y(_02789_));
 sg13g2_a21oi_1 _08295_ (.A1(_01358_),
    .A2(_02531_),
    .Y(_02790_),
    .B1(\i_tinyqv.cpu.instr_data_in[1] ));
 sg13g2_o21ai_1 _08296_ (.B1(net276),
    .Y(_02791_),
    .A1(_02789_),
    .A2(_02790_));
 sg13g2_nand3_1 _08297_ (.B(_02787_),
    .C(_02791_),
    .A(_01144_),
    .Y(_02792_));
 sg13g2_o21ai_1 _08298_ (.B1(_02792_),
    .Y(_02793_),
    .A1(_02575_),
    .A2(_02779_));
 sg13g2_nand2b_1 _08299_ (.Y(_02794_),
    .B(_02521_),
    .A_N(_00204_));
 sg13g2_nand2b_1 _08300_ (.Y(_02795_),
    .B(_02526_),
    .A_N(\i_tinyqv.mem.qspi_data_buf[9] ));
 sg13g2_o21ai_1 _08301_ (.B1(_02795_),
    .Y(_02796_),
    .A1(_02788_),
    .A2(net125));
 sg13g2_a221oi_1 _08302_ (.B2(net230),
    .C1(_01009_),
    .B1(_02796_),
    .A1(_02520_),
    .Y(_02797_),
    .A2(_02794_));
 sg13g2_nor3_1 _08303_ (.A(_02772_),
    .B(_02793_),
    .C(_02797_),
    .Y(_02798_));
 sg13g2_and2_1 _08304_ (.A(net194),
    .B(\i_tinyqv.mem.data_from_read[21] ),
    .X(_02799_));
 sg13g2_a21oi_1 _08305_ (.A1(net223),
    .A2(\i_tinyqv.mem.data_from_read[17] ),
    .Y(_02800_),
    .B1(_02799_));
 sg13g2_mux4_1 _08306_ (.S0(net216),
    .A0(\i_tinyqv.mem.qspi_data_buf[25] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[29] ),
    .A2(_02788_),
    .A3(_02769_),
    .S1(net162),
    .X(_02801_));
 sg13g2_nand2_1 _08307_ (.Y(_02802_),
    .A(net196),
    .B(_02801_));
 sg13g2_o21ai_1 _08308_ (.B1(_02802_),
    .Y(_02803_),
    .A1(net179),
    .A2(_02800_));
 sg13g2_a21oi_1 _08309_ (.A1(net230),
    .A2(_02803_),
    .Y(_02804_),
    .B1(_02599_));
 sg13g2_nor3_1 _08310_ (.A(net156),
    .B(_02798_),
    .C(_02804_),
    .Y(_02805_));
 sg13g2_a21oi_1 _08311_ (.A1(\i_tinyqv.cpu.i_core.load_top_bit ),
    .A2(net156),
    .Y(_02806_),
    .B1(_02805_));
 sg13g2_mux2_1 _08312_ (.A0(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .A1(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .S(net174),
    .X(_02807_));
 sg13g2_buf_1 _08313_ (.A(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .X(_02808_));
 sg13g2_mux2_1 _08314_ (.A0(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .A1(_02808_),
    .S(net255),
    .X(_02809_));
 sg13g2_a22oi_1 _08315_ (.Y(_02810_),
    .B1(_02809_),
    .B2(_02672_),
    .A2(_02807_),
    .A1(_02664_));
 sg13g2_a22oi_1 _08316_ (.Y(_02811_),
    .B1(_02699_),
    .B2(_01361_),
    .A2(_02696_),
    .A1(\i_tinyqv.cpu.i_core.mie[17] ));
 sg13g2_a22oi_1 _08317_ (.Y(_02812_),
    .B1(_02688_),
    .B2(\i_tinyqv.cpu.i_core.mcause[1] ),
    .A2(_02687_),
    .A1(\i_tinyqv.cpu.i_core.mepc[1] ));
 sg13g2_nand3_1 _08318_ (.B(_02811_),
    .C(_02812_),
    .A(_02810_),
    .Y(_02813_));
 sg13g2_nand2_1 _08319_ (.Y(_02814_),
    .A(net260),
    .B(net296));
 sg13g2_nor3_1 _08320_ (.A(_02603_),
    .B(_02605_),
    .C(_02814_),
    .Y(_02815_));
 sg13g2_nand3_1 _08321_ (.B(net259),
    .C(_02815_),
    .A(net261),
    .Y(_02816_));
 sg13g2_xnor2_1 _08322_ (.Y(_02817_),
    .A(_01066_),
    .B(_02816_));
 sg13g2_nor2_1 _08323_ (.A(_02603_),
    .B(_02605_),
    .Y(_02818_));
 sg13g2_xnor2_1 _08324_ (.Y(_02819_),
    .A(net296),
    .B(_02818_));
 sg13g2_nand2_1 _08325_ (.Y(_02820_),
    .A(net261),
    .B(_02610_));
 sg13g2_nor4_2 _08326_ (.A(_02603_),
    .B(_02605_),
    .C(_02814_),
    .Y(_02821_),
    .D(_02820_));
 sg13g2_and3_1 _08327_ (.X(_02822_),
    .A(net262),
    .B(net297),
    .C(_02821_));
 sg13g2_xnor2_1 _08328_ (.Y(_02823_),
    .A(_01058_),
    .B(_02822_));
 sg13g2_mux4_1 _08329_ (.S0(net196),
    .A0(_01438_),
    .A1(_02817_),
    .A2(_02819_),
    .A3(_02823_),
    .S1(net195),
    .X(_02824_));
 sg13g2_nand4_1 _08330_ (.B(net327),
    .C(net324),
    .A(_00829_),
    .Y(_02825_),
    .D(net295));
 sg13g2_nand2_1 _08331_ (.Y(_02826_),
    .A(net334),
    .B(_01175_));
 sg13g2_nor2_1 _08332_ (.A(_02825_),
    .B(_02826_),
    .Y(_02827_));
 sg13g2_and4_1 _08333_ (.A(net262),
    .B(net326),
    .C(_01058_),
    .D(net297),
    .X(_02828_));
 sg13g2_buf_1 _08334_ (.A(_02828_),
    .X(_02829_));
 sg13g2_nor2b_1 _08335_ (.A(_02814_),
    .B_N(_02829_),
    .Y(_02830_));
 sg13g2_nand4_1 _08336_ (.B(_02610_),
    .C(_02827_),
    .A(net261),
    .Y(_02831_),
    .D(_02830_));
 sg13g2_nor3_1 _08337_ (.A(_02603_),
    .B(_02605_),
    .C(_02831_),
    .Y(_02832_));
 sg13g2_xnor2_1 _08338_ (.Y(_02833_),
    .A(net323),
    .B(_02832_));
 sg13g2_nand2_1 _08339_ (.Y(_02834_),
    .A(net258),
    .B(_02625_));
 sg13g2_nand2_1 _08340_ (.Y(_02835_),
    .A(_02821_),
    .B(_02829_));
 sg13g2_nor2_1 _08341_ (.A(_02834_),
    .B(_02835_),
    .Y(_02836_));
 sg13g2_xor2_1 _08342_ (.B(_02836_),
    .A(net324),
    .X(_02837_));
 sg13g2_nor2_1 _08343_ (.A(net194),
    .B(_02837_),
    .Y(_02838_));
 sg13g2_a21oi_1 _08344_ (.A1(net195),
    .A2(_02833_),
    .Y(_02839_),
    .B1(_02838_));
 sg13g2_a21oi_1 _08345_ (.A1(_00093_),
    .A2(_02839_),
    .Y(_02840_),
    .B1(net236));
 sg13g2_a21oi_1 _08346_ (.A1(net236),
    .A2(_02824_),
    .Y(_02841_),
    .B1(_02840_));
 sg13g2_a22oi_1 _08347_ (.Y(_02842_),
    .B1(_02841_),
    .B2(_01545_),
    .A2(_02813_),
    .A1(_02675_));
 sg13g2_nand2_1 _08348_ (.Y(_02843_),
    .A(_01106_),
    .B(_02704_));
 sg13g2_o21ai_1 _08349_ (.B1(_02843_),
    .Y(_02844_),
    .A1(_02704_),
    .A2(_02842_));
 sg13g2_nand2_1 _08350_ (.Y(_02845_),
    .A(net197),
    .B(_02844_));
 sg13g2_o21ai_1 _08351_ (.B1(_02845_),
    .Y(_02846_),
    .A1(net197),
    .A2(_02806_));
 sg13g2_nand2_1 _08352_ (.Y(_02847_),
    .A(_01671_),
    .B(_02846_));
 sg13g2_o21ai_1 _08353_ (.B1(_02847_),
    .Y(_02848_),
    .A1(_01671_),
    .A2(_02768_));
 sg13g2_buf_1 _08354_ (.A(_02848_),
    .X(_02849_));
 sg13g2_buf_1 _08355_ (.A(_02849_),
    .X(\debug_rd[1] ));
 sg13g2_mux2_1 _08356_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .A1(net76),
    .S(_02718_),
    .X(_00053_));
 sg13g2_mux2_1 _08357_ (.A0(_02738_),
    .A1(_02727_),
    .S(net263),
    .X(_02850_));
 sg13g2_xor2_1 _08358_ (.B(_01861_),
    .A(_01843_),
    .X(_02851_));
 sg13g2_xnor2_1 _08359_ (.Y(_02852_),
    .A(_00979_),
    .B(_01269_));
 sg13g2_xnor2_1 _08360_ (.Y(_02853_),
    .A(_01192_),
    .B(_02852_));
 sg13g2_or2_1 _08361_ (.X(_02854_),
    .B(_02488_),
    .A(net203));
 sg13g2_buf_1 _08362_ (.A(_02854_),
    .X(_02855_));
 sg13g2_nand2_1 _08363_ (.Y(_02856_),
    .A(_00976_),
    .B(_02494_));
 sg13g2_o21ai_1 _08364_ (.B1(_02856_),
    .Y(_02857_),
    .A1(_00976_),
    .A2(_02855_));
 sg13g2_a21oi_1 _08365_ (.A1(_00976_),
    .A2(_02855_),
    .Y(_02858_),
    .B1(_01036_));
 sg13g2_a21o_1 _08366_ (.A2(_02857_),
    .A1(_01036_),
    .B1(_02858_),
    .X(_02859_));
 sg13g2_o21ai_1 _08367_ (.B1(_02859_),
    .Y(_02860_),
    .A1(_02487_),
    .A2(_02853_));
 sg13g2_mux2_1 _08368_ (.A0(_02851_),
    .A1(_02860_),
    .S(net198),
    .X(_02861_));
 sg13g2_nor2_1 _08369_ (.A(_02371_),
    .B(_02861_),
    .Y(_02862_));
 sg13g2_a21oi_1 _08370_ (.A1(_02371_),
    .A2(_02850_),
    .Y(_02863_),
    .B1(_02862_));
 sg13g2_nor2_1 _08371_ (.A(_02416_),
    .B(_02766_),
    .Y(_02864_));
 sg13g2_a21oi_1 _08372_ (.A1(_02719_),
    .A2(_02863_),
    .Y(_02865_),
    .B1(_02864_));
 sg13g2_a21oi_1 _08373_ (.A1(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .A2(_02670_),
    .Y(_02866_),
    .B1(_02667_));
 sg13g2_mux2_1 _08374_ (.A0(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .A1(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .S(net174),
    .X(_02867_));
 sg13g2_nand2_1 _08375_ (.Y(_02868_),
    .A(_02664_),
    .B(_02867_));
 sg13g2_nand4_1 _08376_ (.B(net196),
    .C(_01259_),
    .A(net216),
    .Y(_02869_),
    .D(_02667_));
 sg13g2_buf_1 _08377_ (.A(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .X(_02870_));
 sg13g2_mux2_1 _08378_ (.A0(_02870_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .S(net255),
    .X(_02871_));
 sg13g2_a22oi_1 _08379_ (.Y(_02872_),
    .B1(_02871_),
    .B2(_02672_),
    .A2(_02696_),
    .A1(\i_tinyqv.cpu.i_core.mie[18] ));
 sg13g2_nand3_1 _08380_ (.B(_02869_),
    .C(_02872_),
    .A(_02868_),
    .Y(_02873_));
 sg13g2_a221oi_1 _08381_ (.B2(_01374_),
    .C1(_02873_),
    .B1(_02699_),
    .A1(\i_tinyqv.cpu.i_core.mepc[2] ),
    .Y(_02874_),
    .A2(_02687_));
 sg13g2_o21ai_1 _08382_ (.B1(_02874_),
    .Y(_02875_),
    .A1(net170),
    .A2(_02866_));
 sg13g2_inv_1 _08383_ (.Y(_02876_),
    .A(_01433_));
 sg13g2_nand2_1 _08384_ (.Y(_02877_),
    .A(_02613_),
    .B(_01179_));
 sg13g2_nor2_1 _08385_ (.A(_02605_),
    .B(_02877_),
    .Y(_02878_));
 sg13g2_xnor2_1 _08386_ (.Y(_02879_),
    .A(_02612_),
    .B(_02878_));
 sg13g2_nand3_1 _08387_ (.B(_02621_),
    .C(_02616_),
    .A(_01065_),
    .Y(_02880_));
 sg13g2_xor2_1 _08388_ (.B(_02880_),
    .A(_01025_),
    .X(_02881_));
 sg13g2_inv_1 _08389_ (.Y(_02882_),
    .A(_01019_));
 sg13g2_xnor2_1 _08390_ (.Y(_02883_),
    .A(_02882_),
    .B(_02630_));
 sg13g2_mux4_1 _08391_ (.S0(net194),
    .A0(_02876_),
    .A1(_02879_),
    .A2(_02881_),
    .A3(_02883_),
    .S1(_02510_),
    .X(_02884_));
 sg13g2_nand3_1 _08392_ (.B(net323),
    .C(_02827_),
    .A(_01019_),
    .Y(_02885_));
 sg13g2_nor2_1 _08393_ (.A(_02630_),
    .B(_02885_),
    .Y(_02886_));
 sg13g2_xnor2_1 _08394_ (.Y(_02887_),
    .A(_01030_),
    .B(_02886_));
 sg13g2_nor2_1 _08395_ (.A(_02634_),
    .B(_02630_),
    .Y(_02888_));
 sg13g2_xor2_1 _08396_ (.B(_02888_),
    .A(net327),
    .X(_02889_));
 sg13g2_nor2_1 _08397_ (.A(_02592_),
    .B(_02889_),
    .Y(_02890_));
 sg13g2_a21oi_1 _08398_ (.A1(_02574_),
    .A2(_02887_),
    .Y(_02891_),
    .B1(_02890_));
 sg13g2_a21oi_1 _08399_ (.A1(_00093_),
    .A2(_02891_),
    .Y(_02892_),
    .B1(_01104_));
 sg13g2_a21oi_1 _08400_ (.A1(_01104_),
    .A2(_02884_),
    .Y(_02893_),
    .B1(_02892_));
 sg13g2_a22oi_1 _08401_ (.Y(_02894_),
    .B1(_02893_),
    .B2(_01545_),
    .A2(_02875_),
    .A1(_02675_));
 sg13g2_nor2_1 _08402_ (.A(_02704_),
    .B(_02894_),
    .Y(_02895_));
 sg13g2_a21oi_1 _08403_ (.A1(_00926_),
    .A2(_02704_),
    .Y(_02896_),
    .B1(_02895_));
 sg13g2_a21oi_1 _08404_ (.A1(\i_tinyqv.cpu.i_core.load_top_bit ),
    .A2(net156),
    .Y(_02897_),
    .B1(_02508_));
 sg13g2_inv_1 _08405_ (.Y(_02898_),
    .A(\i_tinyqv.cpu.instr_data_in[14] ));
 sg13g2_buf_1 _08406_ (.A(\i_tinyqv.cpu.instr_data_in[6] ),
    .X(_02899_));
 sg13g2_nand2_1 _08407_ (.Y(_02900_),
    .A(_02899_),
    .B(net124));
 sg13g2_o21ai_1 _08408_ (.B1(_02900_),
    .Y(_02901_),
    .A1(_02898_),
    .A2(net124));
 sg13g2_nand2_1 _08409_ (.Y(_02902_),
    .A(\i_tinyqv.mem.qspi_data_buf[14] ),
    .B(net125));
 sg13g2_o21ai_1 _08410_ (.B1(_02902_),
    .Y(_02903_),
    .A1(_02898_),
    .A2(net125));
 sg13g2_buf_2 _08411_ (.A(\i_tinyqv.cpu.instr_data_in[10] ),
    .X(_02904_));
 sg13g2_buf_1 _08412_ (.A(\i_tinyqv.cpu.instr_data_in[2] ),
    .X(_02905_));
 sg13g2_mux2_1 _08413_ (.A0(_02904_),
    .A1(_02905_),
    .S(net124),
    .X(_02906_));
 sg13g2_mux2_1 _08414_ (.A0(_02904_),
    .A1(\i_tinyqv.mem.qspi_data_buf[10] ),
    .S(net125),
    .X(_02907_));
 sg13g2_mux4_1 _08415_ (.S0(net196),
    .A0(_02901_),
    .A1(_02903_),
    .A2(_02906_),
    .A3(_02907_),
    .S1(net223),
    .X(_02908_));
 sg13g2_inv_1 _08416_ (.Y(_02909_),
    .A(_02908_));
 sg13g2_a22oi_1 _08417_ (.Y(_02910_),
    .B1(_02784_),
    .B2(net4),
    .A2(_02568_),
    .A1(\i_uart_rx.recieved_data[2] ));
 sg13g2_nand3_1 _08418_ (.B(_01696_),
    .C(_01709_),
    .A(net30),
    .Y(_02911_));
 sg13g2_a22oi_1 _08419_ (.Y(_02912_),
    .B1(net141),
    .B2(\i_spi.data[2] ),
    .A2(_02521_),
    .A1(\gpio_out_sel[2] ));
 sg13g2_nand4_1 _08420_ (.B(_02910_),
    .C(_02911_),
    .A(_00924_),
    .Y(_02913_),
    .D(_02912_));
 sg13g2_mux2_1 _08421_ (.A0(net6),
    .A1(\gpio_out_sel[6] ),
    .S(net272),
    .X(_02914_));
 sg13g2_a22oi_1 _08422_ (.Y(_02915_),
    .B1(_02914_),
    .B2(net273),
    .A2(_01696_),
    .A1(net34));
 sg13g2_nor2_1 _08423_ (.A(_02541_),
    .B(_02915_),
    .Y(_02916_));
 sg13g2_a221oi_1 _08424_ (.B2(\i_uart_rx.recieved_data[6] ),
    .C1(_02916_),
    .B1(net123),
    .A1(\i_spi.data[6] ),
    .Y(_02917_),
    .A2(_02540_));
 sg13g2_a21oi_1 _08425_ (.A1(_02574_),
    .A2(_02917_),
    .Y(_02918_),
    .B1(_02591_));
 sg13g2_nand2_1 _08426_ (.Y(_02919_),
    .A(_02913_),
    .B(_02918_));
 sg13g2_a22oi_1 _08427_ (.Y(_02920_),
    .B1(_02919_),
    .B2(_02520_),
    .A2(_02909_),
    .A1(_02530_));
 sg13g2_and2_1 _08428_ (.A(net194),
    .B(\i_tinyqv.mem.data_from_read[22] ),
    .X(_02921_));
 sg13g2_a21oi_1 _08429_ (.A1(net223),
    .A2(\i_tinyqv.mem.data_from_read[18] ),
    .Y(_02922_),
    .B1(_02921_));
 sg13g2_mux4_1 _08430_ (.S0(net216),
    .A0(\i_tinyqv.mem.qspi_data_buf[26] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[30] ),
    .A2(_02904_),
    .A3(\i_tinyqv.cpu.instr_data_in[14] ),
    .S1(net162),
    .X(_02923_));
 sg13g2_nand2_1 _08431_ (.Y(_02924_),
    .A(net196),
    .B(_02923_));
 sg13g2_o21ai_1 _08432_ (.B1(_02924_),
    .Y(_02925_),
    .A1(net179),
    .A2(_02922_));
 sg13g2_a21oi_1 _08433_ (.A1(net230),
    .A2(_02925_),
    .Y(_02926_),
    .B1(_02599_));
 sg13g2_nor2_1 _08434_ (.A(_02513_),
    .B(_02926_),
    .Y(_02927_));
 sg13g2_o21ai_1 _08435_ (.B1(_02927_),
    .Y(_02928_),
    .A1(net218),
    .A2(_02920_));
 sg13g2_a22oi_1 _08436_ (.Y(_02929_),
    .B1(_02897_),
    .B2(_02928_),
    .A2(_02896_),
    .A1(_02508_));
 sg13g2_nand2_1 _08437_ (.Y(_02930_),
    .A(_01671_),
    .B(_02929_));
 sg13g2_o21ai_1 _08438_ (.B1(_02930_),
    .Y(_02931_),
    .A1(_01671_),
    .A2(_02865_));
 sg13g2_buf_1 _08439_ (.A(_02931_),
    .X(_02932_));
 sg13g2_buf_1 _08440_ (.A(_02932_),
    .X(\debug_rd[2] ));
 sg13g2_mux2_1 _08441_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .A1(net79),
    .S(_02718_),
    .X(_00054_));
 sg13g2_nor2b_1 _08442_ (.A(_01821_),
    .B_N(_01864_),
    .Y(_02933_));
 sg13g2_xnor2_1 _08443_ (.Y(_02934_),
    .A(_01884_),
    .B(_02933_));
 sg13g2_xnor2_1 _08444_ (.Y(_02935_),
    .A(_01863_),
    .B(_02934_));
 sg13g2_nand2_1 _08445_ (.Y(_02936_),
    .A(_00936_),
    .B(_01036_));
 sg13g2_nand2_1 _08446_ (.Y(_02937_),
    .A(_00936_),
    .B(_01198_));
 sg13g2_mux2_1 _08447_ (.A0(_02936_),
    .A1(_02937_),
    .S(_01192_),
    .X(_02938_));
 sg13g2_nand2_1 _08448_ (.Y(_02939_),
    .A(_00979_),
    .B(_01198_));
 sg13g2_nand2_1 _08449_ (.Y(_02940_),
    .A(_00973_),
    .B(_01036_));
 sg13g2_mux2_1 _08450_ (.A0(_02939_),
    .A1(_02940_),
    .S(_01192_),
    .X(_02941_));
 sg13g2_a21oi_1 _08451_ (.A1(_02938_),
    .A2(_02941_),
    .Y(_02942_),
    .B1(_02487_));
 sg13g2_and2_1 _08452_ (.A(_01266_),
    .B(_01268_),
    .X(_02943_));
 sg13g2_o21ai_1 _08453_ (.B1(_02943_),
    .Y(_02944_),
    .A1(_02855_),
    .A2(_02942_));
 sg13g2_nand3_1 _08454_ (.B(_02938_),
    .C(_02941_),
    .A(_02482_),
    .Y(_02945_));
 sg13g2_or2_1 _08455_ (.X(_02946_),
    .B(_02945_),
    .A(_01266_));
 sg13g2_a21o_1 _08456_ (.A2(_02945_),
    .A1(_02494_),
    .B1(_01268_),
    .X(_02947_));
 sg13g2_nand3_1 _08457_ (.B(_02946_),
    .C(_02947_),
    .A(_02944_),
    .Y(_02948_));
 sg13g2_mux2_1 _08458_ (.A0(_02935_),
    .A1(_02948_),
    .S(net198),
    .X(_02949_));
 sg13g2_mux2_1 _08459_ (.A0(_02474_),
    .A1(_02445_),
    .S(net263),
    .X(_02950_));
 sg13g2_nand2_1 _08460_ (.Y(_02951_),
    .A(_02371_),
    .B(_02950_));
 sg13g2_o21ai_1 _08461_ (.B1(_02951_),
    .Y(_02952_),
    .A1(_02371_),
    .A2(_02949_));
 sg13g2_nand2b_1 _08462_ (.Y(_02953_),
    .B(_02719_),
    .A_N(_02952_));
 sg13g2_o21ai_1 _08463_ (.B1(_02953_),
    .Y(_02954_),
    .A1(_02390_),
    .A2(_02766_));
 sg13g2_a21o_1 _08464_ (.A2(_01661_),
    .A1(_01658_),
    .B1(_01689_),
    .X(_02955_));
 sg13g2_a221oi_1 _08465_ (.B2(\i_spi.data[7] ),
    .C1(_02582_),
    .B1(net141),
    .A1(_01392_),
    .Y(_02956_),
    .A2(_02521_));
 sg13g2_a22oi_1 _08466_ (.Y(_02957_),
    .B1(_02784_),
    .B2(net7),
    .A2(net123),
    .A1(\i_uart_rx.recieved_data[7] ));
 sg13g2_and2_1 _08467_ (.A(_02956_),
    .B(_02957_),
    .X(_02958_));
 sg13g2_inv_1 _08468_ (.Y(_02959_),
    .A(_02958_));
 sg13g2_a21oi_1 _08469_ (.A1(_01428_),
    .A2(_01604_),
    .Y(_02960_),
    .B1(_02959_));
 sg13g2_buf_1 _08470_ (.A(\i_tinyqv.cpu.instr_data_in[15] ),
    .X(_02961_));
 sg13g2_buf_1 _08471_ (.A(\i_tinyqv.cpu.instr_data_in[7] ),
    .X(_02962_));
 sg13g2_mux2_1 _08472_ (.A0(_02961_),
    .A1(_02962_),
    .S(net124),
    .X(_02963_));
 sg13g2_o21ai_1 _08473_ (.B1(_02681_),
    .Y(_02964_),
    .A1(_01350_),
    .A2(_02963_));
 sg13g2_a21o_1 _08474_ (.A2(_02958_),
    .A1(_01710_),
    .B1(_02964_),
    .X(_02965_));
 sg13g2_a21oi_1 _08475_ (.A1(_02955_),
    .A2(_02960_),
    .Y(_02966_),
    .B1(_02965_));
 sg13g2_xnor2_1 _08476_ (.Y(_02967_),
    .A(_00843_),
    .B(_01572_));
 sg13g2_xnor2_1 _08477_ (.Y(_02968_),
    .A(net261),
    .B(_02815_));
 sg13g2_xnor2_1 _08478_ (.Y(_02969_),
    .A(net262),
    .B(_02821_));
 sg13g2_xor2_1 _08479_ (.B(_02835_),
    .A(net258),
    .X(_02970_));
 sg13g2_mux4_1 _08480_ (.S0(_02573_),
    .A0(_02967_),
    .A1(_02968_),
    .A2(_02969_),
    .A3(_02970_),
    .S1(_02510_),
    .X(_02971_));
 sg13g2_nor2_1 _08481_ (.A(_02825_),
    .B(_02835_),
    .Y(_02972_));
 sg13g2_xnor2_1 _08482_ (.Y(_02973_),
    .A(net334),
    .B(_02972_));
 sg13g2_nand3_1 _08483_ (.B(net323),
    .C(_02827_),
    .A(_01030_),
    .Y(_02974_));
 sg13g2_nor2_1 _08484_ (.A(_02835_),
    .B(_02974_),
    .Y(_02975_));
 sg13g2_xnor2_1 _08485_ (.Y(_02976_),
    .A(_00162_),
    .B(_02975_));
 sg13g2_nand2_1 _08486_ (.Y(_02977_),
    .A(_02573_),
    .B(_02976_));
 sg13g2_o21ai_1 _08487_ (.B1(_02977_),
    .Y(_02978_),
    .A1(_02592_),
    .A2(_02973_));
 sg13g2_nand3_1 _08488_ (.B(_00093_),
    .C(_02978_),
    .A(net234),
    .Y(_02979_));
 sg13g2_o21ai_1 _08489_ (.B1(_02979_),
    .Y(_02980_),
    .A1(net234),
    .A2(_02971_));
 sg13g2_a22oi_1 _08490_ (.Y(_02981_),
    .B1(_02683_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .A2(_01261_),
    .A1(_01385_));
 sg13g2_inv_1 _08491_ (.Y(_02982_),
    .A(_02981_));
 sg13g2_mux2_1 _08492_ (.A0(_02698_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .S(_02653_),
    .X(_02983_));
 sg13g2_a22oi_1 _08493_ (.Y(_02984_),
    .B1(_02983_),
    .B2(_02672_),
    .A2(_02982_),
    .A1(_02670_));
 sg13g2_a22oi_1 _08494_ (.Y(_02985_),
    .B1(_02699_),
    .B2(_01382_),
    .A2(_02696_),
    .A1(\i_tinyqv.cpu.i_core.mie[19] ));
 sg13g2_a22oi_1 _08495_ (.Y(_02986_),
    .B1(_02688_),
    .B2(\i_tinyqv.cpu.i_core.mcause[3] ),
    .A2(_02687_),
    .A1(\i_tinyqv.cpu.i_core.mepc[3] ));
 sg13g2_a21oi_1 _08496_ (.A1(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .A2(_02664_),
    .Y(_02987_),
    .B1(_02680_));
 sg13g2_a21oi_1 _08497_ (.A1(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .A2(_02664_),
    .Y(_02988_),
    .B1(net174));
 sg13g2_a21o_1 _08498_ (.A2(_02987_),
    .A1(net174),
    .B1(_02988_),
    .X(_02989_));
 sg13g2_nand4_1 _08499_ (.B(_02985_),
    .C(_02986_),
    .A(_02984_),
    .Y(_02990_),
    .D(_02989_));
 sg13g2_a22oi_1 _08500_ (.Y(_02991_),
    .B1(_02990_),
    .B2(_02675_),
    .A2(_02980_),
    .A1(_01545_));
 sg13g2_nand2_1 _08501_ (.Y(_02992_),
    .A(_00968_),
    .B(_02704_));
 sg13g2_o21ai_1 _08502_ (.B1(_02992_),
    .Y(_02993_),
    .A1(_02704_),
    .A2(_02991_));
 sg13g2_inv_1 _08503_ (.Y(_02994_),
    .A(\i_tinyqv.cpu.i_core.load_top_bit ));
 sg13g2_a21oi_1 _08504_ (.A1(_02994_),
    .A2(net156),
    .Y(_02995_),
    .B1(net197));
 sg13g2_a21oi_1 _08505_ (.A1(net197),
    .A2(_02993_),
    .Y(_02996_),
    .B1(_02995_));
 sg13g2_and2_1 _08506_ (.A(net195),
    .B(\i_tinyqv.mem.data_from_read[23] ),
    .X(_02997_));
 sg13g2_a21oi_1 _08507_ (.A1(net223),
    .A2(\i_tinyqv.mem.data_from_read[19] ),
    .Y(_02998_),
    .B1(_02997_));
 sg13g2_buf_1 _08508_ (.A(\i_tinyqv.cpu.instr_data_in[11] ),
    .X(_02999_));
 sg13g2_mux4_1 _08509_ (.S0(net194),
    .A0(\i_tinyqv.mem.qspi_data_buf[27] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[31] ),
    .A2(_02999_),
    .A3(_02961_),
    .S1(net162),
    .X(_03000_));
 sg13g2_nand2_1 _08510_ (.Y(_03001_),
    .A(net179),
    .B(_03000_));
 sg13g2_o21ai_1 _08511_ (.B1(_03001_),
    .Y(_03002_),
    .A1(net179),
    .A2(_02998_));
 sg13g2_a21oi_1 _08512_ (.A1(net230),
    .A2(_03002_),
    .Y(_03003_),
    .B1(_02599_));
 sg13g2_nor3_1 _08513_ (.A(_02365_),
    .B(_02996_),
    .C(_03003_),
    .Y(_03004_));
 sg13g2_o21ai_1 _08514_ (.B1(_01671_),
    .Y(_03005_),
    .A1(net197),
    .A2(net156));
 sg13g2_mux4_1 _08515_ (.S0(net194),
    .A0(_02999_),
    .A1(_02961_),
    .A2(\i_tinyqv.mem.qspi_data_buf[11] ),
    .A3(\i_tinyqv.mem.qspi_data_buf[15] ),
    .S1(_02526_),
    .X(_03006_));
 sg13g2_nand2b_1 _08516_ (.Y(_03007_),
    .B(net230),
    .A_N(_03006_));
 sg13g2_nor2_1 _08517_ (.A(net238),
    .B(_02520_),
    .Y(_03008_));
 sg13g2_and2_1 _08518_ (.A(\i_spi.data[3] ),
    .B(net141),
    .X(_03009_));
 sg13g2_a221oi_1 _08519_ (.B2(_01332_),
    .C1(_03009_),
    .B1(_02543_),
    .A1(\gpio_out_sel[3] ),
    .Y(_03010_),
    .A2(_02579_));
 sg13g2_a221oi_1 _08520_ (.B2(\i_uart_rx.recieved_data[3] ),
    .C1(_02582_),
    .B1(net123),
    .A1(net31),
    .Y(_03011_),
    .A2(_02544_));
 sg13g2_buf_1 _08521_ (.A(\i_tinyqv.cpu.instr_data_in[3] ),
    .X(_03012_));
 sg13g2_mux2_1 _08522_ (.A0(_02999_),
    .A1(_03012_),
    .S(net124),
    .X(_03013_));
 sg13g2_nor2_1 _08523_ (.A(_01350_),
    .B(_03013_),
    .Y(_03014_));
 sg13g2_a21oi_1 _08524_ (.A1(_03010_),
    .A2(_03011_),
    .Y(_03015_),
    .B1(_03014_));
 sg13g2_a221oi_1 _08525_ (.B2(_01144_),
    .C1(net218),
    .B1(_03015_),
    .A1(_03007_),
    .Y(_03016_),
    .A2(_03008_));
 sg13g2_or3_1 _08526_ (.A(_02365_),
    .B(_03003_),
    .C(_03016_),
    .X(_03017_));
 sg13g2_a21oi_1 _08527_ (.A1(_03005_),
    .A2(_03017_),
    .Y(_03018_),
    .B1(_02996_));
 sg13g2_a221oi_1 _08528_ (.B2(_03004_),
    .C1(_03018_),
    .B1(_02966_),
    .A1(_02365_),
    .Y(_03019_),
    .A2(_02954_));
 sg13g2_buf_2 _08529_ (.A(_03019_),
    .X(_03020_));
 sg13g2_buf_8 _08530_ (.A(_03020_),
    .X(_03021_));
 sg13g2_inv_1 _08531_ (.Y(\debug_rd[3] ),
    .A(net42));
 sg13g2_nor2_1 _08532_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .B(_02718_),
    .Y(_03022_));
 sg13g2_a21oi_1 _08533_ (.A1(_02718_),
    .A2(_03020_),
    .Y(_00055_),
    .B1(_03022_));
 sg13g2_nand2b_1 _08534_ (.Y(_03023_),
    .B(_02711_),
    .A_N(_02712_));
 sg13g2_buf_1 _08535_ (.A(_03023_),
    .X(_03024_));
 sg13g2_nor2_2 _08536_ (.A(_02717_),
    .B(_03024_),
    .Y(_03025_));
 sg13g2_mux2_1 _08537_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .A1(net80),
    .S(_03025_),
    .X(_00048_));
 sg13g2_mux2_1 _08538_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .A1(net76),
    .S(_03025_),
    .X(_00049_));
 sg13g2_mux2_1 _08539_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .A1(net79),
    .S(_03025_),
    .X(_00050_));
 sg13g2_nor2_1 _08540_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .B(_03025_),
    .Y(_03026_));
 sg13g2_a21oi_1 _08541_ (.A1(net42),
    .A2(_03025_),
    .Y(_00051_),
    .B1(_03026_));
 sg13g2_nand2b_1 _08542_ (.Y(_03027_),
    .B(_02712_),
    .A_N(_02711_));
 sg13g2_buf_2 _08543_ (.A(_03027_),
    .X(_03028_));
 sg13g2_nor2_2 _08544_ (.A(_02717_),
    .B(_03028_),
    .Y(_03029_));
 sg13g2_mux2_1 _08545_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .A1(net80),
    .S(_03029_),
    .X(_00044_));
 sg13g2_mux2_1 _08546_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .A1(\debug_rd[1] ),
    .S(_03029_),
    .X(_00045_));
 sg13g2_mux2_1 _08547_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .A1(net79),
    .S(_03029_),
    .X(_00046_));
 sg13g2_nor2_1 _08548_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .B(_03029_),
    .Y(_03030_));
 sg13g2_a21oi_1 _08549_ (.A1(_03021_),
    .A2(_03029_),
    .Y(_00047_),
    .B1(_03030_));
 sg13g2_nor3_2 _08550_ (.A(_02711_),
    .B(_02712_),
    .C(_02717_),
    .Y(_03031_));
 sg13g2_mux2_1 _08551_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .A1(net80),
    .S(_03031_),
    .X(_00040_));
 sg13g2_mux2_1 _08552_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .A1(net76),
    .S(_03031_),
    .X(_00041_));
 sg13g2_mux2_1 _08553_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .A1(net79),
    .S(_03031_),
    .X(_00042_));
 sg13g2_nor2_1 _08554_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .B(_03031_),
    .Y(_03032_));
 sg13g2_a21oi_1 _08555_ (.A1(_03021_),
    .A2(_03031_),
    .Y(_00043_),
    .B1(_03032_));
 sg13g2_nand3b_1 _08556_ (.B(_02715_),
    .C(_01684_),
    .Y(_03033_),
    .A_N(_02714_));
 sg13g2_buf_1 _08557_ (.A(_03033_),
    .X(_03034_));
 sg13g2_nor2_2 _08558_ (.A(_02713_),
    .B(_03034_),
    .Y(_03035_));
 sg13g2_mux2_1 _08559_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .A1(net80),
    .S(_03035_),
    .X(_00036_));
 sg13g2_mux2_1 _08560_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A1(\debug_rd[1] ),
    .S(_03035_),
    .X(_00037_));
 sg13g2_mux2_1 _08561_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .A1(\debug_rd[2] ),
    .S(_03035_),
    .X(_00038_));
 sg13g2_nor2_1 _08562_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .B(_03035_),
    .Y(_03036_));
 sg13g2_a21oi_1 _08563_ (.A1(net42),
    .A2(_03035_),
    .Y(_00039_),
    .B1(_03036_));
 sg13g2_nor2_2 _08564_ (.A(_03024_),
    .B(_03034_),
    .Y(_03037_));
 sg13g2_mux2_1 _08565_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .A1(net80),
    .S(_03037_),
    .X(_00032_));
 sg13g2_mux2_1 _08566_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .A1(net76),
    .S(_03037_),
    .X(_00033_));
 sg13g2_mux2_1 _08567_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .A1(net79),
    .S(_03037_),
    .X(_00034_));
 sg13g2_nor2_1 _08568_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .B(_03037_),
    .Y(_03038_));
 sg13g2_a21oi_1 _08569_ (.A1(net42),
    .A2(_03037_),
    .Y(_00035_),
    .B1(_03038_));
 sg13g2_nor2_2 _08570_ (.A(_03028_),
    .B(_03034_),
    .Y(_03039_));
 sg13g2_mux2_1 _08571_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .A1(_02710_),
    .S(_03039_),
    .X(_00080_));
 sg13g2_mux2_1 _08572_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .A1(_02849_),
    .S(_03039_),
    .X(_00081_));
 sg13g2_mux2_1 _08573_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .A1(_02932_),
    .S(_03039_),
    .X(_00082_));
 sg13g2_nor2_1 _08574_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .B(_03039_),
    .Y(_03040_));
 sg13g2_a21oi_1 _08575_ (.A1(net42),
    .A2(_03039_),
    .Y(_00083_),
    .B1(_03040_));
 sg13g2_or3_1 _08576_ (.A(_02711_),
    .B(_02712_),
    .C(_03034_),
    .X(_03041_));
 sg13g2_buf_2 _08577_ (.A(_03041_),
    .X(_03042_));
 sg13g2_mux2_1 _08578_ (.A0(net80),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .S(_03042_),
    .X(_00076_));
 sg13g2_mux2_1 _08579_ (.A0(net76),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .S(_03042_),
    .X(_00077_));
 sg13g2_mux2_1 _08580_ (.A0(net79),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .S(_03042_),
    .X(_00078_));
 sg13g2_nand2_1 _08581_ (.Y(_03043_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .B(_03042_));
 sg13g2_o21ai_1 _08582_ (.B1(_03043_),
    .Y(_00079_),
    .A1(_03020_),
    .A2(_03042_));
 sg13g2_nand3b_1 _08583_ (.B(_01684_),
    .C(_02714_),
    .Y(_03044_),
    .A_N(_02715_));
 sg13g2_buf_1 _08584_ (.A(_03044_),
    .X(_03045_));
 sg13g2_nor2_2 _08585_ (.A(_02713_),
    .B(_03045_),
    .Y(_03046_));
 sg13g2_mux2_1 _08586_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .A1(_02710_),
    .S(_03046_),
    .X(_00072_));
 sg13g2_mux2_1 _08587_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .A1(_02849_),
    .S(_03046_),
    .X(_00073_));
 sg13g2_mux2_1 _08588_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .A1(_02932_),
    .S(_03046_),
    .X(_00074_));
 sg13g2_nor2_1 _08589_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .B(_03046_),
    .Y(_03047_));
 sg13g2_a21oi_1 _08590_ (.A1(net42),
    .A2(_03046_),
    .Y(_00075_),
    .B1(_03047_));
 sg13g2_nor2_2 _08591_ (.A(_03024_),
    .B(_03045_),
    .Y(_03048_));
 sg13g2_mux2_1 _08592_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .A1(_02710_),
    .S(_03048_),
    .X(_00068_));
 sg13g2_mux2_1 _08593_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .A1(_02849_),
    .S(_03048_),
    .X(_00069_));
 sg13g2_mux2_1 _08594_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .A1(_02932_),
    .S(_03048_),
    .X(_00070_));
 sg13g2_nor2_1 _08595_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .B(_03048_),
    .Y(_03049_));
 sg13g2_a21oi_1 _08596_ (.A1(net42),
    .A2(_03048_),
    .Y(_00071_),
    .B1(_03049_));
 sg13g2_nor2_2 _08597_ (.A(_03028_),
    .B(_03045_),
    .Y(_03050_));
 sg13g2_mux2_1 _08598_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .A1(_02710_),
    .S(_03050_),
    .X(_00064_));
 sg13g2_mux2_1 _08599_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .A1(_02849_),
    .S(_03050_),
    .X(_00065_));
 sg13g2_mux2_1 _08600_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .A1(_02932_),
    .S(_03050_),
    .X(_00066_));
 sg13g2_nor2_1 _08601_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .B(_03050_),
    .Y(_03051_));
 sg13g2_a21oi_1 _08602_ (.A1(net42),
    .A2(_03050_),
    .Y(_00067_),
    .B1(_03051_));
 sg13g2_inv_1 _08603_ (.Y(_03052_),
    .A(_01684_));
 sg13g2_nor3_1 _08604_ (.A(_02714_),
    .B(_02715_),
    .C(_03052_),
    .Y(_03053_));
 sg13g2_nand2b_1 _08605_ (.Y(_03054_),
    .B(_03053_),
    .A_N(_03024_));
 sg13g2_buf_2 _08606_ (.A(_03054_),
    .X(_03055_));
 sg13g2_mux2_1 _08607_ (.A0(net80),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .S(_03055_),
    .X(_00060_));
 sg13g2_mux2_1 _08608_ (.A0(net76),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .S(_03055_),
    .X(_00061_));
 sg13g2_mux2_1 _08609_ (.A0(net79),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .S(_03055_),
    .X(_00062_));
 sg13g2_nand2_1 _08610_ (.Y(_03056_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .B(_03055_));
 sg13g2_o21ai_1 _08611_ (.B1(_03056_),
    .Y(_00063_),
    .A1(_03020_),
    .A2(_03055_));
 sg13g2_nand2b_1 _08612_ (.Y(_03057_),
    .B(_03053_),
    .A_N(_03028_));
 sg13g2_buf_2 _08613_ (.A(_03057_),
    .X(_03058_));
 sg13g2_mux2_1 _08614_ (.A0(\debug_rd[0] ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .S(_03058_),
    .X(_00056_));
 sg13g2_mux2_1 _08615_ (.A0(net76),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .S(_03058_),
    .X(_00057_));
 sg13g2_mux2_1 _08616_ (.A0(net79),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .S(_03058_),
    .X(_00058_));
 sg13g2_nand2_1 _08617_ (.Y(_03059_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .B(_03058_));
 sg13g2_o21ai_1 _08618_ (.B1(_03059_),
    .Y(_00059_),
    .A1(_03020_),
    .A2(_03058_));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_nand2_1 _08620_ (.Y(_03060_),
    .A(net232),
    .B(net309));
 sg13g2_o21ai_1 _08621_ (.B1(_03060_),
    .Y(_03061_),
    .A1(net232),
    .A2(net320));
 sg13g2_buf_1 _08622_ (.A(_00158_),
    .X(_03062_));
 sg13g2_buf_1 _08623_ (.A(_03062_),
    .X(_03063_));
 sg13g2_nor4_1 _08624_ (.A(net273),
    .B(net272),
    .C(_01708_),
    .D(_02516_),
    .Y(_03064_));
 sg13g2_nor2_1 _08625_ (.A(net229),
    .B(_03064_),
    .Y(_03065_));
 sg13g2_mux2_1 _08626_ (.A0(_03061_),
    .A1(net321),
    .S(_03065_),
    .X(_00233_));
 sg13g2_inv_1 _08627_ (.Y(_03066_),
    .A(\i_spi.data[0] ));
 sg13g2_xnor2_1 _08628_ (.Y(_03067_),
    .A(\i_spi.clock_divider[1] ),
    .B(\i_spi.clock_count[1] ));
 sg13g2_buf_1 _08629_ (.A(\i_spi.clock_count[0] ),
    .X(_03068_));
 sg13g2_xnor2_1 _08630_ (.Y(_03069_),
    .A(\i_spi.clock_divider[0] ),
    .B(_03068_));
 sg13g2_nand2_1 _08631_ (.Y(_03070_),
    .A(_03067_),
    .B(_03069_));
 sg13g2_buf_1 _08632_ (.A(_03070_),
    .X(_03071_));
 sg13g2_buf_1 _08633_ (.A(\i_spi.bits_remaining[3] ),
    .X(_03072_));
 sg13g2_inv_1 _08634_ (.Y(_03073_),
    .A(_03072_));
 sg13g2_a21oi_1 _08635_ (.A1(_03073_),
    .A2(\i_spi.read_latency ),
    .Y(_03074_),
    .B1(\i_spi.spi_clk_out ));
 sg13g2_buf_1 _08636_ (.A(\i_spi.busy ),
    .X(_03075_));
 sg13g2_o21ai_1 _08637_ (.B1(_03075_),
    .Y(_03076_),
    .A1(_03071_),
    .A2(_03074_));
 sg13g2_nand2b_1 _08638_ (.Y(_03077_),
    .B(_03076_),
    .A_N(_03062_));
 sg13g2_a21oi_2 _08639_ (.B1(net276),
    .Y(_03078_),
    .A2(_01301_),
    .A1(_01306_));
 sg13g2_nand2_1 _08640_ (.Y(_03079_),
    .A(_03078_),
    .B(net141));
 sg13g2_buf_1 _08641_ (.A(_03079_),
    .X(_03080_));
 sg13g2_nor3_1 _08642_ (.A(_01714_),
    .B(_03080_),
    .C(_03077_),
    .Y(_03081_));
 sg13g2_a21o_1 _08643_ (.A2(_03080_),
    .A1(_03066_),
    .B1(_03081_),
    .X(_03082_));
 sg13g2_inv_1 _08644_ (.Y(_03083_),
    .A(_03075_));
 sg13g2_buf_1 _08645_ (.A(_03083_),
    .X(_03084_));
 sg13g2_nor3_1 _08646_ (.A(_03083_),
    .B(net4),
    .C(_03077_),
    .Y(_03085_));
 sg13g2_a221oi_1 _08647_ (.B2(_03084_),
    .C1(_03085_),
    .B1(_03082_),
    .A1(_03066_),
    .Y(_00277_),
    .A2(_03077_));
 sg13g2_nand2_1 _08648_ (.Y(_03086_),
    .A(_02550_),
    .B(_03080_));
 sg13g2_o21ai_1 _08649_ (.B1(_03075_),
    .Y(_03087_),
    .A1(_01315_),
    .A2(_03071_));
 sg13g2_nand2_1 _08650_ (.Y(_03088_),
    .A(_03086_),
    .B(_03087_));
 sg13g2_or2_1 _08651_ (.X(_03089_),
    .B(_03088_),
    .A(_03062_));
 sg13g2_buf_1 _08652_ (.A(_03089_),
    .X(_03090_));
 sg13g2_buf_1 _08653_ (.A(_03090_),
    .X(_03091_));
 sg13g2_nor2_1 _08654_ (.A(_03083_),
    .B(_03066_),
    .Y(_03092_));
 sg13g2_a21oi_1 _08655_ (.A1(_03084_),
    .A2(_01718_),
    .Y(_03093_),
    .B1(_03092_));
 sg13g2_nand2_1 _08656_ (.Y(_03094_),
    .A(\i_spi.data[1] ),
    .B(net87));
 sg13g2_o21ai_1 _08657_ (.B1(_03094_),
    .Y(_00278_),
    .A1(_03091_),
    .A2(_03093_));
 sg13g2_buf_1 _08658_ (.A(_03075_),
    .X(_03095_));
 sg13g2_and2_1 _08659_ (.A(_03095_),
    .B(\i_spi.data[1] ),
    .X(_03096_));
 sg13g2_a21oi_1 _08660_ (.A1(net228),
    .A2(net307),
    .Y(_03097_),
    .B1(_03096_));
 sg13g2_nand2_1 _08661_ (.Y(_03098_),
    .A(\i_spi.data[2] ),
    .B(_03091_));
 sg13g2_o21ai_1 _08662_ (.B1(_03098_),
    .Y(_00279_),
    .A1(net87),
    .A2(_03097_));
 sg13g2_and2_1 _08663_ (.A(net254),
    .B(\i_spi.data[2] ),
    .X(_03099_));
 sg13g2_a21oi_1 _08664_ (.A1(net228),
    .A2(_01724_),
    .Y(_03100_),
    .B1(_03099_));
 sg13g2_nand2_1 _08665_ (.Y(_03101_),
    .A(\i_spi.data[3] ),
    .B(net87));
 sg13g2_o21ai_1 _08666_ (.B1(_03101_),
    .Y(_00280_),
    .A1(net87),
    .A2(_03100_));
 sg13g2_and2_1 _08667_ (.A(net254),
    .B(\i_spi.data[3] ),
    .X(_03102_));
 sg13g2_a21oi_1 _08668_ (.A1(net228),
    .A2(net306),
    .Y(_03103_),
    .B1(_03102_));
 sg13g2_nand2_1 _08669_ (.Y(_03104_),
    .A(\i_spi.data[4] ),
    .B(_03090_));
 sg13g2_o21ai_1 _08670_ (.B1(_03104_),
    .Y(_00281_),
    .A1(net87),
    .A2(_03103_));
 sg13g2_and2_1 _08671_ (.A(net254),
    .B(\i_spi.data[4] ),
    .X(_03105_));
 sg13g2_a21oi_1 _08672_ (.A1(net228),
    .A2(_01730_),
    .Y(_03106_),
    .B1(_03105_));
 sg13g2_nand2_1 _08673_ (.Y(_03107_),
    .A(\i_spi.data[5] ),
    .B(_03090_));
 sg13g2_o21ai_1 _08674_ (.B1(_03107_),
    .Y(_00282_),
    .A1(net87),
    .A2(_03106_));
 sg13g2_and2_1 _08675_ (.A(_03075_),
    .B(\i_spi.data[5] ),
    .X(_03108_));
 sg13g2_a21oi_1 _08676_ (.A1(net228),
    .A2(_01734_),
    .Y(_03109_),
    .B1(_03108_));
 sg13g2_nand2_1 _08677_ (.Y(_03110_),
    .A(\i_spi.data[6] ),
    .B(_03090_));
 sg13g2_o21ai_1 _08678_ (.B1(_03110_),
    .Y(_00283_),
    .A1(net87),
    .A2(_03109_));
 sg13g2_and2_1 _08679_ (.A(_03075_),
    .B(\i_spi.data[6] ),
    .X(_03111_));
 sg13g2_a21oi_1 _08680_ (.A1(net228),
    .A2(_01737_),
    .Y(_03112_),
    .B1(_03111_));
 sg13g2_nand2_1 _08681_ (.Y(_03113_),
    .A(\i_spi.data[7] ),
    .B(_03090_));
 sg13g2_o21ai_1 _08682_ (.B1(_03113_),
    .Y(_00284_),
    .A1(net87),
    .A2(_03112_));
 sg13g2_nand4_1 _08683_ (.B(_01691_),
    .C(_03078_),
    .A(_02550_),
    .Y(_03114_),
    .D(net141));
 sg13g2_mux2_1 _08684_ (.A0(\data_to_write[8] ),
    .A1(\i_spi.end_txn_reg ),
    .S(_03114_),
    .X(_00285_));
 sg13g2_mux2_1 _08685_ (.A0(\data_to_write[9] ),
    .A1(\i_spi.spi_dc ),
    .S(_03114_),
    .X(_00288_));
 sg13g2_xnor2_1 _08686_ (.Y(_03115_),
    .A(_01557_),
    .B(\i_tinyqv.cpu.i_core.cmp_out ));
 sg13g2_nand4_1 _08687_ (.B(net183),
    .C(_01231_),
    .A(net233),
    .Y(_03116_),
    .D(_01550_));
 sg13g2_a21oi_1 _08688_ (.A1(_00893_),
    .A2(_03115_),
    .Y(_03117_),
    .B1(_03116_));
 sg13g2_o21ai_1 _08689_ (.B1(_01770_),
    .Y(_03118_),
    .A1(net159),
    .A2(_03117_));
 sg13g2_nand2_2 _08690_ (.Y(_03119_),
    .A(_01594_),
    .B(_03118_));
 sg13g2_nor2_1 _08691_ (.A(net159),
    .B(_01326_),
    .Y(_03120_));
 sg13g2_nand2_2 _08692_ (.Y(_03121_),
    .A(_01207_),
    .B(_03120_));
 sg13g2_or2_1 _08693_ (.X(_03122_),
    .B(_03121_),
    .A(_01328_));
 sg13g2_buf_2 _08694_ (.A(_03122_),
    .X(_03123_));
 sg13g2_nand2b_1 _08695_ (.Y(_03124_),
    .B(_03123_),
    .A_N(_03119_));
 sg13g2_buf_2 _08696_ (.A(_03124_),
    .X(_03125_));
 sg13g2_nor2_1 _08697_ (.A(_01767_),
    .B(_03125_),
    .Y(_03126_));
 sg13g2_buf_1 _08698_ (.A(_03126_),
    .X(_03127_));
 sg13g2_buf_1 _08699_ (.A(net56),
    .X(_03128_));
 sg13g2_buf_1 _08700_ (.A(_01585_),
    .X(_03129_));
 sg13g2_buf_1 _08701_ (.A(_01470_),
    .X(_03130_));
 sg13g2_nand3_1 _08702_ (.B(net173),
    .C(net161),
    .A(net155),
    .Y(_03131_));
 sg13g2_inv_1 _08703_ (.Y(_03132_),
    .A(net171));
 sg13g2_nand2_1 _08704_ (.Y(_03133_),
    .A(_01468_),
    .B(_03132_));
 sg13g2_a21oi_1 _08705_ (.A1(_01481_),
    .A2(_03131_),
    .Y(_03134_),
    .B1(_03133_));
 sg13g2_nor3_2 _08706_ (.A(_01534_),
    .B(net100),
    .C(_03134_),
    .Y(_03135_));
 sg13g2_buf_1 _08707_ (.A(net135),
    .X(_03136_));
 sg13g2_nor2_1 _08708_ (.A(net171),
    .B(_01481_),
    .Y(_03137_));
 sg13g2_nor2_1 _08709_ (.A(_01468_),
    .B(_01470_),
    .Y(_03138_));
 sg13g2_a21oi_1 _08710_ (.A1(net160),
    .A2(_01463_),
    .Y(_03139_),
    .B1(_01466_));
 sg13g2_buf_1 _08711_ (.A(_03139_),
    .X(_03140_));
 sg13g2_and2_1 _08712_ (.A(_03132_),
    .B(net161),
    .X(_03141_));
 sg13g2_buf_1 _08713_ (.A(_03141_),
    .X(_03142_));
 sg13g2_nand2_1 _08714_ (.Y(_03143_),
    .A(_01480_),
    .B(_03142_));
 sg13g2_buf_1 _08715_ (.A(net160),
    .X(_03144_));
 sg13g2_mux4_1 _08716_ (.S0(net182),
    .A0(_00145_),
    .A1(_00147_),
    .A2(_00146_),
    .A3(_00144_),
    .S1(net140),
    .X(_03145_));
 sg13g2_nor4_2 _08717_ (.A(net122),
    .B(_01470_),
    .C(_03143_),
    .Y(_03146_),
    .D(_03145_));
 sg13g2_a21o_1 _08718_ (.A2(_03138_),
    .A1(_03137_),
    .B1(_03146_),
    .X(_03147_));
 sg13g2_buf_1 _08719_ (.A(_03147_),
    .X(_03148_));
 sg13g2_a21oi_1 _08720_ (.A1(net140),
    .A2(_01508_),
    .Y(_03149_),
    .B1(_01511_));
 sg13g2_buf_1 _08721_ (.A(_03149_),
    .X(_03150_));
 sg13g2_nor2_1 _08722_ (.A(net112),
    .B(_03148_),
    .Y(_03151_));
 sg13g2_a21oi_1 _08723_ (.A1(net113),
    .A2(_03148_),
    .Y(_03152_),
    .B1(_03151_));
 sg13g2_buf_1 _08724_ (.A(_01455_),
    .X(_03153_));
 sg13g2_nand2_1 _08725_ (.Y(_03154_),
    .A(net111),
    .B(_01498_));
 sg13g2_a21oi_1 _08726_ (.A1(net160),
    .A2(_01450_),
    .Y(_03155_),
    .B1(_01453_));
 sg13g2_buf_1 _08727_ (.A(_03155_),
    .X(_03156_));
 sg13g2_buf_1 _08728_ (.A(net121),
    .X(_03157_));
 sg13g2_buf_1 _08729_ (.A(_01513_),
    .X(_03158_));
 sg13g2_nand2_2 _08730_ (.Y(_03159_),
    .A(net173),
    .B(_03142_));
 sg13g2_nor2_1 _08731_ (.A(net109),
    .B(_03159_),
    .Y(_03160_));
 sg13g2_nor2_1 _08732_ (.A(net112),
    .B(_03138_),
    .Y(_03161_));
 sg13g2_mux4_1 _08733_ (.S0(net182),
    .A0(_00155_),
    .A1(_00154_),
    .A2(_00152_),
    .A3(_00153_),
    .S1(net160),
    .X(_03162_));
 sg13g2_buf_2 _08734_ (.A(_03162_),
    .X(_03163_));
 sg13g2_nor2_1 _08735_ (.A(net147),
    .B(_03163_),
    .Y(_03164_));
 sg13g2_o21ai_1 _08736_ (.B1(_03164_),
    .Y(_03165_),
    .A1(_03160_),
    .A2(_03161_));
 sg13g2_nor2_1 _08737_ (.A(_01584_),
    .B(_01529_),
    .Y(_03166_));
 sg13g2_buf_2 _08738_ (.A(_03166_),
    .X(_03167_));
 sg13g2_nand3_1 _08739_ (.B(_03165_),
    .C(_03167_),
    .A(net110),
    .Y(_03168_));
 sg13g2_nand2_1 _08740_ (.Y(_03169_),
    .A(_03154_),
    .B(_03168_));
 sg13g2_nor2_1 _08741_ (.A(net137),
    .B(_01461_),
    .Y(_03170_));
 sg13g2_a22oi_1 _08742_ (.Y(_03171_),
    .B1(_03169_),
    .B2(_03170_),
    .A2(_03152_),
    .A1(_03135_));
 sg13g2_buf_1 _08743_ (.A(net56),
    .X(_03172_));
 sg13g2_nor2_1 _08744_ (.A(net278),
    .B(net40),
    .Y(_03173_));
 sg13g2_a21oi_1 _08745_ (.A1(net41),
    .A2(_03171_),
    .Y(_00293_),
    .B1(_03173_));
 sg13g2_buf_1 _08746_ (.A(net137),
    .X(_03174_));
 sg13g2_nand2_1 _08747_ (.Y(_03175_),
    .A(_03137_),
    .B(_03138_));
 sg13g2_nor2_1 _08748_ (.A(net108),
    .B(_03175_),
    .Y(_03176_));
 sg13g2_buf_1 _08749_ (.A(_01461_),
    .X(_03177_));
 sg13g2_o21ai_1 _08750_ (.B1(_03135_),
    .Y(_03178_),
    .A1(net107),
    .A2(_03148_));
 sg13g2_nand2_2 _08751_ (.Y(_03179_),
    .A(_01584_),
    .B(_01529_));
 sg13g2_nor2_2 _08752_ (.A(net111),
    .B(_03179_),
    .Y(_03180_));
 sg13g2_a21oi_1 _08753_ (.A1(_01468_),
    .A2(net109),
    .Y(_03181_),
    .B1(_03160_));
 sg13g2_nor2_1 _08754_ (.A(net147),
    .B(_03181_),
    .Y(_03182_));
 sg13g2_nand2_1 _08755_ (.Y(_03183_),
    .A(_01462_),
    .B(_03167_));
 sg13g2_nor3_1 _08756_ (.A(_03163_),
    .B(_03182_),
    .C(_03183_),
    .Y(_03184_));
 sg13g2_a21oi_1 _08757_ (.A1(_01532_),
    .A2(_03180_),
    .Y(_03185_),
    .B1(_03184_));
 sg13g2_o21ai_1 _08758_ (.B1(_03185_),
    .Y(_03186_),
    .A1(_03176_),
    .A2(_03178_));
 sg13g2_buf_1 _08759_ (.A(net56),
    .X(_03187_));
 sg13g2_mux2_1 _08760_ (.A0(_00817_),
    .A1(_03186_),
    .S(net39),
    .X(_00294_));
 sg13g2_a21o_1 _08761_ (.A2(_01442_),
    .A1(net160),
    .B1(_01447_),
    .X(_03188_));
 sg13g2_buf_1 _08762_ (.A(_03188_),
    .X(_03189_));
 sg13g2_buf_1 _08763_ (.A(_03189_),
    .X(_03190_));
 sg13g2_mux2_1 _08764_ (.A0(_00154_),
    .A1(_00152_),
    .S(net182),
    .X(_03191_));
 sg13g2_nand2_1 _08765_ (.Y(_03192_),
    .A(_00153_),
    .B(net184));
 sg13g2_nand2_1 _08766_ (.Y(_03193_),
    .A(_00155_),
    .B(net182));
 sg13g2_a21oi_1 _08767_ (.A1(_03192_),
    .A2(_03193_),
    .Y(_03194_),
    .B1(net140));
 sg13g2_a21oi_2 _08768_ (.B1(_03194_),
    .Y(_03195_),
    .A2(_03191_),
    .A1(net140));
 sg13g2_a21oi_1 _08769_ (.A1(_03146_),
    .A2(_03195_),
    .Y(_03196_),
    .B1(_03176_));
 sg13g2_o21ai_1 _08770_ (.B1(_03196_),
    .Y(_03197_),
    .A1(net106),
    .A2(_03148_));
 sg13g2_inv_1 _08771_ (.Y(_03198_),
    .A(_01470_));
 sg13g2_nor2_1 _08772_ (.A(_03139_),
    .B(_03198_),
    .Y(_03199_));
 sg13g2_and2_1 _08773_ (.A(_01513_),
    .B(_03164_),
    .X(_03200_));
 sg13g2_buf_1 _08774_ (.A(_03200_),
    .X(_03201_));
 sg13g2_nand2_1 _08775_ (.Y(_03202_),
    .A(_03199_),
    .B(_03201_));
 sg13g2_nand2_1 _08776_ (.Y(_03203_),
    .A(_03155_),
    .B(_03170_));
 sg13g2_nand2_1 _08777_ (.Y(_03204_),
    .A(_01490_),
    .B(_01497_));
 sg13g2_buf_1 _08778_ (.A(_03204_),
    .X(_03205_));
 sg13g2_nor2_1 _08779_ (.A(_03203_),
    .B(_03205_),
    .Y(_03206_));
 sg13g2_nand2_1 _08780_ (.Y(_03207_),
    .A(net137),
    .B(net121));
 sg13g2_buf_2 _08781_ (.A(_03207_),
    .X(_03208_));
 sg13g2_nor2_1 _08782_ (.A(_03205_),
    .B(_03208_),
    .Y(_03209_));
 sg13g2_a221oi_1 _08783_ (.B2(_03206_),
    .C1(_03209_),
    .B1(_03202_),
    .A1(_03135_),
    .Y(_03210_),
    .A2(_03197_));
 sg13g2_nor2_1 _08784_ (.A(_02446_),
    .B(net40),
    .Y(_03211_));
 sg13g2_a21oi_1 _08785_ (.A1(net41),
    .A2(_03210_),
    .Y(_00295_),
    .B1(_03211_));
 sg13g2_nand2_1 _08786_ (.Y(_03212_),
    .A(net113),
    .B(net112));
 sg13g2_mux4_1 _08787_ (.S0(net182),
    .A0(_00125_),
    .A1(_00127_),
    .A2(_00126_),
    .A3(_00124_),
    .S1(net140),
    .X(_03213_));
 sg13g2_a21oi_1 _08788_ (.A1(net155),
    .A2(_03212_),
    .Y(_03214_),
    .B1(_03213_));
 sg13g2_o21ai_1 _08789_ (.B1(_03175_),
    .Y(_03215_),
    .A1(_03146_),
    .A2(_03214_));
 sg13g2_inv_1 _08790_ (.Y(_03216_),
    .A(_03215_));
 sg13g2_a21oi_1 _08791_ (.A1(_03199_),
    .A2(net109),
    .Y(_03217_),
    .B1(_03163_));
 sg13g2_nor3_1 _08792_ (.A(net147),
    .B(_03183_),
    .C(_03217_),
    .Y(_03218_));
 sg13g2_a221oi_1 _08793_ (.B2(_03135_),
    .C1(_03218_),
    .B1(_03216_),
    .A1(_01532_),
    .Y(_03219_),
    .A2(_03180_));
 sg13g2_nor2_1 _08794_ (.A(_00888_),
    .B(net40),
    .Y(_03220_));
 sg13g2_a21oi_1 _08795_ (.A1(net41),
    .A2(_03219_),
    .Y(_00296_),
    .B1(_03220_));
 sg13g2_buf_1 _08796_ (.A(_01550_),
    .X(_03221_));
 sg13g2_buf_1 _08797_ (.A(net178),
    .X(_03222_));
 sg13g2_mux2_1 _08798_ (.A0(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A1(net302),
    .S(net169),
    .X(_03223_));
 sg13g2_nor2_1 _08799_ (.A(_01767_),
    .B(_01778_),
    .Y(_03224_));
 sg13g2_buf_2 _08800_ (.A(_03224_),
    .X(_03225_));
 sg13g2_buf_1 _08801_ (.A(_03225_),
    .X(_03226_));
 sg13g2_mux2_1 _08802_ (.A0(\addr[0] ),
    .A1(_03223_),
    .S(net99),
    .X(_00300_));
 sg13g2_buf_1 _08803_ (.A(_02303_),
    .X(_03227_));
 sg13g2_buf_1 _08804_ (.A(net178),
    .X(_03228_));
 sg13g2_mux2_1 _08805_ (.A0(\i_tinyqv.cpu.i_core.mepc[10] ),
    .A1(_03227_),
    .S(net168),
    .X(_03229_));
 sg13g2_mux2_1 _08806_ (.A0(\addr[10] ),
    .A1(_03229_),
    .S(net99),
    .X(_00301_));
 sg13g2_buf_1 _08807_ (.A(_02350_),
    .X(_03230_));
 sg13g2_mux2_1 _08808_ (.A0(\i_tinyqv.cpu.i_core.mepc[11] ),
    .A1(_03230_),
    .S(net178),
    .X(_03231_));
 sg13g2_mux2_1 _08809_ (.A0(\addr[11] ),
    .A1(_03231_),
    .S(net99),
    .X(_00302_));
 sg13g2_mux2_1 _08810_ (.A0(\i_tinyqv.cpu.i_core.mepc[12] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(net178),
    .X(_03232_));
 sg13g2_mux2_1 _08811_ (.A0(\addr[12] ),
    .A1(_03232_),
    .S(net99),
    .X(_00303_));
 sg13g2_mux2_1 _08812_ (.A0(\i_tinyqv.cpu.i_core.mepc[13] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(net168),
    .X(_03233_));
 sg13g2_mux2_1 _08813_ (.A0(\addr[13] ),
    .A1(_03233_),
    .S(net99),
    .X(_00304_));
 sg13g2_mux2_1 _08814_ (.A0(\i_tinyqv.cpu.i_core.mepc[14] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .S(net168),
    .X(_03234_));
 sg13g2_mux2_1 _08815_ (.A0(\addr[14] ),
    .A1(_03234_),
    .S(net99),
    .X(_00305_));
 sg13g2_mux2_1 _08816_ (.A0(\i_tinyqv.cpu.i_core.mepc[15] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .S(net168),
    .X(_03235_));
 sg13g2_mux2_1 _08817_ (.A0(\addr[15] ),
    .A1(_03235_),
    .S(_03226_),
    .X(_00306_));
 sg13g2_mux2_1 _08818_ (.A0(\i_tinyqv.cpu.i_core.mepc[16] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .S(_03221_),
    .X(_03236_));
 sg13g2_mux2_1 _08819_ (.A0(\addr[16] ),
    .A1(_03236_),
    .S(_03226_),
    .X(_00307_));
 sg13g2_mux2_1 _08820_ (.A0(\i_tinyqv.cpu.i_core.mepc[17] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .S(net169),
    .X(_03237_));
 sg13g2_buf_1 _08821_ (.A(_03225_),
    .X(_03238_));
 sg13g2_mux2_1 _08822_ (.A0(\addr[17] ),
    .A1(_03237_),
    .S(net98),
    .X(_00308_));
 sg13g2_mux2_1 _08823_ (.A0(\i_tinyqv.cpu.i_core.mepc[18] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S(_03228_),
    .X(_03239_));
 sg13g2_mux2_1 _08824_ (.A0(\addr[18] ),
    .A1(_03239_),
    .S(net98),
    .X(_00309_));
 sg13g2_mux2_1 _08825_ (.A0(\i_tinyqv.cpu.i_core.mepc[19] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .S(_03221_),
    .X(_03240_));
 sg13g2_mux2_1 _08826_ (.A0(\addr[19] ),
    .A1(_03240_),
    .S(net98),
    .X(_00310_));
 sg13g2_mux2_1 _08827_ (.A0(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A1(_01937_),
    .S(net178),
    .X(_03241_));
 sg13g2_mux2_1 _08828_ (.A0(\addr[1] ),
    .A1(_03241_),
    .S(net98),
    .X(_00311_));
 sg13g2_mux2_1 _08829_ (.A0(\i_tinyqv.cpu.i_core.mepc[20] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .S(net168),
    .X(_03242_));
 sg13g2_mux2_1 _08830_ (.A0(\addr[20] ),
    .A1(_03242_),
    .S(net98),
    .X(_00312_));
 sg13g2_mux2_1 _08831_ (.A0(\i_tinyqv.cpu.i_core.mepc[21] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .S(net169),
    .X(_03243_));
 sg13g2_mux2_1 _08832_ (.A0(\addr[21] ),
    .A1(_03243_),
    .S(_03238_),
    .X(_00313_));
 sg13g2_mux2_1 _08833_ (.A0(\i_tinyqv.cpu.i_core.mepc[22] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .S(net178),
    .X(_03244_));
 sg13g2_mux2_1 _08834_ (.A0(\addr[22] ),
    .A1(_03244_),
    .S(net98),
    .X(_00314_));
 sg13g2_mux2_1 _08835_ (.A0(\i_tinyqv.cpu.i_core.mepc[23] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .S(_03222_),
    .X(_03245_));
 sg13g2_mux2_1 _08836_ (.A0(\addr[23] ),
    .A1(_03245_),
    .S(_03238_),
    .X(_00315_));
 sg13g2_mux2_1 _08837_ (.A0(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A1(_01996_),
    .S(net178),
    .X(_03246_));
 sg13g2_mux2_1 _08838_ (.A0(net273),
    .A1(_03246_),
    .S(net98),
    .X(_00320_));
 sg13g2_mux2_1 _08839_ (.A0(\i_tinyqv.cpu.i_core.mepc[3] ),
    .A1(_02050_),
    .S(net168),
    .X(_03247_));
 sg13g2_nand2_1 _08840_ (.Y(_03248_),
    .A(_03225_),
    .B(_03247_));
 sg13g2_o21ai_1 _08841_ (.B1(_03248_),
    .Y(_00321_),
    .A1(_02517_),
    .A2(net99));
 sg13g2_mux2_1 _08842_ (.A0(\i_tinyqv.cpu.i_core.mepc[4] ),
    .A1(_02083_),
    .S(net178),
    .X(_03249_));
 sg13g2_mux2_1 _08843_ (.A0(net310),
    .A1(_03249_),
    .S(net98),
    .X(_00322_));
 sg13g2_mux2_1 _08844_ (.A0(\i_tinyqv.cpu.i_core.mepc[5] ),
    .A1(_02137_),
    .S(net168),
    .X(_03250_));
 sg13g2_nand2_1 _08845_ (.Y(_03251_),
    .A(_03225_),
    .B(_03250_));
 sg13g2_o21ai_1 _08846_ (.B1(_03251_),
    .Y(_00323_),
    .A1(_02515_),
    .A2(net99));
 sg13g2_mux2_1 _08847_ (.A0(\i_tinyqv.cpu.i_core.mepc[6] ),
    .A1(_02168_),
    .S(_03228_),
    .X(_03252_));
 sg13g2_mux2_1 _08848_ (.A0(\addr[6] ),
    .A1(_03252_),
    .S(_03225_),
    .X(_00324_));
 sg13g2_mux2_1 _08849_ (.A0(\i_tinyqv.cpu.i_core.mepc[7] ),
    .A1(_02204_),
    .S(net169),
    .X(_03253_));
 sg13g2_mux2_1 _08850_ (.A0(\addr[7] ),
    .A1(_03253_),
    .S(_03225_),
    .X(_00325_));
 sg13g2_mux2_1 _08851_ (.A0(\i_tinyqv.cpu.i_core.mepc[8] ),
    .A1(_02248_),
    .S(net168),
    .X(_03254_));
 sg13g2_mux2_1 _08852_ (.A0(\addr[8] ),
    .A1(_03254_),
    .S(_03225_),
    .X(_00326_));
 sg13g2_mux2_1 _08853_ (.A0(\i_tinyqv.cpu.i_core.mepc[9] ),
    .A1(_02283_),
    .S(_01550_),
    .X(_03255_));
 sg13g2_mux2_1 _08854_ (.A0(\addr[9] ),
    .A1(_03255_),
    .S(_03225_),
    .X(_00327_));
 sg13g2_inv_1 _08855_ (.Y(_03256_),
    .A(net309));
 sg13g2_nand2_1 _08856_ (.Y(_03257_),
    .A(_01204_),
    .B(\i_tinyqv.cpu.no_write_in_progress ));
 sg13g2_buf_2 _08857_ (.A(_03257_),
    .X(_03258_));
 sg13g2_nor2_2 _08858_ (.A(net170),
    .B(_03258_),
    .Y(_03259_));
 sg13g2_inv_1 _08859_ (.Y(_03260_),
    .A(net156));
 sg13g2_nand2_1 _08860_ (.Y(_03261_),
    .A(_02477_),
    .B(_03260_));
 sg13g2_inv_1 _08861_ (.Y(_03262_),
    .A(_03261_));
 sg13g2_nand2_1 _08862_ (.Y(_03263_),
    .A(_03262_),
    .B(_03259_));
 sg13g2_o21ai_1 _08863_ (.B1(_03263_),
    .Y(_00328_),
    .A1(_03256_),
    .A2(_03259_));
 sg13g2_and2_1 _08864_ (.A(_00930_),
    .B(_03260_),
    .X(_03264_));
 sg13g2_buf_1 _08865_ (.A(_03264_),
    .X(_03265_));
 sg13g2_nor3_2 _08866_ (.A(net218),
    .B(_01009_),
    .C(_03258_),
    .Y(_03266_));
 sg13g2_mux2_1 _08867_ (.A0(\data_to_write[10] ),
    .A1(_03265_),
    .S(_03266_),
    .X(_00329_));
 sg13g2_and2_1 _08868_ (.A(_00959_),
    .B(_03260_),
    .X(_03267_));
 sg13g2_buf_1 _08869_ (.A(_03267_),
    .X(_03268_));
 sg13g2_mux2_1 _08870_ (.A0(\data_to_write[11] ),
    .A1(_03268_),
    .S(_03266_),
    .X(_00330_));
 sg13g2_buf_1 _08871_ (.A(net195),
    .X(_03269_));
 sg13g2_buf_1 _08872_ (.A(_01261_),
    .X(_03270_));
 sg13g2_nor2_1 _08873_ (.A(_00220_),
    .B(net167),
    .Y(_03271_));
 sg13g2_nor2b_1 _08874_ (.A(_03261_),
    .B_N(_03271_),
    .Y(_03272_));
 sg13g2_buf_1 _08875_ (.A(_03272_),
    .X(_03273_));
 sg13g2_nand2_1 _08876_ (.Y(_03274_),
    .A(net218),
    .B(_01229_));
 sg13g2_buf_2 _08877_ (.A(_03274_),
    .X(_03275_));
 sg13g2_nor2_1 _08878_ (.A(net179),
    .B(_03275_),
    .Y(_03276_));
 sg13g2_a21oi_1 _08879_ (.A1(_03273_),
    .A2(_03276_),
    .Y(_03277_),
    .B1(\data_to_write[12] ));
 sg13g2_nor3_2 _08880_ (.A(net218),
    .B(_01211_),
    .C(_03258_),
    .Y(_03278_));
 sg13g2_nor2_1 _08881_ (.A(_02514_),
    .B(_03258_),
    .Y(_03279_));
 sg13g2_nand2_1 _08882_ (.Y(_03280_),
    .A(_02591_),
    .B(_03279_));
 sg13g2_a22oi_1 _08883_ (.Y(_03281_),
    .B1(_03280_),
    .B2(\data_to_write[12] ),
    .A2(_03278_),
    .A1(_03273_));
 sg13g2_o21ai_1 _08884_ (.B1(_03281_),
    .Y(_00331_),
    .A1(_03269_),
    .A2(_03277_));
 sg13g2_nor2_2 _08885_ (.A(_01095_),
    .B(net156),
    .Y(_03282_));
 sg13g2_and2_1 _08886_ (.A(_03271_),
    .B(_03282_),
    .X(_03283_));
 sg13g2_buf_2 _08887_ (.A(_03283_),
    .X(_03284_));
 sg13g2_a21oi_1 _08888_ (.A1(_03276_),
    .A2(_03284_),
    .Y(_03285_),
    .B1(\data_to_write[13] ));
 sg13g2_a22oi_1 _08889_ (.Y(_03286_),
    .B1(_03284_),
    .B2(_03278_),
    .A2(_03280_),
    .A1(\data_to_write[13] ));
 sg13g2_o21ai_1 _08890_ (.B1(_03286_),
    .Y(_00332_),
    .A1(net177),
    .A2(_03285_));
 sg13g2_and2_1 _08891_ (.A(_03265_),
    .B(_03271_),
    .X(_03287_));
 sg13g2_buf_2 _08892_ (.A(_03287_),
    .X(_03288_));
 sg13g2_a21oi_1 _08893_ (.A1(_03276_),
    .A2(_03288_),
    .Y(_03289_),
    .B1(\data_to_write[14] ));
 sg13g2_a22oi_1 _08894_ (.Y(_03290_),
    .B1(_03288_),
    .B2(_03278_),
    .A2(_03280_),
    .A1(\data_to_write[14] ));
 sg13g2_o21ai_1 _08895_ (.B1(_03290_),
    .Y(_00333_),
    .A1(net177),
    .A2(_03289_));
 sg13g2_and2_1 _08896_ (.A(_03268_),
    .B(_03271_),
    .X(_03291_));
 sg13g2_buf_2 _08897_ (.A(_03291_),
    .X(_03292_));
 sg13g2_a21oi_1 _08898_ (.A1(_03276_),
    .A2(_03292_),
    .Y(_03293_),
    .B1(\data_to_write[15] ));
 sg13g2_a22oi_1 _08899_ (.Y(_03294_),
    .B1(_03292_),
    .B2(_03278_),
    .A2(_03280_),
    .A1(\data_to_write[15] ));
 sg13g2_o21ai_1 _08900_ (.B1(_03294_),
    .Y(_00334_),
    .A1(net177),
    .A2(_03293_));
 sg13g2_nor2_2 _08901_ (.A(_01260_),
    .B(_03275_),
    .Y(_03295_));
 sg13g2_mux2_1 _08902_ (.A0(\data_to_write[16] ),
    .A1(_03262_),
    .S(_03295_),
    .X(_00335_));
 sg13g2_mux2_1 _08903_ (.A0(\data_to_write[17] ),
    .A1(_03282_),
    .S(_03295_),
    .X(_00336_));
 sg13g2_mux2_1 _08904_ (.A0(\data_to_write[18] ),
    .A1(_03265_),
    .S(_03295_),
    .X(_00337_));
 sg13g2_mux2_1 _08905_ (.A0(\data_to_write[19] ),
    .A1(_03268_),
    .S(_03295_),
    .X(_00338_));
 sg13g2_mux2_1 _08906_ (.A0(net308),
    .A1(_03282_),
    .S(_03259_),
    .X(_00339_));
 sg13g2_nor2_1 _08907_ (.A(net238),
    .B(_03275_),
    .Y(_03296_));
 sg13g2_a21oi_1 _08908_ (.A1(_03273_),
    .A2(_03296_),
    .Y(_03297_),
    .B1(\data_to_write[20] ));
 sg13g2_nand2_1 _08909_ (.Y(_03298_),
    .A(_00848_),
    .B(_01229_));
 sg13g2_nor2_2 _08910_ (.A(_02575_),
    .B(_03275_),
    .Y(_03299_));
 sg13g2_a22oi_1 _08911_ (.Y(_03300_),
    .B1(_03299_),
    .B2(_03273_),
    .A2(_03298_),
    .A1(\data_to_write[20] ));
 sg13g2_o21ai_1 _08912_ (.B1(_03300_),
    .Y(_00340_),
    .A1(net177),
    .A2(_03297_));
 sg13g2_a21oi_1 _08913_ (.A1(_03284_),
    .A2(_03296_),
    .Y(_03301_),
    .B1(\data_to_write[21] ));
 sg13g2_a22oi_1 _08914_ (.Y(_03302_),
    .B1(_03284_),
    .B2(_03299_),
    .A2(_03298_),
    .A1(\data_to_write[21] ));
 sg13g2_o21ai_1 _08915_ (.B1(_03302_),
    .Y(_00341_),
    .A1(net177),
    .A2(_03301_));
 sg13g2_a21oi_1 _08916_ (.A1(_03288_),
    .A2(_03296_),
    .Y(_03303_),
    .B1(\data_to_write[22] ));
 sg13g2_a22oi_1 _08917_ (.Y(_03304_),
    .B1(_03288_),
    .B2(_03299_),
    .A2(_03298_),
    .A1(\data_to_write[22] ));
 sg13g2_o21ai_1 _08918_ (.B1(_03304_),
    .Y(_00342_),
    .A1(net177),
    .A2(_03303_));
 sg13g2_a21oi_1 _08919_ (.A1(_03292_),
    .A2(_03296_),
    .Y(_03305_),
    .B1(\data_to_write[23] ));
 sg13g2_a22oi_1 _08920_ (.Y(_03306_),
    .B1(_03292_),
    .B2(_03299_),
    .A2(_03298_),
    .A1(\data_to_write[23] ));
 sg13g2_o21ai_1 _08921_ (.B1(_03306_),
    .Y(_00343_),
    .A1(net177),
    .A2(_03305_));
 sg13g2_nor2_2 _08922_ (.A(_00794_),
    .B(_03258_),
    .Y(_03307_));
 sg13g2_mux2_1 _08923_ (.A0(\data_to_write[24] ),
    .A1(_03262_),
    .S(_03307_),
    .X(_00344_));
 sg13g2_mux2_1 _08924_ (.A0(\data_to_write[25] ),
    .A1(_03282_),
    .S(_03307_),
    .X(_00345_));
 sg13g2_mux2_1 _08925_ (.A0(\data_to_write[26] ),
    .A1(_03265_),
    .S(_03307_),
    .X(_00346_));
 sg13g2_mux2_1 _08926_ (.A0(\data_to_write[27] ),
    .A1(_03268_),
    .S(_03307_),
    .X(_00347_));
 sg13g2_nor2_2 _08927_ (.A(_01211_),
    .B(_03275_),
    .Y(_03308_));
 sg13g2_mux2_1 _08928_ (.A0(\data_to_write[28] ),
    .A1(_03273_),
    .S(_03308_),
    .X(_00348_));
 sg13g2_mux2_1 _08929_ (.A0(\data_to_write[29] ),
    .A1(_03284_),
    .S(_03308_),
    .X(_00349_));
 sg13g2_mux2_1 _08930_ (.A0(net307),
    .A1(_03265_),
    .S(_03259_),
    .X(_00350_));
 sg13g2_mux2_1 _08931_ (.A0(\data_to_write[30] ),
    .A1(_03288_),
    .S(_03308_),
    .X(_00351_));
 sg13g2_mux2_1 _08932_ (.A0(\data_to_write[31] ),
    .A1(_03292_),
    .S(_03308_),
    .X(_00352_));
 sg13g2_mux2_1 _08933_ (.A0(_01724_),
    .A1(_03268_),
    .S(_03259_),
    .X(_00353_));
 sg13g2_nor3_2 _08934_ (.A(net238),
    .B(_02514_),
    .C(_03258_),
    .Y(_03309_));
 sg13g2_a21oi_1 _08935_ (.A1(_03273_),
    .A2(_03309_),
    .Y(_03310_),
    .B1(net306));
 sg13g2_and2_1 _08936_ (.A(_02681_),
    .B(_03279_),
    .X(_03311_));
 sg13g2_buf_1 _08937_ (.A(_03311_),
    .X(_03312_));
 sg13g2_nand2_2 _08938_ (.Y(_03313_),
    .A(net238),
    .B(_03279_));
 sg13g2_a22oi_1 _08939_ (.Y(_03314_),
    .B1(_03313_),
    .B2(net306),
    .A2(_03312_),
    .A1(_03273_));
 sg13g2_o21ai_1 _08940_ (.B1(_03314_),
    .Y(_00354_),
    .A1(_03269_),
    .A2(_03310_));
 sg13g2_a21oi_1 _08941_ (.A1(_03309_),
    .A2(_03284_),
    .Y(_03315_),
    .B1(net305));
 sg13g2_a22oi_1 _08942_ (.Y(_03316_),
    .B1(_03313_),
    .B2(net305),
    .A2(_03312_),
    .A1(_03284_));
 sg13g2_o21ai_1 _08943_ (.B1(_03316_),
    .Y(_00355_),
    .A1(net177),
    .A2(_03315_));
 sg13g2_a21oi_1 _08944_ (.A1(_03309_),
    .A2(_03288_),
    .Y(_03317_),
    .B1(net304));
 sg13g2_a22oi_1 _08945_ (.Y(_03318_),
    .B1(_03313_),
    .B2(net304),
    .A2(_03312_),
    .A1(_03288_));
 sg13g2_o21ai_1 _08946_ (.B1(_03318_),
    .Y(_00356_),
    .A1(net195),
    .A2(_03317_));
 sg13g2_a21oi_1 _08947_ (.A1(_03309_),
    .A2(_03292_),
    .Y(_03319_),
    .B1(_01737_));
 sg13g2_a22oi_1 _08948_ (.Y(_03320_),
    .B1(_03313_),
    .B2(_01737_),
    .A2(_03312_),
    .A1(_03292_));
 sg13g2_o21ai_1 _08949_ (.B1(_03320_),
    .Y(_00357_),
    .A1(net195),
    .A2(_03319_));
 sg13g2_mux2_1 _08950_ (.A0(\data_to_write[8] ),
    .A1(_03262_),
    .S(_03266_),
    .X(_00358_));
 sg13g2_mux2_1 _08951_ (.A0(\data_to_write[9] ),
    .A1(_03282_),
    .S(_03266_),
    .X(_00359_));
 sg13g2_nor3_1 _08952_ (.A(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .B(net170),
    .C(_01225_),
    .Y(_03321_));
 sg13g2_a21o_1 _08953_ (.A2(net170),
    .A1(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .B1(_03321_),
    .X(_00378_));
 sg13g2_nor3_1 _08954_ (.A(_01767_),
    .B(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .C(_03321_),
    .Y(_03322_));
 sg13g2_nor2_1 _08955_ (.A(net236),
    .B(_02575_),
    .Y(_03323_));
 sg13g2_nand2_1 _08956_ (.Y(_03324_),
    .A(_03322_),
    .B(_03323_));
 sg13g2_mux2_1 _08957_ (.A0(\i_tinyqv.cpu.i_core.interrupt_req[0] ),
    .A1(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ),
    .S(_03324_),
    .X(_00379_));
 sg13g2_mux2_1 _08958_ (.A0(\i_tinyqv.cpu.i_core.interrupt_req[1] ),
    .A1(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ),
    .S(_03324_),
    .X(_00380_));
 sg13g2_inv_1 _08959_ (.Y(_03325_),
    .A(\i_tinyqv.cpu.i_core.load_done ));
 sg13g2_nand3_1 _08960_ (.B(\i_tinyqv.cpu.data_ready_core ),
    .C(net167),
    .A(_01774_),
    .Y(_03326_));
 sg13g2_o21ai_1 _08961_ (.B1(_03326_),
    .Y(_00381_),
    .A1(_03325_),
    .A2(net167));
 sg13g2_a21o_1 _08962_ (.A2(_02960_),
    .A1(_02955_),
    .B1(_02965_),
    .X(_03327_));
 sg13g2_a21oi_1 _08963_ (.A1(_03016_),
    .A2(_03327_),
    .Y(_03328_),
    .B1(_03003_));
 sg13g2_nor2_1 _08964_ (.A(_02509_),
    .B(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .Y(_03329_));
 sg13g2_nand3_1 _08965_ (.B(_01209_),
    .C(_03329_),
    .A(net195),
    .Y(_03330_));
 sg13g2_xor2_1 _08966_ (.B(_01556_),
    .A(net179),
    .X(_03331_));
 sg13g2_nor3_1 _08967_ (.A(net197),
    .B(_03330_),
    .C(_03331_),
    .Y(_03332_));
 sg13g2_nor3_1 _08968_ (.A(_02994_),
    .B(net167),
    .C(_03332_),
    .Y(_03333_));
 sg13g2_a21o_1 _08969_ (.A2(_03332_),
    .A1(_03328_),
    .B1(_03333_),
    .X(_00382_));
 sg13g2_nand2_1 _08970_ (.Y(_03334_),
    .A(net233),
    .B(\i_tinyqv.cpu.is_alu_imm ));
 sg13g2_buf_2 _08971_ (.A(_03334_),
    .X(_03335_));
 sg13g2_nand2_1 _08972_ (.Y(_03336_),
    .A(_02477_),
    .B(_03335_));
 sg13g2_o21ai_1 _08973_ (.B1(_03336_),
    .Y(_03337_),
    .A1(_01117_),
    .A2(_03335_));
 sg13g2_nand2_1 _08974_ (.Y(_03338_),
    .A(net167),
    .B(_01775_));
 sg13g2_buf_2 _08975_ (.A(_03338_),
    .X(_03339_));
 sg13g2_mux2_1 _08976_ (.A0(_03337_),
    .A1(net266),
    .S(_03339_),
    .X(_00418_));
 sg13g2_nand2_1 _08977_ (.Y(_03340_),
    .A(_01095_),
    .B(_03335_));
 sg13g2_o21ai_1 _08978_ (.B1(_03340_),
    .Y(_03341_),
    .A1(_01106_),
    .A2(_03335_));
 sg13g2_nand2_1 _08979_ (.Y(_03342_),
    .A(_02397_),
    .B(_03339_));
 sg13g2_o21ai_1 _08980_ (.B1(_03342_),
    .Y(_00419_),
    .A1(_03339_),
    .A2(_03341_));
 sg13g2_nor2b_1 _08981_ (.A(_03335_),
    .B_N(_00926_),
    .Y(_03343_));
 sg13g2_a21oi_1 _08982_ (.A1(_00930_),
    .A2(_03335_),
    .Y(_03344_),
    .B1(_03343_));
 sg13g2_nand2_1 _08983_ (.Y(_03345_),
    .A(_02378_),
    .B(_03339_));
 sg13g2_o21ai_1 _08984_ (.B1(_03345_),
    .Y(_00420_),
    .A1(_03339_),
    .A2(_03344_));
 sg13g2_nor2b_1 _08985_ (.A(_03335_),
    .B_N(_00968_),
    .Y(_03346_));
 sg13g2_a21oi_1 _08986_ (.A1(_00959_),
    .A2(_03335_),
    .Y(_03347_),
    .B1(_03346_));
 sg13g2_nand2_1 _08987_ (.Y(_03348_),
    .A(_02399_),
    .B(_03339_));
 sg13g2_o21ai_1 _08988_ (.B1(_03348_),
    .Y(_00421_),
    .A1(_03339_),
    .A2(_03347_));
 sg13g2_nor4_1 _08989_ (.A(net218),
    .B(net270),
    .C(_01774_),
    .D(_02575_),
    .Y(_03349_));
 sg13g2_mux2_1 _08990_ (.A0(_02428_),
    .A1(_03337_),
    .S(_03349_),
    .X(_00422_));
 sg13g2_buf_1 _08991_ (.A(_01490_),
    .X(_03350_));
 sg13g2_buf_1 _08992_ (.A(_01529_),
    .X(_03351_));
 sg13g2_nor2_1 _08993_ (.A(net105),
    .B(net104),
    .Y(_03352_));
 sg13g2_nand3_1 _08994_ (.B(net173),
    .C(_03142_),
    .A(_01468_),
    .Y(_03353_));
 sg13g2_buf_1 _08995_ (.A(_03353_),
    .X(_03354_));
 sg13g2_nand2_1 _08996_ (.Y(_03355_),
    .A(_03352_),
    .B(_03354_));
 sg13g2_buf_1 _08997_ (.A(_03355_),
    .X(_03356_));
 sg13g2_nor3_2 _08998_ (.A(_03140_),
    .B(_01470_),
    .C(_01483_),
    .Y(_03357_));
 sg13g2_nor2_1 _08999_ (.A(_03130_),
    .B(_01483_),
    .Y(_03358_));
 sg13g2_buf_2 _09000_ (.A(_03358_),
    .X(_03359_));
 sg13g2_mux4_1 _09001_ (.S0(net182),
    .A0(_00109_),
    .A1(_00111_),
    .A2(_00110_),
    .A3(_00108_),
    .S1(net140),
    .X(_03360_));
 sg13g2_nor2_1 _09002_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sg13g2_a22oi_1 _09003_ (.Y(_03362_),
    .B1(_03361_),
    .B2(_01536_),
    .A2(_03357_),
    .A1(net136));
 sg13g2_nor2_1 _09004_ (.A(_03356_),
    .B(_03362_),
    .Y(_03363_));
 sg13g2_nand3_1 _09005_ (.B(_03164_),
    .C(_03206_),
    .A(_03149_),
    .Y(_03364_));
 sg13g2_buf_1 _09006_ (.A(_03364_),
    .X(_03365_));
 sg13g2_o21ai_1 _09007_ (.B1(_03205_),
    .Y(_03366_),
    .A1(net137),
    .A2(_03179_));
 sg13g2_nand2_1 _09008_ (.Y(_03367_),
    .A(net111),
    .B(_03366_));
 sg13g2_o21ai_1 _09009_ (.B1(_03367_),
    .Y(_03368_),
    .A1(_01449_),
    .A2(_03205_));
 sg13g2_nand3_1 _09010_ (.B(net173),
    .C(_03368_),
    .A(net113),
    .Y(_03369_));
 sg13g2_buf_1 _09011_ (.A(net104),
    .X(_03370_));
 sg13g2_buf_1 _09012_ (.A(net105),
    .X(_03371_));
 sg13g2_nor2_1 _09013_ (.A(_01506_),
    .B(net136),
    .Y(_03372_));
 sg13g2_nand3_1 _09014_ (.B(_03163_),
    .C(_03372_),
    .A(_01519_),
    .Y(_03373_));
 sg13g2_nand3_1 _09015_ (.B(net105),
    .C(net147),
    .A(net122),
    .Y(_03374_));
 sg13g2_o21ai_1 _09016_ (.B1(_03374_),
    .Y(_03375_),
    .A1(net96),
    .A2(_03373_));
 sg13g2_nand3_1 _09017_ (.B(net97),
    .C(_03375_),
    .A(_01462_),
    .Y(_03376_));
 sg13g2_nand3_1 _09018_ (.B(_03369_),
    .C(_03376_),
    .A(_03365_),
    .Y(_03377_));
 sg13g2_buf_1 _09019_ (.A(_03126_),
    .X(_03378_));
 sg13g2_o21ai_1 _09020_ (.B1(net55),
    .Y(_03379_),
    .A1(_03363_),
    .A2(_03377_));
 sg13g2_o21ai_1 _09021_ (.B1(_03379_),
    .Y(_00458_),
    .A1(_02651_),
    .A2(net39));
 sg13g2_nand2_1 _09022_ (.Y(_03380_),
    .A(net171),
    .B(_03167_));
 sg13g2_a21oi_1 _09023_ (.A1(_03367_),
    .A2(_03380_),
    .Y(_03381_),
    .B1(net107));
 sg13g2_a21oi_1 _09024_ (.A1(_03164_),
    .A2(_03159_),
    .Y(_03382_),
    .B1(_03183_));
 sg13g2_nor3_1 _09025_ (.A(_03209_),
    .B(_03381_),
    .C(_03382_),
    .Y(_03383_));
 sg13g2_nor2_1 _09026_ (.A(net109),
    .B(_03383_),
    .Y(_03384_));
 sg13g2_nand2_2 _09027_ (.Y(_03385_),
    .A(_01490_),
    .B(_01529_));
 sg13g2_nand2_1 _09028_ (.Y(_03386_),
    .A(net137),
    .B(_01461_));
 sg13g2_buf_2 _09029_ (.A(_03386_),
    .X(_03387_));
 sg13g2_nor3_1 _09030_ (.A(net111),
    .B(_03385_),
    .C(_03387_),
    .Y(_03388_));
 sg13g2_buf_1 _09031_ (.A(_03388_),
    .X(_03389_));
 sg13g2_nor3_1 _09032_ (.A(_03156_),
    .B(_03205_),
    .C(_03387_),
    .Y(_03390_));
 sg13g2_nor3_1 _09033_ (.A(_01506_),
    .B(_01519_),
    .C(net136),
    .Y(_03391_));
 sg13g2_and2_1 _09034_ (.A(_03390_),
    .B(_03391_),
    .X(_03392_));
 sg13g2_nand2_2 _09035_ (.Y(_03393_),
    .A(_03189_),
    .B(_01461_));
 sg13g2_nor2_2 _09036_ (.A(_03393_),
    .B(_03154_),
    .Y(_03394_));
 sg13g2_or2_1 _09037_ (.X(_03395_),
    .B(_03394_),
    .A(_03392_));
 sg13g2_buf_1 _09038_ (.A(_03395_),
    .X(_03396_));
 sg13g2_o21ai_1 _09039_ (.B1(net112),
    .Y(_03397_),
    .A1(net89),
    .A2(_03396_));
 sg13g2_nor2b_1 _09040_ (.A(_03384_),
    .B_N(_03397_),
    .Y(_03398_));
 sg13g2_or2_1 _09041_ (.X(_03399_),
    .B(net90),
    .A(_03213_));
 sg13g2_buf_1 _09042_ (.A(net140),
    .X(_03400_));
 sg13g2_a21oi_1 _09043_ (.A1(net120),
    .A2(_01514_),
    .Y(_03401_),
    .B1(_01517_));
 sg13g2_nand3_1 _09044_ (.B(_01532_),
    .C(_03167_),
    .A(_03401_),
    .Y(_03402_));
 sg13g2_nand3_1 _09045_ (.B(_03399_),
    .C(_03402_),
    .A(_03398_),
    .Y(_03403_));
 sg13g2_buf_1 _09046_ (.A(net56),
    .X(_03404_));
 sg13g2_mux2_1 _09047_ (.A0(net257),
    .A1(_03403_),
    .S(_03404_),
    .X(_00459_));
 sg13g2_nor2_1 _09048_ (.A(_03153_),
    .B(_03387_),
    .Y(_03405_));
 sg13g2_o21ai_1 _09049_ (.B1(_03203_),
    .Y(_03406_),
    .A1(net121),
    .A2(_03387_));
 sg13g2_nor2_1 _09050_ (.A(_01529_),
    .B(_03406_),
    .Y(_03407_));
 sg13g2_o21ai_1 _09051_ (.B1(_01490_),
    .Y(_03408_),
    .A1(_03405_),
    .A2(_03407_));
 sg13g2_nor2_1 _09052_ (.A(net137),
    .B(net121),
    .Y(_03409_));
 sg13g2_nand2_1 _09053_ (.Y(_03410_),
    .A(_01498_),
    .B(_03409_));
 sg13g2_nand3b_1 _09054_ (.B(_03408_),
    .C(_03410_),
    .Y(_03411_),
    .A_N(_03382_));
 sg13g2_or2_1 _09055_ (.X(_03412_),
    .B(_03411_),
    .A(_03392_));
 sg13g2_a21oi_1 _09056_ (.A1(net171),
    .A2(_03206_),
    .Y(_03413_),
    .B1(_03412_));
 sg13g2_nor2_1 _09057_ (.A(net109),
    .B(_03413_),
    .Y(_03414_));
 sg13g2_mux4_1 _09058_ (.S0(_01587_),
    .A0(_00129_),
    .A1(_00131_),
    .A2(_00130_),
    .A3(_00128_),
    .S1(_03144_),
    .X(_03415_));
 sg13g2_buf_1 _09059_ (.A(_03415_),
    .X(_03416_));
 sg13g2_nor2b_1 _09060_ (.A(_01536_),
    .B_N(_03360_),
    .Y(_03417_));
 sg13g2_a21oi_1 _09061_ (.A1(_01536_),
    .A2(_03416_),
    .Y(_03418_),
    .B1(_03417_));
 sg13g2_nor2_1 _09062_ (.A(_03140_),
    .B(_03159_),
    .Y(_03419_));
 sg13g2_nor2_1 _09063_ (.A(_01585_),
    .B(_03419_),
    .Y(_03420_));
 sg13g2_o21ai_1 _09064_ (.B1(_03420_),
    .Y(_03421_),
    .A1(net136),
    .A2(_03175_));
 sg13g2_a21oi_1 _09065_ (.A1(_03357_),
    .A2(_03416_),
    .Y(_03422_),
    .B1(_03421_));
 sg13g2_o21ai_1 _09066_ (.B1(_03422_),
    .Y(_03423_),
    .A1(_03359_),
    .A2(_03418_));
 sg13g2_nor2b_1 _09067_ (.A(_03414_),
    .B_N(_03423_),
    .Y(_03424_));
 sg13g2_nor2_1 _09068_ (.A(net328),
    .B(_03172_),
    .Y(_03425_));
 sg13g2_a21oi_1 _09069_ (.A1(_03128_),
    .A2(_03424_),
    .Y(_00460_),
    .B1(_03425_));
 sg13g2_nor2b_1 _09070_ (.A(_03391_),
    .B_N(_03390_),
    .Y(_03426_));
 sg13g2_buf_1 _09071_ (.A(_03426_),
    .X(_03427_));
 sg13g2_and2_1 _09072_ (.A(_01536_),
    .B(_03354_),
    .X(_03428_));
 sg13g2_buf_1 _09073_ (.A(_03428_),
    .X(_03429_));
 sg13g2_a21oi_1 _09074_ (.A1(_03416_),
    .A2(_03429_),
    .Y(_03430_),
    .B1(net100));
 sg13g2_buf_2 _09075_ (.A(_03430_),
    .X(_03431_));
 sg13g2_nand2_1 _09076_ (.Y(_03432_),
    .A(_01536_),
    .B(_03354_));
 sg13g2_nand2_1 _09077_ (.Y(_03433_),
    .A(net109),
    .B(_03432_));
 sg13g2_a221oi_1 _09078_ (.B2(_03433_),
    .C1(_03414_),
    .B1(_03431_),
    .A1(net173),
    .Y(_03434_),
    .A2(_03427_));
 sg13g2_nor2_1 _09079_ (.A(_01113_),
    .B(net40),
    .Y(_03435_));
 sg13g2_a21oi_1 _09080_ (.A1(net41),
    .A2(_03434_),
    .Y(_00461_),
    .B1(_03435_));
 sg13g2_nand2_1 _09081_ (.Y(_03436_),
    .A(net113),
    .B(_03432_));
 sg13g2_a221oi_1 _09082_ (.B2(_03436_),
    .C1(_03414_),
    .B1(_03431_),
    .A1(_01533_),
    .Y(_03437_),
    .A2(_03427_));
 sg13g2_nor2_1 _09083_ (.A(_01102_),
    .B(_03172_),
    .Y(_03438_));
 sg13g2_a21oi_1 _09084_ (.A1(_03128_),
    .A2(_03437_),
    .Y(_00462_),
    .B1(_03438_));
 sg13g2_nand2_1 _09085_ (.Y(_03439_),
    .A(net106),
    .B(_03432_));
 sg13g2_a221oi_1 _09086_ (.B2(_03439_),
    .C1(_03414_),
    .B1(_03431_),
    .A1(_01477_),
    .Y(_03440_),
    .A2(_03427_));
 sg13g2_buf_1 _09087_ (.A(net56),
    .X(_03441_));
 sg13g2_nor2_1 _09088_ (.A(_00916_),
    .B(net37),
    .Y(_03442_));
 sg13g2_a21oi_1 _09089_ (.A1(net41),
    .A2(_03440_),
    .Y(_00463_),
    .B1(_03442_));
 sg13g2_buf_1 _09090_ (.A(net111),
    .X(_03443_));
 sg13g2_nand2_1 _09091_ (.Y(_03444_),
    .A(net95),
    .B(_03432_));
 sg13g2_a221oi_1 _09092_ (.B2(_03444_),
    .C1(_03414_),
    .B1(_03431_),
    .A1(_03198_),
    .Y(_03445_),
    .A2(_03427_));
 sg13g2_nor2_1 _09093_ (.A(_00961_),
    .B(net37),
    .Y(_03446_));
 sg13g2_a21oi_1 _09094_ (.A1(net41),
    .A2(_03445_),
    .Y(_00464_),
    .B1(_03446_));
 sg13g2_buf_2 _09095_ (.A(net182),
    .X(_03447_));
 sg13g2_mux4_1 _09096_ (.S0(_03447_),
    .A0(\i_tinyqv.cpu.instr_data[0][0] ),
    .A1(\i_tinyqv.cpu.instr_data[3][0] ),
    .A2(\i_tinyqv.cpu.instr_data[2][0] ),
    .A3(\i_tinyqv.cpu.instr_data[1][0] ),
    .S1(net120),
    .X(_03448_));
 sg13g2_o21ai_1 _09097_ (.B1(_03431_),
    .Y(_03449_),
    .A1(_03429_),
    .A2(_03448_));
 sg13g2_inv_1 _09098_ (.Y(_03450_),
    .A(_03449_));
 sg13g2_a221oi_1 _09099_ (.B2(net122),
    .C1(_03450_),
    .B1(_03427_),
    .A1(net112),
    .Y(_03451_),
    .A2(_03412_));
 sg13g2_nor2_1 _09100_ (.A(_01109_),
    .B(_03441_),
    .Y(_03452_));
 sg13g2_a21oi_1 _09101_ (.A1(net41),
    .A2(_03451_),
    .Y(_00465_),
    .B1(_03452_));
 sg13g2_nor2_1 _09102_ (.A(_03390_),
    .B(_03411_),
    .Y(_03453_));
 sg13g2_nor2_2 _09103_ (.A(net109),
    .B(_03453_),
    .Y(_03454_));
 sg13g2_mux4_1 _09104_ (.S0(_03144_),
    .A0(\i_tinyqv.cpu.instr_data[0][1] ),
    .A1(\i_tinyqv.cpu.instr_data[2][1] ),
    .A2(\i_tinyqv.cpu.instr_data[3][1] ),
    .A3(\i_tinyqv.cpu.instr_data[1][1] ),
    .S1(net166),
    .X(_03455_));
 sg13g2_o21ai_1 _09105_ (.B1(_03431_),
    .Y(_03456_),
    .A1(_03429_),
    .A2(_03455_));
 sg13g2_nor2b_1 _09106_ (.A(_03454_),
    .B_N(_03456_),
    .Y(_03457_));
 sg13g2_nor2_1 _09107_ (.A(_01096_),
    .B(net37),
    .Y(_03458_));
 sg13g2_a21oi_1 _09108_ (.A1(net41),
    .A2(_03457_),
    .Y(_00466_),
    .B1(_03458_));
 sg13g2_buf_1 _09109_ (.A(net56),
    .X(_03459_));
 sg13g2_mux4_1 _09110_ (.S0(net166),
    .A0(\i_tinyqv.cpu.instr_data[0][2] ),
    .A1(\i_tinyqv.cpu.instr_data[3][2] ),
    .A2(\i_tinyqv.cpu.instr_data[2][2] ),
    .A3(\i_tinyqv.cpu.instr_data[1][2] ),
    .S1(net120),
    .X(_03460_));
 sg13g2_o21ai_1 _09111_ (.B1(_03431_),
    .Y(_03461_),
    .A1(_03429_),
    .A2(_03460_));
 sg13g2_nor2b_1 _09112_ (.A(_03454_),
    .B_N(_03461_),
    .Y(_03462_));
 sg13g2_nor2_1 _09113_ (.A(_00921_),
    .B(net37),
    .Y(_03463_));
 sg13g2_a21oi_1 _09114_ (.A1(net36),
    .A2(_03462_),
    .Y(_00467_),
    .B1(_03463_));
 sg13g2_mux4_1 _09115_ (.S0(net166),
    .A0(\i_tinyqv.cpu.instr_data[0][3] ),
    .A1(\i_tinyqv.cpu.instr_data[3][3] ),
    .A2(\i_tinyqv.cpu.instr_data[2][3] ),
    .A3(\i_tinyqv.cpu.instr_data[1][3] ),
    .S1(net120),
    .X(_03464_));
 sg13g2_o21ai_1 _09116_ (.B1(_03431_),
    .Y(_03465_),
    .A1(_03429_),
    .A2(_03464_));
 sg13g2_nor2b_1 _09117_ (.A(_03454_),
    .B_N(_03465_),
    .Y(_03466_));
 sg13g2_nor2_1 _09118_ (.A(_00965_),
    .B(_03441_),
    .Y(_03467_));
 sg13g2_a21oi_1 _09119_ (.A1(_03459_),
    .A2(_03466_),
    .Y(_00468_),
    .B1(_03467_));
 sg13g2_mux4_1 _09120_ (.S0(net182),
    .A0(_00113_),
    .A1(_00115_),
    .A2(_00114_),
    .A3(_00112_),
    .S1(net140),
    .X(_03468_));
 sg13g2_nor2b_1 _09121_ (.A(_03359_),
    .B_N(_03468_),
    .Y(_03469_));
 sg13g2_a21oi_1 _09122_ (.A1(_01519_),
    .A2(_03359_),
    .Y(_03470_),
    .B1(_03469_));
 sg13g2_nand2_1 _09123_ (.Y(_03471_),
    .A(net135),
    .B(_03368_));
 sg13g2_a21oi_1 _09124_ (.A1(_03393_),
    .A2(_03208_),
    .Y(_03472_),
    .B1(_03205_));
 sg13g2_inv_1 _09125_ (.Y(_03473_),
    .A(_03472_));
 sg13g2_a22oi_1 _09126_ (.Y(_03474_),
    .B1(_03471_),
    .B2(_03473_),
    .A2(_03365_),
    .A1(_03132_));
 sg13g2_nor3_1 _09127_ (.A(_03203_),
    .B(net155),
    .C(_03385_),
    .Y(_03475_));
 sg13g2_nor2_1 _09128_ (.A(_03474_),
    .B(_03475_),
    .Y(_03476_));
 sg13g2_o21ai_1 _09129_ (.B1(_03476_),
    .Y(_03477_),
    .A1(_03443_),
    .A2(_03393_));
 sg13g2_nand3_1 _09130_ (.B(net107),
    .C(net97),
    .A(_03443_),
    .Y(_03478_));
 sg13g2_buf_1 _09131_ (.A(_01584_),
    .X(_03479_));
 sg13g2_a21oi_1 _09132_ (.A1(_03476_),
    .A2(_03478_),
    .Y(_03480_),
    .B1(net103));
 sg13g2_a221oi_1 _09133_ (.B2(net97),
    .C1(_03480_),
    .B1(_03477_),
    .A1(_03420_),
    .Y(_03481_),
    .A2(_03470_));
 sg13g2_nor2_1 _09134_ (.A(net255),
    .B(net37),
    .Y(_03482_));
 sg13g2_a21oi_1 _09135_ (.A1(net36),
    .A2(_03481_),
    .Y(_00469_),
    .B1(_03482_));
 sg13g2_buf_1 _09136_ (.A(_03352_),
    .X(_03483_));
 sg13g2_nand2_1 _09137_ (.Y(_03484_),
    .A(_03483_),
    .B(_03419_));
 sg13g2_buf_1 _09138_ (.A(_03484_),
    .X(_03485_));
 sg13g2_nor2_1 _09139_ (.A(net90),
    .B(_03416_),
    .Y(_03486_));
 sg13g2_nor2_1 _09140_ (.A(_03454_),
    .B(_03486_),
    .Y(_03487_));
 sg13g2_buf_1 _09141_ (.A(_03487_),
    .X(_03488_));
 sg13g2_o21ai_1 _09142_ (.B1(net85),
    .Y(_03489_),
    .A1(_03360_),
    .A2(net88));
 sg13g2_mux2_1 _09143_ (.A0(_01114_),
    .A1(_03489_),
    .S(net38),
    .X(_00470_));
 sg13g2_o21ai_1 _09144_ (.B1(net85),
    .Y(_03490_),
    .A1(_03468_),
    .A2(net88));
 sg13g2_mux2_1 _09145_ (.A0(_01097_),
    .A1(_03490_),
    .S(net38),
    .X(_00471_));
 sg13g2_mux4_1 _09146_ (.S0(net166),
    .A0(_00117_),
    .A1(_00119_),
    .A2(_00118_),
    .A3(_00116_),
    .S1(net120),
    .X(_03491_));
 sg13g2_o21ai_1 _09147_ (.B1(net85),
    .Y(_03492_),
    .A1(net88),
    .A2(_03491_));
 sg13g2_mux2_1 _09148_ (.A0(_00917_),
    .A1(_03492_),
    .S(net38),
    .X(_00472_));
 sg13g2_mux4_1 _09149_ (.S0(net166),
    .A0(_00133_),
    .A1(_00135_),
    .A2(_00134_),
    .A3(_00132_),
    .S1(net120),
    .X(_03493_));
 sg13g2_o21ai_1 _09150_ (.B1(_03488_),
    .Y(_03494_),
    .A1(_03485_),
    .A2(_03493_));
 sg13g2_mux2_1 _09151_ (.A0(\i_tinyqv.cpu.imm[23] ),
    .A1(_03494_),
    .S(net38),
    .X(_00473_));
 sg13g2_mux4_1 _09152_ (.S0(net166),
    .A0(_00137_),
    .A1(_00139_),
    .A2(_00138_),
    .A3(_00136_),
    .S1(_03400_),
    .X(_03495_));
 sg13g2_o21ai_1 _09153_ (.B1(net85),
    .Y(_03496_),
    .A1(net88),
    .A2(_03495_));
 sg13g2_mux2_1 _09154_ (.A0(\i_tinyqv.cpu.imm[24] ),
    .A1(_03496_),
    .S(net38),
    .X(_00474_));
 sg13g2_mux4_1 _09155_ (.S0(_03447_),
    .A0(_00141_),
    .A1(_00143_),
    .A2(_00142_),
    .A3(_00140_),
    .S1(_03400_),
    .X(_03497_));
 sg13g2_nor2_1 _09156_ (.A(net100),
    .B(_03497_),
    .Y(_03498_));
 sg13g2_inv_1 _09157_ (.Y(_03499_),
    .A(_03487_));
 sg13g2_a21oi_1 _09158_ (.A1(_03419_),
    .A2(_03498_),
    .Y(_03500_),
    .B1(_03499_));
 sg13g2_nor2_1 _09159_ (.A(\i_tinyqv.cpu.imm[25] ),
    .B(net37),
    .Y(_03501_));
 sg13g2_a21oi_1 _09160_ (.A1(_03459_),
    .A2(_03500_),
    .Y(_00475_),
    .B1(_03501_));
 sg13g2_o21ai_1 _09161_ (.B1(net85),
    .Y(_03502_),
    .A1(_03145_),
    .A2(net88));
 sg13g2_mux2_1 _09162_ (.A0(\i_tinyqv.cpu.imm[26] ),
    .A1(_03502_),
    .S(net38),
    .X(_00476_));
 sg13g2_inv_1 _09163_ (.Y(_03503_),
    .A(_03195_));
 sg13g2_o21ai_1 _09164_ (.B1(_03488_),
    .Y(_03504_),
    .A1(_03503_),
    .A2(_03485_));
 sg13g2_mux2_1 _09165_ (.A0(\i_tinyqv.cpu.imm[27] ),
    .A1(_03504_),
    .S(net38),
    .X(_00477_));
 sg13g2_mux4_1 _09166_ (.S0(net166),
    .A0(_00149_),
    .A1(_00151_),
    .A2(_00150_),
    .A3(_00148_),
    .S1(net120),
    .X(_03505_));
 sg13g2_o21ai_1 _09167_ (.B1(net85),
    .Y(_03506_),
    .A1(net88),
    .A2(_03505_));
 sg13g2_mux2_1 _09168_ (.A0(\i_tinyqv.cpu.imm[28] ),
    .A1(_03506_),
    .S(net38),
    .X(_00478_));
 sg13g2_mux4_1 _09169_ (.S0(net166),
    .A0(_00121_),
    .A1(_00123_),
    .A2(_00122_),
    .A3(_00120_),
    .S1(net120),
    .X(_03507_));
 sg13g2_o21ai_1 _09170_ (.B1(net85),
    .Y(_03508_),
    .A1(net88),
    .A2(_03507_));
 sg13g2_mux2_1 _09171_ (.A0(\i_tinyqv.cpu.imm[29] ),
    .A1(_03508_),
    .S(_03404_),
    .X(_00479_));
 sg13g2_buf_1 _09172_ (.A(net108),
    .X(_03509_));
 sg13g2_nand2_1 _09173_ (.Y(_03510_),
    .A(net94),
    .B(_03180_));
 sg13g2_nand2_1 _09174_ (.Y(_03511_),
    .A(_03420_),
    .B(_03359_));
 sg13g2_a21oi_1 _09175_ (.A1(_03510_),
    .A2(_03511_),
    .Y(_03512_),
    .B1(_01505_));
 sg13g2_buf_1 _09176_ (.A(_01497_),
    .X(_03513_));
 sg13g2_nor2_1 _09177_ (.A(net103),
    .B(net102),
    .Y(_03514_));
 sg13g2_nand3_1 _09178_ (.B(net122),
    .C(_03514_),
    .A(net113),
    .Y(_03515_));
 sg13g2_a21oi_1 _09179_ (.A1(net106),
    .A2(net110),
    .Y(_03516_),
    .B1(_03515_));
 sg13g2_nor2b_1 _09180_ (.A(net161),
    .B_N(_03365_),
    .Y(_03517_));
 sg13g2_nor2_1 _09181_ (.A(net106),
    .B(net121),
    .Y(_03518_));
 sg13g2_nor2_1 _09182_ (.A(net108),
    .B(net105),
    .Y(_03519_));
 sg13g2_a21oi_1 _09183_ (.A1(net96),
    .A2(_03518_),
    .Y(_03520_),
    .B1(_03519_));
 sg13g2_nor2_1 _09184_ (.A(net113),
    .B(_03520_),
    .Y(_03521_));
 sg13g2_a21oi_1 _09185_ (.A1(net111),
    .A2(net104),
    .Y(_03522_),
    .B1(_03350_));
 sg13g2_nor4_1 _09186_ (.A(_03514_),
    .B(_03517_),
    .C(_03521_),
    .D(_03522_),
    .Y(_03523_));
 sg13g2_nor3_1 _09187_ (.A(net90),
    .B(_03359_),
    .C(_03491_),
    .Y(_03524_));
 sg13g2_nor4_1 _09188_ (.A(_03512_),
    .B(_03516_),
    .C(_03523_),
    .D(_03524_),
    .Y(_03525_));
 sg13g2_nor2_1 _09189_ (.A(_00919_),
    .B(net37),
    .Y(_03526_));
 sg13g2_a21oi_1 _09190_ (.A1(net36),
    .A2(_03525_),
    .Y(_00480_),
    .B1(_03526_));
 sg13g2_o21ai_1 _09191_ (.B1(net85),
    .Y(_03527_),
    .A1(_03213_),
    .A2(net88));
 sg13g2_mux2_1 _09192_ (.A0(\i_tinyqv.cpu.imm[30] ),
    .A1(_03527_),
    .S(net40),
    .X(_00481_));
 sg13g2_inv_1 _09193_ (.Y(_03528_),
    .A(\i_tinyqv.cpu.imm[31] ));
 sg13g2_buf_1 _09194_ (.A(net100),
    .X(_03529_));
 sg13g2_nor2_1 _09195_ (.A(_03529_),
    .B(_03416_),
    .Y(_03530_));
 sg13g2_o21ai_1 _09196_ (.B1(net56),
    .Y(_03531_),
    .A1(_03454_),
    .A2(_03530_));
 sg13g2_o21ai_1 _09197_ (.B1(_03531_),
    .Y(_00482_),
    .A1(_03528_),
    .A2(_03187_));
 sg13g2_nand2_1 _09198_ (.Y(_03532_),
    .A(_01531_),
    .B(_01529_));
 sg13g2_buf_1 _09199_ (.A(_03532_),
    .X(_03533_));
 sg13g2_nand2_1 _09200_ (.Y(_03534_),
    .A(_03156_),
    .B(_01497_));
 sg13g2_a21oi_1 _09201_ (.A1(_03533_),
    .A2(_03534_),
    .Y(_03535_),
    .B1(_03479_));
 sg13g2_o21ai_1 _09202_ (.B1(_03509_),
    .Y(_03536_),
    .A1(_03180_),
    .A2(_03535_));
 sg13g2_and2_1 _09203_ (.A(_03511_),
    .B(_03536_),
    .X(_03537_));
 sg13g2_nor2_1 _09204_ (.A(net147),
    .B(_03537_),
    .Y(_03538_));
 sg13g2_nor3_1 _09205_ (.A(net90),
    .B(_03359_),
    .C(_03493_),
    .Y(_03539_));
 sg13g2_nor2_1 _09206_ (.A(net110),
    .B(_03179_),
    .Y(_03540_));
 sg13g2_o21ai_1 _09207_ (.B1(net104),
    .Y(_03541_),
    .A1(net108),
    .A2(net155));
 sg13g2_nand3_1 _09208_ (.B(net113),
    .C(_03541_),
    .A(_03153_),
    .Y(_03542_));
 sg13g2_o21ai_1 _09209_ (.B1(_03542_),
    .Y(_03543_),
    .A1(net94),
    .A2(net97));
 sg13g2_a22oi_1 _09210_ (.Y(_03544_),
    .B1(_03543_),
    .B2(net96),
    .A2(_03540_),
    .A1(_03393_));
 sg13g2_a21oi_1 _09211_ (.A1(net155),
    .A2(_03365_),
    .Y(_03545_),
    .B1(_03544_));
 sg13g2_nor3_1 _09212_ (.A(_03538_),
    .B(_03539_),
    .C(_03545_),
    .Y(_03546_));
 sg13g2_nor2_1 _09213_ (.A(net329),
    .B(net37),
    .Y(_03547_));
 sg13g2_a21oi_1 _09214_ (.A1(net36),
    .A2(_03546_),
    .Y(_00483_),
    .B1(_03547_));
 sg13g2_a21oi_1 _09215_ (.A1(net94),
    .A2(_03540_),
    .Y(_03548_),
    .B1(_03396_));
 sg13g2_a22oi_1 _09216_ (.Y(_03549_),
    .B1(_03471_),
    .B2(_03548_),
    .A2(_03365_),
    .A1(_01468_));
 sg13g2_nor3_1 _09217_ (.A(net90),
    .B(_03359_),
    .C(_03495_),
    .Y(_03550_));
 sg13g2_nor2_1 _09218_ (.A(net121),
    .B(_03533_),
    .Y(_03551_));
 sg13g2_a21oi_1 _09219_ (.A1(_01461_),
    .A2(net102),
    .Y(_03552_),
    .B1(_03551_));
 sg13g2_nor2_1 _09220_ (.A(net108),
    .B(_03552_),
    .Y(_03553_));
 sg13g2_nor3_1 _09221_ (.A(net113),
    .B(net102),
    .C(_03208_),
    .Y(_03554_));
 sg13g2_o21ai_1 _09222_ (.B1(net96),
    .Y(_03555_),
    .A1(_03553_),
    .A2(_03554_));
 sg13g2_a21oi_1 _09223_ (.A1(_03537_),
    .A2(_03555_),
    .Y(_03556_),
    .B1(_03163_));
 sg13g2_nor3_1 _09224_ (.A(_03549_),
    .B(_03550_),
    .C(_03556_),
    .Y(_03557_));
 sg13g2_nor2_1 _09225_ (.A(_01112_),
    .B(net55),
    .Y(_03558_));
 sg13g2_a21oi_1 _09226_ (.A1(net36),
    .A2(_03557_),
    .Y(_00484_),
    .B1(_03558_));
 sg13g2_o21ai_1 _09227_ (.B1(net173),
    .Y(_03559_),
    .A1(_03396_),
    .A2(_03472_));
 sg13g2_inv_1 _09228_ (.Y(_03560_),
    .A(net147));
 sg13g2_xnor2_1 _09229_ (.Y(_03561_),
    .A(_03189_),
    .B(net104));
 sg13g2_o21ai_1 _09230_ (.B1(net107),
    .Y(_03562_),
    .A1(net106),
    .A2(net105));
 sg13g2_nand3_1 _09231_ (.B(net100),
    .C(_03562_),
    .A(net112),
    .Y(_03563_));
 sg13g2_a21oi_1 _09232_ (.A1(net110),
    .A2(_03561_),
    .Y(_03564_),
    .B1(_03563_));
 sg13g2_a221oi_1 _09233_ (.B2(_03354_),
    .C1(_03564_),
    .B1(_03498_),
    .A1(_03560_),
    .Y(_03565_),
    .A2(_03389_));
 sg13g2_and2_1 _09234_ (.A(_03559_),
    .B(_03565_),
    .X(_03566_));
 sg13g2_nor2_1 _09235_ (.A(_01100_),
    .B(net55),
    .Y(_03567_));
 sg13g2_a21oi_1 _09236_ (.A1(net36),
    .A2(_03566_),
    .Y(_00485_),
    .B1(_03567_));
 sg13g2_nand2_1 _09237_ (.Y(_03568_),
    .A(_03510_),
    .B(_03555_));
 sg13g2_nand3_1 _09238_ (.B(_03167_),
    .C(_03391_),
    .A(net108),
    .Y(_03569_));
 sg13g2_nand2_1 _09239_ (.Y(_03570_),
    .A(_03410_),
    .B(_03569_));
 sg13g2_a22oi_1 _09240_ (.Y(_03571_),
    .B1(_03570_),
    .B2(net107),
    .A2(_03535_),
    .A1(net94));
 sg13g2_nand3_1 _09241_ (.B(_01498_),
    .C(_03518_),
    .A(net173),
    .Y(_03572_));
 sg13g2_o21ai_1 _09242_ (.B1(_03572_),
    .Y(_03573_),
    .A1(_03145_),
    .A2(net90));
 sg13g2_nand2b_1 _09243_ (.Y(_03574_),
    .B(_03368_),
    .A_N(_03212_));
 sg13g2_nor2b_1 _09244_ (.A(_03573_),
    .B_N(_03574_),
    .Y(_03575_));
 sg13g2_o21ai_1 _09245_ (.B1(_03575_),
    .Y(_03576_),
    .A1(net155),
    .A2(_03571_));
 sg13g2_a21oi_1 _09246_ (.A1(_01525_),
    .A2(_03568_),
    .Y(_03577_),
    .B1(_03576_));
 sg13g2_nor2_1 _09247_ (.A(_02650_),
    .B(net55),
    .Y(_03578_));
 sg13g2_a21oi_1 _09248_ (.A1(net36),
    .A2(_03577_),
    .Y(_00486_),
    .B1(_03578_));
 sg13g2_nor2_1 _09249_ (.A(_03189_),
    .B(net111),
    .Y(_03579_));
 sg13g2_nand2_1 _09250_ (.Y(_03580_),
    .A(net135),
    .B(_03350_));
 sg13g2_nor2_1 _09251_ (.A(_03174_),
    .B(_03580_),
    .Y(_03581_));
 sg13g2_a22oi_1 _09252_ (.Y(_03582_),
    .B1(_03581_),
    .B2(net111),
    .A2(_03580_),
    .A1(_03579_));
 sg13g2_nor3_1 _09253_ (.A(net102),
    .B(_01519_),
    .C(_03582_),
    .Y(_03583_));
 sg13g2_a221oi_1 _09254_ (.B2(net122),
    .C1(_03583_),
    .B1(_03472_),
    .A1(_03195_),
    .Y(_03584_),
    .A2(_03420_));
 sg13g2_and2_1 _09255_ (.A(_03574_),
    .B(_03584_),
    .X(_03585_));
 sg13g2_o21ai_1 _09256_ (.B1(_03585_),
    .Y(_03586_),
    .A1(_03132_),
    .A2(_03548_));
 sg13g2_mux2_1 _09257_ (.A0(_00960_),
    .A1(_03586_),
    .S(net40),
    .X(_00487_));
 sg13g2_nor2_1 _09258_ (.A(net90),
    .B(_03505_),
    .Y(_03587_));
 sg13g2_a21oi_1 _09259_ (.A1(_01477_),
    .A2(_03396_),
    .Y(_03588_),
    .B1(_03587_));
 sg13g2_o21ai_1 _09260_ (.B1(_03588_),
    .Y(_03589_),
    .A1(_01505_),
    .A2(_03555_));
 sg13g2_o21ai_1 _09261_ (.B1(_03127_),
    .Y(_03590_),
    .A1(_03384_),
    .A2(_03589_));
 sg13g2_o21ai_1 _09262_ (.B1(_03590_),
    .Y(_00488_),
    .A1(_01546_),
    .A2(_03187_));
 sg13g2_or2_1 _09263_ (.X(_03591_),
    .B(_03507_),
    .A(net90));
 sg13g2_nand3_1 _09264_ (.B(_03560_),
    .C(_03553_),
    .A(_03371_),
    .Y(_03592_));
 sg13g2_nand3_1 _09265_ (.B(_03591_),
    .C(_03592_),
    .A(_03398_),
    .Y(_03593_));
 sg13g2_mux2_1 _09266_ (.A0(_01101_),
    .A1(_03593_),
    .S(net40),
    .X(_00489_));
 sg13g2_nand4_1 _09267_ (.B(_01564_),
    .C(_01567_),
    .A(_01527_),
    .Y(_03594_),
    .D(_01594_));
 sg13g2_buf_1 _09268_ (.A(_03594_),
    .X(_03595_));
 sg13g2_nand4_1 _09269_ (.B(_01598_),
    .C(_01609_),
    .A(_01541_),
    .Y(_03596_),
    .D(_03595_));
 sg13g2_nor2_1 _09270_ (.A(_01586_),
    .B(_03596_),
    .Y(_03597_));
 sg13g2_nand2b_1 _09271_ (.Y(_03598_),
    .B(_03597_),
    .A_N(net313));
 sg13g2_buf_2 _09272_ (.A(_03598_),
    .X(_03599_));
 sg13g2_buf_1 _09273_ (.A(_03599_),
    .X(_03600_));
 sg13g2_o21ai_1 _09274_ (.B1(_03599_),
    .Y(_03601_),
    .A1(\i_tinyqv.cpu.instr_data[0][0] ),
    .A2(net271));
 sg13g2_o21ai_1 _09275_ (.B1(_03601_),
    .Y(_00490_),
    .A1(_02534_),
    .A2(net54));
 sg13g2_buf_2 _09276_ (.A(_00213_),
    .X(_03602_));
 sg13g2_buf_1 _09277_ (.A(_03599_),
    .X(_03603_));
 sg13g2_nand2_1 _09278_ (.Y(_03604_),
    .A(\i_tinyqv.cpu.instr_data[0][10] ),
    .B(net53));
 sg13g2_o21ai_1 _09279_ (.B1(_03604_),
    .Y(_00491_),
    .A1(_03602_),
    .A2(net54));
 sg13g2_buf_2 _09280_ (.A(_00214_),
    .X(_03605_));
 sg13g2_nand2_1 _09281_ (.Y(_03606_),
    .A(\i_tinyqv.cpu.instr_data[0][11] ),
    .B(net53));
 sg13g2_o21ai_1 _09282_ (.B1(_03606_),
    .Y(_00492_),
    .A1(_03605_),
    .A2(net54));
 sg13g2_buf_2 _09283_ (.A(_00208_),
    .X(_03607_));
 sg13g2_nand2_1 _09284_ (.Y(_03608_),
    .A(\i_tinyqv.cpu.instr_data[0][12] ),
    .B(net53));
 sg13g2_o21ai_1 _09285_ (.B1(_03608_),
    .Y(_00493_),
    .A1(_03607_),
    .A2(net54));
 sg13g2_buf_2 _09286_ (.A(_00209_),
    .X(_03609_));
 sg13g2_nand2_1 _09287_ (.Y(_03610_),
    .A(\i_tinyqv.cpu.instr_data[0][13] ),
    .B(_03603_));
 sg13g2_o21ai_1 _09288_ (.B1(_03610_),
    .Y(_00494_),
    .A1(_03609_),
    .A2(net54));
 sg13g2_buf_2 _09289_ (.A(_00215_),
    .X(_03611_));
 sg13g2_nand2_1 _09290_ (.Y(_03612_),
    .A(\i_tinyqv.cpu.instr_data[0][14] ),
    .B(_03599_));
 sg13g2_o21ai_1 _09291_ (.B1(_03612_),
    .Y(_00495_),
    .A1(_03611_),
    .A2(net54));
 sg13g2_buf_2 _09292_ (.A(_00210_),
    .X(_03613_));
 sg13g2_nand2_1 _09293_ (.Y(_03614_),
    .A(\i_tinyqv.cpu.instr_data[0][15] ),
    .B(_03599_));
 sg13g2_o21ai_1 _09294_ (.B1(_03614_),
    .Y(_00496_),
    .A1(_03613_),
    .A2(_03600_));
 sg13g2_inv_1 _09295_ (.Y(_03615_),
    .A(\i_tinyqv.cpu.instr_data_in[1] ));
 sg13g2_o21ai_1 _09296_ (.B1(_03599_),
    .Y(_03616_),
    .A1(net271),
    .A2(\i_tinyqv.cpu.instr_data[0][1] ));
 sg13g2_o21ai_1 _09297_ (.B1(_03616_),
    .Y(_00497_),
    .A1(_03615_),
    .A2(net54));
 sg13g2_mux2_1 _09298_ (.A0(_02905_),
    .A1(\i_tinyqv.cpu.instr_data[0][2] ),
    .S(net53),
    .X(_00498_));
 sg13g2_mux2_1 _09299_ (.A0(_03012_),
    .A1(\i_tinyqv.cpu.instr_data[0][3] ),
    .S(net53),
    .X(_00499_));
 sg13g2_mux2_1 _09300_ (.A0(_02577_),
    .A1(\i_tinyqv.cpu.instr_data[0][4] ),
    .S(net53),
    .X(_00500_));
 sg13g2_mux2_1 _09301_ (.A0(_02773_),
    .A1(\i_tinyqv.cpu.instr_data[0][5] ),
    .S(net53),
    .X(_00501_));
 sg13g2_mux2_1 _09302_ (.A0(_02899_),
    .A1(\i_tinyqv.cpu.instr_data[0][6] ),
    .S(net53),
    .X(_00502_));
 sg13g2_mux2_1 _09303_ (.A0(_02962_),
    .A1(\i_tinyqv.cpu.instr_data[0][7] ),
    .S(_03603_),
    .X(_00503_));
 sg13g2_buf_2 _09304_ (.A(_00211_),
    .X(_03617_));
 sg13g2_nand2_1 _09305_ (.Y(_03618_),
    .A(\i_tinyqv.cpu.instr_data[0][8] ),
    .B(_03599_));
 sg13g2_o21ai_1 _09306_ (.B1(_03618_),
    .Y(_00504_),
    .A1(_03617_),
    .A2(net54));
 sg13g2_buf_2 _09307_ (.A(_00212_),
    .X(_03619_));
 sg13g2_nand2_1 _09308_ (.Y(_03620_),
    .A(\i_tinyqv.cpu.instr_data[0][9] ),
    .B(_03599_));
 sg13g2_o21ai_1 _09309_ (.B1(_03620_),
    .Y(_00505_),
    .A1(_03619_),
    .A2(_03600_));
 sg13g2_nor2b_1 _09310_ (.A(net313),
    .B_N(_01586_),
    .Y(_03621_));
 sg13g2_nand2b_1 _09311_ (.Y(_03622_),
    .B(_03621_),
    .A_N(_03596_));
 sg13g2_buf_2 _09312_ (.A(_03622_),
    .X(_03623_));
 sg13g2_buf_1 _09313_ (.A(_03623_),
    .X(_03624_));
 sg13g2_o21ai_1 _09314_ (.B1(_03623_),
    .Y(_03625_),
    .A1(\i_tinyqv.cpu.instr_data[1][0] ),
    .A2(net271));
 sg13g2_o21ai_1 _09315_ (.B1(_03625_),
    .Y(_00506_),
    .A1(_02534_),
    .A2(net66));
 sg13g2_buf_1 _09316_ (.A(_03623_),
    .X(_03626_));
 sg13g2_nand2_1 _09317_ (.Y(_03627_),
    .A(\i_tinyqv.cpu.instr_data[1][10] ),
    .B(net65));
 sg13g2_o21ai_1 _09318_ (.B1(_03627_),
    .Y(_00507_),
    .A1(_03602_),
    .A2(net66));
 sg13g2_nand2_1 _09319_ (.Y(_03628_),
    .A(\i_tinyqv.cpu.instr_data[1][11] ),
    .B(net65));
 sg13g2_o21ai_1 _09320_ (.B1(_03628_),
    .Y(_00508_),
    .A1(_03605_),
    .A2(net66));
 sg13g2_nand2_1 _09321_ (.Y(_03629_),
    .A(\i_tinyqv.cpu.instr_data[1][12] ),
    .B(net65));
 sg13g2_o21ai_1 _09322_ (.B1(_03629_),
    .Y(_00509_),
    .A1(_03607_),
    .A2(net66));
 sg13g2_nand2_1 _09323_ (.Y(_03630_),
    .A(\i_tinyqv.cpu.instr_data[1][13] ),
    .B(_03626_));
 sg13g2_o21ai_1 _09324_ (.B1(_03630_),
    .Y(_00510_),
    .A1(_03609_),
    .A2(net66));
 sg13g2_nand2_1 _09325_ (.Y(_03631_),
    .A(\i_tinyqv.cpu.instr_data[1][14] ),
    .B(_03623_));
 sg13g2_o21ai_1 _09326_ (.B1(_03631_),
    .Y(_00511_),
    .A1(_03611_),
    .A2(_03624_));
 sg13g2_nand2_1 _09327_ (.Y(_03632_),
    .A(\i_tinyqv.cpu.instr_data[1][15] ),
    .B(_03623_));
 sg13g2_o21ai_1 _09328_ (.B1(_03632_),
    .Y(_00512_),
    .A1(_03613_),
    .A2(net66));
 sg13g2_o21ai_1 _09329_ (.B1(_03623_),
    .Y(_03633_),
    .A1(net271),
    .A2(\i_tinyqv.cpu.instr_data[1][1] ));
 sg13g2_o21ai_1 _09330_ (.B1(_03633_),
    .Y(_00513_),
    .A1(_03615_),
    .A2(_03624_));
 sg13g2_mux2_1 _09331_ (.A0(_02905_),
    .A1(\i_tinyqv.cpu.instr_data[1][2] ),
    .S(net65),
    .X(_00514_));
 sg13g2_mux2_1 _09332_ (.A0(_03012_),
    .A1(\i_tinyqv.cpu.instr_data[1][3] ),
    .S(net65),
    .X(_00515_));
 sg13g2_mux2_1 _09333_ (.A0(_02577_),
    .A1(\i_tinyqv.cpu.instr_data[1][4] ),
    .S(net65),
    .X(_00516_));
 sg13g2_mux2_1 _09334_ (.A0(_02773_),
    .A1(\i_tinyqv.cpu.instr_data[1][5] ),
    .S(net65),
    .X(_00517_));
 sg13g2_mux2_1 _09335_ (.A0(_02899_),
    .A1(\i_tinyqv.cpu.instr_data[1][6] ),
    .S(net65),
    .X(_00518_));
 sg13g2_mux2_1 _09336_ (.A0(_02962_),
    .A1(\i_tinyqv.cpu.instr_data[1][7] ),
    .S(_03626_),
    .X(_00519_));
 sg13g2_nand2_1 _09337_ (.Y(_03634_),
    .A(\i_tinyqv.cpu.instr_data[1][8] ),
    .B(_03623_));
 sg13g2_o21ai_1 _09338_ (.B1(_03634_),
    .Y(_00520_),
    .A1(_03617_),
    .A2(net66));
 sg13g2_nand2_1 _09339_ (.Y(_03635_),
    .A(\i_tinyqv.cpu.instr_data[1][9] ),
    .B(_03623_));
 sg13g2_o21ai_1 _09340_ (.B1(_03635_),
    .Y(_00521_),
    .A1(_03619_),
    .A2(net66));
 sg13g2_nand2_1 _09341_ (.Y(_03636_),
    .A(net313),
    .B(_03597_));
 sg13g2_buf_2 _09342_ (.A(_03636_),
    .X(_03637_));
 sg13g2_buf_1 _09343_ (.A(_03637_),
    .X(_03638_));
 sg13g2_o21ai_1 _09344_ (.B1(_03637_),
    .Y(_03639_),
    .A1(\i_tinyqv.cpu.instr_data[2][0] ),
    .A2(net271));
 sg13g2_o21ai_1 _09345_ (.B1(_03639_),
    .Y(_00522_),
    .A1(_02534_),
    .A2(net52));
 sg13g2_buf_1 _09346_ (.A(_03637_),
    .X(_03640_));
 sg13g2_nand2_1 _09347_ (.Y(_03641_),
    .A(\i_tinyqv.cpu.instr_data[2][10] ),
    .B(net51));
 sg13g2_o21ai_1 _09348_ (.B1(_03641_),
    .Y(_00523_),
    .A1(_03602_),
    .A2(net52));
 sg13g2_nand2_1 _09349_ (.Y(_03642_),
    .A(\i_tinyqv.cpu.instr_data[2][11] ),
    .B(net51));
 sg13g2_o21ai_1 _09350_ (.B1(_03642_),
    .Y(_00524_),
    .A1(_03605_),
    .A2(net52));
 sg13g2_nand2_1 _09351_ (.Y(_03643_),
    .A(\i_tinyqv.cpu.instr_data[2][12] ),
    .B(net51));
 sg13g2_o21ai_1 _09352_ (.B1(_03643_),
    .Y(_00525_),
    .A1(_03607_),
    .A2(net52));
 sg13g2_nand2_1 _09353_ (.Y(_03644_),
    .A(\i_tinyqv.cpu.instr_data[2][13] ),
    .B(_03640_));
 sg13g2_o21ai_1 _09354_ (.B1(_03644_),
    .Y(_00526_),
    .A1(_03609_),
    .A2(net52));
 sg13g2_nand2_1 _09355_ (.Y(_03645_),
    .A(\i_tinyqv.cpu.instr_data[2][14] ),
    .B(_03637_));
 sg13g2_o21ai_1 _09356_ (.B1(_03645_),
    .Y(_00527_),
    .A1(_03611_),
    .A2(net52));
 sg13g2_nand2_1 _09357_ (.Y(_03646_),
    .A(\i_tinyqv.cpu.instr_data[2][15] ),
    .B(_03637_));
 sg13g2_o21ai_1 _09358_ (.B1(_03646_),
    .Y(_00528_),
    .A1(_03613_),
    .A2(net52));
 sg13g2_o21ai_1 _09359_ (.B1(_03637_),
    .Y(_03647_),
    .A1(net271),
    .A2(\i_tinyqv.cpu.instr_data[2][1] ));
 sg13g2_o21ai_1 _09360_ (.B1(_03647_),
    .Y(_00529_),
    .A1(_03615_),
    .A2(_03638_));
 sg13g2_mux2_1 _09361_ (.A0(_02905_),
    .A1(\i_tinyqv.cpu.instr_data[2][2] ),
    .S(net51),
    .X(_00530_));
 sg13g2_mux2_1 _09362_ (.A0(_03012_),
    .A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .S(net51),
    .X(_00531_));
 sg13g2_mux2_1 _09363_ (.A0(_02577_),
    .A1(\i_tinyqv.cpu.instr_data[2][4] ),
    .S(net51),
    .X(_00532_));
 sg13g2_mux2_1 _09364_ (.A0(_02773_),
    .A1(\i_tinyqv.cpu.instr_data[2][5] ),
    .S(net51),
    .X(_00533_));
 sg13g2_mux2_1 _09365_ (.A0(_02899_),
    .A1(\i_tinyqv.cpu.instr_data[2][6] ),
    .S(net51),
    .X(_00534_));
 sg13g2_mux2_1 _09366_ (.A0(_02962_),
    .A1(\i_tinyqv.cpu.instr_data[2][7] ),
    .S(_03640_),
    .X(_00535_));
 sg13g2_nand2_1 _09367_ (.Y(_03648_),
    .A(\i_tinyqv.cpu.instr_data[2][8] ),
    .B(_03637_));
 sg13g2_o21ai_1 _09368_ (.B1(_03648_),
    .Y(_00536_),
    .A1(_03617_),
    .A2(net52));
 sg13g2_nand2_1 _09369_ (.Y(_03649_),
    .A(\i_tinyqv.cpu.instr_data[2][9] ),
    .B(_03637_));
 sg13g2_o21ai_1 _09370_ (.B1(_03649_),
    .Y(_00537_),
    .A1(_03619_),
    .A2(_03638_));
 sg13g2_buf_1 _09371_ (.A(_01598_),
    .X(_03650_));
 sg13g2_and2_1 _09372_ (.A(net84),
    .B(_03595_),
    .X(_03651_));
 sg13g2_buf_1 _09373_ (.A(_03651_),
    .X(_03652_));
 sg13g2_nand4_1 _09374_ (.B(_01575_),
    .C(_01609_),
    .A(_01586_),
    .Y(_03653_),
    .D(net75));
 sg13g2_buf_1 _09375_ (.A(_03653_),
    .X(_03654_));
 sg13g2_nor2_1 _09376_ (.A(\i_tinyqv.cpu.instr_data_in[0] ),
    .B(_03654_),
    .Y(_03655_));
 sg13g2_nor2b_1 _09377_ (.A(\i_tinyqv.cpu.instr_data[3][0] ),
    .B_N(_03654_),
    .Y(_03656_));
 sg13g2_buf_1 _09378_ (.A(_01541_),
    .X(_03657_));
 sg13g2_o21ai_1 _09379_ (.B1(net251),
    .Y(_00538_),
    .A1(_03655_),
    .A2(_03656_));
 sg13g2_inv_1 _09380_ (.Y(_03658_),
    .A(_03602_));
 sg13g2_nand2_1 _09381_ (.Y(_03659_),
    .A(_01586_),
    .B(net313));
 sg13g2_nor2_1 _09382_ (.A(_03596_),
    .B(_03659_),
    .Y(_03660_));
 sg13g2_buf_2 _09383_ (.A(_03660_),
    .X(_03661_));
 sg13g2_buf_2 _09384_ (.A(_03661_),
    .X(_03662_));
 sg13g2_mux2_1 _09385_ (.A0(\i_tinyqv.cpu.instr_data[3][10] ),
    .A1(_03658_),
    .S(net64),
    .X(_00539_));
 sg13g2_inv_1 _09386_ (.Y(_03663_),
    .A(_03605_));
 sg13g2_mux2_1 _09387_ (.A0(\i_tinyqv.cpu.instr_data[3][11] ),
    .A1(_03663_),
    .S(_03662_),
    .X(_00540_));
 sg13g2_inv_1 _09388_ (.Y(_03664_),
    .A(_03607_));
 sg13g2_mux2_1 _09389_ (.A0(\i_tinyqv.cpu.instr_data[3][12] ),
    .A1(_03664_),
    .S(net64),
    .X(_00541_));
 sg13g2_inv_1 _09390_ (.Y(_03665_),
    .A(_03609_));
 sg13g2_mux2_1 _09391_ (.A0(\i_tinyqv.cpu.instr_data[3][13] ),
    .A1(_03665_),
    .S(net64),
    .X(_00542_));
 sg13g2_inv_1 _09392_ (.Y(_03666_),
    .A(_03611_));
 sg13g2_mux2_1 _09393_ (.A0(\i_tinyqv.cpu.instr_data[3][14] ),
    .A1(_03666_),
    .S(_03662_),
    .X(_00543_));
 sg13g2_inv_1 _09394_ (.Y(_03667_),
    .A(_03613_));
 sg13g2_mux2_1 _09395_ (.A0(\i_tinyqv.cpu.instr_data[3][15] ),
    .A1(_03667_),
    .S(net64),
    .X(_00544_));
 sg13g2_nor2_1 _09396_ (.A(\i_tinyqv.cpu.instr_data_in[1] ),
    .B(_03654_),
    .Y(_03668_));
 sg13g2_nor2b_1 _09397_ (.A(\i_tinyqv.cpu.instr_data[3][1] ),
    .B_N(_03654_),
    .Y(_03669_));
 sg13g2_o21ai_1 _09398_ (.B1(net251),
    .Y(_00545_),
    .A1(_03668_),
    .A2(_03669_));
 sg13g2_mux2_1 _09399_ (.A0(\i_tinyqv.cpu.instr_data[3][2] ),
    .A1(_02905_),
    .S(net64),
    .X(_00546_));
 sg13g2_mux2_1 _09400_ (.A0(\i_tinyqv.cpu.instr_data[3][3] ),
    .A1(_03012_),
    .S(net64),
    .X(_00547_));
 sg13g2_mux2_1 _09401_ (.A0(\i_tinyqv.cpu.instr_data[3][4] ),
    .A1(_02577_),
    .S(net64),
    .X(_00548_));
 sg13g2_mux2_1 _09402_ (.A0(\i_tinyqv.cpu.instr_data[3][5] ),
    .A1(_02773_),
    .S(net64),
    .X(_00549_));
 sg13g2_mux2_1 _09403_ (.A0(\i_tinyqv.cpu.instr_data[3][6] ),
    .A1(_02899_),
    .S(_03661_),
    .X(_00550_));
 sg13g2_mux2_1 _09404_ (.A0(\i_tinyqv.cpu.instr_data[3][7] ),
    .A1(_02962_),
    .S(_03661_),
    .X(_00551_));
 sg13g2_inv_1 _09405_ (.Y(_03670_),
    .A(_03617_));
 sg13g2_mux2_1 _09406_ (.A0(\i_tinyqv.cpu.instr_data[3][8] ),
    .A1(_03670_),
    .S(_03661_),
    .X(_00552_));
 sg13g2_inv_1 _09407_ (.Y(_03671_),
    .A(_03619_));
 sg13g2_mux2_1 _09408_ (.A0(\i_tinyqv.cpu.instr_data[3][9] ),
    .A1(_03671_),
    .S(_03661_),
    .X(_00553_));
 sg13g2_o21ai_1 _09409_ (.B1(net104),
    .Y(_03672_),
    .A1(net121),
    .A2(net135));
 sg13g2_nand2_1 _09410_ (.Y(_03673_),
    .A(net95),
    .B(_03533_));
 sg13g2_a22oi_1 _09411_ (.Y(_03674_),
    .B1(_03673_),
    .B2(_03509_),
    .A2(_03672_),
    .A1(net103));
 sg13g2_nor3_1 _09412_ (.A(_03136_),
    .B(net122),
    .C(_01483_),
    .Y(_03675_));
 sg13g2_nor3_1 _09413_ (.A(_03158_),
    .B(net91),
    .C(_03675_),
    .Y(_03676_));
 sg13g2_a221oi_1 _09414_ (.B2(_03560_),
    .C1(_03676_),
    .B1(_03674_),
    .A1(_03167_),
    .Y(_03677_),
    .A2(_03405_));
 sg13g2_nor2_1 _09415_ (.A(_01556_),
    .B(_03378_),
    .Y(_03678_));
 sg13g2_a21oi_1 _09416_ (.A1(net36),
    .A2(_03677_),
    .Y(_00594_),
    .B1(_03678_));
 sg13g2_nor2_1 _09417_ (.A(net135),
    .B(net105),
    .Y(_03679_));
 sg13g2_o21ai_1 _09418_ (.B1(_03679_),
    .Y(_03680_),
    .A1(net95),
    .A2(net102));
 sg13g2_o21ai_1 _09419_ (.B1(_03680_),
    .Y(_03681_),
    .A1(_03190_),
    .A2(_03672_));
 sg13g2_mux2_1 _09420_ (.A0(_02509_),
    .A1(_03681_),
    .S(net40),
    .X(_00595_));
 sg13g2_nand2_1 _09421_ (.Y(_03682_),
    .A(_03199_),
    .B(_03137_));
 sg13g2_o21ai_1 _09422_ (.B1(_03357_),
    .Y(_03683_),
    .A1(_03174_),
    .A2(net112));
 sg13g2_o21ai_1 _09423_ (.B1(_03683_),
    .Y(_03684_),
    .A1(_03682_),
    .A2(_03158_));
 sg13g2_a21oi_1 _09424_ (.A1(_03177_),
    .A2(_03684_),
    .Y(_03685_),
    .B1(net100));
 sg13g2_o21ai_1 _09425_ (.B1(_03163_),
    .Y(_03686_),
    .A1(_01468_),
    .A2(_01503_));
 sg13g2_inv_1 _09426_ (.Y(_03687_),
    .A(_03686_));
 sg13g2_a22oi_1 _09427_ (.Y(_03688_),
    .B1(_03687_),
    .B2(_03674_),
    .A2(_03685_),
    .A1(net94));
 sg13g2_nor2_1 _09428_ (.A(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .B(_03378_),
    .Y(_03689_));
 sg13g2_a21oi_1 _09429_ (.A1(net39),
    .A2(_03688_),
    .Y(_00596_),
    .B1(_03689_));
 sg13g2_inv_1 _09430_ (.Y(_03690_),
    .A(_03357_));
 sg13g2_nor4_1 _09431_ (.A(_03150_),
    .B(net91),
    .C(_03690_),
    .D(_03387_),
    .Y(_03691_));
 sg13g2_buf_2 _09432_ (.A(\i_tinyqv.cpu.mem_op_increment_reg ),
    .X(_03692_));
 sg13g2_nor2_1 _09433_ (.A(_03692_),
    .B(net55),
    .Y(_03693_));
 sg13g2_a21oi_1 _09434_ (.A1(net39),
    .A2(_03691_),
    .Y(_00597_),
    .B1(_03693_));
 sg13g2_nor2_1 _09435_ (.A(_01328_),
    .B(_03121_),
    .Y(_03694_));
 sg13g2_buf_2 _09436_ (.A(_03694_),
    .X(_03695_));
 sg13g2_buf_1 _09437_ (.A(_03695_),
    .X(_03696_));
 sg13g2_nand2_1 _09438_ (.Y(_03697_),
    .A(net108),
    .B(_01585_));
 sg13g2_o21ai_1 _09439_ (.B1(_03697_),
    .Y(_03698_),
    .A1(_03682_),
    .A2(_03533_));
 sg13g2_o21ai_1 _09440_ (.B1(_03385_),
    .Y(_03699_),
    .A1(_03393_),
    .A2(_03522_));
 sg13g2_a21oi_1 _09441_ (.A1(net110),
    .A2(_03698_),
    .Y(_03700_),
    .B1(_03699_));
 sg13g2_nand4_1 _09442_ (.B(_01484_),
    .C(_01498_),
    .A(net135),
    .Y(_03701_),
    .D(_03150_));
 sg13g2_nand3_1 _09443_ (.B(_03157_),
    .C(_03701_),
    .A(_03190_),
    .Y(_03702_));
 sg13g2_o21ai_1 _09444_ (.B1(_03702_),
    .Y(_03703_),
    .A1(_03157_),
    .A2(_01532_));
 sg13g2_nand2_1 _09445_ (.Y(_03704_),
    .A(_03208_),
    .B(_03385_));
 sg13g2_a22oi_1 _09446_ (.Y(_03705_),
    .B1(_03704_),
    .B2(_01480_),
    .A2(_03703_),
    .A1(net102));
 sg13g2_o21ai_1 _09447_ (.B1(net103),
    .Y(_03706_),
    .A1(net102),
    .A2(_03703_));
 sg13g2_a22oi_1 _09448_ (.Y(_03707_),
    .B1(_03705_),
    .B2(_03706_),
    .A2(_03700_),
    .A1(net136));
 sg13g2_nand2_1 _09449_ (.Y(_03708_),
    .A(_00217_),
    .B(_03695_));
 sg13g2_o21ai_1 _09450_ (.B1(_03708_),
    .Y(_03709_),
    .A1(net74),
    .A2(_03707_));
 sg13g2_a21oi_1 _09451_ (.A1(_03123_),
    .A2(_03119_),
    .Y(_03710_),
    .B1(_01767_));
 sg13g2_buf_1 _09452_ (.A(_03710_),
    .X(_03711_));
 sg13g2_buf_1 _09453_ (.A(_03711_),
    .X(_03712_));
 sg13g2_mux2_1 _09454_ (.A0(_02712_),
    .A1(_03709_),
    .S(net63),
    .X(_00601_));
 sg13g2_buf_1 _09455_ (.A(_03123_),
    .X(_03713_));
 sg13g2_o21ai_1 _09456_ (.B1(_03711_),
    .Y(_03714_),
    .A1(_02712_),
    .A2(net73));
 sg13g2_o21ai_1 _09457_ (.B1(_03385_),
    .Y(_03715_),
    .A1(_03352_),
    .A2(_03208_));
 sg13g2_a221oi_1 _09458_ (.B2(net171),
    .C1(_03695_),
    .B1(_03715_),
    .A1(_03401_),
    .Y(_03716_),
    .A2(_03700_));
 sg13g2_a21oi_1 _09459_ (.A1(_03028_),
    .A2(net74),
    .Y(_03717_),
    .B1(_03716_));
 sg13g2_a22oi_1 _09460_ (.Y(_03718_),
    .B1(_03717_),
    .B2(net63),
    .A2(_03714_),
    .A1(_02711_));
 sg13g2_inv_1 _09461_ (.Y(_00602_),
    .A(_03718_));
 sg13g2_nor3_1 _09462_ (.A(_02714_),
    .B(_02713_),
    .C(net73),
    .Y(_03719_));
 sg13g2_inv_1 _09463_ (.Y(_03720_),
    .A(_01505_));
 sg13g2_a22oi_1 _09464_ (.Y(_03721_),
    .B1(_03715_),
    .B2(net161),
    .A2(_03700_),
    .A1(_03720_));
 sg13g2_nor2_1 _09465_ (.A(net74),
    .B(_03721_),
    .Y(_03722_));
 sg13g2_o21ai_1 _09466_ (.B1(net63),
    .Y(_03723_),
    .A1(_03719_),
    .A2(_03722_));
 sg13g2_and2_1 _09467_ (.A(_02711_),
    .B(_02712_),
    .X(_03724_));
 sg13g2_buf_1 _09468_ (.A(_03724_),
    .X(_03725_));
 sg13g2_o21ai_1 _09469_ (.B1(_03711_),
    .Y(_03726_),
    .A1(_03725_),
    .A2(net73));
 sg13g2_nand2_1 _09470_ (.Y(_03727_),
    .A(_02714_),
    .B(_03726_));
 sg13g2_nand2_1 _09471_ (.Y(_00603_),
    .A(_03723_),
    .B(_03727_));
 sg13g2_o21ai_1 _09472_ (.B1(net106),
    .Y(_03728_),
    .A1(_03177_),
    .A2(_03682_));
 sg13g2_nand2_1 _09473_ (.Y(_03729_),
    .A(_03370_),
    .B(_03728_));
 sg13g2_o21ai_1 _09474_ (.B1(net96),
    .Y(_03730_),
    .A1(net104),
    .A2(_01532_));
 sg13g2_a22oi_1 _09475_ (.Y(_03731_),
    .B1(_03730_),
    .B2(net95),
    .A2(_03729_),
    .A1(net103));
 sg13g2_a21oi_1 _09476_ (.A1(_03580_),
    .A2(_03697_),
    .Y(_03732_),
    .B1(net95));
 sg13g2_nor2_1 _09477_ (.A(_03514_),
    .B(_03732_),
    .Y(_03733_));
 sg13g2_o21ai_1 _09478_ (.B1(_03733_),
    .Y(_03734_),
    .A1(net147),
    .A2(_03731_));
 sg13g2_nand4_1 _09479_ (.B(_02715_),
    .C(_03725_),
    .A(_02714_),
    .Y(_03735_),
    .D(_03695_));
 sg13g2_o21ai_1 _09480_ (.B1(_03735_),
    .Y(_03736_),
    .A1(net74),
    .A2(_03734_));
 sg13g2_a21o_1 _09481_ (.A2(_03725_),
    .A1(_02714_),
    .B1(_03123_),
    .X(_03737_));
 sg13g2_a21oi_1 _09482_ (.A1(net63),
    .A2(_03737_),
    .Y(_03738_),
    .B1(_02715_));
 sg13g2_a21oi_1 _09483_ (.A1(net63),
    .A2(_03736_),
    .Y(_00604_),
    .B1(_03738_));
 sg13g2_nor2_1 _09484_ (.A(net95),
    .B(net91),
    .Y(_03739_));
 sg13g2_nand4_1 _09485_ (.B(net135),
    .C(_03682_),
    .A(net110),
    .Y(_03740_),
    .D(net109));
 sg13g2_nor3_1 _09486_ (.A(net108),
    .B(net105),
    .C(_03672_),
    .Y(_03741_));
 sg13g2_o21ai_1 _09487_ (.B1(_01461_),
    .Y(_03742_),
    .A1(_03189_),
    .A2(net104));
 sg13g2_nand2_1 _09488_ (.Y(_03743_),
    .A(net121),
    .B(_03742_));
 sg13g2_o21ai_1 _09489_ (.B1(_03743_),
    .Y(_03744_),
    .A1(net107),
    .A2(_03561_));
 sg13g2_a22oi_1 _09490_ (.Y(_03745_),
    .B1(_03744_),
    .B2(net96),
    .A2(_03741_),
    .A1(_03740_));
 sg13g2_buf_1 _09491_ (.A(_03745_),
    .X(_03746_));
 sg13g2_nor2b_1 _09492_ (.A(_03746_),
    .B_N(net136),
    .Y(_03747_));
 sg13g2_nor4_1 _09493_ (.A(net89),
    .B(_03394_),
    .C(_03739_),
    .D(_03747_),
    .Y(_03748_));
 sg13g2_nor2_1 _09494_ (.A(net289),
    .B(net55),
    .Y(_03749_));
 sg13g2_a21oi_1 _09495_ (.A1(net39),
    .A2(_03748_),
    .Y(_00605_),
    .B1(_03749_));
 sg13g2_nor2_1 _09496_ (.A(_01531_),
    .B(_01584_),
    .Y(_03750_));
 sg13g2_nand2_1 _09497_ (.Y(_03751_),
    .A(net110),
    .B(_03750_));
 sg13g2_o21ai_1 _09498_ (.B1(_03751_),
    .Y(_03752_),
    .A1(net107),
    .A2(net96));
 sg13g2_xnor2_1 _09499_ (.Y(_03753_),
    .A(net107),
    .B(net103));
 sg13g2_a22oi_1 _09500_ (.Y(_03754_),
    .B1(_03753_),
    .B2(_03409_),
    .A2(_03752_),
    .A1(net94));
 sg13g2_a221oi_1 _09501_ (.B2(_03750_),
    .C1(net97),
    .B1(_03518_),
    .A1(net103),
    .Y(_03755_),
    .A2(_03448_));
 sg13g2_a21oi_1 _09502_ (.A1(net97),
    .A2(_03754_),
    .Y(_03756_),
    .B1(_03755_));
 sg13g2_nor2_1 _09503_ (.A(_01519_),
    .B(_03746_),
    .Y(_03757_));
 sg13g2_o21ai_1 _09504_ (.B1(net56),
    .Y(_03758_),
    .A1(_03756_),
    .A2(_03757_));
 sg13g2_o21ai_1 _09505_ (.B1(_03758_),
    .Y(_00606_),
    .A1(_00788_),
    .A2(net39));
 sg13g2_nand2_1 _09506_ (.Y(_03759_),
    .A(_03513_),
    .B(_03455_));
 sg13g2_o21ai_1 _09507_ (.B1(_03759_),
    .Y(_03760_),
    .A1(net102),
    .A2(_03387_));
 sg13g2_nor2_1 _09508_ (.A(_01505_),
    .B(_03746_),
    .Y(_03761_));
 sg13g2_a21oi_1 _09509_ (.A1(net103),
    .A2(_03760_),
    .Y(_03762_),
    .B1(_03761_));
 sg13g2_nor2_1 _09510_ (.A(net287),
    .B(net55),
    .Y(_03763_));
 sg13g2_a21oi_1 _09511_ (.A1(net39),
    .A2(_03762_),
    .Y(_00607_),
    .B1(_03763_));
 sg13g2_o21ai_1 _09512_ (.B1(_03743_),
    .Y(_03764_),
    .A1(net106),
    .A2(_03533_));
 sg13g2_a21oi_1 _09513_ (.A1(_03371_),
    .A2(_03764_),
    .Y(_03765_),
    .B1(_03560_));
 sg13g2_nor2_1 _09514_ (.A(_03746_),
    .B(_03765_),
    .Y(_03766_));
 sg13g2_a21oi_1 _09515_ (.A1(net92),
    .A2(_03460_),
    .Y(_03767_),
    .B1(_03766_));
 sg13g2_nor2_1 _09516_ (.A(net286),
    .B(net55),
    .Y(_03768_));
 sg13g2_a21oi_1 _09517_ (.A1(net39),
    .A2(_03767_),
    .Y(_00608_),
    .B1(_03768_));
 sg13g2_o21ai_1 _09518_ (.B1(_03711_),
    .Y(_03769_),
    .A1(_03692_),
    .A2(net73));
 sg13g2_nand2_1 _09519_ (.Y(_03770_),
    .A(_03167_),
    .B(_03579_));
 sg13g2_a221oi_1 _09520_ (.B2(_01479_),
    .C1(net89),
    .B1(_03770_),
    .A1(_03479_),
    .Y(_03771_),
    .A2(_03513_));
 sg13g2_a21oi_1 _09521_ (.A1(net92),
    .A2(_03360_),
    .Y(_03772_),
    .B1(_03771_));
 sg13g2_nand3_1 _09522_ (.B(_03692_),
    .C(net74),
    .A(net281),
    .Y(_03773_));
 sg13g2_o21ai_1 _09523_ (.B1(_03773_),
    .Y(_03774_),
    .A1(net74),
    .A2(_03772_));
 sg13g2_a22oi_1 _09524_ (.Y(_00609_),
    .B1(_03774_),
    .B2(net63),
    .A2(_03769_),
    .A1(_00856_));
 sg13g2_nor2_1 _09525_ (.A(_03209_),
    .B(net89),
    .Y(_03775_));
 sg13g2_a21oi_1 _09526_ (.A1(net171),
    .A2(_03775_),
    .Y(_03776_),
    .B1(net92));
 sg13g2_a21oi_1 _09527_ (.A1(net92),
    .A2(_03468_),
    .Y(_03777_),
    .B1(_03776_));
 sg13g2_nand3_1 _09528_ (.B(_00902_),
    .C(_03695_),
    .A(_03692_),
    .Y(_03778_));
 sg13g2_o21ai_1 _09529_ (.B1(_03778_),
    .Y(_03779_),
    .A1(net74),
    .A2(_03777_));
 sg13g2_a21o_1 _09530_ (.A2(_03692_),
    .A1(net281),
    .B1(_03123_),
    .X(_03780_));
 sg13g2_a21oi_1 _09531_ (.A1(net63),
    .A2(_03780_),
    .Y(_03781_),
    .B1(_00874_));
 sg13g2_a21oi_1 _09532_ (.A1(net63),
    .A2(_03779_),
    .Y(_00610_),
    .B1(_03781_));
 sg13g2_a21o_1 _09533_ (.A2(_00902_),
    .A1(_03692_),
    .B1(net73),
    .X(_03782_));
 sg13g2_a21oi_1 _09534_ (.A1(_03712_),
    .A2(_03782_),
    .Y(_03783_),
    .B1(net237));
 sg13g2_nand3_1 _09535_ (.B(net100),
    .C(_03775_),
    .A(net161),
    .Y(_03784_));
 sg13g2_o21ai_1 _09536_ (.B1(_03784_),
    .Y(_03785_),
    .A1(net91),
    .A2(_03491_));
 sg13g2_nand3_1 _09537_ (.B(_03692_),
    .C(_00902_),
    .A(net237),
    .Y(_03786_));
 sg13g2_nand2_1 _09538_ (.Y(_03787_),
    .A(_03695_),
    .B(_03786_));
 sg13g2_nand2_1 _09539_ (.Y(_03788_),
    .A(_03711_),
    .B(_03787_));
 sg13g2_a21oi_1 _09540_ (.A1(net73),
    .A2(_03785_),
    .Y(_03789_),
    .B1(_03788_));
 sg13g2_nor2_1 _09541_ (.A(_03783_),
    .B(_03789_),
    .Y(_00611_));
 sg13g2_or2_1 _09542_ (.X(_03790_),
    .B(net89),
    .A(_03180_));
 sg13g2_a221oi_1 _09543_ (.B2(net155),
    .C1(_03209_),
    .B1(_03790_),
    .A1(_03483_),
    .Y(_03791_),
    .A2(_03493_));
 sg13g2_nand4_1 _09544_ (.B(_00902_),
    .C(_00869_),
    .A(_03692_),
    .Y(_03792_),
    .D(_03695_));
 sg13g2_o21ai_1 _09545_ (.B1(_03792_),
    .Y(_03793_),
    .A1(net74),
    .A2(_03791_));
 sg13g2_a22oi_1 _09546_ (.Y(_00612_),
    .B1(_03793_),
    .B2(_03712_),
    .A2(_03788_),
    .A1(_00938_));
 sg13g2_and2_1 _09547_ (.A(net230),
    .B(_01637_),
    .X(_03794_));
 sg13g2_a21oi_1 _09548_ (.A1(_01659_),
    .A2(_01596_),
    .Y(_03795_),
    .B1(_03794_));
 sg13g2_nor2_1 _09549_ (.A(_01654_),
    .B(_03795_),
    .Y(_03796_));
 sg13g2_buf_1 _09550_ (.A(_03796_),
    .X(_03797_));
 sg13g2_inv_1 _09551_ (.Y(_03798_),
    .A(_01654_));
 sg13g2_and4_1 _09552_ (.A(_01659_),
    .B(_01596_),
    .C(_03798_),
    .D(_01638_),
    .X(_03799_));
 sg13g2_buf_1 _09553_ (.A(_03799_),
    .X(_03800_));
 sg13g2_nor2_1 _09554_ (.A(_01356_),
    .B(_03800_),
    .Y(_03801_));
 sg13g2_buf_1 _09555_ (.A(_03801_),
    .X(_03802_));
 sg13g2_buf_1 _09556_ (.A(_03802_),
    .X(_03803_));
 sg13g2_nand3_1 _09557_ (.B(net69),
    .C(net50),
    .A(\addr[0] ),
    .Y(_03804_));
 sg13g2_nand2b_1 _09558_ (.Y(_03805_),
    .B(_03798_),
    .A_N(_03795_));
 sg13g2_buf_1 _09559_ (.A(_03805_),
    .X(_03806_));
 sg13g2_buf_1 _09560_ (.A(net68),
    .X(_03807_));
 sg13g2_buf_2 _09561_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .X(_03808_));
 sg13g2_inv_1 _09562_ (.Y(_03809_),
    .A(net311));
 sg13g2_nor3_1 _09563_ (.A(net275),
    .B(net312),
    .C(_03809_),
    .Y(_03810_));
 sg13g2_buf_1 _09564_ (.A(_03810_),
    .X(_03811_));
 sg13g2_nand2_1 _09565_ (.Y(_03812_),
    .A(_03808_),
    .B(_03811_));
 sg13g2_buf_2 _09566_ (.A(_03812_),
    .X(_03813_));
 sg13g2_buf_1 _09567_ (.A(_03813_),
    .X(_03814_));
 sg13g2_nand3_1 _09568_ (.B(net62),
    .C(net165),
    .A(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .Y(_03815_));
 sg13g2_nand2_1 _09569_ (.Y(_00618_),
    .A(_03804_),
    .B(_03815_));
 sg13g2_and2_1 _09570_ (.A(_03808_),
    .B(_03811_),
    .X(_03816_));
 sg13g2_buf_1 _09571_ (.A(_03816_),
    .X(_03817_));
 sg13g2_nor2_1 _09572_ (.A(net69),
    .B(_03817_),
    .Y(_03818_));
 sg13g2_buf_1 _09573_ (.A(_03818_),
    .X(_03819_));
 sg13g2_buf_1 _09574_ (.A(\i_tinyqv.cpu.was_early_branch ),
    .X(_03820_));
 sg13g2_buf_1 _09575_ (.A(net294),
    .X(_03821_));
 sg13g2_and2_1 _09576_ (.A(net333),
    .B(net329),
    .X(_03822_));
 sg13g2_a22oi_1 _09577_ (.Y(_03823_),
    .B1(_01067_),
    .B2(_01099_),
    .A2(net330),
    .A1(_01026_));
 sg13g2_nor2_1 _09578_ (.A(_01026_),
    .B(net330),
    .Y(_03824_));
 sg13g2_nor2_1 _09579_ (.A(net333),
    .B(net329),
    .Y(_03825_));
 sg13g2_nor3_1 _09580_ (.A(_03823_),
    .B(_03824_),
    .C(_03825_),
    .Y(_03826_));
 sg13g2_or2_1 _09581_ (.X(_03827_),
    .B(_01112_),
    .A(_01179_));
 sg13g2_o21ai_1 _09582_ (.B1(_03827_),
    .Y(_03828_),
    .A1(_03822_),
    .A2(_03826_));
 sg13g2_nand2_1 _09583_ (.Y(_03829_),
    .A(_01179_),
    .B(_01112_));
 sg13g2_nor2_1 _09584_ (.A(net296),
    .B(_01100_),
    .Y(_03830_));
 sg13g2_nor2_1 _09585_ (.A(_00831_),
    .B(_00960_),
    .Y(_03831_));
 sg13g2_nor2_1 _09586_ (.A(_03830_),
    .B(_03831_),
    .Y(_03832_));
 sg13g2_nand2_1 _09587_ (.Y(_03833_),
    .A(_00915_),
    .B(_03832_));
 sg13g2_nand2_1 _09588_ (.Y(_03834_),
    .A(net260),
    .B(_03832_));
 sg13g2_a22oi_1 _09589_ (.Y(_03835_),
    .B1(_03833_),
    .B2(_03834_),
    .A2(_03829_),
    .A1(_03828_));
 sg13g2_buf_1 _09590_ (.A(_03835_),
    .X(_03836_));
 sg13g2_nand2_1 _09591_ (.Y(_03837_),
    .A(net260),
    .B(_00915_));
 sg13g2_nand2_1 _09592_ (.Y(_03838_),
    .A(net296),
    .B(_01100_));
 sg13g2_nor2_1 _09593_ (.A(_03838_),
    .B(_03831_),
    .Y(_03839_));
 sg13g2_o21ai_1 _09594_ (.B1(_03839_),
    .Y(_03840_),
    .A1(_01021_),
    .A2(_00915_));
 sg13g2_o21ai_1 _09595_ (.B1(_03840_),
    .Y(_03841_),
    .A1(_03831_),
    .A2(_03837_));
 sg13g2_buf_1 _09596_ (.A(_03841_),
    .X(_03842_));
 sg13g2_nor2_1 _09597_ (.A(_01547_),
    .B(_01066_),
    .Y(_03843_));
 sg13g2_and2_1 _09598_ (.A(net261),
    .B(_00960_),
    .X(_03844_));
 sg13g2_buf_1 _09599_ (.A(_03844_),
    .X(_03845_));
 sg13g2_or2_1 _09600_ (.X(_03846_),
    .B(_03845_),
    .A(_03843_));
 sg13g2_or4_1 _09601_ (.A(net259),
    .B(_03836_),
    .C(_03842_),
    .D(_03846_),
    .X(_03847_));
 sg13g2_or4_1 _09602_ (.A(_01110_),
    .B(_03836_),
    .C(_03842_),
    .D(_03846_),
    .X(_03848_));
 sg13g2_nor3_1 _09603_ (.A(_01110_),
    .B(net259),
    .C(_03843_),
    .Y(_03849_));
 sg13g2_a21oi_1 _09604_ (.A1(_01547_),
    .A2(_01066_),
    .Y(_03850_),
    .B1(_03849_));
 sg13g2_and3_1 _09605_ (.X(_03851_),
    .A(_03847_),
    .B(_03848_),
    .C(_03850_));
 sg13g2_buf_1 _09606_ (.A(_03851_),
    .X(_03852_));
 sg13g2_xor2_1 _09607_ (.B(net257),
    .A(net325),
    .X(_03853_));
 sg13g2_xnor2_1 _09608_ (.Y(_03854_),
    .A(_03852_),
    .B(_03853_));
 sg13g2_nand2_1 _09609_ (.Y(_03855_),
    .A(net333),
    .B(_01568_));
 sg13g2_buf_2 _09610_ (.A(_03855_),
    .X(_03856_));
 sg13g2_nor2_2 _09611_ (.A(_02615_),
    .B(_03856_),
    .Y(_03857_));
 sg13g2_nand3_1 _09612_ (.B(_02621_),
    .C(_03857_),
    .A(_01065_),
    .Y(_03858_));
 sg13g2_xnor2_1 _09613_ (.Y(_03859_),
    .A(net325),
    .B(_03858_));
 sg13g2_nor2_1 _09614_ (.A(net294),
    .B(_03859_),
    .Y(_03860_));
 sg13g2_a21oi_1 _09615_ (.A1(net250),
    .A2(_03854_),
    .Y(_03861_),
    .B1(_03860_));
 sg13g2_nand4_1 _09616_ (.B(_01596_),
    .C(_03798_),
    .A(_01659_),
    .Y(_03862_),
    .D(_01638_));
 sg13g2_buf_1 _09617_ (.A(_03862_),
    .X(_03863_));
 sg13g2_nand2_1 _09618_ (.Y(_03864_),
    .A(_01355_),
    .B(net72));
 sg13g2_buf_1 _09619_ (.A(_03864_),
    .X(_03865_));
 sg13g2_mux2_1 _09620_ (.A0(\addr[10] ),
    .A1(_03861_),
    .S(net61),
    .X(_03866_));
 sg13g2_buf_1 _09621_ (.A(_03817_),
    .X(_03867_));
 sg13g2_and2_1 _09622_ (.A(\i_tinyqv.mem.q_ctrl.addr[6] ),
    .B(net164),
    .X(_03868_));
 sg13g2_a221oi_1 _09623_ (.B2(net69),
    .C1(_03868_),
    .B1(_03866_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .Y(_03869_),
    .A2(net49));
 sg13g2_inv_1 _09624_ (.Y(_00619_),
    .A(_03869_));
 sg13g2_buf_1 _09625_ (.A(net68),
    .X(_03870_));
 sg13g2_nor2_1 _09626_ (.A(net257),
    .B(_03852_),
    .Y(_03871_));
 sg13g2_a21oi_1 _09627_ (.A1(net257),
    .A2(_03852_),
    .Y(_03872_),
    .B1(net325));
 sg13g2_nor2_1 _09628_ (.A(_03871_),
    .B(_03872_),
    .Y(_03873_));
 sg13g2_xor2_1 _09629_ (.B(net328),
    .A(net262),
    .X(_03874_));
 sg13g2_xnor2_1 _09630_ (.Y(_03875_),
    .A(_03873_),
    .B(_03874_));
 sg13g2_buf_1 _09631_ (.A(net294),
    .X(_03876_));
 sg13g2_buf_1 _09632_ (.A(net249),
    .X(_03877_));
 sg13g2_nor3_1 _09633_ (.A(_02603_),
    .B(_02814_),
    .C(_03856_),
    .Y(_03878_));
 sg13g2_nor2b_1 _09634_ (.A(_02820_),
    .B_N(_03878_),
    .Y(_03879_));
 sg13g2_xnor2_1 _09635_ (.Y(_03880_),
    .A(_00841_),
    .B(_03879_));
 sg13g2_nor2_1 _09636_ (.A(net250),
    .B(_03880_),
    .Y(_03881_));
 sg13g2_a221oi_1 _09637_ (.B2(net227),
    .C1(_03881_),
    .B1(_03875_),
    .A1(_01355_),
    .Y(_03882_),
    .A2(net72));
 sg13g2_a21oi_1 _09638_ (.A1(\addr[11] ),
    .A2(net50),
    .Y(_03883_),
    .B1(_03882_));
 sg13g2_a22oi_1 _09639_ (.Y(_03884_),
    .B1(net49),
    .B2(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .A2(net164),
    .A1(\i_tinyqv.mem.q_ctrl.addr[7] ));
 sg13g2_o21ai_1 _09640_ (.B1(_03884_),
    .Y(_00620_),
    .A1(net60),
    .A2(_03883_));
 sg13g2_xnor2_1 _09641_ (.Y(_03885_),
    .A(net297),
    .B(_01113_));
 sg13g2_a21o_1 _09642_ (.A2(_03873_),
    .A1(net328),
    .B1(net262),
    .X(_03886_));
 sg13g2_o21ai_1 _09643_ (.B1(_03886_),
    .Y(_03887_),
    .A1(net328),
    .A2(_03873_));
 sg13g2_xnor2_1 _09644_ (.Y(_03888_),
    .A(_03885_),
    .B(_03887_));
 sg13g2_nand3_1 _09645_ (.B(_02610_),
    .C(_03857_),
    .A(_02608_),
    .Y(_03889_));
 sg13g2_xnor2_1 _09646_ (.Y(_03890_),
    .A(_02607_),
    .B(_03889_));
 sg13g2_nor2_1 _09647_ (.A(_03820_),
    .B(_03890_),
    .Y(_03891_));
 sg13g2_a21oi_1 _09648_ (.A1(net250),
    .A2(_03888_),
    .Y(_03892_),
    .B1(_03891_));
 sg13g2_mux2_1 _09649_ (.A0(\addr[12] ),
    .A1(_03892_),
    .S(net61),
    .X(_03893_));
 sg13g2_and2_1 _09650_ (.A(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .B(net164),
    .X(_03894_));
 sg13g2_a221oi_1 _09651_ (.B2(net69),
    .C1(_03894_),
    .B1(_03893_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .Y(_03895_),
    .A2(net49));
 sg13g2_inv_1 _09652_ (.Y(_00621_),
    .A(_03895_));
 sg13g2_buf_1 _09653_ (.A(_03802_),
    .X(_03896_));
 sg13g2_buf_1 _09654_ (.A(_03820_),
    .X(_03897_));
 sg13g2_nor2_1 _09655_ (.A(net297),
    .B(_01113_),
    .Y(_03898_));
 sg13g2_or2_1 _09656_ (.X(_03899_),
    .B(net257),
    .A(net325));
 sg13g2_nor3_1 _09657_ (.A(_01101_),
    .B(_00920_),
    .C(_01065_),
    .Y(_03900_));
 sg13g2_nor3_1 _09658_ (.A(_00841_),
    .B(_03900_),
    .C(_03898_),
    .Y(_03901_));
 sg13g2_a21oi_1 _09659_ (.A1(net328),
    .A2(_03899_),
    .Y(_03902_),
    .B1(_03901_));
 sg13g2_nor3_1 _09660_ (.A(_02647_),
    .B(_03898_),
    .C(_03902_),
    .Y(_03903_));
 sg13g2_nand4_1 _09661_ (.B(_03848_),
    .C(_03850_),
    .A(_03847_),
    .Y(_03904_),
    .D(_03903_));
 sg13g2_nand2_1 _09662_ (.Y(_03905_),
    .A(net325),
    .B(_03901_));
 sg13g2_or3_1 _09663_ (.A(net257),
    .B(_01178_),
    .C(_03843_),
    .X(_03906_));
 sg13g2_nor4_1 _09664_ (.A(_03845_),
    .B(_03836_),
    .C(_03842_),
    .D(_03906_),
    .Y(_03907_));
 sg13g2_or3_1 _09665_ (.A(_01110_),
    .B(net257),
    .C(_03843_),
    .X(_03908_));
 sg13g2_nor4_1 _09666_ (.A(_03845_),
    .B(_03836_),
    .C(_03842_),
    .D(_03908_),
    .Y(_03909_));
 sg13g2_nor2_1 _09667_ (.A(net259),
    .B(_03908_),
    .Y(_03910_));
 sg13g2_or4_1 _09668_ (.A(_03905_),
    .B(_03907_),
    .C(_03909_),
    .D(_03910_),
    .X(_03911_));
 sg13g2_buf_1 _09669_ (.A(_03911_),
    .X(_03912_));
 sg13g2_a21o_1 _09670_ (.A2(_02646_),
    .A1(net325),
    .B1(_00840_),
    .X(_03913_));
 sg13g2_a22oi_1 _09671_ (.Y(_03914_),
    .B1(_03913_),
    .B2(_00964_),
    .A2(_01113_),
    .A1(net297));
 sg13g2_or2_1 _09672_ (.X(_03915_),
    .B(_03914_),
    .A(_03898_));
 sg13g2_buf_1 _09673_ (.A(_03915_),
    .X(_03916_));
 sg13g2_nand3_1 _09674_ (.B(_03912_),
    .C(_03916_),
    .A(_03904_),
    .Y(_03917_));
 sg13g2_xnor2_1 _09675_ (.Y(_03918_),
    .A(_01058_),
    .B(_01102_));
 sg13g2_xnor2_1 _09676_ (.Y(_03919_),
    .A(_03917_),
    .B(_03918_));
 sg13g2_inv_1 _09677_ (.Y(_03920_),
    .A(_01058_));
 sg13g2_nand3_1 _09678_ (.B(net297),
    .C(_03879_),
    .A(net262),
    .Y(_03921_));
 sg13g2_xnor2_1 _09679_ (.Y(_03922_),
    .A(_03920_),
    .B(_03921_));
 sg13g2_nor2_1 _09680_ (.A(net249),
    .B(_03922_),
    .Y(_03923_));
 sg13g2_a21oi_1 _09681_ (.A1(net248),
    .A2(_03919_),
    .Y(_03924_),
    .B1(_03923_));
 sg13g2_nor2_1 _09682_ (.A(net48),
    .B(_03924_),
    .Y(_03925_));
 sg13g2_a21oi_1 _09683_ (.A1(\addr[13] ),
    .A2(net50),
    .Y(_03926_),
    .B1(_03925_));
 sg13g2_buf_1 _09684_ (.A(net68),
    .X(_03927_));
 sg13g2_mux2_1 _09685_ (.A0(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .S(net165),
    .X(_03928_));
 sg13g2_nand2_1 _09686_ (.Y(_03929_),
    .A(net59),
    .B(_03928_));
 sg13g2_o21ai_1 _09687_ (.B1(_03929_),
    .Y(_00622_),
    .A1(net60),
    .A2(_03926_));
 sg13g2_buf_1 _09688_ (.A(_03802_),
    .X(_03930_));
 sg13g2_xor2_1 _09689_ (.B(_00916_),
    .A(net326),
    .X(_03931_));
 sg13g2_nand4_1 _09690_ (.B(_03904_),
    .C(_03912_),
    .A(_03920_),
    .Y(_03932_),
    .D(_03916_));
 sg13g2_inv_1 _09691_ (.Y(_03933_),
    .A(_01102_));
 sg13g2_nand2_1 _09692_ (.Y(_03934_),
    .A(_03920_),
    .B(_03933_));
 sg13g2_nand4_1 _09693_ (.B(_03904_),
    .C(_03912_),
    .A(_03933_),
    .Y(_03935_),
    .D(_03916_));
 sg13g2_nand3_1 _09694_ (.B(_03934_),
    .C(_03935_),
    .A(_03932_),
    .Y(_03936_));
 sg13g2_xnor2_1 _09695_ (.Y(_03937_),
    .A(_03931_),
    .B(_03936_));
 sg13g2_nand2_1 _09696_ (.Y(_03938_),
    .A(_02629_),
    .B(_03857_));
 sg13g2_xnor2_1 _09697_ (.Y(_03939_),
    .A(_02882_),
    .B(_03938_));
 sg13g2_nor2_1 _09698_ (.A(net249),
    .B(_03939_),
    .Y(_03940_));
 sg13g2_a21oi_1 _09699_ (.A1(net248),
    .A2(_03937_),
    .Y(_03941_),
    .B1(_03940_));
 sg13g2_nor2_1 _09700_ (.A(net47),
    .B(_03941_),
    .Y(_03942_));
 sg13g2_a21oi_1 _09701_ (.A1(\addr[14] ),
    .A2(net50),
    .Y(_03943_),
    .B1(_03942_));
 sg13g2_mux2_1 _09702_ (.A0(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .S(net165),
    .X(_03944_));
 sg13g2_nand2_1 _09703_ (.Y(_03945_),
    .A(net62),
    .B(_03944_));
 sg13g2_o21ai_1 _09704_ (.B1(_03945_),
    .Y(_00623_),
    .A1(net60),
    .A2(_03943_));
 sg13g2_nand2_1 _09705_ (.Y(_03946_),
    .A(_02829_),
    .B(_03879_));
 sg13g2_nand2_1 _09706_ (.Y(_03947_),
    .A(net326),
    .B(_00916_));
 sg13g2_nor2_1 _09707_ (.A(net326),
    .B(_00916_),
    .Y(_03948_));
 sg13g2_a21oi_1 _09708_ (.A1(_03936_),
    .A2(_03947_),
    .Y(_03949_),
    .B1(_03948_));
 sg13g2_xnor2_1 _09709_ (.Y(_03950_),
    .A(_00961_),
    .B(_03949_));
 sg13g2_mux2_1 _09710_ (.A0(_03946_),
    .A1(_03950_),
    .S(net294),
    .X(_03951_));
 sg13g2_xnor2_1 _09711_ (.Y(_03952_),
    .A(_02626_),
    .B(_03951_));
 sg13g2_and2_1 _09712_ (.A(\addr[15] ),
    .B(_03802_),
    .X(_03953_));
 sg13g2_a21oi_1 _09713_ (.A1(net61),
    .A2(_03952_),
    .Y(_03954_),
    .B1(_03953_));
 sg13g2_mux2_1 _09714_ (.A0(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .S(_03814_),
    .X(_03955_));
 sg13g2_nand2_1 _09715_ (.Y(_03956_),
    .A(net62),
    .B(_03955_));
 sg13g2_o21ai_1 _09716_ (.B1(_03956_),
    .Y(_00624_),
    .A1(net60),
    .A2(_03954_));
 sg13g2_nor2b_1 _09717_ (.A(_03948_),
    .B_N(_00961_),
    .Y(_03957_));
 sg13g2_nand4_1 _09718_ (.B(_03934_),
    .C(_03935_),
    .A(_03932_),
    .Y(_03958_),
    .D(_03957_));
 sg13g2_nor2b_1 _09719_ (.A(_03948_),
    .B_N(net258),
    .Y(_03959_));
 sg13g2_nand4_1 _09720_ (.B(_03934_),
    .C(_03935_),
    .A(_03932_),
    .Y(_03960_),
    .D(_03959_));
 sg13g2_nand2_1 _09721_ (.Y(_03961_),
    .A(net258),
    .B(_00961_));
 sg13g2_and2_1 _09722_ (.A(net326),
    .B(_00916_),
    .X(_03962_));
 sg13g2_o21ai_1 _09723_ (.B1(_03962_),
    .Y(_03963_),
    .A1(net258),
    .A2(_00961_));
 sg13g2_and2_1 _09724_ (.A(_03961_),
    .B(_03963_),
    .X(_03964_));
 sg13g2_buf_1 _09725_ (.A(_03964_),
    .X(_03965_));
 sg13g2_nand3_1 _09726_ (.B(_03960_),
    .C(_03965_),
    .A(_03958_),
    .Y(_03966_));
 sg13g2_buf_1 _09727_ (.A(_03966_),
    .X(_03967_));
 sg13g2_xnor2_1 _09728_ (.Y(_03968_),
    .A(net295),
    .B(_01109_));
 sg13g2_xnor2_1 _09729_ (.Y(_03969_),
    .A(_03967_),
    .B(_03968_));
 sg13g2_nor2_1 _09730_ (.A(_02627_),
    .B(_03938_),
    .Y(_03970_));
 sg13g2_xnor2_1 _09731_ (.Y(_03971_),
    .A(_02625_),
    .B(_03970_));
 sg13g2_nor2_1 _09732_ (.A(net249),
    .B(_03971_),
    .Y(_03972_));
 sg13g2_a21oi_1 _09733_ (.A1(net248),
    .A2(_03969_),
    .Y(_03973_),
    .B1(_03972_));
 sg13g2_nor2_1 _09734_ (.A(net47),
    .B(_03973_),
    .Y(_03974_));
 sg13g2_a21oi_1 _09735_ (.A1(\addr[16] ),
    .A2(net50),
    .Y(_03975_),
    .B1(_03974_));
 sg13g2_mux2_1 _09736_ (.A0(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .S(_03814_),
    .X(_03976_));
 sg13g2_nand2_1 _09737_ (.Y(_03977_),
    .A(_03807_),
    .B(_03976_));
 sg13g2_o21ai_1 _09738_ (.B1(_03977_),
    .Y(_00625_),
    .A1(_03870_),
    .A2(_03975_));
 sg13g2_nor2_1 _09739_ (.A(net295),
    .B(_01109_),
    .Y(_03978_));
 sg13g2_and2_1 _09740_ (.A(net295),
    .B(_01109_),
    .X(_03979_));
 sg13g2_nor2_1 _09741_ (.A(_03967_),
    .B(_03979_),
    .Y(_03980_));
 sg13g2_nor2_1 _09742_ (.A(_03978_),
    .B(_03980_),
    .Y(_03981_));
 sg13g2_xnor2_1 _09743_ (.Y(_03982_),
    .A(_01096_),
    .B(_03981_));
 sg13g2_nor2b_1 _09744_ (.A(_03982_),
    .B_N(\i_tinyqv.cpu.was_early_branch ),
    .Y(_03983_));
 sg13g2_nor3_1 _09745_ (.A(net294),
    .B(_02834_),
    .C(_03946_),
    .Y(_03984_));
 sg13g2_nor2_1 _09746_ (.A(_03983_),
    .B(_03984_),
    .Y(_03985_));
 sg13g2_xor2_1 _09747_ (.B(_03985_),
    .A(_01062_),
    .X(_03986_));
 sg13g2_nor2_1 _09748_ (.A(net47),
    .B(_03986_),
    .Y(_03987_));
 sg13g2_a21oi_1 _09749_ (.A1(\addr[17] ),
    .A2(net50),
    .Y(_03988_),
    .B1(_03987_));
 sg13g2_mux2_1 _09750_ (.A0(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .S(_03813_),
    .X(_03989_));
 sg13g2_nand2_1 _09751_ (.Y(_03990_),
    .A(net62),
    .B(_03989_));
 sg13g2_o21ai_1 _09752_ (.B1(_03990_),
    .Y(_00626_),
    .A1(net60),
    .A2(_03988_));
 sg13g2_xor2_1 _09753_ (.B(_00921_),
    .A(net327),
    .X(_03991_));
 sg13g2_a21o_1 _09754_ (.A2(_03981_),
    .A1(net324),
    .B1(_01096_),
    .X(_03992_));
 sg13g2_o21ai_1 _09755_ (.B1(_03992_),
    .Y(_03993_),
    .A1(net324),
    .A2(_03981_));
 sg13g2_xnor2_1 _09756_ (.Y(_03994_),
    .A(_03991_),
    .B(_03993_));
 sg13g2_nor2_1 _09757_ (.A(_02634_),
    .B(_03938_),
    .Y(_03995_));
 sg13g2_xnor2_1 _09758_ (.Y(_03996_),
    .A(_01017_),
    .B(_03995_));
 sg13g2_nor2_1 _09759_ (.A(net249),
    .B(_03996_),
    .Y(_03997_));
 sg13g2_a21oi_1 _09760_ (.A1(net248),
    .A2(_03994_),
    .Y(_03998_),
    .B1(_03997_));
 sg13g2_nor2_1 _09761_ (.A(net47),
    .B(_03998_),
    .Y(_03999_));
 sg13g2_a21oi_1 _09762_ (.A1(\addr[18] ),
    .A2(_03803_),
    .Y(_04000_),
    .B1(_03999_));
 sg13g2_mux2_1 _09763_ (.A0(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .S(_03813_),
    .X(_04001_));
 sg13g2_nand2_1 _09764_ (.Y(_04002_),
    .A(_03807_),
    .B(_04001_));
 sg13g2_o21ai_1 _09765_ (.B1(_04002_),
    .Y(_00627_),
    .A1(_03870_),
    .A2(_04000_));
 sg13g2_a221oi_1 _09766_ (.B2(_03979_),
    .C1(net324),
    .B1(_01096_),
    .A1(net327),
    .Y(_04003_),
    .A2(_00921_));
 sg13g2_nor2b_1 _09767_ (.A(_03978_),
    .B_N(_01096_),
    .Y(_04004_));
 sg13g2_nand2_1 _09768_ (.Y(_04005_),
    .A(_03967_),
    .B(_04004_));
 sg13g2_nand2_1 _09769_ (.Y(_04006_),
    .A(net295),
    .B(_01109_));
 sg13g2_nor2_1 _09770_ (.A(_00921_),
    .B(_01096_),
    .Y(_04007_));
 sg13g2_and2_1 _09771_ (.A(_04006_),
    .B(_04007_),
    .X(_04008_));
 sg13g2_nand4_1 _09772_ (.B(_03960_),
    .C(_03965_),
    .A(_03958_),
    .Y(_04009_),
    .D(_04008_));
 sg13g2_nor2_1 _09773_ (.A(net327),
    .B(_01096_),
    .Y(_04010_));
 sg13g2_and2_1 _09774_ (.A(_04006_),
    .B(_04010_),
    .X(_04011_));
 sg13g2_nand4_1 _09775_ (.B(_03960_),
    .C(_03965_),
    .A(_03958_),
    .Y(_04012_),
    .D(_04011_));
 sg13g2_o21ai_1 _09776_ (.B1(_03978_),
    .Y(_04013_),
    .A1(_04007_),
    .A2(_04010_));
 sg13g2_or2_1 _09777_ (.X(_04014_),
    .B(_00921_),
    .A(net327));
 sg13g2_nand4_1 _09778_ (.B(_04012_),
    .C(_04013_),
    .A(_04009_),
    .Y(_04015_),
    .D(_04014_));
 sg13g2_a21oi_2 _09779_ (.B1(_04015_),
    .Y(_04016_),
    .A2(_04005_),
    .A1(_04003_));
 sg13g2_xnor2_1 _09780_ (.Y(_04017_),
    .A(net334),
    .B(_00965_));
 sg13g2_xnor2_1 _09781_ (.Y(_04018_),
    .A(_04016_),
    .B(_04017_));
 sg13g2_nor2_1 _09782_ (.A(_02825_),
    .B(_03946_),
    .Y(_04019_));
 sg13g2_xnor2_1 _09783_ (.Y(_04020_),
    .A(_00836_),
    .B(_04019_));
 sg13g2_nor2_1 _09784_ (.A(_03876_),
    .B(_04020_),
    .Y(_04021_));
 sg13g2_a21oi_1 _09785_ (.A1(_03897_),
    .A2(_04018_),
    .Y(_04022_),
    .B1(_04021_));
 sg13g2_nor2_1 _09786_ (.A(net47),
    .B(_04022_),
    .Y(_04023_));
 sg13g2_a21oi_1 _09787_ (.A1(\addr[19] ),
    .A2(net48),
    .Y(_04024_),
    .B1(_04023_));
 sg13g2_mux2_1 _09788_ (.A0(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .S(_03813_),
    .X(_04025_));
 sg13g2_nand2_1 _09789_ (.Y(_04026_),
    .A(net62),
    .B(_04025_));
 sg13g2_o21ai_1 _09790_ (.B1(_04026_),
    .Y(_00628_),
    .A1(_03927_),
    .A2(_04024_));
 sg13g2_xnor2_1 _09791_ (.Y(_04027_),
    .A(_01067_),
    .B(net255));
 sg13g2_nor2_1 _09792_ (.A(_01586_),
    .B(net250),
    .Y(_04028_));
 sg13g2_a221oi_1 _09793_ (.B2(net227),
    .C1(_04028_),
    .B1(_04027_),
    .A1(_01355_),
    .Y(_04029_),
    .A2(net72));
 sg13g2_a21oi_1 _09794_ (.A1(\addr[1] ),
    .A2(net48),
    .Y(_04030_),
    .B1(_04029_));
 sg13g2_nand3_1 _09795_ (.B(net68),
    .C(net165),
    .A(\i_tinyqv.mem.q_ctrl.addr[1] ),
    .Y(_04031_));
 sg13g2_o21ai_1 _09796_ (.B1(_04031_),
    .Y(_00629_),
    .A1(net59),
    .A2(_04030_));
 sg13g2_and2_1 _09797_ (.A(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .B(_03817_),
    .X(_04032_));
 sg13g2_a21oi_1 _09798_ (.A1(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .A2(net165),
    .Y(_04033_),
    .B1(_04032_));
 sg13g2_a21oi_1 _09799_ (.A1(\addr[20] ),
    .A2(net50),
    .Y(_04034_),
    .B1(net62));
 sg13g2_nor2_1 _09800_ (.A(_02636_),
    .B(_03856_),
    .Y(_04035_));
 sg13g2_xnor2_1 _09801_ (.Y(_04036_),
    .A(_01175_),
    .B(_04035_));
 sg13g2_xnor2_1 _09802_ (.Y(_04037_),
    .A(_01175_),
    .B(_01114_));
 sg13g2_a21oi_1 _09803_ (.A1(_00965_),
    .A2(_04016_),
    .Y(_04038_),
    .B1(net334));
 sg13g2_nor2_1 _09804_ (.A(_00965_),
    .B(_04016_),
    .Y(_04039_));
 sg13g2_nor2_1 _09805_ (.A(_04038_),
    .B(_04039_),
    .Y(_04040_));
 sg13g2_xnor2_1 _09806_ (.Y(_04041_),
    .A(_04037_),
    .B(_04040_));
 sg13g2_nand2_1 _09807_ (.Y(_04042_),
    .A(net227),
    .B(_04041_));
 sg13g2_o21ai_1 _09808_ (.B1(_04042_),
    .Y(_04043_),
    .A1(net227),
    .A2(_04036_));
 sg13g2_nand2_1 _09809_ (.Y(_04044_),
    .A(net61),
    .B(_04043_));
 sg13g2_a22oi_1 _09810_ (.Y(_00630_),
    .B1(_04034_),
    .B2(_04044_),
    .A2(_04033_),
    .A1(net60));
 sg13g2_and2_1 _09811_ (.A(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .B(_03817_),
    .X(_04045_));
 sg13g2_a21oi_1 _09812_ (.A1(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .A2(net165),
    .Y(_04046_),
    .B1(_04045_));
 sg13g2_a21oi_1 _09813_ (.A1(\addr[21] ),
    .A2(net50),
    .Y(_04047_),
    .B1(net68));
 sg13g2_nor2_1 _09814_ (.A(_02603_),
    .B(_03856_),
    .Y(_04048_));
 sg13g2_nand2b_1 _09815_ (.Y(_04049_),
    .B(_04048_),
    .A_N(_02831_));
 sg13g2_nand2_1 _09816_ (.Y(_04050_),
    .A(_00961_),
    .B(_04004_));
 sg13g2_nand2_1 _09817_ (.Y(_04051_),
    .A(net258),
    .B(_04004_));
 sg13g2_a221oi_1 _09818_ (.B2(_04051_),
    .C1(_03948_),
    .B1(_04050_),
    .A1(_03936_),
    .Y(_04052_),
    .A2(_03947_));
 sg13g2_nand2b_1 _09819_ (.Y(_04053_),
    .B(_04004_),
    .A_N(_03961_));
 sg13g2_nand2_1 _09820_ (.Y(_04054_),
    .A(_04003_),
    .B(_04053_));
 sg13g2_nor2_1 _09821_ (.A(_01175_),
    .B(_01114_),
    .Y(_04055_));
 sg13g2_nor2b_1 _09822_ (.A(_04055_),
    .B_N(_00965_),
    .Y(_04056_));
 sg13g2_o21ai_1 _09823_ (.B1(_04056_),
    .Y(_04057_),
    .A1(_04052_),
    .A2(_04054_));
 sg13g2_nor2b_1 _09824_ (.A(_04055_),
    .B_N(net334),
    .Y(_04058_));
 sg13g2_o21ai_1 _09825_ (.B1(_04058_),
    .Y(_04059_),
    .A1(_04052_),
    .A2(_04054_));
 sg13g2_a21oi_1 _09826_ (.A1(_04057_),
    .A2(_04059_),
    .Y(_04060_),
    .B1(_04015_));
 sg13g2_nand2_1 _09827_ (.Y(_04061_),
    .A(net334),
    .B(_00965_));
 sg13g2_nand2_1 _09828_ (.Y(_04062_),
    .A(_01175_),
    .B(_01114_));
 sg13g2_o21ai_1 _09829_ (.B1(_04062_),
    .Y(_04063_),
    .A1(_04055_),
    .A2(_04061_));
 sg13g2_nor2_1 _09830_ (.A(_04060_),
    .B(_04063_),
    .Y(_04064_));
 sg13g2_xor2_1 _09831_ (.B(_04064_),
    .A(_01097_),
    .X(_04065_));
 sg13g2_nand2b_1 _09832_ (.Y(_04066_),
    .B(net294),
    .A_N(_04065_));
 sg13g2_o21ai_1 _09833_ (.B1(_04066_),
    .Y(_04067_),
    .A1(net249),
    .A2(_04049_));
 sg13g2_o21ai_1 _09834_ (.B1(_03865_),
    .Y(_04068_),
    .A1(_01071_),
    .A2(_04067_));
 sg13g2_a21o_1 _09835_ (.A2(_04067_),
    .A1(_01071_),
    .B1(_04068_),
    .X(_04069_));
 sg13g2_a22oi_1 _09836_ (.Y(_00631_),
    .B1(_04047_),
    .B2(_04069_),
    .A2(_04046_),
    .A1(net60));
 sg13g2_nand2b_1 _09837_ (.Y(_04070_),
    .B(net164),
    .A_N(\i_tinyqv.mem.q_ctrl.addr[18] ));
 sg13g2_o21ai_1 _09838_ (.B1(_04070_),
    .Y(_04071_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .A2(net164));
 sg13g2_nand2_1 _09839_ (.Y(_04072_),
    .A(net323),
    .B(_01097_));
 sg13g2_nor2_1 _09840_ (.A(net323),
    .B(_01097_),
    .Y(_04073_));
 sg13g2_a21oi_1 _09841_ (.A1(_04064_),
    .A2(_04072_),
    .Y(_04074_),
    .B1(_04073_));
 sg13g2_xor2_1 _09842_ (.B(_04074_),
    .A(_00917_),
    .X(_04075_));
 sg13g2_nor3_1 _09843_ (.A(net294),
    .B(_02885_),
    .C(_03938_),
    .Y(_04076_));
 sg13g2_a21oi_1 _09844_ (.A1(_03821_),
    .A2(_04075_),
    .Y(_04077_),
    .B1(_04076_));
 sg13g2_xnor2_1 _09845_ (.Y(_04078_),
    .A(_01030_),
    .B(_04077_));
 sg13g2_nand2_1 _09846_ (.Y(_04079_),
    .A(_03865_),
    .B(_04078_));
 sg13g2_a21oi_1 _09847_ (.A1(\addr[22] ),
    .A2(_03803_),
    .Y(_04080_),
    .B1(net62));
 sg13g2_a22oi_1 _09848_ (.Y(_00632_),
    .B1(_04079_),
    .B2(_04080_),
    .A2(_04071_),
    .A1(net60));
 sg13g2_nand2_1 _09849_ (.Y(_04081_),
    .A(net69),
    .B(net61));
 sg13g2_xor2_1 _09850_ (.B(\i_tinyqv.cpu.imm[23] ),
    .A(\i_tinyqv.cpu.instr_data_start[23] ),
    .X(_04082_));
 sg13g2_a21o_1 _09851_ (.A2(_00917_),
    .A1(_01030_),
    .B1(_04074_),
    .X(_04083_));
 sg13g2_o21ai_1 _09852_ (.B1(_04083_),
    .Y(_04084_),
    .A1(_01030_),
    .A2(_00917_));
 sg13g2_xnor2_1 _09853_ (.Y(_04085_),
    .A(_04082_),
    .B(_04084_));
 sg13g2_nor2_1 _09854_ (.A(_02974_),
    .B(_03946_),
    .Y(_04086_));
 sg13g2_xor2_1 _09855_ (.B(_04086_),
    .A(_00162_),
    .X(_04087_));
 sg13g2_nor2_1 _09856_ (.A(net227),
    .B(_04087_),
    .Y(_04088_));
 sg13g2_a21oi_1 _09857_ (.A1(net227),
    .A2(_04085_),
    .Y(_04089_),
    .B1(_04088_));
 sg13g2_buf_1 _09858_ (.A(_00161_),
    .X(_04090_));
 sg13g2_nor3_1 _09859_ (.A(_04090_),
    .B(_03806_),
    .C(net61),
    .Y(_04091_));
 sg13g2_a221oi_1 _09860_ (.B2(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .C1(_04091_),
    .B1(net49),
    .A1(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .Y(_04092_),
    .A2(net164));
 sg13g2_o21ai_1 _09861_ (.B1(_04092_),
    .Y(_00633_),
    .A1(_04081_),
    .A2(_04089_));
 sg13g2_nand2_1 _09862_ (.Y(_04093_),
    .A(_01067_),
    .B(net255));
 sg13g2_xor2_1 _09863_ (.B(net330),
    .A(_01026_),
    .X(_04094_));
 sg13g2_xnor2_1 _09864_ (.Y(_04095_),
    .A(_04093_),
    .B(_04094_));
 sg13g2_nor2b_1 _09865_ (.A(net250),
    .B_N(net313),
    .Y(_04096_));
 sg13g2_a21oi_1 _09866_ (.A1(net248),
    .A2(_04095_),
    .Y(_04097_),
    .B1(_04096_));
 sg13g2_nor2_1 _09867_ (.A(net47),
    .B(_04097_),
    .Y(_04098_));
 sg13g2_a21oi_1 _09868_ (.A1(net273),
    .A2(net48),
    .Y(_04099_),
    .B1(_04098_));
 sg13g2_nand3_1 _09869_ (.B(net68),
    .C(net165),
    .A(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .Y(_04100_));
 sg13g2_o21ai_1 _09870_ (.B1(_04100_),
    .Y(_00634_),
    .A1(net59),
    .A2(_04099_));
 sg13g2_or2_1 _09871_ (.X(_04101_),
    .B(_03824_),
    .A(_03823_));
 sg13g2_xor2_1 _09872_ (.B(_00963_),
    .A(net333),
    .X(_04102_));
 sg13g2_xnor2_1 _09873_ (.Y(_04103_),
    .A(_04101_),
    .B(_04102_));
 sg13g2_xnor2_1 _09874_ (.Y(_04104_),
    .A(net333),
    .B(_01568_));
 sg13g2_nor2_1 _09875_ (.A(net249),
    .B(_04104_),
    .Y(_04105_));
 sg13g2_a21oi_1 _09876_ (.A1(net248),
    .A2(_04103_),
    .Y(_04106_),
    .B1(_04105_));
 sg13g2_nor2_1 _09877_ (.A(net47),
    .B(_04106_),
    .Y(_04107_));
 sg13g2_a21oi_1 _09878_ (.A1(net272),
    .A2(net48),
    .Y(_04108_),
    .B1(_04107_));
 sg13g2_nand3_1 _09879_ (.B(net68),
    .C(net165),
    .A(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .Y(_04109_));
 sg13g2_o21ai_1 _09880_ (.B1(_04109_),
    .Y(_00635_),
    .A1(net59),
    .A2(_04108_));
 sg13g2_nor2_1 _09881_ (.A(_03822_),
    .B(_03826_),
    .Y(_04110_));
 sg13g2_xnor2_1 _09882_ (.Y(_04111_),
    .A(_01179_),
    .B(_01112_));
 sg13g2_xnor2_1 _09883_ (.Y(_04112_),
    .A(_04110_),
    .B(_04111_));
 sg13g2_xnor2_1 _09884_ (.Y(_04113_),
    .A(_01179_),
    .B(_03856_));
 sg13g2_nor2_1 _09885_ (.A(net250),
    .B(_04113_),
    .Y(_04114_));
 sg13g2_a221oi_1 _09886_ (.B2(_03877_),
    .C1(_04114_),
    .B1(_04112_),
    .A1(_01355_),
    .Y(_04115_),
    .A2(net72));
 sg13g2_a21oi_1 _09887_ (.A1(_01697_),
    .A2(net48),
    .Y(_04116_),
    .B1(_04115_));
 sg13g2_a22oi_1 _09888_ (.Y(_04117_),
    .B1(net49),
    .B2(\i_tinyqv.mem.q_ctrl.addr[4] ),
    .A2(_03867_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[0] ));
 sg13g2_o21ai_1 _09889_ (.B1(_04117_),
    .Y(_00636_),
    .A1(net59),
    .A2(_04116_));
 sg13g2_nand2_1 _09890_ (.Y(_04118_),
    .A(_03828_),
    .B(_03829_));
 sg13g2_xor2_1 _09891_ (.B(_01100_),
    .A(net296),
    .X(_04119_));
 sg13g2_xnor2_1 _09892_ (.Y(_04120_),
    .A(_04118_),
    .B(_04119_));
 sg13g2_xor2_1 _09893_ (.B(_04048_),
    .A(_02613_),
    .X(_04121_));
 sg13g2_nor2_1 _09894_ (.A(net250),
    .B(_04121_),
    .Y(_04122_));
 sg13g2_a221oi_1 _09895_ (.B2(_03877_),
    .C1(_04122_),
    .B1(_04120_),
    .A1(_01355_),
    .Y(_04123_),
    .A2(net72));
 sg13g2_a21oi_1 _09896_ (.A1(_01698_),
    .A2(net48),
    .Y(_04124_),
    .B1(_04123_));
 sg13g2_a22oi_1 _09897_ (.Y(_04125_),
    .B1(net49),
    .B2(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .A2(net164),
    .A1(\i_tinyqv.mem.q_ctrl.addr[1] ));
 sg13g2_o21ai_1 _09898_ (.B1(_04125_),
    .Y(_00637_),
    .A1(net59),
    .A2(_04124_));
 sg13g2_o21ai_1 _09899_ (.B1(_04118_),
    .Y(_04126_),
    .A1(net296),
    .A2(_01100_));
 sg13g2_nand2_1 _09900_ (.Y(_04127_),
    .A(_04126_),
    .B(_03838_));
 sg13g2_xor2_1 _09901_ (.B(net256),
    .A(net260),
    .X(_04128_));
 sg13g2_xnor2_1 _09902_ (.Y(_04129_),
    .A(_04127_),
    .B(_04128_));
 sg13g2_or2_1 _09903_ (.X(_04130_),
    .B(_03856_),
    .A(_02877_));
 sg13g2_xnor2_1 _09904_ (.Y(_04131_),
    .A(net260),
    .B(_04130_));
 sg13g2_nor2_1 _09905_ (.A(net294),
    .B(_04131_),
    .Y(_04132_));
 sg13g2_a21oi_1 _09906_ (.A1(net250),
    .A2(_04129_),
    .Y(_04133_),
    .B1(_04132_));
 sg13g2_mux2_1 _09907_ (.A0(\addr[6] ),
    .A1(_04133_),
    .S(_03864_),
    .X(_04134_));
 sg13g2_and2_1 _09908_ (.A(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .B(_03817_),
    .X(_04135_));
 sg13g2_a221oi_1 _09909_ (.B2(_03797_),
    .C1(_04135_),
    .B1(_04134_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[6] ),
    .Y(_04136_),
    .A2(_03819_));
 sg13g2_inv_1 _09910_ (.Y(_00638_),
    .A(_04136_));
 sg13g2_a21o_1 _09911_ (.A2(_04127_),
    .A1(net260),
    .B1(net256),
    .X(_04137_));
 sg13g2_o21ai_1 _09912_ (.B1(_04137_),
    .Y(_04138_),
    .A1(net260),
    .A2(_04127_));
 sg13g2_xor2_1 _09913_ (.B(_00960_),
    .A(net261),
    .X(_04139_));
 sg13g2_xnor2_1 _09914_ (.Y(_04140_),
    .A(_04138_),
    .B(_04139_));
 sg13g2_xnor2_1 _09915_ (.Y(_04141_),
    .A(_02611_),
    .B(_03878_));
 sg13g2_nor2_1 _09916_ (.A(net249),
    .B(_04141_),
    .Y(_04142_));
 sg13g2_a21oi_1 _09917_ (.A1(net248),
    .A2(_04140_),
    .Y(_04143_),
    .B1(_04142_));
 sg13g2_nor2_1 _09918_ (.A(net47),
    .B(_04143_),
    .Y(_04144_));
 sg13g2_a21oi_1 _09919_ (.A1(\addr[7] ),
    .A2(net48),
    .Y(_04145_),
    .B1(_04144_));
 sg13g2_a22oi_1 _09920_ (.Y(_04146_),
    .B1(net49),
    .B2(\i_tinyqv.mem.q_ctrl.addr[7] ),
    .A2(net164),
    .A1(\i_tinyqv.mem.q_ctrl.addr[3] ));
 sg13g2_o21ai_1 _09921_ (.B1(_04146_),
    .Y(_00639_),
    .A1(net59),
    .A2(_04145_));
 sg13g2_nor3_2 _09922_ (.A(_03845_),
    .B(_03836_),
    .C(_03842_),
    .Y(_04147_));
 sg13g2_xnor2_1 _09923_ (.Y(_04148_),
    .A(_01110_),
    .B(net259));
 sg13g2_xnor2_1 _09924_ (.Y(_04149_),
    .A(_04147_),
    .B(_04148_));
 sg13g2_xnor2_1 _09925_ (.Y(_04150_),
    .A(_02622_),
    .B(_03857_));
 sg13g2_nor2_1 _09926_ (.A(_03821_),
    .B(_04150_),
    .Y(_04151_));
 sg13g2_a221oi_1 _09927_ (.B2(net248),
    .C1(_04151_),
    .B1(_04149_),
    .A1(_01355_),
    .Y(_04152_),
    .A2(net72));
 sg13g2_a21oi_1 _09928_ (.A1(\addr[8] ),
    .A2(_03896_),
    .Y(_04153_),
    .B1(_04152_));
 sg13g2_a22oi_1 _09929_ (.Y(_04154_),
    .B1(net49),
    .B2(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .A2(_03867_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[4] ));
 sg13g2_o21ai_1 _09930_ (.B1(_04154_),
    .Y(_00640_),
    .A1(_03927_),
    .A2(_04153_));
 sg13g2_nor2_1 _09931_ (.A(_02622_),
    .B(_04147_),
    .Y(_04155_));
 sg13g2_nand2_1 _09932_ (.Y(_04156_),
    .A(_02622_),
    .B(_04147_));
 sg13g2_o21ai_1 _09933_ (.B1(_04156_),
    .Y(_04157_),
    .A1(_01110_),
    .A2(_04155_));
 sg13g2_xor2_1 _09934_ (.B(_01065_),
    .A(_01101_),
    .X(_04158_));
 sg13g2_xnor2_1 _09935_ (.Y(_04159_),
    .A(_04157_),
    .B(_04158_));
 sg13g2_nand3_1 _09936_ (.B(net259),
    .C(_03878_),
    .A(net261),
    .Y(_04160_));
 sg13g2_xnor2_1 _09937_ (.Y(_04161_),
    .A(_01066_),
    .B(_04160_));
 sg13g2_nor2_1 _09938_ (.A(_03876_),
    .B(_04161_),
    .Y(_04162_));
 sg13g2_a21oi_1 _09939_ (.A1(_03897_),
    .A2(_04159_),
    .Y(_04163_),
    .B1(_04162_));
 sg13g2_nor2_1 _09940_ (.A(_03930_),
    .B(_04163_),
    .Y(_04164_));
 sg13g2_a21oi_1 _09941_ (.A1(\addr[9] ),
    .A2(_03896_),
    .Y(_04165_),
    .B1(_04164_));
 sg13g2_mux2_1 _09942_ (.A0(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .S(_03813_),
    .X(_04166_));
 sg13g2_nand2_1 _09943_ (.Y(_04167_),
    .A(net62),
    .B(_04166_));
 sg13g2_o21ai_1 _09944_ (.B1(_04167_),
    .Y(_00641_),
    .A1(net59),
    .A2(_04165_));
 sg13g2_buf_1 _09945_ (.A(\i_tinyqv.mem.q_ctrl.is_writing ),
    .X(_04168_));
 sg13g2_buf_1 _09946_ (.A(_04168_),
    .X(_04169_));
 sg13g2_buf_2 _09947_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .X(_04170_));
 sg13g2_nor2_1 _09948_ (.A(net275),
    .B(net312),
    .Y(_04171_));
 sg13g2_nand2_1 _09949_ (.Y(_04172_),
    .A(_04170_),
    .B(_04171_));
 sg13g2_buf_1 _09950_ (.A(_04172_),
    .X(_04173_));
 sg13g2_buf_1 _09951_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .X(_04174_));
 sg13g2_nor3_2 _09952_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .B(_04174_),
    .C(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .Y(_04175_));
 sg13g2_inv_2 _09953_ (.Y(_04176_),
    .A(net312));
 sg13g2_inv_2 _09954_ (.Y(_04177_),
    .A(_04170_));
 sg13g2_nor2_1 _09955_ (.A(_04176_),
    .B(_04177_),
    .Y(_04178_));
 sg13g2_nand2_2 _09956_ (.Y(_04179_),
    .A(net275),
    .B(_04178_));
 sg13g2_inv_1 _09957_ (.Y(_04180_),
    .A(_04179_));
 sg13g2_o21ai_1 _09958_ (.B1(_03808_),
    .Y(_04181_),
    .A1(_04175_),
    .A2(_04180_));
 sg13g2_nand2_1 _09959_ (.Y(_04182_),
    .A(net193),
    .B(_04181_));
 sg13g2_buf_1 _09960_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .X(_04183_));
 sg13g2_buf_2 _09961_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ),
    .X(_04184_));
 sg13g2_nand2_1 _09962_ (.Y(_04185_),
    .A(net312),
    .B(_04170_));
 sg13g2_nor3_1 _09963_ (.A(_04183_),
    .B(_04184_),
    .C(_04185_),
    .Y(_04186_));
 sg13g2_buf_2 _09964_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .X(_04187_));
 sg13g2_a21oi_1 _09965_ (.A1(net275),
    .A2(_04187_),
    .Y(_04188_),
    .B1(_04168_));
 sg13g2_a22oi_1 _09966_ (.Y(_04189_),
    .B1(_04186_),
    .B2(_04188_),
    .A2(_04182_),
    .A1(net247));
 sg13g2_buf_2 _09967_ (.A(_04189_),
    .X(_04190_));
 sg13g2_buf_1 _09968_ (.A(_04190_),
    .X(_04191_));
 sg13g2_inv_2 _09969_ (.Y(_04192_),
    .A(_04168_));
 sg13g2_nand3_1 _09970_ (.B(_04187_),
    .C(_04186_),
    .A(_01648_),
    .Y(_04193_));
 sg13g2_buf_1 _09971_ (.A(_04193_),
    .X(_04194_));
 sg13g2_mux2_1 _09972_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .S(_04194_),
    .X(_04195_));
 sg13g2_nor3_1 _09973_ (.A(_04183_),
    .B(_04187_),
    .C(_04184_),
    .Y(_04196_));
 sg13g2_inv_1 _09974_ (.Y(_04197_),
    .A(_04196_));
 sg13g2_nor2_2 _09975_ (.A(_04179_),
    .B(_04197_),
    .Y(_04198_));
 sg13g2_mux2_1 _09976_ (.A0(_04195_),
    .A1(net8),
    .S(_04198_),
    .X(_04199_));
 sg13g2_xnor2_1 _09977_ (.Y(_04200_),
    .A(_01337_),
    .B(_01296_));
 sg13g2_buf_4 _09978_ (.X(_04201_),
    .A(_04200_));
 sg13g2_nand2_1 _09979_ (.Y(_04202_),
    .A(_01337_),
    .B(_01296_));
 sg13g2_xor2_1 _09980_ (.B(_04202_),
    .A(_01298_),
    .X(_04203_));
 sg13g2_buf_4 _09981_ (.X(_04204_),
    .A(_04203_));
 sg13g2_mux4_1 _09982_ (.S0(_04201_),
    .A0(\data_to_write[24] ),
    .A1(\data_to_write[16] ),
    .A2(\data_to_write[8] ),
    .A3(net309),
    .S1(_04204_),
    .X(_04205_));
 sg13g2_inv_1 _09983_ (.Y(_04206_),
    .A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ));
 sg13g2_inv_1 _09984_ (.Y(_04207_),
    .A(_04174_));
 sg13g2_inv_1 _09985_ (.Y(_04208_),
    .A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ));
 sg13g2_nand3_1 _09986_ (.B(_04207_),
    .C(_04208_),
    .A(_04206_),
    .Y(_04209_));
 sg13g2_buf_1 _09987_ (.A(_04209_),
    .X(_04210_));
 sg13g2_nand2_2 _09988_ (.Y(_04211_),
    .A(net193),
    .B(_04210_));
 sg13g2_mux2_1 _09989_ (.A0(net8),
    .A1(_04205_),
    .S(_04211_),
    .X(_04212_));
 sg13g2_and2_1 _09990_ (.A(net247),
    .B(_04212_),
    .X(_04213_));
 sg13g2_a21oi_1 _09991_ (.A1(_04192_),
    .A2(_04199_),
    .Y(_04214_),
    .B1(_04213_));
 sg13g2_nand2_1 _09992_ (.Y(_04215_),
    .A(_02523_),
    .B(net119));
 sg13g2_o21ai_1 _09993_ (.B1(_04215_),
    .Y(_00642_),
    .A1(_04191_),
    .A2(_04214_));
 sg13g2_mux2_1 _09994_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .S(_04194_),
    .X(_04216_));
 sg13g2_mux2_1 _09995_ (.A0(_04216_),
    .A1(net9),
    .S(_04198_),
    .X(_04217_));
 sg13g2_mux4_1 _09996_ (.S0(_04201_),
    .A0(\data_to_write[25] ),
    .A1(\data_to_write[17] ),
    .A2(\data_to_write[9] ),
    .A3(net308),
    .S1(_04204_),
    .X(_04218_));
 sg13g2_mux2_1 _09997_ (.A0(net9),
    .A1(_04218_),
    .S(_04211_),
    .X(_04219_));
 sg13g2_and2_1 _09998_ (.A(net247),
    .B(_04219_),
    .X(_04220_));
 sg13g2_a21oi_1 _09999_ (.A1(_04192_),
    .A2(_04217_),
    .Y(_04221_),
    .B1(_04220_));
 sg13g2_nand2_1 _10000_ (.Y(_04222_),
    .A(_02788_),
    .B(net119));
 sg13g2_o21ai_1 _10001_ (.B1(_04222_),
    .Y(_00643_),
    .A1(net119),
    .A2(_04221_));
 sg13g2_mux2_1 _10002_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .S(_04194_),
    .X(_04223_));
 sg13g2_mux2_1 _10003_ (.A0(_04223_),
    .A1(net10),
    .S(_04198_),
    .X(_04224_));
 sg13g2_mux4_1 _10004_ (.S0(_04201_),
    .A0(\data_to_write[26] ),
    .A1(\data_to_write[18] ),
    .A2(\data_to_write[10] ),
    .A3(net307),
    .S1(_04204_),
    .X(_04225_));
 sg13g2_mux2_1 _10005_ (.A0(net10),
    .A1(_04225_),
    .S(_04211_),
    .X(_04226_));
 sg13g2_and2_1 _10006_ (.A(net247),
    .B(_04226_),
    .X(_04227_));
 sg13g2_a21oi_1 _10007_ (.A1(_04192_),
    .A2(_04224_),
    .Y(_04228_),
    .B1(_04227_));
 sg13g2_nand2_1 _10008_ (.Y(_04229_),
    .A(_02904_),
    .B(_04190_));
 sg13g2_o21ai_1 _10009_ (.B1(_04229_),
    .Y(_00644_),
    .A1(net119),
    .A2(_04228_));
 sg13g2_mux2_1 _10010_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .S(_04194_),
    .X(_04230_));
 sg13g2_mux2_1 _10011_ (.A0(_04230_),
    .A1(net11),
    .S(_04198_),
    .X(_04231_));
 sg13g2_mux4_1 _10012_ (.S0(_04201_),
    .A0(\data_to_write[27] ),
    .A1(\data_to_write[19] ),
    .A2(\data_to_write[11] ),
    .A3(_01724_),
    .S1(_04204_),
    .X(_04232_));
 sg13g2_mux2_1 _10013_ (.A0(net11),
    .A1(_04232_),
    .S(_04211_),
    .X(_04233_));
 sg13g2_and2_1 _10014_ (.A(net247),
    .B(_04233_),
    .X(_04234_));
 sg13g2_a21oi_1 _10015_ (.A1(_04192_),
    .A2(_04231_),
    .Y(_04235_),
    .B1(_04234_));
 sg13g2_nand2_1 _10016_ (.Y(_04236_),
    .A(_02999_),
    .B(_04190_));
 sg13g2_o21ai_1 _10017_ (.B1(_04236_),
    .Y(_00645_),
    .A1(net119),
    .A2(_04235_));
 sg13g2_mux4_1 _10018_ (.S0(_04201_),
    .A0(\data_to_write[28] ),
    .A1(\data_to_write[20] ),
    .A2(\data_to_write[12] ),
    .A3(net306),
    .S1(_04204_),
    .X(_04237_));
 sg13g2_a21oi_1 _10019_ (.A1(net193),
    .A2(_04210_),
    .Y(_04238_),
    .B1(_04192_));
 sg13g2_buf_2 _10020_ (.A(_04238_),
    .X(_04239_));
 sg13g2_nor2b_1 _10021_ (.A(_04239_),
    .B_N(_02523_),
    .Y(_04240_));
 sg13g2_a21oi_1 _10022_ (.A1(_04237_),
    .A2(_04239_),
    .Y(_04241_),
    .B1(_04240_));
 sg13g2_nand2_1 _10023_ (.Y(_04242_),
    .A(_02576_),
    .B(_04190_));
 sg13g2_o21ai_1 _10024_ (.B1(_04242_),
    .Y(_00646_),
    .A1(net119),
    .A2(_04241_));
 sg13g2_mux4_1 _10025_ (.S0(_04201_),
    .A0(\data_to_write[29] ),
    .A1(\data_to_write[21] ),
    .A2(\data_to_write[13] ),
    .A3(net305),
    .S1(_04204_),
    .X(_04243_));
 sg13g2_nor2b_1 _10026_ (.A(_04239_),
    .B_N(_02788_),
    .Y(_04244_));
 sg13g2_a21oi_1 _10027_ (.A1(_04239_),
    .A2(_04243_),
    .Y(_04245_),
    .B1(_04244_));
 sg13g2_nand2_1 _10028_ (.Y(_04246_),
    .A(_02769_),
    .B(_04190_));
 sg13g2_o21ai_1 _10029_ (.B1(_04246_),
    .Y(_00647_),
    .A1(net119),
    .A2(_04245_));
 sg13g2_mux4_1 _10030_ (.S0(_04201_),
    .A0(\data_to_write[30] ),
    .A1(\data_to_write[22] ),
    .A2(\data_to_write[14] ),
    .A3(net304),
    .S1(_04204_),
    .X(_04247_));
 sg13g2_mux2_1 _10031_ (.A0(_02904_),
    .A1(_04247_),
    .S(_04239_),
    .X(_04248_));
 sg13g2_nor2_1 _10032_ (.A(_04190_),
    .B(_04248_),
    .Y(_04249_));
 sg13g2_a21oi_1 _10033_ (.A1(_02898_),
    .A2(_04191_),
    .Y(_00648_),
    .B1(_04249_));
 sg13g2_mux4_1 _10034_ (.S0(_04201_),
    .A0(\data_to_write[31] ),
    .A1(\data_to_write[23] ),
    .A2(\data_to_write[15] ),
    .A3(_01737_),
    .S1(_04204_),
    .X(_04250_));
 sg13g2_nor2b_1 _10035_ (.A(_04239_),
    .B_N(_02999_),
    .Y(_04251_));
 sg13g2_a21oi_1 _10036_ (.A1(_04239_),
    .A2(_04250_),
    .Y(_04252_),
    .B1(_04251_));
 sg13g2_nand2_1 _10037_ (.Y(_04253_),
    .A(_02961_),
    .B(_04190_));
 sg13g2_o21ai_1 _10038_ (.B1(_04253_),
    .Y(_00649_),
    .A1(net119),
    .A2(_04252_));
 sg13g2_or2_1 _10039_ (.X(_04254_),
    .B(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .A(_03062_));
 sg13g2_inv_1 _10040_ (.Y(_04255_),
    .A(_03808_));
 sg13g2_nor2_1 _10041_ (.A(_01641_),
    .B(_01644_),
    .Y(_04256_));
 sg13g2_nand3_1 _10042_ (.B(_01596_),
    .C(_01660_),
    .A(_01659_),
    .Y(_04257_));
 sg13g2_a221oi_1 _10043_ (.B2(_04257_),
    .C1(_01655_),
    .B1(_04256_),
    .A1(_04168_),
    .Y(_04258_),
    .A2(_04255_));
 sg13g2_or3_1 _10044_ (.A(_01653_),
    .B(_04254_),
    .C(_04258_),
    .X(_04259_));
 sg13g2_buf_2 _10045_ (.A(_04259_),
    .X(_04260_));
 sg13g2_buf_1 _10046_ (.A(\i_tinyqv.mem.data_stall ),
    .X(_04261_));
 sg13g2_nor4_2 _10047_ (.A(_04187_),
    .B(_04184_),
    .C(_04261_),
    .Y(_04262_),
    .D(_01634_));
 sg13g2_inv_1 _10048_ (.Y(_04263_),
    .A(_04262_));
 sg13g2_nor3_1 _10049_ (.A(net247),
    .B(_04173_),
    .C(_04263_),
    .Y(_04264_));
 sg13g2_or2_1 _10050_ (.X(_04265_),
    .B(_04196_),
    .A(_00167_));
 sg13g2_buf_1 _10051_ (.A(_00164_),
    .X(_04266_));
 sg13g2_o21ai_1 _10052_ (.B1(_04178_),
    .Y(_04267_),
    .A1(_01648_),
    .A2(_04266_));
 sg13g2_mux2_1 _10053_ (.A0(_04196_),
    .A1(_03808_),
    .S(_04267_),
    .X(_04268_));
 sg13g2_buf_2 _10054_ (.A(_04268_),
    .X(_04269_));
 sg13g2_buf_1 _10055_ (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ),
    .X(_04270_));
 sg13g2_nand3_1 _10056_ (.B(_04270_),
    .C(_04178_),
    .A(_01648_),
    .Y(_04271_));
 sg13g2_buf_1 _10057_ (.A(_04271_),
    .X(_04272_));
 sg13g2_nand2_1 _10058_ (.Y(_04273_),
    .A(_04210_),
    .B(_04272_));
 sg13g2_and2_1 _10059_ (.A(_04269_),
    .B(_04273_),
    .X(_04274_));
 sg13g2_buf_1 _10060_ (.A(_04274_),
    .X(_04275_));
 sg13g2_and2_1 _10061_ (.A(_04170_),
    .B(_04275_),
    .X(_04276_));
 sg13g2_buf_1 _10062_ (.A(_01648_),
    .X(_04277_));
 sg13g2_nor2b_1 _10063_ (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .B_N(_04275_),
    .Y(_04278_));
 sg13g2_nor2_1 _10064_ (.A(net312),
    .B(_04177_),
    .Y(_04279_));
 sg13g2_o21ai_1 _10065_ (.B1(_04279_),
    .Y(_04280_),
    .A1(_04277_),
    .A2(_04278_));
 sg13g2_o21ai_1 _10066_ (.B1(_04280_),
    .Y(_04281_),
    .A1(_04265_),
    .A2(_04276_));
 sg13g2_o21ai_1 _10067_ (.B1(_04281_),
    .Y(_04282_),
    .A1(net193),
    .A2(_04262_));
 sg13g2_nor3_1 _10068_ (.A(_04261_),
    .B(_01634_),
    .C(_04185_),
    .Y(_04283_));
 sg13g2_nor2_1 _10069_ (.A(_04281_),
    .B(_04283_),
    .Y(_04284_));
 sg13g2_a221oi_1 _10070_ (.B2(_04282_),
    .C1(_04284_),
    .B1(_04265_),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .Y(_04285_),
    .A2(_04264_));
 sg13g2_nand2_1 _10071_ (.Y(_04286_),
    .A(_04183_),
    .B(_04260_));
 sg13g2_o21ai_1 _10072_ (.B1(_04286_),
    .Y(_00664_),
    .A1(_04260_),
    .A2(_04285_));
 sg13g2_buf_1 _10073_ (.A(_01647_),
    .X(_04287_));
 sg13g2_nor2_1 _10074_ (.A(_04261_),
    .B(_01634_),
    .Y(_04288_));
 sg13g2_nand2b_1 _10075_ (.Y(_04289_),
    .B(_04276_),
    .A_N(_04171_));
 sg13g2_a21oi_2 _10076_ (.B1(_04289_),
    .Y(_04290_),
    .A2(_04288_),
    .A1(net245));
 sg13g2_nor2_1 _10077_ (.A(_04183_),
    .B(_04187_),
    .Y(_04291_));
 sg13g2_nand2_1 _10078_ (.Y(_04292_),
    .A(_04184_),
    .B(_04291_));
 sg13g2_nand2_1 _10079_ (.Y(_04293_),
    .A(_04183_),
    .B(_04187_));
 sg13g2_a21oi_1 _10080_ (.A1(_04292_),
    .A2(_04293_),
    .Y(_04294_),
    .B1(_04290_));
 sg13g2_a221oi_1 _10081_ (.B2(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .C1(_04294_),
    .B1(_04290_),
    .A1(_04270_),
    .Y(_04295_),
    .A2(_04264_));
 sg13g2_nand2_1 _10082_ (.Y(_04296_),
    .A(_04187_),
    .B(_04260_));
 sg13g2_o21ai_1 _10083_ (.B1(_04296_),
    .Y(_00665_),
    .A1(_04260_),
    .A2(_04295_));
 sg13g2_nand2_1 _10084_ (.Y(_04297_),
    .A(_04270_),
    .B(_04290_));
 sg13g2_nor2_1 _10085_ (.A(_04290_),
    .B(_04291_),
    .Y(_04298_));
 sg13g2_o21ai_1 _10086_ (.B1(_04184_),
    .Y(_04299_),
    .A1(_04260_),
    .A2(_04298_));
 sg13g2_o21ai_1 _10087_ (.B1(_04299_),
    .Y(_00666_),
    .A1(_04260_),
    .A2(_04297_));
 sg13g2_nor2_1 _10088_ (.A(_04187_),
    .B(_04184_),
    .Y(_04300_));
 sg13g2_nand2_1 _10089_ (.Y(_04301_),
    .A(_04266_),
    .B(_00167_));
 sg13g2_nor3_1 _10090_ (.A(net193),
    .B(_04300_),
    .C(_04301_),
    .Y(_04302_));
 sg13g2_buf_4 _10091_ (.X(_04303_),
    .A(_04302_));
 sg13g2_mux2_1 _10092_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .A1(net8),
    .S(_04303_),
    .X(_00670_));
 sg13g2_mux2_1 _10093_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .A1(net9),
    .S(_04303_),
    .X(_00671_));
 sg13g2_mux2_1 _10094_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .A1(net10),
    .S(_04303_),
    .X(_00672_));
 sg13g2_mux2_1 _10095_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .A1(net11),
    .S(_04303_),
    .X(_00673_));
 sg13g2_mux2_1 _10096_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .S(_04303_),
    .X(_00674_));
 sg13g2_mux2_1 _10097_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .S(_04303_),
    .X(_00675_));
 sg13g2_mux2_1 _10098_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .S(_04303_),
    .X(_00676_));
 sg13g2_mux2_1 _10099_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .S(_04303_),
    .X(_00677_));
 sg13g2_nor2_1 _10100_ (.A(net322),
    .B(net318),
    .Y(_04304_));
 sg13g2_nand2_1 _10101_ (.Y(_04305_),
    .A(net319),
    .B(_04304_));
 sg13g2_buf_1 _10102_ (.A(_04305_),
    .X(_04306_));
 sg13g2_mux2_1 _10103_ (.A0(_02523_),
    .A1(\i_tinyqv.cpu.instr_data_in[0] ),
    .S(net215),
    .X(_00681_));
 sg13g2_nor2b_1 _10104_ (.A(net318),
    .B_N(net322),
    .Y(_04307_));
 sg13g2_buf_1 _10105_ (.A(_01303_),
    .X(_04308_));
 sg13g2_nor2b_1 _10106_ (.A(_04308_),
    .B_N(net319),
    .Y(_04309_));
 sg13g2_o21ai_1 _10107_ (.B1(_04309_),
    .Y(_04310_),
    .A1(_01339_),
    .A2(_04307_));
 sg13g2_buf_2 _10108_ (.A(_04310_),
    .X(_04311_));
 sg13g2_nand2_1 _10109_ (.Y(_04312_),
    .A(\i_tinyqv.mem.qspi_data_buf[10] ),
    .B(net199));
 sg13g2_o21ai_1 _10110_ (.B1(_04312_),
    .Y(_00682_),
    .A1(_03602_),
    .A2(_04311_));
 sg13g2_nand2_1 _10111_ (.Y(_04313_),
    .A(\i_tinyqv.mem.qspi_data_buf[11] ),
    .B(net199));
 sg13g2_o21ai_1 _10112_ (.B1(_04313_),
    .Y(_00683_),
    .A1(_03605_),
    .A2(_04311_));
 sg13g2_nand2_1 _10113_ (.Y(_04314_),
    .A(\i_tinyqv.mem.qspi_data_buf[12] ),
    .B(net199));
 sg13g2_o21ai_1 _10114_ (.B1(_04314_),
    .Y(_00684_),
    .A1(_03607_),
    .A2(_04311_));
 sg13g2_nand2_1 _10115_ (.Y(_04315_),
    .A(\i_tinyqv.mem.qspi_data_buf[13] ),
    .B(net199));
 sg13g2_o21ai_1 _10116_ (.B1(_04315_),
    .Y(_00685_),
    .A1(_03609_),
    .A2(_04311_));
 sg13g2_nand2_1 _10117_ (.Y(_04316_),
    .A(\i_tinyqv.mem.qspi_data_buf[14] ),
    .B(net199));
 sg13g2_o21ai_1 _10118_ (.B1(_04316_),
    .Y(_00686_),
    .A1(_03611_),
    .A2(_04311_));
 sg13g2_nand2_1 _10119_ (.Y(_04317_),
    .A(\i_tinyqv.mem.qspi_data_buf[15] ),
    .B(net199));
 sg13g2_o21ai_1 _10120_ (.B1(_04317_),
    .Y(_00687_),
    .A1(_03613_),
    .A2(_04311_));
 sg13g2_nand3b_1 _10121_ (.B(net322),
    .C(net319),
    .Y(_04318_),
    .A_N(net318));
 sg13g2_buf_2 _10122_ (.A(_04318_),
    .X(_04319_));
 sg13g2_buf_1 _10123_ (.A(_04319_),
    .X(_04320_));
 sg13g2_nand2_1 _10124_ (.Y(_04321_),
    .A(\i_tinyqv.mem.data_from_read[16] ),
    .B(net214));
 sg13g2_o21ai_1 _10125_ (.B1(_04321_),
    .Y(_00688_),
    .A1(_03617_),
    .A2(net214));
 sg13g2_nand2_1 _10126_ (.Y(_04322_),
    .A(\i_tinyqv.mem.data_from_read[17] ),
    .B(net214));
 sg13g2_o21ai_1 _10127_ (.B1(_04322_),
    .Y(_00689_),
    .A1(_03619_),
    .A2(net214));
 sg13g2_nand2_1 _10128_ (.Y(_04323_),
    .A(\i_tinyqv.mem.data_from_read[18] ),
    .B(_04319_));
 sg13g2_o21ai_1 _10129_ (.B1(_04323_),
    .Y(_00690_),
    .A1(_03602_),
    .A2(net214));
 sg13g2_nand2_1 _10130_ (.Y(_04324_),
    .A(\i_tinyqv.mem.data_from_read[19] ),
    .B(_04319_));
 sg13g2_o21ai_1 _10131_ (.B1(_04324_),
    .Y(_00691_),
    .A1(_03605_),
    .A2(_04320_));
 sg13g2_mux2_1 _10132_ (.A0(_02788_),
    .A1(\i_tinyqv.cpu.instr_data_in[1] ),
    .S(_04306_),
    .X(_00692_));
 sg13g2_nand2_1 _10133_ (.Y(_04325_),
    .A(\i_tinyqv.mem.data_from_read[20] ),
    .B(_04319_));
 sg13g2_o21ai_1 _10134_ (.B1(_04325_),
    .Y(_00693_),
    .A1(_03607_),
    .A2(net214));
 sg13g2_nand2_1 _10135_ (.Y(_04326_),
    .A(\i_tinyqv.mem.data_from_read[21] ),
    .B(_04319_));
 sg13g2_o21ai_1 _10136_ (.B1(_04326_),
    .Y(_00694_),
    .A1(_03609_),
    .A2(net214));
 sg13g2_nand2_1 _10137_ (.Y(_04327_),
    .A(\i_tinyqv.mem.data_from_read[22] ),
    .B(_04319_));
 sg13g2_o21ai_1 _10138_ (.B1(_04327_),
    .Y(_00695_),
    .A1(_03611_),
    .A2(net214));
 sg13g2_nand2_1 _10139_ (.Y(_04328_),
    .A(\i_tinyqv.mem.data_from_read[23] ),
    .B(_04319_));
 sg13g2_o21ai_1 _10140_ (.B1(_04328_),
    .Y(_00696_),
    .A1(_03613_),
    .A2(_04320_));
 sg13g2_and2_1 _10141_ (.A(net322),
    .B(net318),
    .X(_04329_));
 sg13g2_nand2_1 _10142_ (.Y(_04330_),
    .A(net319),
    .B(_04329_));
 sg13g2_buf_1 _10143_ (.A(_04330_),
    .X(_04331_));
 sg13g2_buf_1 _10144_ (.A(_04331_),
    .X(_04332_));
 sg13g2_nor3_1 _10145_ (.A(net244),
    .B(_03617_),
    .C(net192),
    .Y(_04333_));
 sg13g2_a21o_1 _10146_ (.A2(net192),
    .A1(\i_tinyqv.mem.qspi_data_buf[24] ),
    .B1(_04333_),
    .X(_00697_));
 sg13g2_nor3_1 _10147_ (.A(net244),
    .B(_03619_),
    .C(net192),
    .Y(_04334_));
 sg13g2_a21o_1 _10148_ (.A2(net192),
    .A1(\i_tinyqv.mem.qspi_data_buf[25] ),
    .B1(_04334_),
    .X(_00698_));
 sg13g2_nor3_1 _10149_ (.A(net244),
    .B(_03602_),
    .C(_04331_),
    .Y(_04335_));
 sg13g2_a21o_1 _10150_ (.A2(net192),
    .A1(\i_tinyqv.mem.qspi_data_buf[26] ),
    .B1(_04335_),
    .X(_00699_));
 sg13g2_nor3_1 _10151_ (.A(net244),
    .B(_03605_),
    .C(_04331_),
    .Y(_04336_));
 sg13g2_a21o_1 _10152_ (.A2(_04332_),
    .A1(\i_tinyqv.mem.qspi_data_buf[27] ),
    .B1(_04336_),
    .X(_00700_));
 sg13g2_nor3_1 _10153_ (.A(net244),
    .B(_03607_),
    .C(_04331_),
    .Y(_04337_));
 sg13g2_a21o_1 _10154_ (.A2(_04332_),
    .A1(\i_tinyqv.mem.qspi_data_buf[28] ),
    .B1(_04337_),
    .X(_00701_));
 sg13g2_nor3_1 _10155_ (.A(net244),
    .B(_03609_),
    .C(_04331_),
    .Y(_04338_));
 sg13g2_a21o_1 _10156_ (.A2(net192),
    .A1(\i_tinyqv.mem.qspi_data_buf[29] ),
    .B1(_04338_),
    .X(_00702_));
 sg13g2_mux2_1 _10157_ (.A0(_02904_),
    .A1(_02905_),
    .S(net215),
    .X(_00703_));
 sg13g2_nor3_1 _10158_ (.A(net244),
    .B(_03611_),
    .C(_04331_),
    .Y(_04339_));
 sg13g2_a21o_1 _10159_ (.A2(net192),
    .A1(\i_tinyqv.mem.qspi_data_buf[30] ),
    .B1(_04339_),
    .X(_00704_));
 sg13g2_nor3_1 _10160_ (.A(net244),
    .B(_03613_),
    .C(_04331_),
    .Y(_04340_));
 sg13g2_a21o_1 _10161_ (.A2(net192),
    .A1(\i_tinyqv.mem.qspi_data_buf[31] ),
    .B1(_04340_),
    .X(_00705_));
 sg13g2_mux2_1 _10162_ (.A0(_02999_),
    .A1(_03012_),
    .S(net215),
    .X(_00706_));
 sg13g2_mux2_1 _10163_ (.A0(_02576_),
    .A1(_02577_),
    .S(net215),
    .X(_00707_));
 sg13g2_mux2_1 _10164_ (.A0(_02769_),
    .A1(_02773_),
    .S(net215),
    .X(_00708_));
 sg13g2_nand2_1 _10165_ (.Y(_04341_),
    .A(_02899_),
    .B(net215));
 sg13g2_o21ai_1 _10166_ (.B1(_04341_),
    .Y(_00709_),
    .A1(_02898_),
    .A2(net215));
 sg13g2_mux2_1 _10167_ (.A0(_02961_),
    .A1(_02962_),
    .S(net215),
    .X(_00710_));
 sg13g2_nand2_1 _10168_ (.Y(_04342_),
    .A(\i_tinyqv.mem.qspi_data_buf[8] ),
    .B(net199));
 sg13g2_o21ai_1 _10169_ (.B1(_04342_),
    .Y(_00711_),
    .A1(_03617_),
    .A2(_04311_));
 sg13g2_nand2_1 _10170_ (.Y(_04343_),
    .A(\i_tinyqv.mem.qspi_data_buf[9] ),
    .B(net199));
 sg13g2_o21ai_1 _10171_ (.B1(_04343_),
    .Y(_00712_),
    .A1(_03619_),
    .A2(_04311_));
 sg13g2_buf_1 _10172_ (.A(\i_uart_rx.cycle_counter[5] ),
    .X(_04344_));
 sg13g2_buf_1 _10173_ (.A(\i_uart_rx.cycle_counter[1] ),
    .X(_04345_));
 sg13g2_buf_1 _10174_ (.A(\i_uart_rx.cycle_counter[0] ),
    .X(_04346_));
 sg13g2_and3_1 _10175_ (.X(_04347_),
    .A(_04345_),
    .B(_04346_),
    .C(\i_uart_rx.cycle_counter[3] ));
 sg13g2_buf_1 _10176_ (.A(_04347_),
    .X(_04348_));
 sg13g2_buf_1 _10177_ (.A(\i_uart_rx.cycle_counter[7] ),
    .X(_04349_));
 sg13g2_nor3_1 _10178_ (.A(_04349_),
    .B(\i_uart_rx.cycle_counter[6] ),
    .C(\i_uart_rx.cycle_counter[10] ),
    .Y(_04350_));
 sg13g2_buf_2 _10179_ (.A(\i_uart_rx.cycle_counter[2] ),
    .X(_04351_));
 sg13g2_buf_1 _10180_ (.A(\i_uart_rx.cycle_counter[4] ),
    .X(_04352_));
 sg13g2_inv_1 _10181_ (.Y(_04353_),
    .A(\i_uart_rx.cycle_counter[9] ));
 sg13g2_nor4_1 _10182_ (.A(_04351_),
    .B(_04352_),
    .C(_04353_),
    .D(\i_uart_rx.cycle_counter[8] ),
    .Y(_04354_));
 sg13g2_and4_1 _10183_ (.A(_04344_),
    .B(_04348_),
    .C(_04350_),
    .D(_04354_),
    .X(_04355_));
 sg13g2_buf_1 _10184_ (.A(_04355_),
    .X(_04356_));
 sg13g2_nor2_1 _10185_ (.A(net316),
    .B(_01368_),
    .Y(_04357_));
 sg13g2_xnor2_1 _10186_ (.Y(_04358_),
    .A(net315),
    .B(_04357_));
 sg13g2_nand2_1 _10187_ (.Y(_04359_),
    .A(_04356_),
    .B(_04358_));
 sg13g2_buf_4 _10188_ (.X(_04360_),
    .A(_04359_));
 sg13g2_mux2_1 _10189_ (.A0(\i_uart_rx.recieved_data[1] ),
    .A1(\i_uart_rx.recieved_data[0] ),
    .S(_04360_),
    .X(_00731_));
 sg13g2_mux2_1 _10190_ (.A0(\i_uart_rx.recieved_data[2] ),
    .A1(\i_uart_rx.recieved_data[1] ),
    .S(_04360_),
    .X(_00732_));
 sg13g2_mux2_1 _10191_ (.A0(\i_uart_rx.recieved_data[3] ),
    .A1(\i_uart_rx.recieved_data[2] ),
    .S(_04360_),
    .X(_00733_));
 sg13g2_mux2_1 _10192_ (.A0(\i_uart_rx.recieved_data[4] ),
    .A1(\i_uart_rx.recieved_data[3] ),
    .S(_04360_),
    .X(_00734_));
 sg13g2_mux2_1 _10193_ (.A0(\i_uart_rx.recieved_data[5] ),
    .A1(\i_uart_rx.recieved_data[4] ),
    .S(_04360_),
    .X(_00735_));
 sg13g2_mux2_1 _10194_ (.A0(\i_uart_rx.recieved_data[6] ),
    .A1(\i_uart_rx.recieved_data[5] ),
    .S(_04360_),
    .X(_00736_));
 sg13g2_mux2_1 _10195_ (.A0(\i_uart_rx.recieved_data[7] ),
    .A1(\i_uart_rx.recieved_data[6] ),
    .S(_04360_),
    .X(_00737_));
 sg13g2_mux2_1 _10196_ (.A0(\i_uart_rx.bit_sample ),
    .A1(\i_uart_rx.recieved_data[7] ),
    .S(_04360_),
    .X(_00738_));
 sg13g2_nand2_1 _10197_ (.Y(_04361_),
    .A(net179),
    .B(net218));
 sg13g2_buf_1 _10198_ (.A(_04361_),
    .X(_04362_));
 sg13g2_buf_1 _10199_ (.A(_04362_),
    .X(_04363_));
 sg13g2_mux2_1 _10200_ (.A0(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[4] ),
    .S(net139),
    .X(_00387_));
 sg13g2_mux2_1 _10201_ (.A0(\i_tinyqv.cpu.i_core.mepc[10] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[14] ),
    .S(net139),
    .X(_00388_));
 sg13g2_mux2_1 _10202_ (.A0(\i_tinyqv.cpu.i_core.mepc[11] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[15] ),
    .S(net139),
    .X(_00389_));
 sg13g2_mux2_1 _10203_ (.A0(\i_tinyqv.cpu.i_core.mepc[12] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[16] ),
    .S(net139),
    .X(_00390_));
 sg13g2_mux2_1 _10204_ (.A0(\i_tinyqv.cpu.i_core.mepc[13] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[17] ),
    .S(net139),
    .X(_00391_));
 sg13g2_mux2_1 _10205_ (.A0(\i_tinyqv.cpu.i_core.mepc[14] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[18] ),
    .S(_04363_),
    .X(_00392_));
 sg13g2_mux2_1 _10206_ (.A0(\i_tinyqv.cpu.i_core.mepc[15] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[19] ),
    .S(net139),
    .X(_00393_));
 sg13g2_mux2_1 _10207_ (.A0(\i_tinyqv.cpu.i_core.mepc[16] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[20] ),
    .S(net139),
    .X(_00394_));
 sg13g2_mux2_1 _10208_ (.A0(\i_tinyqv.cpu.i_core.mepc[17] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[21] ),
    .S(net139),
    .X(_00395_));
 sg13g2_mux2_1 _10209_ (.A0(\i_tinyqv.cpu.i_core.mepc[18] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[22] ),
    .S(_04363_),
    .X(_00396_));
 sg13g2_buf_1 _10210_ (.A(_04362_),
    .X(_04364_));
 sg13g2_mux2_1 _10211_ (.A0(\i_tinyqv.cpu.i_core.mepc[19] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[23] ),
    .S(net138),
    .X(_00397_));
 sg13g2_mux2_1 _10212_ (.A0(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[5] ),
    .S(net138),
    .X(_00398_));
 sg13g2_nor2_2 _10213_ (.A(_01677_),
    .B(_02369_),
    .Y(_04365_));
 sg13g2_nor2b_1 _10214_ (.A(_02686_),
    .B_N(_04365_),
    .Y(_04366_));
 sg13g2_buf_2 _10215_ (.A(_04366_),
    .X(_04367_));
 sg13g2_nor2_1 _10216_ (.A(\i_tinyqv.cpu.i_core.mepc[0] ),
    .B(_04367_),
    .Y(_04368_));
 sg13g2_a21oi_1 _10217_ (.A1(net158),
    .A2(_04367_),
    .Y(_04369_),
    .B1(_04368_));
 sg13g2_nor3_1 _10218_ (.A(_01177_),
    .B(_01181_),
    .C(net183),
    .Y(_04370_));
 sg13g2_a21oi_1 _10219_ (.A1(net183),
    .A2(_04369_),
    .Y(_04371_),
    .B1(_04370_));
 sg13g2_buf_1 _10220_ (.A(_01541_),
    .X(_04372_));
 sg13g2_nand2_1 _10221_ (.Y(_04373_),
    .A(net243),
    .B(_04362_));
 sg13g2_nand2_1 _10222_ (.Y(_04374_),
    .A(\i_tinyqv.cpu.i_core.mepc[20] ),
    .B(_02685_));
 sg13g2_o21ai_1 _10223_ (.B1(_04374_),
    .Y(_00399_),
    .A1(_04371_),
    .A2(_04373_));
 sg13g2_inv_1 _10224_ (.Y(_04375_),
    .A(_01057_));
 sg13g2_nor2_1 _10225_ (.A(\i_tinyqv.cpu.i_core.mepc[1] ),
    .B(_04367_),
    .Y(_04376_));
 sg13g2_a21oi_1 _10226_ (.A1(_04375_),
    .A2(_04367_),
    .Y(_04377_),
    .B1(_04376_));
 sg13g2_a21oi_1 _10227_ (.A1(_01070_),
    .A2(_01073_),
    .Y(_04378_),
    .B1(net183));
 sg13g2_a21oi_1 _10228_ (.A1(net183),
    .A2(_04377_),
    .Y(_04379_),
    .B1(_04378_));
 sg13g2_nand2_1 _10229_ (.Y(_04380_),
    .A(\i_tinyqv.cpu.i_core.mepc[21] ),
    .B(_02685_));
 sg13g2_o21ai_1 _10230_ (.B1(_04380_),
    .Y(_00400_),
    .A1(_04373_),
    .A2(_04379_));
 sg13g2_nor2_1 _10231_ (.A(\i_tinyqv.cpu.i_core.mepc[2] ),
    .B(_04367_),
    .Y(_04381_));
 sg13g2_and2_1 _10232_ (.A(_01014_),
    .B(_04367_),
    .X(_04382_));
 sg13g2_nor3_1 _10233_ (.A(net186),
    .B(_04381_),
    .C(_04382_),
    .Y(_04383_));
 sg13g2_a21oi_1 _10234_ (.A1(_01033_),
    .A2(net186),
    .Y(_04384_),
    .B1(_04383_));
 sg13g2_nand2_1 _10235_ (.Y(_04385_),
    .A(\i_tinyqv.cpu.i_core.mepc[22] ),
    .B(_02685_));
 sg13g2_o21ai_1 _10236_ (.B1(_04385_),
    .Y(_00401_),
    .A1(_04373_),
    .A2(_04384_));
 sg13g2_nand2_1 _10237_ (.Y(_04386_),
    .A(_01893_),
    .B(_04367_));
 sg13g2_o21ai_1 _10238_ (.B1(_04386_),
    .Y(_04387_),
    .A1(\i_tinyqv.cpu.i_core.mepc[3] ),
    .A2(_04367_));
 sg13g2_nor2_1 _10239_ (.A(_01227_),
    .B(_04387_),
    .Y(_04388_));
 sg13g2_a21oi_1 _10240_ (.A1(_00852_),
    .A2(_01227_),
    .Y(_04389_),
    .B1(_04388_));
 sg13g2_nand2_1 _10241_ (.Y(_04390_),
    .A(\i_tinyqv.cpu.i_core.mepc[23] ),
    .B(_02685_));
 sg13g2_o21ai_1 _10242_ (.B1(_04390_),
    .Y(_00402_),
    .A1(_04373_),
    .A2(_04389_));
 sg13g2_mux2_1 _10243_ (.A0(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[6] ),
    .S(net138),
    .X(_00403_));
 sg13g2_mux2_1 _10244_ (.A0(\i_tinyqv.cpu.i_core.mepc[3] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[7] ),
    .S(net138),
    .X(_00404_));
 sg13g2_mux2_1 _10245_ (.A0(\i_tinyqv.cpu.i_core.mepc[4] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[8] ),
    .S(net138),
    .X(_00405_));
 sg13g2_mux2_1 _10246_ (.A0(\i_tinyqv.cpu.i_core.mepc[5] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[9] ),
    .S(net138),
    .X(_00406_));
 sg13g2_mux2_1 _10247_ (.A0(\i_tinyqv.cpu.i_core.mepc[6] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[10] ),
    .S(net138),
    .X(_00407_));
 sg13g2_mux2_1 _10248_ (.A0(\i_tinyqv.cpu.i_core.mepc[7] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[11] ),
    .S(net138),
    .X(_00408_));
 sg13g2_mux2_1 _10249_ (.A0(\i_tinyqv.cpu.i_core.mepc[8] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[12] ),
    .S(_04364_),
    .X(_00409_));
 sg13g2_mux2_1 _10250_ (.A0(\i_tinyqv.cpu.i_core.mepc[9] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[13] ),
    .S(_04364_),
    .X(_00410_));
 sg13g2_a21oi_1 _10251_ (.A1(net198),
    .A2(_02369_),
    .Y(_04391_),
    .B1(_02367_));
 sg13g2_buf_1 _10252_ (.A(_04391_),
    .X(_04392_));
 sg13g2_buf_1 _10253_ (.A(_04392_),
    .X(_04393_));
 sg13g2_mux2_1 _10254_ (.A0(net302),
    .A1(net269),
    .S(net154),
    .X(_00426_));
 sg13g2_inv_1 _10255_ (.Y(_04394_),
    .A(_02303_));
 sg13g2_buf_1 _10256_ (.A(_04392_),
    .X(_04395_));
 sg13g2_nand2_1 _10257_ (.Y(_04396_),
    .A(_02168_),
    .B(net153));
 sg13g2_o21ai_1 _10258_ (.B1(_04396_),
    .Y(_00427_),
    .A1(_04394_),
    .A2(net154));
 sg13g2_inv_1 _10259_ (.Y(_04397_),
    .A(_02350_));
 sg13g2_nand2_1 _10260_ (.Y(_04398_),
    .A(_02204_),
    .B(net153));
 sg13g2_o21ai_1 _10261_ (.B1(_04398_),
    .Y(_00428_),
    .A1(_04397_),
    .A2(net154));
 sg13g2_mux2_1 _10262_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .A1(_02248_),
    .S(_04393_),
    .X(_00429_));
 sg13g2_mux2_1 _10263_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .A1(net299),
    .S(_04393_),
    .X(_00430_));
 sg13g2_buf_1 _10264_ (.A(_04392_),
    .X(_04399_));
 sg13g2_mux2_1 _10265_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .A1(_03227_),
    .S(net152),
    .X(_00431_));
 sg13g2_mux2_1 _10266_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A1(_03230_),
    .S(net152),
    .X(_00432_));
 sg13g2_mux2_1 _10267_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(net152),
    .X(_00433_));
 sg13g2_mux2_1 _10268_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(net152),
    .X(_00434_));
 sg13g2_mux2_1 _10269_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .S(net152),
    .X(_00435_));
 sg13g2_mux2_1 _10270_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .S(net152),
    .X(_00436_));
 sg13g2_mux2_1 _10271_ (.A0(_01937_),
    .A1(_01794_),
    .S(_04399_),
    .X(_00437_));
 sg13g2_mux2_1 _10272_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .S(_04399_),
    .X(_00438_));
 sg13g2_mux2_1 _10273_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .S(net152),
    .X(_00439_));
 sg13g2_mux2_1 _10274_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S(net152),
    .X(_00440_));
 sg13g2_buf_1 _10275_ (.A(_04392_),
    .X(_04400_));
 sg13g2_mux2_1 _10276_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .S(net151),
    .X(_00441_));
 sg13g2_mux2_1 _10277_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .S(net151),
    .X(_00442_));
 sg13g2_mux2_1 _10278_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .S(net151),
    .X(_00443_));
 sg13g2_mux2_1 _10279_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .S(_04400_),
    .X(_00444_));
 sg13g2_mux2_1 _10280_ (.A0(_02407_),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .S(_04400_),
    .X(_00445_));
 sg13g2_nand2_1 _10281_ (.Y(_04401_),
    .A(_01174_),
    .B(_02369_));
 sg13g2_buf_2 _10282_ (.A(_04401_),
    .X(_04402_));
 sg13g2_nand2_1 _10283_ (.Y(_04403_),
    .A(_01675_),
    .B(_01775_));
 sg13g2_buf_2 _10284_ (.A(_04403_),
    .X(_04404_));
 sg13g2_nand2_1 _10285_ (.Y(_04405_),
    .A(_02477_),
    .B(_04404_));
 sg13g2_o21ai_1 _10286_ (.B1(_04405_),
    .Y(_04406_),
    .A1(_02496_),
    .A2(_04404_));
 sg13g2_nand2_1 _10287_ (.Y(_04407_),
    .A(net158),
    .B(_04402_));
 sg13g2_o21ai_1 _10288_ (.B1(_04407_),
    .Y(_04408_),
    .A1(_04402_),
    .A2(_04406_));
 sg13g2_nand2b_1 _10289_ (.Y(_04409_),
    .B(net183),
    .A_N(net153));
 sg13g2_nand2_1 _10290_ (.Y(_04410_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .B(net153));
 sg13g2_o21ai_1 _10291_ (.B1(_04410_),
    .Y(_00446_),
    .A1(_04408_),
    .A2(_04409_));
 sg13g2_mux2_1 _10292_ (.A0(_02752_),
    .A1(_01095_),
    .S(_04404_),
    .X(_04411_));
 sg13g2_nor2_1 _10293_ (.A(_04402_),
    .B(_04411_),
    .Y(_04412_));
 sg13g2_a21oi_1 _10294_ (.A1(_01057_),
    .A2(_04402_),
    .Y(_04413_),
    .B1(_04412_));
 sg13g2_nand2_1 _10295_ (.Y(_04414_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .B(net153));
 sg13g2_o21ai_1 _10296_ (.B1(_04414_),
    .Y(_00447_),
    .A1(_04409_),
    .A2(_04413_));
 sg13g2_nand2_1 _10297_ (.Y(_04415_),
    .A(_01796_),
    .B(net153));
 sg13g2_o21ai_1 _10298_ (.B1(_04415_),
    .Y(_00448_),
    .A1(_01997_),
    .A2(net154));
 sg13g2_nor2_1 _10299_ (.A(net170),
    .B(_01225_),
    .Y(_04416_));
 sg13g2_mux2_1 _10300_ (.A0(_02860_),
    .A1(_00930_),
    .S(_04404_),
    .X(_04417_));
 sg13g2_nor2_1 _10301_ (.A(_04402_),
    .B(_04417_),
    .Y(_04418_));
 sg13g2_a21oi_1 _10302_ (.A1(net163),
    .A2(_04402_),
    .Y(_04419_),
    .B1(_04418_));
 sg13g2_a22oi_1 _10303_ (.Y(_04420_),
    .B1(_04419_),
    .B2(_01544_),
    .A2(_04416_),
    .A1(\i_tinyqv.cpu.i_core.mstatus_mte ));
 sg13g2_nand2_1 _10304_ (.Y(_04421_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .B(net153));
 sg13g2_o21ai_1 _10305_ (.B1(_04421_),
    .Y(_00449_),
    .A1(net154),
    .A2(_04420_));
 sg13g2_nand2b_1 _10306_ (.Y(_04422_),
    .B(_04404_),
    .A_N(_00959_));
 sg13g2_o21ai_1 _10307_ (.B1(_04422_),
    .Y(_04423_),
    .A1(_02948_),
    .A2(_04404_));
 sg13g2_nand2_1 _10308_ (.Y(_04424_),
    .A(_01968_),
    .B(_04402_));
 sg13g2_o21ai_1 _10309_ (.B1(_04424_),
    .Y(_04425_),
    .A1(_04402_),
    .A2(_04423_));
 sg13g2_nor2_1 _10310_ (.A(_00089_),
    .B(net170),
    .Y(_04426_));
 sg13g2_a21oi_1 _10311_ (.A1(_01544_),
    .A2(_04425_),
    .Y(_04427_),
    .B1(_04426_));
 sg13g2_nand2_1 _10312_ (.Y(_04428_),
    .A(_02407_),
    .B(net153));
 sg13g2_o21ai_1 _10313_ (.B1(_04428_),
    .Y(_00450_),
    .A1(net154),
    .A2(_04427_));
 sg13g2_mux2_1 _10314_ (.A0(net300),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .S(net151),
    .X(_00451_));
 sg13g2_mux2_1 _10315_ (.A0(_02083_),
    .A1(_01897_),
    .S(net151),
    .X(_00452_));
 sg13g2_nand2_1 _10316_ (.Y(_04429_),
    .A(_01937_),
    .B(_04395_));
 sg13g2_o21ai_1 _10317_ (.B1(_04429_),
    .Y(_00453_),
    .A1(_02138_),
    .A2(net154));
 sg13g2_nand2_1 _10318_ (.Y(_04430_),
    .A(_01996_),
    .B(_04395_));
 sg13g2_o21ai_1 _10319_ (.B1(_04430_),
    .Y(_00454_),
    .A1(_02215_),
    .A2(net154));
 sg13g2_mux2_1 _10320_ (.A0(_02204_),
    .A1(_02050_),
    .S(net151),
    .X(_00455_));
 sg13g2_mux2_1 _10321_ (.A0(_02248_),
    .A1(_02083_),
    .S(net151),
    .X(_00456_));
 sg13g2_mux2_1 _10322_ (.A0(net299),
    .A1(_02137_),
    .S(net151),
    .X(_00457_));
 sg13g2_buf_1 _10323_ (.A(net232),
    .X(_04431_));
 sg13g2_mux2_1 _10324_ (.A0(net8),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .S(net213),
    .X(_00652_));
 sg13g2_mux2_1 _10325_ (.A0(net9),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .S(net231),
    .X(_00653_));
 sg13g2_mux2_1 _10326_ (.A0(net10),
    .A1(_04270_),
    .S(net231),
    .X(_00654_));
 sg13g2_or3_1 _10327_ (.A(_01768_),
    .B(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .C(_03321_),
    .X(_04432_));
 sg13g2_buf_2 _10328_ (.A(_04432_),
    .X(_04433_));
 sg13g2_a21o_1 _10329_ (.A2(_02699_),
    .A1(_01678_),
    .B1(_03323_),
    .X(_04434_));
 sg13g2_buf_1 _10330_ (.A(_04434_),
    .X(_04435_));
 sg13g2_nand2b_1 _10331_ (.Y(_04436_),
    .B(_00817_),
    .A_N(net278));
 sg13g2_a21o_1 _10332_ (.A2(_04436_),
    .A1(_02369_),
    .B1(_01677_),
    .X(_04437_));
 sg13g2_buf_1 _10333_ (.A(_04437_),
    .X(_04438_));
 sg13g2_o21ai_1 _10334_ (.B1(_02693_),
    .Y(_04439_),
    .A1(_04375_),
    .A2(_04438_));
 sg13g2_o21ai_1 _10335_ (.B1(_04435_),
    .Y(_04440_),
    .A1(_01057_),
    .A2(_04365_));
 sg13g2_a22oi_1 _10336_ (.Y(_04441_),
    .B1(_04440_),
    .B2(_01361_),
    .A2(_04439_),
    .A1(_04435_));
 sg13g2_nor2b_1 _10337_ (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ),
    .B_N(\i_tinyqv.cpu.i_core.interrupt_req[1] ),
    .Y(_04442_));
 sg13g2_nor3_1 _10338_ (.A(_01361_),
    .B(_02693_),
    .C(_04442_),
    .Y(_04443_));
 sg13g2_nor3_1 _10339_ (.A(_04433_),
    .B(_04441_),
    .C(_04443_),
    .Y(_00227_));
 sg13g2_o21ai_1 _10340_ (.B1(_02693_),
    .Y(_04444_),
    .A1(net158),
    .A2(_04438_));
 sg13g2_nand2b_1 _10341_ (.Y(_04445_),
    .B(net158),
    .A_N(_04365_));
 sg13g2_nand2_1 _10342_ (.Y(_04446_),
    .A(_04435_),
    .B(_04445_));
 sg13g2_a22oi_1 _10343_ (.Y(_04447_),
    .B1(_04446_),
    .B2(_01363_),
    .A2(_04444_),
    .A1(_04435_));
 sg13g2_nor2b_1 _10344_ (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ),
    .B_N(\i_tinyqv.cpu.i_core.interrupt_req[0] ),
    .Y(_04448_));
 sg13g2_nor3_1 _10345_ (.A(_01363_),
    .B(_02693_),
    .C(_04448_),
    .Y(_04449_));
 sg13g2_nor3_1 _10346_ (.A(_04433_),
    .B(_04447_),
    .C(_04449_),
    .Y(_00228_));
 sg13g2_and2_1 _10347_ (.A(_01678_),
    .B(_02696_),
    .X(_04450_));
 sg13g2_buf_1 _10348_ (.A(_04450_),
    .X(_04451_));
 sg13g2_o21ai_1 _10349_ (.B1(_04451_),
    .Y(_04452_),
    .A1(_01968_),
    .A2(_04365_));
 sg13g2_nor4_2 _10350_ (.A(net256),
    .B(_02649_),
    .C(_02695_),
    .Y(_04453_),
    .D(_04438_));
 sg13g2_a22oi_1 _10351_ (.Y(_04454_),
    .B1(_04453_),
    .B2(_01968_),
    .A2(_04452_),
    .A1(\i_tinyqv.cpu.i_core.mie[19] ));
 sg13g2_nor2_1 _10352_ (.A(_04433_),
    .B(_04454_),
    .Y(_00229_));
 sg13g2_o21ai_1 _10353_ (.B1(_04451_),
    .Y(_04455_),
    .A1(net128),
    .A2(_04365_));
 sg13g2_a22oi_1 _10354_ (.Y(_04456_),
    .B1(_04455_),
    .B2(\i_tinyqv.cpu.i_core.mie[18] ),
    .A2(_04453_),
    .A1(net128));
 sg13g2_nor2_1 _10355_ (.A(_04433_),
    .B(_04456_),
    .Y(_00230_));
 sg13g2_o21ai_1 _10356_ (.B1(_04451_),
    .Y(_04457_),
    .A1(_01057_),
    .A2(_04365_));
 sg13g2_a22oi_1 _10357_ (.Y(_04458_),
    .B1(_04457_),
    .B2(\i_tinyqv.cpu.i_core.mie[17] ),
    .A2(_04453_),
    .A1(_01057_));
 sg13g2_nor2_1 _10358_ (.A(_04433_),
    .B(_04458_),
    .Y(_00231_));
 sg13g2_nand2_1 _10359_ (.Y(_04459_),
    .A(_04445_),
    .B(_04451_));
 sg13g2_a22oi_1 _10360_ (.Y(_04460_),
    .B1(_04459_),
    .B2(\i_tinyqv.cpu.i_core.mie[16] ),
    .A2(_04453_),
    .A1(_01831_));
 sg13g2_nor2_1 _10361_ (.A(_04433_),
    .B(_04460_),
    .Y(_00232_));
 sg13g2_inv_1 _10362_ (.Y(_04461_),
    .A(_00168_));
 sg13g2_buf_1 _10363_ (.A(\i_debug_uart_tx.cycle_counter[1] ),
    .X(_04462_));
 sg13g2_nand4_1 _10364_ (.B(\i_debug_uart_tx.cycle_counter[0] ),
    .C(\i_debug_uart_tx.cycle_counter[2] ),
    .A(_04462_),
    .Y(_04463_),
    .D(\i_debug_uart_tx.cycle_counter[3] ));
 sg13g2_nor2_1 _10365_ (.A(_04461_),
    .B(_04463_),
    .Y(_04464_));
 sg13g2_buf_1 _10366_ (.A(_04464_),
    .X(_04465_));
 sg13g2_nor2b_1 _10367_ (.A(net217),
    .B_N(_00222_),
    .Y(_04466_));
 sg13g2_a21oi_1 _10368_ (.A1(\i_debug_uart_tx.cycle_counter[0] ),
    .A2(net217),
    .Y(_04467_),
    .B1(_04466_));
 sg13g2_nor3_1 _10369_ (.A(net229),
    .B(_04465_),
    .C(_04467_),
    .Y(_00234_));
 sg13g2_nor2b_1 _10370_ (.A(net217),
    .B_N(\i_debug_uart_tx.cycle_counter[0] ),
    .Y(_04468_));
 sg13g2_xnor2_1 _10371_ (.Y(_04469_),
    .A(_04462_),
    .B(_04468_));
 sg13g2_nor3_1 _10372_ (.A(net229),
    .B(_04465_),
    .C(_04469_),
    .Y(_00235_));
 sg13g2_nand2_1 _10373_ (.Y(_04470_),
    .A(_04462_),
    .B(_04468_));
 sg13g2_xor2_1 _10374_ (.B(_04470_),
    .A(\i_debug_uart_tx.cycle_counter[2] ),
    .X(_04471_));
 sg13g2_nor3_1 _10375_ (.A(net229),
    .B(net212),
    .C(_04471_),
    .Y(_00236_));
 sg13g2_nand3_1 _10376_ (.B(\i_debug_uart_tx.cycle_counter[0] ),
    .C(\i_debug_uart_tx.cycle_counter[2] ),
    .A(_04462_),
    .Y(_04472_));
 sg13g2_and2_1 _10377_ (.A(_04461_),
    .B(net217),
    .X(_04473_));
 sg13g2_o21ai_1 _10378_ (.B1(\i_debug_uart_tx.cycle_counter[3] ),
    .Y(_04474_),
    .A1(_04472_),
    .A2(_04473_));
 sg13g2_or3_1 _10379_ (.A(\i_debug_uart_tx.cycle_counter[3] ),
    .B(net217),
    .C(_04472_),
    .X(_04475_));
 sg13g2_a21oi_1 _10380_ (.A1(_04474_),
    .A2(_04475_),
    .Y(_00237_),
    .B1(_03063_));
 sg13g2_nand2_1 _10381_ (.Y(_04476_),
    .A(\i_debug_uart_tx.cycle_counter[4] ),
    .B(net217));
 sg13g2_o21ai_1 _10382_ (.B1(_04476_),
    .Y(_04477_),
    .A1(_00168_),
    .A2(_02561_));
 sg13g2_a22oi_1 _10383_ (.Y(_04478_),
    .B1(_04477_),
    .B2(_04463_),
    .A2(_04473_),
    .A1(\i_debug_uart_tx.cycle_counter[4] ));
 sg13g2_nor2_1 _10384_ (.A(_03063_),
    .B(_04478_),
    .Y(_00238_));
 sg13g2_inv_1 _10385_ (.Y(_04479_),
    .A(_00221_));
 sg13g2_and4_1 _10386_ (.A(_01407_),
    .B(_01404_),
    .C(_01415_),
    .D(_01401_),
    .X(_04480_));
 sg13g2_buf_1 _10387_ (.A(_04480_),
    .X(_04481_));
 sg13g2_nand3_1 _10388_ (.B(_01398_),
    .C(_04481_),
    .A(_01400_),
    .Y(_04482_));
 sg13g2_nor3_1 _10389_ (.A(net314),
    .B(_01396_),
    .C(_04482_),
    .Y(_04483_));
 sg13g2_or2_1 _10390_ (.X(_04484_),
    .B(_04483_),
    .A(net229));
 sg13g2_buf_2 _10391_ (.A(_04484_),
    .X(_04485_));
 sg13g2_nor2_1 _10392_ (.A(_04479_),
    .B(_04485_),
    .Y(_00252_));
 sg13g2_xnor2_1 _10393_ (.Y(_04486_),
    .A(net314),
    .B(_01407_));
 sg13g2_nor2_1 _10394_ (.A(_04485_),
    .B(_04486_),
    .Y(_00253_));
 sg13g2_nand2_1 _10395_ (.Y(_04487_),
    .A(net314),
    .B(_01407_));
 sg13g2_xnor2_1 _10396_ (.Y(_04488_),
    .A(_01406_),
    .B(_04487_));
 sg13g2_nor2_1 _10397_ (.A(_04485_),
    .B(_04488_),
    .Y(_00254_));
 sg13g2_nand3_1 _10398_ (.B(_01407_),
    .C(_01404_),
    .A(_01409_),
    .Y(_04489_));
 sg13g2_xor2_1 _10399_ (.B(_04489_),
    .A(_01415_),
    .X(_04490_));
 sg13g2_nor2_1 _10400_ (.A(_04485_),
    .B(_04490_),
    .Y(_00255_));
 sg13g2_nand4_1 _10401_ (.B(_01407_),
    .C(_01404_),
    .A(net314),
    .Y(_04491_),
    .D(_01415_));
 sg13g2_xor2_1 _10402_ (.B(_04491_),
    .A(_01401_),
    .X(_04492_));
 sg13g2_nor2_1 _10403_ (.A(_04485_),
    .B(_04492_),
    .Y(_00256_));
 sg13g2_nand2_1 _10404_ (.Y(_04493_),
    .A(net314),
    .B(_04481_));
 sg13g2_xor2_1 _10405_ (.B(_04493_),
    .A(_01400_),
    .X(_04494_));
 sg13g2_nor2_1 _10406_ (.A(_04485_),
    .B(_04494_),
    .Y(_00257_));
 sg13g2_nand3_1 _10407_ (.B(_01400_),
    .C(_04481_),
    .A(net314),
    .Y(_04495_));
 sg13g2_xor2_1 _10408_ (.B(_04495_),
    .A(_01398_),
    .X(_04496_));
 sg13g2_nor2_1 _10409_ (.A(_04485_),
    .B(_04496_),
    .Y(_00258_));
 sg13g2_inv_1 _10410_ (.Y(_04497_),
    .A(net314));
 sg13g2_nor3_1 _10411_ (.A(_04497_),
    .B(\i_pwm.pwm_count[7] ),
    .C(_04482_),
    .Y(_04498_));
 sg13g2_a21oi_1 _10412_ (.A1(\i_pwm.pwm_count[7] ),
    .A2(_04482_),
    .Y(_04499_),
    .B1(_04498_));
 sg13g2_nor2_1 _10413_ (.A(net229),
    .B(_04499_),
    .Y(_00259_));
 sg13g2_a21oi_1 _10414_ (.A1(\i_tinyqv.cpu.load_started ),
    .A2(_01360_),
    .Y(_04500_),
    .B1(_01771_));
 sg13g2_buf_1 _10415_ (.A(_01778_),
    .X(_04501_));
 sg13g2_nor2_1 _10416_ (.A(_01557_),
    .B(net118),
    .Y(_04502_));
 sg13g2_a21oi_1 _10417_ (.A1(\i_tinyqv.cpu.data_read_n[0] ),
    .A2(net118),
    .Y(_04503_),
    .B1(_04502_));
 sg13g2_nand2_1 _10418_ (.Y(_00360_),
    .A(_04500_),
    .B(_04503_));
 sg13g2_nand2b_1 _10419_ (.Y(_04504_),
    .B(net118),
    .A_N(\i_tinyqv.cpu.data_read_n[1] ));
 sg13g2_o21ai_1 _10420_ (.B1(_04504_),
    .Y(_04505_),
    .A1(_02509_),
    .A2(net118));
 sg13g2_nand2_1 _10421_ (.Y(_00361_),
    .A(_04500_),
    .B(_04505_));
 sg13g2_nor2_1 _10422_ (.A(\i_tinyqv.cpu.data_ready_latch ),
    .B(_01360_),
    .Y(_04506_));
 sg13g2_nor3_1 _10423_ (.A(net271),
    .B(_01213_),
    .C(_04506_),
    .Y(_00363_));
 sg13g2_nand2_1 _10424_ (.Y(_04507_),
    .A(_01678_),
    .B(_02670_));
 sg13g2_a21oi_1 _10425_ (.A1(_00817_),
    .A2(_01893_),
    .Y(_04508_),
    .B1(_04507_));
 sg13g2_nor4_1 _10426_ (.A(_01893_),
    .B(_02502_),
    .C(net186),
    .D(_04438_),
    .Y(_04509_));
 sg13g2_o21ai_1 _10427_ (.B1(net167),
    .Y(_04510_),
    .A1(net186),
    .A2(_04508_));
 sg13g2_a22oi_1 _10428_ (.Y(_04511_),
    .B1(_04510_),
    .B2(_01385_),
    .A2(_04509_),
    .A1(_04508_));
 sg13g2_nand2_2 _10429_ (.Y(_04512_),
    .A(_03270_),
    .B(net186));
 sg13g2_a21oi_1 _10430_ (.A1(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .A2(_04512_),
    .Y(_04513_),
    .B1(net169));
 sg13g2_a21oi_1 _10431_ (.A1(net169),
    .A2(_04511_),
    .Y(_04514_),
    .B1(_04513_));
 sg13g2_nand2b_1 _10432_ (.Y(_00411_),
    .B(_03322_),
    .A_N(_04514_));
 sg13g2_nor2_1 _10433_ (.A(_01385_),
    .B(_04512_),
    .Y(_04515_));
 sg13g2_nand3_1 _10434_ (.B(_02683_),
    .C(_04508_),
    .A(net169),
    .Y(_04516_));
 sg13g2_nor3_1 _10435_ (.A(_01893_),
    .B(_04438_),
    .C(_04516_),
    .Y(_04517_));
 sg13g2_a221oi_1 _10436_ (.B2(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .C1(_04517_),
    .B1(_04516_),
    .A1(_03270_),
    .Y(_04518_),
    .A2(net186));
 sg13g2_nor3_1 _10437_ (.A(_04433_),
    .B(_04515_),
    .C(_04518_),
    .Y(_00412_));
 sg13g2_nor2_1 _10438_ (.A(_02502_),
    .B(net183),
    .Y(_04519_));
 sg13g2_nor2b_1 _10439_ (.A(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .B_N(net169),
    .Y(_04520_));
 sg13g2_o21ai_1 _10440_ (.B1(_03322_),
    .Y(_00413_),
    .A1(_04519_),
    .A2(_04520_));
 sg13g2_a21oi_1 _10441_ (.A1(_02340_),
    .A2(_02362_),
    .Y(_04521_),
    .B1(_02361_));
 sg13g2_nand2_1 _10442_ (.Y(_04522_),
    .A(_02357_),
    .B(_02354_));
 sg13g2_o21ai_1 _10443_ (.B1(_02358_),
    .Y(_04523_),
    .A1(_02357_),
    .A2(_02354_));
 sg13g2_nand2_1 _10444_ (.Y(_04524_),
    .A(_04522_),
    .B(_04523_));
 sg13g2_nand2_1 _10445_ (.Y(_04525_),
    .A(_02346_),
    .B(_02352_));
 sg13g2_nor2_1 _10446_ (.A(_02346_),
    .B(_02352_),
    .Y(_04526_));
 sg13g2_a21o_1 _10447_ (.A2(_04525_),
    .A1(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .B1(_04526_),
    .X(_04527_));
 sg13g2_and2_1 _10448_ (.A(net299),
    .B(net114),
    .X(_04528_));
 sg13g2_nand2_1 _10449_ (.Y(_04529_),
    .A(net129),
    .B(net144));
 sg13g2_nand3_1 _10450_ (.B(_02350_),
    .C(net130),
    .A(_02303_),
    .Y(_04530_));
 sg13g2_o21ai_1 _10451_ (.B1(_04530_),
    .Y(_04531_),
    .A1(_02303_),
    .A2(_04529_));
 sg13g2_a22oi_1 _10452_ (.Y(_04532_),
    .B1(_04531_),
    .B2(net299),
    .A2(_01857_),
    .A1(net253));
 sg13g2_inv_1 _10453_ (.Y(_04533_),
    .A(_04532_));
 sg13g2_nand2_1 _10454_ (.Y(_04534_),
    .A(_02303_),
    .B(net129));
 sg13g2_nor3_1 _10455_ (.A(_04397_),
    .B(net130),
    .C(_04534_),
    .Y(_04535_));
 sg13g2_a22oi_1 _10456_ (.Y(_04536_),
    .B1(_04535_),
    .B2(_01833_),
    .A2(net130),
    .A1(_04394_));
 sg13g2_o21ai_1 _10457_ (.B1(_02350_),
    .Y(_04537_),
    .A1(net115),
    .A2(net144));
 sg13g2_a21oi_1 _10458_ (.A1(_01868_),
    .A2(_02305_),
    .Y(_04538_),
    .B1(_02350_));
 sg13g2_a221oi_1 _10459_ (.B2(_04394_),
    .C1(_04538_),
    .B1(_04537_),
    .A1(_01857_),
    .Y(_04539_),
    .A2(net130));
 sg13g2_o21ai_1 _10460_ (.B1(_04539_),
    .Y(_04540_),
    .A1(net299),
    .A2(_04536_));
 sg13g2_a21oi_1 _10461_ (.A1(net115),
    .A2(_04533_),
    .Y(_04541_),
    .B1(_04540_));
 sg13g2_xor2_1 _10462_ (.B(_04541_),
    .A(_04528_),
    .X(_04542_));
 sg13g2_xnor2_1 _10463_ (.Y(_04543_),
    .A(_04527_),
    .B(_04542_));
 sg13g2_xnor2_1 _10464_ (.Y(_04544_),
    .A(_04524_),
    .B(_04543_));
 sg13g2_xor2_1 _10465_ (.B(_04544_),
    .A(_04521_),
    .X(_00414_));
 sg13g2_nand2_1 _10466_ (.Y(_04545_),
    .A(_04524_),
    .B(_04543_));
 sg13g2_and2_1 _10467_ (.A(_02362_),
    .B(_04545_),
    .X(_04546_));
 sg13g2_and3_1 _10468_ (.X(_04547_),
    .A(_02332_),
    .B(_02339_),
    .C(_04546_));
 sg13g2_nand2_1 _10469_ (.Y(_04548_),
    .A(_02361_),
    .B(_04545_));
 sg13g2_o21ai_1 _10470_ (.B1(_04548_),
    .Y(_04549_),
    .A1(_04524_),
    .A2(_04543_));
 sg13g2_nor2_2 _10471_ (.A(_04547_),
    .B(_04549_),
    .Y(_04550_));
 sg13g2_nand2_2 _10472_ (.Y(_04551_),
    .A(_04527_),
    .B(_04542_));
 sg13g2_nand2_1 _10473_ (.Y(_04552_),
    .A(net253),
    .B(_01857_));
 sg13g2_nand3_1 _10474_ (.B(_02284_),
    .C(_01829_),
    .A(_02350_),
    .Y(_04553_));
 sg13g2_nand3_1 _10475_ (.B(_02284_),
    .C(net130),
    .A(net252),
    .Y(_04554_));
 sg13g2_o21ai_1 _10476_ (.B1(_04554_),
    .Y(_04555_),
    .A1(net252),
    .A2(net130));
 sg13g2_nor2_1 _10477_ (.A(net253),
    .B(_04553_),
    .Y(_04556_));
 sg13g2_a21oi_1 _10478_ (.A1(net253),
    .A2(_04555_),
    .Y(_04557_),
    .B1(_04556_));
 sg13g2_or2_1 _10479_ (.X(_04558_),
    .B(_04557_),
    .A(_02347_));
 sg13g2_o21ai_1 _10480_ (.B1(_04558_),
    .Y(_04559_),
    .A1(_04552_),
    .A2(_04553_));
 sg13g2_a21oi_2 _10481_ (.B1(_04559_),
    .Y(_04560_),
    .A2(_04541_),
    .A1(_04528_));
 sg13g2_nand2_1 _10482_ (.Y(_04561_),
    .A(net252),
    .B(_01868_));
 sg13g2_nand2_1 _10483_ (.Y(_04562_),
    .A(_01837_),
    .B(net114));
 sg13g2_nand2b_1 _10484_ (.Y(_04563_),
    .B(_01829_),
    .A_N(net114));
 sg13g2_o21ai_1 _10485_ (.B1(_04563_),
    .Y(_04564_),
    .A1(_04561_),
    .A2(_04562_));
 sg13g2_nand2_1 _10486_ (.Y(_04565_),
    .A(net253),
    .B(net114));
 sg13g2_a22oi_1 _10487_ (.Y(_04566_),
    .B1(_04565_),
    .B2(_04561_),
    .A2(_04564_),
    .A1(net253));
 sg13g2_nand2b_1 _10488_ (.Y(_04567_),
    .B(_04566_),
    .A_N(_04560_));
 sg13g2_inv_1 _10489_ (.Y(_04568_),
    .A(_04567_));
 sg13g2_nor2b_1 _10490_ (.A(_04566_),
    .B_N(_04560_),
    .Y(_04569_));
 sg13g2_nor2_1 _10491_ (.A(_04568_),
    .B(_04569_),
    .Y(_04570_));
 sg13g2_xnor2_1 _10492_ (.Y(_04571_),
    .A(_04551_),
    .B(_04570_));
 sg13g2_xnor2_1 _10493_ (.Y(_00415_),
    .A(_04550_),
    .B(_04571_));
 sg13g2_nand2_1 _10494_ (.Y(_04572_),
    .A(net114),
    .B(_04534_));
 sg13g2_o21ai_1 _10495_ (.B1(_04572_),
    .Y(_04573_),
    .A1(_04534_),
    .A2(_04563_));
 sg13g2_nand2_1 _10496_ (.Y(_04574_),
    .A(net252),
    .B(_04573_));
 sg13g2_inv_1 _10497_ (.Y(_04575_),
    .A(_04551_));
 sg13g2_nor2_1 _10498_ (.A(_04575_),
    .B(_04568_),
    .Y(_04576_));
 sg13g2_nand2_1 _10499_ (.Y(_04577_),
    .A(_04548_),
    .B(_04569_));
 sg13g2_nor2_1 _10500_ (.A(_04551_),
    .B(_04567_),
    .Y(_04578_));
 sg13g2_nand4_1 _10501_ (.B(_02339_),
    .C(_04546_),
    .A(_02332_),
    .Y(_04579_),
    .D(_04578_));
 sg13g2_o21ai_1 _10502_ (.B1(_04579_),
    .Y(_04580_),
    .A1(_04547_),
    .A2(_04577_));
 sg13g2_a221oi_1 _10503_ (.B2(_04550_),
    .C1(_04580_),
    .B1(_04576_),
    .A1(_04551_),
    .Y(_04581_),
    .A2(_04569_));
 sg13g2_xnor2_1 _10504_ (.Y(_00416_),
    .A(_04574_),
    .B(_04581_));
 sg13g2_or4_1 _10505_ (.A(_01286_),
    .B(net252),
    .C(_01893_),
    .D(_04560_),
    .X(_04582_));
 sg13g2_o21ai_1 _10506_ (.B1(_04582_),
    .Y(_04583_),
    .A1(_04563_),
    .A2(_04561_));
 sg13g2_nor2_1 _10507_ (.A(_01857_),
    .B(_04560_),
    .Y(_04584_));
 sg13g2_nand2_1 _10508_ (.Y(_04585_),
    .A(_04562_),
    .B(_04584_));
 sg13g2_nand2_1 _10509_ (.Y(_04586_),
    .A(_04572_),
    .B(_04585_));
 sg13g2_a22oi_1 _10510_ (.Y(_04587_),
    .B1(_04586_),
    .B2(net252),
    .A2(_04583_),
    .A1(net253));
 sg13g2_inv_1 _10511_ (.Y(_04588_),
    .A(_04563_));
 sg13g2_a22oi_1 _10512_ (.Y(_04589_),
    .B1(_04588_),
    .B2(_04584_),
    .A2(net114),
    .A1(_01857_));
 sg13g2_nand2_1 _10513_ (.Y(_04590_),
    .A(_01857_),
    .B(_04560_));
 sg13g2_nand3_1 _10514_ (.B(net114),
    .C(_04590_),
    .A(_04394_),
    .Y(_04591_));
 sg13g2_o21ai_1 _10515_ (.B1(_04591_),
    .Y(_04592_),
    .A1(_04394_),
    .A2(_04589_));
 sg13g2_nand2_1 _10516_ (.Y(_04593_),
    .A(net252),
    .B(_04592_));
 sg13g2_o21ai_1 _10517_ (.B1(_04593_),
    .Y(_04594_),
    .A1(_04550_),
    .A2(_04587_));
 sg13g2_a21o_1 _10518_ (.A2(_04590_),
    .A1(net253),
    .B1(_04584_),
    .X(_04595_));
 sg13g2_nand3_1 _10519_ (.B(net114),
    .C(_04595_),
    .A(net252),
    .Y(_04596_));
 sg13g2_o21ai_1 _10520_ (.B1(_04596_),
    .Y(_04597_),
    .A1(_04550_),
    .A2(_04593_));
 sg13g2_a21o_1 _10521_ (.A2(_04594_),
    .A1(_04575_),
    .B1(_04597_),
    .X(_00417_));
 sg13g2_xnor2_1 _10522_ (.Y(_04598_),
    .A(_01621_),
    .B(_01632_));
 sg13g2_buf_1 _10523_ (.A(_03595_),
    .X(_04599_));
 sg13g2_nand2_1 _10524_ (.Y(_04600_),
    .A(net84),
    .B(_04599_));
 sg13g2_nor3_1 _10525_ (.A(_01768_),
    .B(_04598_),
    .C(_04600_),
    .Y(_00581_));
 sg13g2_a21oi_1 _10526_ (.A1(_04256_),
    .A2(_04257_),
    .Y(_04601_),
    .B1(_01655_));
 sg13g2_nand3_1 _10527_ (.B(_04176_),
    .C(net311),
    .A(_01649_),
    .Y(_04602_));
 sg13g2_buf_1 _10528_ (.A(_04602_),
    .X(_04603_));
 sg13g2_buf_1 _10529_ (.A(_04603_),
    .X(_04604_));
 sg13g2_nand2_1 _10530_ (.Y(_04605_),
    .A(_01336_),
    .B(_04604_));
 sg13g2_a21oi_1 _10531_ (.A1(net72),
    .A2(_04605_),
    .Y(_04606_),
    .B1(net229));
 sg13g2_nor2b_1 _10532_ (.A(_04601_),
    .B_N(_04606_),
    .Y(_00615_));
 sg13g2_or2_1 _10533_ (.X(_04607_),
    .B(_04258_),
    .A(_04254_));
 sg13g2_buf_2 _10534_ (.A(_04607_),
    .X(_04608_));
 sg13g2_buf_1 _10535_ (.A(_04608_),
    .X(_04609_));
 sg13g2_nand3_1 _10536_ (.B(_04175_),
    .C(_04180_),
    .A(net247),
    .Y(_04610_));
 sg13g2_nor3_1 _10537_ (.A(net46),
    .B(_04269_),
    .C(_04610_),
    .Y(_00651_));
 sg13g2_inv_1 _10538_ (.Y(_04611_),
    .A(\addr[24] ));
 sg13g2_mux2_1 _10539_ (.A0(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ),
    .A1(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ),
    .S(_04090_),
    .X(_04612_));
 sg13g2_or4_1 _10540_ (.A(_01356_),
    .B(_04611_),
    .C(_03800_),
    .D(_04612_),
    .X(_04613_));
 sg13g2_and2_1 _10541_ (.A(net69),
    .B(_04613_),
    .X(_04614_));
 sg13g2_buf_8 _10542_ (.A(_04614_),
    .X(_04615_));
 sg13g2_nand2_1 _10543_ (.Y(_04616_),
    .A(net246),
    .B(_04170_));
 sg13g2_a22oi_1 _10544_ (.Y(_04617_),
    .B1(_04616_),
    .B2(_04603_),
    .A2(_04197_),
    .A1(_04287_));
 sg13g2_a21o_1 _10545_ (.A2(_04269_),
    .A1(_04175_),
    .B1(_04617_),
    .X(_04618_));
 sg13g2_buf_1 _10546_ (.A(_04618_),
    .X(_04619_));
 sg13g2_o21ai_1 _10547_ (.B1(_04619_),
    .Y(_04620_),
    .A1(_01651_),
    .A2(net45));
 sg13g2_nor3_1 _10548_ (.A(_01356_),
    .B(_04611_),
    .C(_03800_),
    .Y(_04621_));
 sg13g2_buf_2 _10549_ (.A(_04621_),
    .X(_04622_));
 sg13g2_inv_1 _10550_ (.Y(_04623_),
    .A(_04273_));
 sg13g2_nor2_1 _10551_ (.A(_04623_),
    .B(_04283_),
    .Y(_04624_));
 sg13g2_buf_1 _10552_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .X(_04625_));
 sg13g2_o21ai_1 _10553_ (.B1(_04192_),
    .Y(_04626_),
    .A1(net245),
    .A2(_04625_));
 sg13g2_mux2_1 _10554_ (.A0(_00165_),
    .A1(_04626_),
    .S(_03811_),
    .X(_04627_));
 sg13g2_nand2_1 _10555_ (.Y(_04628_),
    .A(_04603_),
    .B(_04172_));
 sg13g2_a21oi_1 _10556_ (.A1(_04185_),
    .A2(_04627_),
    .Y(_04629_),
    .B1(_04628_));
 sg13g2_nor2_1 _10557_ (.A(_04173_),
    .B(_04262_),
    .Y(_04630_));
 sg13g2_a21oi_1 _10558_ (.A1(_04624_),
    .A2(_04629_),
    .Y(_04631_),
    .B1(_04630_));
 sg13g2_o21ai_1 _10559_ (.B1(_04631_),
    .Y(_04632_),
    .A1(net191),
    .A2(_04622_));
 sg13g2_a221oi_1 _10560_ (.B2(_04619_),
    .C1(net46),
    .B1(_04632_),
    .A1(_04176_),
    .Y(_00655_),
    .A2(_04620_));
 sg13g2_nor2_1 _10561_ (.A(net191),
    .B(net45),
    .Y(_04633_));
 sg13g2_nor2_1 _10562_ (.A(net246),
    .B(_04619_),
    .Y(_04634_));
 sg13g2_nor2_1 _10563_ (.A(net191),
    .B(_04622_),
    .Y(_04635_));
 sg13g2_inv_1 _10564_ (.Y(_04636_),
    .A(_04625_));
 sg13g2_a21oi_1 _10565_ (.A1(_04192_),
    .A2(_04636_),
    .Y(_04637_),
    .B1(_03809_));
 sg13g2_nor2_1 _10566_ (.A(net312),
    .B(_04170_),
    .Y(_04638_));
 sg13g2_nand2_1 _10567_ (.Y(_04639_),
    .A(net246),
    .B(_04638_));
 sg13g2_nand2_1 _10568_ (.Y(_04640_),
    .A(net246),
    .B(_04177_));
 sg13g2_nand2_1 _10569_ (.Y(_04641_),
    .A(net245),
    .B(_04640_));
 sg13g2_o21ai_1 _10570_ (.B1(_04641_),
    .Y(_04642_),
    .A1(_04637_),
    .A2(_04639_));
 sg13g2_o21ai_1 _10571_ (.B1(_04266_),
    .Y(_04643_),
    .A1(_04270_),
    .A2(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ));
 sg13g2_a21oi_1 _10572_ (.A1(_04262_),
    .A2(_04643_),
    .Y(_04644_),
    .B1(net193));
 sg13g2_a21oi_1 _10573_ (.A1(_04624_),
    .A2(_04642_),
    .Y(_04645_),
    .B1(_04644_));
 sg13g2_nand2_1 _10574_ (.Y(_04646_),
    .A(_04619_),
    .B(_04645_));
 sg13g2_nor2_1 _10575_ (.A(_04635_),
    .B(_04646_),
    .Y(_04647_));
 sg13g2_nor4_1 _10576_ (.A(_04608_),
    .B(_04633_),
    .C(_04634_),
    .D(_04647_),
    .Y(_00656_));
 sg13g2_nand2_2 _10577_ (.Y(_04648_),
    .A(_04177_),
    .B(_04175_));
 sg13g2_nor4_1 _10578_ (.A(net245),
    .B(net247),
    .C(_04625_),
    .D(_04648_),
    .Y(_04649_));
 sg13g2_a21oi_1 _10579_ (.A1(net245),
    .A2(_04648_),
    .Y(_04650_),
    .B1(net246));
 sg13g2_or2_1 _10580_ (.X(_04651_),
    .B(_04650_),
    .A(_04649_));
 sg13g2_nor4_1 _10581_ (.A(net275),
    .B(_04176_),
    .C(net311),
    .D(_04648_),
    .Y(_04652_));
 sg13g2_a21oi_1 _10582_ (.A1(net311),
    .A2(_04651_),
    .Y(_04653_),
    .B1(_04652_));
 sg13g2_nor2_1 _10583_ (.A(_04177_),
    .B(_04619_),
    .Y(_04654_));
 sg13g2_a21oi_1 _10584_ (.A1(_04619_),
    .A2(_04653_),
    .Y(_04655_),
    .B1(_04654_));
 sg13g2_nand3b_1 _10585_ (.B(_01653_),
    .C(_04170_),
    .Y(_04656_),
    .A_N(net45));
 sg13g2_a21oi_1 _10586_ (.A1(_04655_),
    .A2(_04656_),
    .Y(_00657_),
    .B1(net46));
 sg13g2_nand3_1 _10587_ (.B(_01351_),
    .C(_03798_),
    .A(net230),
    .Y(_04657_));
 sg13g2_nand4_1 _10588_ (.B(_04622_),
    .C(net45),
    .A(net72),
    .Y(_04658_),
    .D(_04657_));
 sg13g2_nand2b_1 _10589_ (.Y(_04659_),
    .B(_04169_),
    .A_N(_04615_));
 sg13g2_a21oi_1 _10590_ (.A1(_04658_),
    .A2(_04659_),
    .Y(_00658_),
    .B1(_04609_));
 sg13g2_inv_1 _10591_ (.Y(_04660_),
    .A(_04628_));
 sg13g2_a21o_1 _10592_ (.A2(_04613_),
    .A1(net69),
    .B1(_04660_),
    .X(_04661_));
 sg13g2_buf_1 _10593_ (.A(_04661_),
    .X(_04662_));
 sg13g2_a21o_1 _10594_ (.A2(_04648_),
    .A1(_04269_),
    .B1(net246),
    .X(_04663_));
 sg13g2_o21ai_1 _10595_ (.B1(_04663_),
    .Y(_04664_),
    .A1(_04176_),
    .A2(_04648_));
 sg13g2_a21oi_1 _10596_ (.A1(_04176_),
    .A2(_04640_),
    .Y(_04665_),
    .B1(_04269_));
 sg13g2_a21oi_2 _10597_ (.B1(_04665_),
    .Y(_04666_),
    .A2(_04664_),
    .A1(_03809_));
 sg13g2_nand2_1 _10598_ (.Y(_04667_),
    .A(_04662_),
    .B(_04666_));
 sg13g2_and4_1 _10599_ (.A(_04174_),
    .B(net191),
    .C(_04272_),
    .D(_04666_),
    .X(_04668_));
 sg13g2_a221oi_1 _10600_ (.B2(_04662_),
    .C1(net46),
    .B1(_04668_),
    .A1(_04207_),
    .Y(_00661_),
    .A2(_04667_));
 sg13g2_nand2_1 _10601_ (.Y(_04669_),
    .A(net246),
    .B(net311));
 sg13g2_nor2_1 _10602_ (.A(net312),
    .B(_04168_),
    .Y(_04670_));
 sg13g2_a22oi_1 _10603_ (.Y(_04671_),
    .B1(_04625_),
    .B2(_04670_),
    .A2(_04177_),
    .A1(net245));
 sg13g2_o21ai_1 _10604_ (.B1(_04208_),
    .Y(_04672_),
    .A1(_04669_),
    .A2(_04671_));
 sg13g2_nand3_1 _10605_ (.B(_04207_),
    .C(_04672_),
    .A(_04206_),
    .Y(_04673_));
 sg13g2_o21ai_1 _10606_ (.B1(_04673_),
    .Y(_04674_),
    .A1(_04206_),
    .A2(_04207_));
 sg13g2_nand3_1 _10607_ (.B(_04272_),
    .C(_04674_),
    .A(net191),
    .Y(_04675_));
 sg13g2_nor2_1 _10608_ (.A(_04608_),
    .B(_04675_),
    .Y(_04676_));
 sg13g2_nor2_1 _10609_ (.A(_04206_),
    .B(_04608_),
    .Y(_04677_));
 sg13g2_mux2_1 _10610_ (.A0(_04676_),
    .A1(_04677_),
    .S(_04667_),
    .X(_00662_));
 sg13g2_a21o_1 _10611_ (.A2(_04666_),
    .A1(_04662_),
    .B1(_04208_),
    .X(_04678_));
 sg13g2_nor2_1 _10612_ (.A(_01651_),
    .B(_04648_),
    .Y(_04679_));
 sg13g2_o21ai_1 _10613_ (.B1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .Y(_04680_),
    .A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .A2(_04174_));
 sg13g2_nor2b_1 _10614_ (.A(_04680_),
    .B_N(_04272_),
    .Y(_04681_));
 sg13g2_o21ai_1 _10615_ (.B1(net191),
    .Y(_04682_),
    .A1(_04679_),
    .A2(_04681_));
 sg13g2_o21ai_1 _10616_ (.B1(_04682_),
    .Y(_04683_),
    .A1(net191),
    .A2(_04622_));
 sg13g2_nand3_1 _10617_ (.B(_04666_),
    .C(_04683_),
    .A(_04662_),
    .Y(_04684_));
 sg13g2_a21oi_1 _10618_ (.A1(_04678_),
    .A2(_04684_),
    .Y(_00663_),
    .B1(net46));
 sg13g2_nand3b_1 _10619_ (.B(_01653_),
    .C(_03808_),
    .Y(_04685_),
    .A_N(net45));
 sg13g2_nand2_1 _10620_ (.Y(_04686_),
    .A(_04255_),
    .B(_04660_));
 sg13g2_a21oi_1 _10621_ (.A1(_04685_),
    .A2(_04686_),
    .Y(_00667_),
    .B1(net46));
 sg13g2_o21ai_1 _10622_ (.B1(_04177_),
    .Y(_04687_),
    .A1(net311),
    .A2(_00165_));
 sg13g2_nand2b_1 _10623_ (.Y(_04688_),
    .B(_01650_),
    .A_N(_04266_));
 sg13g2_nand3_1 _10624_ (.B(_00165_),
    .C(_04688_),
    .A(_04176_),
    .Y(_04689_));
 sg13g2_o21ai_1 _10625_ (.B1(_04689_),
    .Y(_04690_),
    .A1(_04176_),
    .A2(_04687_));
 sg13g2_a21oi_1 _10626_ (.A1(_01648_),
    .A2(_04690_),
    .Y(_04691_),
    .B1(_01653_));
 sg13g2_nand2_1 _10627_ (.Y(_04692_),
    .A(_04273_),
    .B(_04691_));
 sg13g2_o21ai_1 _10628_ (.B1(_04692_),
    .Y(_04693_),
    .A1(_04273_),
    .A2(_04638_));
 sg13g2_a21oi_1 _10629_ (.A1(_04269_),
    .A2(_04623_),
    .Y(_04694_),
    .B1(_04279_));
 sg13g2_nand2b_1 _10630_ (.Y(_04695_),
    .B(net191),
    .A_N(_04269_));
 sg13g2_o21ai_1 _10631_ (.B1(_04695_),
    .Y(_04696_),
    .A1(net275),
    .A2(_04694_));
 sg13g2_a21oi_1 _10632_ (.A1(_04269_),
    .A2(_04693_),
    .Y(_04697_),
    .B1(_04696_));
 sg13g2_a21oi_1 _10633_ (.A1(net45),
    .A2(_04697_),
    .Y(_04698_),
    .B1(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ));
 sg13g2_nor4_1 _10634_ (.A(net275),
    .B(net245),
    .C(_03809_),
    .D(_04625_),
    .Y(_04699_));
 sg13g2_nand4_1 _10635_ (.B(net193),
    .C(_04275_),
    .A(_04266_),
    .Y(_04700_),
    .D(_04699_));
 sg13g2_nand3_1 _10636_ (.B(_04697_),
    .C(_04700_),
    .A(_04604_),
    .Y(_04701_));
 sg13g2_o21ai_1 _10637_ (.B1(_04701_),
    .Y(_04702_),
    .A1(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .A2(_01653_));
 sg13g2_nor3_1 _10638_ (.A(net46),
    .B(_04698_),
    .C(_04702_),
    .Y(_00668_));
 sg13g2_mux2_1 _10639_ (.A0(_04625_),
    .A1(_04622_),
    .S(net45),
    .X(_04703_));
 sg13g2_or2_1 _10640_ (.X(_00669_),
    .B(_04703_),
    .A(net46));
 sg13g2_nand4_1 _10641_ (.B(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ),
    .C(net69),
    .A(_04090_),
    .Y(_04704_),
    .D(_04622_));
 sg13g2_o21ai_1 _10642_ (.B1(_04704_),
    .Y(_04705_),
    .A1(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .A2(_04615_));
 sg13g2_nand2b_1 _10643_ (.Y(_00678_),
    .B(_04705_),
    .A_N(_04609_));
 sg13g2_nand2b_1 _10644_ (.Y(_04706_),
    .B(_04622_),
    .A_N(_04090_));
 sg13g2_mux2_1 _10645_ (.A0(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .A1(_04706_),
    .S(net45),
    .X(_04707_));
 sg13g2_or2_1 _10646_ (.X(_00679_),
    .B(_04707_),
    .A(_04608_));
 sg13g2_nand2_1 _10647_ (.Y(_04708_),
    .A(net318),
    .B(_01645_));
 sg13g2_or2_1 _10648_ (.X(_04709_),
    .B(_01296_),
    .A(_01335_));
 sg13g2_a22oi_1 _10649_ (.Y(_04710_),
    .B1(_04329_),
    .B2(_01305_),
    .A2(_04304_),
    .A1(_02531_));
 sg13g2_nand2b_1 _10650_ (.Y(_04711_),
    .B(_03930_),
    .A_N(_04710_));
 sg13g2_o21ai_1 _10651_ (.B1(_01339_),
    .Y(_04712_),
    .A1(_02524_),
    .A2(net61));
 sg13g2_nand4_1 _10652_ (.B(_04709_),
    .C(_04711_),
    .A(_04308_),
    .Y(_04713_),
    .D(_04712_));
 sg13g2_nand2b_1 _10653_ (.Y(_04714_),
    .B(net68),
    .A_N(net229));
 sg13g2_a21oi_1 _10654_ (.A1(_04708_),
    .A2(_04713_),
    .Y(_00713_),
    .B1(_04714_));
 sg13g2_nand2_1 _10655_ (.Y(_04715_),
    .A(net318),
    .B(_04709_));
 sg13g2_nor4_1 _10656_ (.A(net322),
    .B(_02524_),
    .C(net61),
    .D(_04715_),
    .Y(_04716_));
 sg13g2_a21oi_1 _10657_ (.A1(_01298_),
    .A2(_04715_),
    .Y(_04717_),
    .B1(_04716_));
 sg13g2_nor2_1 _10658_ (.A(_04714_),
    .B(_04717_),
    .Y(_00714_));
 sg13g2_inv_1 _10659_ (.Y(_04718_),
    .A(_00225_));
 sg13g2_inv_1 _10660_ (.Y(_04719_),
    .A(net316));
 sg13g2_nor2_1 _10661_ (.A(net317),
    .B(net315),
    .Y(_04720_));
 sg13g2_nand2_1 _10662_ (.Y(_04721_),
    .A(_04719_),
    .B(_04720_));
 sg13g2_nand3_1 _10663_ (.B(net317),
    .C(_01370_),
    .A(net316),
    .Y(_04722_));
 sg13g2_a21oi_1 _10664_ (.A1(_04721_),
    .A2(_04722_),
    .Y(_04723_),
    .B1(_01368_));
 sg13g2_or3_1 _10665_ (.A(_03062_),
    .B(_04356_),
    .C(_04723_),
    .X(_04724_));
 sg13g2_buf_1 _10666_ (.A(_04724_),
    .X(_04725_));
 sg13g2_buf_1 _10667_ (.A(_04725_),
    .X(_04726_));
 sg13g2_nor2_1 _10668_ (.A(_04718_),
    .B(net150),
    .Y(_00716_));
 sg13g2_and4_1 _10669_ (.A(_04351_),
    .B(_04344_),
    .C(_04352_),
    .D(_04348_),
    .X(_04727_));
 sg13g2_and2_1 _10670_ (.A(\i_uart_rx.cycle_counter[6] ),
    .B(_04727_),
    .X(_04728_));
 sg13g2_buf_1 _10671_ (.A(_04728_),
    .X(_04729_));
 sg13g2_nand3_1 _10672_ (.B(\i_uart_rx.cycle_counter[8] ),
    .C(_04729_),
    .A(_04349_),
    .Y(_04730_));
 sg13g2_nor2_1 _10673_ (.A(_04353_),
    .B(_04730_),
    .Y(_04731_));
 sg13g2_xnor2_1 _10674_ (.Y(_04732_),
    .A(\i_uart_rx.cycle_counter[10] ),
    .B(_04731_));
 sg13g2_nor2_1 _10675_ (.A(net150),
    .B(_04732_),
    .Y(_00717_));
 sg13g2_xnor2_1 _10676_ (.Y(_04733_),
    .A(_04345_),
    .B(_04346_));
 sg13g2_nor2_1 _10677_ (.A(net150),
    .B(_04733_),
    .Y(_00718_));
 sg13g2_nand2_1 _10678_ (.Y(_04734_),
    .A(_04345_),
    .B(_04346_));
 sg13g2_xor2_1 _10679_ (.B(_04734_),
    .A(_04351_),
    .X(_04735_));
 sg13g2_nor2_1 _10680_ (.A(net150),
    .B(_04735_),
    .Y(_00719_));
 sg13g2_nand3_1 _10681_ (.B(_04346_),
    .C(_04351_),
    .A(_04345_),
    .Y(_04736_));
 sg13g2_xor2_1 _10682_ (.B(_04736_),
    .A(\i_uart_rx.cycle_counter[3] ),
    .X(_04737_));
 sg13g2_nor2_1 _10683_ (.A(net150),
    .B(_04737_),
    .Y(_00720_));
 sg13g2_nand2_1 _10684_ (.Y(_04738_),
    .A(_04351_),
    .B(_04348_));
 sg13g2_xor2_1 _10685_ (.B(_04738_),
    .A(_04352_),
    .X(_04739_));
 sg13g2_nor2_1 _10686_ (.A(net150),
    .B(_04739_),
    .Y(_00721_));
 sg13g2_nand3_1 _10687_ (.B(_04352_),
    .C(_04348_),
    .A(_04351_),
    .Y(_04740_));
 sg13g2_xor2_1 _10688_ (.B(_04740_),
    .A(_04344_),
    .X(_04741_));
 sg13g2_nor2_1 _10689_ (.A(_04726_),
    .B(_04741_),
    .Y(_00722_));
 sg13g2_xnor2_1 _10690_ (.Y(_04742_),
    .A(\i_uart_rx.cycle_counter[6] ),
    .B(_04727_));
 sg13g2_nor2_1 _10691_ (.A(net150),
    .B(_04742_),
    .Y(_00723_));
 sg13g2_xnor2_1 _10692_ (.Y(_04743_),
    .A(_04349_),
    .B(_04729_));
 sg13g2_nor2_1 _10693_ (.A(_04726_),
    .B(_04743_),
    .Y(_00724_));
 sg13g2_inv_1 _10694_ (.Y(_04744_),
    .A(\i_uart_rx.cycle_counter[8] ));
 sg13g2_nand2_1 _10695_ (.Y(_04745_),
    .A(_04349_),
    .B(_04729_));
 sg13g2_xnor2_1 _10696_ (.Y(_04746_),
    .A(_04744_),
    .B(_04745_));
 sg13g2_nor2_1 _10697_ (.A(net150),
    .B(_04746_),
    .Y(_00725_));
 sg13g2_xnor2_1 _10698_ (.Y(_04747_),
    .A(_04353_),
    .B(_04730_));
 sg13g2_nor2_1 _10699_ (.A(_04725_),
    .B(_04747_),
    .Y(_00726_));
 sg13g2_nand2_1 _10700_ (.Y(_04748_),
    .A(\i_uart_tx.cycle_counter[0] ),
    .B(_01382_));
 sg13g2_nand2_1 _10701_ (.Y(_04749_),
    .A(_00224_),
    .B(_02547_));
 sg13g2_inv_1 _10702_ (.Y(_04750_),
    .A(\i_uart_tx.cycle_counter[4] ));
 sg13g2_buf_1 _10703_ (.A(\i_uart_tx.cycle_counter[5] ),
    .X(_04751_));
 sg13g2_buf_1 _10704_ (.A(\i_uart_tx.cycle_counter[2] ),
    .X(_04752_));
 sg13g2_buf_1 _10705_ (.A(\i_uart_tx.cycle_counter[8] ),
    .X(_04753_));
 sg13g2_inv_1 _10706_ (.Y(_04754_),
    .A(\i_uart_tx.cycle_counter[9] ));
 sg13g2_or4_1 _10707_ (.A(\i_uart_tx.cycle_counter[7] ),
    .B(\i_uart_tx.cycle_counter[6] ),
    .C(_04753_),
    .D(_04754_),
    .X(_04755_));
 sg13g2_nand2_1 _10708_ (.Y(_04756_),
    .A(\i_uart_tx.cycle_counter[0] ),
    .B(\i_uart_tx.cycle_counter[1] ));
 sg13g2_nor4_1 _10709_ (.A(_04752_),
    .B(\i_uart_tx.cycle_counter[10] ),
    .C(_04755_),
    .D(_04756_),
    .Y(_04757_));
 sg13g2_and4_1 _10710_ (.A(\i_uart_tx.cycle_counter[3] ),
    .B(_04750_),
    .C(_04751_),
    .D(_04757_),
    .X(_04758_));
 sg13g2_buf_1 _10711_ (.A(_04758_),
    .X(_04759_));
 sg13g2_or2_1 _10712_ (.X(_04760_),
    .B(net190),
    .A(_03062_));
 sg13g2_buf_1 _10713_ (.A(_04760_),
    .X(_04761_));
 sg13g2_a21oi_1 _10714_ (.A1(_04748_),
    .A2(_04749_),
    .Y(_00742_),
    .B1(_04761_));
 sg13g2_buf_1 _10715_ (.A(_04761_),
    .X(_04762_));
 sg13g2_inv_1 _10716_ (.Y(_04763_),
    .A(\i_uart_tx.cycle_counter[7] ));
 sg13g2_nor2_1 _10717_ (.A(_01382_),
    .B(_04756_),
    .Y(_04764_));
 sg13g2_nand3_1 _10718_ (.B(\i_uart_tx.cycle_counter[3] ),
    .C(_04764_),
    .A(_04752_),
    .Y(_04765_));
 sg13g2_nor2_1 _10719_ (.A(_04750_),
    .B(_04765_),
    .Y(_04766_));
 sg13g2_nand3_1 _10720_ (.B(\i_uart_tx.cycle_counter[6] ),
    .C(_04766_),
    .A(_04751_),
    .Y(_04767_));
 sg13g2_nor2_1 _10721_ (.A(_04763_),
    .B(_04767_),
    .Y(_04768_));
 sg13g2_nand3_1 _10722_ (.B(\i_uart_tx.cycle_counter[9] ),
    .C(_04768_),
    .A(_04753_),
    .Y(_04769_));
 sg13g2_xor2_1 _10723_ (.B(_04769_),
    .A(\i_uart_tx.cycle_counter[10] ),
    .X(_04770_));
 sg13g2_nor2_1 _10724_ (.A(net149),
    .B(_04770_),
    .Y(_00743_));
 sg13g2_and2_1 _10725_ (.A(\i_uart_tx.cycle_counter[0] ),
    .B(_02547_),
    .X(_04771_));
 sg13g2_xnor2_1 _10726_ (.Y(_04772_),
    .A(\i_uart_tx.cycle_counter[1] ),
    .B(_04771_));
 sg13g2_nor2_1 _10727_ (.A(net149),
    .B(_04772_),
    .Y(_00744_));
 sg13g2_xnor2_1 _10728_ (.Y(_04773_),
    .A(_04752_),
    .B(_04764_));
 sg13g2_nor2_1 _10729_ (.A(_04762_),
    .B(_04773_),
    .Y(_00745_));
 sg13g2_nand2_1 _10730_ (.Y(_04774_),
    .A(_04752_),
    .B(_04764_));
 sg13g2_xor2_1 _10731_ (.B(_04774_),
    .A(\i_uart_tx.cycle_counter[3] ),
    .X(_04775_));
 sg13g2_nor2_1 _10732_ (.A(net149),
    .B(_04775_),
    .Y(_00746_));
 sg13g2_xnor2_1 _10733_ (.Y(_04776_),
    .A(_04750_),
    .B(_04765_));
 sg13g2_nor2_1 _10734_ (.A(_04762_),
    .B(_04776_),
    .Y(_00747_));
 sg13g2_xnor2_1 _10735_ (.Y(_04777_),
    .A(_04751_),
    .B(_04766_));
 sg13g2_nor2_1 _10736_ (.A(net149),
    .B(_04777_),
    .Y(_00748_));
 sg13g2_nand2_1 _10737_ (.Y(_04778_),
    .A(_04751_),
    .B(_04766_));
 sg13g2_xor2_1 _10738_ (.B(_04778_),
    .A(\i_uart_tx.cycle_counter[6] ),
    .X(_04779_));
 sg13g2_nor2_1 _10739_ (.A(net149),
    .B(_04779_),
    .Y(_00749_));
 sg13g2_xnor2_1 _10740_ (.Y(_04780_),
    .A(_04763_),
    .B(_04767_));
 sg13g2_nor2_1 _10741_ (.A(net149),
    .B(_04780_),
    .Y(_00750_));
 sg13g2_xnor2_1 _10742_ (.Y(_04781_),
    .A(_04753_),
    .B(_04768_));
 sg13g2_nor2_1 _10743_ (.A(net149),
    .B(_04781_),
    .Y(_00751_));
 sg13g2_nand2_1 _10744_ (.Y(_04782_),
    .A(_04753_),
    .B(_04768_));
 sg13g2_xnor2_1 _10745_ (.Y(_04783_),
    .A(_04754_),
    .B(_04782_));
 sg13g2_nor2_1 _10746_ (.A(net149),
    .B(_04783_),
    .Y(_00752_));
 sg13g2_nor2_1 _10747_ (.A(net273),
    .B(_01348_),
    .Y(_04784_));
 sg13g2_nand4_1 _10748_ (.B(_02549_),
    .C(net217),
    .A(net272),
    .Y(_04785_),
    .D(_04784_));
 sg13g2_buf_1 _10749_ (.A(_04785_),
    .X(_04786_));
 sg13g2_inv_2 _10750_ (.Y(_04787_),
    .A(net117));
 sg13g2_nand2_1 _10751_ (.Y(_04788_),
    .A(net309),
    .B(_04787_));
 sg13g2_xnor2_1 _10752_ (.Y(_04789_),
    .A(_02558_),
    .B(_02556_));
 sg13g2_nand2_1 _10753_ (.Y(_04790_),
    .A(_04464_),
    .B(_04789_));
 sg13g2_buf_2 _10754_ (.A(_04790_),
    .X(_04791_));
 sg13g2_mux2_1 _10755_ (.A0(\i_debug_uart_tx.data_to_send[1] ),
    .A1(\i_debug_uart_tx.data_to_send[0] ),
    .S(_04791_),
    .X(_04792_));
 sg13g2_nand2_1 _10756_ (.Y(_04793_),
    .A(net117),
    .B(_04792_));
 sg13g2_inv_1 _10757_ (.Y(_04794_),
    .A(_01691_));
 sg13g2_buf_1 _10758_ (.A(_04794_),
    .X(_04795_));
 sg13g2_a21oi_1 _10759_ (.A1(_04788_),
    .A2(_04793_),
    .Y(_00239_),
    .B1(net211));
 sg13g2_nand2_1 _10760_ (.Y(_04796_),
    .A(net308),
    .B(_04787_));
 sg13g2_mux2_1 _10761_ (.A0(\i_debug_uart_tx.data_to_send[2] ),
    .A1(\i_debug_uart_tx.data_to_send[1] ),
    .S(_04791_),
    .X(_04797_));
 sg13g2_nand2_1 _10762_ (.Y(_04798_),
    .A(net117),
    .B(_04797_));
 sg13g2_a21oi_1 _10763_ (.A1(_04796_),
    .A2(_04798_),
    .Y(_00240_),
    .B1(net211));
 sg13g2_nand2_1 _10764_ (.Y(_04799_),
    .A(net307),
    .B(_04787_));
 sg13g2_mux2_1 _10765_ (.A0(\i_debug_uart_tx.data_to_send[3] ),
    .A1(\i_debug_uart_tx.data_to_send[2] ),
    .S(_04791_),
    .X(_04800_));
 sg13g2_nand2_1 _10766_ (.Y(_04801_),
    .A(net117),
    .B(_04800_));
 sg13g2_a21oi_1 _10767_ (.A1(_04799_),
    .A2(_04801_),
    .Y(_00241_),
    .B1(net211));
 sg13g2_nand2_1 _10768_ (.Y(_04802_),
    .A(_01724_),
    .B(_04787_));
 sg13g2_mux2_1 _10769_ (.A0(\i_debug_uart_tx.data_to_send[4] ),
    .A1(\i_debug_uart_tx.data_to_send[3] ),
    .S(_04791_),
    .X(_04803_));
 sg13g2_nand2_1 _10770_ (.Y(_04804_),
    .A(_04786_),
    .B(_04803_));
 sg13g2_a21oi_1 _10771_ (.A1(_04802_),
    .A2(_04804_),
    .Y(_00242_),
    .B1(net211));
 sg13g2_nand2_1 _10772_ (.Y(_04805_),
    .A(net306),
    .B(_04787_));
 sg13g2_mux2_1 _10773_ (.A0(\i_debug_uart_tx.data_to_send[5] ),
    .A1(\i_debug_uart_tx.data_to_send[4] ),
    .S(_04791_),
    .X(_04806_));
 sg13g2_nand2_1 _10774_ (.Y(_04807_),
    .A(_04786_),
    .B(_04806_));
 sg13g2_a21oi_1 _10775_ (.A1(_04805_),
    .A2(_04807_),
    .Y(_00243_),
    .B1(net211));
 sg13g2_nand2_1 _10776_ (.Y(_04808_),
    .A(net305),
    .B(_04787_));
 sg13g2_mux2_1 _10777_ (.A0(\i_debug_uart_tx.data_to_send[6] ),
    .A1(\i_debug_uart_tx.data_to_send[5] ),
    .S(_04791_),
    .X(_04809_));
 sg13g2_nand2_1 _10778_ (.Y(_04810_),
    .A(net117),
    .B(_04809_));
 sg13g2_a21oi_1 _10779_ (.A1(_04808_),
    .A2(_04810_),
    .Y(_00244_),
    .B1(net211));
 sg13g2_nand2_1 _10780_ (.Y(_04811_),
    .A(net304),
    .B(_04787_));
 sg13g2_mux2_1 _10781_ (.A0(\i_debug_uart_tx.data_to_send[7] ),
    .A1(\i_debug_uart_tx.data_to_send[6] ),
    .S(_04791_),
    .X(_04812_));
 sg13g2_nand2_1 _10782_ (.Y(_04813_),
    .A(net117),
    .B(_04812_));
 sg13g2_a21oi_1 _10783_ (.A1(_04811_),
    .A2(_04813_),
    .Y(_00245_),
    .B1(net211));
 sg13g2_or2_1 _10784_ (.X(_04814_),
    .B(net117),
    .A(_00205_));
 sg13g2_nand3_1 _10785_ (.B(net117),
    .C(_04791_),
    .A(\i_debug_uart_tx.data_to_send[7] ),
    .Y(_04815_));
 sg13g2_buf_1 _10786_ (.A(_04794_),
    .X(_04816_));
 sg13g2_a21oi_1 _10787_ (.A1(_04814_),
    .A2(_04815_),
    .Y(_00246_),
    .B1(net210));
 sg13g2_buf_1 _10788_ (.A(_04794_),
    .X(_04817_));
 sg13g2_a21oi_1 _10789_ (.A1(_02558_),
    .A2(net212),
    .Y(_04818_),
    .B1(_04787_));
 sg13g2_inv_1 _10790_ (.Y(_04819_),
    .A(_02558_));
 sg13g2_a21oi_1 _10791_ (.A1(_02554_),
    .A2(_04819_),
    .Y(_04820_),
    .B1(_02555_));
 sg13g2_nand2b_1 _10792_ (.Y(_04821_),
    .B(net212),
    .A_N(_04820_));
 sg13g2_o21ai_1 _10793_ (.B1(_04821_),
    .Y(_04822_),
    .A1(_02554_),
    .A2(_04818_));
 sg13g2_nand2_1 _10794_ (.Y(_04823_),
    .A(_02557_),
    .B(net212));
 sg13g2_o21ai_1 _10795_ (.B1(_04823_),
    .Y(_04824_),
    .A1(_02557_),
    .A2(_04822_));
 sg13g2_nor2_1 _10796_ (.A(net209),
    .B(_04824_),
    .Y(_00247_));
 sg13g2_nor2_1 _10797_ (.A(_04819_),
    .B(_02555_),
    .Y(_04825_));
 sg13g2_o21ai_1 _10798_ (.B1(net212),
    .Y(_04826_),
    .A1(_02557_),
    .A2(_04825_));
 sg13g2_nor2_1 _10799_ (.A(_02554_),
    .B(_04823_),
    .Y(_04827_));
 sg13g2_a21oi_1 _10800_ (.A1(_02554_),
    .A2(_04826_),
    .Y(_04828_),
    .B1(_04827_));
 sg13g2_nor2_1 _10801_ (.A(net209),
    .B(_04828_),
    .Y(_00248_));
 sg13g2_nand3_1 _10802_ (.B(_02554_),
    .C(net212),
    .A(_02557_),
    .Y(_04829_));
 sg13g2_xor2_1 _10803_ (.B(_04829_),
    .A(_02555_),
    .X(_04830_));
 sg13g2_nor2_1 _10804_ (.A(net209),
    .B(_04830_),
    .Y(_00249_));
 sg13g2_nand2b_1 _10805_ (.Y(_04831_),
    .B(_02555_),
    .A_N(_02557_));
 sg13g2_nand3_1 _10806_ (.B(net212),
    .C(_04831_),
    .A(_02554_),
    .Y(_04832_));
 sg13g2_nand4_1 _10807_ (.B(_04819_),
    .C(_02555_),
    .A(_02554_),
    .Y(_04833_),
    .D(net212));
 sg13g2_nand2b_1 _10808_ (.Y(_04834_),
    .B(_04833_),
    .A_N(_04825_));
 sg13g2_a22oi_1 _10809_ (.Y(_04835_),
    .B1(_04834_),
    .B2(_02557_),
    .A2(_04832_),
    .A1(_02558_));
 sg13g2_nor2_1 _10810_ (.A(_04817_),
    .B(_04835_),
    .Y(_00250_));
 sg13g2_a21oi_1 _10811_ (.A1(_02558_),
    .A2(\i_debug_uart_tx.data_to_send[0] ),
    .Y(_04836_),
    .B1(_02559_));
 sg13g2_nor3_1 _10812_ (.A(_02558_),
    .B(\i_debug_uart_tx.data_to_send[0] ),
    .C(_02556_),
    .Y(_04837_));
 sg13g2_a21oi_1 _10813_ (.A1(_02556_),
    .A2(_04836_),
    .Y(_04838_),
    .B1(_04837_));
 sg13g2_buf_1 _10814_ (.A(net232),
    .X(_04839_));
 sg13g2_nand2b_1 _10815_ (.Y(_00251_),
    .B(net208),
    .A_N(_04838_));
 sg13g2_nand4_1 _10816_ (.B(_01698_),
    .C(_02537_),
    .A(net272),
    .Y(_04840_),
    .D(_04784_));
 sg13g2_buf_1 _10817_ (.A(_04840_),
    .X(_04841_));
 sg13g2_nand2_1 _10818_ (.Y(_04842_),
    .A(\i_pwm.pwm_level[0] ),
    .B(net148));
 sg13g2_o21ai_1 _10819_ (.B1(_04842_),
    .Y(_04843_),
    .A1(_03256_),
    .A2(net148));
 sg13g2_and2_1 _10820_ (.A(net208),
    .B(_04843_),
    .X(_00260_));
 sg13g2_mux2_1 _10821_ (.A0(net308),
    .A1(\i_pwm.pwm_level[1] ),
    .S(net148),
    .X(_04844_));
 sg13g2_and2_1 _10822_ (.A(net208),
    .B(_04844_),
    .X(_00261_));
 sg13g2_mux2_1 _10823_ (.A0(net307),
    .A1(\i_pwm.pwm_level[2] ),
    .S(net148),
    .X(_04845_));
 sg13g2_and2_1 _10824_ (.A(net213),
    .B(_04845_),
    .X(_00262_));
 sg13g2_mux2_1 _10825_ (.A0(_01724_),
    .A1(\i_pwm.pwm_level[3] ),
    .S(net148),
    .X(_04846_));
 sg13g2_and2_1 _10826_ (.A(net213),
    .B(_04846_),
    .X(_00263_));
 sg13g2_mux2_1 _10827_ (.A0(net306),
    .A1(\i_pwm.pwm_level[4] ),
    .S(_04841_),
    .X(_04847_));
 sg13g2_and2_1 _10828_ (.A(net213),
    .B(_04847_),
    .X(_00264_));
 sg13g2_mux2_1 _10829_ (.A0(net305),
    .A1(\i_pwm.pwm_level[5] ),
    .S(net148),
    .X(_04848_));
 sg13g2_and2_1 _10830_ (.A(net213),
    .B(_04848_),
    .X(_00265_));
 sg13g2_mux2_1 _10831_ (.A0(net304),
    .A1(\i_pwm.pwm_level[6] ),
    .S(net148),
    .X(_04849_));
 sg13g2_and2_1 _10832_ (.A(net213),
    .B(_04849_),
    .X(_00266_));
 sg13g2_mux2_1 _10833_ (.A0(_01737_),
    .A1(\i_pwm.pwm_level[7] ),
    .S(net148),
    .X(_04850_));
 sg13g2_and2_1 _10834_ (.A(net213),
    .B(_04850_),
    .X(_00267_));
 sg13g2_inv_1 _10835_ (.Y(_04851_),
    .A(\i_spi.bits_remaining[0] ));
 sg13g2_or2_1 _10836_ (.X(_04852_),
    .B(\i_spi.bits_remaining[1] ),
    .A(\i_spi.bits_remaining[0] ));
 sg13g2_buf_1 _10837_ (.A(_04852_),
    .X(_04853_));
 sg13g2_nor2_2 _10838_ (.A(\i_spi.bits_remaining[2] ),
    .B(_04853_),
    .Y(_04854_));
 sg13g2_nor2_1 _10839_ (.A(_03083_),
    .B(_03072_),
    .Y(_04855_));
 sg13g2_nand2_1 _10840_ (.Y(_04856_),
    .A(_04854_),
    .B(_04855_));
 sg13g2_nand4_1 _10841_ (.B(_03086_),
    .C(_03087_),
    .A(_04851_),
    .Y(_04857_),
    .D(_04856_));
 sg13g2_nand2_1 _10842_ (.Y(_04858_),
    .A(\i_spi.bits_remaining[0] ),
    .B(_03088_));
 sg13g2_a21o_1 _10843_ (.A2(_03086_),
    .A1(_03083_),
    .B1(_04794_),
    .X(_04859_));
 sg13g2_a21oi_1 _10844_ (.A1(_04857_),
    .A2(_04858_),
    .Y(_00268_),
    .B1(_04859_));
 sg13g2_xor2_1 _10845_ (.B(_04857_),
    .A(\i_spi.bits_remaining[1] ),
    .X(_04860_));
 sg13g2_nor2_1 _10846_ (.A(_04859_),
    .B(_04860_),
    .Y(_00269_));
 sg13g2_or4_1 _10847_ (.A(\i_spi.bits_remaining[2] ),
    .B(_03088_),
    .C(_04853_),
    .D(_04855_),
    .X(_04861_));
 sg13g2_o21ai_1 _10848_ (.B1(\i_spi.bits_remaining[2] ),
    .Y(_04862_),
    .A1(_03088_),
    .A2(_04853_));
 sg13g2_a21oi_1 _10849_ (.A1(_04861_),
    .A2(_04862_),
    .Y(_00270_),
    .B1(_04859_));
 sg13g2_inv_1 _10850_ (.Y(_04863_),
    .A(_02550_));
 sg13g2_nand4_1 _10851_ (.B(_03086_),
    .C(_03087_),
    .A(_03072_),
    .Y(_04864_),
    .D(_04854_));
 sg13g2_o21ai_1 _10852_ (.B1(_04864_),
    .Y(_04865_),
    .A1(_03072_),
    .A2(_04854_));
 sg13g2_a21oi_1 _10853_ (.A1(_03095_),
    .A2(_04854_),
    .Y(_04866_),
    .B1(_03088_));
 sg13g2_o21ai_1 _10854_ (.B1(net231),
    .Y(_04867_),
    .A1(_03072_),
    .A2(_04866_));
 sg13g2_a21oi_1 _10855_ (.A1(_04863_),
    .A2(_04865_),
    .Y(_00271_),
    .B1(_04867_));
 sg13g2_inv_1 _10856_ (.Y(_04868_),
    .A(_03071_));
 sg13g2_nand2_1 _10857_ (.Y(_04869_),
    .A(_01315_),
    .B(_04868_));
 sg13g2_o21ai_1 _10858_ (.B1(_01716_),
    .Y(_04870_),
    .A1(_04856_),
    .A2(_04869_));
 sg13g2_a21oi_1 _10859_ (.A1(net228),
    .A2(_03080_),
    .Y(_00272_),
    .B1(_04870_));
 sg13g2_nand2_1 _10860_ (.Y(_04871_),
    .A(_03068_),
    .B(net228));
 sg13g2_nand3b_1 _10861_ (.B(net254),
    .C(_03071_),
    .Y(_04872_),
    .A_N(_03068_));
 sg13g2_a21oi_1 _10862_ (.A1(_04871_),
    .A2(_04872_),
    .Y(_00273_),
    .B1(net210));
 sg13g2_o21ai_1 _10863_ (.B1(net254),
    .Y(_04873_),
    .A1(_03068_),
    .A2(_04868_));
 sg13g2_nand3_1 _10864_ (.B(_03075_),
    .C(_03071_),
    .A(_03068_),
    .Y(_04874_));
 sg13g2_nor2_1 _10865_ (.A(\i_spi.clock_count[1] ),
    .B(_04874_),
    .Y(_04875_));
 sg13g2_a21oi_1 _10866_ (.A1(\i_spi.clock_count[1] ),
    .A2(_04873_),
    .Y(_04876_),
    .B1(_04875_));
 sg13g2_nor2_1 _10867_ (.A(net209),
    .B(_04876_),
    .Y(_00274_));
 sg13g2_or3_1 _10868_ (.A(_01348_),
    .B(_02538_),
    .C(_02542_),
    .X(_04877_));
 sg13g2_buf_1 _10869_ (.A(_04877_),
    .X(_04878_));
 sg13g2_nor2_1 _10870_ (.A(net309),
    .B(_04878_),
    .Y(_04879_));
 sg13g2_nor2b_1 _10871_ (.A(\i_spi.clock_divider[0] ),
    .B_N(_04878_),
    .Y(_04880_));
 sg13g2_o21ai_1 _10872_ (.B1(net208),
    .Y(_00275_),
    .A1(_04879_),
    .A2(_04880_));
 sg13g2_mux2_1 _10873_ (.A0(net308),
    .A1(\i_spi.clock_divider[1] ),
    .S(_04878_),
    .X(_04881_));
 sg13g2_and2_1 _10874_ (.A(_04431_),
    .B(_04881_),
    .X(_00276_));
 sg13g2_mux2_1 _10875_ (.A0(net307),
    .A1(\i_spi.read_latency ),
    .S(_04878_),
    .X(_04882_));
 sg13g2_and2_1 _10876_ (.A(_04431_),
    .B(_04882_),
    .X(_00286_));
 sg13g2_a21oi_1 _10877_ (.A1(_03073_),
    .A2(_04854_),
    .Y(_04883_),
    .B1(_04869_));
 sg13g2_a21o_1 _10878_ (.A2(_03071_),
    .A1(\i_spi.spi_clk_out ),
    .B1(_04883_),
    .X(_04884_));
 sg13g2_nor2_1 _10879_ (.A(net254),
    .B(_01315_),
    .Y(_04885_));
 sg13g2_a22oi_1 _10880_ (.Y(_04886_),
    .B1(_04885_),
    .B2(_03080_),
    .A2(_04884_),
    .A1(net254));
 sg13g2_nor2_1 _10881_ (.A(net209),
    .B(_04886_),
    .Y(_00287_));
 sg13g2_nor2_1 _10882_ (.A(_04856_),
    .B(_04869_),
    .Y(_04887_));
 sg13g2_o21ai_1 _10883_ (.B1(\i_spi.spi_select ),
    .Y(_04888_),
    .A1(net254),
    .A2(_03080_));
 sg13g2_a21oi_1 _10884_ (.A1(\i_spi.end_txn_reg ),
    .A2(_04887_),
    .Y(_04889_),
    .B1(_04794_));
 sg13g2_o21ai_1 _10885_ (.B1(_04889_),
    .Y(_00289_),
    .A1(_04887_),
    .A2(_04888_));
 sg13g2_buf_1 _10886_ (.A(_01542_),
    .X(_04890_));
 sg13g2_buf_1 _10887_ (.A(net226),
    .X(_04891_));
 sg13g2_nor2_1 _10888_ (.A(_00216_),
    .B(net73),
    .Y(_04892_));
 sg13g2_a221oi_1 _10889_ (.B2(net136),
    .C1(net92),
    .B1(_03394_),
    .A1(_01479_),
    .Y(_04893_),
    .A2(net89));
 sg13g2_nor3_1 _10890_ (.A(_03119_),
    .B(_03685_),
    .C(_04893_),
    .Y(_04894_));
 sg13g2_and2_1 _10891_ (.A(_01327_),
    .B(_03119_),
    .X(_04895_));
 sg13g2_nor3_1 _10892_ (.A(_03696_),
    .B(_04894_),
    .C(_04895_),
    .Y(_04896_));
 sg13g2_nor3_1 _10893_ (.A(net207),
    .B(_04892_),
    .C(_04896_),
    .Y(_00290_));
 sg13g2_nand2_1 _10894_ (.Y(_04897_),
    .A(_03123_),
    .B(_03119_));
 sg13g2_a21oi_1 _10895_ (.A1(_01484_),
    .A2(net112),
    .Y(_04898_),
    .B1(_03357_));
 sg13g2_nor3_1 _10896_ (.A(_03129_),
    .B(_03387_),
    .C(_04898_),
    .Y(_04899_));
 sg13g2_a221oi_1 _10897_ (.B2(_03401_),
    .C1(_04899_),
    .B1(_03394_),
    .A1(net171),
    .Y(_04900_),
    .A2(net89));
 sg13g2_inv_1 _10898_ (.Y(_04901_),
    .A(\i_tinyqv.cpu.additional_mem_ops[1] ));
 sg13g2_nor3_1 _10899_ (.A(_01327_),
    .B(_04901_),
    .C(_03121_),
    .Y(_04902_));
 sg13g2_a21o_1 _10900_ (.A2(_04900_),
    .A1(net73),
    .B1(_04902_),
    .X(_04903_));
 sg13g2_inv_1 _10901_ (.Y(_04904_),
    .A(_01327_));
 sg13g2_o21ai_1 _10902_ (.B1(_04897_),
    .Y(_04905_),
    .A1(_04904_),
    .A2(_03121_));
 sg13g2_a221oi_1 _10903_ (.B2(_04901_),
    .C1(net207),
    .B1(_04905_),
    .A1(_04897_),
    .Y(_00291_),
    .A2(_04903_));
 sg13g2_buf_1 _10904_ (.A(net226),
    .X(_04906_));
 sg13g2_nor2_1 _10905_ (.A(_01327_),
    .B(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .Y(_04907_));
 sg13g2_o21ai_1 _10906_ (.B1(_04897_),
    .Y(_04908_),
    .A1(_04907_),
    .A2(_03121_));
 sg13g2_buf_1 _10907_ (.A(_03125_),
    .X(_04909_));
 sg13g2_a22oi_1 _10908_ (.Y(_04910_),
    .B1(_03394_),
    .B2(_03720_),
    .A2(net89),
    .A1(net161));
 sg13g2_nor2_1 _10909_ (.A(net58),
    .B(_04910_),
    .Y(_04911_));
 sg13g2_a21oi_1 _10910_ (.A1(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .A2(_04908_),
    .Y(_04912_),
    .B1(_04911_));
 sg13g2_nor2_1 _10911_ (.A(net206),
    .B(_04912_),
    .Y(_00292_));
 sg13g2_and2_1 _10912_ (.A(net251),
    .B(_00220_),
    .X(_00297_));
 sg13g2_o21ai_1 _10913_ (.B1(_03657_),
    .Y(_04913_),
    .A1(_00900_),
    .A2(_02681_));
 sg13g2_inv_1 _10914_ (.Y(_00298_),
    .A(_04913_));
 sg13g2_xnor2_1 _10915_ (.Y(_04914_),
    .A(net236),
    .B(_01211_));
 sg13g2_nor2_1 _10916_ (.A(net206),
    .B(_04914_),
    .Y(_00299_));
 sg13g2_nor2b_2 _10917_ (.A(net118),
    .B_N(_03222_),
    .Y(_04915_));
 sg13g2_a22oi_1 _10918_ (.Y(_04916_),
    .B1(_04915_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A2(net118),
    .A1(\addr[24] ));
 sg13g2_nor2_1 _10919_ (.A(net206),
    .B(_04916_),
    .Y(_00316_));
 sg13g2_a22oi_1 _10920_ (.Y(_04917_),
    .B1(_04915_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .A2(net118),
    .A1(\addr[25] ));
 sg13g2_nor2_1 _10921_ (.A(net206),
    .B(_04917_),
    .Y(_00317_));
 sg13g2_a22oi_1 _10922_ (.Y(_04918_),
    .B1(_04915_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A2(_04501_),
    .A1(\addr[26] ));
 sg13g2_nor2_1 _10923_ (.A(_04906_),
    .B(_04918_),
    .Y(_00318_));
 sg13g2_a22oi_1 _10924_ (.Y(_04919_),
    .B1(_04915_),
    .B2(_02407_),
    .A2(_04501_),
    .A1(\addr[27] ));
 sg13g2_nor2_1 _10925_ (.A(_04906_),
    .B(_04919_),
    .Y(_00319_));
 sg13g2_nor2_1 _10926_ (.A(net159),
    .B(_04506_),
    .Y(_04920_));
 sg13g2_a21oi_1 _10927_ (.A1(\i_tinyqv.cpu.data_ready_core ),
    .A2(net159),
    .Y(_04921_),
    .B1(_04920_));
 sg13g2_nor2_1 _10928_ (.A(net206),
    .B(_04921_),
    .Y(_00362_));
 sg13g2_or2_1 _10929_ (.X(_04922_),
    .B(_01778_),
    .A(_01769_));
 sg13g2_buf_1 _10930_ (.A(_04922_),
    .X(_04923_));
 sg13g2_nor2_1 _10931_ (.A(_01556_),
    .B(_04923_),
    .Y(_04924_));
 sg13g2_nor2_1 _10932_ (.A(_01769_),
    .B(_01778_),
    .Y(_04925_));
 sg13g2_nor3_1 _10933_ (.A(_01306_),
    .B(_01360_),
    .C(_04925_),
    .Y(_04926_));
 sg13g2_o21ai_1 _10934_ (.B1(net251),
    .Y(_00364_),
    .A1(_04924_),
    .A2(_04926_));
 sg13g2_nor2_1 _10935_ (.A(_02509_),
    .B(_04923_),
    .Y(_04927_));
 sg13g2_nor3_1 _10936_ (.A(_01301_),
    .B(_01360_),
    .C(_04925_),
    .Y(_04928_));
 sg13g2_o21ai_1 _10937_ (.B1(net251),
    .Y(_00365_),
    .A1(_04927_),
    .A2(_04928_));
 sg13g2_nand2_1 _10938_ (.Y(_04929_),
    .A(net270),
    .B(net159));
 sg13g2_nand3_1 _10939_ (.B(_01326_),
    .C(_02367_),
    .A(net174),
    .Y(_04930_));
 sg13g2_buf_1 _10940_ (.A(net226),
    .X(_04931_));
 sg13g2_a21oi_1 _10941_ (.A1(_04929_),
    .A2(_04930_),
    .Y(_00366_),
    .B1(_04931_));
 sg13g2_a21oi_1 _10942_ (.A1(net270),
    .A2(net174),
    .Y(_04932_),
    .B1(_01774_));
 sg13g2_nor3_1 _10943_ (.A(net207),
    .B(_03120_),
    .C(_04932_),
    .Y(_00367_));
 sg13g2_nor2_1 _10944_ (.A(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .B(_01261_),
    .Y(_04933_));
 sg13g2_nor2b_1 _10945_ (.A(_04933_),
    .B_N(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .Y(_04934_));
 sg13g2_and2_1 _10946_ (.A(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .B(_04934_),
    .X(_04935_));
 sg13g2_buf_1 _10947_ (.A(_04935_),
    .X(_04936_));
 sg13g2_nand3_1 _10948_ (.B(_02698_),
    .C(_04936_),
    .A(_02870_),
    .Y(_04937_));
 sg13g2_nor2_1 _10949_ (.A(net206),
    .B(_04937_),
    .Y(_00368_));
 sg13g2_buf_1 _10950_ (.A(_01542_),
    .X(_04938_));
 sg13g2_nor3_1 _10951_ (.A(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .B(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .C(net167),
    .Y(_04939_));
 sg13g2_nor3_1 _10952_ (.A(net225),
    .B(_04934_),
    .C(_04939_),
    .Y(_00369_));
 sg13g2_xor2_1 _10953_ (.B(_04934_),
    .A(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .X(_04940_));
 sg13g2_and2_1 _10954_ (.A(net251),
    .B(_04940_),
    .X(_00370_));
 sg13g2_xnor2_1 _10955_ (.Y(_04941_),
    .A(_02870_),
    .B(_04936_));
 sg13g2_nor2_1 _10956_ (.A(net206),
    .B(_04941_),
    .Y(_00371_));
 sg13g2_nand2_1 _10957_ (.Y(_04942_),
    .A(_02870_),
    .B(_04936_));
 sg13g2_xor2_1 _10958_ (.B(_04942_),
    .A(_02698_),
    .X(_04943_));
 sg13g2_nor2_1 _10959_ (.A(net206),
    .B(_04943_),
    .Y(_00372_));
 sg13g2_inv_1 _10960_ (.Y(_04944_),
    .A(\i_tinyqv.cpu.i_core.i_instrret.data[3] ));
 sg13g2_and2_1 _10961_ (.A(_00218_),
    .B(net167),
    .X(_04945_));
 sg13g2_a21oi_1 _10962_ (.A1(_00219_),
    .A2(net170),
    .Y(_04946_),
    .B1(_04945_));
 sg13g2_and2_1 _10963_ (.A(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .B(_04946_),
    .X(_04947_));
 sg13g2_buf_1 _10964_ (.A(_04947_),
    .X(_04948_));
 sg13g2_nand3_1 _10965_ (.B(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .C(_04948_),
    .A(_02808_),
    .Y(_04949_));
 sg13g2_nor3_1 _10966_ (.A(net225),
    .B(_04944_),
    .C(_04949_),
    .Y(_00373_));
 sg13g2_buf_1 _10967_ (.A(_04890_),
    .X(_04950_));
 sg13g2_xor2_1 _10968_ (.B(_04946_),
    .A(_00170_),
    .X(_04951_));
 sg13g2_nor2_1 _10969_ (.A(net204),
    .B(_04951_),
    .Y(_00374_));
 sg13g2_xnor2_1 _10970_ (.Y(_04952_),
    .A(_02808_),
    .B(_04948_));
 sg13g2_nor2_1 _10971_ (.A(net204),
    .B(_04952_),
    .Y(_00375_));
 sg13g2_nand2_1 _10972_ (.Y(_04953_),
    .A(_02808_),
    .B(_04948_));
 sg13g2_xor2_1 _10973_ (.B(_04953_),
    .A(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .X(_04954_));
 sg13g2_nor2_1 _10974_ (.A(net204),
    .B(_04954_),
    .Y(_00376_));
 sg13g2_xnor2_1 _10975_ (.Y(_04955_),
    .A(_04944_),
    .B(_04949_));
 sg13g2_nor2_1 _10976_ (.A(net204),
    .B(_04955_),
    .Y(_00377_));
 sg13g2_buf_1 _10977_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .X(_04956_));
 sg13g2_nor4_1 _10978_ (.A(_04956_),
    .B(_00926_),
    .C(_00968_),
    .D(_01106_),
    .Y(_04957_));
 sg13g2_nor2_1 _10979_ (.A(_04512_),
    .B(_04957_),
    .Y(_04958_));
 sg13g2_nand2_1 _10980_ (.Y(_04959_),
    .A(\i_tinyqv.cpu.i_core.mie[18] ),
    .B(_01374_));
 sg13g2_nand3_1 _10981_ (.B(_04959_),
    .C(_01382_),
    .A(\i_tinyqv.cpu.i_core.mie[19] ),
    .Y(_04960_));
 sg13g2_nand2_1 _10982_ (.Y(_04961_),
    .A(_01362_),
    .B(_04960_));
 sg13g2_nand3_1 _10983_ (.B(_01364_),
    .C(_04961_),
    .A(_04956_),
    .Y(_04962_));
 sg13g2_o21ai_1 _10984_ (.B1(_03657_),
    .Y(_04963_),
    .A1(\i_tinyqv.cpu.i_core.mcause[0] ),
    .A2(_04519_));
 sg13g2_a21oi_1 _10985_ (.A1(_04958_),
    .A2(_04962_),
    .Y(_00383_),
    .B1(_04963_));
 sg13g2_o21ai_1 _10986_ (.B1(_04426_),
    .Y(_04964_),
    .A1(_01365_),
    .A2(_01383_));
 sg13g2_nor3_1 _10987_ (.A(\i_tinyqv.cpu.i_core.mcause[1] ),
    .B(_04416_),
    .C(_04426_),
    .Y(_04965_));
 sg13g2_nor2_1 _10988_ (.A(_04890_),
    .B(_04965_),
    .Y(_04966_));
 sg13g2_and2_1 _10989_ (.A(_04964_),
    .B(_04966_),
    .X(_00384_));
 sg13g2_and2_1 _10990_ (.A(_01117_),
    .B(_04519_),
    .X(_04967_));
 sg13g2_a21oi_1 _10991_ (.A1(\i_tinyqv.cpu.i_core.mcause[3] ),
    .A2(_04512_),
    .Y(_04968_),
    .B1(_04967_));
 sg13g2_nor3_1 _10992_ (.A(net225),
    .B(_04958_),
    .C(_04968_),
    .Y(_00385_));
 sg13g2_nand2_1 _10993_ (.Y(_04969_),
    .A(_04956_),
    .B(_04519_));
 sg13g2_nand2_1 _10994_ (.Y(_04970_),
    .A(\i_tinyqv.cpu.i_core.mcause[4] ),
    .B(_04512_));
 sg13g2_a21oi_1 _10995_ (.A1(_04969_),
    .A2(_04970_),
    .Y(_00386_),
    .B1(net205));
 sg13g2_nor2_1 _10996_ (.A(net159),
    .B(_04937_),
    .Y(_04971_));
 sg13g2_nand2_1 _10997_ (.Y(_04972_),
    .A(_00223_),
    .B(_04971_));
 sg13g2_o21ai_1 _10998_ (.B1(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .Y(_04973_),
    .A1(net159),
    .A2(_04937_));
 sg13g2_a21oi_1 _10999_ (.A1(_04972_),
    .A2(_04973_),
    .Y(_00423_),
    .B1(net205));
 sg13g2_nand2_1 _11000_ (.Y(_04974_),
    .A(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .B(_04971_));
 sg13g2_xor2_1 _11001_ (.B(_04974_),
    .A(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .X(_04975_));
 sg13g2_nor2_1 _11002_ (.A(net204),
    .B(_04975_),
    .Y(_00424_));
 sg13g2_nand3_1 _11003_ (.B(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .C(_04971_),
    .A(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .Y(_04976_));
 sg13g2_xor2_1 _11004_ (.B(_04976_),
    .A(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .X(_04977_));
 sg13g2_nor2_1 _11005_ (.A(net204),
    .B(_04977_),
    .Y(_00425_));
 sg13g2_nor2_2 _11006_ (.A(_01326_),
    .B(_01331_),
    .Y(_04978_));
 sg13g2_nor2_1 _11007_ (.A(_04978_),
    .B(_04600_),
    .Y(_04979_));
 sg13g2_buf_2 _11008_ (.A(_04979_),
    .X(_04980_));
 sg13g2_and2_1 _11009_ (.A(_01527_),
    .B(_01663_),
    .X(_04981_));
 sg13g2_buf_1 _11010_ (.A(_04981_),
    .X(_04982_));
 sg13g2_buf_1 _11011_ (.A(_04982_),
    .X(_04983_));
 sg13g2_buf_1 _11012_ (.A(_01770_),
    .X(_04984_));
 sg13g2_nor3_1 _11013_ (.A(net83),
    .B(_02967_),
    .C(_04982_),
    .Y(_04985_));
 sg13g2_a21o_1 _11014_ (.A2(net67),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .B1(_04985_),
    .X(_04986_));
 sg13g2_buf_1 _11015_ (.A(net84),
    .X(_04987_));
 sg13g2_buf_1 _11016_ (.A(_01559_),
    .X(_04988_));
 sg13g2_buf_1 _11017_ (.A(net189),
    .X(_04989_));
 sg13g2_nand2_1 _11018_ (.Y(_04990_),
    .A(net176),
    .B(_03247_));
 sg13g2_and2_1 _11019_ (.A(net233),
    .B(_00893_),
    .X(_04991_));
 sg13g2_buf_1 _11020_ (.A(_04991_),
    .X(_04992_));
 sg13g2_buf_1 _11021_ (.A(net188),
    .X(_04993_));
 sg13g2_nand2_1 _11022_ (.Y(_04994_),
    .A(net175),
    .B(_04103_));
 sg13g2_a21oi_1 _11023_ (.A1(_04990_),
    .A2(_04994_),
    .Y(_04995_),
    .B1(net82));
 sg13g2_a221oi_1 _11024_ (.B2(net82),
    .C1(_04995_),
    .B1(_04986_),
    .A1(net333),
    .Y(_04996_),
    .A2(_04980_));
 sg13g2_nor2_1 _11025_ (.A(_04950_),
    .B(_04996_),
    .Y(_00554_));
 sg13g2_buf_1 _11026_ (.A(_04980_),
    .X(_04997_));
 sg13g2_buf_1 _11027_ (.A(net77),
    .X(_04998_));
 sg13g2_nand3_1 _11028_ (.B(_02823_),
    .C(net71),
    .A(_04978_),
    .Y(_04999_));
 sg13g2_o21ai_1 _11029_ (.B1(_04999_),
    .Y(_05000_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .A2(net71));
 sg13g2_buf_1 _11030_ (.A(net84),
    .X(_05001_));
 sg13g2_buf_1 _11031_ (.A(net81),
    .X(_05002_));
 sg13g2_mux2_1 _11032_ (.A0(_03233_),
    .A1(_03919_),
    .S(_04993_),
    .X(_05003_));
 sg13g2_o21ai_1 _11033_ (.B1(net243),
    .Y(_05004_),
    .A1(net78),
    .A2(_05003_));
 sg13g2_a221oi_1 _11034_ (.B2(net78),
    .C1(_05004_),
    .B1(_05000_),
    .A1(_03920_),
    .Y(_00555_),
    .A2(net44));
 sg13g2_nand3_1 _11035_ (.B(_02883_),
    .C(net71),
    .A(_04978_),
    .Y(_05005_));
 sg13g2_o21ai_1 _11036_ (.B1(_05005_),
    .Y(_05006_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .A2(net71));
 sg13g2_mux2_1 _11037_ (.A0(_03234_),
    .A1(_03937_),
    .S(net188),
    .X(_05007_));
 sg13g2_o21ai_1 _11038_ (.B1(net243),
    .Y(_05008_),
    .A1(net78),
    .A2(_05007_));
 sg13g2_a221oi_1 _11039_ (.B2(_05002_),
    .C1(_05008_),
    .B1(_05006_),
    .A1(_02882_),
    .Y(_00556_),
    .A2(net44));
 sg13g2_nand2_1 _11040_ (.Y(_05009_),
    .A(_01770_),
    .B(net75));
 sg13g2_buf_2 _11041_ (.A(_05009_),
    .X(_05010_));
 sg13g2_buf_1 _11042_ (.A(_05010_),
    .X(_05011_));
 sg13g2_nor2_1 _11043_ (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .B(_04998_),
    .Y(_05012_));
 sg13g2_a21oi_1 _11044_ (.A1(_02970_),
    .A2(_04998_),
    .Y(_05013_),
    .B1(_05012_));
 sg13g2_nand2_1 _11045_ (.Y(_05014_),
    .A(net176),
    .B(_03235_));
 sg13g2_xnor2_1 _11046_ (.Y(_05015_),
    .A(net258),
    .B(_03950_));
 sg13g2_nand2_1 _11047_ (.Y(_05016_),
    .A(_04992_),
    .B(_05015_));
 sg13g2_a21oi_1 _11048_ (.A1(_05014_),
    .A2(_05016_),
    .Y(_05017_),
    .B1(_04987_));
 sg13g2_a21oi_1 _11049_ (.A1(_05002_),
    .A2(_05013_),
    .Y(_05018_),
    .B1(_05017_));
 sg13g2_o21ai_1 _11050_ (.B1(net243),
    .Y(_05019_),
    .A1(_02626_),
    .A2(_05011_));
 sg13g2_a21oi_1 _11051_ (.A1(net43),
    .A2(_05018_),
    .Y(_00557_),
    .B1(_05019_));
 sg13g2_nand2_1 _11052_ (.Y(_05020_),
    .A(net188),
    .B(_03969_));
 sg13g2_a21oi_1 _11053_ (.A1(net189),
    .A2(_03236_),
    .Y(_05021_),
    .B1(net84));
 sg13g2_buf_1 _11054_ (.A(net77),
    .X(_05022_));
 sg13g2_nand2_1 _11055_ (.Y(_05023_),
    .A(_02632_),
    .B(net77));
 sg13g2_o21ai_1 _11056_ (.B1(_05023_),
    .Y(_05024_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .A2(net70));
 sg13g2_a221oi_1 _11057_ (.B2(net81),
    .C1(_04980_),
    .B1(_05024_),
    .A1(_05020_),
    .Y(_05025_),
    .A2(_05021_));
 sg13g2_a21oi_1 _11058_ (.A1(net295),
    .A2(net44),
    .Y(_05026_),
    .B1(_05025_));
 sg13g2_nor2_1 _11059_ (.A(_04950_),
    .B(_05026_),
    .Y(_00558_));
 sg13g2_or3_1 _11060_ (.A(net83),
    .B(_02837_),
    .C(net67),
    .X(_05027_));
 sg13g2_o21ai_1 _11061_ (.B1(_05027_),
    .Y(_05028_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .A2(net71));
 sg13g2_a21oi_1 _11062_ (.A1(net176),
    .A2(_03237_),
    .Y(_05029_),
    .B1(_04987_));
 sg13g2_xnor2_1 _11063_ (.Y(_05030_),
    .A(net324),
    .B(_03982_));
 sg13g2_nand2_1 _11064_ (.Y(_05031_),
    .A(net175),
    .B(_05030_));
 sg13g2_o21ai_1 _11065_ (.B1(net243),
    .Y(_05032_),
    .A1(_01062_),
    .A2(_05010_));
 sg13g2_a221oi_1 _11066_ (.B2(_05031_),
    .C1(_05032_),
    .B1(_05029_),
    .A1(net78),
    .Y(_00559_),
    .A2(_05028_));
 sg13g2_nor2_1 _11067_ (.A(_01017_),
    .B(_05011_),
    .Y(_05033_));
 sg13g2_mux2_1 _11068_ (.A0(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .A1(_02889_),
    .S(_05022_),
    .X(_05034_));
 sg13g2_nor2_1 _11069_ (.A(net176),
    .B(_03994_),
    .Y(_05035_));
 sg13g2_nor2_1 _11070_ (.A(net188),
    .B(_03239_),
    .Y(_05036_));
 sg13g2_nor3_1 _11071_ (.A(net81),
    .B(_05035_),
    .C(_05036_),
    .Y(_05037_));
 sg13g2_a221oi_1 _11072_ (.B2(net82),
    .C1(_05037_),
    .B1(_05034_),
    .A1(net83),
    .Y(_05038_),
    .A2(net75));
 sg13g2_nor3_1 _11073_ (.A(net225),
    .B(_05033_),
    .C(_05038_),
    .Y(_00560_));
 sg13g2_nor2_1 _11074_ (.A(_00836_),
    .B(net43),
    .Y(_05039_));
 sg13g2_mux2_1 _11075_ (.A0(_03240_),
    .A1(_04018_),
    .S(_04992_),
    .X(_05040_));
 sg13g2_nor2_1 _11076_ (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .B(net77),
    .Y(_05041_));
 sg13g2_a21oi_1 _11077_ (.A1(_02973_),
    .A2(net70),
    .Y(_05042_),
    .B1(_05041_));
 sg13g2_mux2_1 _11078_ (.A0(_05040_),
    .A1(_05042_),
    .S(net81),
    .X(_05043_));
 sg13g2_nor2_1 _11079_ (.A(net44),
    .B(_05043_),
    .Y(_05044_));
 sg13g2_nor3_1 _11080_ (.A(net225),
    .B(_05039_),
    .C(_05044_),
    .Y(_00561_));
 sg13g2_mux2_1 _11081_ (.A0(_03242_),
    .A1(_04041_),
    .S(net175),
    .X(_05045_));
 sg13g2_nor2_1 _11082_ (.A(net78),
    .B(_05045_),
    .Y(_05046_));
 sg13g2_mux2_1 _11083_ (.A0(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .A1(_02638_),
    .S(net70),
    .X(_05047_));
 sg13g2_nor4_1 _11084_ (.A(net146),
    .B(net86),
    .C(_04980_),
    .D(_05047_),
    .Y(_05048_));
 sg13g2_o21ai_1 _11085_ (.B1(_04372_),
    .Y(_05049_),
    .A1(_01175_),
    .A2(_05010_));
 sg13g2_nor3_1 _11086_ (.A(_05046_),
    .B(_05048_),
    .C(_05049_),
    .Y(_00562_));
 sg13g2_xor2_1 _11087_ (.B(_04065_),
    .A(net323),
    .X(_05050_));
 sg13g2_nor2_1 _11088_ (.A(net176),
    .B(_05050_),
    .Y(_05051_));
 sg13g2_a21oi_1 _11089_ (.A1(net176),
    .A2(_03243_),
    .Y(_05052_),
    .B1(_05051_));
 sg13g2_nand3_1 _11090_ (.B(_02833_),
    .C(net70),
    .A(_04978_),
    .Y(_05053_));
 sg13g2_o21ai_1 _11091_ (.B1(_05053_),
    .Y(_05054_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .A2(net71));
 sg13g2_mux2_1 _11092_ (.A0(_05052_),
    .A1(_05054_),
    .S(net82),
    .X(_05055_));
 sg13g2_o21ai_1 _11093_ (.B1(net251),
    .Y(_05056_),
    .A1(net323),
    .A2(net43));
 sg13g2_nor2_1 _11094_ (.A(_05055_),
    .B(_05056_),
    .Y(_00563_));
 sg13g2_inv_1 _11095_ (.Y(_05057_),
    .A(_01030_));
 sg13g2_nand2_1 _11096_ (.Y(_05058_),
    .A(net189),
    .B(_03244_));
 sg13g2_nand3_1 _11097_ (.B(_02887_),
    .C(net77),
    .A(_04978_),
    .Y(_05059_));
 sg13g2_or2_1 _11098_ (.X(_05060_),
    .B(_04599_),
    .A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_nand3_1 _11099_ (.B(_05059_),
    .C(_05060_),
    .A(net84),
    .Y(_05061_));
 sg13g2_o21ai_1 _11100_ (.B1(_05061_),
    .Y(_05062_),
    .A1(net84),
    .A2(_05058_));
 sg13g2_o21ai_1 _11101_ (.B1(_05010_),
    .Y(_05063_),
    .A1(_04075_),
    .A2(_05062_));
 sg13g2_nand2b_1 _11102_ (.Y(_05064_),
    .B(net70),
    .A_N(_02887_));
 sg13g2_a221oi_1 _11103_ (.B2(net81),
    .C1(net176),
    .B1(_05064_),
    .A1(_01030_),
    .Y(_05065_),
    .A2(_04075_));
 sg13g2_o21ai_1 _11104_ (.B1(_04372_),
    .Y(_05066_),
    .A1(_05062_),
    .A2(_05065_));
 sg13g2_a21oi_1 _11105_ (.A1(_05057_),
    .A2(_05063_),
    .Y(_00564_),
    .B1(_05066_));
 sg13g2_nand2_1 _11106_ (.Y(_05067_),
    .A(_01179_),
    .B(net44));
 sg13g2_nor2_1 _11107_ (.A(net188),
    .B(_03249_),
    .Y(_05068_));
 sg13g2_a21oi_1 _11108_ (.A1(net188),
    .A2(_04112_),
    .Y(_05069_),
    .B1(_05068_));
 sg13g2_nand3_1 _11109_ (.B(_01527_),
    .C(_01663_),
    .A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Y(_05070_));
 sg13g2_o21ai_1 _11110_ (.B1(_05070_),
    .Y(_05071_),
    .A1(_02606_),
    .A2(_04983_));
 sg13g2_mux2_1 _11111_ (.A0(_05069_),
    .A1(_05071_),
    .S(_05001_),
    .X(_05072_));
 sg13g2_nand2_1 _11112_ (.Y(_05073_),
    .A(net43),
    .B(_05072_));
 sg13g2_a21oi_1 _11113_ (.A1(_05067_),
    .A2(_05073_),
    .Y(_00565_),
    .B1(net205));
 sg13g2_nor3_1 _11114_ (.A(net176),
    .B(net82),
    .C(_04085_),
    .Y(_05074_));
 sg13g2_nor2_1 _11115_ (.A(net175),
    .B(_03245_),
    .Y(_05075_));
 sg13g2_nand3b_1 _11116_ (.B(net70),
    .C(_04978_),
    .Y(_05076_),
    .A_N(_02976_));
 sg13g2_o21ai_1 _11117_ (.B1(_05076_),
    .Y(_05077_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .A2(net71));
 sg13g2_mux2_1 _11118_ (.A0(_05075_),
    .A1(_05077_),
    .S(net82),
    .X(_05078_));
 sg13g2_o21ai_1 _11119_ (.B1(net243),
    .Y(_05079_),
    .A1(\i_tinyqv.cpu.instr_data_start[23] ),
    .A2(_05010_));
 sg13g2_nor3_1 _11120_ (.A(_05074_),
    .B(_05078_),
    .C(_05079_),
    .Y(_00566_));
 sg13g2_nor2_1 _11121_ (.A(net175),
    .B(_03250_),
    .Y(_05080_));
 sg13g2_a21oi_1 _11122_ (.A1(net175),
    .A2(_04120_),
    .Y(_05081_),
    .B1(_05080_));
 sg13g2_o21ai_1 _11123_ (.B1(_05081_),
    .Y(_05082_),
    .A1(net146),
    .A2(net86));
 sg13g2_nor3_1 _11124_ (.A(net83),
    .B(_02819_),
    .C(net67),
    .Y(_05083_));
 sg13g2_a21o_1 _11125_ (.A2(net67),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .B1(_05083_),
    .X(_05084_));
 sg13g2_a22oi_1 _11126_ (.Y(_05085_),
    .B1(_05084_),
    .B2(net78),
    .A2(net44),
    .A1(net296));
 sg13g2_a21oi_1 _11127_ (.A1(_05082_),
    .A2(_05085_),
    .Y(_00567_),
    .B1(_04931_));
 sg13g2_nor2_1 _11128_ (.A(_04993_),
    .B(_03252_),
    .Y(_05086_));
 sg13g2_a21oi_1 _11129_ (.A1(net175),
    .A2(_04129_),
    .Y(_05087_),
    .B1(_05086_));
 sg13g2_o21ai_1 _11130_ (.B1(_05087_),
    .Y(_05088_),
    .A1(_01555_),
    .A2(_01563_));
 sg13g2_nor3_1 _11131_ (.A(net83),
    .B(_02879_),
    .C(net67),
    .Y(_05089_));
 sg13g2_a21o_1 _11132_ (.A2(net67),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .B1(_05089_),
    .X(_05090_));
 sg13g2_a22oi_1 _11133_ (.Y(_05091_),
    .B1(_05090_),
    .B2(net78),
    .A2(_04980_),
    .A1(_02612_));
 sg13g2_a21oi_1 _11134_ (.A1(_05088_),
    .A2(_05091_),
    .Y(_00568_),
    .B1(net205));
 sg13g2_mux2_1 _11135_ (.A0(_03253_),
    .A1(_04140_),
    .S(net175),
    .X(_05092_));
 sg13g2_o21ai_1 _11136_ (.B1(_05092_),
    .Y(_05093_),
    .A1(_01555_),
    .A2(_01563_));
 sg13g2_nor3_1 _11137_ (.A(net83),
    .B(_02968_),
    .C(_04983_),
    .Y(_05094_));
 sg13g2_a21o_1 _11138_ (.A2(net67),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .B1(_05094_),
    .X(_05095_));
 sg13g2_a22oi_1 _11139_ (.Y(_05096_),
    .B1(_05095_),
    .B2(net78),
    .A2(_04980_),
    .A1(net261));
 sg13g2_a21oi_1 _11140_ (.A1(_05093_),
    .A2(_05096_),
    .Y(_00569_),
    .B1(_04891_));
 sg13g2_nor2_1 _11141_ (.A(net259),
    .B(net43),
    .Y(_05097_));
 sg13g2_mux2_1 _11142_ (.A0(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .A1(_02623_),
    .S(net70),
    .X(_05098_));
 sg13g2_nor2_1 _11143_ (.A(_04988_),
    .B(_04149_),
    .Y(_05099_));
 sg13g2_a21oi_1 _11144_ (.A1(_04989_),
    .A2(_03254_),
    .Y(_05100_),
    .B1(_05099_));
 sg13g2_nor2_1 _11145_ (.A(net81),
    .B(_05100_),
    .Y(_05101_));
 sg13g2_a221oi_1 _11146_ (.B2(net82),
    .C1(_05101_),
    .B1(_05098_),
    .A1(_04984_),
    .Y(_05102_),
    .A2(net75));
 sg13g2_nor3_1 _11147_ (.A(net225),
    .B(_05097_),
    .C(_05102_),
    .Y(_00570_));
 sg13g2_and2_1 _11148_ (.A(_01559_),
    .B(_03255_),
    .X(_05103_));
 sg13g2_a21oi_1 _11149_ (.A1(net188),
    .A2(_04159_),
    .Y(_05104_),
    .B1(_05103_));
 sg13g2_inv_1 _11150_ (.Y(_05105_),
    .A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_mux2_1 _11151_ (.A0(_05105_),
    .A1(_02817_),
    .S(net77),
    .X(_05106_));
 sg13g2_mux2_1 _11152_ (.A0(_05104_),
    .A1(_05106_),
    .S(_03650_),
    .X(_05107_));
 sg13g2_nor2_1 _11153_ (.A(_04980_),
    .B(_05107_),
    .Y(_05108_));
 sg13g2_a21oi_1 _11154_ (.A1(_01065_),
    .A2(_04997_),
    .Y(_05109_),
    .B1(_05108_));
 sg13g2_nor2_1 _11155_ (.A(net204),
    .B(_05109_),
    .Y(_00571_));
 sg13g2_nor2_1 _11156_ (.A(net325),
    .B(net43),
    .Y(_05110_));
 sg13g2_nor2_1 _11157_ (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .B(net70),
    .Y(_05111_));
 sg13g2_a21oi_1 _11158_ (.A1(_02881_),
    .A2(net71),
    .Y(_05112_),
    .B1(_05111_));
 sg13g2_nor2_1 _11159_ (.A(net189),
    .B(_03854_),
    .Y(_05113_));
 sg13g2_a21oi_1 _11160_ (.A1(_04989_),
    .A2(_03229_),
    .Y(_05114_),
    .B1(_05113_));
 sg13g2_nor2_1 _11161_ (.A(net81),
    .B(_05114_),
    .Y(_05115_));
 sg13g2_a221oi_1 _11162_ (.B2(net82),
    .C1(_05115_),
    .B1(_05112_),
    .A1(_04984_),
    .Y(_05116_),
    .A2(_03652_));
 sg13g2_nor3_1 _11163_ (.A(_04938_),
    .B(_05110_),
    .C(_05116_),
    .Y(_00572_));
 sg13g2_nand2_1 _11164_ (.Y(_05117_),
    .A(net262),
    .B(net44));
 sg13g2_nor2_1 _11165_ (.A(net189),
    .B(_03875_),
    .Y(_05118_));
 sg13g2_a21oi_1 _11166_ (.A1(net189),
    .A2(_03231_),
    .Y(_05119_),
    .B1(_05118_));
 sg13g2_nand2_1 _11167_ (.Y(_05120_),
    .A(_02969_),
    .B(_05022_));
 sg13g2_or2_1 _11168_ (.X(_05121_),
    .B(net77),
    .A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_nand3_1 _11169_ (.B(_05120_),
    .C(_05121_),
    .A(_03650_),
    .Y(_05122_));
 sg13g2_o21ai_1 _11170_ (.B1(_05122_),
    .Y(_05123_),
    .A1(net81),
    .A2(_05119_));
 sg13g2_nand2_1 _11171_ (.Y(_05124_),
    .A(net43),
    .B(_05123_));
 sg13g2_a21oi_1 _11172_ (.A1(_05117_),
    .A2(_05124_),
    .Y(_00573_),
    .B1(_04891_));
 sg13g2_nor2_1 _11173_ (.A(net297),
    .B(net43),
    .Y(_05125_));
 sg13g2_nand2_1 _11174_ (.Y(_05126_),
    .A(net189),
    .B(_03232_));
 sg13g2_o21ai_1 _11175_ (.B1(_05126_),
    .Y(_05127_),
    .A1(net189),
    .A2(_03888_));
 sg13g2_mux2_1 _11176_ (.A0(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .A1(_02618_),
    .S(net77),
    .X(_05128_));
 sg13g2_mux2_1 _11177_ (.A0(_05127_),
    .A1(_05128_),
    .S(_05001_),
    .X(_05129_));
 sg13g2_nor2_1 _11178_ (.A(_04997_),
    .B(_05129_),
    .Y(_05130_));
 sg13g2_nor3_1 _11179_ (.A(_04938_),
    .B(_05125_),
    .C(_05130_),
    .Y(_00574_));
 sg13g2_nand2_1 _11180_ (.Y(_05131_),
    .A(_01539_),
    .B(_01663_));
 sg13g2_and2_1 _11181_ (.A(net75),
    .B(_05131_),
    .X(_05132_));
 sg13g2_nor3_1 _11182_ (.A(\i_tinyqv.cpu.instr_fetch_started ),
    .B(\i_tinyqv.cpu.instr_fetch_stopped ),
    .C(\i_tinyqv.cpu.instr_fetch_running ),
    .Y(_05133_));
 sg13g2_o21ai_1 _11183_ (.B1(net227),
    .Y(_05134_),
    .A1(net146),
    .A2(net86));
 sg13g2_inv_1 _11184_ (.Y(_05135_),
    .A(\i_tinyqv.cpu.instr_fetch_stopped ));
 sg13g2_o21ai_1 _11185_ (.B1(_05132_),
    .Y(_05136_),
    .A1(\i_tinyqv.cpu.instr_fetch_started ),
    .A2(_05135_));
 sg13g2_a221oi_1 _11186_ (.B2(_05136_),
    .C1(net207),
    .B1(_05134_),
    .A1(_05132_),
    .Y(_00575_),
    .A2(_05133_));
 sg13g2_inv_1 _11187_ (.Y(_05137_),
    .A(_01429_));
 sg13g2_buf_1 _11188_ (.A(_03125_),
    .X(_05138_));
 sg13g2_o21ai_1 _11189_ (.B1(net243),
    .Y(_05139_),
    .A1(_03529_),
    .A2(_03125_));
 sg13g2_a21oi_1 _11190_ (.A1(_05137_),
    .A2(net57),
    .Y(_00576_),
    .B1(_05139_));
 sg13g2_a21o_1 _11191_ (.A2(_05138_),
    .A1(_01431_),
    .B1(_05139_),
    .X(_00577_));
 sg13g2_nor2_1 _11192_ (.A(_01295_),
    .B(_01386_),
    .Y(_05140_));
 sg13g2_nor2_1 _11193_ (.A(_05140_),
    .B(_03118_),
    .Y(_05141_));
 sg13g2_o21ai_1 _11194_ (.B1(net233),
    .Y(_05142_),
    .A1(_03696_),
    .A2(_05141_));
 sg13g2_or4_1 _11195_ (.A(net146),
    .B(net86),
    .C(_01527_),
    .D(_03125_),
    .X(_05143_));
 sg13g2_a21oi_1 _11196_ (.A1(_05142_),
    .A2(_05143_),
    .Y(_00578_),
    .B1(net207));
 sg13g2_nor2_1 _11197_ (.A(_01559_),
    .B(_04027_),
    .Y(_05144_));
 sg13g2_a21oi_1 _11198_ (.A1(_04988_),
    .A2(_03241_),
    .Y(_05145_),
    .B1(_05144_));
 sg13g2_nand2_1 _11199_ (.Y(_05146_),
    .A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .B(_04982_));
 sg13g2_o21ai_1 _11200_ (.B1(_05146_),
    .Y(_05147_),
    .A1(net84),
    .A2(_05145_));
 sg13g2_a21oi_1 _11201_ (.A1(_01614_),
    .A2(net75),
    .Y(_05148_),
    .B1(_05147_));
 sg13g2_nor2_1 _11202_ (.A(net204),
    .B(_05148_),
    .Y(_00579_));
 sg13g2_mux2_1 _11203_ (.A0(_03246_),
    .A1(_04095_),
    .S(net188),
    .X(_05149_));
 sg13g2_o21ai_1 _11204_ (.B1(_05149_),
    .Y(_05150_),
    .A1(net146),
    .A2(net86));
 sg13g2_nand2_1 _11205_ (.Y(_05151_),
    .A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .B(net67));
 sg13g2_and2_1 _11206_ (.A(_05150_),
    .B(_05151_),
    .X(_05152_));
 sg13g2_xnor2_1 _11207_ (.Y(_05153_),
    .A(_00160_),
    .B(_01611_));
 sg13g2_nand2_1 _11208_ (.Y(_05154_),
    .A(net75),
    .B(_05153_));
 sg13g2_a21oi_1 _11209_ (.A1(_05152_),
    .A2(_05154_),
    .Y(_00580_),
    .B1(net207));
 sg13g2_nand2_1 _11210_ (.Y(_05155_),
    .A(_03713_),
    .B(_03118_));
 sg13g2_a22oi_1 _11211_ (.Y(_05156_),
    .B1(_05155_),
    .B2(_04956_),
    .A2(_03713_),
    .A1(_05140_));
 sg13g2_nor2_1 _11212_ (.A(net205),
    .B(_05156_),
    .Y(_00582_));
 sg13g2_nor2b_1 _11213_ (.A(\i_tinyqv.cpu.is_alu_imm ),
    .B_N(net58),
    .Y(_05157_));
 sg13g2_nor2_1 _11214_ (.A(net100),
    .B(_03143_),
    .Y(_05158_));
 sg13g2_a21oi_1 _11215_ (.A1(net94),
    .A2(_03351_),
    .Y(_05159_),
    .B1(net110));
 sg13g2_nor3_1 _11216_ (.A(net94),
    .B(_03370_),
    .C(_03201_),
    .Y(_05160_));
 sg13g2_o21ai_1 _11217_ (.B1(_03136_),
    .Y(_05161_),
    .A1(_05159_),
    .A2(_05160_));
 sg13g2_nand2b_1 _11218_ (.Y(_05162_),
    .B(_05161_),
    .A_N(_03392_));
 sg13g2_a221oi_1 _11219_ (.B2(net91),
    .C1(net57),
    .B1(_05162_),
    .A1(_03199_),
    .Y(_05163_),
    .A2(_05158_));
 sg13g2_nor3_1 _11220_ (.A(net225),
    .B(_05157_),
    .C(_05163_),
    .Y(_00583_));
 sg13g2_nor2_1 _11221_ (.A(net122),
    .B(net155),
    .Y(_05164_));
 sg13g2_nor3_1 _11222_ (.A(net95),
    .B(_03179_),
    .C(_03728_),
    .Y(_05165_));
 sg13g2_a221oi_1 _11223_ (.B2(_05164_),
    .C1(_05165_),
    .B1(_05158_),
    .A1(_03206_),
    .Y(_05166_),
    .A2(_03201_));
 sg13g2_nor2_1 _11224_ (.A(_04909_),
    .B(_05166_),
    .Y(_05167_));
 sg13g2_a21oi_1 _11225_ (.A1(_00894_),
    .A2(net57),
    .Y(_05168_),
    .B1(_05167_));
 sg13g2_nor2_1 _11226_ (.A(net205),
    .B(_05168_),
    .Y(_00584_));
 sg13g2_nor4_1 _11227_ (.A(_01471_),
    .B(net91),
    .C(_03125_),
    .D(_03159_),
    .Y(_05169_));
 sg13g2_a21oi_1 _11228_ (.A1(\i_tinyqv.cpu.is_auipc ),
    .A2(_05138_),
    .Y(_05170_),
    .B1(_05169_));
 sg13g2_nor2_1 _11229_ (.A(net205),
    .B(_05170_),
    .Y(_00585_));
 sg13g2_nor2b_1 _11230_ (.A(_00893_),
    .B_N(net58),
    .Y(_05171_));
 sg13g2_o21ai_1 _11231_ (.B1(_03770_),
    .Y(_05172_),
    .A1(net91),
    .A2(_03175_));
 sg13g2_nor2_1 _11232_ (.A(net57),
    .B(_05172_),
    .Y(_05173_));
 sg13g2_nor3_1 _11233_ (.A(net225),
    .B(_05171_),
    .C(_05173_),
    .Y(_00586_));
 sg13g2_mux2_1 _11234_ (.A0(_01539_),
    .A1(\i_tinyqv.cpu.is_jal ),
    .S(_03125_),
    .X(_05174_));
 sg13g2_and2_1 _11235_ (.A(net251),
    .B(_05174_),
    .X(_00587_));
 sg13g2_nor2b_1 _11236_ (.A(\i_tinyqv.cpu.is_jalr ),
    .B_N(net58),
    .Y(_05175_));
 sg13g2_inv_1 _11237_ (.Y(_05176_),
    .A(_01500_));
 sg13g2_nor2_1 _11238_ (.A(net171),
    .B(net91),
    .Y(_05177_));
 sg13g2_a221oi_1 _11239_ (.B2(_01534_),
    .C1(net57),
    .B1(_05177_),
    .A1(_05176_),
    .Y(_05178_),
    .A2(_03373_));
 sg13g2_nor3_1 _11240_ (.A(net226),
    .B(_05175_),
    .C(_05178_),
    .Y(_00588_));
 sg13g2_nand4_1 _11241_ (.B(net105),
    .C(_03351_),
    .A(_01462_),
    .Y(_05179_),
    .D(_03163_));
 sg13g2_nor2_1 _11242_ (.A(net106),
    .B(_03533_),
    .Y(_05180_));
 sg13g2_o21ai_1 _11243_ (.B1(net95),
    .Y(_05181_),
    .A1(_03679_),
    .A2(_05180_));
 sg13g2_a21oi_1 _11244_ (.A1(_05179_),
    .A2(_05181_),
    .Y(_05182_),
    .B1(net92));
 sg13g2_a21oi_1 _11245_ (.A1(_01484_),
    .A2(net92),
    .Y(_05183_),
    .B1(_05182_));
 sg13g2_nor2_1 _11246_ (.A(net58),
    .B(_05183_),
    .Y(_05184_));
 sg13g2_a21oi_1 _11247_ (.A1(_01203_),
    .A2(net57),
    .Y(_05185_),
    .B1(_05184_));
 sg13g2_nor2_1 _11248_ (.A(net205),
    .B(_05185_),
    .Y(_00589_));
 sg13g2_nor2b_1 _11249_ (.A(\i_tinyqv.cpu.is_lui ),
    .B_N(net58),
    .Y(_05186_));
 sg13g2_nor4_1 _11250_ (.A(net122),
    .B(_03130_),
    .C(_03129_),
    .D(_03159_),
    .Y(_05187_));
 sg13g2_nor3_1 _11251_ (.A(net58),
    .B(_03427_),
    .C(_05187_),
    .Y(_05188_));
 sg13g2_nor3_1 _11252_ (.A(net226),
    .B(_05186_),
    .C(_05188_),
    .Y(_00590_));
 sg13g2_and2_1 _11253_ (.A(_01769_),
    .B(_04909_),
    .X(_05189_));
 sg13g2_nand2b_1 _11254_ (.Y(_05190_),
    .B(net96),
    .A_N(_03163_));
 sg13g2_o21ai_1 _11255_ (.B1(_03208_),
    .Y(_05191_),
    .A1(_03203_),
    .A2(_05190_));
 sg13g2_a221oi_1 _11256_ (.B2(net97),
    .C1(net57),
    .B1(_05191_),
    .A1(net92),
    .Y(_05192_),
    .A2(_03357_));
 sg13g2_nor3_1 _11257_ (.A(net226),
    .B(_05189_),
    .C(_05192_),
    .Y(_00591_));
 sg13g2_nor2b_1 _11258_ (.A(_01219_),
    .B_N(net58),
    .Y(_05193_));
 sg13g2_and2_1 _11259_ (.A(_03208_),
    .B(_03750_),
    .X(_05194_));
 sg13g2_a22oi_1 _11260_ (.Y(_05195_),
    .B1(_05194_),
    .B2(net97),
    .A2(_05158_),
    .A1(_03138_));
 sg13g2_o21ai_1 _11261_ (.B1(_05195_),
    .Y(_05196_),
    .A1(_01500_),
    .A2(_03373_));
 sg13g2_nor2_1 _11262_ (.A(net57),
    .B(_05196_),
    .Y(_05197_));
 sg13g2_nor3_1 _11263_ (.A(net226),
    .B(_05193_),
    .C(_05197_),
    .Y(_00592_));
 sg13g2_inv_1 _11264_ (.Y(_05198_),
    .A(\i_tinyqv.cpu.load_started ));
 sg13g2_a21oi_1 _11265_ (.A1(_05198_),
    .A2(net118),
    .Y(_00593_),
    .B1(_01771_));
 sg13g2_a21oi_1 _11266_ (.A1(_01306_),
    .A2(_01301_),
    .Y(_05199_),
    .B1(_01360_));
 sg13g2_nand2_1 _11267_ (.Y(_05200_),
    .A(_01213_),
    .B(_04923_));
 sg13g2_a21oi_1 _11268_ (.A1(\i_tinyqv.cpu.no_write_in_progress ),
    .A2(_01590_),
    .Y(_05201_),
    .B1(net226));
 sg13g2_o21ai_1 _11269_ (.B1(_05201_),
    .Y(_00598_),
    .A1(_05199_),
    .A2(_05200_));
 sg13g2_o21ai_1 _11270_ (.B1(_05010_),
    .Y(_05202_),
    .A1(_01429_),
    .A2(_05147_));
 sg13g2_nor2_1 _11271_ (.A(net83),
    .B(_01430_),
    .Y(_05203_));
 sg13g2_nor2_1 _11272_ (.A(_04600_),
    .B(_05203_),
    .Y(_05204_));
 sg13g2_o21ai_1 _11273_ (.B1(net243),
    .Y(_05205_),
    .A1(_05147_),
    .A2(_05204_));
 sg13g2_a21oi_1 _11274_ (.A1(_01068_),
    .A2(_05202_),
    .Y(_00599_),
    .B1(_05205_));
 sg13g2_o21ai_1 _11275_ (.B1(net75),
    .Y(_05206_),
    .A1(net83),
    .A2(_01433_));
 sg13g2_a221oi_1 _11276_ (.B2(_05206_),
    .C1(net207),
    .B1(_05152_),
    .A1(_01027_),
    .Y(_00600_),
    .A2(net44));
 sg13g2_nand2_1 _11277_ (.Y(_05207_),
    .A(net227),
    .B(_01590_));
 sg13g2_a21oi_1 _11278_ (.A1(_05131_),
    .A2(_05207_),
    .Y(_00613_),
    .B1(net207));
 sg13g2_nand3b_1 _11279_ (.B(_03794_),
    .C(_04304_),
    .Y(_05208_),
    .A_N(net162));
 sg13g2_mux2_1 _11280_ (.A0(_01305_),
    .A1(_02531_),
    .S(net318),
    .X(_05209_));
 sg13g2_a22oi_1 _11281_ (.Y(_05210_),
    .B1(_05209_),
    .B2(net322),
    .A2(_04304_),
    .A1(_02524_));
 sg13g2_o21ai_1 _11282_ (.B1(_01354_),
    .Y(_05211_),
    .A1(_01297_),
    .A2(_05210_));
 sg13g2_a21oi_1 _11283_ (.A1(_04261_),
    .A2(_05208_),
    .Y(_05212_),
    .B1(_05211_));
 sg13g2_nor2b_1 _11284_ (.A(_05212_),
    .B_N(debug_data_continue),
    .Y(_00614_));
 sg13g2_nor2_1 _11285_ (.A(net209),
    .B(_03863_),
    .Y(_00616_));
 sg13g2_and2_1 _11286_ (.A(net232),
    .B(_04601_),
    .X(_00617_));
 sg13g2_nand4_1 _11287_ (.B(net193),
    .C(_04275_),
    .A(_04266_),
    .Y(_05213_),
    .D(_04283_));
 sg13g2_nor2b_1 _11288_ (.A(_04264_),
    .B_N(_05213_),
    .Y(_05214_));
 sg13g2_nor2_1 _11289_ (.A(_04260_),
    .B(_05214_),
    .Y(_00650_));
 sg13g2_nand2b_1 _11290_ (.Y(_00659_),
    .B(net208),
    .A_N(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ));
 sg13g2_nand2b_1 _11291_ (.Y(_00660_),
    .B(net208),
    .A_N(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ));
 sg13g2_nor3_1 _11292_ (.A(_04192_),
    .B(_03808_),
    .C(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .Y(_05215_));
 sg13g2_and2_1 _11293_ (.A(_00617_),
    .B(_05215_),
    .X(_00680_));
 sg13g2_inv_1 _11294_ (.Y(_05216_),
    .A(_04345_));
 sg13g2_and4_1 _11295_ (.A(_05216_),
    .B(_04346_),
    .C(_04351_),
    .D(_04352_),
    .X(_05217_));
 sg13g2_nor4_1 _11296_ (.A(\i_uart_rx.cycle_counter[3] ),
    .B(_04344_),
    .C(\i_uart_rx.cycle_counter[9] ),
    .D(_04744_),
    .Y(_05218_));
 sg13g2_nand3_1 _11297_ (.B(_05217_),
    .C(_05218_),
    .A(_04350_),
    .Y(_05219_));
 sg13g2_mux2_1 _11298_ (.A0(\i_uart_rx.rxd_reg[0] ),
    .A1(\i_uart_rx.bit_sample ),
    .S(_05219_),
    .X(_05220_));
 sg13g2_and2_1 _11299_ (.A(net213),
    .B(_05220_),
    .X(_00715_));
 sg13g2_a21oi_1 _11300_ (.A1(_01371_),
    .A2(_04721_),
    .Y(_05221_),
    .B1(_01368_));
 sg13g2_or2_1 _11301_ (.X(_05222_),
    .B(_05221_),
    .A(_04356_));
 sg13g2_buf_1 _11302_ (.A(_05222_),
    .X(_05223_));
 sg13g2_nand3_1 _11303_ (.B(_01351_),
    .C(net123),
    .A(_01350_),
    .Y(_05224_));
 sg13g2_and2_1 _11304_ (.A(_01374_),
    .B(_05224_),
    .X(_05225_));
 sg13g2_nor2_1 _11305_ (.A(net317),
    .B(\i_uart_rx.rxd_reg[0] ),
    .Y(_05226_));
 sg13g2_a22oi_1 _11306_ (.Y(_05227_),
    .B1(_04357_),
    .B2(_05226_),
    .A2(_00206_),
    .A1(net316));
 sg13g2_nor2_1 _11307_ (.A(net316),
    .B(_04720_),
    .Y(_05228_));
 sg13g2_o21ai_1 _11308_ (.B1(_00206_),
    .Y(_05229_),
    .A1(_01368_),
    .A2(_05228_));
 sg13g2_o21ai_1 _11309_ (.B1(_05229_),
    .Y(_05230_),
    .A1(net315),
    .A2(_05227_));
 sg13g2_nor4_1 _11310_ (.A(net317),
    .B(_00207_),
    .C(_01373_),
    .D(_05219_),
    .Y(_05231_));
 sg13g2_nor3_1 _11311_ (.A(_05225_),
    .B(_05230_),
    .C(_05231_),
    .Y(_05232_));
 sg13g2_o21ai_1 _11312_ (.B1(net231),
    .Y(_05233_),
    .A1(net317),
    .A2(_05223_));
 sg13g2_a21oi_1 _11313_ (.A1(_05223_),
    .A2(_05232_),
    .Y(_00727_),
    .B1(_05233_));
 sg13g2_o21ai_1 _11314_ (.B1(_05223_),
    .Y(_05234_),
    .A1(_01366_),
    .A2(_01372_));
 sg13g2_nor2_1 _11315_ (.A(net317),
    .B(_01373_),
    .Y(_05235_));
 sg13g2_nand4_1 _11316_ (.B(_04350_),
    .C(_05217_),
    .A(_00207_),
    .Y(_05236_),
    .D(_05218_));
 sg13g2_a21oi_1 _11317_ (.A1(_05235_),
    .A2(_05236_),
    .Y(_05237_),
    .B1(_05225_));
 sg13g2_o21ai_1 _11318_ (.B1(_05237_),
    .Y(_05238_),
    .A1(net316),
    .A2(_01367_));
 sg13g2_a22oi_1 _11319_ (.Y(_05239_),
    .B1(_05238_),
    .B2(_05223_),
    .A2(_05234_),
    .A1(_01369_));
 sg13g2_nor2_1 _11320_ (.A(net209),
    .B(_05239_),
    .Y(_00728_));
 sg13g2_nand3_1 _11321_ (.B(net317),
    .C(_04356_),
    .A(net316),
    .Y(_05240_));
 sg13g2_nor3_1 _11322_ (.A(_01368_),
    .B(net315),
    .C(_05240_),
    .Y(_05241_));
 sg13g2_a21oi_1 _11323_ (.A1(_01368_),
    .A2(_05240_),
    .Y(_05242_),
    .B1(_05241_));
 sg13g2_nor2_1 _11324_ (.A(net209),
    .B(_05242_),
    .Y(_00729_));
 sg13g2_inv_1 _11325_ (.Y(_05243_),
    .A(_04356_));
 sg13g2_o21ai_1 _11326_ (.B1(net315),
    .Y(_05244_),
    .A1(_01367_),
    .A2(_05243_));
 sg13g2_o21ai_1 _11327_ (.B1(_05244_),
    .Y(_05245_),
    .A1(net315),
    .A2(_05240_));
 sg13g2_a22oi_1 _11328_ (.Y(_05246_),
    .B1(_05245_),
    .B2(_01368_),
    .A2(_01370_),
    .A1(_04719_));
 sg13g2_a21oi_1 _11329_ (.A1(_05237_),
    .A2(_05246_),
    .Y(_00730_),
    .B1(net210));
 sg13g2_nand2b_1 _11330_ (.Y(_00739_),
    .B(net208),
    .A_N(\i_uart_rx.rxd_reg[1] ));
 sg13g2_nand2b_1 _11331_ (.Y(_00740_),
    .B(_04839_),
    .A_N(net7));
 sg13g2_nand3b_1 _11332_ (.B(_04839_),
    .C(_04357_),
    .Y(_00741_),
    .A_N(net315));
 sg13g2_nand3_1 _11333_ (.B(_03078_),
    .C(net123),
    .A(_01382_),
    .Y(_05247_));
 sg13g2_buf_1 _11334_ (.A(_05247_),
    .X(_05248_));
 sg13g2_inv_2 _11335_ (.Y(_05249_),
    .A(_05248_));
 sg13g2_nand2_1 _11336_ (.Y(_05250_),
    .A(net309),
    .B(_05249_));
 sg13g2_xnor2_1 _11337_ (.Y(_05251_),
    .A(_01379_),
    .B(_01377_));
 sg13g2_and2_1 _11338_ (.A(net190),
    .B(_05251_),
    .X(_05252_));
 sg13g2_buf_2 _11339_ (.A(_05252_),
    .X(_05253_));
 sg13g2_mux2_1 _11340_ (.A0(\i_uart_tx.data_to_send[0] ),
    .A1(\i_uart_tx.data_to_send[1] ),
    .S(_05253_),
    .X(_05254_));
 sg13g2_nand2_1 _11341_ (.Y(_05255_),
    .A(net93),
    .B(_05254_));
 sg13g2_a21oi_1 _11342_ (.A1(_05250_),
    .A2(_05255_),
    .Y(_00753_),
    .B1(net210));
 sg13g2_nand2_1 _11343_ (.Y(_05256_),
    .A(net308),
    .B(_05249_));
 sg13g2_mux2_1 _11344_ (.A0(\i_uart_tx.data_to_send[1] ),
    .A1(\i_uart_tx.data_to_send[2] ),
    .S(_05253_),
    .X(_05257_));
 sg13g2_nand2_1 _11345_ (.Y(_05258_),
    .A(net93),
    .B(_05257_));
 sg13g2_a21oi_1 _11346_ (.A1(_05256_),
    .A2(_05258_),
    .Y(_00754_),
    .B1(net210));
 sg13g2_nand2_1 _11347_ (.Y(_05259_),
    .A(_01721_),
    .B(_05249_));
 sg13g2_mux2_1 _11348_ (.A0(\i_uart_tx.data_to_send[2] ),
    .A1(\i_uart_tx.data_to_send[3] ),
    .S(_05253_),
    .X(_05260_));
 sg13g2_nand2_1 _11349_ (.Y(_05261_),
    .A(net93),
    .B(_05260_));
 sg13g2_a21oi_1 _11350_ (.A1(_05259_),
    .A2(_05261_),
    .Y(_00755_),
    .B1(net210));
 sg13g2_nand2_1 _11351_ (.Y(_05262_),
    .A(_01724_),
    .B(_05249_));
 sg13g2_mux2_1 _11352_ (.A0(\i_uart_tx.data_to_send[3] ),
    .A1(\i_uart_tx.data_to_send[4] ),
    .S(_05253_),
    .X(_05263_));
 sg13g2_nand2_1 _11353_ (.Y(_05264_),
    .A(net93),
    .B(_05263_));
 sg13g2_a21oi_1 _11354_ (.A1(_05262_),
    .A2(_05264_),
    .Y(_00756_),
    .B1(_04816_));
 sg13g2_nand2_1 _11355_ (.Y(_05265_),
    .A(_01727_),
    .B(_05249_));
 sg13g2_mux2_1 _11356_ (.A0(\i_uart_tx.data_to_send[4] ),
    .A1(\i_uart_tx.data_to_send[5] ),
    .S(_05253_),
    .X(_05266_));
 sg13g2_nand2_1 _11357_ (.Y(_05267_),
    .A(_05248_),
    .B(_05266_));
 sg13g2_a21oi_1 _11358_ (.A1(_05265_),
    .A2(_05267_),
    .Y(_00757_),
    .B1(_04816_));
 sg13g2_nand2_1 _11359_ (.Y(_05268_),
    .A(net305),
    .B(_05249_));
 sg13g2_mux2_1 _11360_ (.A0(\i_uart_tx.data_to_send[5] ),
    .A1(\i_uart_tx.data_to_send[6] ),
    .S(_05253_),
    .X(_05269_));
 sg13g2_nand2_1 _11361_ (.Y(_05270_),
    .A(net93),
    .B(_05269_));
 sg13g2_a21oi_1 _11362_ (.A1(_05268_),
    .A2(_05270_),
    .Y(_00758_),
    .B1(net210));
 sg13g2_nand2_1 _11363_ (.Y(_05271_),
    .A(net304),
    .B(_05249_));
 sg13g2_mux2_1 _11364_ (.A0(\i_uart_tx.data_to_send[6] ),
    .A1(\i_uart_tx.data_to_send[7] ),
    .S(_05253_),
    .X(_05272_));
 sg13g2_nand2_1 _11365_ (.Y(_05273_),
    .A(net93),
    .B(_05272_));
 sg13g2_a21oi_1 _11366_ (.A1(_05271_),
    .A2(_05273_),
    .Y(_00759_),
    .B1(net210));
 sg13g2_or2_1 _11367_ (.X(_05274_),
    .B(net93),
    .A(_00205_));
 sg13g2_nand3b_1 _11368_ (.B(\i_uart_tx.data_to_send[7] ),
    .C(net93),
    .Y(_05275_),
    .A_N(_05253_));
 sg13g2_a21oi_1 _11369_ (.A1(_05274_),
    .A2(_05275_),
    .Y(_00760_),
    .B1(_04794_));
 sg13g2_a21oi_1 _11370_ (.A1(_01379_),
    .A2(net190),
    .Y(_05276_),
    .B1(_05249_));
 sg13g2_inv_1 _11371_ (.Y(_05277_),
    .A(_01379_));
 sg13g2_a21oi_1 _11372_ (.A1(_01375_),
    .A2(_05277_),
    .Y(_05278_),
    .B1(_01376_));
 sg13g2_nand2b_1 _11373_ (.Y(_05279_),
    .B(net190),
    .A_N(_05278_));
 sg13g2_o21ai_1 _11374_ (.B1(_05279_),
    .Y(_05280_),
    .A1(_01375_),
    .A2(_05276_));
 sg13g2_nand2_1 _11375_ (.Y(_05281_),
    .A(_01378_),
    .B(net190));
 sg13g2_o21ai_1 _11376_ (.B1(_05281_),
    .Y(_05282_),
    .A1(_01378_),
    .A2(_05280_));
 sg13g2_nor2_1 _11377_ (.A(_04817_),
    .B(_05282_),
    .Y(_00761_));
 sg13g2_nor2_1 _11378_ (.A(_05277_),
    .B(_01376_),
    .Y(_05283_));
 sg13g2_o21ai_1 _11379_ (.B1(net190),
    .Y(_05284_),
    .A1(_01378_),
    .A2(_05283_));
 sg13g2_nor2_1 _11380_ (.A(_01375_),
    .B(_05281_),
    .Y(_05285_));
 sg13g2_a21oi_1 _11381_ (.A1(_01375_),
    .A2(_05284_),
    .Y(_05286_),
    .B1(_05285_));
 sg13g2_nor2_1 _11382_ (.A(_04795_),
    .B(_05286_),
    .Y(_00762_));
 sg13g2_nand3_1 _11383_ (.B(_01375_),
    .C(net190),
    .A(_01378_),
    .Y(_05287_));
 sg13g2_xor2_1 _11384_ (.B(_05287_),
    .A(_01376_),
    .X(_05288_));
 sg13g2_nor2_1 _11385_ (.A(_04795_),
    .B(_05288_),
    .Y(_00763_));
 sg13g2_nand2b_1 _11386_ (.Y(_05289_),
    .B(_01376_),
    .A_N(_01378_));
 sg13g2_nand3_1 _11387_ (.B(net190),
    .C(_05289_),
    .A(_01375_),
    .Y(_05290_));
 sg13g2_nand4_1 _11388_ (.B(_05277_),
    .C(_01376_),
    .A(_01375_),
    .Y(_05291_),
    .D(_04759_));
 sg13g2_nand2b_1 _11389_ (.Y(_05292_),
    .B(_05291_),
    .A_N(_05283_));
 sg13g2_a22oi_1 _11390_ (.Y(_05293_),
    .B1(_05292_),
    .B2(_01378_),
    .A2(_05290_),
    .A1(_01379_));
 sg13g2_nor2_1 _11391_ (.A(net211),
    .B(_05293_),
    .Y(_00764_));
 sg13g2_a21oi_1 _11392_ (.A1(_01379_),
    .A2(\i_uart_tx.data_to_send[0] ),
    .Y(_05294_),
    .B1(_01380_));
 sg13g2_nor3_1 _11393_ (.A(_01379_),
    .B(\i_uart_tx.data_to_send[0] ),
    .C(_01377_),
    .Y(_05295_));
 sg13g2_a21oi_1 _11394_ (.A1(_01377_),
    .A2(_05294_),
    .Y(_05296_),
    .B1(_05295_));
 sg13g2_nand2b_1 _11395_ (.Y(_00765_),
    .B(net208),
    .A_N(_05296_));
 sg13g2_and2_1 _11396_ (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .B(net1),
    .X(net17));
 sg13g2_nor2_1 _11397_ (.A(\gpio_out_sel[9] ),
    .B(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .Y(_05297_));
 sg13g2_a21oi_1 _11398_ (.A1(\gpio_out_sel[9] ),
    .A2(_01425_),
    .Y(uio_out7),
    .B1(_05297_));
 sg13g2_nand2_1 _11399_ (.Y(_05298_),
    .A(net245),
    .B(_04207_));
 sg13g2_nor3_1 _11400_ (.A(_04169_),
    .B(_01651_),
    .C(_05298_),
    .Y(_05299_));
 sg13g2_nand2_1 _11401_ (.Y(_05300_),
    .A(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .B(_03811_));
 sg13g2_o21ai_1 _11402_ (.B1(_05300_),
    .Y(_05301_),
    .A1(_03607_),
    .A2(_04179_));
 sg13g2_o21ai_1 _11403_ (.B1(_04287_),
    .Y(_05302_),
    .A1(net311),
    .A2(_04170_));
 sg13g2_o21ai_1 _11404_ (.B1(_04639_),
    .Y(_05303_),
    .A1(net246),
    .A2(_05302_));
 sg13g2_buf_1 _11405_ (.A(_05303_),
    .X(_05304_));
 sg13g2_o21ai_1 _11406_ (.B1(_05304_),
    .Y(_05305_),
    .A1(_05299_),
    .A2(_05301_));
 sg13g2_inv_1 _11407_ (.Y(net21),
    .A(_05305_));
 sg13g2_nand2_1 _11408_ (.Y(_05306_),
    .A(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .B(_04171_));
 sg13g2_o21ai_1 _11409_ (.B1(_05306_),
    .Y(_05307_),
    .A1(_04277_),
    .A2(_05298_));
 sg13g2_a22oi_1 _11410_ (.Y(_05308_),
    .B1(_05307_),
    .B2(_01650_),
    .A2(_04180_),
    .A1(_03665_));
 sg13g2_nand2_1 _11411_ (.Y(net22),
    .A(_05304_),
    .B(_05308_));
 sg13g2_nand3_1 _11412_ (.B(_03811_),
    .C(_05304_),
    .A(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .Y(_05309_));
 sg13g2_o21ai_1 _11413_ (.B1(_05309_),
    .Y(net24),
    .A1(_02898_),
    .A2(_04179_));
 sg13g2_nand2_1 _11414_ (.Y(_05310_),
    .A(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .B(_03811_));
 sg13g2_a21oi_1 _11415_ (.A1(_03667_),
    .A2(_04180_),
    .Y(_05311_),
    .B1(_05299_));
 sg13g2_nand3_1 _11416_ (.B(_05310_),
    .C(_05311_),
    .A(_05304_),
    .Y(net25));
 sg13g2_dfrbp_1 _11417_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net342),
    .D(_00227_),
    .Q_N(_05717_),
    .Q(\i_tinyqv.cpu.i_core.mip[17] ));
 sg13g2_dfrbp_1 _11418_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net343),
    .D(_00228_),
    .Q_N(_05716_),
    .Q(\i_tinyqv.cpu.i_core.mip[16] ));
 sg13g2_dfrbp_1 _11419_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net344),
    .D(_00229_),
    .Q_N(_05715_),
    .Q(\i_tinyqv.cpu.i_core.mie[19] ));
 sg13g2_dfrbp_1 _11420_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net345),
    .D(_00230_),
    .Q_N(_05714_),
    .Q(\i_tinyqv.cpu.i_core.mie[18] ));
 sg13g2_dfrbp_1 _11421_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net346),
    .D(_00231_),
    .Q_N(_05713_),
    .Q(\i_tinyqv.cpu.i_core.mie[17] ));
 sg13g2_dfrbp_1 _11422_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net347),
    .D(_00232_),
    .Q_N(_05718_),
    .Q(\i_tinyqv.cpu.i_core.mie[16] ));
 sg13g2_inv_1 _08619__1 (.Y(net1396),
    .A(clknet_leaf_49_clk));
 sg13g2_buf_1 _11424_ (.A(net1),
    .X(net12));
 sg13g2_buf_1 _11425_ (.A(net17),
    .X(net13));
 sg13g2_buf_1 _11426_ (.A(net17),
    .X(net14));
 sg13g2_buf_1 _11427_ (.A(net1),
    .X(net15));
 sg13g2_buf_1 _11428_ (.A(net17),
    .X(net16));
 sg13g2_buf_1 _11429_ (.A(net1),
    .X(net18));
 sg13g2_buf_1 _11430_ (.A(net1),
    .X(net19));
 sg13g2_buf_1 _11431_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .X(net20));
 sg13g2_buf_1 _11432_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .X(net23));
 sg13g2_buf_1 _11433_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .X(net26));
 sg13g2_buf_1 _11434_ (.A(uio_out7),
    .X(net27));
 sg13g2_dfrbp_1 \debug_rd_r[0]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net348),
    .D(\debug_rd[0] ),
    .Q_N(_05719_),
    .Q(\debug_rd_r[0] ));
 sg13g2_dfrbp_1 \debug_rd_r[1]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net349),
    .D(net76),
    .Q_N(_05720_),
    .Q(\debug_rd_r[1] ));
 sg13g2_dfrbp_1 \debug_rd_r[2]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net350),
    .D(\debug_rd[2] ),
    .Q_N(_05721_),
    .Q(\debug_rd_r[2] ));
 sg13g2_dfrbp_1 \debug_rd_r[3]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net351),
    .D(\debug_rd[3] ),
    .Q_N(_05712_),
    .Q(\debug_rd_r[3] ));
 sg13g2_dfrbp_1 \debug_register_data$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net352),
    .D(_00233_),
    .Q_N(_05722_),
    .Q(debug_register_data));
 sg13g2_dfrbp_1 \gpio_out[0]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net353),
    .D(_00000_),
    .Q_N(_05723_),
    .Q(\gpio_out[0] ));
 sg13g2_dfrbp_1 \gpio_out[1]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net354),
    .D(_00001_),
    .Q_N(_05724_),
    .Q(\gpio_out[1] ));
 sg13g2_dfrbp_1 \gpio_out[2]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net355),
    .D(_00002_),
    .Q_N(_05725_),
    .Q(\gpio_out[2] ));
 sg13g2_dfrbp_1 \gpio_out[3]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net356),
    .D(_00003_),
    .Q_N(_05726_),
    .Q(\gpio_out[3] ));
 sg13g2_dfrbp_1 \gpio_out[4]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net357),
    .D(_00004_),
    .Q_N(_05727_),
    .Q(\gpio_out[4] ));
 sg13g2_dfrbp_1 \gpio_out[5]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net358),
    .D(_00005_),
    .Q_N(_05728_),
    .Q(\gpio_out[5] ));
 sg13g2_dfrbp_1 \gpio_out[6]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net359),
    .D(_00006_),
    .Q_N(_05729_),
    .Q(\gpio_out[6] ));
 sg13g2_dfrbp_1 \gpio_out[7]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net360),
    .D(_00007_),
    .Q_N(_05730_),
    .Q(\gpio_out[7] ));
 sg13g2_dfrbp_1 \gpio_out_sel[0]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net361),
    .D(_00008_),
    .Q_N(_05731_),
    .Q(\gpio_out_sel[0] ));
 sg13g2_dfrbp_1 \gpio_out_sel[1]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net362),
    .D(_00009_),
    .Q_N(_05732_),
    .Q(\gpio_out_sel[1] ));
 sg13g2_dfrbp_1 \gpio_out_sel[2]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net363),
    .D(_00010_),
    .Q_N(_05733_),
    .Q(\gpio_out_sel[2] ));
 sg13g2_dfrbp_1 \gpio_out_sel[3]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net364),
    .D(_00011_),
    .Q_N(_05734_),
    .Q(\gpio_out_sel[3] ));
 sg13g2_dfrbp_1 \gpio_out_sel[4]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net365),
    .D(_00012_),
    .Q_N(_05735_),
    .Q(\gpio_out_sel[4] ));
 sg13g2_dfrbp_1 \gpio_out_sel[5]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net366),
    .D(_00013_),
    .Q_N(_05736_),
    .Q(\gpio_out_sel[5] ));
 sg13g2_dfrbp_1 \gpio_out_sel[6]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net367),
    .D(_00014_),
    .Q_N(_05737_),
    .Q(\gpio_out_sel[6] ));
 sg13g2_dfrbp_1 \gpio_out_sel[7]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net368),
    .D(_00015_),
    .Q_N(_05738_),
    .Q(\gpio_out_sel[7] ));
 sg13g2_dfrbp_1 \gpio_out_sel[8]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net369),
    .D(_00016_),
    .Q_N(_00171_),
    .Q(\gpio_out_sel[8] ));
 sg13g2_dfrbp_1 \gpio_out_sel[9]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net370),
    .D(_00017_),
    .Q_N(_00204_),
    .Q(\gpio_out_sel[9] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net371),
    .D(_00234_),
    .Q_N(_00222_),
    .Q(\i_debug_uart_tx.cycle_counter[0] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net372),
    .D(_00235_),
    .Q_N(_05711_),
    .Q(\i_debug_uart_tx.cycle_counter[1] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net373),
    .D(_00236_),
    .Q_N(_05710_),
    .Q(\i_debug_uart_tx.cycle_counter[2] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net374),
    .D(_00237_),
    .Q_N(_05709_),
    .Q(\i_debug_uart_tx.cycle_counter[3] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.cycle_counter[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net375),
    .D(_00238_),
    .Q_N(_00168_),
    .Q(\i_debug_uart_tx.cycle_counter[4] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net376),
    .D(_00239_),
    .Q_N(_05708_),
    .Q(\i_debug_uart_tx.data_to_send[0] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net377),
    .D(_00240_),
    .Q_N(_05707_),
    .Q(\i_debug_uart_tx.data_to_send[1] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net378),
    .D(_00241_),
    .Q_N(_05706_),
    .Q(\i_debug_uart_tx.data_to_send[2] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net379),
    .D(_00242_),
    .Q_N(_05705_),
    .Q(\i_debug_uart_tx.data_to_send[3] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net380),
    .D(_00243_),
    .Q_N(_05704_),
    .Q(\i_debug_uart_tx.data_to_send[4] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net381),
    .D(_00244_),
    .Q_N(_05703_),
    .Q(\i_debug_uart_tx.data_to_send[5] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net382),
    .D(_00245_),
    .Q_N(_05702_),
    .Q(\i_debug_uart_tx.data_to_send[6] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.data_to_send[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net383),
    .D(_00246_),
    .Q_N(_05701_),
    .Q(\i_debug_uart_tx.data_to_send[7] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.fsm_state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net384),
    .D(_00247_),
    .Q_N(_05700_),
    .Q(\i_debug_uart_tx.fsm_state[0] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.fsm_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net385),
    .D(_00248_),
    .Q_N(_05699_),
    .Q(\i_debug_uart_tx.fsm_state[1] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.fsm_state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net386),
    .D(_00249_),
    .Q_N(_05698_),
    .Q(\i_debug_uart_tx.fsm_state[2] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.fsm_state[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net387),
    .D(_00250_),
    .Q_N(_05697_),
    .Q(\i_debug_uart_tx.fsm_state[3] ));
 sg13g2_dfrbp_1 \i_debug_uart_tx.txd_reg$_SDFF_PN1_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net388),
    .D(_00251_),
    .Q_N(_05696_),
    .Q(debug_uart_txd));
 sg13g2_dfrbp_1 \i_pwm.pwm_count[0]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net389),
    .D(_00252_),
    .Q_N(_00221_),
    .Q(\i_pwm.pwm_count[0] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_count[1]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net390),
    .D(_00253_),
    .Q_N(_05695_),
    .Q(\i_pwm.pwm_count[1] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_count[2]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net391),
    .D(_00254_),
    .Q_N(_05694_),
    .Q(\i_pwm.pwm_count[2] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_count[3]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net392),
    .D(_00255_),
    .Q_N(_05693_),
    .Q(\i_pwm.pwm_count[3] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_count[4]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net393),
    .D(_00256_),
    .Q_N(_05692_),
    .Q(\i_pwm.pwm_count[4] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_count[5]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net394),
    .D(_00257_),
    .Q_N(_05691_),
    .Q(\i_pwm.pwm_count[5] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_count[6]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net395),
    .D(_00258_),
    .Q_N(_05690_),
    .Q(\i_pwm.pwm_count[6] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_count[7]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net396),
    .D(_00259_),
    .Q_N(_05689_),
    .Q(\i_pwm.pwm_count[7] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_level[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net397),
    .D(_00260_),
    .Q_N(_05688_),
    .Q(\i_pwm.pwm_level[0] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_level[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net398),
    .D(_00261_),
    .Q_N(_05687_),
    .Q(\i_pwm.pwm_level[1] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_level[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net399),
    .D(_00262_),
    .Q_N(_05686_),
    .Q(\i_pwm.pwm_level[2] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_level[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net400),
    .D(_00263_),
    .Q_N(_05685_),
    .Q(\i_pwm.pwm_level[3] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_level[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net401),
    .D(_00264_),
    .Q_N(_05684_),
    .Q(\i_pwm.pwm_level[4] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_level[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net402),
    .D(_00265_),
    .Q_N(_05683_),
    .Q(\i_pwm.pwm_level[5] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_level[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net403),
    .D(_00266_),
    .Q_N(_05682_),
    .Q(\i_pwm.pwm_level[6] ));
 sg13g2_dfrbp_1 \i_pwm.pwm_level[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net404),
    .D(_00267_),
    .Q_N(_05681_),
    .Q(\i_pwm.pwm_level[7] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net405),
    .D(_00268_),
    .Q_N(_05680_),
    .Q(\i_spi.bits_remaining[0] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net406),
    .D(_00269_),
    .Q_N(_05679_),
    .Q(\i_spi.bits_remaining[1] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net407),
    .D(_00270_),
    .Q_N(_05678_),
    .Q(\i_spi.bits_remaining[2] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net408),
    .D(_00271_),
    .Q_N(_05677_),
    .Q(\i_spi.bits_remaining[3] ));
 sg13g2_dfrbp_1 \i_spi.busy$_SDFF_PN0_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net409),
    .D(_00272_),
    .Q_N(_00169_),
    .Q(\i_spi.busy ));
 sg13g2_dfrbp_1 \i_spi.clock_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net410),
    .D(_00273_),
    .Q_N(_05676_),
    .Q(\i_spi.clock_count[0] ));
 sg13g2_dfrbp_1 \i_spi.clock_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net411),
    .D(_00274_),
    .Q_N(_05675_),
    .Q(\i_spi.clock_count[1] ));
 sg13g2_dfrbp_1 \i_spi.clock_divider[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net412),
    .D(_00275_),
    .Q_N(_05674_),
    .Q(\i_spi.clock_divider[0] ));
 sg13g2_dfrbp_1 \i_spi.clock_divider[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net413),
    .D(_00276_),
    .Q_N(_05673_),
    .Q(\i_spi.clock_divider[1] ));
 sg13g2_dfrbp_1 \i_spi.data[0]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net414),
    .D(_00277_),
    .Q_N(_05672_),
    .Q(\i_spi.data[0] ));
 sg13g2_dfrbp_1 \i_spi.data[1]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net415),
    .D(_00278_),
    .Q_N(_05671_),
    .Q(\i_spi.data[1] ));
 sg13g2_dfrbp_1 \i_spi.data[2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net416),
    .D(_00279_),
    .Q_N(_05670_),
    .Q(\i_spi.data[2] ));
 sg13g2_dfrbp_1 \i_spi.data[3]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net417),
    .D(_00280_),
    .Q_N(_05669_),
    .Q(\i_spi.data[3] ));
 sg13g2_dfrbp_1 \i_spi.data[4]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net418),
    .D(_00281_),
    .Q_N(_05668_),
    .Q(\i_spi.data[4] ));
 sg13g2_dfrbp_1 \i_spi.data[5]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net419),
    .D(_00282_),
    .Q_N(_05667_),
    .Q(\i_spi.data[5] ));
 sg13g2_dfrbp_1 \i_spi.data[6]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net420),
    .D(_00283_),
    .Q_N(_05666_),
    .Q(\i_spi.data[6] ));
 sg13g2_dfrbp_1 \i_spi.data[7]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net421),
    .D(_00284_),
    .Q_N(_05665_),
    .Q(\i_spi.data[7] ));
 sg13g2_dfrbp_1 \i_spi.end_txn_reg$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net422),
    .D(_00285_),
    .Q_N(_05664_),
    .Q(\i_spi.end_txn_reg ));
 sg13g2_dfrbp_1 \i_spi.read_latency$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net423),
    .D(_00286_),
    .Q_N(_05663_),
    .Q(\i_spi.read_latency ));
 sg13g2_dfrbp_1 \i_spi.spi_clk_out$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net424),
    .D(_00287_),
    .Q_N(_05662_),
    .Q(\i_spi.spi_clk_out ));
 sg13g2_dfrbp_1 \i_spi.spi_dc$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net425),
    .D(_00288_),
    .Q_N(_05661_),
    .Q(\i_spi.spi_dc ));
 sg13g2_dfrbp_1 \i_spi.spi_select$_SDFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net426),
    .D(_00289_),
    .Q_N(_05660_),
    .Q(\i_spi.spi_select ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.additional_mem_ops[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net427),
    .D(_00290_),
    .Q_N(_00216_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.additional_mem_ops[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net428),
    .D(_00291_),
    .Q_N(_05659_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.additional_mem_ops[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net429),
    .D(_00292_),
    .Q_N(_05658_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.alu_op[0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net430),
    .D(_00293_),
    .Q_N(_05657_),
    .Q(\i_tinyqv.cpu.alu_op[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.alu_op[1]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net431),
    .D(_00294_),
    .Q_N(_00094_),
    .Q(\i_tinyqv.cpu.alu_op[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.alu_op[2]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net432),
    .D(_00295_),
    .Q_N(_00090_),
    .Q(\i_tinyqv.cpu.alu_op[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.alu_op[3]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net433),
    .D(_00296_),
    .Q_N(_00091_),
    .Q(\i_tinyqv.cpu.alu_op[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.counter_hi[0]$_SDFF_PN0_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net434),
    .D(_00297_),
    .Q_N(_00220_),
    .Q(\i_tinyqv.cpu.counter[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.counter_hi[1]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net435),
    .D(_00298_),
    .Q_N(_00093_),
    .Q(\i_tinyqv.cpu.counter[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.counter_hi[2]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net436),
    .D(_00299_),
    .Q_N(_00088_),
    .Q(\i_tinyqv.cpu.counter[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net437),
    .D(_00300_),
    .Q_N(_05656_),
    .Q(\addr[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[10]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net438),
    .D(_00301_),
    .Q_N(_05655_),
    .Q(\addr[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[11]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net439),
    .D(_00302_),
    .Q_N(_05654_),
    .Q(\addr[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[12]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net440),
    .D(_00303_),
    .Q_N(_05653_),
    .Q(\addr[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[13]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net441),
    .D(_00304_),
    .Q_N(_05652_),
    .Q(\addr[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[14]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net442),
    .D(_00305_),
    .Q_N(_05651_),
    .Q(\addr[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[15]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net443),
    .D(_00306_),
    .Q_N(_05650_),
    .Q(\addr[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[16]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net444),
    .D(_00307_),
    .Q_N(_05649_),
    .Q(\addr[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[17]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net445),
    .D(_00308_),
    .Q_N(_05648_),
    .Q(\addr[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[18]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net446),
    .D(_00309_),
    .Q_N(_05647_),
    .Q(\addr[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[19]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net447),
    .D(_00310_),
    .Q_N(_05646_),
    .Q(\addr[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net448),
    .D(_00311_),
    .Q_N(_05645_),
    .Q(\addr[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[20]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net449),
    .D(_00312_),
    .Q_N(_05644_),
    .Q(\addr[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[21]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net450),
    .D(_00313_),
    .Q_N(_05643_),
    .Q(\addr[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[22]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net451),
    .D(_00314_),
    .Q_N(_05642_),
    .Q(\addr[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[23]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net452),
    .D(_00315_),
    .Q_N(_00161_),
    .Q(\addr[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net453),
    .D(_00316_),
    .Q_N(_05641_),
    .Q(\addr[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net454),
    .D(_00317_),
    .Q_N(_05640_),
    .Q(\addr[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net455),
    .D(_00318_),
    .Q_N(_05639_),
    .Q(\addr[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net456),
    .D(_00319_),
    .Q_N(_05638_),
    .Q(\addr[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[2]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net457),
    .D(_00320_),
    .Q_N(_05637_),
    .Q(\addr[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[3]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net458),
    .D(_00321_),
    .Q_N(_05636_),
    .Q(\addr[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[4]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net459),
    .D(_00322_),
    .Q_N(_05635_),
    .Q(\addr[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[5]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net460),
    .D(_00323_),
    .Q_N(_05634_),
    .Q(\addr[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[6]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net461),
    .D(_00324_),
    .Q_N(_05633_),
    .Q(\addr[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[7]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net462),
    .D(_00325_),
    .Q_N(_05632_),
    .Q(\addr[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[8]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net463),
    .D(_00326_),
    .Q_N(_05631_),
    .Q(\addr[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_addr[9]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net464),
    .D(_00327_),
    .Q_N(_05739_),
    .Q(\addr[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_continue$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net465),
    .D(_00030_),
    .Q_N(_05630_),
    .Q(debug_data_continue));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net466),
    .D(_00328_),
    .Q_N(_05629_),
    .Q(\data_to_write[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[10]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net467),
    .D(_00329_),
    .Q_N(_05628_),
    .Q(\data_to_write[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[11]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net468),
    .D(_00330_),
    .Q_N(_05627_),
    .Q(\data_to_write[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[12]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net469),
    .D(_00331_),
    .Q_N(_05626_),
    .Q(\data_to_write[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[13]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net470),
    .D(_00332_),
    .Q_N(_05625_),
    .Q(\data_to_write[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[14]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net471),
    .D(_00333_),
    .Q_N(_05624_),
    .Q(\data_to_write[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[15]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net472),
    .D(_00334_),
    .Q_N(_05623_),
    .Q(\data_to_write[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[16]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net473),
    .D(_00335_),
    .Q_N(_05622_),
    .Q(\data_to_write[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net474),
    .D(_00336_),
    .Q_N(_05621_),
    .Q(\data_to_write[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[18]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net475),
    .D(_00337_),
    .Q_N(_05620_),
    .Q(\data_to_write[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[19]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net476),
    .D(_00338_),
    .Q_N(_05619_),
    .Q(\data_to_write[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net477),
    .D(_00339_),
    .Q_N(_05618_),
    .Q(\data_to_write[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[20]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net478),
    .D(_00340_),
    .Q_N(_05617_),
    .Q(\data_to_write[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[21]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net479),
    .D(_00341_),
    .Q_N(_05616_),
    .Q(\data_to_write[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[22]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net480),
    .D(_00342_),
    .Q_N(_05615_),
    .Q(\data_to_write[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[23]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net481),
    .D(_00343_),
    .Q_N(_05614_),
    .Q(\data_to_write[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[24]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net482),
    .D(_00344_),
    .Q_N(_05613_),
    .Q(\data_to_write[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[25]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net483),
    .D(_00345_),
    .Q_N(_05612_),
    .Q(\data_to_write[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[26]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net484),
    .D(_00346_),
    .Q_N(_05611_),
    .Q(\data_to_write[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[27]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net485),
    .D(_00347_),
    .Q_N(_05610_),
    .Q(\data_to_write[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[28]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net486),
    .D(_00348_),
    .Q_N(_05609_),
    .Q(\data_to_write[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[29]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net487),
    .D(_00349_),
    .Q_N(_05608_),
    .Q(\data_to_write[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net488),
    .D(_00350_),
    .Q_N(_05607_),
    .Q(\data_to_write[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[30]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net489),
    .D(_00351_),
    .Q_N(_05606_),
    .Q(\data_to_write[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[31]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net490),
    .D(_00352_),
    .Q_N(_05605_),
    .Q(\data_to_write[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net491),
    .D(_00353_),
    .Q_N(_05604_),
    .Q(\data_to_write[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net492),
    .D(_00354_),
    .Q_N(_05603_),
    .Q(\data_to_write[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net493),
    .D(_00355_),
    .Q_N(_05602_),
    .Q(\data_to_write[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net494),
    .D(_00356_),
    .Q_N(_05601_),
    .Q(\data_to_write[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net495),
    .D(_00357_),
    .Q_N(_00205_),
    .Q(\data_to_write[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[8]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net496),
    .D(_00358_),
    .Q_N(_05600_),
    .Q(\data_to_write[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_out[9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net497),
    .D(_00359_),
    .Q_N(_05599_),
    .Q(\data_to_write[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_read_n[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net498),
    .D(_00360_),
    .Q_N(_05598_),
    .Q(\i_tinyqv.cpu.data_read_n[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_read_n[1]$_SDFFE_PP1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net499),
    .D(_00361_),
    .Q_N(_05597_),
    .Q(\i_tinyqv.cpu.data_read_n[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_ready_core$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net500),
    .D(_00362_),
    .Q_N(_05596_),
    .Q(\i_tinyqv.cpu.data_ready_core ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_ready_latch$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net501),
    .D(_00363_),
    .Q_N(_05595_),
    .Q(\i_tinyqv.cpu.data_ready_latch ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_write_n[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net502),
    .D(_00364_),
    .Q_N(_05594_),
    .Q(\i_tinyqv.cpu.data_write_n[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.data_write_n[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net503),
    .D(_00365_),
    .Q_N(_05740_),
    .Q(\i_tinyqv.cpu.data_write_n[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.cmp$_DFF_P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net504),
    .D(\i_tinyqv.cpu.i_core.cmp_out ),
    .Q_N(_05741_),
    .Q(\i_tinyqv.cpu.i_core.cmp ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.cy$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net505),
    .D(\i_tinyqv.cpu.i_core.cy_out ),
    .Q_N(_00097_),
    .Q(\i_tinyqv.cpu.i_core.cy ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.cycle[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net506),
    .D(_00366_),
    .Q_N(_00099_),
    .Q(\i_tinyqv.cpu.i_core.cycle[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.cycle[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net507),
    .D(_00367_),
    .Q_N(_05593_),
    .Q(\i_tinyqv.cpu.i_core.cycle[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.cy$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net508),
    .D(_00368_),
    .Q_N(_05592_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.cy ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[0]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net509),
    .D(_00369_),
    .Q_N(_05742_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[10]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net510),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ),
    .Q_N(_05743_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[11]$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net511),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ),
    .Q_N(_05744_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[12]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net512),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ),
    .Q_N(_05745_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[13]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net513),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ),
    .Q_N(_05746_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[14]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net514),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ),
    .Q_N(_05747_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[15]$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net515),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ),
    .Q_N(_05748_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[16]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net516),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ),
    .Q_N(_05749_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[17]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net517),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ),
    .Q_N(_05750_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[18]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net518),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ),
    .Q_N(_05751_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[19]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net519),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ),
    .Q_N(_05591_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[1]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net520),
    .D(_00370_),
    .Q_N(_05752_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[20]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net521),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ),
    .Q_N(_05753_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[21]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net522),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ),
    .Q_N(_05754_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[22]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net523),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ),
    .Q_N(_05755_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[23]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net524),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ),
    .Q_N(_05756_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[24]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net525),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ),
    .Q_N(_05757_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[25]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net526),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ),
    .Q_N(_05758_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[26]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net527),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ),
    .Q_N(_05759_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[27]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net528),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ),
    .Q_N(_05760_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[28]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net529),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ),
    .Q_N(_05761_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[29]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net530),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ),
    .Q_N(_05590_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[2]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net531),
    .D(_00371_),
    .Q_N(_05762_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[30]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net532),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ),
    .Q_N(_05763_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[31]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net533),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ),
    .Q_N(_05589_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[3]$_SDFF_PN0_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net534),
    .D(_00372_),
    .Q_N(_05764_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[4]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net535),
    .D(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .Q_N(_05765_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[5]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net536),
    .D(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .Q_N(_05766_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[6]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net537),
    .D(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .Q_N(_05767_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[7]$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net538),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ),
    .Q_N(_05768_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[8]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net539),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ),
    .Q_N(_05769_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_cycles.register[9]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net540),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ),
    .Q_N(_05588_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.cy$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net541),
    .D(_00373_),
    .Q_N(_00219_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.cy ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[0]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net542),
    .D(_00374_),
    .Q_N(_05770_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[10]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net543),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ),
    .Q_N(_05771_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[11]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net544),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ),
    .Q_N(_05772_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[12]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net545),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ),
    .Q_N(_05773_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[13]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net546),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ),
    .Q_N(_05774_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[14]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net547),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ),
    .Q_N(_05775_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[15]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net548),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ),
    .Q_N(_05776_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[16]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net549),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ),
    .Q_N(_05777_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[17]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net550),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ),
    .Q_N(_05778_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[18]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net551),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ),
    .Q_N(_05779_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[19]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net552),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ),
    .Q_N(_05587_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[1]$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net553),
    .D(_00375_),
    .Q_N(_05780_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[20]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net554),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ),
    .Q_N(_05781_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[21]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net555),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ),
    .Q_N(_05782_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[22]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net556),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ),
    .Q_N(_05783_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[23]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net557),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ),
    .Q_N(_05784_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[24]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net558),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ),
    .Q_N(_05785_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[25]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net559),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ),
    .Q_N(_05786_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[26]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net560),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ),
    .Q_N(_05787_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[27]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net561),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ),
    .Q_N(_05788_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[28]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net562),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ),
    .Q_N(_05789_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[29]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net563),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ),
    .Q_N(_05586_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[2]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net564),
    .D(_00376_),
    .Q_N(_05790_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[30]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net565),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ),
    .Q_N(_05791_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[31]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net566),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ),
    .Q_N(_05585_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[3]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net567),
    .D(_00377_),
    .Q_N(_05792_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[4]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net568),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ),
    .Q_N(_00170_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[5]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net569),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ),
    .Q_N(_05793_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[6]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net570),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ),
    .Q_N(_05794_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[7]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net571),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ),
    .Q_N(_05795_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[8]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net572),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ),
    .Q_N(_05796_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_instrret.register[9]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net573),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ),
    .Q_N(_05797_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][0]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net574),
    .D(_00032_),
    .Q_N(_05798_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][10]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net575),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05799_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][11]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net576),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05800_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][12]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net577),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05801_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][13]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net578),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05802_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][14]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net579),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05803_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][15]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net580),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05804_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][16]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net581),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05805_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][17]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net582),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05806_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][18]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net583),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05807_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][19]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net584),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05808_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][1]$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net585),
    .D(_00033_),
    .Q_N(_05809_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][20]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net586),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05810_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][21]$_DFF_P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net587),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05811_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][22]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net588),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05812_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][23]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net589),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05813_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][24]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net590),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05814_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][25]$_DFF_P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net591),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05815_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][26]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net592),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05816_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][27]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net593),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05817_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][28]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net594),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05818_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][29]$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net595),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05819_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][2]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net596),
    .D(_00034_),
    .Q_N(_05820_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][30]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net597),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05821_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][31]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net598),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05822_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][3]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net599),
    .D(_00035_),
    .Q_N(_05823_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][4]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net600),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05824_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][5]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net601),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05825_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][6]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net602),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05826_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][7]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net603),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05827_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][8]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net604),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05828_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[10][9]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net605),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05829_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][0]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net606),
    .D(_00036_),
    .Q_N(_05830_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][10]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net607),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05831_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][11]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net608),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05832_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][12]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net609),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05833_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][13]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net610),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05834_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][14]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net611),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05835_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][15]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net612),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05836_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][16]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net613),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05837_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][17]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net614),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05838_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][18]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net615),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05839_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][19]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net616),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05840_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][1]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net617),
    .D(_00037_),
    .Q_N(_05841_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][20]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net618),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05842_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][21]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net619),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05843_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][22]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net620),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05844_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][23]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net621),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05845_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][24]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net622),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05846_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][25]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net623),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05847_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][26]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net624),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05848_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][27]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net625),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05849_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][28]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net626),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05850_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][29]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net627),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05851_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][2]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net628),
    .D(_00038_),
    .Q_N(_05852_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][30]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net629),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05853_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][31]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net630),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05854_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][3]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net631),
    .D(_00039_),
    .Q_N(_05855_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][4]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net632),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05856_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][5]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net633),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05857_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][6]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net634),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05858_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][7]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net635),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05859_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][8]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net636),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05860_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[11][9]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net637),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05861_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][0]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net638),
    .D(_00040_),
    .Q_N(_05862_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][10]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net639),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05863_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][11]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net640),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05864_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][12]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net641),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05865_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][13]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net642),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05866_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][14]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net643),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05867_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][15]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net644),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05868_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][16]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net645),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05869_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][17]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net646),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05870_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][18]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net647),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05871_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][19]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net648),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05872_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][1]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net649),
    .D(_00041_),
    .Q_N(_05873_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][20]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net650),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05874_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][21]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net651),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05875_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][22]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net652),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05876_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][23]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net653),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05877_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][24]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net654),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05878_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][25]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net655),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05879_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][26]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net656),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05880_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][27]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net657),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05881_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][28]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net658),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05882_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][29]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net659),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05883_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][2]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net660),
    .D(_00042_),
    .Q_N(_05884_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][30]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net661),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05885_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][31]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net662),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05886_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][3]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net663),
    .D(_00043_),
    .Q_N(_05887_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][4]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net664),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05888_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][5]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net665),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05889_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][6]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net666),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05890_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][7]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net667),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05891_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][8]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net668),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05892_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[12][9]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net669),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05893_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][0]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net670),
    .D(_00044_),
    .Q_N(_05894_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][10]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net671),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05895_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][11]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net672),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05896_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][12]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net673),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05897_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][13]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net674),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05898_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][14]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net675),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05899_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][15]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net676),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05900_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][16]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net677),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05901_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][17]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net678),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05902_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][18]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net679),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05903_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][19]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net680),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05904_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][1]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net681),
    .D(_00045_),
    .Q_N(_05905_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][20]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net682),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05906_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][21]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net683),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05907_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][22]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net684),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05908_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][23]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net685),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05909_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][24]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net686),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05910_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][25]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net687),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05911_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][26]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net688),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05912_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][27]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net689),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05913_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][28]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net690),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05914_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][29]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net691),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05915_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][2]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net692),
    .D(_00046_),
    .Q_N(_05916_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][30]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net693),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05917_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][31]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net694),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05918_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][3]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net695),
    .D(_00047_),
    .Q_N(_05919_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][4]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net696),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05920_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][5]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net697),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05921_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][6]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net698),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05922_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][7]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net699),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05923_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][8]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net700),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05924_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[13][9]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net701),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05925_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][0]$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net702),
    .D(_00048_),
    .Q_N(_05926_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][10]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net703),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05927_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][11]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net704),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05928_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][12]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net705),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05929_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][13]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net706),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05930_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][14]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net707),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05931_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][15]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net708),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05932_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][16]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net709),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05933_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][17]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net710),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05934_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][18]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net711),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05935_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][19]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net712),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05936_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][1]$_DFF_P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net713),
    .D(_00049_),
    .Q_N(_05937_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][20]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net714),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05938_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][21]$_DFF_P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net715),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05939_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][22]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net716),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05940_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][23]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net717),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05941_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][24]$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net718),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05942_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][25]$_DFF_P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net719),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05943_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][26]$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net720),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05944_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][27]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net721),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05945_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][28]$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net722),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05946_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][29]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net723),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05947_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][2]$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net724),
    .D(_00050_),
    .Q_N(_05948_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][30]$_DFF_P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net725),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05949_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][31]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net726),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05950_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][3]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net727),
    .D(_00051_),
    .Q_N(_05951_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][4]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net728),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05952_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][5]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net729),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_05953_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][6]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net730),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_05954_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][7]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net731),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_05955_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][8]$_DFF_P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net732),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05956_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[14][9]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net733),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05957_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][0]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net734),
    .D(_00052_),
    .Q_N(_05958_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][10]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net735),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05959_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][11]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net736),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05960_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][12]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net737),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05961_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][13]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net738),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05962_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][14]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net739),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05963_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][15]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net740),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05964_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][16]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net741),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05965_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][17]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net742),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05966_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][18]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net743),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05967_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][19]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net744),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05968_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][1]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net745),
    .D(_00053_),
    .Q_N(_05969_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][20]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net746),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05970_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][21]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net747),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_05971_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][22]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net748),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_05972_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][23]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net749),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_05973_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][24]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net750),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_05974_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][25]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net751),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_05975_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][26]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net752),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_05976_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][27]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net753),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_05977_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][28]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net754),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_05978_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][29]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net755),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_05979_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][2]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net756),
    .D(_00054_),
    .Q_N(_05980_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][30]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net757),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_05981_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][31]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net758),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_05982_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][3]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net759),
    .D(_00055_),
    .Q_N(_05983_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][4]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net760),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_05984_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][5]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net761),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_00096_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][6]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net762),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_00095_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][7]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net763),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_00092_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][8]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net764),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_05985_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[15][9]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net765),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_05986_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][0]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net766),
    .D(_00056_),
    .Q_N(_05987_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][10]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net767),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_05988_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][11]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net768),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_05989_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][12]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net769),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_05990_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][13]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net770),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_05991_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][14]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net771),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_05992_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][15]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net772),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_05993_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][16]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net773),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_05994_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][17]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net774),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_05995_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][18]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net775),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_05996_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][19]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net776),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_05997_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][1]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net777),
    .D(_00057_),
    .Q_N(_05998_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][20]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net778),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_05999_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][21]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net779),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_06000_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][22]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net780),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_06001_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][23]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net781),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_06002_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][24]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net782),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_06003_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][25]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net783),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_06004_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][26]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net784),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_06005_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][27]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net785),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_06006_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][28]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net786),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_06007_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][29]$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net787),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_06008_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][2]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net788),
    .D(_00058_),
    .Q_N(_06009_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][30]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net789),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_06010_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][31]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net790),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_06011_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][3]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net791),
    .D(_00059_),
    .Q_N(_06012_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][4]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net792),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_06013_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][5]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net793),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_06014_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][6]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net794),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_06015_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][7]$_DFF_P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net795),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_06016_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][8]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net796),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_06017_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[1][9]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net797),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_06018_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][0]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net798),
    .D(_00060_),
    .Q_N(_06019_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][10]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net799),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_06020_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][11]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net800),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_06021_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][12]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net801),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_06022_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][13]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net802),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_06023_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][14]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net803),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_06024_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][15]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net804),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_06025_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][16]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net805),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_06026_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][17]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net806),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_06027_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][18]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net807),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_06028_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][19]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net808),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_06029_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][1]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net809),
    .D(_00061_),
    .Q_N(_06030_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][20]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net810),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_06031_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][21]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net811),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_06032_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][22]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net812),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_06033_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][23]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net813),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_06034_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][24]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net814),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_06035_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][25]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net815),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_06036_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][26]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net816),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_06037_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][27]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net817),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_06038_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][28]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net818),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_06039_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][29]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net819),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_06040_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][2]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net820),
    .D(_00062_),
    .Q_N(_06041_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][30]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net821),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_06042_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][31]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net822),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_06043_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][3]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net823),
    .D(_00063_),
    .Q_N(_06044_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][4]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net824),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_06045_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][5]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net825),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_06046_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][6]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net826),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_06047_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][7]$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net827),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_06048_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][8]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net828),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_06049_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[2][9]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net829),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_06050_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][0]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net830),
    .D(_00064_),
    .Q_N(_06051_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][10]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net831),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_06052_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][11]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net832),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_06053_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][12]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net833),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_06054_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][13]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net834),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_06055_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][14]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net835),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_06056_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][15]$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net836),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_06057_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][16]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net837),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_06058_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][17]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net838),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_06059_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][18]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net839),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_06060_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][19]$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net840),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_06061_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][1]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net841),
    .D(_00065_),
    .Q_N(_06062_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][20]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net842),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_06063_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][21]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net843),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_06064_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][22]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net844),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_06065_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][23]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net845),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_06066_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][24]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net846),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_06067_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][25]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net847),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_06068_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][26]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net848),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_06069_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][27]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net849),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_06070_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][28]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net850),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_06071_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][29]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net851),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_06072_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][2]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net852),
    .D(_00066_),
    .Q_N(_06073_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][30]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net853),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_06074_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][31]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net854),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_06075_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][3]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net855),
    .D(_00067_),
    .Q_N(_06076_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][4]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net856),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_06077_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][5]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net857),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_06078_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][6]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net858),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_06079_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][7]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net859),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_06080_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][8]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net860),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_06081_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[5][9]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net861),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_06082_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][0]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net862),
    .D(_00068_),
    .Q_N(_06083_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][10]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net863),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_06084_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][11]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net864),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_06085_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][12]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net865),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_06086_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][13]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net866),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_06087_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][14]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net867),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_06088_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][15]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net868),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_06089_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][16]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net869),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_06090_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][17]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net870),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_06091_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][18]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net871),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_06092_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][19]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net872),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_06093_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][1]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net873),
    .D(_00069_),
    .Q_N(_06094_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][20]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net874),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_06095_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][21]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net875),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_06096_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][22]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net876),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_06097_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][23]$_DFF_P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net877),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_06098_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][24]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net878),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_06099_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][25]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net879),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_06100_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][26]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net880),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_06101_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][27]$_DFF_P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net881),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_06102_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][28]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net882),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_06103_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][29]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net883),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_06104_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][2]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net884),
    .D(_00070_),
    .Q_N(_06105_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][30]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net885),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_06106_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][31]$_DFF_P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net886),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_06107_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][3]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net887),
    .D(_00071_),
    .Q_N(_06108_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][4]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net888),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_06109_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][5]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net889),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_06110_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][6]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net890),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_06111_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][7]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net891),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_06112_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][8]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net892),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_06113_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[6][9]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net893),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_06114_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][0]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net894),
    .D(_00072_),
    .Q_N(_06115_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][10]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net895),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_06116_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][11]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net896),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_06117_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][12]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net897),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_06118_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][13]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net898),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_06119_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][14]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net899),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_06120_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][15]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net900),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_06121_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][16]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net901),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_06122_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][17]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net902),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_06123_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][18]$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net903),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_06124_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][19]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net904),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_06125_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][1]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net905),
    .D(_00073_),
    .Q_N(_06126_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][20]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net906),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_06127_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][21]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net907),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_06128_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][22]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net908),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_06129_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][23]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net909),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_06130_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][24]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net910),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_06131_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][25]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net911),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_06132_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][26]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net912),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_06133_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][27]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net913),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_06134_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][28]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net914),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_06135_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][29]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net915),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_06136_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][2]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net916),
    .D(_00074_),
    .Q_N(_06137_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][30]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net917),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_06138_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][31]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net918),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_06139_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][3]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net919),
    .D(_00075_),
    .Q_N(_06140_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][4]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net920),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_06141_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][5]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net921),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_06142_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][6]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net922),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_06143_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][7]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net923),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_06144_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][8]$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net924),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_06145_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[7][9]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net925),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_06146_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][0]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net926),
    .D(_00076_),
    .Q_N(_06147_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][10]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net927),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_06148_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][11]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net928),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_06149_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][12]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net929),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_06150_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][13]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net930),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_06151_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][14]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net931),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_06152_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][15]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net932),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_06153_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][16]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net933),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_06154_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][17]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net934),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_06155_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][18]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net935),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_06156_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][19]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net936),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_06157_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][1]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net937),
    .D(_00077_),
    .Q_N(_06158_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][20]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net938),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_06159_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][21]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net939),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_06160_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][22]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net940),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_06161_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][23]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net941),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_06162_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][24]$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net942),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_06163_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][25]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net943),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_06164_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][26]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net944),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_06165_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][27]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net945),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_06166_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][28]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net946),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_06167_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][29]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net947),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_06168_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][2]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net948),
    .D(_00078_),
    .Q_N(_06169_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][30]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net949),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_06170_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][31]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net950),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_06171_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][3]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net951),
    .D(_00079_),
    .Q_N(_06172_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][4]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net952),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_06173_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][5]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net953),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_06174_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][6]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net954),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_06175_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][7]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net955),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_06176_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][8]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net956),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_06177_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[8][9]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net957),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_06178_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][0]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net958),
    .D(_00080_),
    .Q_N(_06179_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][10]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net959),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .Q_N(_06180_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][11]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net960),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .Q_N(_06181_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][12]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net961),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .Q_N(_06182_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][13]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net962),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .Q_N(_06183_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][14]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net963),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .Q_N(_06184_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][15]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net964),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .Q_N(_06185_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][16]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net965),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .Q_N(_06186_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][17]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net966),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .Q_N(_06187_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][18]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net967),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .Q_N(_06188_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][19]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net968),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .Q_N(_06189_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][1]$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net969),
    .D(_00081_),
    .Q_N(_06190_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][20]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net970),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .Q_N(_06191_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][21]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net971),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .Q_N(_06192_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][22]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net972),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .Q_N(_06193_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][23]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net973),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .Q_N(_06194_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][24]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net974),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .Q_N(_06195_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][25]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net975),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .Q_N(_06196_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][26]$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net976),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .Q_N(_06197_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][27]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net977),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .Q_N(_06198_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][28]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net978),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .Q_N(_06199_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][29]$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net979),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .Q_N(_06200_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][2]$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net980),
    .D(_00082_),
    .Q_N(_06201_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][30]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net981),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .Q_N(_06202_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][31]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net982),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .Q_N(_06203_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][3]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net983),
    .D(_00083_),
    .Q_N(_06204_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][4]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net984),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .Q_N(_06205_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][5]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net985),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .Q_N(_06206_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][6]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net986),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .Q_N(_06207_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][7]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net987),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .Q_N(_06208_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][8]$_DFF_P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net988),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .Q_N(_06209_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.i_registers.registers[9][9]$_DFF_P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net989),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .Q_N(_06210_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.instr_retired$_DFF_P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net990),
    .D(_00031_),
    .Q_N(_00218_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.add ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.is_double_fault_r$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net991),
    .D(_00378_),
    .Q_N(_05584_),
    .Q(\i_tinyqv.cpu.i_core.is_double_fault_r ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.last_interrupt_req[0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net992),
    .D(_00379_),
    .Q_N(_05583_),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.last_interrupt_req[1]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net993),
    .D(_00380_),
    .Q_N(_05582_),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.load_done$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net994),
    .D(_00381_),
    .Q_N(_05581_),
    .Q(\i_tinyqv.cpu.i_core.load_done ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.load_top_bit$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net995),
    .D(_00382_),
    .Q_N(_05580_),
    .Q(\i_tinyqv.cpu.i_core.load_top_bit ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mcause[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net996),
    .D(_00383_),
    .Q_N(_05579_),
    .Q(\i_tinyqv.cpu.i_core.mcause[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mcause[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net997),
    .D(_00384_),
    .Q_N(_05578_),
    .Q(\i_tinyqv.cpu.i_core.mcause[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mcause[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net998),
    .D(_00385_),
    .Q_N(_05577_),
    .Q(\i_tinyqv.cpu.i_core.mcause[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mcause[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net999),
    .D(_00386_),
    .Q_N(_05576_),
    .Q(\i_tinyqv.cpu.i_core.mcause[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[0]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1000),
    .D(_00387_),
    .Q_N(_05575_),
    .Q(\i_tinyqv.cpu.i_core.mepc[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[10]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1001),
    .D(_00388_),
    .Q_N(_05574_),
    .Q(\i_tinyqv.cpu.i_core.mepc[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[11]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1002),
    .D(_00389_),
    .Q_N(_05573_),
    .Q(\i_tinyqv.cpu.i_core.mepc[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[12]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1003),
    .D(_00390_),
    .Q_N(_05572_),
    .Q(\i_tinyqv.cpu.i_core.mepc[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[13]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1004),
    .D(_00391_),
    .Q_N(_05571_),
    .Q(\i_tinyqv.cpu.i_core.mepc[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[14]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1005),
    .D(_00392_),
    .Q_N(_05570_),
    .Q(\i_tinyqv.cpu.i_core.mepc[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[15]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1006),
    .D(_00393_),
    .Q_N(_05569_),
    .Q(\i_tinyqv.cpu.i_core.mepc[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[16]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1007),
    .D(_00394_),
    .Q_N(_05568_),
    .Q(\i_tinyqv.cpu.i_core.mepc[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[17]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1008),
    .D(_00395_),
    .Q_N(_05567_),
    .Q(\i_tinyqv.cpu.i_core.mepc[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[18]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1009),
    .D(_00396_),
    .Q_N(_05566_),
    .Q(\i_tinyqv.cpu.i_core.mepc[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[19]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1010),
    .D(_00397_),
    .Q_N(_05565_),
    .Q(\i_tinyqv.cpu.i_core.mepc[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[1]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1011),
    .D(_00398_),
    .Q_N(_05564_),
    .Q(\i_tinyqv.cpu.i_core.mepc[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[20]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1012),
    .D(_00399_),
    .Q_N(_05563_),
    .Q(\i_tinyqv.cpu.i_core.mepc[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[21]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1013),
    .D(_00400_),
    .Q_N(_05562_),
    .Q(\i_tinyqv.cpu.i_core.mepc[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[22]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1014),
    .D(_00401_),
    .Q_N(_05561_),
    .Q(\i_tinyqv.cpu.i_core.mepc[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[23]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1015),
    .D(_00402_),
    .Q_N(_05560_),
    .Q(\i_tinyqv.cpu.i_core.mepc[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[2]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1016),
    .D(_00403_),
    .Q_N(_05559_),
    .Q(\i_tinyqv.cpu.i_core.mepc[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[3]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1017),
    .D(_00404_),
    .Q_N(_05558_),
    .Q(\i_tinyqv.cpu.i_core.mepc[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[4]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1018),
    .D(_00405_),
    .Q_N(_05557_),
    .Q(\i_tinyqv.cpu.i_core.mepc[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[5]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1019),
    .D(_00406_),
    .Q_N(_05556_),
    .Q(\i_tinyqv.cpu.i_core.mepc[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[6]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1020),
    .D(_00407_),
    .Q_N(_05555_),
    .Q(\i_tinyqv.cpu.i_core.mepc[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[7]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1021),
    .D(_00408_),
    .Q_N(_05554_),
    .Q(\i_tinyqv.cpu.i_core.mepc[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[8]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1022),
    .D(_00409_),
    .Q_N(_05553_),
    .Q(\i_tinyqv.cpu.i_core.mepc[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mepc[9]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1023),
    .D(_00410_),
    .Q_N(_05552_),
    .Q(\i_tinyqv.cpu.i_core.mepc[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mstatus_mie$_SDFFE_PP1P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1024),
    .D(_00411_),
    .Q_N(_05551_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mie ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mstatus_mpie$_SDFFE_PP0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1025),
    .D(_00412_),
    .Q_N(_05550_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mpie ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.mstatus_mte$_SDFFE_PP1P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1026),
    .D(_00413_),
    .Q_N(_06211_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mte ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[0]$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1027),
    .D(_00018_),
    .Q_N(_06212_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[10]$_DFF_P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1028),
    .D(_00019_),
    .Q_N(_06213_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[11]$_DFF_P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1029),
    .D(_00020_),
    .Q_N(_05549_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[12]$_SDFF_PP0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1030),
    .D(_00414_),
    .Q_N(_05548_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[13]$_SDFF_PP0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1031),
    .D(_00415_),
    .Q_N(_05547_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[14]$_SDFF_PP0_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1032),
    .D(_00416_),
    .Q_N(_05546_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[15]$_SDFF_PP0_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1033),
    .D(_00417_),
    .Q_N(_06214_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[1]$_DFF_P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1034),
    .D(_00021_),
    .Q_N(_06215_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[2]$_DFF_P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1035),
    .D(_00022_),
    .Q_N(_06216_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[3]$_DFF_P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1036),
    .D(_00023_),
    .Q_N(_06217_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[4]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1037),
    .D(_00024_),
    .Q_N(_06218_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[5]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1038),
    .D(_00025_),
    .Q_N(_06219_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[6]$_DFF_P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1039),
    .D(_00026_),
    .Q_N(_06220_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[7]$_DFF_P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1040),
    .D(_00027_),
    .Q_N(_06221_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[8]$_DFF_P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1041),
    .D(_00028_),
    .Q_N(_06222_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.multiplier.accum[9]$_DFF_P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1042),
    .D(_00029_),
    .Q_N(_05545_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[0]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1043),
    .D(_00418_),
    .Q_N(_05544_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[1]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1044),
    .D(_00419_),
    .Q_N(_05543_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[2]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1045),
    .D(_00420_),
    .Q_N(_05542_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[3]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1046),
    .D(_00421_),
    .Q_N(_05541_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.shift_amt[4]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1047),
    .D(_00422_),
    .Q_N(_05540_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.time_hi[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1048),
    .D(_00423_),
    .Q_N(_00223_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.time_hi[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1049),
    .D(_00424_),
    .Q_N(_05539_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.time_hi[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1050),
    .D(_00425_),
    .Q_N(_05538_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[0]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1051),
    .D(_00426_),
    .Q_N(_00172_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[10]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1052),
    .D(_00427_),
    .Q_N(_00187_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[11]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1053),
    .D(_00428_),
    .Q_N(_00189_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[12]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1054),
    .D(_00429_),
    .Q_N(_00191_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[13]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1055),
    .D(_00430_),
    .Q_N(_00193_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[14]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1056),
    .D(_00431_),
    .Q_N(_00195_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[15]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1057),
    .D(_00432_),
    .Q_N(_00197_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[16]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1058),
    .D(_00433_),
    .Q_N(_00198_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[17]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1059),
    .D(_00434_),
    .Q_N(_00196_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[18]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1060),
    .D(_00435_),
    .Q_N(_00194_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[19]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1061),
    .D(_00436_),
    .Q_N(_00192_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[1]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1062),
    .D(_00437_),
    .Q_N(_00201_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[20]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1063),
    .D(_00438_),
    .Q_N(_00190_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[21]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1064),
    .D(_00439_),
    .Q_N(_00188_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[22]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1065),
    .D(_00440_),
    .Q_N(_00186_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[23]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1066),
    .D(_00441_),
    .Q_N(_00184_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[24]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1067),
    .D(_00442_),
    .Q_N(_00182_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[25]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1068),
    .D(_00443_),
    .Q_N(_00180_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[26]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1069),
    .D(_00444_),
    .Q_N(_00178_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[27]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1070),
    .D(_00445_),
    .Q_N(_00176_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[28]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1071),
    .D(_00446_),
    .Q_N(_00174_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[29]$_SDFFCE_PN0N_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1072),
    .D(_00447_),
    .Q_N(_00200_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[2]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1073),
    .D(_00448_),
    .Q_N(_00199_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[30]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1074),
    .D(_00449_),
    .Q_N(_00202_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[31]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1075),
    .D(_00450_),
    .Q_N(_00203_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[3]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1076),
    .D(_00451_),
    .Q_N(_00173_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[4]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1077),
    .D(_00452_),
    .Q_N(_00175_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[5]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1078),
    .D(_00453_),
    .Q_N(_00177_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[6]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1079),
    .D(_00454_),
    .Q_N(_00179_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[7]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1080),
    .D(_00455_),
    .Q_N(_00181_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[8]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1081),
    .D(_00456_),
    .Q_N(_00183_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.i_core.tmp_data[9]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1082),
    .D(_00457_),
    .Q_N(_00185_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1083),
    .D(_00458_),
    .Q_N(_05537_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1084),
    .D(_00459_),
    .Q_N(_05536_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1085),
    .D(_00460_),
    .Q_N(_05535_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1086),
    .D(_00461_),
    .Q_N(_05534_),
    .Q(\i_tinyqv.cpu.imm[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1087),
    .D(_00462_),
    .Q_N(_05533_),
    .Q(\i_tinyqv.cpu.imm[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1088),
    .D(_00463_),
    .Q_N(_05532_),
    .Q(\i_tinyqv.cpu.imm[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1089),
    .D(_00464_),
    .Q_N(_05531_),
    .Q(\i_tinyqv.cpu.imm[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[16]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1090),
    .D(_00465_),
    .Q_N(_05530_),
    .Q(\i_tinyqv.cpu.imm[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[17]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1091),
    .D(_00466_),
    .Q_N(_05529_),
    .Q(\i_tinyqv.cpu.imm[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[18]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1092),
    .D(_00467_),
    .Q_N(_05528_),
    .Q(\i_tinyqv.cpu.imm[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[19]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1093),
    .D(_00468_),
    .Q_N(_05527_),
    .Q(\i_tinyqv.cpu.imm[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1094),
    .D(_00469_),
    .Q_N(_05526_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[20]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1095),
    .D(_00470_),
    .Q_N(_05525_),
    .Q(\i_tinyqv.cpu.imm[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[21]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1096),
    .D(_00471_),
    .Q_N(_05524_),
    .Q(\i_tinyqv.cpu.imm[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[22]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1097),
    .D(_00472_),
    .Q_N(_05523_),
    .Q(\i_tinyqv.cpu.imm[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1098),
    .D(_00473_),
    .Q_N(_05522_),
    .Q(\i_tinyqv.cpu.imm[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[24]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1099),
    .D(_00474_),
    .Q_N(_05521_),
    .Q(\i_tinyqv.cpu.imm[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[25]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1100),
    .D(_00475_),
    .Q_N(_05520_),
    .Q(\i_tinyqv.cpu.imm[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[26]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1101),
    .D(_00476_),
    .Q_N(_05519_),
    .Q(\i_tinyqv.cpu.imm[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[27]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1102),
    .D(_00477_),
    .Q_N(_05518_),
    .Q(\i_tinyqv.cpu.imm[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[28]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1103),
    .D(_00478_),
    .Q_N(_05517_),
    .Q(\i_tinyqv.cpu.imm[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[29]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1104),
    .D(_00479_),
    .Q_N(_05516_),
    .Q(\i_tinyqv.cpu.imm[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1105),
    .D(_00480_),
    .Q_N(_05515_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[30]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1106),
    .D(_00481_),
    .Q_N(_05514_),
    .Q(\i_tinyqv.cpu.imm[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[31]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1107),
    .D(_00482_),
    .Q_N(_05513_),
    .Q(\i_tinyqv.cpu.imm[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1108),
    .D(_00483_),
    .Q_N(_05512_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1109),
    .D(_00484_),
    .Q_N(_05511_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1110),
    .D(_00485_),
    .Q_N(_05510_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1111),
    .D(_00486_),
    .Q_N(_05509_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1112),
    .D(_00487_),
    .Q_N(_05508_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1113),
    .D(_00488_),
    .Q_N(_05507_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1114),
    .D(_00489_),
    .Q_N(_05506_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][0]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1115),
    .D(_00490_),
    .Q_N(_05505_),
    .Q(\i_tinyqv.cpu.instr_data[0][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1116),
    .D(_00491_),
    .Q_N(_00145_),
    .Q(\i_tinyqv.cpu.instr_data[0][10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1117),
    .D(_00492_),
    .Q_N(_00153_),
    .Q(\i_tinyqv.cpu.instr_data[0][11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1118),
    .D(_00493_),
    .Q_N(_00149_),
    .Q(\i_tinyqv.cpu.instr_data[0][12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1119),
    .D(_00494_),
    .Q_N(_00121_),
    .Q(\i_tinyqv.cpu.instr_data[0][13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1120),
    .D(_00495_),
    .Q_N(_00125_),
    .Q(\i_tinyqv.cpu.instr_data[0][14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1121),
    .D(_00496_),
    .Q_N(_00129_),
    .Q(\i_tinyqv.cpu.instr_data[0][15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1122),
    .D(_00497_),
    .Q_N(_00104_),
    .Q(\i_tinyqv.cpu.instr_data[0][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1123),
    .D(_00498_),
    .Q_N(_05504_),
    .Q(\i_tinyqv.cpu.instr_data[0][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1124),
    .D(_00499_),
    .Q_N(_05503_),
    .Q(\i_tinyqv.cpu.instr_data[0][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1125),
    .D(_00500_),
    .Q_N(_00109_),
    .Q(\i_tinyqv.cpu.instr_data[0][4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1126),
    .D(_00501_),
    .Q_N(_00113_),
    .Q(\i_tinyqv.cpu.instr_data[0][5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1127),
    .D(_00502_),
    .Q_N(_00117_),
    .Q(\i_tinyqv.cpu.instr_data[0][6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1128),
    .D(_00503_),
    .Q_N(_00133_),
    .Q(\i_tinyqv.cpu.instr_data[0][7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1129),
    .D(_00504_),
    .Q_N(_00137_),
    .Q(\i_tinyqv.cpu.instr_data[0][8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1130),
    .D(_00505_),
    .Q_N(_00141_),
    .Q(\i_tinyqv.cpu.instr_data[0][9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][0]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1131),
    .D(_00506_),
    .Q_N(_05502_),
    .Q(\i_tinyqv.cpu.instr_data[1][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1132),
    .D(_00507_),
    .Q_N(_00144_),
    .Q(\i_tinyqv.cpu.instr_data[1][10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1133),
    .D(_00508_),
    .Q_N(_00152_),
    .Q(\i_tinyqv.cpu.instr_data[1][11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1134),
    .D(_00509_),
    .Q_N(_00148_),
    .Q(\i_tinyqv.cpu.instr_data[1][12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1135),
    .D(_00510_),
    .Q_N(_00120_),
    .Q(\i_tinyqv.cpu.instr_data[1][13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1136),
    .D(_00511_),
    .Q_N(_00124_),
    .Q(\i_tinyqv.cpu.instr_data[1][14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1137),
    .D(_00512_),
    .Q_N(_00128_),
    .Q(\i_tinyqv.cpu.instr_data[1][15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1138),
    .D(_00513_),
    .Q_N(_00103_),
    .Q(\i_tinyqv.cpu.instr_data[1][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1139),
    .D(_00514_),
    .Q_N(_05501_),
    .Q(\i_tinyqv.cpu.instr_data[1][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1140),
    .D(_00515_),
    .Q_N(_05500_),
    .Q(\i_tinyqv.cpu.instr_data[1][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1141),
    .D(_00516_),
    .Q_N(_00108_),
    .Q(\i_tinyqv.cpu.instr_data[1][4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1142),
    .D(_00517_),
    .Q_N(_00112_),
    .Q(\i_tinyqv.cpu.instr_data[1][5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1143),
    .D(_00518_),
    .Q_N(_00116_),
    .Q(\i_tinyqv.cpu.instr_data[1][6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1144),
    .D(_00519_),
    .Q_N(_00132_),
    .Q(\i_tinyqv.cpu.instr_data[1][7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1145),
    .D(_00520_),
    .Q_N(_00136_),
    .Q(\i_tinyqv.cpu.instr_data[1][8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1146),
    .D(_00521_),
    .Q_N(_00140_),
    .Q(\i_tinyqv.cpu.instr_data[1][9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][0]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1147),
    .D(_00522_),
    .Q_N(_05499_),
    .Q(\i_tinyqv.cpu.instr_data[2][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1148),
    .D(_00523_),
    .Q_N(_00146_),
    .Q(\i_tinyqv.cpu.instr_data[2][10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1149),
    .D(_00524_),
    .Q_N(_00154_),
    .Q(\i_tinyqv.cpu.instr_data[2][11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1150),
    .D(_00525_),
    .Q_N(_00150_),
    .Q(\i_tinyqv.cpu.instr_data[2][12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1151),
    .D(_00526_),
    .Q_N(_00122_),
    .Q(\i_tinyqv.cpu.instr_data[2][13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1152),
    .D(_00527_),
    .Q_N(_00126_),
    .Q(\i_tinyqv.cpu.instr_data[2][14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1153),
    .D(_00528_),
    .Q_N(_00130_),
    .Q(\i_tinyqv.cpu.instr_data[2][15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1154),
    .D(_00529_),
    .Q_N(_00105_),
    .Q(\i_tinyqv.cpu.instr_data[2][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1155),
    .D(_00530_),
    .Q_N(_05498_),
    .Q(\i_tinyqv.cpu.instr_data[2][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1156),
    .D(_00531_),
    .Q_N(_05497_),
    .Q(\i_tinyqv.cpu.instr_data[2][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1157),
    .D(_00532_),
    .Q_N(_00110_),
    .Q(\i_tinyqv.cpu.instr_data[2][4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1158),
    .D(_00533_),
    .Q_N(_00114_),
    .Q(\i_tinyqv.cpu.instr_data[2][5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1159),
    .D(_00534_),
    .Q_N(_00118_),
    .Q(\i_tinyqv.cpu.instr_data[2][6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1160),
    .D(_00535_),
    .Q_N(_00134_),
    .Q(\i_tinyqv.cpu.instr_data[2][7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1161),
    .D(_00536_),
    .Q_N(_00138_),
    .Q(\i_tinyqv.cpu.instr_data[2][8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1162),
    .D(_00537_),
    .Q_N(_00142_),
    .Q(\i_tinyqv.cpu.instr_data[2][9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1163),
    .D(_00538_),
    .Q_N(_05496_),
    .Q(\i_tinyqv.cpu.instr_data[3][0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1164),
    .D(_00539_),
    .Q_N(_00147_),
    .Q(\i_tinyqv.cpu.instr_data[3][10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1165),
    .D(_00540_),
    .Q_N(_00155_),
    .Q(\i_tinyqv.cpu.instr_data[3][11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1166),
    .D(_00541_),
    .Q_N(_00151_),
    .Q(\i_tinyqv.cpu.instr_data[3][12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1167),
    .D(_00542_),
    .Q_N(_00123_),
    .Q(\i_tinyqv.cpu.instr_data[3][13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1168),
    .D(_00543_),
    .Q_N(_00127_),
    .Q(\i_tinyqv.cpu.instr_data[3][14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1169),
    .D(_00544_),
    .Q_N(_00131_),
    .Q(\i_tinyqv.cpu.instr_data[3][15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1170),
    .D(_00545_),
    .Q_N(_00106_),
    .Q(\i_tinyqv.cpu.instr_data[3][1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1171),
    .D(_00546_),
    .Q_N(_05495_),
    .Q(\i_tinyqv.cpu.instr_data[3][2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1172),
    .D(_00547_),
    .Q_N(_05494_),
    .Q(\i_tinyqv.cpu.instr_data[3][3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1173),
    .D(_00548_),
    .Q_N(_00111_),
    .Q(\i_tinyqv.cpu.instr_data[3][4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1174),
    .D(_00549_),
    .Q_N(_00115_),
    .Q(\i_tinyqv.cpu.instr_data[3][5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1175),
    .D(_00550_),
    .Q_N(_00119_),
    .Q(\i_tinyqv.cpu.instr_data[3][6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1176),
    .D(_00551_),
    .Q_N(_00135_),
    .Q(\i_tinyqv.cpu.instr_data[3][7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1177),
    .D(_00552_),
    .Q_N(_00139_),
    .Q(\i_tinyqv.cpu.instr_data[3][8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1178),
    .D(_00553_),
    .Q_N(_00143_),
    .Q(\i_tinyqv.cpu.instr_data[3][9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1179),
    .D(_00554_),
    .Q_N(_05493_),
    .Q(\i_tinyqv.cpu.instr_data_start[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1180),
    .D(_00555_),
    .Q_N(_05492_),
    .Q(\i_tinyqv.cpu.instr_data_start[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1181),
    .D(_00556_),
    .Q_N(_05491_),
    .Q(\i_tinyqv.cpu.instr_data_start[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1182),
    .D(_00557_),
    .Q_N(_05490_),
    .Q(\i_tinyqv.cpu.instr_data_start[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1183),
    .D(_00558_),
    .Q_N(_05489_),
    .Q(\i_tinyqv.cpu.instr_data_start[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1184),
    .D(_00559_),
    .Q_N(_05488_),
    .Q(\i_tinyqv.cpu.instr_data_start[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1185),
    .D(_00560_),
    .Q_N(_05487_),
    .Q(\i_tinyqv.cpu.instr_data_start[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1186),
    .D(_00561_),
    .Q_N(_05486_),
    .Q(\i_tinyqv.cpu.instr_data_start[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1187),
    .D(_00562_),
    .Q_N(_05485_),
    .Q(\i_tinyqv.cpu.instr_data_start[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1188),
    .D(_00563_),
    .Q_N(_05484_),
    .Q(\i_tinyqv.cpu.instr_data_start[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1189),
    .D(_00564_),
    .Q_N(_05483_),
    .Q(\i_tinyqv.cpu.instr_data_start[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1190),
    .D(_00565_),
    .Q_N(_00163_),
    .Q(\i_tinyqv.cpu.instr_data_start[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1191),
    .D(_00566_),
    .Q_N(_00162_),
    .Q(\i_tinyqv.cpu.instr_data_start[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1192),
    .D(_00567_),
    .Q_N(_05482_),
    .Q(\i_tinyqv.cpu.instr_data_start[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1193),
    .D(_00568_),
    .Q_N(_05481_),
    .Q(\i_tinyqv.cpu.instr_data_start[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1194),
    .D(_00569_),
    .Q_N(_05480_),
    .Q(\i_tinyqv.cpu.instr_data_start[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1195),
    .D(_00570_),
    .Q_N(_05479_),
    .Q(\i_tinyqv.cpu.instr_data_start[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1196),
    .D(_00571_),
    .Q_N(_05478_),
    .Q(\i_tinyqv.cpu.instr_data_start[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1197),
    .D(_00572_),
    .Q_N(_05477_),
    .Q(\i_tinyqv.cpu.instr_data_start[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1198),
    .D(_00573_),
    .Q_N(_05476_),
    .Q(\i_tinyqv.cpu.instr_data_start[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_data_start[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1199),
    .D(_00574_),
    .Q_N(_05475_),
    .Q(\i_tinyqv.cpu.instr_data_start[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_fetch_running$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1200),
    .D(_00575_),
    .Q_N(_00086_),
    .Q(\i_tinyqv.cpu.instr_fetch_running ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_len[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1201),
    .D(_00576_),
    .Q_N(_05474_),
    .Q(\i_tinyqv.cpu.instr_len[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_len[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1202),
    .D(_00577_),
    .Q_N(_05473_),
    .Q(\i_tinyqv.cpu.instr_len[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_valid$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1203),
    .D(_00578_),
    .Q_N(_00100_),
    .Q(debug_instr_valid));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_write_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1204),
    .D(_00579_),
    .Q_N(_00107_),
    .Q(\i_tinyqv.cpu.instr_write_offset[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_write_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1205),
    .D(_00580_),
    .Q_N(_00160_),
    .Q(\i_tinyqv.cpu.instr_write_offset[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.instr_write_offset[2]$_SDFF_PP0_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1206),
    .D(_00581_),
    .Q_N(_05472_),
    .Q(\i_tinyqv.cpu.instr_write_offset[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.interrupt_core$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1207),
    .D(_00582_),
    .Q_N(_00089_),
    .Q(\i_tinyqv.cpu.i_core.is_interrupt ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_alu_imm$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1208),
    .D(_00583_),
    .Q_N(_05471_),
    .Q(\i_tinyqv.cpu.is_alu_imm ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_alu_reg$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1209),
    .D(_00584_),
    .Q_N(_05470_),
    .Q(\i_tinyqv.cpu.is_alu_reg ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_auipc$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1210),
    .D(_00585_),
    .Q_N(_05469_),
    .Q(\i_tinyqv.cpu.is_auipc ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_branch$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1211),
    .D(_00586_),
    .Q_N(_05468_),
    .Q(\i_tinyqv.cpu.is_branch ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_jal$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1212),
    .D(_00587_),
    .Q_N(_05467_),
    .Q(\i_tinyqv.cpu.is_jal ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_jalr$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1213),
    .D(_00588_),
    .Q_N(_05466_),
    .Q(\i_tinyqv.cpu.is_jalr ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_load$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1214),
    .D(_00589_),
    .Q_N(_05465_),
    .Q(\i_tinyqv.cpu.is_load ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_lui$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1215),
    .D(_00590_),
    .Q_N(_05464_),
    .Q(\i_tinyqv.cpu.is_lui ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_store$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1216),
    .D(_00591_),
    .Q_N(_05463_),
    .Q(\i_tinyqv.cpu.is_store ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.is_system$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1217),
    .D(_00592_),
    .Q_N(_05462_),
    .Q(\i_tinyqv.cpu.is_system ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.load_started$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1218),
    .D(_00593_),
    .Q_N(_05461_),
    .Q(\i_tinyqv.cpu.load_started ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.mem_op[0]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1219),
    .D(_00594_),
    .Q_N(_05460_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.mem_op[1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1220),
    .D(_00595_),
    .Q_N(_05459_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.mem_op[2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1221),
    .D(_00596_),
    .Q_N(_05458_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.mem_op_increment_reg$_SDFFCE_PN1P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1222),
    .D(_00597_),
    .Q_N(_05457_),
    .Q(\i_tinyqv.cpu.mem_op_increment_reg ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.no_write_in_progress$_SDFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1223),
    .D(_00598_),
    .Q_N(_00098_),
    .Q(\i_tinyqv.cpu.no_write_in_progress ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.pc_offset[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1224),
    .D(_00599_),
    .Q_N(_00101_),
    .Q(\i_tinyqv.cpu.pc[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.pc_offset[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1225),
    .D(_00600_),
    .Q_N(_00102_),
    .Q(\i_tinyqv.cpu.pc[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1226),
    .D(_00601_),
    .Q_N(_00217_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1227),
    .D(_00602_),
    .Q_N(_05456_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1228),
    .D(_00603_),
    .Q_N(_05455_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1229),
    .D(_00604_),
    .Q_N(_05454_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1230),
    .D(_00605_),
    .Q_N(_05453_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1231),
    .D(_00606_),
    .Q_N(_05452_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1232),
    .D(_00607_),
    .Q_N(_05451_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1233),
    .D(_00608_),
    .Q_N(_05450_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1234),
    .D(_00609_),
    .Q_N(_05449_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1235),
    .D(_00610_),
    .Q_N(_05448_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1236),
    .D(_00611_),
    .Q_N(_05447_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1237),
    .D(_00612_),
    .Q_N(_05446_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.cpu.was_early_branch$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1238),
    .D(_00613_),
    .Q_N(_00087_),
    .Q(\i_tinyqv.cpu.was_early_branch ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.data_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1239),
    .D(_00614_),
    .Q_N(_05445_),
    .Q(\i_tinyqv.mem.data_stall ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.instr_active$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1240),
    .D(_00615_),
    .Q_N(_00085_),
    .Q(\i_tinyqv.mem.instr_active ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.instr_fetch_started$_SDFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1241),
    .D(_00616_),
    .Q_N(_05444_),
    .Q(\i_tinyqv.cpu.instr_fetch_started ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.instr_fetch_stopped$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1242),
    .D(_00617_),
    .Q_N(_05443_),
    .Q(\i_tinyqv.cpu.instr_fetch_stopped ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1243),
    .D(_00618_),
    .Q_N(_05442_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[10]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1244),
    .D(_00619_),
    .Q_N(_05441_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[11]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1245),
    .D(_00620_),
    .Q_N(_05440_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[12]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1246),
    .D(_00621_),
    .Q_N(_05439_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[13]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1247),
    .D(_00622_),
    .Q_N(_05438_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[14]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1248),
    .D(_00623_),
    .Q_N(_05437_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[15]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1249),
    .D(_00624_),
    .Q_N(_05436_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[16]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1250),
    .D(_00625_),
    .Q_N(_05435_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[17]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1251),
    .D(_00626_),
    .Q_N(_05434_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[18]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1252),
    .D(_00627_),
    .Q_N(_05433_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[19]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1253),
    .D(_00628_),
    .Q_N(_05432_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1254),
    .D(_00629_),
    .Q_N(_05431_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[20]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1255),
    .D(_00630_),
    .Q_N(_05430_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[21]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1256),
    .D(_00631_),
    .Q_N(_05429_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[22]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1257),
    .D(_00632_),
    .Q_N(_05428_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[23]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1258),
    .D(_00633_),
    .Q_N(_05427_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1259),
    .D(_00634_),
    .Q_N(_05426_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1260),
    .D(_00635_),
    .Q_N(_05425_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[4]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1261),
    .D(_00636_),
    .Q_N(_05424_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[5]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1262),
    .D(_00637_),
    .Q_N(_05423_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[6]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1263),
    .D(_00638_),
    .Q_N(_05422_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[7]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1264),
    .D(_00639_),
    .Q_N(_05421_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[8]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1265),
    .D(_00640_),
    .Q_N(_05420_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.addr[9]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1266),
    .D(_00641_),
    .Q_N(_05419_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[0]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1267),
    .D(_00642_),
    .Q_N(_00211_),
    .Q(\i_tinyqv.cpu.instr_data_in[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[1]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1268),
    .D(_00643_),
    .Q_N(_00212_),
    .Q(\i_tinyqv.cpu.instr_data_in[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[2]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1269),
    .D(_00644_),
    .Q_N(_00213_),
    .Q(\i_tinyqv.cpu.instr_data_in[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[3]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1270),
    .D(_00645_),
    .Q_N(_00214_),
    .Q(\i_tinyqv.cpu.instr_data_in[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1271),
    .D(_00646_),
    .Q_N(_00208_),
    .Q(\i_tinyqv.cpu.instr_data_in[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1272),
    .D(_00647_),
    .Q_N(_00209_),
    .Q(\i_tinyqv.cpu.instr_data_in[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1273),
    .D(_00648_),
    .Q_N(_00215_),
    .Q(\i_tinyqv.cpu.instr_data_in[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data[7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1274),
    .D(_00649_),
    .Q_N(_00210_),
    .Q(\i_tinyqv.cpu.instr_data_in[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data_ready$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1275),
    .D(_00650_),
    .Q_N(_05418_),
    .Q(\i_tinyqv.mem.q_ctrl.data_ready ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.data_req$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1276),
    .D(_00651_),
    .Q_N(_05417_),
    .Q(\i_tinyqv.mem.q_ctrl.data_req ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1277),
    .D(_00652_),
    .Q_N(_05416_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1278),
    .D(_00653_),
    .Q_N(_05415_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1279),
    .D(_00654_),
    .Q_N(_05414_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.fsm_state[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1280),
    .D(_00655_),
    .Q_N(_00165_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.fsm_state[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1281),
    .D(_00656_),
    .Q_N(_05413_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.fsm_state[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1282),
    .D(_00657_),
    .Q_N(_00157_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.is_writing$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1283),
    .D(_00658_),
    .Q_N(_00164_),
    .Q(\i_tinyqv.mem.q_ctrl.is_writing ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.last_ram_a_sel$_SDFF_PN1_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1284),
    .D(_00659_),
    .Q_N(_05412_),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.last_ram_b_sel$_SDFF_PN1_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1285),
    .D(_00660_),
    .Q_N(_05411_),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.nibbles_remaining[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1286),
    .D(_00661_),
    .Q_N(_05410_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.nibbles_remaining[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1287),
    .D(_00662_),
    .Q_N(_05409_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.nibbles_remaining[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1288),
    .D(_00663_),
    .Q_N(_05408_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.read_cycles_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1289),
    .D(_00664_),
    .Q_N(_00167_),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.read_cycles_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1290),
    .D(_00665_),
    .Q_N(_05407_),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.read_cycles_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1291),
    .D(_00666_),
    .Q_N(_05406_),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_clk_out$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1292),
    .D(_00667_),
    .Q_N(_05405_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_out ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_data_oe[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1293),
    .D(_00668_),
    .Q_N(_05404_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_flash_select$_SDFFE_PP1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1294),
    .D(_00669_),
    .Q_N(_05403_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_flash_select ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1295),
    .D(_00670_),
    .Q_N(_05402_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[1]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1296),
    .D(_00671_),
    .Q_N(_05401_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1297),
    .D(_00672_),
    .Q_N(_05400_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[3]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1298),
    .D(_00673_),
    .Q_N(_05399_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[4]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1299),
    .D(_00674_),
    .Q_N(_05398_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1300),
    .D(_00675_),
    .Q_N(_05397_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[6]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1301),
    .D(_00676_),
    .Q_N(_05396_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_in_buffer[7]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1302),
    .D(_00677_),
    .Q_N(_05395_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_ram_a_select$_SDFFE_PP1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1303),
    .D(_00678_),
    .Q_N(_05394_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.spi_ram_b_select$_SDFFE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1304),
    .D(_00679_),
    .Q_N(_05393_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.q_ctrl.stop_txn_reg$_SDFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1305),
    .D(_00680_),
    .Q_N(_05392_),
    .Q(\i_tinyqv.mem.q_ctrl.stop_txn_reg ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[0]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1306),
    .D(_00681_),
    .Q_N(_05391_),
    .Q(\i_tinyqv.cpu.instr_data_in[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1307),
    .D(_00682_),
    .Q_N(_05390_),
    .Q(\i_tinyqv.mem.qspi_data_buf[10] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[11]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1308),
    .D(_00683_),
    .Q_N(_05389_),
    .Q(\i_tinyqv.mem.qspi_data_buf[11] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[12]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1309),
    .D(_00684_),
    .Q_N(_05388_),
    .Q(\i_tinyqv.mem.qspi_data_buf[12] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1310),
    .D(_00685_),
    .Q_N(_05387_),
    .Q(\i_tinyqv.mem.qspi_data_buf[13] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1311),
    .D(_00686_),
    .Q_N(_05386_),
    .Q(\i_tinyqv.mem.qspi_data_buf[14] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[15]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1312),
    .D(_00687_),
    .Q_N(_05385_),
    .Q(\i_tinyqv.mem.qspi_data_buf[15] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[16]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1313),
    .D(_00688_),
    .Q_N(_05384_),
    .Q(\i_tinyqv.mem.data_from_read[16] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[17]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1314),
    .D(_00689_),
    .Q_N(_05383_),
    .Q(\i_tinyqv.mem.data_from_read[17] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[18]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1315),
    .D(_00690_),
    .Q_N(_05382_),
    .Q(\i_tinyqv.mem.data_from_read[18] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[19]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1316),
    .D(_00691_),
    .Q_N(_05381_),
    .Q(\i_tinyqv.mem.data_from_read[19] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[1]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1317),
    .D(_00692_),
    .Q_N(_05380_),
    .Q(\i_tinyqv.cpu.instr_data_in[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[20]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1318),
    .D(_00693_),
    .Q_N(_05379_),
    .Q(\i_tinyqv.mem.data_from_read[20] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[21]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1319),
    .D(_00694_),
    .Q_N(_05378_),
    .Q(\i_tinyqv.mem.data_from_read[21] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[22]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1320),
    .D(_00695_),
    .Q_N(_05377_),
    .Q(\i_tinyqv.mem.data_from_read[22] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[23]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1321),
    .D(_00696_),
    .Q_N(_05376_),
    .Q(\i_tinyqv.mem.data_from_read[23] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[24]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1322),
    .D(_00697_),
    .Q_N(_05375_),
    .Q(\i_tinyqv.mem.qspi_data_buf[24] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[25]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1323),
    .D(_00698_),
    .Q_N(_05374_),
    .Q(\i_tinyqv.mem.qspi_data_buf[25] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[26]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1324),
    .D(_00699_),
    .Q_N(_05373_),
    .Q(\i_tinyqv.mem.qspi_data_buf[26] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[27]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1325),
    .D(_00700_),
    .Q_N(_05372_),
    .Q(\i_tinyqv.mem.qspi_data_buf[27] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[28]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1326),
    .D(_00701_),
    .Q_N(_05371_),
    .Q(\i_tinyqv.mem.qspi_data_buf[28] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[29]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1327),
    .D(_00702_),
    .Q_N(_05370_),
    .Q(\i_tinyqv.mem.qspi_data_buf[29] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1328),
    .D(_00703_),
    .Q_N(_05369_),
    .Q(\i_tinyqv.cpu.instr_data_in[2] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[30]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1329),
    .D(_00704_),
    .Q_N(_05368_),
    .Q(\i_tinyqv.mem.qspi_data_buf[30] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[31]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1330),
    .D(_00705_),
    .Q_N(_05367_),
    .Q(\i_tinyqv.mem.qspi_data_buf[31] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[3]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1331),
    .D(_00706_),
    .Q_N(_05366_),
    .Q(\i_tinyqv.cpu.instr_data_in[3] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1332),
    .D(_00707_),
    .Q_N(_05365_),
    .Q(\i_tinyqv.cpu.instr_data_in[4] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1333),
    .D(_00708_),
    .Q_N(_05364_),
    .Q(\i_tinyqv.cpu.instr_data_in[5] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[6]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1334),
    .D(_00709_),
    .Q_N(_05363_),
    .Q(\i_tinyqv.cpu.instr_data_in[6] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[7]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1335),
    .D(_00710_),
    .Q_N(_05362_),
    .Q(\i_tinyqv.cpu.instr_data_in[7] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[8]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1336),
    .D(_00711_),
    .Q_N(_05361_),
    .Q(\i_tinyqv.mem.qspi_data_buf[8] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_buf[9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1337),
    .D(_00712_),
    .Q_N(_05360_),
    .Q(\i_tinyqv.mem.qspi_data_buf[9] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_byte_idx[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1338),
    .D(_00713_),
    .Q_N(_00159_),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[0] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_data_byte_idx[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1339),
    .D(_00714_),
    .Q_N(_06223_),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[1] ));
 sg13g2_dfrbp_1 \i_tinyqv.mem.qspi_write_done$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1340),
    .D(_00084_),
    .Q_N(_00156_),
    .Q(\i_tinyqv.mem.qspi_write_done ));
 sg13g2_dfrbp_1 \i_tinyqv.rst_reg_n$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1341),
    .D(\i_debug_uart_tx.resetn ),
    .Q_N(_00166_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.rstn ));
 sg13g2_dfrbp_1 \i_uart_rx.bit_sample$_SDFFE_PN0N_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1342),
    .D(_00715_),
    .Q_N(_05359_),
    .Q(\i_uart_rx.bit_sample ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1343),
    .D(_00716_),
    .Q_N(_00225_),
    .Q(\i_uart_rx.cycle_counter[0] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[10]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1344),
    .D(_00717_),
    .Q_N(_05358_),
    .Q(\i_uart_rx.cycle_counter[10] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1345),
    .D(_00718_),
    .Q_N(_05357_),
    .Q(\i_uart_rx.cycle_counter[1] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1346),
    .D(_00719_),
    .Q_N(_05356_),
    .Q(\i_uart_rx.cycle_counter[2] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1347),
    .D(_00720_),
    .Q_N(_05355_),
    .Q(\i_uart_rx.cycle_counter[3] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1348),
    .D(_00721_),
    .Q_N(_05354_),
    .Q(\i_uart_rx.cycle_counter[4] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[5]$_SDFF_PP0_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1349),
    .D(_00722_),
    .Q_N(_05353_),
    .Q(\i_uart_rx.cycle_counter[5] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1350),
    .D(_00723_),
    .Q_N(_05352_),
    .Q(\i_uart_rx.cycle_counter[6] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1351),
    .D(_00724_),
    .Q_N(_05351_),
    .Q(\i_uart_rx.cycle_counter[7] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[8]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1352),
    .D(_00725_),
    .Q_N(_05350_),
    .Q(\i_uart_rx.cycle_counter[8] ));
 sg13g2_dfrbp_1 \i_uart_rx.cycle_counter[9]$_SDFF_PP0_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1353),
    .D(_00726_),
    .Q_N(_05349_),
    .Q(\i_uart_rx.cycle_counter[9] ));
 sg13g2_dfrbp_1 \i_uart_rx.fsm_state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1354),
    .D(_00727_),
    .Q_N(_00206_),
    .Q(\i_uart_rx.fsm_state[0] ));
 sg13g2_dfrbp_1 \i_uart_rx.fsm_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1355),
    .D(_00728_),
    .Q_N(_05348_),
    .Q(\i_uart_rx.fsm_state[1] ));
 sg13g2_dfrbp_1 \i_uart_rx.fsm_state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1356),
    .D(_00729_),
    .Q_N(_05347_),
    .Q(\i_uart_rx.fsm_state[2] ));
 sg13g2_dfrbp_1 \i_uart_rx.fsm_state[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1357),
    .D(_00730_),
    .Q_N(_05346_),
    .Q(\i_uart_rx.fsm_state[3] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1358),
    .D(_00731_),
    .Q_N(_05345_),
    .Q(\i_uart_rx.recieved_data[0] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[1]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1359),
    .D(_00732_),
    .Q_N(_05344_),
    .Q(\i_uart_rx.recieved_data[1] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[2]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1360),
    .D(_00733_),
    .Q_N(_05343_),
    .Q(\i_uart_rx.recieved_data[2] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[3]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1361),
    .D(_00734_),
    .Q_N(_05342_),
    .Q(\i_uart_rx.recieved_data[3] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1362),
    .D(_00735_),
    .Q_N(_05341_),
    .Q(\i_uart_rx.recieved_data[4] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[5]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1363),
    .D(_00736_),
    .Q_N(_05340_),
    .Q(\i_uart_rx.recieved_data[5] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[6]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1364),
    .D(_00737_),
    .Q_N(_05339_),
    .Q(\i_uart_rx.recieved_data[6] ));
 sg13g2_dfrbp_1 \i_uart_rx.recieved_data[7]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1365),
    .D(_00738_),
    .Q_N(_05338_),
    .Q(\i_uart_rx.recieved_data[7] ));
 sg13g2_dfrbp_1 \i_uart_rx.rxd_reg[0]$_SDFF_PN1_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1366),
    .D(_00739_),
    .Q_N(_00207_),
    .Q(\i_uart_rx.rxd_reg[0] ));
 sg13g2_dfrbp_1 \i_uart_rx.rxd_reg[1]$_SDFF_PN1_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1367),
    .D(_00740_),
    .Q_N(_05337_),
    .Q(\i_uart_rx.rxd_reg[1] ));
 sg13g2_dfrbp_1 \i_uart_rx.uart_rts$_SDFF_PN1_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1368),
    .D(_00741_),
    .Q_N(_05336_),
    .Q(\i_uart_rx.uart_rts ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1369),
    .D(_00742_),
    .Q_N(_00224_),
    .Q(\i_uart_tx.cycle_counter[0] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1370),
    .D(_00743_),
    .Q_N(_05335_),
    .Q(\i_uart_tx.cycle_counter[10] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1371),
    .D(_00744_),
    .Q_N(_05334_),
    .Q(\i_uart_tx.cycle_counter[1] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1372),
    .D(_00745_),
    .Q_N(_05333_),
    .Q(\i_uart_tx.cycle_counter[2] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1373),
    .D(_00746_),
    .Q_N(_05332_),
    .Q(\i_uart_tx.cycle_counter[3] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1374),
    .D(_00747_),
    .Q_N(_05331_),
    .Q(\i_uart_tx.cycle_counter[4] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1375),
    .D(_00748_),
    .Q_N(_05330_),
    .Q(\i_uart_tx.cycle_counter[5] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1376),
    .D(_00749_),
    .Q_N(_05329_),
    .Q(\i_uart_tx.cycle_counter[6] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1377),
    .D(_00750_),
    .Q_N(_05328_),
    .Q(\i_uart_tx.cycle_counter[7] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1378),
    .D(_00751_),
    .Q_N(_05327_),
    .Q(\i_uart_tx.cycle_counter[8] ));
 sg13g2_dfrbp_1 \i_uart_tx.cycle_counter[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1379),
    .D(_00752_),
    .Q_N(_05326_),
    .Q(\i_uart_tx.cycle_counter[9] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1380),
    .D(_00753_),
    .Q_N(_05325_),
    .Q(\i_uart_tx.data_to_send[0] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1381),
    .D(_00754_),
    .Q_N(_05324_),
    .Q(\i_uart_tx.data_to_send[1] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1382),
    .D(_00755_),
    .Q_N(_05323_),
    .Q(\i_uart_tx.data_to_send[2] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1383),
    .D(_00756_),
    .Q_N(_05322_),
    .Q(\i_uart_tx.data_to_send[3] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1384),
    .D(_00757_),
    .Q_N(_05321_),
    .Q(\i_uart_tx.data_to_send[4] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1385),
    .D(_00758_),
    .Q_N(_05320_),
    .Q(\i_uart_tx.data_to_send[5] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1386),
    .D(_00759_),
    .Q_N(_05319_),
    .Q(\i_uart_tx.data_to_send[6] ));
 sg13g2_dfrbp_1 \i_uart_tx.data_to_send[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1387),
    .D(_00760_),
    .Q_N(_05318_),
    .Q(\i_uart_tx.data_to_send[7] ));
 sg13g2_dfrbp_1 \i_uart_tx.fsm_state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1388),
    .D(_00761_),
    .Q_N(_05317_),
    .Q(\i_uart_tx.fsm_state[0] ));
 sg13g2_dfrbp_1 \i_uart_tx.fsm_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1389),
    .D(_00762_),
    .Q_N(_05316_),
    .Q(\i_uart_tx.fsm_state[1] ));
 sg13g2_dfrbp_1 \i_uart_tx.fsm_state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1390),
    .D(_00763_),
    .Q_N(_05315_),
    .Q(\i_uart_tx.fsm_state[2] ));
 sg13g2_dfrbp_1 \i_uart_tx.fsm_state[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1391),
    .D(_00764_),
    .Q_N(_05314_),
    .Q(\i_uart_tx.fsm_state[3] ));
 sg13g2_dfrbp_1 \i_uart_tx.txd_reg$_SDFF_PN1_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1392),
    .D(_00765_),
    .Q_N(_05313_),
    .Q(\i_uart_tx.txd_reg ));
 sg13g2_dfrbp_1 \rst_reg_n$_DFF_N_  (.CLK(net1396),
    .RESET_B(net1393),
    .D(net1),
    .Q_N(_00158_),
    .Q(\i_debug_uart_tx.resetn ));
 sg13g2_dfrbp_1 \ui_in_reg[0]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1394),
    .D(net2),
    .Q_N(_06224_),
    .Q(\i_tinyqv.cpu.i_core.interrupt_req[0] ));
 sg13g2_dfrbp_1 \ui_in_reg[1]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1395),
    .D(net3),
    .Q_N(_05312_),
    .Q(\i_tinyqv.cpu.i_core.interrupt_req[1] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[0]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[1]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[2]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[4]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[5]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[6]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[7]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[0]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[1]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[2]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[3]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[4]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_out[5]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[6]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[7]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[0]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[1]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[2]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[3]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[4]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uo_out[5]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[6]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout36 (.A(_03459_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_03441_),
    .X(net37));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(_03404_));
 sg13g2_buf_2 fanout39 (.A(_03187_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_03172_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_03128_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_03021_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_05011_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_04997_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_04615_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_04609_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_03930_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_03896_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_03819_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_03803_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_03640_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_03638_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_03603_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_03600_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_03378_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_03127_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_05138_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_04909_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_03927_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_03870_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_03865_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_03807_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_03712_),
    .X(net63));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(_03662_));
 sg13g2_buf_2 fanout65 (.A(_03626_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_03624_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_04983_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_03806_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_03797_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_05022_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_04998_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_03863_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_03713_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_03696_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_03652_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(\debug_rd[1] ),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_04599_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_05002_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(\debug_rd[2] ),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(\debug_rd[0] ),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_05001_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_04987_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_04984_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_03650_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_03488_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_01563_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_03091_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_03485_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_03389_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_03356_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_03529_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_03483_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_05248_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_03509_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_03443_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_03371_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_03370_),
    .X(net97));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(_03238_));
 sg13g2_buf_2 fanout99 (.A(_03226_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_03129_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_02090_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_03513_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_03479_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_03351_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_03350_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_03190_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_03177_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_03174_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_03158_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_03157_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_03153_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_03150_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_03136_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_02292_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_02284_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_02213_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_04786_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_04501_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_04191_),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(_03400_));
 sg13g2_buf_2 fanout121 (.A(_03156_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_03140_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_02568_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_02533_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_02526_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_02052_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_01960_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_01877_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_01868_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_01837_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_01824_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_01786_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_01747_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_01713_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_01531_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_01525_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_01449_),
    .X(net137));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(_04364_));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(_04363_));
 sg13g2_buf_2 fanout140 (.A(_03144_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_02540_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_01846_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_01831_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_01829_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_01746_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_01555_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_01503_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_04841_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_04762_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_04726_),
    .X(net150));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(_04400_));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_04399_));
 sg13g2_buf_2 fanout153 (.A(_04395_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_04393_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_03130_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_02513_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_01828_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_01807_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_01590_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_01507_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_01477_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_01358_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_01014_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03867_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03814_),
    .X(net165));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(_03447_));
 sg13g2_buf_2 fanout167 (.A(_03270_),
    .X(net167));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(_03228_));
 sg13g2_buf_2 fanout169 (.A(_03222_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_02502_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_01533_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_01501_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_01479_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_01213_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_04993_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_04989_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_03269_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_03221_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_02591_),
    .X(net179));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(_02406_));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(_02382_));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(_01587_));
 sg13g2_buf_2 fanout183 (.A(_01544_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_01444_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_01437_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_01227_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_00979_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_04992_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_04988_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_04759_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_04604_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_04332_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_04173_),
    .X(net193));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(_02592_));
 sg13g2_buf_2 fanout195 (.A(_02574_),
    .X(net195));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(_02510_));
 sg13g2_buf_2 fanout197 (.A(_02508_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_01675_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_01643_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_01491_),
    .X(net200));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(_01441_));
 sg13g2_buf_2 fanout202 (.A(_01436_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_00822_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_04950_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_04931_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_04906_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_04891_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_04839_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_04817_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_04816_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_04795_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_04465_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_04431_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_04320_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_04306_),
    .X(net215));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(_02573_));
 sg13g2_buf_2 fanout217 (.A(_02561_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_02514_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_02398_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_01732_),
    .X(net220));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(_01440_));
 sg13g2_buf_2 fanout222 (.A(_01217_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_00924_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_00897_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_04938_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_04890_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_03877_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_03084_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_03063_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_02530_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_01716_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_01692_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_01565_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_01259_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_01216_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_01104_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_01082_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_01016_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_00874_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_00847_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_00839_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_00779_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_04372_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_04308_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_04287_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_04277_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_04169_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_03897_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_03876_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_03821_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_03657_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_03230_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_03227_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_03095_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_02653_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_02650_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_02646_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_02626_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_02621_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_02612_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_02611_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_02608_),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_02446_));
 sg13g2_buf_2 fanout264 (.A(_02391_),
    .X(net264));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_02388_));
 sg13g2_buf_2 fanout266 (.A(_02384_),
    .X(net266));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_02376_));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_02375_));
 sg13g2_buf_2 fanout269 (.A(_01784_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_01773_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_01768_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_01743_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_01742_),
    .X(net273));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_01672_));
 sg13g2_buf_2 fanout275 (.A(_01649_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_01300_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_01286_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_01236_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_01202_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_00879_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_00877_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_00863_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_00858_),
    .X(net283));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_00835_));
 sg13g2_buf_2 fanout285 (.A(_00833_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_00804_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_00801_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_00790_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_00783_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_00780_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_00775_),
    .X(net291));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(_00773_));
 sg13g2_buf_2 fanout293 (.A(_00767_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_03820_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_02625_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_02613_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_02607_),
    .X(net297));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(_02397_));
 sg13g2_buf_2 fanout299 (.A(_02283_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_02050_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_02049_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_01897_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_01794_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_01734_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_01730_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_01727_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_01721_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_01718_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_01714_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_01697_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_01650_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_01647_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_01575_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_01409_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_01370_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_01369_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_01366_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_01337_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_01335_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_01334_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_01311_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_01298_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_01071_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_01062_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_01025_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_01019_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_01017_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_00964_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_00963_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_00919_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_00857_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_00855_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_00843_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_00836_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_00818_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_00792_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_00791_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_00769_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_00766_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_01343_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_01332_),
    .X(net341));
 sg13g2_tiehi _11417__342 (.L_HI(net342));
 sg13g2_tiehi _11418__343 (.L_HI(net343));
 sg13g2_tiehi _11419__344 (.L_HI(net344));
 sg13g2_tiehi _11420__345 (.L_HI(net345));
 sg13g2_tiehi _11421__346 (.L_HI(net346));
 sg13g2_tiehi _11422__347 (.L_HI(net347));
 sg13g2_tiehi \debug_rd_r[0]$_DFF_P__348  (.L_HI(net348));
 sg13g2_tiehi \debug_rd_r[1]$_DFF_P__349  (.L_HI(net349));
 sg13g2_tiehi \debug_rd_r[2]$_DFF_P__350  (.L_HI(net350));
 sg13g2_tiehi \debug_rd_r[3]$_DFF_P__351  (.L_HI(net351));
 sg13g2_tiehi \debug_register_data$_DFFE_PP__352  (.L_HI(net352));
 sg13g2_tiehi \gpio_out[0]$_DFF_P__353  (.L_HI(net353));
 sg13g2_tiehi \gpio_out[1]$_DFF_P__354  (.L_HI(net354));
 sg13g2_tiehi \gpio_out[2]$_DFF_P__355  (.L_HI(net355));
 sg13g2_tiehi \gpio_out[3]$_DFF_P__356  (.L_HI(net356));
 sg13g2_tiehi \gpio_out[4]$_DFF_P__357  (.L_HI(net357));
 sg13g2_tiehi \gpio_out[5]$_DFF_P__358  (.L_HI(net358));
 sg13g2_tiehi \gpio_out[6]$_DFF_P__359  (.L_HI(net359));
 sg13g2_tiehi \gpio_out[7]$_DFF_P__360  (.L_HI(net360));
 sg13g2_tiehi \gpio_out_sel[0]$_DFF_P__361  (.L_HI(net361));
 sg13g2_tiehi \gpio_out_sel[1]$_DFF_P__362  (.L_HI(net362));
 sg13g2_tiehi \gpio_out_sel[2]$_DFF_P__363  (.L_HI(net363));
 sg13g2_tiehi \gpio_out_sel[3]$_DFF_P__364  (.L_HI(net364));
 sg13g2_tiehi \gpio_out_sel[4]$_DFF_P__365  (.L_HI(net365));
 sg13g2_tiehi \gpio_out_sel[5]$_DFF_P__366  (.L_HI(net366));
 sg13g2_tiehi \gpio_out_sel[6]$_DFF_P__367  (.L_HI(net367));
 sg13g2_tiehi \gpio_out_sel[7]$_DFF_P__368  (.L_HI(net368));
 sg13g2_tiehi \gpio_out_sel[8]$_DFF_P__369  (.L_HI(net369));
 sg13g2_tiehi \gpio_out_sel[9]$_DFF_P__370  (.L_HI(net370));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[0]$_SDFFE_PP0N__371  (.L_HI(net371));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[1]$_SDFFE_PP0N__372  (.L_HI(net372));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[2]$_SDFFE_PP0N__373  (.L_HI(net373));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[3]$_SDFFE_PP0N__374  (.L_HI(net374));
 sg13g2_tiehi \i_debug_uart_tx.cycle_counter[4]$_SDFFE_PP0N__375  (.L_HI(net375));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[0]$_SDFFE_PN0P__376  (.L_HI(net376));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[1]$_SDFFE_PN0P__377  (.L_HI(net377));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[2]$_SDFFE_PN0P__378  (.L_HI(net378));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[3]$_SDFFE_PN0P__379  (.L_HI(net379));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[4]$_SDFFE_PN0P__380  (.L_HI(net380));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[5]$_SDFFE_PN0P__381  (.L_HI(net381));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[6]$_SDFFE_PN0P__382  (.L_HI(net382));
 sg13g2_tiehi \i_debug_uart_tx.data_to_send[7]$_SDFFE_PN0P__383  (.L_HI(net383));
 sg13g2_tiehi \i_debug_uart_tx.fsm_state[0]$_SDFFE_PN0P__384  (.L_HI(net384));
 sg13g2_tiehi \i_debug_uart_tx.fsm_state[1]$_SDFFE_PN0P__385  (.L_HI(net385));
 sg13g2_tiehi \i_debug_uart_tx.fsm_state[2]$_SDFFE_PN0P__386  (.L_HI(net386));
 sg13g2_tiehi \i_debug_uart_tx.fsm_state[3]$_SDFFE_PN0P__387  (.L_HI(net387));
 sg13g2_tiehi \i_debug_uart_tx.txd_reg$_SDFF_PN1__388  (.L_HI(net388));
 sg13g2_tiehi \i_pwm.pwm_count[0]$_SDFF_PP0__389  (.L_HI(net389));
 sg13g2_tiehi \i_pwm.pwm_count[1]$_SDFF_PP0__390  (.L_HI(net390));
 sg13g2_tiehi \i_pwm.pwm_count[2]$_SDFF_PP0__391  (.L_HI(net391));
 sg13g2_tiehi \i_pwm.pwm_count[3]$_SDFF_PP0__392  (.L_HI(net392));
 sg13g2_tiehi \i_pwm.pwm_count[4]$_SDFF_PP0__393  (.L_HI(net393));
 sg13g2_tiehi \i_pwm.pwm_count[5]$_SDFF_PP0__394  (.L_HI(net394));
 sg13g2_tiehi \i_pwm.pwm_count[6]$_SDFF_PP0__395  (.L_HI(net395));
 sg13g2_tiehi \i_pwm.pwm_count[7]$_SDFF_PP0__396  (.L_HI(net396));
 sg13g2_tiehi \i_pwm.pwm_level[0]$_SDFFE_PN0P__397  (.L_HI(net397));
 sg13g2_tiehi \i_pwm.pwm_level[1]$_SDFFE_PN0P__398  (.L_HI(net398));
 sg13g2_tiehi \i_pwm.pwm_level[2]$_SDFFE_PN0P__399  (.L_HI(net399));
 sg13g2_tiehi \i_pwm.pwm_level[3]$_SDFFE_PN0P__400  (.L_HI(net400));
 sg13g2_tiehi \i_pwm.pwm_level[4]$_SDFFE_PN0P__401  (.L_HI(net401));
 sg13g2_tiehi \i_pwm.pwm_level[5]$_SDFFE_PN0P__402  (.L_HI(net402));
 sg13g2_tiehi \i_pwm.pwm_level[6]$_SDFFE_PN0P__403  (.L_HI(net403));
 sg13g2_tiehi \i_pwm.pwm_level[7]$_SDFFE_PN0P__404  (.L_HI(net404));
 sg13g2_tiehi \i_spi.bits_remaining[0]$_SDFFE_PN0P__405  (.L_HI(net405));
 sg13g2_tiehi \i_spi.bits_remaining[1]$_SDFFE_PN0P__406  (.L_HI(net406));
 sg13g2_tiehi \i_spi.bits_remaining[2]$_SDFFE_PN0P__407  (.L_HI(net407));
 sg13g2_tiehi \i_spi.bits_remaining[3]$_SDFFE_PN0P__408  (.L_HI(net408));
 sg13g2_tiehi \i_spi.busy$_SDFF_PN0__409  (.L_HI(net409));
 sg13g2_tiehi \i_spi.clock_count[0]$_SDFFE_PN0P__410  (.L_HI(net410));
 sg13g2_tiehi \i_spi.clock_count[1]$_SDFFE_PN0P__411  (.L_HI(net411));
 sg13g2_tiehi \i_spi.clock_divider[0]$_SDFFE_PN1P__412  (.L_HI(net412));
 sg13g2_tiehi \i_spi.clock_divider[1]$_SDFFE_PN0P__413  (.L_HI(net413));
 sg13g2_tiehi \i_spi.data[0]$_DFFE_PP__414  (.L_HI(net414));
 sg13g2_tiehi \i_spi.data[1]$_DFFE_PP__415  (.L_HI(net415));
 sg13g2_tiehi \i_spi.data[2]$_DFFE_PP__416  (.L_HI(net416));
 sg13g2_tiehi \i_spi.data[3]$_DFFE_PP__417  (.L_HI(net417));
 sg13g2_tiehi \i_spi.data[4]$_DFFE_PP__418  (.L_HI(net418));
 sg13g2_tiehi \i_spi.data[5]$_DFFE_PP__419  (.L_HI(net419));
 sg13g2_tiehi \i_spi.data[6]$_DFFE_PP__420  (.L_HI(net420));
 sg13g2_tiehi \i_spi.data[7]$_DFFE_PP__421  (.L_HI(net421));
 sg13g2_tiehi \i_spi.end_txn_reg$_DFFE_PP__422  (.L_HI(net422));
 sg13g2_tiehi \i_spi.read_latency$_SDFFE_PN0P__423  (.L_HI(net423));
 sg13g2_tiehi \i_spi.spi_clk_out$_SDFFE_PN0P__424  (.L_HI(net424));
 sg13g2_tiehi \i_spi.spi_dc$_DFFE_PP__425  (.L_HI(net425));
 sg13g2_tiehi \i_spi.spi_select$_SDFFE_PN1P__426  (.L_HI(net426));
 sg13g2_tiehi \i_tinyqv.cpu.additional_mem_ops[0]$_SDFFE_PN0P__427  (.L_HI(net427));
 sg13g2_tiehi \i_tinyqv.cpu.additional_mem_ops[1]$_SDFFE_PN0P__428  (.L_HI(net428));
 sg13g2_tiehi \i_tinyqv.cpu.additional_mem_ops[2]$_SDFFE_PN0P__429  (.L_HI(net429));
 sg13g2_tiehi \i_tinyqv.cpu.alu_op[0]$_DFFE_PP__430  (.L_HI(net430));
 sg13g2_tiehi \i_tinyqv.cpu.alu_op[1]$_DFFE_PP__431  (.L_HI(net431));
 sg13g2_tiehi \i_tinyqv.cpu.alu_op[2]$_DFFE_PP__432  (.L_HI(net432));
 sg13g2_tiehi \i_tinyqv.cpu.alu_op[3]$_DFFE_PP__433  (.L_HI(net433));
 sg13g2_tiehi \i_tinyqv.cpu.counter_hi[0]$_SDFF_PN0__434  (.L_HI(net434));
 sg13g2_tiehi \i_tinyqv.cpu.counter_hi[1]$_SDFF_PN0__435  (.L_HI(net435));
 sg13g2_tiehi \i_tinyqv.cpu.counter_hi[2]$_SDFF_PN0__436  (.L_HI(net436));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[0]$_DFFE_PP__437  (.L_HI(net437));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[10]$_DFFE_PP__438  (.L_HI(net438));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[11]$_DFFE_PP__439  (.L_HI(net439));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[12]$_DFFE_PP__440  (.L_HI(net440));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[13]$_DFFE_PP__441  (.L_HI(net441));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[14]$_DFFE_PP__442  (.L_HI(net442));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[15]$_DFFE_PP__443  (.L_HI(net443));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[16]$_DFFE_PP__444  (.L_HI(net444));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[17]$_DFFE_PP__445  (.L_HI(net445));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[18]$_DFFE_PP__446  (.L_HI(net446));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[19]$_DFFE_PP__447  (.L_HI(net447));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[1]$_DFFE_PP__448  (.L_HI(net448));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[20]$_DFFE_PP__449  (.L_HI(net449));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[21]$_DFFE_PP__450  (.L_HI(net450));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[22]$_DFFE_PP__451  (.L_HI(net451));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[23]$_DFFE_PP__452  (.L_HI(net452));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[24]$_SDFFE_PN0P__453  (.L_HI(net453));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[25]$_SDFFE_PN0P__454  (.L_HI(net454));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[26]$_SDFFE_PN0P__455  (.L_HI(net455));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[27]$_SDFFE_PN0P__456  (.L_HI(net456));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[2]$_DFFE_PP__457  (.L_HI(net457));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[3]$_DFFE_PP__458  (.L_HI(net458));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[4]$_DFFE_PP__459  (.L_HI(net459));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[5]$_DFFE_PP__460  (.L_HI(net460));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[6]$_DFFE_PP__461  (.L_HI(net461));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[7]$_DFFE_PP__462  (.L_HI(net462));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[8]$_DFFE_PP__463  (.L_HI(net463));
 sg13g2_tiehi \i_tinyqv.cpu.data_addr[9]$_DFFE_PP__464  (.L_HI(net464));
 sg13g2_tiehi \i_tinyqv.cpu.data_continue$_DFF_P__465  (.L_HI(net465));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[0]$_DFFE_PP__466  (.L_HI(net466));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[10]$_DFFE_PP__467  (.L_HI(net467));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[11]$_DFFE_PP__468  (.L_HI(net468));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[12]$_DFFE_PP__469  (.L_HI(net469));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[13]$_DFFE_PP__470  (.L_HI(net470));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[14]$_DFFE_PP__471  (.L_HI(net471));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[15]$_DFFE_PP__472  (.L_HI(net472));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[16]$_DFFE_PP__473  (.L_HI(net473));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[17]$_DFFE_PP__474  (.L_HI(net474));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[18]$_DFFE_PP__475  (.L_HI(net475));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[19]$_DFFE_PP__476  (.L_HI(net476));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[1]$_DFFE_PP__477  (.L_HI(net477));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[20]$_DFFE_PP__478  (.L_HI(net478));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[21]$_DFFE_PP__479  (.L_HI(net479));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[22]$_DFFE_PP__480  (.L_HI(net480));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[23]$_DFFE_PP__481  (.L_HI(net481));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[24]$_DFFE_PP__482  (.L_HI(net482));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[25]$_DFFE_PP__483  (.L_HI(net483));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[26]$_DFFE_PP__484  (.L_HI(net484));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[27]$_DFFE_PP__485  (.L_HI(net485));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[28]$_DFFE_PP__486  (.L_HI(net486));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[29]$_DFFE_PP__487  (.L_HI(net487));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[2]$_DFFE_PP__488  (.L_HI(net488));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[30]$_DFFE_PP__489  (.L_HI(net489));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[31]$_DFFE_PP__490  (.L_HI(net490));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[3]$_DFFE_PP__491  (.L_HI(net491));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[4]$_DFFE_PP__492  (.L_HI(net492));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[5]$_DFFE_PP__493  (.L_HI(net493));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[6]$_DFFE_PP__494  (.L_HI(net494));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[7]$_DFFE_PP__495  (.L_HI(net495));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[8]$_DFFE_PP__496  (.L_HI(net496));
 sg13g2_tiehi \i_tinyqv.cpu.data_out[9]$_DFFE_PP__497  (.L_HI(net497));
 sg13g2_tiehi \i_tinyqv.cpu.data_read_n[0]$_SDFFE_PP1P__498  (.L_HI(net498));
 sg13g2_tiehi \i_tinyqv.cpu.data_read_n[1]$_SDFFE_PP1P__499  (.L_HI(net499));
 sg13g2_tiehi \i_tinyqv.cpu.data_ready_core$_SDFFE_PN0P__500  (.L_HI(net500));
 sg13g2_tiehi \i_tinyqv.cpu.data_ready_latch$_SDFF_PP0__501  (.L_HI(net501));
 sg13g2_tiehi \i_tinyqv.cpu.data_write_n[0]$_SDFFE_PN1P__502  (.L_HI(net502));
 sg13g2_tiehi \i_tinyqv.cpu.data_write_n[1]$_SDFFE_PN1P__503  (.L_HI(net503));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.cmp$_DFF_P__504  (.L_HI(net504));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.cy$_DFF_P__505  (.L_HI(net505));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.cycle[0]$_SDFFE_PN0P__506  (.L_HI(net506));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.cycle[1]$_SDFFE_PN0P__507  (.L_HI(net507));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.cy$_SDFF_PN0__508  (.L_HI(net508));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[0]$_SDFF_PN0__509  (.L_HI(net509));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[10]$_DFF_P__510  (.L_HI(net510));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[11]$_DFF_P__511  (.L_HI(net511));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[12]$_DFF_P__512  (.L_HI(net512));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[13]$_DFF_P__513  (.L_HI(net513));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[14]$_DFF_P__514  (.L_HI(net514));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[15]$_DFF_P__515  (.L_HI(net515));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[16]$_DFF_P__516  (.L_HI(net516));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[17]$_DFF_P__517  (.L_HI(net517));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[18]$_DFF_P__518  (.L_HI(net518));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[19]$_DFF_P__519  (.L_HI(net519));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[1]$_SDFF_PN0__520  (.L_HI(net520));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[20]$_DFF_P__521  (.L_HI(net521));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[21]$_DFF_P__522  (.L_HI(net522));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[22]$_DFF_P__523  (.L_HI(net523));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[23]$_DFF_P__524  (.L_HI(net524));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[24]$_DFF_P__525  (.L_HI(net525));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[25]$_DFF_P__526  (.L_HI(net526));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[26]$_DFF_P__527  (.L_HI(net527));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[27]$_DFF_P__528  (.L_HI(net528));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[28]$_DFF_P__529  (.L_HI(net529));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[29]$_DFF_P__530  (.L_HI(net530));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[2]$_SDFF_PN0__531  (.L_HI(net531));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[30]$_DFF_P__532  (.L_HI(net532));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[31]$_DFF_P__533  (.L_HI(net533));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[3]$_SDFF_PN0__534  (.L_HI(net534));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[4]$_DFF_P__535  (.L_HI(net535));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[5]$_DFF_P__536  (.L_HI(net536));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[6]$_DFF_P__537  (.L_HI(net537));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[7]$_DFF_P__538  (.L_HI(net538));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[8]$_DFF_P__539  (.L_HI(net539));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_cycles.register[9]$_DFF_P__540  (.L_HI(net540));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.cy$_SDFF_PN0__541  (.L_HI(net541));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[0]$_SDFF_PN0__542  (.L_HI(net542));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[10]$_DFF_P__543  (.L_HI(net543));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[11]$_DFF_P__544  (.L_HI(net544));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[12]$_DFF_P__545  (.L_HI(net545));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[13]$_DFF_P__546  (.L_HI(net546));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[14]$_DFF_P__547  (.L_HI(net547));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[15]$_DFF_P__548  (.L_HI(net548));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[16]$_DFF_P__549  (.L_HI(net549));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[17]$_DFF_P__550  (.L_HI(net550));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[18]$_DFF_P__551  (.L_HI(net551));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[19]$_DFF_P__552  (.L_HI(net552));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[1]$_SDFF_PN0__553  (.L_HI(net553));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[20]$_DFF_P__554  (.L_HI(net554));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[21]$_DFF_P__555  (.L_HI(net555));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[22]$_DFF_P__556  (.L_HI(net556));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[23]$_DFF_P__557  (.L_HI(net557));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[24]$_DFF_P__558  (.L_HI(net558));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[25]$_DFF_P__559  (.L_HI(net559));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[26]$_DFF_P__560  (.L_HI(net560));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[27]$_DFF_P__561  (.L_HI(net561));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[28]$_DFF_P__562  (.L_HI(net562));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[29]$_DFF_P__563  (.L_HI(net563));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[2]$_SDFF_PN0__564  (.L_HI(net564));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[30]$_DFF_P__565  (.L_HI(net565));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[31]$_DFF_P__566  (.L_HI(net566));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[3]$_SDFF_PN0__567  (.L_HI(net567));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[4]$_DFF_P__568  (.L_HI(net568));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[5]$_DFF_P__569  (.L_HI(net569));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[6]$_DFF_P__570  (.L_HI(net570));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[7]$_DFF_P__571  (.L_HI(net571));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[8]$_DFF_P__572  (.L_HI(net572));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_instrret.register[9]$_DFF_P__573  (.L_HI(net573));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][0]$_DFF_P__574  (.L_HI(net574));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][10]$_DFF_P__575  (.L_HI(net575));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][11]$_DFF_P__576  (.L_HI(net576));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][12]$_DFF_P__577  (.L_HI(net577));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][13]$_DFF_P__578  (.L_HI(net578));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][14]$_DFF_P__579  (.L_HI(net579));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][15]$_DFF_P__580  (.L_HI(net580));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][16]$_DFF_P__581  (.L_HI(net581));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][17]$_DFF_P__582  (.L_HI(net582));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][18]$_DFF_P__583  (.L_HI(net583));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][19]$_DFF_P__584  (.L_HI(net584));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][1]$_DFF_P__585  (.L_HI(net585));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][20]$_DFF_P__586  (.L_HI(net586));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][21]$_DFF_P__587  (.L_HI(net587));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][22]$_DFF_P__588  (.L_HI(net588));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][23]$_DFF_P__589  (.L_HI(net589));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][24]$_DFF_P__590  (.L_HI(net590));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][25]$_DFF_P__591  (.L_HI(net591));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][26]$_DFF_P__592  (.L_HI(net592));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][27]$_DFF_P__593  (.L_HI(net593));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][28]$_DFF_P__594  (.L_HI(net594));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][29]$_DFF_P__595  (.L_HI(net595));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][2]$_DFF_P__596  (.L_HI(net596));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][30]$_DFF_P__597  (.L_HI(net597));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][31]$_DFF_P__598  (.L_HI(net598));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][3]$_DFF_P__599  (.L_HI(net599));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][4]$_DFF_P__600  (.L_HI(net600));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][5]$_DFF_P__601  (.L_HI(net601));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][6]$_DFF_P__602  (.L_HI(net602));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][7]$_DFF_P__603  (.L_HI(net603));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][8]$_DFF_P__604  (.L_HI(net604));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[10][9]$_DFF_P__605  (.L_HI(net605));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][0]$_DFF_P__606  (.L_HI(net606));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][10]$_DFF_P__607  (.L_HI(net607));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][11]$_DFF_P__608  (.L_HI(net608));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][12]$_DFF_P__609  (.L_HI(net609));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][13]$_DFF_P__610  (.L_HI(net610));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][14]$_DFF_P__611  (.L_HI(net611));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][15]$_DFF_P__612  (.L_HI(net612));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][16]$_DFF_P__613  (.L_HI(net613));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][17]$_DFF_P__614  (.L_HI(net614));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][18]$_DFF_P__615  (.L_HI(net615));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][19]$_DFF_P__616  (.L_HI(net616));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][1]$_DFF_P__617  (.L_HI(net617));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][20]$_DFF_P__618  (.L_HI(net618));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][21]$_DFF_P__619  (.L_HI(net619));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][22]$_DFF_P__620  (.L_HI(net620));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][23]$_DFF_P__621  (.L_HI(net621));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][24]$_DFF_P__622  (.L_HI(net622));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][25]$_DFF_P__623  (.L_HI(net623));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][26]$_DFF_P__624  (.L_HI(net624));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][27]$_DFF_P__625  (.L_HI(net625));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][28]$_DFF_P__626  (.L_HI(net626));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][29]$_DFF_P__627  (.L_HI(net627));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][2]$_DFF_P__628  (.L_HI(net628));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][30]$_DFF_P__629  (.L_HI(net629));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][31]$_DFF_P__630  (.L_HI(net630));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][3]$_DFF_P__631  (.L_HI(net631));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][4]$_DFF_P__632  (.L_HI(net632));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][5]$_DFF_P__633  (.L_HI(net633));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][6]$_DFF_P__634  (.L_HI(net634));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][7]$_DFF_P__635  (.L_HI(net635));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][8]$_DFF_P__636  (.L_HI(net636));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[11][9]$_DFF_P__637  (.L_HI(net637));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][0]$_DFF_P__638  (.L_HI(net638));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][10]$_DFF_P__639  (.L_HI(net639));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][11]$_DFF_P__640  (.L_HI(net640));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][12]$_DFF_P__641  (.L_HI(net641));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][13]$_DFF_P__642  (.L_HI(net642));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][14]$_DFF_P__643  (.L_HI(net643));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][15]$_DFF_P__644  (.L_HI(net644));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][16]$_DFF_P__645  (.L_HI(net645));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][17]$_DFF_P__646  (.L_HI(net646));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][18]$_DFF_P__647  (.L_HI(net647));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][19]$_DFF_P__648  (.L_HI(net648));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][1]$_DFF_P__649  (.L_HI(net649));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][20]$_DFF_P__650  (.L_HI(net650));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][21]$_DFF_P__651  (.L_HI(net651));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][22]$_DFF_P__652  (.L_HI(net652));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][23]$_DFF_P__653  (.L_HI(net653));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][24]$_DFF_P__654  (.L_HI(net654));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][25]$_DFF_P__655  (.L_HI(net655));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][26]$_DFF_P__656  (.L_HI(net656));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][27]$_DFF_P__657  (.L_HI(net657));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][28]$_DFF_P__658  (.L_HI(net658));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][29]$_DFF_P__659  (.L_HI(net659));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][2]$_DFF_P__660  (.L_HI(net660));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][30]$_DFF_P__661  (.L_HI(net661));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][31]$_DFF_P__662  (.L_HI(net662));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][3]$_DFF_P__663  (.L_HI(net663));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][4]$_DFF_P__664  (.L_HI(net664));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][5]$_DFF_P__665  (.L_HI(net665));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][6]$_DFF_P__666  (.L_HI(net666));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][7]$_DFF_P__667  (.L_HI(net667));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][8]$_DFF_P__668  (.L_HI(net668));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[12][9]$_DFF_P__669  (.L_HI(net669));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][0]$_DFF_P__670  (.L_HI(net670));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][10]$_DFF_P__671  (.L_HI(net671));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][11]$_DFF_P__672  (.L_HI(net672));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][12]$_DFF_P__673  (.L_HI(net673));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][13]$_DFF_P__674  (.L_HI(net674));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][14]$_DFF_P__675  (.L_HI(net675));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][15]$_DFF_P__676  (.L_HI(net676));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][16]$_DFF_P__677  (.L_HI(net677));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][17]$_DFF_P__678  (.L_HI(net678));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][18]$_DFF_P__679  (.L_HI(net679));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][19]$_DFF_P__680  (.L_HI(net680));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][1]$_DFF_P__681  (.L_HI(net681));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][20]$_DFF_P__682  (.L_HI(net682));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][21]$_DFF_P__683  (.L_HI(net683));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][22]$_DFF_P__684  (.L_HI(net684));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][23]$_DFF_P__685  (.L_HI(net685));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][24]$_DFF_P__686  (.L_HI(net686));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][25]$_DFF_P__687  (.L_HI(net687));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][26]$_DFF_P__688  (.L_HI(net688));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][27]$_DFF_P__689  (.L_HI(net689));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][28]$_DFF_P__690  (.L_HI(net690));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][29]$_DFF_P__691  (.L_HI(net691));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][2]$_DFF_P__692  (.L_HI(net692));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][30]$_DFF_P__693  (.L_HI(net693));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][31]$_DFF_P__694  (.L_HI(net694));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][3]$_DFF_P__695  (.L_HI(net695));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][4]$_DFF_P__696  (.L_HI(net696));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][5]$_DFF_P__697  (.L_HI(net697));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][6]$_DFF_P__698  (.L_HI(net698));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][7]$_DFF_P__699  (.L_HI(net699));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][8]$_DFF_P__700  (.L_HI(net700));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[13][9]$_DFF_P__701  (.L_HI(net701));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][0]$_DFF_P__702  (.L_HI(net702));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][10]$_DFF_P__703  (.L_HI(net703));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][11]$_DFF_P__704  (.L_HI(net704));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][12]$_DFF_P__705  (.L_HI(net705));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][13]$_DFF_P__706  (.L_HI(net706));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][14]$_DFF_P__707  (.L_HI(net707));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][15]$_DFF_P__708  (.L_HI(net708));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][16]$_DFF_P__709  (.L_HI(net709));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][17]$_DFF_P__710  (.L_HI(net710));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][18]$_DFF_P__711  (.L_HI(net711));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][19]$_DFF_P__712  (.L_HI(net712));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][1]$_DFF_P__713  (.L_HI(net713));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][20]$_DFF_P__714  (.L_HI(net714));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][21]$_DFF_P__715  (.L_HI(net715));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][22]$_DFF_P__716  (.L_HI(net716));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][23]$_DFF_P__717  (.L_HI(net717));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][24]$_DFF_P__718  (.L_HI(net718));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][25]$_DFF_P__719  (.L_HI(net719));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][26]$_DFF_P__720  (.L_HI(net720));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][27]$_DFF_P__721  (.L_HI(net721));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][28]$_DFF_P__722  (.L_HI(net722));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][29]$_DFF_P__723  (.L_HI(net723));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][2]$_DFF_P__724  (.L_HI(net724));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][30]$_DFF_P__725  (.L_HI(net725));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][31]$_DFF_P__726  (.L_HI(net726));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][3]$_DFF_P__727  (.L_HI(net727));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][4]$_DFF_P__728  (.L_HI(net728));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][5]$_DFF_P__729  (.L_HI(net729));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][6]$_DFF_P__730  (.L_HI(net730));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][7]$_DFF_P__731  (.L_HI(net731));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][8]$_DFF_P__732  (.L_HI(net732));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[14][9]$_DFF_P__733  (.L_HI(net733));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][0]$_DFF_P__734  (.L_HI(net734));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][10]$_DFF_P__735  (.L_HI(net735));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][11]$_DFF_P__736  (.L_HI(net736));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][12]$_DFF_P__737  (.L_HI(net737));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][13]$_DFF_P__738  (.L_HI(net738));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][14]$_DFF_P__739  (.L_HI(net739));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][15]$_DFF_P__740  (.L_HI(net740));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][16]$_DFF_P__741  (.L_HI(net741));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][17]$_DFF_P__742  (.L_HI(net742));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][18]$_DFF_P__743  (.L_HI(net743));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][19]$_DFF_P__744  (.L_HI(net744));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][1]$_DFF_P__745  (.L_HI(net745));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][20]$_DFF_P__746  (.L_HI(net746));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][21]$_DFF_P__747  (.L_HI(net747));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][22]$_DFF_P__748  (.L_HI(net748));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][23]$_DFF_P__749  (.L_HI(net749));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][24]$_DFF_P__750  (.L_HI(net750));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][25]$_DFF_P__751  (.L_HI(net751));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][26]$_DFF_P__752  (.L_HI(net752));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][27]$_DFF_P__753  (.L_HI(net753));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][28]$_DFF_P__754  (.L_HI(net754));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][29]$_DFF_P__755  (.L_HI(net755));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][2]$_DFF_P__756  (.L_HI(net756));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][30]$_DFF_P__757  (.L_HI(net757));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][31]$_DFF_P__758  (.L_HI(net758));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][3]$_DFF_P__759  (.L_HI(net759));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][4]$_DFF_P__760  (.L_HI(net760));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][5]$_DFF_P__761  (.L_HI(net761));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][6]$_DFF_P__762  (.L_HI(net762));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][7]$_DFF_P__763  (.L_HI(net763));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][8]$_DFF_P__764  (.L_HI(net764));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[15][9]$_DFF_P__765  (.L_HI(net765));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][0]$_DFF_P__766  (.L_HI(net766));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][10]$_DFF_P__767  (.L_HI(net767));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][11]$_DFF_P__768  (.L_HI(net768));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][12]$_DFF_P__769  (.L_HI(net769));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][13]$_DFF_P__770  (.L_HI(net770));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][14]$_DFF_P__771  (.L_HI(net771));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][15]$_DFF_P__772  (.L_HI(net772));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][16]$_DFF_P__773  (.L_HI(net773));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][17]$_DFF_P__774  (.L_HI(net774));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][18]$_DFF_P__775  (.L_HI(net775));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][19]$_DFF_P__776  (.L_HI(net776));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][1]$_DFF_P__777  (.L_HI(net777));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][20]$_DFF_P__778  (.L_HI(net778));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][21]$_DFF_P__779  (.L_HI(net779));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][22]$_DFF_P__780  (.L_HI(net780));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][23]$_DFF_P__781  (.L_HI(net781));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][24]$_DFF_P__782  (.L_HI(net782));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][25]$_DFF_P__783  (.L_HI(net783));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][26]$_DFF_P__784  (.L_HI(net784));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][27]$_DFF_P__785  (.L_HI(net785));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][28]$_DFF_P__786  (.L_HI(net786));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][29]$_DFF_P__787  (.L_HI(net787));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][2]$_DFF_P__788  (.L_HI(net788));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][30]$_DFF_P__789  (.L_HI(net789));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][31]$_DFF_P__790  (.L_HI(net790));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][3]$_DFF_P__791  (.L_HI(net791));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][4]$_DFF_P__792  (.L_HI(net792));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][5]$_DFF_P__793  (.L_HI(net793));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][6]$_DFF_P__794  (.L_HI(net794));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][7]$_DFF_P__795  (.L_HI(net795));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][8]$_DFF_P__796  (.L_HI(net796));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[1][9]$_DFF_P__797  (.L_HI(net797));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][0]$_DFF_P__798  (.L_HI(net798));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][10]$_DFF_P__799  (.L_HI(net799));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][11]$_DFF_P__800  (.L_HI(net800));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][12]$_DFF_P__801  (.L_HI(net801));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][13]$_DFF_P__802  (.L_HI(net802));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][14]$_DFF_P__803  (.L_HI(net803));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][15]$_DFF_P__804  (.L_HI(net804));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][16]$_DFF_P__805  (.L_HI(net805));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][17]$_DFF_P__806  (.L_HI(net806));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][18]$_DFF_P__807  (.L_HI(net807));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][19]$_DFF_P__808  (.L_HI(net808));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][1]$_DFF_P__809  (.L_HI(net809));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][20]$_DFF_P__810  (.L_HI(net810));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][21]$_DFF_P__811  (.L_HI(net811));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][22]$_DFF_P__812  (.L_HI(net812));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][23]$_DFF_P__813  (.L_HI(net813));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][24]$_DFF_P__814  (.L_HI(net814));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][25]$_DFF_P__815  (.L_HI(net815));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][26]$_DFF_P__816  (.L_HI(net816));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][27]$_DFF_P__817  (.L_HI(net817));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][28]$_DFF_P__818  (.L_HI(net818));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][29]$_DFF_P__819  (.L_HI(net819));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][2]$_DFF_P__820  (.L_HI(net820));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][30]$_DFF_P__821  (.L_HI(net821));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][31]$_DFF_P__822  (.L_HI(net822));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][3]$_DFF_P__823  (.L_HI(net823));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][4]$_DFF_P__824  (.L_HI(net824));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][5]$_DFF_P__825  (.L_HI(net825));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][6]$_DFF_P__826  (.L_HI(net826));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][7]$_DFF_P__827  (.L_HI(net827));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][8]$_DFF_P__828  (.L_HI(net828));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[2][9]$_DFF_P__829  (.L_HI(net829));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][0]$_DFF_P__830  (.L_HI(net830));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][10]$_DFF_P__831  (.L_HI(net831));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][11]$_DFF_P__832  (.L_HI(net832));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][12]$_DFF_P__833  (.L_HI(net833));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][13]$_DFF_P__834  (.L_HI(net834));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][14]$_DFF_P__835  (.L_HI(net835));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][15]$_DFF_P__836  (.L_HI(net836));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][16]$_DFF_P__837  (.L_HI(net837));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][17]$_DFF_P__838  (.L_HI(net838));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][18]$_DFF_P__839  (.L_HI(net839));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][19]$_DFF_P__840  (.L_HI(net840));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][1]$_DFF_P__841  (.L_HI(net841));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][20]$_DFF_P__842  (.L_HI(net842));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][21]$_DFF_P__843  (.L_HI(net843));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][22]$_DFF_P__844  (.L_HI(net844));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][23]$_DFF_P__845  (.L_HI(net845));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][24]$_DFF_P__846  (.L_HI(net846));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][25]$_DFF_P__847  (.L_HI(net847));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][26]$_DFF_P__848  (.L_HI(net848));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][27]$_DFF_P__849  (.L_HI(net849));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][28]$_DFF_P__850  (.L_HI(net850));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][29]$_DFF_P__851  (.L_HI(net851));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][2]$_DFF_P__852  (.L_HI(net852));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][30]$_DFF_P__853  (.L_HI(net853));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][31]$_DFF_P__854  (.L_HI(net854));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][3]$_DFF_P__855  (.L_HI(net855));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][4]$_DFF_P__856  (.L_HI(net856));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][5]$_DFF_P__857  (.L_HI(net857));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][6]$_DFF_P__858  (.L_HI(net858));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][7]$_DFF_P__859  (.L_HI(net859));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][8]$_DFF_P__860  (.L_HI(net860));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[5][9]$_DFF_P__861  (.L_HI(net861));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][0]$_DFF_P__862  (.L_HI(net862));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][10]$_DFF_P__863  (.L_HI(net863));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][11]$_DFF_P__864  (.L_HI(net864));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][12]$_DFF_P__865  (.L_HI(net865));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][13]$_DFF_P__866  (.L_HI(net866));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][14]$_DFF_P__867  (.L_HI(net867));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][15]$_DFF_P__868  (.L_HI(net868));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][16]$_DFF_P__869  (.L_HI(net869));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][17]$_DFF_P__870  (.L_HI(net870));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][18]$_DFF_P__871  (.L_HI(net871));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][19]$_DFF_P__872  (.L_HI(net872));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][1]$_DFF_P__873  (.L_HI(net873));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][20]$_DFF_P__874  (.L_HI(net874));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][21]$_DFF_P__875  (.L_HI(net875));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][22]$_DFF_P__876  (.L_HI(net876));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][23]$_DFF_P__877  (.L_HI(net877));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][24]$_DFF_P__878  (.L_HI(net878));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][25]$_DFF_P__879  (.L_HI(net879));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][26]$_DFF_P__880  (.L_HI(net880));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][27]$_DFF_P__881  (.L_HI(net881));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][28]$_DFF_P__882  (.L_HI(net882));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][29]$_DFF_P__883  (.L_HI(net883));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][2]$_DFF_P__884  (.L_HI(net884));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][30]$_DFF_P__885  (.L_HI(net885));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][31]$_DFF_P__886  (.L_HI(net886));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][3]$_DFF_P__887  (.L_HI(net887));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][4]$_DFF_P__888  (.L_HI(net888));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][5]$_DFF_P__889  (.L_HI(net889));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][6]$_DFF_P__890  (.L_HI(net890));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][7]$_DFF_P__891  (.L_HI(net891));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][8]$_DFF_P__892  (.L_HI(net892));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[6][9]$_DFF_P__893  (.L_HI(net893));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][0]$_DFF_P__894  (.L_HI(net894));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][10]$_DFF_P__895  (.L_HI(net895));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][11]$_DFF_P__896  (.L_HI(net896));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][12]$_DFF_P__897  (.L_HI(net897));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][13]$_DFF_P__898  (.L_HI(net898));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][14]$_DFF_P__899  (.L_HI(net899));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][15]$_DFF_P__900  (.L_HI(net900));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][16]$_DFF_P__901  (.L_HI(net901));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][17]$_DFF_P__902  (.L_HI(net902));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][18]$_DFF_P__903  (.L_HI(net903));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][19]$_DFF_P__904  (.L_HI(net904));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][1]$_DFF_P__905  (.L_HI(net905));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][20]$_DFF_P__906  (.L_HI(net906));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][21]$_DFF_P__907  (.L_HI(net907));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][22]$_DFF_P__908  (.L_HI(net908));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][23]$_DFF_P__909  (.L_HI(net909));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][24]$_DFF_P__910  (.L_HI(net910));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][25]$_DFF_P__911  (.L_HI(net911));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][26]$_DFF_P__912  (.L_HI(net912));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][27]$_DFF_P__913  (.L_HI(net913));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][28]$_DFF_P__914  (.L_HI(net914));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][29]$_DFF_P__915  (.L_HI(net915));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][2]$_DFF_P__916  (.L_HI(net916));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][30]$_DFF_P__917  (.L_HI(net917));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][31]$_DFF_P__918  (.L_HI(net918));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][3]$_DFF_P__919  (.L_HI(net919));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][4]$_DFF_P__920  (.L_HI(net920));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][5]$_DFF_P__921  (.L_HI(net921));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][6]$_DFF_P__922  (.L_HI(net922));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][7]$_DFF_P__923  (.L_HI(net923));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][8]$_DFF_P__924  (.L_HI(net924));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[7][9]$_DFF_P__925  (.L_HI(net925));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][0]$_DFF_P__926  (.L_HI(net926));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][10]$_DFF_P__927  (.L_HI(net927));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][11]$_DFF_P__928  (.L_HI(net928));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][12]$_DFF_P__929  (.L_HI(net929));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][13]$_DFF_P__930  (.L_HI(net930));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][14]$_DFF_P__931  (.L_HI(net931));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][15]$_DFF_P__932  (.L_HI(net932));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][16]$_DFF_P__933  (.L_HI(net933));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][17]$_DFF_P__934  (.L_HI(net934));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][18]$_DFF_P__935  (.L_HI(net935));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][19]$_DFF_P__936  (.L_HI(net936));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][1]$_DFF_P__937  (.L_HI(net937));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][20]$_DFF_P__938  (.L_HI(net938));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][21]$_DFF_P__939  (.L_HI(net939));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][22]$_DFF_P__940  (.L_HI(net940));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][23]$_DFF_P__941  (.L_HI(net941));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][24]$_DFF_P__942  (.L_HI(net942));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][25]$_DFF_P__943  (.L_HI(net943));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][26]$_DFF_P__944  (.L_HI(net944));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][27]$_DFF_P__945  (.L_HI(net945));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][28]$_DFF_P__946  (.L_HI(net946));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][29]$_DFF_P__947  (.L_HI(net947));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][2]$_DFF_P__948  (.L_HI(net948));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][30]$_DFF_P__949  (.L_HI(net949));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][31]$_DFF_P__950  (.L_HI(net950));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][3]$_DFF_P__951  (.L_HI(net951));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][4]$_DFF_P__952  (.L_HI(net952));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][5]$_DFF_P__953  (.L_HI(net953));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][6]$_DFF_P__954  (.L_HI(net954));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][7]$_DFF_P__955  (.L_HI(net955));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][8]$_DFF_P__956  (.L_HI(net956));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[8][9]$_DFF_P__957  (.L_HI(net957));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][0]$_DFF_P__958  (.L_HI(net958));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][10]$_DFF_P__959  (.L_HI(net959));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][11]$_DFF_P__960  (.L_HI(net960));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][12]$_DFF_P__961  (.L_HI(net961));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][13]$_DFF_P__962  (.L_HI(net962));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][14]$_DFF_P__963  (.L_HI(net963));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][15]$_DFF_P__964  (.L_HI(net964));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][16]$_DFF_P__965  (.L_HI(net965));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][17]$_DFF_P__966  (.L_HI(net966));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][18]$_DFF_P__967  (.L_HI(net967));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][19]$_DFF_P__968  (.L_HI(net968));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][1]$_DFF_P__969  (.L_HI(net969));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][20]$_DFF_P__970  (.L_HI(net970));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][21]$_DFF_P__971  (.L_HI(net971));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][22]$_DFF_P__972  (.L_HI(net972));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][23]$_DFF_P__973  (.L_HI(net973));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][24]$_DFF_P__974  (.L_HI(net974));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][25]$_DFF_P__975  (.L_HI(net975));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][26]$_DFF_P__976  (.L_HI(net976));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][27]$_DFF_P__977  (.L_HI(net977));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][28]$_DFF_P__978  (.L_HI(net978));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][29]$_DFF_P__979  (.L_HI(net979));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][2]$_DFF_P__980  (.L_HI(net980));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][30]$_DFF_P__981  (.L_HI(net981));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][31]$_DFF_P__982  (.L_HI(net982));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][3]$_DFF_P__983  (.L_HI(net983));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][4]$_DFF_P__984  (.L_HI(net984));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][5]$_DFF_P__985  (.L_HI(net985));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][6]$_DFF_P__986  (.L_HI(net986));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][7]$_DFF_P__987  (.L_HI(net987));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][8]$_DFF_P__988  (.L_HI(net988));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.i_registers.registers[9][9]$_DFF_P__989  (.L_HI(net989));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.instr_retired$_DFF_P__990  (.L_HI(net990));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.is_double_fault_r$_DFFE_PP__991  (.L_HI(net991));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.last_interrupt_req[0]$_DFFE_PP__992  (.L_HI(net992));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.last_interrupt_req[1]$_DFFE_PP__993  (.L_HI(net993));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.load_done$_DFFE_PP__994  (.L_HI(net994));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.load_top_bit$_SDFFCE_PN0P__995  (.L_HI(net995));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mcause[0]$_SDFFE_PN0P__996  (.L_HI(net996));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mcause[1]$_SDFFE_PN0P__997  (.L_HI(net997));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mcause[3]$_SDFFE_PN0P__998  (.L_HI(net998));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mcause[4]$_SDFFE_PN0P__999  (.L_HI(net999));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[0]$_DFFE_PN__1000  (.L_HI(net1000));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[10]$_DFFE_PN__1001  (.L_HI(net1001));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[11]$_DFFE_PN__1002  (.L_HI(net1002));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[12]$_DFFE_PN__1003  (.L_HI(net1003));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[13]$_DFFE_PN__1004  (.L_HI(net1004));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[14]$_DFFE_PN__1005  (.L_HI(net1005));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[15]$_DFFE_PN__1006  (.L_HI(net1006));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[16]$_DFFE_PN__1007  (.L_HI(net1007));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[17]$_DFFE_PN__1008  (.L_HI(net1008));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[18]$_DFFE_PN__1009  (.L_HI(net1009));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[19]$_DFFE_PN__1010  (.L_HI(net1010));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[1]$_DFFE_PN__1011  (.L_HI(net1011));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[20]$_SDFFCE_PN0N__1012  (.L_HI(net1012));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[21]$_SDFFCE_PN0N__1013  (.L_HI(net1013));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[22]$_SDFFCE_PN0N__1014  (.L_HI(net1014));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[23]$_SDFFCE_PN0N__1015  (.L_HI(net1015));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[2]$_DFFE_PN__1016  (.L_HI(net1016));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[3]$_DFFE_PN__1017  (.L_HI(net1017));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[4]$_DFFE_PN__1018  (.L_HI(net1018));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[5]$_DFFE_PN__1019  (.L_HI(net1019));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[6]$_DFFE_PN__1020  (.L_HI(net1020));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[7]$_DFFE_PN__1021  (.L_HI(net1021));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[8]$_DFFE_PN__1022  (.L_HI(net1022));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mepc[9]$_DFFE_PN__1023  (.L_HI(net1023));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mstatus_mie$_SDFFE_PP1P__1024  (.L_HI(net1024));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mstatus_mpie$_SDFFE_PP0P__1025  (.L_HI(net1025));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.mstatus_mte$_SDFFE_PP1P__1026  (.L_HI(net1026));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[0]$_DFF_P__1027  (.L_HI(net1027));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[10]$_DFF_P__1028  (.L_HI(net1028));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[11]$_DFF_P__1029  (.L_HI(net1029));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[12]$_SDFF_PP0__1030  (.L_HI(net1030));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[13]$_SDFF_PP0__1031  (.L_HI(net1031));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[14]$_SDFF_PP0__1032  (.L_HI(net1032));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[15]$_SDFF_PP0__1033  (.L_HI(net1033));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[1]$_DFF_P__1034  (.L_HI(net1034));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[2]$_DFF_P__1035  (.L_HI(net1035));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[3]$_DFF_P__1036  (.L_HI(net1036));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[4]$_DFF_P__1037  (.L_HI(net1037));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[5]$_DFF_P__1038  (.L_HI(net1038));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[6]$_DFF_P__1039  (.L_HI(net1039));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[7]$_DFF_P__1040  (.L_HI(net1040));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[8]$_DFF_P__1041  (.L_HI(net1041));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.multiplier.accum[9]$_DFF_P__1042  (.L_HI(net1042));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[0]$_DFFE_PP__1043  (.L_HI(net1043));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[1]$_DFFE_PP__1044  (.L_HI(net1044));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[2]$_DFFE_PP__1045  (.L_HI(net1045));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[3]$_DFFE_PP__1046  (.L_HI(net1046));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.shift_amt[4]$_DFFE_PP__1047  (.L_HI(net1047));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.time_hi[0]$_SDFFE_PN0P__1048  (.L_HI(net1048));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.time_hi[1]$_SDFFE_PN0P__1049  (.L_HI(net1049));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.time_hi[2]$_SDFFE_PN0P__1050  (.L_HI(net1050));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[0]$_DFFE_PN__1051  (.L_HI(net1051));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[10]$_DFFE_PN__1052  (.L_HI(net1052));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[11]$_DFFE_PN__1053  (.L_HI(net1053));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[12]$_DFFE_PN__1054  (.L_HI(net1054));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[13]$_DFFE_PN__1055  (.L_HI(net1055));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[14]$_DFFE_PN__1056  (.L_HI(net1056));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[15]$_DFFE_PN__1057  (.L_HI(net1057));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[16]$_DFFE_PN__1058  (.L_HI(net1058));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[17]$_DFFE_PN__1059  (.L_HI(net1059));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[18]$_DFFE_PN__1060  (.L_HI(net1060));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[19]$_DFFE_PN__1061  (.L_HI(net1061));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[1]$_DFFE_PN__1062  (.L_HI(net1062));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[20]$_DFFE_PN__1063  (.L_HI(net1063));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[21]$_DFFE_PN__1064  (.L_HI(net1064));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[22]$_DFFE_PN__1065  (.L_HI(net1065));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[23]$_DFFE_PN__1066  (.L_HI(net1066));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[24]$_DFFE_PN__1067  (.L_HI(net1067));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[25]$_DFFE_PN__1068  (.L_HI(net1068));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[26]$_DFFE_PN__1069  (.L_HI(net1069));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[27]$_DFFE_PN__1070  (.L_HI(net1070));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[28]$_SDFFCE_PN0N__1071  (.L_HI(net1071));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[29]$_SDFFCE_PN0N__1072  (.L_HI(net1072));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[2]$_DFFE_PN__1073  (.L_HI(net1073));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[30]$_DFFE_PN__1074  (.L_HI(net1074));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[31]$_DFFE_PN__1075  (.L_HI(net1075));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[3]$_DFFE_PN__1076  (.L_HI(net1076));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[4]$_DFFE_PN__1077  (.L_HI(net1077));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[5]$_DFFE_PN__1078  (.L_HI(net1078));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[6]$_DFFE_PN__1079  (.L_HI(net1079));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[7]$_DFFE_PN__1080  (.L_HI(net1080));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[8]$_DFFE_PN__1081  (.L_HI(net1081));
 sg13g2_tiehi \i_tinyqv.cpu.i_core.tmp_data[9]$_DFFE_PN__1082  (.L_HI(net1082));
 sg13g2_tiehi \i_tinyqv.cpu.imm[0]$_DFFE_PP__1083  (.L_HI(net1083));
 sg13g2_tiehi \i_tinyqv.cpu.imm[10]$_DFFE_PP__1084  (.L_HI(net1084));
 sg13g2_tiehi \i_tinyqv.cpu.imm[11]$_DFFE_PP__1085  (.L_HI(net1085));
 sg13g2_tiehi \i_tinyqv.cpu.imm[12]$_DFFE_PP__1086  (.L_HI(net1086));
 sg13g2_tiehi \i_tinyqv.cpu.imm[13]$_DFFE_PP__1087  (.L_HI(net1087));
 sg13g2_tiehi \i_tinyqv.cpu.imm[14]$_DFFE_PP__1088  (.L_HI(net1088));
 sg13g2_tiehi \i_tinyqv.cpu.imm[15]$_DFFE_PP__1089  (.L_HI(net1089));
 sg13g2_tiehi \i_tinyqv.cpu.imm[16]$_DFFE_PP__1090  (.L_HI(net1090));
 sg13g2_tiehi \i_tinyqv.cpu.imm[17]$_DFFE_PP__1091  (.L_HI(net1091));
 sg13g2_tiehi \i_tinyqv.cpu.imm[18]$_DFFE_PP__1092  (.L_HI(net1092));
 sg13g2_tiehi \i_tinyqv.cpu.imm[19]$_DFFE_PP__1093  (.L_HI(net1093));
 sg13g2_tiehi \i_tinyqv.cpu.imm[1]$_DFFE_PP__1094  (.L_HI(net1094));
 sg13g2_tiehi \i_tinyqv.cpu.imm[20]$_DFFE_PP__1095  (.L_HI(net1095));
 sg13g2_tiehi \i_tinyqv.cpu.imm[21]$_DFFE_PP__1096  (.L_HI(net1096));
 sg13g2_tiehi \i_tinyqv.cpu.imm[22]$_DFFE_PP__1097  (.L_HI(net1097));
 sg13g2_tiehi \i_tinyqv.cpu.imm[23]$_DFFE_PP__1098  (.L_HI(net1098));
 sg13g2_tiehi \i_tinyqv.cpu.imm[24]$_DFFE_PP__1099  (.L_HI(net1099));
 sg13g2_tiehi \i_tinyqv.cpu.imm[25]$_DFFE_PP__1100  (.L_HI(net1100));
 sg13g2_tiehi \i_tinyqv.cpu.imm[26]$_DFFE_PP__1101  (.L_HI(net1101));
 sg13g2_tiehi \i_tinyqv.cpu.imm[27]$_DFFE_PP__1102  (.L_HI(net1102));
 sg13g2_tiehi \i_tinyqv.cpu.imm[28]$_DFFE_PP__1103  (.L_HI(net1103));
 sg13g2_tiehi \i_tinyqv.cpu.imm[29]$_DFFE_PP__1104  (.L_HI(net1104));
 sg13g2_tiehi \i_tinyqv.cpu.imm[2]$_DFFE_PP__1105  (.L_HI(net1105));
 sg13g2_tiehi \i_tinyqv.cpu.imm[30]$_DFFE_PP__1106  (.L_HI(net1106));
 sg13g2_tiehi \i_tinyqv.cpu.imm[31]$_DFFE_PP__1107  (.L_HI(net1107));
 sg13g2_tiehi \i_tinyqv.cpu.imm[3]$_DFFE_PP__1108  (.L_HI(net1108));
 sg13g2_tiehi \i_tinyqv.cpu.imm[4]$_DFFE_PP__1109  (.L_HI(net1109));
 sg13g2_tiehi \i_tinyqv.cpu.imm[5]$_DFFE_PP__1110  (.L_HI(net1110));
 sg13g2_tiehi \i_tinyqv.cpu.imm[6]$_DFFE_PP__1111  (.L_HI(net1111));
 sg13g2_tiehi \i_tinyqv.cpu.imm[7]$_DFFE_PP__1112  (.L_HI(net1112));
 sg13g2_tiehi \i_tinyqv.cpu.imm[8]$_DFFE_PP__1113  (.L_HI(net1113));
 sg13g2_tiehi \i_tinyqv.cpu.imm[9]$_DFFE_PP__1114  (.L_HI(net1114));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][0]$_SDFFCE_PN1P__1115  (.L_HI(net1115));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][10]$_DFFE_PP__1116  (.L_HI(net1116));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][11]$_DFFE_PP__1117  (.L_HI(net1117));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][12]$_DFFE_PP__1118  (.L_HI(net1118));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][13]$_DFFE_PP__1119  (.L_HI(net1119));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][14]$_DFFE_PP__1120  (.L_HI(net1120));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][15]$_DFFE_PP__1121  (.L_HI(net1121));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][1]$_SDFFCE_PN1P__1122  (.L_HI(net1122));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][2]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][3]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][4]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][5]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][6]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][7]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][8]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[0][9]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][0]$_SDFFCE_PN1P__1131  (.L_HI(net1131));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][10]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][11]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][12]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][13]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][14]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][15]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][1]$_SDFFCE_PN1P__1138  (.L_HI(net1138));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][2]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][3]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][4]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][5]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][6]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][7]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][8]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[1][9]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][0]$_SDFFCE_PN1P__1147  (.L_HI(net1147));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][10]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][11]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][12]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][13]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][14]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][15]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][1]$_SDFFCE_PN1P__1154  (.L_HI(net1154));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][2]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][3]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][4]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][5]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][6]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][7]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][8]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[2][9]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][0]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][10]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][11]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][12]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][13]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][14]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][15]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][1]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][2]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][3]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][4]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][5]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][6]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][7]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][8]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data[3][9]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[0]$_SDFFE_PN0P__1179  (.L_HI(net1179));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[10]$_SDFFE_PN0P__1180  (.L_HI(net1180));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[11]$_SDFFE_PN0P__1181  (.L_HI(net1181));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[12]$_SDFFE_PN0P__1182  (.L_HI(net1182));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[13]$_SDFFE_PN0P__1183  (.L_HI(net1183));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[14]$_SDFFE_PN0P__1184  (.L_HI(net1184));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[15]$_SDFFE_PN0P__1185  (.L_HI(net1185));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[16]$_SDFFE_PN0P__1186  (.L_HI(net1186));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[17]$_SDFFE_PN0P__1187  (.L_HI(net1187));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[18]$_SDFFE_PN0P__1188  (.L_HI(net1188));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[19]$_SDFFE_PN0P__1189  (.L_HI(net1189));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[1]$_SDFFE_PN0P__1190  (.L_HI(net1190));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[20]$_SDFFE_PN0P__1191  (.L_HI(net1191));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[2]$_SDFFE_PN0P__1192  (.L_HI(net1192));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[3]$_SDFFE_PN0P__1193  (.L_HI(net1193));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[4]$_SDFFE_PN0P__1194  (.L_HI(net1194));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[5]$_SDFFE_PN0P__1195  (.L_HI(net1195));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[6]$_SDFFE_PN0P__1196  (.L_HI(net1196));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[7]$_SDFFE_PN0P__1197  (.L_HI(net1197));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[8]$_SDFFE_PN0P__1198  (.L_HI(net1198));
 sg13g2_tiehi \i_tinyqv.cpu.instr_data_start[9]$_SDFFE_PN0P__1199  (.L_HI(net1199));
 sg13g2_tiehi \i_tinyqv.cpu.instr_fetch_running$_SDFFE_PN0P__1200  (.L_HI(net1200));
 sg13g2_tiehi \i_tinyqv.cpu.instr_len[0]$_SDFFE_PN0P__1201  (.L_HI(net1201));
 sg13g2_tiehi \i_tinyqv.cpu.instr_len[1]$_SDFFE_PN1P__1202  (.L_HI(net1202));
 sg13g2_tiehi \i_tinyqv.cpu.instr_valid$_SDFFE_PN0P__1203  (.L_HI(net1203));
 sg13g2_tiehi \i_tinyqv.cpu.instr_write_offset[0]$_SDFF_PN0__1204  (.L_HI(net1204));
 sg13g2_tiehi \i_tinyqv.cpu.instr_write_offset[1]$_SDFF_PN0__1205  (.L_HI(net1205));
 sg13g2_tiehi \i_tinyqv.cpu.instr_write_offset[2]$_SDFF_PP0__1206  (.L_HI(net1206));
 sg13g2_tiehi \i_tinyqv.cpu.interrupt_core$_SDFFE_PN0P__1207  (.L_HI(net1207));
 sg13g2_tiehi \i_tinyqv.cpu.is_alu_imm$_SDFFE_PN0P__1208  (.L_HI(net1208));
 sg13g2_tiehi \i_tinyqv.cpu.is_alu_reg$_SDFFE_PN0P__1209  (.L_HI(net1209));
 sg13g2_tiehi \i_tinyqv.cpu.is_auipc$_SDFFE_PN0P__1210  (.L_HI(net1210));
 sg13g2_tiehi \i_tinyqv.cpu.is_branch$_SDFFE_PN0P__1211  (.L_HI(net1211));
 sg13g2_tiehi \i_tinyqv.cpu.is_jal$_SDFFE_PN0P__1212  (.L_HI(net1212));
 sg13g2_tiehi \i_tinyqv.cpu.is_jalr$_SDFFE_PN0P__1213  (.L_HI(net1213));
 sg13g2_tiehi \i_tinyqv.cpu.is_load$_SDFFE_PN0P__1214  (.L_HI(net1214));
 sg13g2_tiehi \i_tinyqv.cpu.is_lui$_SDFFE_PN0P__1215  (.L_HI(net1215));
 sg13g2_tiehi \i_tinyqv.cpu.is_store$_SDFFE_PN0P__1216  (.L_HI(net1216));
 sg13g2_tiehi \i_tinyqv.cpu.is_system$_SDFFE_PN0P__1217  (.L_HI(net1217));
 sg13g2_tiehi \i_tinyqv.cpu.load_started$_SDFFE_PN0P__1218  (.L_HI(net1218));
 sg13g2_tiehi \i_tinyqv.cpu.mem_op[0]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \i_tinyqv.cpu.mem_op[1]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \i_tinyqv.cpu.mem_op[2]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \i_tinyqv.cpu.mem_op_increment_reg$_SDFFCE_PN1P__1222  (.L_HI(net1222));
 sg13g2_tiehi \i_tinyqv.cpu.no_write_in_progress$_SDFFE_PN1P__1223  (.L_HI(net1223));
 sg13g2_tiehi \i_tinyqv.cpu.pc_offset[0]$_SDFFE_PN0P__1224  (.L_HI(net1224));
 sg13g2_tiehi \i_tinyqv.cpu.pc_offset[1]$_SDFFE_PN0P__1225  (.L_HI(net1225));
 sg13g2_tiehi \i_tinyqv.cpu.rd[0]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \i_tinyqv.cpu.rd[1]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \i_tinyqv.cpu.rd[2]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \i_tinyqv.cpu.rd[3]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \i_tinyqv.cpu.rs1[0]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \i_tinyqv.cpu.rs1[1]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \i_tinyqv.cpu.rs1[2]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \i_tinyqv.cpu.rs1[3]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \i_tinyqv.cpu.rs2[0]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \i_tinyqv.cpu.rs2[1]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \i_tinyqv.cpu.rs2[2]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \i_tinyqv.cpu.rs2[3]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \i_tinyqv.cpu.was_early_branch$_SDFFE_PN0P__1238  (.L_HI(net1238));
 sg13g2_tiehi \i_tinyqv.mem.data_stall$_SDFFE_PN0P__1239  (.L_HI(net1239));
 sg13g2_tiehi \i_tinyqv.mem.instr_active$_SDFFE_PP0P__1240  (.L_HI(net1240));
 sg13g2_tiehi \i_tinyqv.mem.instr_fetch_started$_SDFF_PN0__1241  (.L_HI(net1241));
 sg13g2_tiehi \i_tinyqv.mem.instr_fetch_stopped$_SDFF_PN0__1242  (.L_HI(net1242));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[0]$_SDFFCE_PP0P__1243  (.L_HI(net1243));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[10]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[11]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[12]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[13]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[14]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[15]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[16]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[17]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[18]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[19]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[1]$_SDFFCE_PN0P__1254  (.L_HI(net1254));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[20]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[21]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[22]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[23]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[2]$_SDFFCE_PN0P__1259  (.L_HI(net1259));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[3]$_SDFFCE_PN0P__1260  (.L_HI(net1260));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[4]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[5]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[6]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[7]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[8]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.addr[9]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[0]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[1]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[2]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[3]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[4]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[5]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[6]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data[7]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data_ready$_SDFF_PN0__1275  (.L_HI(net1275));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.data_req$_SDFF_PP0__1276  (.L_HI(net1276));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0]$_DFFE_PN__1277  (.L_HI(net1277));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1]$_DFFE_PN__1278  (.L_HI(net1278));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2]$_DFFE_PN__1279  (.L_HI(net1279));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.fsm_state[0]$_SDFFE_PP0P__1280  (.L_HI(net1280));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.fsm_state[1]$_SDFFE_PP0P__1281  (.L_HI(net1281));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.fsm_state[2]$_SDFFE_PP0P__1282  (.L_HI(net1282));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.is_writing$_SDFFE_PP0P__1283  (.L_HI(net1283));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.last_ram_a_sel$_SDFF_PN1__1284  (.L_HI(net1284));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.last_ram_b_sel$_SDFF_PN1__1285  (.L_HI(net1285));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.nibbles_remaining[0]$_SDFFE_PP0P__1286  (.L_HI(net1286));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.nibbles_remaining[1]$_SDFFE_PP0P__1287  (.L_HI(net1287));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.nibbles_remaining[2]$_SDFFE_PP0P__1288  (.L_HI(net1288));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.read_cycles_count[0]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.read_cycles_count[1]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.read_cycles_count[2]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_clk_out$_SDFFE_PP0P__1292  (.L_HI(net1292));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_data_oe[2]$_SDFFE_PP0P__1293  (.L_HI(net1293));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_flash_select$_SDFFE_PP1P__1294  (.L_HI(net1294));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[0]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[1]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[2]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[3]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[4]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[5]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[6]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_in_buffer[7]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_ram_a_select$_SDFFE_PP1P__1303  (.L_HI(net1303));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.spi_ram_b_select$_SDFFE_PP1P__1304  (.L_HI(net1304));
 sg13g2_tiehi \i_tinyqv.mem.q_ctrl.stop_txn_reg$_SDFF_PN0__1305  (.L_HI(net1305));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[0]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[10]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[11]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[12]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[13]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[14]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[15]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[16]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[17]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[18]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[19]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[1]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[20]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[21]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[22]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[23]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[24]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[25]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[26]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[27]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[28]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[29]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[2]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[30]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[31]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[3]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[4]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[5]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[6]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[7]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[8]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_buf[9]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_byte_idx[0]$_SDFFE_PP0N__1338  (.L_HI(net1338));
 sg13g2_tiehi \i_tinyqv.mem.qspi_data_byte_idx[1]$_SDFFE_PP0N__1339  (.L_HI(net1339));
 sg13g2_tiehi \i_tinyqv.mem.qspi_write_done$_DFF_P__1340  (.L_HI(net1340));
 sg13g2_tiehi \i_tinyqv.rst_reg_n$_DFF_P__1341  (.L_HI(net1341));
 sg13g2_tiehi \i_uart_rx.bit_sample$_SDFFE_PN0N__1342  (.L_HI(net1342));
 sg13g2_tiehi \i_uart_rx.cycle_counter[0]$_SDFF_PP0__1343  (.L_HI(net1343));
 sg13g2_tiehi \i_uart_rx.cycle_counter[10]$_SDFF_PP0__1344  (.L_HI(net1344));
 sg13g2_tiehi \i_uart_rx.cycle_counter[1]$_SDFF_PP0__1345  (.L_HI(net1345));
 sg13g2_tiehi \i_uart_rx.cycle_counter[2]$_SDFF_PP0__1346  (.L_HI(net1346));
 sg13g2_tiehi \i_uart_rx.cycle_counter[3]$_SDFF_PP0__1347  (.L_HI(net1347));
 sg13g2_tiehi \i_uart_rx.cycle_counter[4]$_SDFF_PP0__1348  (.L_HI(net1348));
 sg13g2_tiehi \i_uart_rx.cycle_counter[5]$_SDFF_PP0__1349  (.L_HI(net1349));
 sg13g2_tiehi \i_uart_rx.cycle_counter[6]$_SDFF_PP0__1350  (.L_HI(net1350));
 sg13g2_tiehi \i_uart_rx.cycle_counter[7]$_SDFF_PP0__1351  (.L_HI(net1351));
 sg13g2_tiehi \i_uart_rx.cycle_counter[8]$_SDFF_PP0__1352  (.L_HI(net1352));
 sg13g2_tiehi \i_uart_rx.cycle_counter[9]$_SDFF_PP0__1353  (.L_HI(net1353));
 sg13g2_tiehi \i_uart_rx.fsm_state[0]$_SDFFE_PN0P__1354  (.L_HI(net1354));
 sg13g2_tiehi \i_uart_rx.fsm_state[1]$_SDFFE_PN0P__1355  (.L_HI(net1355));
 sg13g2_tiehi \i_uart_rx.fsm_state[2]$_SDFFE_PN0P__1356  (.L_HI(net1356));
 sg13g2_tiehi \i_uart_rx.fsm_state[3]$_SDFFE_PN0P__1357  (.L_HI(net1357));
 sg13g2_tiehi \i_uart_rx.recieved_data[0]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \i_uart_rx.recieved_data[1]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \i_uart_rx.recieved_data[2]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \i_uart_rx.recieved_data[3]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \i_uart_rx.recieved_data[4]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \i_uart_rx.recieved_data[5]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \i_uart_rx.recieved_data[6]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \i_uart_rx.recieved_data[7]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \i_uart_rx.rxd_reg[0]$_SDFF_PN1__1366  (.L_HI(net1366));
 sg13g2_tiehi \i_uart_rx.rxd_reg[1]$_SDFF_PN1__1367  (.L_HI(net1367));
 sg13g2_tiehi \i_uart_rx.uart_rts$_SDFF_PN1__1368  (.L_HI(net1368));
 sg13g2_tiehi \i_uart_tx.cycle_counter[0]$_SDFFE_PP0N__1369  (.L_HI(net1369));
 sg13g2_tiehi \i_uart_tx.cycle_counter[10]$_SDFFE_PP0N__1370  (.L_HI(net1370));
 sg13g2_tiehi \i_uart_tx.cycle_counter[1]$_SDFFE_PP0N__1371  (.L_HI(net1371));
 sg13g2_tiehi \i_uart_tx.cycle_counter[2]$_SDFFE_PP0N__1372  (.L_HI(net1372));
 sg13g2_tiehi \i_uart_tx.cycle_counter[3]$_SDFFE_PP0N__1373  (.L_HI(net1373));
 sg13g2_tiehi \i_uart_tx.cycle_counter[4]$_SDFFE_PP0N__1374  (.L_HI(net1374));
 sg13g2_tiehi \i_uart_tx.cycle_counter[5]$_SDFFE_PP0N__1375  (.L_HI(net1375));
 sg13g2_tiehi \i_uart_tx.cycle_counter[6]$_SDFFE_PP0N__1376  (.L_HI(net1376));
 sg13g2_tiehi \i_uart_tx.cycle_counter[7]$_SDFFE_PP0N__1377  (.L_HI(net1377));
 sg13g2_tiehi \i_uart_tx.cycle_counter[8]$_SDFFE_PP0N__1378  (.L_HI(net1378));
 sg13g2_tiehi \i_uart_tx.cycle_counter[9]$_SDFFE_PP0N__1379  (.L_HI(net1379));
 sg13g2_tiehi \i_uart_tx.data_to_send[0]$_SDFFE_PN0P__1380  (.L_HI(net1380));
 sg13g2_tiehi \i_uart_tx.data_to_send[1]$_SDFFE_PN0P__1381  (.L_HI(net1381));
 sg13g2_tiehi \i_uart_tx.data_to_send[2]$_SDFFE_PN0P__1382  (.L_HI(net1382));
 sg13g2_tiehi \i_uart_tx.data_to_send[3]$_SDFFE_PN0P__1383  (.L_HI(net1383));
 sg13g2_tiehi \i_uart_tx.data_to_send[4]$_SDFFE_PN0P__1384  (.L_HI(net1384));
 sg13g2_tiehi \i_uart_tx.data_to_send[5]$_SDFFE_PN0P__1385  (.L_HI(net1385));
 sg13g2_tiehi \i_uart_tx.data_to_send[6]$_SDFFE_PN0P__1386  (.L_HI(net1386));
 sg13g2_tiehi \i_uart_tx.data_to_send[7]$_SDFFE_PN0P__1387  (.L_HI(net1387));
 sg13g2_tiehi \i_uart_tx.fsm_state[0]$_SDFFE_PN0P__1388  (.L_HI(net1388));
 sg13g2_tiehi \i_uart_tx.fsm_state[1]$_SDFFE_PN0P__1389  (.L_HI(net1389));
 sg13g2_tiehi \i_uart_tx.fsm_state[2]$_SDFFE_PN0P__1390  (.L_HI(net1390));
 sg13g2_tiehi \i_uart_tx.fsm_state[3]$_SDFFE_PN0P__1391  (.L_HI(net1391));
 sg13g2_tiehi \i_uart_tx.txd_reg$_SDFF_PN1__1392  (.L_HI(net1392));
 sg13g2_tiehi \rst_reg_n$_DFF_N__1393  (.L_HI(net1393));
 sg13g2_tiehi \ui_in_reg[0]$_DFF_P__1394  (.L_HI(net1394));
 sg13g2_tiehi \ui_in_reg[1]$_DFF_P__1395  (.L_HI(net1395));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_62_clk (.X(clknet_leaf_62_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_63_clk (.X(clknet_leaf_63_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_64_clk (.X(clknet_leaf_64_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_65_clk (.X(clknet_leaf_65_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_66_clk (.X(clknet_leaf_66_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_67_clk (.X(clknet_leaf_67_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_68_clk (.X(clknet_leaf_68_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_69_clk (.X(clknet_leaf_69_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_70_clk (.X(clknet_leaf_70_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_71_clk (.X(clknet_leaf_71_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_72_clk (.X(clknet_leaf_72_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_73_clk (.X(clknet_leaf_73_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_74_clk (.X(clknet_leaf_74_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_75_clk (.X(clknet_leaf_75_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_76_clk (.X(clknet_leaf_76_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_77_clk (.X(clknet_leaf_77_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_78_clk (.X(clknet_leaf_78_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_79_clk (.X(clknet_leaf_79_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_80_clk (.X(clknet_leaf_80_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_81_clk (.X(clknet_leaf_81_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_82_clk (.X(clknet_leaf_82_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_83_clk (.X(clknet_leaf_83_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_84_clk (.X(clknet_leaf_84_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_85_clk (.X(clknet_leaf_85_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_86_clk (.X(clknet_leaf_86_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_87_clk (.X(clknet_leaf_87_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_88_clk (.X(clknet_leaf_88_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_89_clk (.X(clknet_leaf_89_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_90_clk (.X(clknet_leaf_90_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_91_clk (.X(clknet_leaf_91_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_92_clk (.X(clknet_leaf_92_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_93_clk (.X(clknet_leaf_93_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_94_clk (.X(clknet_leaf_94_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_95_clk (.X(clknet_leaf_95_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_96_clk (.X(clknet_leaf_96_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_97_clk (.X(clknet_leaf_97_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_98_clk (.X(clknet_leaf_98_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_99_clk (.X(clknet_leaf_99_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_100_clk (.X(clknet_leaf_100_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_101_clk (.X(clknet_leaf_101_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_102_clk (.X(clknet_leaf_102_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_103_clk (.X(clknet_leaf_103_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_104_clk (.X(clknet_leaf_104_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_105_clk (.X(clknet_leaf_105_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_106_clk (.X(clknet_leaf_106_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_107_clk (.X(clknet_leaf_107_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_108_clk (.X(clknet_leaf_108_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_109_clk (.X(clknet_leaf_109_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_110_clk (.X(clknet_leaf_110_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_111_clk (.X(clknet_leaf_111_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_112_clk (.X(clknet_leaf_112_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_113_clk (.X(clknet_leaf_113_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_114_clk (.X(clknet_leaf_114_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_115_clk (.X(clknet_leaf_115_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_116_clk (.X(clknet_leaf_116_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_117_clk (.X(clknet_leaf_117_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_118_clk (.X(clknet_leaf_118_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_119_clk (.X(clknet_leaf_119_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_120_clk (.X(clknet_leaf_120_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_121_clk (.X(clknet_leaf_121_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_122_clk (.X(clknet_leaf_122_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_123_clk (.X(clknet_leaf_123_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_124_clk (.X(clknet_leaf_124_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_125_clk (.X(clknet_leaf_125_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_126_clk (.X(clknet_leaf_126_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_127_clk (.X(clknet_leaf_127_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_128_clk (.X(clknet_leaf_128_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_129_clk (.X(clknet_leaf_129_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_130_clk (.X(clknet_leaf_130_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_131_clk (.X(clknet_leaf_131_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_132_clk (.X(clknet_leaf_132_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_133_clk (.X(clknet_leaf_133_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_134_clk (.X(clknet_leaf_134_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_135_clk (.X(clknet_leaf_135_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_136_clk (.X(clknet_leaf_136_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_137_clk (.X(clknet_leaf_137_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_138_clk (.X(clknet_leaf_138_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_139_clk (.X(clknet_leaf_139_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkload6 (.A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkload8 (.A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkload9 (.A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkload10 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkload11 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_139_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_leaf_117_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_118_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_17_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_29_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_21_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_51_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_116_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_85_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_113_clk));
 sg13g2_buf_16 clkload22 (.A(clknet_leaf_111_clk));
 sg13g2_buf_16 clkload23 (.A(clknet_leaf_94_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_95_clk));
 sg13g2_buf_16 clkload25 (.A(clknet_leaf_97_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_87_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_92_clk));
 sg13g2_buf_8 clkload28 (.A(clknet_leaf_93_clk));
 sg13g2_inv_2 clkload29 (.A(clknet_leaf_53_clk));
 sg13g2_buf_8 clkload30 (.A(clknet_leaf_54_clk));
 sg13g2_buf_8 clkload31 (.A(clknet_leaf_56_clk));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_75_clk));
 sg13g2_inv_2 clkload33 (.A(clknet_leaf_82_clk));
 sg13g2_buf_16 clkload34 (.A(clknet_leaf_83_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_70_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00052_));
 sg13g2_antennanp ANTENNA_2 (.A(_00052_));
 sg13g2_antennanp ANTENNA_3 (.A(_00369_));
 sg13g2_antennanp ANTENNA_4 (.A(_00370_));
 sg13g2_antennanp ANTENNA_5 (.A(_04271_));
 sg13g2_antennanp ANTENNA_6 (.A(\debug_rd[3] ));
 sg13g2_antennanp ANTENNA_7 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_antennanp ANTENNA_8 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_antennanp ANTENNA_9 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_antennanp ANTENNA_10 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_antennanp ANTENNA_11 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_antennanp ANTENNA_12 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_antennanp ANTENNA_13 (.A(\i_tinyqv.mem.q_ctrl.addr[21] ));
 sg13g2_antennanp ANTENNA_14 (.A(\i_tinyqv.mem.q_ctrl.addr[21] ));
 sg13g2_antennanp ANTENNA_15 (.A(net12));
 sg13g2_antennanp ANTENNA_16 (.A(_00369_));
 sg13g2_antennanp ANTENNA_17 (.A(_00370_));
 sg13g2_antennanp ANTENNA_18 (.A(_04271_));
 sg13g2_antennanp ANTENNA_19 (.A(\debug_rd[3] ));
 sg13g2_antennanp ANTENNA_20 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_antennanp ANTENNA_21 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_antennanp ANTENNA_22 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_antennanp ANTENNA_23 (.A(net12));
 sg13g2_antennanp ANTENNA_24 (.A(_00369_));
 sg13g2_antennanp ANTENNA_25 (.A(_00370_));
 sg13g2_antennanp ANTENNA_26 (.A(\debug_rd[3] ));
 sg13g2_antennanp ANTENNA_27 (.A(net12));
 sg13g2_antennanp ANTENNA_28 (.A(_00369_));
 sg13g2_antennanp ANTENNA_29 (.A(\debug_rd[3] ));
 sg13g2_antennanp ANTENNA_30 (.A(net12));
 sg13g2_antennanp ANTENNA_31 (.A(_00369_));
 sg13g2_antennanp ANTENNA_32 (.A(\debug_rd[3] ));
 sg13g2_antennanp ANTENNA_33 (.A(net12));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_fill_2 FILLER_0_56 ();
 sg13g2_fill_1 FILLER_0_58 ();
 sg13g2_fill_2 FILLER_0_233 ();
 sg13g2_fill_2 FILLER_0_317 ();
 sg13g2_fill_1 FILLER_0_319 ();
 sg13g2_fill_1 FILLER_0_526 ();
 sg13g2_fill_2 FILLER_0_587 ();
 sg13g2_fill_1 FILLER_0_589 ();
 sg13g2_decap_8 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_663 ();
 sg13g2_decap_8 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_684 ();
 sg13g2_decap_8 FILLER_0_691 ();
 sg13g2_decap_8 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_decap_8 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_719 ();
 sg13g2_decap_8 FILLER_0_726 ();
 sg13g2_decap_8 FILLER_0_733 ();
 sg13g2_decap_8 FILLER_0_740 ();
 sg13g2_decap_8 FILLER_0_747 ();
 sg13g2_decap_8 FILLER_0_754 ();
 sg13g2_decap_8 FILLER_0_761 ();
 sg13g2_decap_8 FILLER_0_768 ();
 sg13g2_decap_8 FILLER_0_775 ();
 sg13g2_decap_8 FILLER_0_782 ();
 sg13g2_decap_8 FILLER_0_789 ();
 sg13g2_decap_8 FILLER_0_796 ();
 sg13g2_decap_8 FILLER_0_803 ();
 sg13g2_decap_8 FILLER_0_810 ();
 sg13g2_decap_8 FILLER_0_817 ();
 sg13g2_decap_8 FILLER_0_824 ();
 sg13g2_decap_8 FILLER_0_831 ();
 sg13g2_decap_8 FILLER_0_838 ();
 sg13g2_decap_8 FILLER_0_845 ();
 sg13g2_decap_8 FILLER_0_852 ();
 sg13g2_decap_8 FILLER_0_859 ();
 sg13g2_decap_8 FILLER_0_866 ();
 sg13g2_decap_4 FILLER_0_873 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_2 FILLER_1_49 ();
 sg13g2_fill_1 FILLER_1_51 ();
 sg13g2_fill_2 FILLER_1_166 ();
 sg13g2_fill_1 FILLER_1_168 ();
 sg13g2_fill_2 FILLER_1_211 ();
 sg13g2_fill_2 FILLER_1_307 ();
 sg13g2_fill_2 FILLER_1_339 ();
 sg13g2_fill_1 FILLER_1_561 ();
 sg13g2_fill_2 FILLER_1_604 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_fill_2 FILLER_1_875 ();
 sg13g2_fill_1 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_fill_1 FILLER_2_49 ();
 sg13g2_fill_2 FILLER_2_156 ();
 sg13g2_fill_1 FILLER_2_278 ();
 sg13g2_fill_2 FILLER_2_309 ();
 sg13g2_fill_1 FILLER_2_311 ();
 sg13g2_fill_1 FILLER_2_342 ();
 sg13g2_fill_2 FILLER_2_353 ();
 sg13g2_fill_2 FILLER_2_397 ();
 sg13g2_fill_1 FILLER_2_399 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_fill_1 FILLER_2_435 ();
 sg13g2_fill_1 FILLER_2_462 ();
 sg13g2_fill_2 FILLER_2_543 ();
 sg13g2_fill_2 FILLER_2_631 ();
 sg13g2_decap_8 FILLER_2_667 ();
 sg13g2_decap_8 FILLER_2_674 ();
 sg13g2_decap_8 FILLER_2_681 ();
 sg13g2_decap_8 FILLER_2_688 ();
 sg13g2_decap_8 FILLER_2_695 ();
 sg13g2_decap_8 FILLER_2_702 ();
 sg13g2_decap_8 FILLER_2_709 ();
 sg13g2_decap_8 FILLER_2_716 ();
 sg13g2_decap_8 FILLER_2_723 ();
 sg13g2_decap_8 FILLER_2_730 ();
 sg13g2_decap_8 FILLER_2_737 ();
 sg13g2_decap_8 FILLER_2_744 ();
 sg13g2_decap_8 FILLER_2_751 ();
 sg13g2_decap_8 FILLER_2_758 ();
 sg13g2_decap_8 FILLER_2_765 ();
 sg13g2_decap_8 FILLER_2_772 ();
 sg13g2_decap_8 FILLER_2_779 ();
 sg13g2_decap_8 FILLER_2_786 ();
 sg13g2_decap_8 FILLER_2_793 ();
 sg13g2_decap_8 FILLER_2_800 ();
 sg13g2_decap_8 FILLER_2_807 ();
 sg13g2_decap_8 FILLER_2_814 ();
 sg13g2_decap_8 FILLER_2_821 ();
 sg13g2_decap_8 FILLER_2_828 ();
 sg13g2_decap_8 FILLER_2_835 ();
 sg13g2_decap_8 FILLER_2_842 ();
 sg13g2_decap_8 FILLER_2_849 ();
 sg13g2_decap_8 FILLER_2_856 ();
 sg13g2_decap_8 FILLER_2_863 ();
 sg13g2_decap_8 FILLER_2_870 ();
 sg13g2_fill_1 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_fill_1 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_141 ();
 sg13g2_fill_2 FILLER_3_202 ();
 sg13g2_fill_1 FILLER_3_204 ();
 sg13g2_fill_2 FILLER_3_327 ();
 sg13g2_fill_1 FILLER_3_329 ();
 sg13g2_fill_2 FILLER_3_446 ();
 sg13g2_fill_2 FILLER_3_552 ();
 sg13g2_fill_1 FILLER_3_580 ();
 sg13g2_fill_2 FILLER_3_607 ();
 sg13g2_fill_2 FILLER_3_639 ();
 sg13g2_decap_8 FILLER_3_675 ();
 sg13g2_decap_8 FILLER_3_682 ();
 sg13g2_decap_8 FILLER_3_689 ();
 sg13g2_decap_8 FILLER_3_696 ();
 sg13g2_decap_8 FILLER_3_703 ();
 sg13g2_decap_8 FILLER_3_710 ();
 sg13g2_decap_8 FILLER_3_717 ();
 sg13g2_decap_8 FILLER_3_724 ();
 sg13g2_decap_8 FILLER_3_731 ();
 sg13g2_decap_8 FILLER_3_738 ();
 sg13g2_decap_8 FILLER_3_745 ();
 sg13g2_decap_8 FILLER_3_752 ();
 sg13g2_decap_8 FILLER_3_759 ();
 sg13g2_decap_8 FILLER_3_766 ();
 sg13g2_decap_8 FILLER_3_773 ();
 sg13g2_decap_8 FILLER_3_780 ();
 sg13g2_decap_8 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_794 ();
 sg13g2_decap_8 FILLER_3_801 ();
 sg13g2_decap_8 FILLER_3_808 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_decap_8 FILLER_3_829 ();
 sg13g2_decap_8 FILLER_3_836 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_850 ();
 sg13g2_decap_8 FILLER_3_857 ();
 sg13g2_decap_8 FILLER_3_864 ();
 sg13g2_decap_8 FILLER_3_871 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_21 ();
 sg13g2_fill_1 FILLER_4_218 ();
 sg13g2_fill_2 FILLER_4_263 ();
 sg13g2_fill_1 FILLER_4_275 ();
 sg13g2_fill_1 FILLER_4_354 ();
 sg13g2_fill_2 FILLER_4_365 ();
 sg13g2_fill_1 FILLER_4_384 ();
 sg13g2_fill_1 FILLER_4_411 ();
 sg13g2_fill_1 FILLER_4_426 ();
 sg13g2_fill_1 FILLER_4_453 ();
 sg13g2_fill_1 FILLER_4_458 ();
 sg13g2_fill_1 FILLER_4_653 ();
 sg13g2_decap_8 FILLER_4_688 ();
 sg13g2_decap_8 FILLER_4_695 ();
 sg13g2_decap_8 FILLER_4_702 ();
 sg13g2_decap_8 FILLER_4_709 ();
 sg13g2_decap_8 FILLER_4_716 ();
 sg13g2_decap_8 FILLER_4_723 ();
 sg13g2_decap_8 FILLER_4_730 ();
 sg13g2_decap_8 FILLER_4_737 ();
 sg13g2_decap_8 FILLER_4_744 ();
 sg13g2_decap_8 FILLER_4_751 ();
 sg13g2_decap_8 FILLER_4_758 ();
 sg13g2_decap_8 FILLER_4_765 ();
 sg13g2_decap_8 FILLER_4_772 ();
 sg13g2_decap_8 FILLER_4_779 ();
 sg13g2_decap_8 FILLER_4_786 ();
 sg13g2_decap_8 FILLER_4_793 ();
 sg13g2_decap_8 FILLER_4_800 ();
 sg13g2_decap_8 FILLER_4_807 ();
 sg13g2_decap_8 FILLER_4_814 ();
 sg13g2_decap_8 FILLER_4_821 ();
 sg13g2_decap_8 FILLER_4_828 ();
 sg13g2_decap_8 FILLER_4_835 ();
 sg13g2_decap_8 FILLER_4_842 ();
 sg13g2_decap_8 FILLER_4_849 ();
 sg13g2_decap_8 FILLER_4_856 ();
 sg13g2_decap_8 FILLER_4_863 ();
 sg13g2_decap_8 FILLER_4_870 ();
 sg13g2_fill_1 FILLER_4_877 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_10 ();
 sg13g2_fill_1 FILLER_5_26 ();
 sg13g2_fill_2 FILLER_5_69 ();
 sg13g2_fill_2 FILLER_5_156 ();
 sg13g2_fill_1 FILLER_5_162 ();
 sg13g2_fill_1 FILLER_5_223 ();
 sg13g2_fill_2 FILLER_5_250 ();
 sg13g2_fill_2 FILLER_5_334 ();
 sg13g2_fill_2 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_436 ();
 sg13g2_fill_2 FILLER_5_441 ();
 sg13g2_fill_2 FILLER_5_503 ();
 sg13g2_fill_1 FILLER_5_505 ();
 sg13g2_fill_2 FILLER_5_558 ();
 sg13g2_fill_2 FILLER_5_598 ();
 sg13g2_decap_8 FILLER_5_704 ();
 sg13g2_decap_8 FILLER_5_711 ();
 sg13g2_decap_8 FILLER_5_718 ();
 sg13g2_decap_8 FILLER_5_725 ();
 sg13g2_decap_8 FILLER_5_732 ();
 sg13g2_decap_8 FILLER_5_739 ();
 sg13g2_decap_8 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_decap_8 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_8 FILLER_5_830 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_decap_8 FILLER_5_865 ();
 sg13g2_decap_4 FILLER_5_872 ();
 sg13g2_fill_2 FILLER_5_876 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_10 ();
 sg13g2_fill_1 FILLER_6_19 ();
 sg13g2_fill_2 FILLER_6_40 ();
 sg13g2_fill_1 FILLER_6_128 ();
 sg13g2_fill_1 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_216 ();
 sg13g2_fill_1 FILLER_6_248 ();
 sg13g2_fill_1 FILLER_6_301 ();
 sg13g2_fill_2 FILLER_6_389 ();
 sg13g2_fill_1 FILLER_6_417 ();
 sg13g2_fill_2 FILLER_6_452 ();
 sg13g2_fill_2 FILLER_6_458 ();
 sg13g2_fill_1 FILLER_6_460 ();
 sg13g2_fill_1 FILLER_6_471 ();
 sg13g2_fill_2 FILLER_6_486 ();
 sg13g2_fill_1 FILLER_6_488 ();
 sg13g2_fill_2 FILLER_6_523 ();
 sg13g2_fill_1 FILLER_6_525 ();
 sg13g2_fill_1 FILLER_6_552 ();
 sg13g2_decap_8 FILLER_6_715 ();
 sg13g2_decap_8 FILLER_6_722 ();
 sg13g2_decap_8 FILLER_6_729 ();
 sg13g2_decap_8 FILLER_6_736 ();
 sg13g2_decap_8 FILLER_6_743 ();
 sg13g2_decap_8 FILLER_6_750 ();
 sg13g2_decap_8 FILLER_6_757 ();
 sg13g2_decap_8 FILLER_6_764 ();
 sg13g2_decap_8 FILLER_6_771 ();
 sg13g2_decap_8 FILLER_6_778 ();
 sg13g2_decap_8 FILLER_6_785 ();
 sg13g2_decap_8 FILLER_6_792 ();
 sg13g2_decap_8 FILLER_6_799 ();
 sg13g2_decap_8 FILLER_6_806 ();
 sg13g2_decap_8 FILLER_6_813 ();
 sg13g2_decap_8 FILLER_6_820 ();
 sg13g2_decap_8 FILLER_6_827 ();
 sg13g2_decap_8 FILLER_6_834 ();
 sg13g2_decap_8 FILLER_6_841 ();
 sg13g2_decap_8 FILLER_6_848 ();
 sg13g2_decap_8 FILLER_6_855 ();
 sg13g2_decap_8 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_869 ();
 sg13g2_fill_2 FILLER_6_876 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_fill_1 FILLER_7_18 ();
 sg13g2_fill_1 FILLER_7_53 ();
 sg13g2_fill_2 FILLER_7_182 ();
 sg13g2_fill_1 FILLER_7_184 ();
 sg13g2_fill_2 FILLER_7_313 ();
 sg13g2_fill_2 FILLER_7_397 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_fill_2 FILLER_7_460 ();
 sg13g2_fill_2 FILLER_7_518 ();
 sg13g2_fill_2 FILLER_7_678 ();
 sg13g2_fill_1 FILLER_7_680 ();
 sg13g2_fill_1 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_fill_2 FILLER_7_875 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_200 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_339 ();
 sg13g2_fill_2 FILLER_8_367 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_1 FILLER_8_375 ();
 sg13g2_fill_2 FILLER_8_380 ();
 sg13g2_fill_1 FILLER_8_382 ();
 sg13g2_fill_2 FILLER_8_465 ();
 sg13g2_fill_2 FILLER_8_487 ();
 sg13g2_fill_1 FILLER_8_649 ();
 sg13g2_decap_8 FILLER_8_750 ();
 sg13g2_decap_8 FILLER_8_757 ();
 sg13g2_decap_8 FILLER_8_764 ();
 sg13g2_decap_8 FILLER_8_771 ();
 sg13g2_decap_8 FILLER_8_778 ();
 sg13g2_decap_8 FILLER_8_785 ();
 sg13g2_decap_8 FILLER_8_792 ();
 sg13g2_decap_8 FILLER_8_799 ();
 sg13g2_decap_8 FILLER_8_806 ();
 sg13g2_decap_8 FILLER_8_813 ();
 sg13g2_decap_8 FILLER_8_820 ();
 sg13g2_decap_8 FILLER_8_827 ();
 sg13g2_decap_8 FILLER_8_834 ();
 sg13g2_decap_8 FILLER_8_841 ();
 sg13g2_decap_8 FILLER_8_848 ();
 sg13g2_decap_8 FILLER_8_855 ();
 sg13g2_decap_8 FILLER_8_862 ();
 sg13g2_decap_8 FILLER_8_869 ();
 sg13g2_fill_2 FILLER_8_876 ();
 sg13g2_fill_2 FILLER_9_30 ();
 sg13g2_fill_1 FILLER_9_32 ();
 sg13g2_fill_2 FILLER_9_94 ();
 sg13g2_fill_1 FILLER_9_96 ();
 sg13g2_fill_1 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_228 ();
 sg13g2_fill_2 FILLER_9_259 ();
 sg13g2_fill_1 FILLER_9_331 ();
 sg13g2_fill_2 FILLER_9_426 ();
 sg13g2_fill_1 FILLER_9_428 ();
 sg13g2_fill_2 FILLER_9_437 ();
 sg13g2_fill_1 FILLER_9_439 ();
 sg13g2_fill_1 FILLER_9_448 ();
 sg13g2_decap_4 FILLER_9_459 ();
 sg13g2_fill_1 FILLER_9_463 ();
 sg13g2_fill_1 FILLER_9_542 ();
 sg13g2_fill_2 FILLER_9_593 ();
 sg13g2_fill_2 FILLER_9_681 ();
 sg13g2_fill_1 FILLER_9_683 ();
 sg13g2_fill_1 FILLER_9_708 ();
 sg13g2_fill_1 FILLER_9_747 ();
 sg13g2_fill_1 FILLER_9_753 ();
 sg13g2_decap_4 FILLER_9_766 ();
 sg13g2_fill_1 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_775 ();
 sg13g2_decap_8 FILLER_9_782 ();
 sg13g2_decap_8 FILLER_9_789 ();
 sg13g2_decap_8 FILLER_9_796 ();
 sg13g2_decap_8 FILLER_9_803 ();
 sg13g2_decap_8 FILLER_9_814 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_decap_8 FILLER_9_828 ();
 sg13g2_decap_8 FILLER_9_835 ();
 sg13g2_decap_8 FILLER_9_842 ();
 sg13g2_decap_8 FILLER_9_849 ();
 sg13g2_decap_8 FILLER_9_856 ();
 sg13g2_decap_8 FILLER_9_863 ();
 sg13g2_decap_8 FILLER_9_870 ();
 sg13g2_fill_1 FILLER_9_877 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_fill_1 FILLER_10_13 ();
 sg13g2_fill_2 FILLER_10_52 ();
 sg13g2_fill_1 FILLER_10_54 ();
 sg13g2_fill_2 FILLER_10_107 ();
 sg13g2_fill_1 FILLER_10_213 ();
 sg13g2_fill_2 FILLER_10_240 ();
 sg13g2_fill_2 FILLER_10_294 ();
 sg13g2_fill_1 FILLER_10_382 ();
 sg13g2_decap_4 FILLER_10_387 ();
 sg13g2_fill_2 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_449 ();
 sg13g2_fill_1 FILLER_10_456 ();
 sg13g2_fill_2 FILLER_10_561 ();
 sg13g2_fill_1 FILLER_10_563 ();
 sg13g2_fill_2 FILLER_10_568 ();
 sg13g2_fill_1 FILLER_10_570 ();
 sg13g2_fill_1 FILLER_10_597 ();
 sg13g2_fill_2 FILLER_10_624 ();
 sg13g2_fill_1 FILLER_10_668 ();
 sg13g2_fill_2 FILLER_10_694 ();
 sg13g2_fill_1 FILLER_10_696 ();
 sg13g2_fill_1 FILLER_10_716 ();
 sg13g2_fill_1 FILLER_10_775 ();
 sg13g2_fill_2 FILLER_10_801 ();
 sg13g2_fill_1 FILLER_10_803 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_8 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_865 ();
 sg13g2_decap_4 FILLER_10_872 ();
 sg13g2_fill_2 FILLER_10_876 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_27 ();
 sg13g2_fill_1 FILLER_11_80 ();
 sg13g2_fill_1 FILLER_11_107 ();
 sg13g2_fill_2 FILLER_11_134 ();
 sg13g2_fill_2 FILLER_11_246 ();
 sg13g2_fill_1 FILLER_11_248 ();
 sg13g2_fill_1 FILLER_11_257 ();
 sg13g2_fill_2 FILLER_11_322 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_fill_2 FILLER_11_442 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_fill_1 FILLER_11_469 ();
 sg13g2_decap_4 FILLER_11_474 ();
 sg13g2_fill_1 FILLER_11_588 ();
 sg13g2_fill_2 FILLER_11_609 ();
 sg13g2_fill_2 FILLER_11_645 ();
 sg13g2_fill_1 FILLER_11_655 ();
 sg13g2_fill_1 FILLER_11_661 ();
 sg13g2_fill_2 FILLER_11_668 ();
 sg13g2_fill_1 FILLER_11_685 ();
 sg13g2_fill_1 FILLER_11_691 ();
 sg13g2_decap_4 FILLER_11_779 ();
 sg13g2_fill_2 FILLER_11_793 ();
 sg13g2_fill_1 FILLER_11_795 ();
 sg13g2_fill_1 FILLER_11_804 ();
 sg13g2_fill_1 FILLER_11_809 ();
 sg13g2_fill_1 FILLER_11_815 ();
 sg13g2_fill_1 FILLER_11_824 ();
 sg13g2_decap_4 FILLER_11_829 ();
 sg13g2_fill_1 FILLER_11_836 ();
 sg13g2_decap_4 FILLER_11_840 ();
 sg13g2_fill_2 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_849 ();
 sg13g2_decap_8 FILLER_11_856 ();
 sg13g2_decap_8 FILLER_11_863 ();
 sg13g2_decap_8 FILLER_11_870 ();
 sg13g2_fill_1 FILLER_11_877 ();
 sg13g2_fill_1 FILLER_12_12 ();
 sg13g2_fill_2 FILLER_12_17 ();
 sg13g2_fill_1 FILLER_12_19 ();
 sg13g2_fill_1 FILLER_12_46 ();
 sg13g2_fill_2 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_185 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_fill_2 FILLER_12_240 ();
 sg13g2_fill_1 FILLER_12_242 ();
 sg13g2_fill_1 FILLER_12_364 ();
 sg13g2_fill_2 FILLER_12_373 ();
 sg13g2_fill_2 FILLER_12_383 ();
 sg13g2_fill_2 FILLER_12_519 ();
 sg13g2_fill_1 FILLER_12_521 ();
 sg13g2_fill_1 FILLER_12_578 ();
 sg13g2_fill_1 FILLER_12_643 ();
 sg13g2_fill_2 FILLER_12_669 ();
 sg13g2_fill_1 FILLER_12_679 ();
 sg13g2_fill_1 FILLER_12_690 ();
 sg13g2_fill_2 FILLER_12_698 ();
 sg13g2_fill_1 FILLER_12_700 ();
 sg13g2_fill_2 FILLER_12_738 ();
 sg13g2_fill_1 FILLER_12_740 ();
 sg13g2_fill_2 FILLER_12_793 ();
 sg13g2_fill_2 FILLER_12_805 ();
 sg13g2_fill_1 FILLER_12_844 ();
 sg13g2_fill_2 FILLER_13_29 ();
 sg13g2_fill_1 FILLER_13_31 ();
 sg13g2_fill_2 FILLER_13_148 ();
 sg13g2_fill_1 FILLER_13_214 ();
 sg13g2_fill_1 FILLER_13_284 ();
 sg13g2_fill_2 FILLER_13_299 ();
 sg13g2_fill_1 FILLER_13_331 ();
 sg13g2_fill_2 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_432 ();
 sg13g2_fill_1 FILLER_13_443 ();
 sg13g2_fill_1 FILLER_13_598 ();
 sg13g2_fill_1 FILLER_13_613 ();
 sg13g2_fill_1 FILLER_13_629 ();
 sg13g2_fill_1 FILLER_13_647 ();
 sg13g2_fill_1 FILLER_13_653 ();
 sg13g2_fill_2 FILLER_13_671 ();
 sg13g2_fill_1 FILLER_13_673 ();
 sg13g2_fill_2 FILLER_13_745 ();
 sg13g2_fill_2 FILLER_13_767 ();
 sg13g2_fill_2 FILLER_13_788 ();
 sg13g2_fill_1 FILLER_13_790 ();
 sg13g2_fill_1 FILLER_13_804 ();
 sg13g2_fill_1 FILLER_13_818 ();
 sg13g2_fill_1 FILLER_13_829 ();
 sg13g2_fill_2 FILLER_13_838 ();
 sg13g2_fill_1 FILLER_14_67 ();
 sg13g2_fill_1 FILLER_14_98 ();
 sg13g2_fill_2 FILLER_14_125 ();
 sg13g2_fill_2 FILLER_14_157 ();
 sg13g2_fill_2 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_fill_1 FILLER_14_451 ();
 sg13g2_fill_2 FILLER_14_456 ();
 sg13g2_fill_1 FILLER_14_462 ();
 sg13g2_fill_2 FILLER_14_467 ();
 sg13g2_fill_1 FILLER_14_495 ();
 sg13g2_fill_2 FILLER_14_500 ();
 sg13g2_fill_1 FILLER_14_506 ();
 sg13g2_fill_2 FILLER_14_625 ();
 sg13g2_fill_2 FILLER_14_656 ();
 sg13g2_fill_1 FILLER_14_687 ();
 sg13g2_fill_2 FILLER_14_701 ();
 sg13g2_fill_1 FILLER_14_703 ();
 sg13g2_fill_1 FILLER_14_712 ();
 sg13g2_fill_1 FILLER_14_738 ();
 sg13g2_fill_1 FILLER_14_747 ();
 sg13g2_fill_1 FILLER_14_761 ();
 sg13g2_fill_1 FILLER_14_770 ();
 sg13g2_fill_1 FILLER_14_781 ();
 sg13g2_fill_2 FILLER_14_795 ();
 sg13g2_fill_1 FILLER_14_797 ();
 sg13g2_decap_8 FILLER_14_802 ();
 sg13g2_fill_1 FILLER_14_839 ();
 sg13g2_fill_1 FILLER_15_16 ();
 sg13g2_fill_1 FILLER_15_73 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_170 ();
 sg13g2_fill_1 FILLER_15_197 ();
 sg13g2_fill_2 FILLER_15_234 ();
 sg13g2_fill_1 FILLER_15_236 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_fill_1 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_338 ();
 sg13g2_fill_1 FILLER_15_340 ();
 sg13g2_fill_2 FILLER_15_345 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_fill_2 FILLER_15_355 ();
 sg13g2_decap_4 FILLER_15_364 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_fill_2 FILLER_15_392 ();
 sg13g2_fill_2 FILLER_15_417 ();
 sg13g2_decap_4 FILLER_15_436 ();
 sg13g2_fill_1 FILLER_15_440 ();
 sg13g2_fill_2 FILLER_15_493 ();
 sg13g2_fill_1 FILLER_15_495 ();
 sg13g2_fill_1 FILLER_15_527 ();
 sg13g2_fill_1 FILLER_15_580 ();
 sg13g2_fill_1 FILLER_15_602 ();
 sg13g2_fill_1 FILLER_15_644 ();
 sg13g2_fill_2 FILLER_15_650 ();
 sg13g2_fill_2 FILLER_15_664 ();
 sg13g2_fill_1 FILLER_15_739 ();
 sg13g2_fill_2 FILLER_15_765 ();
 sg13g2_fill_1 FILLER_15_772 ();
 sg13g2_fill_1 FILLER_15_789 ();
 sg13g2_fill_2 FILLER_15_797 ();
 sg13g2_fill_1 FILLER_15_807 ();
 sg13g2_fill_2 FILLER_15_812 ();
 sg13g2_fill_2 FILLER_15_842 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_1 FILLER_16_15 ();
 sg13g2_fill_1 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_107 ();
 sg13g2_fill_2 FILLER_16_173 ();
 sg13g2_fill_2 FILLER_16_281 ();
 sg13g2_fill_1 FILLER_16_283 ();
 sg13g2_fill_2 FILLER_16_374 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_fill_2 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_441 ();
 sg13g2_fill_2 FILLER_16_447 ();
 sg13g2_decap_8 FILLER_16_460 ();
 sg13g2_fill_2 FILLER_16_467 ();
 sg13g2_fill_1 FILLER_16_469 ();
 sg13g2_fill_2 FILLER_16_474 ();
 sg13g2_fill_2 FILLER_16_480 ();
 sg13g2_fill_1 FILLER_16_482 ();
 sg13g2_decap_4 FILLER_16_509 ();
 sg13g2_fill_1 FILLER_16_513 ();
 sg13g2_fill_2 FILLER_16_522 ();
 sg13g2_fill_2 FILLER_16_554 ();
 sg13g2_fill_1 FILLER_16_556 ();
 sg13g2_fill_1 FILLER_16_573 ();
 sg13g2_fill_2 FILLER_16_605 ();
 sg13g2_fill_2 FILLER_16_620 ();
 sg13g2_fill_1 FILLER_16_622 ();
 sg13g2_fill_1 FILLER_16_665 ();
 sg13g2_fill_2 FILLER_16_683 ();
 sg13g2_fill_1 FILLER_16_693 ();
 sg13g2_fill_1 FILLER_16_715 ();
 sg13g2_fill_1 FILLER_16_746 ();
 sg13g2_fill_1 FILLER_16_755 ();
 sg13g2_fill_1 FILLER_16_775 ();
 sg13g2_fill_1 FILLER_16_785 ();
 sg13g2_fill_1 FILLER_16_839 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_346 ();
 sg13g2_fill_2 FILLER_17_376 ();
 sg13g2_fill_2 FILLER_17_405 ();
 sg13g2_fill_1 FILLER_17_412 ();
 sg13g2_fill_1 FILLER_17_449 ();
 sg13g2_fill_1 FILLER_17_455 ();
 sg13g2_fill_1 FILLER_17_604 ();
 sg13g2_fill_2 FILLER_17_615 ();
 sg13g2_fill_1 FILLER_17_622 ();
 sg13g2_fill_1 FILLER_17_628 ();
 sg13g2_fill_1 FILLER_17_640 ();
 sg13g2_fill_2 FILLER_17_649 ();
 sg13g2_fill_2 FILLER_17_675 ();
 sg13g2_fill_2 FILLER_17_720 ();
 sg13g2_fill_1 FILLER_17_825 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_fill_2 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_128 ();
 sg13g2_fill_1 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_139 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_fill_1 FILLER_18_259 ();
 sg13g2_fill_2 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_331 ();
 sg13g2_fill_1 FILLER_18_338 ();
 sg13g2_fill_1 FILLER_18_346 ();
 sg13g2_fill_1 FILLER_18_365 ();
 sg13g2_fill_1 FILLER_18_380 ();
 sg13g2_fill_1 FILLER_18_386 ();
 sg13g2_fill_1 FILLER_18_391 ();
 sg13g2_fill_2 FILLER_18_397 ();
 sg13g2_fill_1 FILLER_18_414 ();
 sg13g2_fill_1 FILLER_18_432 ();
 sg13g2_fill_1 FILLER_18_457 ();
 sg13g2_fill_2 FILLER_18_468 ();
 sg13g2_fill_2 FILLER_18_474 ();
 sg13g2_fill_1 FILLER_18_476 ();
 sg13g2_fill_2 FILLER_18_558 ();
 sg13g2_fill_1 FILLER_18_560 ();
 sg13g2_fill_2 FILLER_18_566 ();
 sg13g2_fill_1 FILLER_18_580 ();
 sg13g2_fill_1 FILLER_18_618 ();
 sg13g2_fill_2 FILLER_18_633 ();
 sg13g2_fill_1 FILLER_18_635 ();
 sg13g2_fill_1 FILLER_18_644 ();
 sg13g2_fill_1 FILLER_18_657 ();
 sg13g2_fill_1 FILLER_18_663 ();
 sg13g2_fill_2 FILLER_18_732 ();
 sg13g2_fill_2 FILLER_18_775 ();
 sg13g2_fill_1 FILLER_18_794 ();
 sg13g2_fill_1 FILLER_18_824 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_45 ();
 sg13g2_fill_2 FILLER_19_85 ();
 sg13g2_fill_1 FILLER_19_87 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_fill_1 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_190 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_fill_2 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_331 ();
 sg13g2_fill_1 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_348 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_414 ();
 sg13g2_decap_4 FILLER_19_466 ();
 sg13g2_fill_1 FILLER_19_470 ();
 sg13g2_decap_4 FILLER_19_479 ();
 sg13g2_fill_2 FILLER_19_483 ();
 sg13g2_fill_2 FILLER_19_519 ();
 sg13g2_decap_8 FILLER_19_526 ();
 sg13g2_fill_1 FILLER_19_533 ();
 sg13g2_fill_2 FILLER_19_551 ();
 sg13g2_fill_2 FILLER_19_562 ();
 sg13g2_fill_1 FILLER_19_564 ();
 sg13g2_fill_1 FILLER_19_598 ();
 sg13g2_fill_2 FILLER_19_626 ();
 sg13g2_fill_2 FILLER_19_647 ();
 sg13g2_fill_1 FILLER_19_682 ();
 sg13g2_fill_1 FILLER_19_726 ();
 sg13g2_fill_2 FILLER_19_736 ();
 sg13g2_fill_1 FILLER_19_748 ();
 sg13g2_fill_1 FILLER_19_769 ();
 sg13g2_fill_1 FILLER_19_783 ();
 sg13g2_fill_2 FILLER_19_804 ();
 sg13g2_fill_1 FILLER_19_813 ();
 sg13g2_fill_1 FILLER_19_877 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_9 ();
 sg13g2_fill_2 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_65 ();
 sg13g2_fill_1 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_fill_1 FILLER_20_298 ();
 sg13g2_fill_1 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_319 ();
 sg13g2_fill_1 FILLER_20_358 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_388 ();
 sg13g2_fill_1 FILLER_20_394 ();
 sg13g2_fill_2 FILLER_20_424 ();
 sg13g2_fill_2 FILLER_20_432 ();
 sg13g2_fill_1 FILLER_20_439 ();
 sg13g2_fill_1 FILLER_20_453 ();
 sg13g2_decap_4 FILLER_20_482 ();
 sg13g2_fill_1 FILLER_20_520 ();
 sg13g2_fill_1 FILLER_20_563 ();
 sg13g2_fill_2 FILLER_20_578 ();
 sg13g2_fill_2 FILLER_20_609 ();
 sg13g2_fill_1 FILLER_20_647 ();
 sg13g2_fill_1 FILLER_20_680 ();
 sg13g2_fill_1 FILLER_20_693 ();
 sg13g2_fill_1 FILLER_20_721 ();
 sg13g2_fill_1 FILLER_20_749 ();
 sg13g2_fill_2 FILLER_20_755 ();
 sg13g2_fill_2 FILLER_20_762 ();
 sg13g2_fill_1 FILLER_20_780 ();
 sg13g2_fill_2 FILLER_20_801 ();
 sg13g2_fill_2 FILLER_20_841 ();
 sg13g2_fill_2 FILLER_20_876 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_2 FILLER_21_190 ();
 sg13g2_fill_1 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_321 ();
 sg13g2_fill_1 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_360 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_397 ();
 sg13g2_fill_1 FILLER_21_403 ();
 sg13g2_fill_1 FILLER_21_409 ();
 sg13g2_fill_1 FILLER_21_414 ();
 sg13g2_fill_1 FILLER_21_425 ();
 sg13g2_fill_2 FILLER_21_433 ();
 sg13g2_fill_1 FILLER_21_435 ();
 sg13g2_fill_2 FILLER_21_451 ();
 sg13g2_fill_2 FILLER_21_468 ();
 sg13g2_fill_1 FILLER_21_474 ();
 sg13g2_fill_2 FILLER_21_526 ();
 sg13g2_fill_1 FILLER_21_528 ();
 sg13g2_fill_2 FILLER_21_559 ();
 sg13g2_fill_1 FILLER_21_565 ();
 sg13g2_fill_1 FILLER_21_571 ();
 sg13g2_fill_1 FILLER_21_582 ();
 sg13g2_fill_1 FILLER_21_593 ();
 sg13g2_fill_1 FILLER_21_606 ();
 sg13g2_fill_2 FILLER_21_619 ();
 sg13g2_fill_1 FILLER_21_621 ();
 sg13g2_fill_1 FILLER_21_633 ();
 sg13g2_fill_1 FILLER_21_639 ();
 sg13g2_fill_2 FILLER_21_680 ();
 sg13g2_fill_2 FILLER_21_714 ();
 sg13g2_fill_1 FILLER_21_736 ();
 sg13g2_fill_1 FILLER_21_784 ();
 sg13g2_fill_2 FILLER_21_790 ();
 sg13g2_fill_2 FILLER_21_809 ();
 sg13g2_fill_2 FILLER_21_847 ();
 sg13g2_fill_2 FILLER_21_870 ();
 sg13g2_fill_2 FILLER_21_876 ();
 sg13g2_fill_2 FILLER_22_77 ();
 sg13g2_fill_2 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_255 ();
 sg13g2_fill_1 FILLER_22_286 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_2 FILLER_22_358 ();
 sg13g2_fill_2 FILLER_22_365 ();
 sg13g2_decap_4 FILLER_22_372 ();
 sg13g2_fill_1 FILLER_22_376 ();
 sg13g2_fill_1 FILLER_22_415 ();
 sg13g2_decap_4 FILLER_22_436 ();
 sg13g2_fill_1 FILLER_22_440 ();
 sg13g2_fill_2 FILLER_22_564 ();
 sg13g2_fill_1 FILLER_22_566 ();
 sg13g2_fill_1 FILLER_22_578 ();
 sg13g2_fill_2 FILLER_22_625 ();
 sg13g2_fill_1 FILLER_22_627 ();
 sg13g2_fill_2 FILLER_22_641 ();
 sg13g2_fill_1 FILLER_22_658 ();
 sg13g2_fill_1 FILLER_22_683 ();
 sg13g2_fill_1 FILLER_22_689 ();
 sg13g2_fill_1 FILLER_22_695 ();
 sg13g2_fill_1 FILLER_22_707 ();
 sg13g2_fill_1 FILLER_22_725 ();
 sg13g2_fill_2 FILLER_22_755 ();
 sg13g2_fill_1 FILLER_22_769 ();
 sg13g2_fill_1 FILLER_22_799 ();
 sg13g2_fill_2 FILLER_22_852 ();
 sg13g2_fill_1 FILLER_22_859 ();
 sg13g2_fill_2 FILLER_22_876 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_36 ();
 sg13g2_fill_2 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_130 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_fill_2 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_229 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_2 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_fill_1 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_327 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_354 ();
 sg13g2_fill_1 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_389 ();
 sg13g2_fill_1 FILLER_23_394 ();
 sg13g2_fill_1 FILLER_23_418 ();
 sg13g2_fill_2 FILLER_23_424 ();
 sg13g2_fill_1 FILLER_23_426 ();
 sg13g2_fill_2 FILLER_23_458 ();
 sg13g2_decap_4 FILLER_23_470 ();
 sg13g2_decap_4 FILLER_23_511 ();
 sg13g2_fill_1 FILLER_23_515 ();
 sg13g2_fill_1 FILLER_23_520 ();
 sg13g2_fill_1 FILLER_23_532 ();
 sg13g2_fill_1 FILLER_23_538 ();
 sg13g2_fill_1 FILLER_23_642 ();
 sg13g2_fill_2 FILLER_23_688 ();
 sg13g2_fill_2 FILLER_23_745 ();
 sg13g2_fill_1 FILLER_23_800 ();
 sg13g2_fill_1 FILLER_23_815 ();
 sg13g2_fill_1 FILLER_23_835 ();
 sg13g2_fill_2 FILLER_23_856 ();
 sg13g2_fill_2 FILLER_23_875 ();
 sg13g2_fill_1 FILLER_23_877 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_fill_1 FILLER_24_20 ();
 sg13g2_fill_2 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_fill_2 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_254 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_350 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_decap_4 FILLER_24_395 ();
 sg13g2_fill_1 FILLER_24_404 ();
 sg13g2_fill_2 FILLER_24_421 ();
 sg13g2_fill_1 FILLER_24_423 ();
 sg13g2_fill_2 FILLER_24_429 ();
 sg13g2_fill_1 FILLER_24_431 ();
 sg13g2_fill_2 FILLER_24_446 ();
 sg13g2_fill_1 FILLER_24_448 ();
 sg13g2_fill_1 FILLER_24_454 ();
 sg13g2_fill_1 FILLER_24_459 ();
 sg13g2_fill_1 FILLER_24_465 ();
 sg13g2_decap_4 FILLER_24_494 ();
 sg13g2_fill_2 FILLER_24_498 ();
 sg13g2_fill_1 FILLER_24_517 ();
 sg13g2_fill_1 FILLER_24_526 ();
 sg13g2_decap_4 FILLER_24_549 ();
 sg13g2_decap_4 FILLER_24_557 ();
 sg13g2_decap_4 FILLER_24_565 ();
 sg13g2_fill_2 FILLER_24_595 ();
 sg13g2_fill_1 FILLER_24_597 ();
 sg13g2_decap_4 FILLER_24_628 ();
 sg13g2_fill_1 FILLER_24_632 ();
 sg13g2_fill_2 FILLER_24_646 ();
 sg13g2_fill_1 FILLER_24_670 ();
 sg13g2_fill_1 FILLER_24_758 ();
 sg13g2_fill_2 FILLER_24_793 ();
 sg13g2_fill_1 FILLER_24_817 ();
 sg13g2_fill_2 FILLER_24_826 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_6 ();
 sg13g2_fill_2 FILLER_25_16 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_157 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_fill_2 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_287 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_475 ();
 sg13g2_fill_2 FILLER_25_486 ();
 sg13g2_fill_1 FILLER_25_493 ();
 sg13g2_fill_2 FILLER_25_499 ();
 sg13g2_fill_1 FILLER_25_506 ();
 sg13g2_fill_2 FILLER_25_532 ();
 sg13g2_fill_1 FILLER_25_544 ();
 sg13g2_fill_1 FILLER_25_555 ();
 sg13g2_fill_2 FILLER_25_566 ();
 sg13g2_decap_8 FILLER_25_624 ();
 sg13g2_decap_4 FILLER_25_631 ();
 sg13g2_fill_1 FILLER_25_635 ();
 sg13g2_fill_1 FILLER_25_644 ();
 sg13g2_fill_1 FILLER_25_653 ();
 sg13g2_fill_1 FILLER_25_715 ();
 sg13g2_fill_2 FILLER_25_743 ();
 sg13g2_fill_1 FILLER_25_800 ();
 sg13g2_fill_2 FILLER_25_836 ();
 sg13g2_fill_2 FILLER_25_859 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_376 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_fill_1 FILLER_26_400 ();
 sg13g2_fill_1 FILLER_26_427 ();
 sg13g2_fill_2 FILLER_26_432 ();
 sg13g2_fill_1 FILLER_26_434 ();
 sg13g2_fill_2 FILLER_26_439 ();
 sg13g2_decap_4 FILLER_26_449 ();
 sg13g2_fill_1 FILLER_26_453 ();
 sg13g2_fill_1 FILLER_26_459 ();
 sg13g2_fill_1 FILLER_26_465 ();
 sg13g2_fill_1 FILLER_26_470 ();
 sg13g2_fill_2 FILLER_26_498 ();
 sg13g2_fill_1 FILLER_26_505 ();
 sg13g2_fill_2 FILLER_26_542 ();
 sg13g2_fill_2 FILLER_26_580 ();
 sg13g2_fill_1 FILLER_26_582 ();
 sg13g2_decap_8 FILLER_26_587 ();
 sg13g2_decap_4 FILLER_26_594 ();
 sg13g2_fill_1 FILLER_26_602 ();
 sg13g2_fill_2 FILLER_26_607 ();
 sg13g2_fill_1 FILLER_26_609 ();
 sg13g2_fill_1 FILLER_26_636 ();
 sg13g2_fill_2 FILLER_26_645 ();
 sg13g2_fill_2 FILLER_26_743 ();
 sg13g2_fill_2 FILLER_26_781 ();
 sg13g2_fill_1 FILLER_26_787 ();
 sg13g2_fill_2 FILLER_26_820 ();
 sg13g2_fill_1 FILLER_26_863 ();
 sg13g2_fill_2 FILLER_26_876 ();
 sg13g2_fill_1 FILLER_27_26 ();
 sg13g2_fill_2 FILLER_27_61 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_220 ();
 sg13g2_fill_2 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_276 ();
 sg13g2_fill_2 FILLER_27_290 ();
 sg13g2_decap_4 FILLER_27_346 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_decap_4 FILLER_27_361 ();
 sg13g2_fill_2 FILLER_27_383 ();
 sg13g2_fill_1 FILLER_27_385 ();
 sg13g2_fill_2 FILLER_27_447 ();
 sg13g2_fill_1 FILLER_27_449 ();
 sg13g2_decap_4 FILLER_27_496 ();
 sg13g2_fill_2 FILLER_27_500 ();
 sg13g2_decap_4 FILLER_27_511 ();
 sg13g2_fill_2 FILLER_27_528 ();
 sg13g2_fill_1 FILLER_27_546 ();
 sg13g2_fill_1 FILLER_27_551 ();
 sg13g2_fill_1 FILLER_27_616 ();
 sg13g2_fill_1 FILLER_27_625 ();
 sg13g2_fill_2 FILLER_27_645 ();
 sg13g2_fill_2 FILLER_27_671 ();
 sg13g2_fill_2 FILLER_27_700 ();
 sg13g2_fill_1 FILLER_27_742 ();
 sg13g2_fill_1 FILLER_27_769 ();
 sg13g2_fill_1 FILLER_27_814 ();
 sg13g2_fill_2 FILLER_27_871 ();
 sg13g2_fill_1 FILLER_27_873 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_17 ();
 sg13g2_fill_1 FILLER_28_19 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_fill_1 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_284 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_331 ();
 sg13g2_fill_1 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_402 ();
 sg13g2_fill_1 FILLER_28_404 ();
 sg13g2_decap_4 FILLER_28_417 ();
 sg13g2_fill_2 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_decap_8 FILLER_28_438 ();
 sg13g2_decap_8 FILLER_28_445 ();
 sg13g2_fill_2 FILLER_28_452 ();
 sg13g2_fill_1 FILLER_28_454 ();
 sg13g2_fill_2 FILLER_28_470 ();
 sg13g2_fill_1 FILLER_28_501 ();
 sg13g2_fill_1 FILLER_28_507 ();
 sg13g2_fill_1 FILLER_28_513 ();
 sg13g2_fill_2 FILLER_28_519 ();
 sg13g2_fill_2 FILLER_28_526 ();
 sg13g2_fill_1 FILLER_28_537 ();
 sg13g2_fill_1 FILLER_28_561 ();
 sg13g2_fill_1 FILLER_28_567 ();
 sg13g2_fill_2 FILLER_28_575 ();
 sg13g2_fill_2 FILLER_28_622 ();
 sg13g2_fill_1 FILLER_28_708 ();
 sg13g2_fill_1 FILLER_28_723 ();
 sg13g2_fill_1 FILLER_28_728 ();
 sg13g2_fill_1 FILLER_28_733 ();
 sg13g2_fill_2 FILLER_28_828 ();
 sg13g2_fill_2 FILLER_28_834 ();
 sg13g2_fill_1 FILLER_28_836 ();
 sg13g2_fill_2 FILLER_28_841 ();
 sg13g2_fill_2 FILLER_28_847 ();
 sg13g2_fill_2 FILLER_28_859 ();
 sg13g2_decap_8 FILLER_28_871 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_15 ();
 sg13g2_fill_1 FILLER_29_43 ();
 sg13g2_fill_2 FILLER_29_156 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_fill_1 FILLER_29_304 ();
 sg13g2_fill_2 FILLER_29_385 ();
 sg13g2_fill_1 FILLER_29_418 ();
 sg13g2_decap_8 FILLER_29_423 ();
 sg13g2_decap_4 FILLER_29_430 ();
 sg13g2_fill_1 FILLER_29_446 ();
 sg13g2_fill_2 FILLER_29_481 ();
 sg13g2_fill_1 FILLER_29_491 ();
 sg13g2_fill_2 FILLER_29_526 ();
 sg13g2_fill_1 FILLER_29_564 ();
 sg13g2_fill_1 FILLER_29_570 ();
 sg13g2_fill_1 FILLER_29_599 ();
 sg13g2_fill_2 FILLER_29_604 ();
 sg13g2_fill_2 FILLER_29_610 ();
 sg13g2_fill_1 FILLER_29_612 ();
 sg13g2_fill_1 FILLER_29_617 ();
 sg13g2_fill_2 FILLER_29_641 ();
 sg13g2_fill_2 FILLER_29_701 ();
 sg13g2_fill_1 FILLER_29_840 ();
 sg13g2_decap_4 FILLER_29_872 ();
 sg13g2_fill_2 FILLER_29_876 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_27 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_89 ();
 sg13g2_fill_1 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_130 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_fill_2 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_211 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_fill_2 FILLER_30_247 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_336 ();
 sg13g2_fill_1 FILLER_30_342 ();
 sg13g2_fill_1 FILLER_30_347 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_fill_2 FILLER_30_383 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_425 ();
 sg13g2_fill_2 FILLER_30_429 ();
 sg13g2_fill_2 FILLER_30_451 ();
 sg13g2_fill_1 FILLER_30_492 ();
 sg13g2_fill_2 FILLER_30_538 ();
 sg13g2_fill_2 FILLER_30_590 ();
 sg13g2_fill_1 FILLER_30_610 ();
 sg13g2_fill_2 FILLER_30_635 ();
 sg13g2_fill_2 FILLER_30_667 ();
 sg13g2_fill_1 FILLER_30_844 ();
 sg13g2_fill_2 FILLER_30_855 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_117 ();
 sg13g2_fill_2 FILLER_31_149 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_303 ();
 sg13g2_decap_4 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_390 ();
 sg13g2_fill_1 FILLER_31_425 ();
 sg13g2_fill_1 FILLER_31_436 ();
 sg13g2_fill_1 FILLER_31_441 ();
 sg13g2_fill_1 FILLER_31_524 ();
 sg13g2_fill_1 FILLER_31_530 ();
 sg13g2_fill_1 FILLER_31_537 ();
 sg13g2_fill_2 FILLER_31_560 ();
 sg13g2_fill_1 FILLER_31_566 ();
 sg13g2_fill_2 FILLER_31_585 ();
 sg13g2_fill_1 FILLER_31_592 ();
 sg13g2_fill_1 FILLER_31_597 ();
 sg13g2_fill_1 FILLER_31_603 ();
 sg13g2_fill_1 FILLER_31_609 ();
 sg13g2_fill_1 FILLER_31_638 ();
 sg13g2_fill_2 FILLER_31_685 ();
 sg13g2_fill_2 FILLER_31_742 ();
 sg13g2_fill_1 FILLER_31_765 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_fill_1 FILLER_31_833 ();
 sg13g2_decap_4 FILLER_31_872 ();
 sg13g2_fill_2 FILLER_31_876 ();
 sg13g2_fill_1 FILLER_32_26 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_fill_1 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_255 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_1 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_284 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_fill_2 FILLER_32_296 ();
 sg13g2_fill_1 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_371 ();
 sg13g2_fill_1 FILLER_32_376 ();
 sg13g2_fill_2 FILLER_32_401 ();
 sg13g2_fill_2 FILLER_32_452 ();
 sg13g2_fill_2 FILLER_32_512 ();
 sg13g2_fill_2 FILLER_32_606 ();
 sg13g2_fill_1 FILLER_32_630 ();
 sg13g2_fill_2 FILLER_32_635 ();
 sg13g2_fill_1 FILLER_32_642 ();
 sg13g2_fill_1 FILLER_32_667 ();
 sg13g2_fill_1 FILLER_32_672 ();
 sg13g2_fill_1 FILLER_32_717 ();
 sg13g2_fill_1 FILLER_32_747 ();
 sg13g2_fill_1 FILLER_32_779 ();
 sg13g2_fill_2 FILLER_32_801 ();
 sg13g2_fill_1 FILLER_32_803 ();
 sg13g2_decap_4 FILLER_32_845 ();
 sg13g2_decap_8 FILLER_32_870 ();
 sg13g2_fill_1 FILLER_32_877 ();
 sg13g2_fill_2 FILLER_33_29 ();
 sg13g2_fill_1 FILLER_33_124 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_fill_2 FILLER_33_228 ();
 sg13g2_fill_1 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_281 ();
 sg13g2_fill_1 FILLER_33_288 ();
 sg13g2_fill_2 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_2 FILLER_33_409 ();
 sg13g2_fill_2 FILLER_33_451 ();
 sg13g2_fill_1 FILLER_33_458 ();
 sg13g2_fill_1 FILLER_33_463 ();
 sg13g2_fill_1 FILLER_33_473 ();
 sg13g2_fill_1 FILLER_33_494 ();
 sg13g2_fill_2 FILLER_33_563 ();
 sg13g2_fill_1 FILLER_33_565 ();
 sg13g2_fill_2 FILLER_33_592 ();
 sg13g2_fill_2 FILLER_33_599 ();
 sg13g2_fill_2 FILLER_33_606 ();
 sg13g2_fill_2 FILLER_33_613 ();
 sg13g2_fill_2 FILLER_33_654 ();
 sg13g2_fill_2 FILLER_33_670 ();
 sg13g2_fill_2 FILLER_33_744 ();
 sg13g2_fill_1 FILLER_33_801 ();
 sg13g2_fill_1 FILLER_33_823 ();
 sg13g2_fill_2 FILLER_33_834 ();
 sg13g2_decap_4 FILLER_33_856 ();
 sg13g2_fill_1 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_33_871 ();
 sg13g2_fill_2 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_fill_1 FILLER_34_340 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_1 FILLER_34_352 ();
 sg13g2_fill_2 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_fill_2 FILLER_34_393 ();
 sg13g2_fill_1 FILLER_34_395 ();
 sg13g2_fill_1 FILLER_34_427 ();
 sg13g2_fill_2 FILLER_34_446 ();
 sg13g2_fill_1 FILLER_34_484 ();
 sg13g2_fill_2 FILLER_34_490 ();
 sg13g2_fill_1 FILLER_34_501 ();
 sg13g2_fill_2 FILLER_34_590 ();
 sg13g2_fill_1 FILLER_34_602 ();
 sg13g2_fill_1 FILLER_34_629 ();
 sg13g2_fill_2 FILLER_34_643 ();
 sg13g2_fill_1 FILLER_34_645 ();
 sg13g2_fill_2 FILLER_34_656 ();
 sg13g2_fill_2 FILLER_34_698 ();
 sg13g2_fill_2 FILLER_34_704 ();
 sg13g2_fill_1 FILLER_34_706 ();
 sg13g2_fill_2 FILLER_34_730 ();
 sg13g2_fill_1 FILLER_34_732 ();
 sg13g2_fill_1 FILLER_34_745 ();
 sg13g2_fill_1 FILLER_34_751 ();
 sg13g2_fill_1 FILLER_34_794 ();
 sg13g2_fill_1 FILLER_34_799 ();
 sg13g2_decap_8 FILLER_34_842 ();
 sg13g2_fill_1 FILLER_34_849 ();
 sg13g2_decap_8 FILLER_34_871 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_34 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_decap_4 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_320 ();
 sg13g2_fill_2 FILLER_35_331 ();
 sg13g2_fill_2 FILLER_35_367 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_fill_2 FILLER_35_384 ();
 sg13g2_fill_1 FILLER_35_386 ();
 sg13g2_fill_2 FILLER_35_464 ();
 sg13g2_fill_1 FILLER_35_470 ();
 sg13g2_fill_2 FILLER_35_476 ();
 sg13g2_fill_1 FILLER_35_488 ();
 sg13g2_fill_1 FILLER_35_494 ();
 sg13g2_fill_2 FILLER_35_572 ();
 sg13g2_fill_1 FILLER_35_574 ();
 sg13g2_decap_4 FILLER_35_588 ();
 sg13g2_fill_1 FILLER_35_592 ();
 sg13g2_fill_2 FILLER_35_597 ();
 sg13g2_decap_8 FILLER_35_603 ();
 sg13g2_decap_4 FILLER_35_618 ();
 sg13g2_fill_1 FILLER_35_622 ();
 sg13g2_fill_1 FILLER_35_670 ();
 sg13g2_fill_2 FILLER_35_681 ();
 sg13g2_fill_2 FILLER_35_717 ();
 sg13g2_fill_1 FILLER_35_719 ();
 sg13g2_fill_2 FILLER_35_746 ();
 sg13g2_fill_2 FILLER_35_769 ();
 sg13g2_fill_1 FILLER_35_771 ();
 sg13g2_decap_4 FILLER_35_814 ();
 sg13g2_decap_8 FILLER_35_870 ();
 sg13g2_fill_1 FILLER_35_877 ();
 sg13g2_fill_2 FILLER_36_82 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_191 ();
 sg13g2_fill_2 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_341 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_decap_4 FILLER_36_407 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_2 FILLER_36_439 ();
 sg13g2_fill_1 FILLER_36_451 ();
 sg13g2_fill_1 FILLER_36_513 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_fill_1 FILLER_36_554 ();
 sg13g2_fill_2 FILLER_36_601 ();
 sg13g2_fill_1 FILLER_36_641 ();
 sg13g2_fill_2 FILLER_36_673 ();
 sg13g2_fill_1 FILLER_36_675 ();
 sg13g2_fill_1 FILLER_36_684 ();
 sg13g2_fill_1 FILLER_36_702 ();
 sg13g2_fill_2 FILLER_36_744 ();
 sg13g2_fill_2 FILLER_36_754 ();
 sg13g2_decap_8 FILLER_36_760 ();
 sg13g2_decap_4 FILLER_36_767 ();
 sg13g2_fill_2 FILLER_36_783 ();
 sg13g2_fill_2 FILLER_36_798 ();
 sg13g2_fill_1 FILLER_36_810 ();
 sg13g2_fill_1 FILLER_36_821 ();
 sg13g2_fill_1 FILLER_36_843 ();
 sg13g2_fill_2 FILLER_36_865 ();
 sg13g2_fill_1 FILLER_36_877 ();
 sg13g2_fill_2 FILLER_37_108 ();
 sg13g2_fill_1 FILLER_37_110 ();
 sg13g2_fill_1 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_157 ();
 sg13g2_fill_1 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_fill_2 FILLER_37_177 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_189 ();
 sg13g2_fill_2 FILLER_37_219 ();
 sg13g2_fill_1 FILLER_37_229 ();
 sg13g2_fill_1 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_253 ();
 sg13g2_fill_2 FILLER_37_265 ();
 sg13g2_fill_2 FILLER_37_280 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_298 ();
 sg13g2_fill_2 FILLER_37_339 ();
 sg13g2_fill_2 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_414 ();
 sg13g2_fill_1 FILLER_37_421 ();
 sg13g2_fill_1 FILLER_37_432 ();
 sg13g2_fill_1 FILLER_37_452 ();
 sg13g2_fill_2 FILLER_37_462 ();
 sg13g2_fill_1 FILLER_37_474 ();
 sg13g2_fill_1 FILLER_37_479 ();
 sg13g2_fill_1 FILLER_37_484 ();
 sg13g2_fill_1 FILLER_37_489 ();
 sg13g2_fill_1 FILLER_37_494 ();
 sg13g2_fill_1 FILLER_37_501 ();
 sg13g2_fill_2 FILLER_37_506 ();
 sg13g2_fill_1 FILLER_37_517 ();
 sg13g2_fill_2 FILLER_37_524 ();
 sg13g2_fill_1 FILLER_37_547 ();
 sg13g2_fill_2 FILLER_37_557 ();
 sg13g2_fill_2 FILLER_37_586 ();
 sg13g2_fill_2 FILLER_37_644 ();
 sg13g2_fill_2 FILLER_37_676 ();
 sg13g2_fill_2 FILLER_37_721 ();
 sg13g2_fill_1 FILLER_37_723 ();
 sg13g2_fill_2 FILLER_37_846 ();
 sg13g2_fill_1 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_138 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_fill_1 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_245 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_1 FILLER_38_296 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_2 FILLER_38_336 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_384 ();
 sg13g2_fill_2 FILLER_38_421 ();
 sg13g2_fill_1 FILLER_38_440 ();
 sg13g2_fill_1 FILLER_38_456 ();
 sg13g2_fill_2 FILLER_38_462 ();
 sg13g2_fill_2 FILLER_38_471 ();
 sg13g2_fill_1 FILLER_38_473 ();
 sg13g2_decap_4 FILLER_38_478 ();
 sg13g2_fill_2 FILLER_38_482 ();
 sg13g2_fill_2 FILLER_38_506 ();
 sg13g2_fill_1 FILLER_38_569 ();
 sg13g2_fill_1 FILLER_38_587 ();
 sg13g2_decap_4 FILLER_38_603 ();
 sg13g2_fill_1 FILLER_38_646 ();
 sg13g2_fill_1 FILLER_38_652 ();
 sg13g2_fill_2 FILLER_38_693 ();
 sg13g2_fill_2 FILLER_38_715 ();
 sg13g2_fill_2 FILLER_38_763 ();
 sg13g2_fill_1 FILLER_38_801 ();
 sg13g2_fill_2 FILLER_38_834 ();
 sg13g2_fill_2 FILLER_38_876 ();
 sg13g2_fill_2 FILLER_39_65 ();
 sg13g2_fill_2 FILLER_39_71 ();
 sg13g2_fill_1 FILLER_39_129 ();
 sg13g2_fill_1 FILLER_39_165 ();
 sg13g2_fill_2 FILLER_39_178 ();
 sg13g2_fill_1 FILLER_39_184 ();
 sg13g2_fill_2 FILLER_39_193 ();
 sg13g2_fill_1 FILLER_39_199 ();
 sg13g2_fill_2 FILLER_39_220 ();
 sg13g2_fill_1 FILLER_39_263 ();
 sg13g2_fill_1 FILLER_39_277 ();
 sg13g2_fill_1 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_365 ();
 sg13g2_fill_2 FILLER_39_389 ();
 sg13g2_fill_2 FILLER_39_396 ();
 sg13g2_fill_2 FILLER_39_402 ();
 sg13g2_fill_1 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_410 ();
 sg13g2_fill_1 FILLER_39_461 ();
 sg13g2_fill_1 FILLER_39_470 ();
 sg13g2_fill_1 FILLER_39_492 ();
 sg13g2_fill_2 FILLER_39_561 ();
 sg13g2_fill_2 FILLER_39_567 ();
 sg13g2_decap_4 FILLER_39_583 ();
 sg13g2_fill_1 FILLER_39_587 ();
 sg13g2_fill_2 FILLER_39_603 ();
 sg13g2_fill_1 FILLER_39_649 ();
 sg13g2_fill_2 FILLER_39_659 ();
 sg13g2_fill_2 FILLER_39_704 ();
 sg13g2_fill_1 FILLER_39_754 ();
 sg13g2_fill_2 FILLER_39_809 ();
 sg13g2_fill_1 FILLER_39_837 ();
 sg13g2_fill_1 FILLER_39_865 ();
 sg13g2_fill_2 FILLER_39_875 ();
 sg13g2_fill_1 FILLER_39_877 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_13 ();
 sg13g2_fill_1 FILLER_40_24 ();
 sg13g2_fill_1 FILLER_40_29 ();
 sg13g2_fill_1 FILLER_40_44 ();
 sg13g2_fill_1 FILLER_40_53 ();
 sg13g2_fill_2 FILLER_40_86 ();
 sg13g2_fill_2 FILLER_40_99 ();
 sg13g2_fill_1 FILLER_40_153 ();
 sg13g2_fill_1 FILLER_40_159 ();
 sg13g2_fill_1 FILLER_40_169 ();
 sg13g2_fill_1 FILLER_40_175 ();
 sg13g2_fill_2 FILLER_40_207 ();
 sg13g2_fill_1 FILLER_40_213 ();
 sg13g2_fill_1 FILLER_40_273 ();
 sg13g2_fill_1 FILLER_40_278 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_4 FILLER_40_294 ();
 sg13g2_decap_4 FILLER_40_302 ();
 sg13g2_decap_4 FILLER_40_311 ();
 sg13g2_fill_2 FILLER_40_335 ();
 sg13g2_fill_2 FILLER_40_356 ();
 sg13g2_fill_2 FILLER_40_384 ();
 sg13g2_fill_2 FILLER_40_424 ();
 sg13g2_fill_2 FILLER_40_441 ();
 sg13g2_fill_2 FILLER_40_480 ();
 sg13g2_fill_2 FILLER_40_494 ();
 sg13g2_fill_1 FILLER_40_526 ();
 sg13g2_fill_1 FILLER_40_532 ();
 sg13g2_fill_1 FILLER_40_546 ();
 sg13g2_fill_1 FILLER_40_556 ();
 sg13g2_fill_1 FILLER_40_569 ();
 sg13g2_decap_4 FILLER_40_604 ();
 sg13g2_fill_2 FILLER_40_608 ();
 sg13g2_fill_2 FILLER_40_632 ();
 sg13g2_decap_4 FILLER_40_658 ();
 sg13g2_fill_1 FILLER_40_676 ();
 sg13g2_fill_1 FILLER_40_713 ();
 sg13g2_fill_1 FILLER_40_728 ();
 sg13g2_fill_2 FILLER_40_755 ();
 sg13g2_fill_1 FILLER_40_757 ();
 sg13g2_fill_2 FILLER_40_766 ();
 sg13g2_fill_2 FILLER_40_850 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_162 ();
 sg13g2_fill_2 FILLER_41_210 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_fill_1 FILLER_41_273 ();
 sg13g2_fill_2 FILLER_41_278 ();
 sg13g2_fill_1 FILLER_41_280 ();
 sg13g2_fill_2 FILLER_41_317 ();
 sg13g2_fill_2 FILLER_41_364 ();
 sg13g2_fill_1 FILLER_41_401 ();
 sg13g2_fill_1 FILLER_41_454 ();
 sg13g2_fill_2 FILLER_41_475 ();
 sg13g2_fill_1 FILLER_41_477 ();
 sg13g2_fill_1 FILLER_41_498 ();
 sg13g2_fill_2 FILLER_41_507 ();
 sg13g2_decap_8 FILLER_41_516 ();
 sg13g2_fill_1 FILLER_41_557 ();
 sg13g2_fill_1 FILLER_41_563 ();
 sg13g2_fill_1 FILLER_41_578 ();
 sg13g2_fill_1 FILLER_41_583 ();
 sg13g2_fill_2 FILLER_41_610 ();
 sg13g2_fill_1 FILLER_41_697 ();
 sg13g2_fill_1 FILLER_41_712 ();
 sg13g2_fill_2 FILLER_41_732 ();
 sg13g2_fill_1 FILLER_41_734 ();
 sg13g2_fill_1 FILLER_41_745 ();
 sg13g2_fill_1 FILLER_41_802 ();
 sg13g2_fill_1 FILLER_41_863 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_fill_2 FILLER_41_875 ();
 sg13g2_fill_1 FILLER_41_877 ();
 sg13g2_fill_1 FILLER_42_26 ();
 sg13g2_fill_1 FILLER_42_74 ();
 sg13g2_fill_1 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_121 ();
 sg13g2_fill_1 FILLER_42_131 ();
 sg13g2_fill_1 FILLER_42_136 ();
 sg13g2_fill_1 FILLER_42_148 ();
 sg13g2_fill_1 FILLER_42_154 ();
 sg13g2_fill_2 FILLER_42_232 ();
 sg13g2_fill_1 FILLER_42_247 ();
 sg13g2_fill_2 FILLER_42_264 ();
 sg13g2_fill_2 FILLER_42_271 ();
 sg13g2_fill_1 FILLER_42_273 ();
 sg13g2_fill_2 FILLER_42_280 ();
 sg13g2_fill_1 FILLER_42_282 ();
 sg13g2_fill_1 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_326 ();
 sg13g2_fill_1 FILLER_42_336 ();
 sg13g2_fill_2 FILLER_42_342 ();
 sg13g2_fill_1 FILLER_42_344 ();
 sg13g2_fill_2 FILLER_42_349 ();
 sg13g2_fill_1 FILLER_42_351 ();
 sg13g2_fill_2 FILLER_42_429 ();
 sg13g2_fill_2 FILLER_42_436 ();
 sg13g2_fill_1 FILLER_42_451 ();
 sg13g2_fill_1 FILLER_42_456 ();
 sg13g2_decap_4 FILLER_42_476 ();
 sg13g2_fill_1 FILLER_42_480 ();
 sg13g2_fill_1 FILLER_42_511 ();
 sg13g2_fill_2 FILLER_42_517 ();
 sg13g2_decap_4 FILLER_42_523 ();
 sg13g2_fill_1 FILLER_42_532 ();
 sg13g2_fill_2 FILLER_42_564 ();
 sg13g2_fill_2 FILLER_42_592 ();
 sg13g2_decap_4 FILLER_42_598 ();
 sg13g2_fill_2 FILLER_42_606 ();
 sg13g2_decap_4 FILLER_42_643 ();
 sg13g2_decap_8 FILLER_42_655 ();
 sg13g2_fill_2 FILLER_42_662 ();
 sg13g2_fill_1 FILLER_42_664 ();
 sg13g2_fill_2 FILLER_42_678 ();
 sg13g2_fill_1 FILLER_42_680 ();
 sg13g2_fill_2 FILLER_42_717 ();
 sg13g2_fill_2 FILLER_42_759 ();
 sg13g2_fill_1 FILLER_42_761 ();
 sg13g2_fill_2 FILLER_42_772 ();
 sg13g2_fill_2 FILLER_42_814 ();
 sg13g2_fill_1 FILLER_42_816 ();
 sg13g2_fill_2 FILLER_42_875 ();
 sg13g2_fill_1 FILLER_42_877 ();
 sg13g2_fill_1 FILLER_43_4 ();
 sg13g2_fill_1 FILLER_43_13 ();
 sg13g2_fill_2 FILLER_43_24 ();
 sg13g2_fill_1 FILLER_43_36 ();
 sg13g2_fill_1 FILLER_43_41 ();
 sg13g2_fill_1 FILLER_43_85 ();
 sg13g2_fill_1 FILLER_43_96 ();
 sg13g2_fill_1 FILLER_43_122 ();
 sg13g2_fill_1 FILLER_43_155 ();
 sg13g2_fill_1 FILLER_43_161 ();
 sg13g2_fill_2 FILLER_43_196 ();
 sg13g2_fill_2 FILLER_43_203 ();
 sg13g2_fill_1 FILLER_43_215 ();
 sg13g2_fill_2 FILLER_43_252 ();
 sg13g2_fill_1 FILLER_43_254 ();
 sg13g2_fill_1 FILLER_43_297 ();
 sg13g2_fill_2 FILLER_43_306 ();
 sg13g2_fill_1 FILLER_43_308 ();
 sg13g2_fill_1 FILLER_43_314 ();
 sg13g2_fill_1 FILLER_43_319 ();
 sg13g2_fill_1 FILLER_43_324 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_fill_2 FILLER_43_334 ();
 sg13g2_fill_2 FILLER_43_385 ();
 sg13g2_fill_2 FILLER_43_391 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_decap_4 FILLER_43_413 ();
 sg13g2_fill_2 FILLER_43_456 ();
 sg13g2_fill_1 FILLER_43_462 ();
 sg13g2_decap_4 FILLER_43_467 ();
 sg13g2_fill_2 FILLER_43_475 ();
 sg13g2_fill_1 FILLER_43_477 ();
 sg13g2_fill_1 FILLER_43_500 ();
 sg13g2_decap_4 FILLER_43_506 ();
 sg13g2_fill_2 FILLER_43_510 ();
 sg13g2_fill_2 FILLER_43_535 ();
 sg13g2_fill_1 FILLER_43_544 ();
 sg13g2_fill_1 FILLER_43_549 ();
 sg13g2_fill_1 FILLER_43_554 ();
 sg13g2_fill_1 FILLER_43_563 ();
 sg13g2_fill_1 FILLER_43_568 ();
 sg13g2_fill_1 FILLER_43_595 ();
 sg13g2_fill_1 FILLER_43_664 ();
 sg13g2_fill_1 FILLER_43_695 ();
 sg13g2_decap_4 FILLER_43_802 ();
 sg13g2_fill_1 FILLER_44_61 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_fill_2 FILLER_44_132 ();
 sg13g2_fill_1 FILLER_44_176 ();
 sg13g2_fill_1 FILLER_44_260 ();
 sg13g2_fill_1 FILLER_44_316 ();
 sg13g2_fill_2 FILLER_44_418 ();
 sg13g2_fill_2 FILLER_44_428 ();
 sg13g2_fill_2 FILLER_44_453 ();
 sg13g2_fill_1 FILLER_44_493 ();
 sg13g2_decap_4 FILLER_44_511 ();
 sg13g2_fill_2 FILLER_44_515 ();
 sg13g2_fill_2 FILLER_44_529 ();
 sg13g2_fill_1 FILLER_44_531 ();
 sg13g2_fill_1 FILLER_44_547 ();
 sg13g2_fill_2 FILLER_44_589 ();
 sg13g2_fill_1 FILLER_44_591 ();
 sg13g2_fill_1 FILLER_44_600 ();
 sg13g2_fill_2 FILLER_44_639 ();
 sg13g2_fill_1 FILLER_44_641 ();
 sg13g2_fill_2 FILLER_44_653 ();
 sg13g2_fill_2 FILLER_44_687 ();
 sg13g2_fill_2 FILLER_44_745 ();
 sg13g2_fill_1 FILLER_44_747 ();
 sg13g2_fill_1 FILLER_44_836 ();
 sg13g2_fill_1 FILLER_44_851 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_174 ();
 sg13g2_fill_1 FILLER_45_185 ();
 sg13g2_fill_2 FILLER_45_190 ();
 sg13g2_fill_1 FILLER_45_229 ();
 sg13g2_fill_2 FILLER_45_280 ();
 sg13g2_fill_1 FILLER_45_287 ();
 sg13g2_fill_2 FILLER_45_297 ();
 sg13g2_fill_2 FILLER_45_308 ();
 sg13g2_fill_1 FILLER_45_310 ();
 sg13g2_fill_1 FILLER_45_329 ();
 sg13g2_fill_1 FILLER_45_344 ();
 sg13g2_fill_1 FILLER_45_355 ();
 sg13g2_fill_1 FILLER_45_366 ();
 sg13g2_fill_2 FILLER_45_397 ();
 sg13g2_fill_1 FILLER_45_420 ();
 sg13g2_fill_1 FILLER_45_426 ();
 sg13g2_fill_1 FILLER_45_434 ();
 sg13g2_fill_1 FILLER_45_481 ();
 sg13g2_fill_1 FILLER_45_499 ();
 sg13g2_fill_1 FILLER_45_515 ();
 sg13g2_fill_2 FILLER_45_532 ();
 sg13g2_fill_1 FILLER_45_539 ();
 sg13g2_fill_1 FILLER_45_543 ();
 sg13g2_fill_1 FILLER_45_557 ();
 sg13g2_fill_1 FILLER_45_566 ();
 sg13g2_fill_1 FILLER_45_580 ();
 sg13g2_fill_2 FILLER_45_585 ();
 sg13g2_fill_1 FILLER_45_587 ();
 sg13g2_fill_2 FILLER_45_625 ();
 sg13g2_fill_1 FILLER_45_627 ();
 sg13g2_fill_1 FILLER_45_633 ();
 sg13g2_fill_1 FILLER_45_639 ();
 sg13g2_fill_1 FILLER_45_652 ();
 sg13g2_fill_2 FILLER_45_669 ();
 sg13g2_fill_1 FILLER_45_671 ();
 sg13g2_fill_2 FILLER_45_688 ();
 sg13g2_fill_1 FILLER_45_690 ();
 sg13g2_decap_4 FILLER_45_715 ();
 sg13g2_fill_2 FILLER_45_724 ();
 sg13g2_fill_2 FILLER_45_737 ();
 sg13g2_fill_1 FILLER_45_755 ();
 sg13g2_fill_2 FILLER_45_800 ();
 sg13g2_fill_2 FILLER_45_876 ();
 sg13g2_fill_1 FILLER_46_56 ();
 sg13g2_fill_1 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_96 ();
 sg13g2_fill_1 FILLER_46_101 ();
 sg13g2_fill_1 FILLER_46_112 ();
 sg13g2_fill_2 FILLER_46_176 ();
 sg13g2_fill_2 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_218 ();
 sg13g2_fill_2 FILLER_46_266 ();
 sg13g2_fill_2 FILLER_46_273 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_fill_1 FILLER_46_287 ();
 sg13g2_fill_2 FILLER_46_319 ();
 sg13g2_fill_2 FILLER_46_386 ();
 sg13g2_fill_1 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_462 ();
 sg13g2_fill_2 FILLER_46_472 ();
 sg13g2_fill_1 FILLER_46_478 ();
 sg13g2_fill_1 FILLER_46_482 ();
 sg13g2_fill_1 FILLER_46_536 ();
 sg13g2_fill_2 FILLER_46_542 ();
 sg13g2_fill_1 FILLER_46_548 ();
 sg13g2_fill_1 FILLER_46_593 ();
 sg13g2_fill_1 FILLER_46_626 ();
 sg13g2_fill_1 FILLER_46_631 ();
 sg13g2_decap_4 FILLER_46_668 ();
 sg13g2_fill_2 FILLER_46_689 ();
 sg13g2_fill_1 FILLER_46_726 ();
 sg13g2_fill_2 FILLER_46_756 ();
 sg13g2_fill_1 FILLER_46_772 ();
 sg13g2_fill_2 FILLER_46_777 ();
 sg13g2_fill_1 FILLER_46_779 ();
 sg13g2_fill_2 FILLER_46_798 ();
 sg13g2_fill_2 FILLER_46_810 ();
 sg13g2_fill_2 FILLER_46_826 ();
 sg13g2_fill_1 FILLER_46_828 ();
 sg13g2_fill_2 FILLER_46_875 ();
 sg13g2_fill_1 FILLER_46_877 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_27 ();
 sg13g2_fill_1 FILLER_47_38 ();
 sg13g2_fill_2 FILLER_47_59 ();
 sg13g2_fill_1 FILLER_47_155 ();
 sg13g2_fill_1 FILLER_47_213 ();
 sg13g2_fill_2 FILLER_47_227 ();
 sg13g2_fill_2 FILLER_47_257 ();
 sg13g2_fill_1 FILLER_47_269 ();
 sg13g2_fill_2 FILLER_47_326 ();
 sg13g2_fill_1 FILLER_47_328 ();
 sg13g2_fill_1 FILLER_47_386 ();
 sg13g2_fill_2 FILLER_47_408 ();
 sg13g2_decap_4 FILLER_47_432 ();
 sg13g2_fill_2 FILLER_47_436 ();
 sg13g2_fill_2 FILLER_47_441 ();
 sg13g2_fill_1 FILLER_47_443 ();
 sg13g2_fill_2 FILLER_47_448 ();
 sg13g2_fill_1 FILLER_47_450 ();
 sg13g2_fill_1 FILLER_47_455 ();
 sg13g2_fill_2 FILLER_47_461 ();
 sg13g2_fill_1 FILLER_47_467 ();
 sg13g2_decap_8 FILLER_47_472 ();
 sg13g2_fill_1 FILLER_47_479 ();
 sg13g2_fill_1 FILLER_47_484 ();
 sg13g2_fill_2 FILLER_47_489 ();
 sg13g2_fill_2 FILLER_47_495 ();
 sg13g2_fill_1 FILLER_47_497 ();
 sg13g2_fill_1 FILLER_47_515 ();
 sg13g2_fill_1 FILLER_47_521 ();
 sg13g2_fill_2 FILLER_47_566 ();
 sg13g2_fill_1 FILLER_47_568 ();
 sg13g2_fill_1 FILLER_47_574 ();
 sg13g2_fill_2 FILLER_47_610 ();
 sg13g2_fill_1 FILLER_47_612 ();
 sg13g2_fill_1 FILLER_47_633 ();
 sg13g2_fill_2 FILLER_47_674 ();
 sg13g2_fill_1 FILLER_47_676 ();
 sg13g2_fill_1 FILLER_47_688 ();
 sg13g2_fill_1 FILLER_47_693 ();
 sg13g2_fill_1 FILLER_47_699 ();
 sg13g2_fill_2 FILLER_47_717 ();
 sg13g2_fill_2 FILLER_47_727 ();
 sg13g2_fill_1 FILLER_47_729 ();
 sg13g2_fill_2 FILLER_47_789 ();
 sg13g2_fill_2 FILLER_47_817 ();
 sg13g2_fill_1 FILLER_47_849 ();
 sg13g2_fill_2 FILLER_47_876 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_1 FILLER_48_70 ();
 sg13g2_fill_1 FILLER_48_115 ();
 sg13g2_fill_1 FILLER_48_120 ();
 sg13g2_fill_2 FILLER_48_125 ();
 sg13g2_fill_1 FILLER_48_153 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_279 ();
 sg13g2_fill_1 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_313 ();
 sg13g2_fill_1 FILLER_48_319 ();
 sg13g2_fill_1 FILLER_48_325 ();
 sg13g2_fill_1 FILLER_48_336 ();
 sg13g2_fill_1 FILLER_48_345 ();
 sg13g2_fill_1 FILLER_48_350 ();
 sg13g2_fill_2 FILLER_48_361 ();
 sg13g2_fill_1 FILLER_48_370 ();
 sg13g2_fill_2 FILLER_48_375 ();
 sg13g2_decap_4 FILLER_48_384 ();
 sg13g2_fill_2 FILLER_48_418 ();
 sg13g2_fill_1 FILLER_48_424 ();
 sg13g2_fill_1 FILLER_48_446 ();
 sg13g2_fill_1 FILLER_48_457 ();
 sg13g2_fill_2 FILLER_48_466 ();
 sg13g2_fill_1 FILLER_48_468 ();
 sg13g2_decap_4 FILLER_48_474 ();
 sg13g2_fill_2 FILLER_48_517 ();
 sg13g2_fill_1 FILLER_48_595 ();
 sg13g2_fill_1 FILLER_48_601 ();
 sg13g2_fill_1 FILLER_48_610 ();
 sg13g2_fill_2 FILLER_48_624 ();
 sg13g2_fill_1 FILLER_48_626 ();
 sg13g2_fill_2 FILLER_48_635 ();
 sg13g2_fill_1 FILLER_48_637 ();
 sg13g2_fill_2 FILLER_48_710 ();
 sg13g2_fill_1 FILLER_48_712 ();
 sg13g2_fill_2 FILLER_48_751 ();
 sg13g2_fill_1 FILLER_48_770 ();
 sg13g2_fill_2 FILLER_48_776 ();
 sg13g2_fill_1 FILLER_48_778 ();
 sg13g2_fill_1 FILLER_48_829 ();
 sg13g2_fill_1 FILLER_48_840 ();
 sg13g2_fill_1 FILLER_48_877 ();
 sg13g2_fill_2 FILLER_49_81 ();
 sg13g2_fill_1 FILLER_49_127 ();
 sg13g2_fill_1 FILLER_49_190 ();
 sg13g2_fill_1 FILLER_49_241 ();
 sg13g2_fill_1 FILLER_49_353 ();
 sg13g2_fill_2 FILLER_49_395 ();
 sg13g2_fill_2 FILLER_49_446 ();
 sg13g2_fill_1 FILLER_49_448 ();
 sg13g2_fill_2 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_461 ();
 sg13g2_fill_2 FILLER_49_484 ();
 sg13g2_fill_1 FILLER_49_520 ();
 sg13g2_fill_1 FILLER_49_530 ();
 sg13g2_fill_1 FILLER_49_535 ();
 sg13g2_fill_1 FILLER_49_541 ();
 sg13g2_fill_1 FILLER_49_546 ();
 sg13g2_fill_2 FILLER_49_646 ();
 sg13g2_fill_1 FILLER_49_674 ();
 sg13g2_fill_2 FILLER_49_679 ();
 sg13g2_fill_1 FILLER_49_695 ();
 sg13g2_fill_1 FILLER_49_709 ();
 sg13g2_fill_1 FILLER_49_718 ();
 sg13g2_fill_2 FILLER_49_738 ();
 sg13g2_fill_2 FILLER_49_750 ();
 sg13g2_fill_1 FILLER_49_756 ();
 sg13g2_fill_1 FILLER_49_813 ();
 sg13g2_fill_1 FILLER_49_840 ();
 sg13g2_fill_2 FILLER_49_875 ();
 sg13g2_fill_1 FILLER_49_877 ();
 sg13g2_fill_1 FILLER_50_61 ();
 sg13g2_fill_2 FILLER_50_94 ();
 sg13g2_fill_1 FILLER_50_101 ();
 sg13g2_fill_1 FILLER_50_106 ();
 sg13g2_fill_1 FILLER_50_111 ();
 sg13g2_fill_2 FILLER_50_122 ();
 sg13g2_fill_2 FILLER_50_167 ();
 sg13g2_fill_1 FILLER_50_305 ();
 sg13g2_fill_1 FILLER_50_310 ();
 sg13g2_fill_1 FILLER_50_321 ();
 sg13g2_fill_2 FILLER_50_326 ();
 sg13g2_fill_2 FILLER_50_332 ();
 sg13g2_decap_4 FILLER_50_370 ();
 sg13g2_fill_1 FILLER_50_374 ();
 sg13g2_fill_1 FILLER_50_396 ();
 sg13g2_fill_2 FILLER_50_418 ();
 sg13g2_fill_1 FILLER_50_420 ();
 sg13g2_fill_2 FILLER_50_424 ();
 sg13g2_fill_1 FILLER_50_479 ();
 sg13g2_fill_2 FILLER_50_491 ();
 sg13g2_fill_1 FILLER_50_518 ();
 sg13g2_fill_1 FILLER_50_566 ();
 sg13g2_fill_1 FILLER_50_572 ();
 sg13g2_fill_1 FILLER_50_583 ();
 sg13g2_fill_2 FILLER_50_611 ();
 sg13g2_fill_1 FILLER_50_618 ();
 sg13g2_fill_2 FILLER_50_624 ();
 sg13g2_fill_2 FILLER_50_631 ();
 sg13g2_fill_2 FILLER_50_638 ();
 sg13g2_fill_1 FILLER_50_645 ();
 sg13g2_fill_1 FILLER_50_651 ();
 sg13g2_fill_1 FILLER_50_659 ();
 sg13g2_fill_1 FILLER_50_676 ();
 sg13g2_fill_1 FILLER_50_711 ();
 sg13g2_fill_2 FILLER_50_716 ();
 sg13g2_fill_1 FILLER_50_760 ();
 sg13g2_fill_2 FILLER_50_770 ();
 sg13g2_fill_2 FILLER_50_827 ();
 sg13g2_fill_2 FILLER_50_875 ();
 sg13g2_fill_1 FILLER_50_877 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_102 ();
 sg13g2_fill_1 FILLER_51_124 ();
 sg13g2_fill_1 FILLER_51_129 ();
 sg13g2_fill_2 FILLER_51_135 ();
 sg13g2_fill_2 FILLER_51_163 ();
 sg13g2_fill_2 FILLER_51_226 ();
 sg13g2_fill_1 FILLER_51_241 ();
 sg13g2_fill_1 FILLER_51_278 ();
 sg13g2_decap_8 FILLER_51_440 ();
 sg13g2_decap_4 FILLER_51_447 ();
 sg13g2_fill_1 FILLER_51_451 ();
 sg13g2_fill_1 FILLER_51_488 ();
 sg13g2_decap_4 FILLER_51_493 ();
 sg13g2_fill_2 FILLER_51_497 ();
 sg13g2_fill_1 FILLER_51_587 ();
 sg13g2_fill_1 FILLER_51_593 ();
 sg13g2_fill_1 FILLER_51_604 ();
 sg13g2_fill_2 FILLER_51_617 ();
 sg13g2_fill_1 FILLER_51_636 ();
 sg13g2_fill_2 FILLER_51_686 ();
 sg13g2_fill_1 FILLER_51_688 ();
 sg13g2_fill_1 FILLER_51_707 ();
 sg13g2_fill_1 FILLER_51_723 ();
 sg13g2_fill_1 FILLER_51_752 ();
 sg13g2_fill_1 FILLER_51_770 ();
 sg13g2_fill_2 FILLER_51_789 ();
 sg13g2_fill_2 FILLER_51_865 ();
 sg13g2_fill_2 FILLER_51_875 ();
 sg13g2_fill_1 FILLER_51_877 ();
 sg13g2_fill_2 FILLER_52_32 ();
 sg13g2_fill_1 FILLER_52_43 ();
 sg13g2_fill_2 FILLER_52_58 ();
 sg13g2_fill_1 FILLER_52_91 ();
 sg13g2_fill_1 FILLER_52_123 ();
 sg13g2_fill_1 FILLER_52_131 ();
 sg13g2_fill_1 FILLER_52_159 ();
 sg13g2_fill_1 FILLER_52_169 ();
 sg13g2_fill_1 FILLER_52_177 ();
 sg13g2_fill_1 FILLER_52_241 ();
 sg13g2_fill_1 FILLER_52_250 ();
 sg13g2_fill_2 FILLER_52_367 ();
 sg13g2_fill_2 FILLER_52_390 ();
 sg13g2_fill_1 FILLER_52_392 ();
 sg13g2_fill_2 FILLER_52_406 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_fill_1 FILLER_52_414 ();
 sg13g2_fill_2 FILLER_52_436 ();
 sg13g2_fill_2 FILLER_52_451 ();
 sg13g2_fill_1 FILLER_52_457 ();
 sg13g2_fill_2 FILLER_52_480 ();
 sg13g2_fill_1 FILLER_52_508 ();
 sg13g2_fill_1 FILLER_52_513 ();
 sg13g2_fill_1 FILLER_52_518 ();
 sg13g2_fill_2 FILLER_52_524 ();
 sg13g2_fill_2 FILLER_52_531 ();
 sg13g2_fill_2 FILLER_52_566 ();
 sg13g2_fill_1 FILLER_52_576 ();
 sg13g2_fill_2 FILLER_52_603 ();
 sg13g2_fill_2 FILLER_52_614 ();
 sg13g2_fill_2 FILLER_52_624 ();
 sg13g2_fill_1 FILLER_52_626 ();
 sg13g2_fill_1 FILLER_52_630 ();
 sg13g2_fill_1 FILLER_52_639 ();
 sg13g2_fill_2 FILLER_52_669 ();
 sg13g2_fill_2 FILLER_52_694 ();
 sg13g2_fill_2 FILLER_52_708 ();
 sg13g2_fill_1 FILLER_52_710 ();
 sg13g2_fill_1 FILLER_52_727 ();
 sg13g2_fill_1 FILLER_52_738 ();
 sg13g2_fill_1 FILLER_52_747 ();
 sg13g2_fill_1 FILLER_52_775 ();
 sg13g2_fill_1 FILLER_52_877 ();
 sg13g2_fill_2 FILLER_53_66 ();
 sg13g2_fill_2 FILLER_53_76 ();
 sg13g2_fill_1 FILLER_53_78 ();
 sg13g2_fill_2 FILLER_53_100 ();
 sg13g2_fill_1 FILLER_53_102 ();
 sg13g2_fill_1 FILLER_53_107 ();
 sg13g2_fill_1 FILLER_53_166 ();
 sg13g2_fill_1 FILLER_53_211 ();
 sg13g2_fill_1 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_fill_1 FILLER_53_317 ();
 sg13g2_fill_2 FILLER_53_323 ();
 sg13g2_fill_1 FILLER_53_344 ();
 sg13g2_fill_1 FILLER_53_361 ();
 sg13g2_fill_1 FILLER_53_367 ();
 sg13g2_fill_2 FILLER_53_383 ();
 sg13g2_fill_1 FILLER_53_398 ();
 sg13g2_fill_1 FILLER_53_404 ();
 sg13g2_fill_1 FILLER_53_410 ();
 sg13g2_fill_2 FILLER_53_415 ();
 sg13g2_fill_1 FILLER_53_422 ();
 sg13g2_fill_1 FILLER_53_427 ();
 sg13g2_fill_1 FILLER_53_434 ();
 sg13g2_fill_2 FILLER_53_470 ();
 sg13g2_fill_1 FILLER_53_490 ();
 sg13g2_fill_1 FILLER_53_552 ();
 sg13g2_fill_1 FILLER_53_557 ();
 sg13g2_fill_1 FILLER_53_562 ();
 sg13g2_fill_2 FILLER_53_568 ();
 sg13g2_fill_1 FILLER_53_616 ();
 sg13g2_fill_2 FILLER_53_632 ();
 sg13g2_fill_1 FILLER_53_653 ();
 sg13g2_fill_1 FILLER_53_667 ();
 sg13g2_fill_2 FILLER_53_687 ();
 sg13g2_fill_1 FILLER_53_715 ();
 sg13g2_fill_1 FILLER_53_747 ();
 sg13g2_fill_1 FILLER_53_753 ();
 sg13g2_fill_2 FILLER_53_790 ();
 sg13g2_fill_2 FILLER_53_818 ();
 sg13g2_fill_2 FILLER_53_850 ();
 sg13g2_fill_1 FILLER_54_144 ();
 sg13g2_fill_1 FILLER_54_204 ();
 sg13g2_fill_2 FILLER_54_266 ();
 sg13g2_fill_1 FILLER_54_278 ();
 sg13g2_fill_1 FILLER_54_289 ();
 sg13g2_fill_1 FILLER_54_301 ();
 sg13g2_fill_1 FILLER_54_306 ();
 sg13g2_fill_1 FILLER_54_344 ();
 sg13g2_fill_1 FILLER_54_371 ();
 sg13g2_fill_1 FILLER_54_398 ();
 sg13g2_fill_1 FILLER_54_407 ();
 sg13g2_fill_2 FILLER_54_414 ();
 sg13g2_fill_1 FILLER_54_416 ();
 sg13g2_fill_2 FILLER_54_437 ();
 sg13g2_fill_1 FILLER_54_549 ();
 sg13g2_fill_1 FILLER_54_555 ();
 sg13g2_fill_1 FILLER_54_569 ();
 sg13g2_fill_1 FILLER_54_575 ();
 sg13g2_fill_1 FILLER_54_584 ();
 sg13g2_fill_1 FILLER_54_589 ();
 sg13g2_fill_2 FILLER_54_598 ();
 sg13g2_fill_1 FILLER_54_618 ();
 sg13g2_fill_2 FILLER_54_640 ();
 sg13g2_fill_1 FILLER_54_667 ();
 sg13g2_fill_1 FILLER_54_698 ();
 sg13g2_fill_2 FILLER_54_716 ();
 sg13g2_fill_2 FILLER_54_739 ();
 sg13g2_fill_2 FILLER_54_803 ();
 sg13g2_fill_1 FILLER_54_813 ();
 sg13g2_fill_2 FILLER_54_844 ();
 sg13g2_fill_2 FILLER_54_875 ();
 sg13g2_fill_1 FILLER_54_877 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_6 ();
 sg13g2_fill_1 FILLER_55_8 ();
 sg13g2_fill_1 FILLER_55_64 ();
 sg13g2_fill_2 FILLER_55_101 ();
 sg13g2_fill_2 FILLER_55_112 ();
 sg13g2_fill_1 FILLER_55_114 ();
 sg13g2_fill_2 FILLER_55_175 ();
 sg13g2_fill_1 FILLER_55_181 ();
 sg13g2_fill_1 FILLER_55_222 ();
 sg13g2_fill_2 FILLER_55_233 ();
 sg13g2_fill_2 FILLER_55_258 ();
 sg13g2_fill_1 FILLER_55_260 ();
 sg13g2_fill_1 FILLER_55_295 ();
 sg13g2_fill_1 FILLER_55_301 ();
 sg13g2_fill_2 FILLER_55_334 ();
 sg13g2_fill_2 FILLER_55_353 ();
 sg13g2_fill_1 FILLER_55_355 ();
 sg13g2_fill_1 FILLER_55_361 ();
 sg13g2_fill_1 FILLER_55_392 ();
 sg13g2_fill_1 FILLER_55_419 ();
 sg13g2_fill_1 FILLER_55_454 ();
 sg13g2_fill_2 FILLER_55_459 ();
 sg13g2_fill_2 FILLER_55_465 ();
 sg13g2_fill_1 FILLER_55_467 ();
 sg13g2_fill_2 FILLER_55_504 ();
 sg13g2_fill_2 FILLER_55_518 ();
 sg13g2_fill_1 FILLER_55_520 ();
 sg13g2_fill_2 FILLER_55_533 ();
 sg13g2_fill_2 FILLER_55_540 ();
 sg13g2_fill_2 FILLER_55_558 ();
 sg13g2_fill_2 FILLER_55_602 ();
 sg13g2_fill_2 FILLER_55_675 ();
 sg13g2_fill_1 FILLER_55_677 ();
 sg13g2_fill_2 FILLER_55_699 ();
 sg13g2_fill_1 FILLER_55_701 ();
 sg13g2_fill_1 FILLER_55_707 ();
 sg13g2_fill_1 FILLER_55_717 ();
 sg13g2_fill_2 FILLER_55_744 ();
 sg13g2_fill_1 FILLER_55_746 ();
 sg13g2_fill_2 FILLER_55_755 ();
 sg13g2_fill_1 FILLER_55_786 ();
 sg13g2_fill_2 FILLER_56_26 ();
 sg13g2_fill_1 FILLER_56_28 ();
 sg13g2_fill_2 FILLER_56_59 ();
 sg13g2_fill_1 FILLER_56_61 ();
 sg13g2_fill_1 FILLER_56_150 ();
 sg13g2_fill_2 FILLER_56_155 ();
 sg13g2_fill_1 FILLER_56_212 ();
 sg13g2_fill_1 FILLER_56_239 ();
 sg13g2_fill_1 FILLER_56_245 ();
 sg13g2_fill_1 FILLER_56_251 ();
 sg13g2_fill_2 FILLER_56_257 ();
 sg13g2_fill_1 FILLER_56_263 ();
 sg13g2_fill_1 FILLER_56_272 ();
 sg13g2_fill_2 FILLER_56_303 ();
 sg13g2_fill_1 FILLER_56_338 ();
 sg13g2_fill_1 FILLER_56_361 ();
 sg13g2_fill_2 FILLER_56_400 ();
 sg13g2_fill_1 FILLER_56_434 ();
 sg13g2_fill_1 FILLER_56_448 ();
 sg13g2_fill_1 FILLER_56_453 ();
 sg13g2_fill_2 FILLER_56_517 ();
 sg13g2_fill_1 FILLER_56_519 ();
 sg13g2_fill_1 FILLER_56_525 ();
 sg13g2_fill_2 FILLER_56_539 ();
 sg13g2_fill_1 FILLER_56_541 ();
 sg13g2_fill_2 FILLER_56_561 ();
 sg13g2_fill_1 FILLER_56_624 ();
 sg13g2_fill_2 FILLER_56_762 ();
 sg13g2_fill_2 FILLER_56_809 ();
 sg13g2_fill_1 FILLER_56_811 ();
 sg13g2_fill_1 FILLER_56_822 ();
 sg13g2_fill_2 FILLER_56_833 ();
 sg13g2_decap_8 FILLER_56_869 ();
 sg13g2_fill_2 FILLER_56_876 ();
 sg13g2_fill_1 FILLER_57_61 ();
 sg13g2_fill_1 FILLER_57_88 ();
 sg13g2_fill_1 FILLER_57_127 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_fill_1 FILLER_57_157 ();
 sg13g2_fill_1 FILLER_57_162 ();
 sg13g2_fill_2 FILLER_57_182 ();
 sg13g2_fill_1 FILLER_57_188 ();
 sg13g2_fill_2 FILLER_57_239 ();
 sg13g2_fill_1 FILLER_57_241 ();
 sg13g2_fill_1 FILLER_57_281 ();
 sg13g2_fill_1 FILLER_57_330 ();
 sg13g2_decap_4 FILLER_57_374 ();
 sg13g2_fill_1 FILLER_57_382 ();
 sg13g2_fill_2 FILLER_57_396 ();
 sg13g2_fill_2 FILLER_57_428 ();
 sg13g2_fill_1 FILLER_57_435 ();
 sg13g2_decap_4 FILLER_57_461 ();
 sg13g2_fill_2 FILLER_57_476 ();
 sg13g2_fill_1 FILLER_57_483 ();
 sg13g2_fill_1 FILLER_57_501 ();
 sg13g2_fill_2 FILLER_57_515 ();
 sg13g2_fill_1 FILLER_57_517 ();
 sg13g2_fill_1 FILLER_57_538 ();
 sg13g2_fill_1 FILLER_57_552 ();
 sg13g2_fill_2 FILLER_57_567 ();
 sg13g2_fill_2 FILLER_57_578 ();
 sg13g2_fill_2 FILLER_57_626 ();
 sg13g2_fill_1 FILLER_57_645 ();
 sg13g2_fill_2 FILLER_57_650 ();
 sg13g2_fill_1 FILLER_57_652 ();
 sg13g2_fill_2 FILLER_57_673 ();
 sg13g2_fill_1 FILLER_57_675 ();
 sg13g2_fill_2 FILLER_57_680 ();
 sg13g2_fill_1 FILLER_57_732 ();
 sg13g2_fill_1 FILLER_57_784 ();
 sg13g2_fill_2 FILLER_57_795 ();
 sg13g2_fill_2 FILLER_57_807 ();
 sg13g2_decap_8 FILLER_57_871 ();
 sg13g2_fill_2 FILLER_58_14 ();
 sg13g2_fill_1 FILLER_58_34 ();
 sg13g2_fill_1 FILLER_58_96 ();
 sg13g2_fill_1 FILLER_58_101 ();
 sg13g2_fill_2 FILLER_58_135 ();
 sg13g2_fill_2 FILLER_58_141 ();
 sg13g2_fill_1 FILLER_58_147 ();
 sg13g2_fill_1 FILLER_58_200 ();
 sg13g2_fill_1 FILLER_58_206 ();
 sg13g2_fill_1 FILLER_58_212 ();
 sg13g2_fill_1 FILLER_58_223 ();
 sg13g2_fill_1 FILLER_58_298 ();
 sg13g2_fill_2 FILLER_58_385 ();
 sg13g2_fill_1 FILLER_58_387 ();
 sg13g2_fill_2 FILLER_58_412 ();
 sg13g2_fill_2 FILLER_58_475 ();
 sg13g2_fill_2 FILLER_58_552 ();
 sg13g2_fill_1 FILLER_58_587 ();
 sg13g2_fill_2 FILLER_58_593 ();
 sg13g2_fill_1 FILLER_58_595 ();
 sg13g2_fill_1 FILLER_58_627 ();
 sg13g2_fill_1 FILLER_58_659 ();
 sg13g2_fill_2 FILLER_58_686 ();
 sg13g2_fill_2 FILLER_58_696 ();
 sg13g2_fill_2 FILLER_58_711 ();
 sg13g2_fill_2 FILLER_58_836 ();
 sg13g2_fill_1 FILLER_58_848 ();
 sg13g2_fill_2 FILLER_58_875 ();
 sg13g2_fill_1 FILLER_58_877 ();
 sg13g2_fill_2 FILLER_59_64 ();
 sg13g2_fill_2 FILLER_59_119 ();
 sg13g2_fill_1 FILLER_59_121 ();
 sg13g2_fill_1 FILLER_59_252 ();
 sg13g2_fill_1 FILLER_59_283 ();
 sg13g2_fill_1 FILLER_59_289 ();
 sg13g2_fill_2 FILLER_59_346 ();
 sg13g2_fill_2 FILLER_59_352 ();
 sg13g2_fill_2 FILLER_59_360 ();
 sg13g2_fill_2 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_435 ();
 sg13g2_fill_1 FILLER_59_446 ();
 sg13g2_decap_4 FILLER_59_450 ();
 sg13g2_fill_2 FILLER_59_454 ();
 sg13g2_fill_2 FILLER_59_460 ();
 sg13g2_decap_8 FILLER_59_470 ();
 sg13g2_fill_2 FILLER_59_481 ();
 sg13g2_fill_1 FILLER_59_483 ();
 sg13g2_fill_1 FILLER_59_502 ();
 sg13g2_fill_1 FILLER_59_511 ();
 sg13g2_fill_1 FILLER_59_520 ();
 sg13g2_fill_1 FILLER_59_533 ();
 sg13g2_fill_2 FILLER_59_568 ();
 sg13g2_fill_1 FILLER_59_570 ();
 sg13g2_fill_1 FILLER_59_599 ();
 sg13g2_fill_1 FILLER_59_626 ();
 sg13g2_fill_1 FILLER_59_640 ();
 sg13g2_fill_2 FILLER_59_665 ();
 sg13g2_fill_1 FILLER_59_698 ();
 sg13g2_fill_1 FILLER_59_704 ();
 sg13g2_fill_1 FILLER_59_774 ();
 sg13g2_fill_1 FILLER_59_793 ();
 sg13g2_fill_2 FILLER_59_825 ();
 sg13g2_decap_8 FILLER_59_867 ();
 sg13g2_decap_4 FILLER_59_874 ();
 sg13g2_fill_2 FILLER_60_30 ();
 sg13g2_fill_1 FILLER_60_32 ();
 sg13g2_fill_1 FILLER_60_84 ();
 sg13g2_fill_1 FILLER_60_122 ();
 sg13g2_fill_1 FILLER_60_128 ();
 sg13g2_fill_1 FILLER_60_183 ();
 sg13g2_fill_1 FILLER_60_189 ();
 sg13g2_fill_1 FILLER_60_195 ();
 sg13g2_fill_2 FILLER_60_209 ();
 sg13g2_fill_1 FILLER_60_224 ();
 sg13g2_fill_2 FILLER_60_235 ();
 sg13g2_fill_1 FILLER_60_237 ();
 sg13g2_fill_1 FILLER_60_325 ();
 sg13g2_fill_1 FILLER_60_379 ();
 sg13g2_fill_1 FILLER_60_389 ();
 sg13g2_fill_2 FILLER_60_451 ();
 sg13g2_decap_4 FILLER_60_465 ();
 sg13g2_fill_2 FILLER_60_469 ();
 sg13g2_decap_4 FILLER_60_476 ();
 sg13g2_fill_1 FILLER_60_480 ();
 sg13g2_fill_2 FILLER_60_527 ();
 sg13g2_fill_2 FILLER_60_567 ();
 sg13g2_fill_1 FILLER_60_569 ();
 sg13g2_fill_2 FILLER_60_582 ();
 sg13g2_fill_1 FILLER_60_584 ();
 sg13g2_fill_1 FILLER_60_624 ();
 sg13g2_fill_1 FILLER_60_632 ();
 sg13g2_fill_2 FILLER_60_688 ();
 sg13g2_fill_1 FILLER_60_748 ();
 sg13g2_decap_8 FILLER_60_863 ();
 sg13g2_decap_8 FILLER_60_870 ();
 sg13g2_fill_1 FILLER_60_877 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_31 ();
 sg13g2_fill_1 FILLER_61_33 ();
 sg13g2_fill_1 FILLER_61_38 ();
 sg13g2_fill_2 FILLER_61_55 ();
 sg13g2_fill_1 FILLER_61_151 ();
 sg13g2_fill_1 FILLER_61_178 ();
 sg13g2_fill_1 FILLER_61_205 ();
 sg13g2_fill_2 FILLER_61_213 ();
 sg13g2_fill_1 FILLER_61_242 ();
 sg13g2_fill_1 FILLER_61_309 ();
 sg13g2_fill_2 FILLER_61_338 ();
 sg13g2_fill_2 FILLER_61_378 ();
 sg13g2_fill_1 FILLER_61_380 ();
 sg13g2_fill_1 FILLER_61_419 ();
 sg13g2_fill_1 FILLER_61_494 ();
 sg13g2_fill_1 FILLER_61_499 ();
 sg13g2_fill_2 FILLER_61_557 ();
 sg13g2_fill_2 FILLER_61_573 ();
 sg13g2_fill_1 FILLER_61_575 ();
 sg13g2_fill_1 FILLER_61_581 ();
 sg13g2_fill_1 FILLER_61_587 ();
 sg13g2_fill_2 FILLER_61_593 ();
 sg13g2_fill_1 FILLER_61_619 ();
 sg13g2_fill_2 FILLER_61_689 ();
 sg13g2_fill_1 FILLER_61_697 ();
 sg13g2_fill_1 FILLER_61_760 ();
 sg13g2_fill_1 FILLER_61_851 ();
 sg13g2_fill_1 FILLER_62_34 ();
 sg13g2_fill_1 FILLER_62_61 ();
 sg13g2_fill_1 FILLER_62_90 ();
 sg13g2_fill_1 FILLER_62_149 ();
 sg13g2_fill_2 FILLER_62_155 ();
 sg13g2_fill_1 FILLER_62_162 ();
 sg13g2_fill_2 FILLER_62_167 ();
 sg13g2_fill_2 FILLER_62_174 ();
 sg13g2_fill_2 FILLER_62_220 ();
 sg13g2_fill_2 FILLER_62_301 ();
 sg13g2_fill_1 FILLER_62_307 ();
 sg13g2_fill_1 FILLER_62_321 ();
 sg13g2_fill_1 FILLER_62_332 ();
 sg13g2_fill_2 FILLER_62_383 ();
 sg13g2_fill_1 FILLER_62_385 ();
 sg13g2_decap_4 FILLER_62_398 ();
 sg13g2_fill_1 FILLER_62_412 ();
 sg13g2_fill_1 FILLER_62_433 ();
 sg13g2_fill_1 FILLER_62_444 ();
 sg13g2_fill_1 FILLER_62_450 ();
 sg13g2_fill_2 FILLER_62_456 ();
 sg13g2_fill_2 FILLER_62_462 ();
 sg13g2_fill_2 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_498 ();
 sg13g2_fill_1 FILLER_62_514 ();
 sg13g2_fill_1 FILLER_62_520 ();
 sg13g2_fill_1 FILLER_62_614 ();
 sg13g2_fill_1 FILLER_62_652 ();
 sg13g2_fill_1 FILLER_62_663 ();
 sg13g2_fill_2 FILLER_62_669 ();
 sg13g2_fill_1 FILLER_62_676 ();
 sg13g2_fill_1 FILLER_62_703 ();
 sg13g2_fill_1 FILLER_62_709 ();
 sg13g2_fill_1 FILLER_62_720 ();
 sg13g2_fill_2 FILLER_62_762 ();
 sg13g2_fill_1 FILLER_62_800 ();
 sg13g2_fill_1 FILLER_62_849 ();
 sg13g2_decap_8 FILLER_62_857 ();
 sg13g2_decap_4 FILLER_62_864 ();
 sg13g2_fill_2 FILLER_62_876 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_20 ();
 sg13g2_fill_1 FILLER_63_71 ();
 sg13g2_fill_1 FILLER_63_106 ();
 sg13g2_fill_2 FILLER_63_112 ();
 sg13g2_fill_2 FILLER_63_119 ();
 sg13g2_fill_2 FILLER_63_125 ();
 sg13g2_fill_1 FILLER_63_127 ();
 sg13g2_fill_2 FILLER_63_192 ();
 sg13g2_fill_2 FILLER_63_207 ();
 sg13g2_fill_2 FILLER_63_233 ();
 sg13g2_fill_1 FILLER_63_313 ();
 sg13g2_fill_1 FILLER_63_324 ();
 sg13g2_fill_2 FILLER_63_343 ();
 sg13g2_fill_2 FILLER_63_351 ();
 sg13g2_fill_2 FILLER_63_385 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_1 FILLER_63_417 ();
 sg13g2_fill_2 FILLER_63_435 ();
 sg13g2_fill_1 FILLER_63_437 ();
 sg13g2_fill_1 FILLER_63_443 ();
 sg13g2_fill_2 FILLER_63_450 ();
 sg13g2_fill_2 FILLER_63_478 ();
 sg13g2_fill_2 FILLER_63_506 ();
 sg13g2_fill_1 FILLER_63_573 ();
 sg13g2_fill_1 FILLER_63_579 ();
 sg13g2_fill_1 FILLER_63_585 ();
 sg13g2_fill_1 FILLER_63_595 ();
 sg13g2_fill_2 FILLER_63_668 ();
 sg13g2_fill_2 FILLER_63_744 ();
 sg13g2_fill_2 FILLER_63_772 ();
 sg13g2_fill_2 FILLER_63_804 ();
 sg13g2_fill_1 FILLER_63_806 ();
 sg13g2_fill_1 FILLER_63_851 ();
 sg13g2_fill_1 FILLER_64_112 ();
 sg13g2_fill_2 FILLER_64_159 ();
 sg13g2_fill_2 FILLER_64_199 ();
 sg13g2_fill_1 FILLER_64_245 ();
 sg13g2_fill_1 FILLER_64_254 ();
 sg13g2_fill_1 FILLER_64_281 ();
 sg13g2_fill_2 FILLER_64_287 ();
 sg13g2_fill_1 FILLER_64_360 ();
 sg13g2_fill_2 FILLER_64_366 ();
 sg13g2_decap_8 FILLER_64_408 ();
 sg13g2_fill_1 FILLER_64_432 ();
 sg13g2_decap_4 FILLER_64_469 ();
 sg13g2_fill_2 FILLER_64_473 ();
 sg13g2_fill_2 FILLER_64_484 ();
 sg13g2_fill_2 FILLER_64_490 ();
 sg13g2_fill_1 FILLER_64_549 ();
 sg13g2_fill_1 FILLER_64_554 ();
 sg13g2_fill_2 FILLER_64_616 ();
 sg13g2_fill_2 FILLER_64_622 ();
 sg13g2_fill_1 FILLER_64_624 ();
 sg13g2_fill_1 FILLER_64_649 ();
 sg13g2_fill_2 FILLER_64_668 ();
 sg13g2_fill_1 FILLER_64_722 ();
 sg13g2_fill_2 FILLER_64_759 ();
 sg13g2_fill_1 FILLER_64_771 ();
 sg13g2_fill_1 FILLER_64_798 ();
 sg13g2_fill_1 FILLER_64_841 ();
 sg13g2_fill_1 FILLER_64_855 ();
 sg13g2_fill_2 FILLER_64_876 ();
 sg13g2_fill_1 FILLER_65_57 ();
 sg13g2_fill_1 FILLER_65_98 ();
 sg13g2_fill_1 FILLER_65_103 ();
 sg13g2_fill_1 FILLER_65_109 ();
 sg13g2_fill_1 FILLER_65_114 ();
 sg13g2_fill_2 FILLER_65_156 ();
 sg13g2_fill_2 FILLER_65_168 ();
 sg13g2_fill_1 FILLER_65_170 ();
 sg13g2_fill_1 FILLER_65_197 ();
 sg13g2_fill_1 FILLER_65_203 ();
 sg13g2_fill_1 FILLER_65_235 ();
 sg13g2_fill_1 FILLER_65_297 ();
 sg13g2_fill_2 FILLER_65_325 ();
 sg13g2_fill_1 FILLER_65_342 ();
 sg13g2_fill_1 FILLER_65_357 ();
 sg13g2_fill_2 FILLER_65_399 ();
 sg13g2_fill_1 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_426 ();
 sg13g2_fill_1 FILLER_65_432 ();
 sg13g2_fill_1 FILLER_65_469 ();
 sg13g2_fill_2 FILLER_65_501 ();
 sg13g2_fill_1 FILLER_65_510 ();
 sg13g2_fill_1 FILLER_65_541 ();
 sg13g2_fill_2 FILLER_65_582 ();
 sg13g2_fill_1 FILLER_65_589 ();
 sg13g2_fill_1 FILLER_65_595 ();
 sg13g2_fill_2 FILLER_65_604 ();
 sg13g2_fill_1 FILLER_65_615 ();
 sg13g2_fill_2 FILLER_65_640 ();
 sg13g2_fill_1 FILLER_65_647 ();
 sg13g2_fill_1 FILLER_65_653 ();
 sg13g2_fill_1 FILLER_65_664 ();
 sg13g2_fill_1 FILLER_65_695 ();
 sg13g2_fill_1 FILLER_65_752 ();
 sg13g2_fill_1 FILLER_65_791 ();
 sg13g2_fill_1 FILLER_65_850 ();
 sg13g2_fill_1 FILLER_65_877 ();
 sg13g2_fill_1 FILLER_66_73 ();
 sg13g2_fill_1 FILLER_66_79 ();
 sg13g2_fill_2 FILLER_66_85 ();
 sg13g2_fill_1 FILLER_66_97 ();
 sg13g2_fill_1 FILLER_66_103 ();
 sg13g2_fill_1 FILLER_66_109 ();
 sg13g2_fill_2 FILLER_66_180 ();
 sg13g2_fill_1 FILLER_66_182 ();
 sg13g2_fill_2 FILLER_66_239 ();
 sg13g2_fill_1 FILLER_66_331 ();
 sg13g2_fill_1 FILLER_66_355 ();
 sg13g2_fill_2 FILLER_66_440 ();
 sg13g2_fill_1 FILLER_66_472 ();
 sg13g2_fill_2 FILLER_66_477 ();
 sg13g2_fill_1 FILLER_66_483 ();
 sg13g2_fill_2 FILLER_66_489 ();
 sg13g2_fill_2 FILLER_66_500 ();
 sg13g2_fill_1 FILLER_66_512 ();
 sg13g2_fill_2 FILLER_66_522 ();
 sg13g2_fill_2 FILLER_66_568 ();
 sg13g2_fill_2 FILLER_66_610 ();
 sg13g2_fill_1 FILLER_66_612 ();
 sg13g2_fill_2 FILLER_66_666 ();
 sg13g2_fill_2 FILLER_66_684 ();
 sg13g2_fill_1 FILLER_66_691 ();
 sg13g2_fill_1 FILLER_66_700 ();
 sg13g2_fill_2 FILLER_66_765 ();
 sg13g2_fill_1 FILLER_66_767 ();
 sg13g2_fill_1 FILLER_66_799 ();
 sg13g2_fill_2 FILLER_66_820 ();
 sg13g2_fill_1 FILLER_66_822 ();
 sg13g2_fill_2 FILLER_66_832 ();
 sg13g2_fill_2 FILLER_67_43 ();
 sg13g2_fill_1 FILLER_67_127 ();
 sg13g2_fill_2 FILLER_67_141 ();
 sg13g2_fill_1 FILLER_67_143 ();
 sg13g2_fill_2 FILLER_67_165 ();
 sg13g2_fill_1 FILLER_67_251 ();
 sg13g2_fill_1 FILLER_67_260 ();
 sg13g2_fill_1 FILLER_67_291 ();
 sg13g2_fill_1 FILLER_67_303 ();
 sg13g2_fill_2 FILLER_67_320 ();
 sg13g2_fill_1 FILLER_67_422 ();
 sg13g2_fill_1 FILLER_67_427 ();
 sg13g2_fill_1 FILLER_67_441 ();
 sg13g2_fill_1 FILLER_67_447 ();
 sg13g2_fill_1 FILLER_67_452 ();
 sg13g2_fill_2 FILLER_67_494 ();
 sg13g2_fill_1 FILLER_67_502 ();
 sg13g2_fill_1 FILLER_67_508 ();
 sg13g2_fill_1 FILLER_67_518 ();
 sg13g2_fill_1 FILLER_67_523 ();
 sg13g2_fill_1 FILLER_67_529 ();
 sg13g2_fill_2 FILLER_67_535 ();
 sg13g2_fill_2 FILLER_67_581 ();
 sg13g2_fill_2 FILLER_67_596 ();
 sg13g2_fill_2 FILLER_67_634 ();
 sg13g2_fill_1 FILLER_67_636 ();
 sg13g2_fill_2 FILLER_67_729 ();
 sg13g2_fill_2 FILLER_67_761 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_5 ();
 sg13g2_fill_1 FILLER_68_31 ();
 sg13g2_fill_2 FILLER_68_61 ();
 sg13g2_fill_2 FILLER_68_73 ();
 sg13g2_fill_2 FILLER_68_89 ();
 sg13g2_fill_1 FILLER_68_121 ();
 sg13g2_fill_2 FILLER_68_152 ();
 sg13g2_fill_2 FILLER_68_188 ();
 sg13g2_fill_1 FILLER_68_270 ();
 sg13g2_fill_2 FILLER_68_302 ();
 sg13g2_fill_2 FILLER_68_309 ();
 sg13g2_fill_2 FILLER_68_347 ();
 sg13g2_fill_1 FILLER_68_375 ();
 sg13g2_fill_2 FILLER_68_380 ();
 sg13g2_fill_1 FILLER_68_422 ();
 sg13g2_fill_1 FILLER_68_433 ();
 sg13g2_fill_1 FILLER_68_438 ();
 sg13g2_fill_1 FILLER_68_448 ();
 sg13g2_fill_1 FILLER_68_453 ();
 sg13g2_fill_1 FILLER_68_458 ();
 sg13g2_fill_1 FILLER_68_469 ();
 sg13g2_fill_1 FILLER_68_504 ();
 sg13g2_fill_1 FILLER_68_612 ();
 sg13g2_fill_2 FILLER_68_676 ();
 sg13g2_fill_2 FILLER_68_690 ();
 sg13g2_fill_1 FILLER_68_705 ();
 sg13g2_fill_1 FILLER_68_741 ();
 sg13g2_fill_1 FILLER_68_778 ();
 sg13g2_fill_1 FILLER_68_818 ();
 sg13g2_fill_1 FILLER_68_827 ();
 sg13g2_fill_1 FILLER_68_840 ();
 sg13g2_fill_1 FILLER_69_34 ();
 sg13g2_fill_1 FILLER_69_91 ();
 sg13g2_fill_2 FILLER_69_105 ();
 sg13g2_fill_2 FILLER_69_133 ();
 sg13g2_fill_2 FILLER_69_169 ();
 sg13g2_fill_1 FILLER_69_197 ();
 sg13g2_fill_2 FILLER_69_243 ();
 sg13g2_fill_1 FILLER_69_285 ();
 sg13g2_fill_1 FILLER_69_312 ();
 sg13g2_fill_2 FILLER_69_353 ();
 sg13g2_fill_1 FILLER_69_364 ();
 sg13g2_fill_2 FILLER_69_370 ();
 sg13g2_fill_1 FILLER_69_372 ();
 sg13g2_fill_1 FILLER_69_391 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_fill_2 FILLER_69_418 ();
 sg13g2_fill_1 FILLER_69_438 ();
 sg13g2_fill_1 FILLER_69_443 ();
 sg13g2_fill_1 FILLER_69_449 ();
 sg13g2_fill_1 FILLER_69_476 ();
 sg13g2_fill_1 FILLER_69_501 ();
 sg13g2_fill_1 FILLER_69_532 ();
 sg13g2_fill_1 FILLER_69_538 ();
 sg13g2_fill_2 FILLER_69_578 ();
 sg13g2_fill_1 FILLER_69_580 ();
 sg13g2_fill_2 FILLER_69_757 ();
 sg13g2_fill_1 FILLER_69_759 ();
 sg13g2_fill_1 FILLER_69_770 ();
 sg13g2_fill_2 FILLER_69_815 ();
 sg13g2_fill_1 FILLER_69_847 ();
 sg13g2_fill_1 FILLER_70_93 ();
 sg13g2_fill_1 FILLER_70_104 ();
 sg13g2_fill_1 FILLER_70_110 ();
 sg13g2_fill_1 FILLER_70_116 ();
 sg13g2_fill_2 FILLER_70_124 ();
 sg13g2_fill_1 FILLER_70_131 ();
 sg13g2_fill_1 FILLER_70_141 ();
 sg13g2_fill_1 FILLER_70_147 ();
 sg13g2_fill_1 FILLER_70_226 ();
 sg13g2_fill_1 FILLER_70_232 ();
 sg13g2_fill_2 FILLER_70_242 ();
 sg13g2_fill_2 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_70_401 ();
 sg13g2_fill_2 FILLER_70_433 ();
 sg13g2_decap_8 FILLER_70_464 ();
 sg13g2_decap_4 FILLER_70_471 ();
 sg13g2_fill_1 FILLER_70_475 ();
 sg13g2_fill_1 FILLER_70_526 ();
 sg13g2_fill_1 FILLER_70_567 ();
 sg13g2_fill_1 FILLER_70_590 ();
 sg13g2_fill_2 FILLER_70_604 ();
 sg13g2_fill_1 FILLER_70_606 ();
 sg13g2_fill_2 FILLER_70_624 ();
 sg13g2_fill_1 FILLER_70_626 ();
 sg13g2_fill_2 FILLER_70_650 ();
 sg13g2_fill_1 FILLER_70_672 ();
 sg13g2_fill_1 FILLER_70_692 ();
 sg13g2_fill_2 FILLER_70_707 ();
 sg13g2_fill_2 FILLER_70_723 ();
 sg13g2_fill_1 FILLER_70_730 ();
 sg13g2_fill_2 FILLER_70_741 ();
 sg13g2_fill_1 FILLER_70_757 ();
 sg13g2_fill_1 FILLER_70_768 ();
 sg13g2_fill_2 FILLER_70_785 ();
 sg13g2_fill_1 FILLER_70_787 ();
 sg13g2_fill_1 FILLER_70_819 ();
 sg13g2_fill_1 FILLER_70_829 ();
 sg13g2_fill_2 FILLER_70_859 ();
 sg13g2_fill_1 FILLER_71_162 ();
 sg13g2_fill_2 FILLER_71_304 ();
 sg13g2_fill_1 FILLER_71_306 ();
 sg13g2_fill_2 FILLER_71_311 ();
 sg13g2_fill_1 FILLER_71_378 ();
 sg13g2_fill_2 FILLER_71_405 ();
 sg13g2_fill_1 FILLER_71_407 ();
 sg13g2_decap_4 FILLER_71_479 ();
 sg13g2_fill_2 FILLER_71_522 ();
 sg13g2_fill_2 FILLER_71_569 ();
 sg13g2_fill_1 FILLER_71_623 ();
 sg13g2_fill_2 FILLER_71_629 ();
 sg13g2_fill_1 FILLER_71_631 ();
 sg13g2_fill_1 FILLER_71_677 ();
 sg13g2_fill_2 FILLER_71_704 ();
 sg13g2_fill_2 FILLER_71_767 ();
 sg13g2_fill_1 FILLER_71_769 ();
 sg13g2_fill_2 FILLER_71_784 ();
 sg13g2_fill_1 FILLER_71_786 ();
 sg13g2_fill_2 FILLER_71_805 ();
 sg13g2_fill_1 FILLER_71_816 ();
 sg13g2_fill_1 FILLER_71_822 ();
 sg13g2_fill_2 FILLER_71_876 ();
 sg13g2_fill_2 FILLER_72_54 ();
 sg13g2_fill_1 FILLER_72_79 ();
 sg13g2_fill_1 FILLER_72_94 ();
 sg13g2_fill_2 FILLER_72_108 ();
 sg13g2_fill_1 FILLER_72_163 ();
 sg13g2_fill_1 FILLER_72_204 ();
 sg13g2_fill_1 FILLER_72_215 ();
 sg13g2_fill_1 FILLER_72_221 ();
 sg13g2_fill_1 FILLER_72_232 ();
 sg13g2_fill_1 FILLER_72_259 ();
 sg13g2_fill_1 FILLER_72_295 ();
 sg13g2_fill_2 FILLER_72_306 ();
 sg13g2_fill_1 FILLER_72_343 ();
 sg13g2_fill_1 FILLER_72_348 ();
 sg13g2_fill_1 FILLER_72_353 ();
 sg13g2_fill_1 FILLER_72_359 ();
 sg13g2_fill_1 FILLER_72_364 ();
 sg13g2_fill_1 FILLER_72_419 ();
 sg13g2_fill_1 FILLER_72_425 ();
 sg13g2_fill_1 FILLER_72_438 ();
 sg13g2_fill_1 FILLER_72_444 ();
 sg13g2_fill_1 FILLER_72_449 ();
 sg13g2_fill_2 FILLER_72_454 ();
 sg13g2_fill_2 FILLER_72_461 ();
 sg13g2_fill_1 FILLER_72_508 ();
 sg13g2_fill_1 FILLER_72_535 ();
 sg13g2_fill_1 FILLER_72_541 ();
 sg13g2_fill_2 FILLER_72_568 ();
 sg13g2_fill_2 FILLER_72_579 ();
 sg13g2_fill_1 FILLER_72_581 ();
 sg13g2_fill_1 FILLER_72_589 ();
 sg13g2_fill_2 FILLER_72_670 ();
 sg13g2_fill_1 FILLER_72_672 ();
 sg13g2_fill_1 FILLER_72_682 ();
 sg13g2_fill_2 FILLER_72_704 ();
 sg13g2_fill_1 FILLER_72_706 ();
 sg13g2_fill_2 FILLER_72_716 ();
 sg13g2_fill_1 FILLER_72_718 ();
 sg13g2_fill_1 FILLER_72_727 ();
 sg13g2_fill_1 FILLER_72_838 ();
 sg13g2_fill_1 FILLER_72_844 ();
 sg13g2_fill_1 FILLER_73_31 ();
 sg13g2_fill_1 FILLER_73_37 ();
 sg13g2_fill_1 FILLER_73_52 ();
 sg13g2_fill_1 FILLER_73_115 ();
 sg13g2_fill_2 FILLER_73_195 ();
 sg13g2_fill_1 FILLER_73_273 ();
 sg13g2_fill_2 FILLER_73_328 ();
 sg13g2_fill_1 FILLER_73_330 ();
 sg13g2_fill_1 FILLER_73_341 ();
 sg13g2_fill_1 FILLER_73_347 ();
 sg13g2_fill_2 FILLER_73_374 ();
 sg13g2_fill_1 FILLER_73_376 ();
 sg13g2_fill_2 FILLER_73_386 ();
 sg13g2_fill_2 FILLER_73_397 ();
 sg13g2_fill_1 FILLER_73_399 ();
 sg13g2_fill_2 FILLER_73_408 ();
 sg13g2_fill_2 FILLER_73_438 ();
 sg13g2_fill_1 FILLER_73_440 ();
 sg13g2_fill_1 FILLER_73_452 ();
 sg13g2_fill_1 FILLER_73_463 ();
 sg13g2_fill_1 FILLER_73_470 ();
 sg13g2_fill_1 FILLER_73_475 ();
 sg13g2_fill_1 FILLER_73_522 ();
 sg13g2_fill_1 FILLER_73_528 ();
 sg13g2_fill_1 FILLER_73_580 ();
 sg13g2_fill_1 FILLER_73_608 ();
 sg13g2_fill_1 FILLER_73_622 ();
 sg13g2_fill_2 FILLER_73_714 ();
 sg13g2_fill_1 FILLER_73_748 ();
 sg13g2_fill_2 FILLER_73_771 ();
 sg13g2_fill_1 FILLER_73_787 ();
 sg13g2_fill_1 FILLER_73_819 ();
 sg13g2_fill_1 FILLER_74_76 ();
 sg13g2_fill_1 FILLER_74_87 ();
 sg13g2_fill_1 FILLER_74_117 ();
 sg13g2_fill_2 FILLER_74_123 ();
 sg13g2_fill_2 FILLER_74_130 ();
 sg13g2_fill_2 FILLER_74_167 ();
 sg13g2_fill_1 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_216 ();
 sg13g2_fill_1 FILLER_74_253 ();
 sg13g2_fill_2 FILLER_74_305 ();
 sg13g2_fill_1 FILLER_74_376 ();
 sg13g2_fill_1 FILLER_74_382 ();
 sg13g2_fill_1 FILLER_74_409 ();
 sg13g2_fill_1 FILLER_74_414 ();
 sg13g2_fill_1 FILLER_74_441 ();
 sg13g2_fill_2 FILLER_74_478 ();
 sg13g2_fill_1 FILLER_74_480 ();
 sg13g2_fill_1 FILLER_74_488 ();
 sg13g2_fill_1 FILLER_74_494 ();
 sg13g2_fill_1 FILLER_74_499 ();
 sg13g2_fill_2 FILLER_74_578 ();
 sg13g2_fill_2 FILLER_74_620 ();
 sg13g2_fill_1 FILLER_74_622 ();
 sg13g2_fill_2 FILLER_74_660 ();
 sg13g2_fill_1 FILLER_74_662 ();
 sg13g2_fill_2 FILLER_74_672 ();
 sg13g2_fill_1 FILLER_74_684 ();
 sg13g2_fill_1 FILLER_74_700 ();
 sg13g2_fill_1 FILLER_74_711 ();
 sg13g2_fill_1 FILLER_74_782 ();
 sg13g2_fill_2 FILLER_74_801 ();
 sg13g2_fill_1 FILLER_74_808 ();
 sg13g2_fill_1 FILLER_74_814 ();
 sg13g2_fill_2 FILLER_74_820 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_fill_1 FILLER_75_44 ();
 sg13g2_fill_1 FILLER_75_65 ();
 sg13g2_fill_1 FILLER_75_81 ();
 sg13g2_fill_1 FILLER_75_92 ();
 sg13g2_fill_1 FILLER_75_98 ();
 sg13g2_fill_1 FILLER_75_104 ();
 sg13g2_fill_2 FILLER_75_110 ();
 sg13g2_fill_2 FILLER_75_121 ();
 sg13g2_fill_1 FILLER_75_251 ();
 sg13g2_fill_2 FILLER_75_257 ();
 sg13g2_fill_2 FILLER_75_319 ();
 sg13g2_fill_2 FILLER_75_329 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_fill_2 FILLER_75_353 ();
 sg13g2_fill_2 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_380 ();
 sg13g2_fill_2 FILLER_75_389 ();
 sg13g2_fill_1 FILLER_75_400 ();
 sg13g2_fill_1 FILLER_75_427 ();
 sg13g2_fill_1 FILLER_75_433 ();
 sg13g2_fill_1 FILLER_75_439 ();
 sg13g2_fill_2 FILLER_75_448 ();
 sg13g2_fill_1 FILLER_75_455 ();
 sg13g2_fill_1 FILLER_75_460 ();
 sg13g2_fill_1 FILLER_75_487 ();
 sg13g2_fill_1 FILLER_75_493 ();
 sg13g2_fill_1 FILLER_75_499 ();
 sg13g2_fill_1 FILLER_75_505 ();
 sg13g2_fill_2 FILLER_75_511 ();
 sg13g2_fill_2 FILLER_75_623 ();
 sg13g2_fill_1 FILLER_75_630 ();
 sg13g2_fill_1 FILLER_75_657 ();
 sg13g2_fill_1 FILLER_75_692 ();
 sg13g2_fill_1 FILLER_75_732 ();
 sg13g2_fill_2 FILLER_75_842 ();
 sg13g2_fill_1 FILLER_76_36 ();
 sg13g2_fill_1 FILLER_76_47 ();
 sg13g2_fill_1 FILLER_76_84 ();
 sg13g2_fill_1 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_143 ();
 sg13g2_fill_1 FILLER_76_149 ();
 sg13g2_fill_1 FILLER_76_159 ();
 sg13g2_fill_1 FILLER_76_199 ();
 sg13g2_fill_1 FILLER_76_226 ();
 sg13g2_fill_1 FILLER_76_305 ();
 sg13g2_fill_2 FILLER_76_314 ();
 sg13g2_fill_1 FILLER_76_404 ();
 sg13g2_fill_1 FILLER_76_413 ();
 sg13g2_fill_2 FILLER_76_418 ();
 sg13g2_fill_2 FILLER_76_485 ();
 sg13g2_fill_1 FILLER_76_487 ();
 sg13g2_fill_2 FILLER_76_605 ();
 sg13g2_fill_1 FILLER_76_607 ();
 sg13g2_fill_2 FILLER_76_790 ();
 sg13g2_fill_1 FILLER_76_827 ();
 sg13g2_fill_2 FILLER_76_833 ();
 sg13g2_fill_2 FILLER_76_875 ();
 sg13g2_fill_1 FILLER_76_877 ();
 sg13g2_fill_1 FILLER_77_56 ();
 sg13g2_fill_1 FILLER_77_78 ();
 sg13g2_fill_1 FILLER_77_89 ();
 sg13g2_fill_2 FILLER_77_129 ();
 sg13g2_fill_2 FILLER_77_135 ();
 sg13g2_fill_1 FILLER_77_146 ();
 sg13g2_fill_1 FILLER_77_173 ();
 sg13g2_fill_1 FILLER_77_255 ();
 sg13g2_fill_1 FILLER_77_299 ();
 sg13g2_fill_1 FILLER_77_326 ();
 sg13g2_fill_1 FILLER_77_337 ();
 sg13g2_fill_2 FILLER_77_348 ();
 sg13g2_fill_2 FILLER_77_380 ();
 sg13g2_fill_1 FILLER_77_433 ();
 sg13g2_fill_1 FILLER_77_597 ();
 sg13g2_fill_1 FILLER_77_639 ();
 sg13g2_fill_2 FILLER_77_651 ();
 sg13g2_fill_1 FILLER_77_851 ();
 sg13g2_fill_2 FILLER_77_856 ();
 sg13g2_decap_8 FILLER_77_862 ();
 sg13g2_fill_1 FILLER_77_869 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_27 ();
 sg13g2_fill_1 FILLER_78_64 ();
 sg13g2_fill_2 FILLER_78_105 ();
 sg13g2_fill_1 FILLER_78_351 ();
 sg13g2_fill_2 FILLER_78_369 ();
 sg13g2_fill_1 FILLER_78_371 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_fill_2 FILLER_78_413 ();
 sg13g2_fill_1 FILLER_78_446 ();
 sg13g2_fill_1 FILLER_78_451 ();
 sg13g2_fill_1 FILLER_78_460 ();
 sg13g2_fill_2 FILLER_78_495 ();
 sg13g2_fill_2 FILLER_78_523 ();
 sg13g2_fill_1 FILLER_78_564 ();
 sg13g2_fill_1 FILLER_78_623 ();
 sg13g2_fill_2 FILLER_78_731 ();
 sg13g2_fill_2 FILLER_78_737 ();
 sg13g2_fill_2 FILLER_78_747 ();
 sg13g2_fill_1 FILLER_78_782 ();
 sg13g2_fill_1 FILLER_78_788 ();
 sg13g2_decap_8 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_853 ();
 sg13g2_decap_8 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_78_867 ();
 sg13g2_fill_1 FILLER_79_110 ();
 sg13g2_fill_1 FILLER_79_121 ();
 sg13g2_fill_2 FILLER_79_169 ();
 sg13g2_fill_1 FILLER_79_379 ();
 sg13g2_fill_1 FILLER_79_426 ();
 sg13g2_fill_1 FILLER_79_437 ();
 sg13g2_fill_1 FILLER_79_474 ();
 sg13g2_fill_1 FILLER_79_485 ();
 sg13g2_fill_1 FILLER_79_512 ();
 sg13g2_fill_1 FILLER_79_681 ();
 sg13g2_fill_2 FILLER_79_711 ();
 sg13g2_fill_1 FILLER_79_750 ();
 sg13g2_fill_1 FILLER_79_756 ();
 sg13g2_fill_2 FILLER_79_794 ();
 sg13g2_decap_8 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_decap_8 FILLER_79_862 ();
 sg13g2_decap_8 FILLER_79_869 ();
 sg13g2_fill_2 FILLER_79_876 ();
 sg13g2_fill_2 FILLER_80_62 ();
 sg13g2_fill_1 FILLER_80_131 ();
 sg13g2_fill_1 FILLER_80_189 ();
 sg13g2_fill_1 FILLER_80_258 ();
 sg13g2_fill_1 FILLER_80_331 ();
 sg13g2_fill_2 FILLER_80_337 ();
 sg13g2_fill_1 FILLER_80_423 ();
 sg13g2_fill_1 FILLER_80_454 ();
 sg13g2_fill_2 FILLER_80_468 ();
 sg13g2_fill_1 FILLER_80_478 ();
 sg13g2_fill_1 FILLER_80_489 ();
 sg13g2_fill_1 FILLER_80_504 ();
 sg13g2_fill_1 FILLER_80_519 ();
 sg13g2_fill_2 FILLER_80_541 ();
 sg13g2_fill_1 FILLER_80_633 ();
 sg13g2_fill_1 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_838 ();
 sg13g2_decap_8 FILLER_80_845 ();
 sg13g2_decap_8 FILLER_80_852 ();
 sg13g2_decap_8 FILLER_80_859 ();
 sg13g2_decap_8 FILLER_80_866 ();
 sg13g2_decap_4 FILLER_80_873 ();
 sg13g2_fill_1 FILLER_80_877 ();
endmodule
