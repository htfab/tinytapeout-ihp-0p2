module tt_um_algofoogle_vga_fun_wrapper (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire clknet_0_clk;
 wire net86;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[1] ;
 wire \counter[20] ;
 wire \counter[21] ;
 wire \counter[22] ;
 wire \counter[23] ;
 wire \counter[24] ;
 wire \counter[25] ;
 wire \counter[26] ;
 wire \counter[27] ;
 wire \counter[28] ;
 wire \counter[29] ;
 wire \counter[2] ;
 wire \counter[30] ;
 wire \counter[31] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \depth[0] ;
 wire \depth[1] ;
 wire \depth[2] ;
 wire \dither_threshold[0] ;
 wire \dither_threshold[1] ;
 wire \dither_threshold[2] ;
 wire \dither_threshold[3] ;
 wire \dither_threshold[4] ;
 wire \frame_counter[0] ;
 wire \frame_counter[1] ;
 wire hsync;
 wire \i_project.controller_0.divider[0] ;
 wire \i_project.controller_0.divider[1] ;
 wire \i_project.controller_0.grey_pass[10] ;
 wire \i_project.controller_0.grey_pass[11] ;
 wire \i_project.controller_0.grey_pass[12] ;
 wire \i_project.controller_0.grey_pass[13] ;
 wire \i_project.controller_0.grey_pass[14] ;
 wire \i_project.controller_0.grey_pass[15] ;
 wire \i_project.controller_0.h[0] ;
 wire \i_project.controller_0.h[1] ;
 wire \i_project.controller_0.h[2] ;
 wire \i_project.controller_0.h[3] ;
 wire \i_project.controller_0.h[4] ;
 wire \i_project.controller_0.h[5] ;
 wire \i_project.controller_0.h[6] ;
 wire \i_project.controller_0.h[7] ;
 wire \i_project.controller_0.h[8] ;
 wire \i_project.controller_0.h[9] ;
 wire \i_project.controller_0.mode[0] ;
 wire \i_project.controller_0.mode[1] ;
 wire \i_project.controller_0.mode[2] ;
 wire \i_project.controller_0.mode_ramp_base[0] ;
 wire \i_project.controller_0.mode_ramp_base[1] ;
 wire \i_project.controller_0.mode_ramp_base[2] ;
 wire \i_project.controller_0.mode_ramp_base[3] ;
 wire \i_project.controller_0.mode_ramp_base[4] ;
 wire \i_project.controller_0.mode_ramp_base[5] ;
 wire \i_project.controller_0.mode_ramp_base[6] ;
 wire \i_project.controller_0.mode_ramp_base[7] ;
 wire \i_project.controller_0.rst_n ;
 wire \i_project.controller_0.t[10] ;
 wire \i_project.controller_0.t[11] ;
 wire \i_project.controller_0.t[8] ;
 wire \i_project.controller_0.t[9] ;
 wire \i_project.controller_0.v[0] ;
 wire \i_project.controller_0.v[1] ;
 wire \i_project.controller_0.v[2] ;
 wire \i_project.controller_0.v[3] ;
 wire \i_project.controller_0.v[4] ;
 wire \i_project.controller_0.v[5] ;
 wire \i_project.controller_0.v[6] ;
 wire \i_project.controller_0.v[7] ;
 wire \i_project.controller_0.v[8] ;
 wire \i_project.controller_0.v[9] ;
 wire \i_project.controller_0.vga_sync.hsync ;
 wire \i_project.controller_0.vga_sync.mode ;
 wire \i_project.controller_0.vga_sync.o_vsync ;
 wire \i_project.controller_0.vga_sync.vsync ;
 wire \i_project.controller_0.voffset[0] ;
 wire \i_project.controller_0.voffset[1] ;
 wire \i_project.controller_0.voffset[2] ;
 wire \i_project.controller_0.voffset[3] ;
 wire \i_project.controller_0.voffset[4] ;
 wire \i_project.controller_0.voffset[5] ;
 wire \i_project.controller_0.voffset[6] ;
 wire \i_project.controller_0.voffset[7] ;
 wire prev_vsync;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_nor2b_1 _2123_ (.A(_0479_),
    .B_N(_0481_),
    .Y(_0482_));
 sg13g2_a21oi_1 _2124_ (.A1(_1982_),
    .A2(net41),
    .Y(_0483_),
    .B1(net30));
 sg13g2_o21ai_1 _2125_ (.B1(_0483_),
    .Y(_0484_),
    .A1(_0468_),
    .A2(_0482_));
 sg13g2_a21oi_1 _2126_ (.A1(_0220_),
    .A2(_0484_),
    .Y(_0485_),
    .B1(net56));
 sg13g2_a221oi_1 _2127_ (.B2(_0251_),
    .C1(_0299_),
    .B1(_0420_),
    .A1(_0052_),
    .Y(_0486_),
    .A2(net56));
 sg13g2_nand2b_1 _2128_ (.Y(_0487_),
    .B(_0486_),
    .A_N(_0485_));
 sg13g2_nand2_1 _2129_ (.Y(_0488_),
    .A(_0449_),
    .B(_0487_));
 sg13g2_a21oi_1 _2130_ (.A1(_0228_),
    .A2(net23),
    .Y(_0489_),
    .B1(_0488_));
 sg13g2_nand2_1 _2131_ (.Y(_0490_),
    .A(net22),
    .B(_0343_));
 sg13g2_nand3_1 _2132_ (.B(_0489_),
    .C(_0490_),
    .A(_0466_),
    .Y(_0491_));
 sg13g2_nor2_1 _2133_ (.A(net54),
    .B(_0243_),
    .Y(_0492_));
 sg13g2_inv_1 _2134_ (.Y(_0493_),
    .A(_0492_));
 sg13g2_inv_1 _2135_ (.Y(_0494_),
    .A(_0238_));
 sg13g2_o21ai_1 _2136_ (.B1(_0494_),
    .Y(_0495_),
    .A1(_0242_),
    .A2(_0493_));
 sg13g2_nand2_1 _2137_ (.Y(_0496_),
    .A(_0466_),
    .B(_0495_));
 sg13g2_nand2_2 _2138_ (.Y(_0497_),
    .A(_0496_),
    .B(_0455_));
 sg13g2_nor2_1 _2139_ (.A(_0491_),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_nor2_1 _2140_ (.A(_0465_),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_nand2_1 _2141_ (.Y(_0500_),
    .A(_0464_),
    .B(_0499_));
 sg13g2_inv_4 _2142_ (.A(_0497_),
    .Y(_0501_));
 sg13g2_nand2_2 _2143_ (.Y(_0502_),
    .A(_0491_),
    .B(_0455_));
 sg13g2_nor2_1 _2144_ (.A(_0501_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_xnor2_1 _2145_ (.Y(_0504_),
    .A(_1540_),
    .B(net33));
 sg13g2_a21oi_1 _2146_ (.A1(_0504_),
    .A2(net53),
    .Y(_0505_),
    .B1(net47));
 sg13g2_nor2_1 _2147_ (.A(_1504_),
    .B(_0357_),
    .Y(_0506_));
 sg13g2_a21oi_2 _2148_ (.B1(_0506_),
    .Y(_0507_),
    .A2(_0429_),
    .A1(_1504_));
 sg13g2_nand2_1 _2149_ (.Y(_0508_),
    .A(_0507_),
    .B(net48));
 sg13g2_xnor2_1 _2150_ (.Y(_0509_),
    .A(_2018_),
    .B(_0267_));
 sg13g2_xnor2_1 _2151_ (.Y(_0510_),
    .A(_1979_),
    .B(_0261_));
 sg13g2_xnor2_1 _2152_ (.Y(_0511_),
    .A(_0509_),
    .B(_0510_));
 sg13g2_a22oi_1 _2153_ (.Y(_0512_),
    .B1(net40),
    .B2(_0511_),
    .A2(_0508_),
    .A1(_0505_));
 sg13g2_o21ai_1 _2154_ (.B1(_0323_),
    .Y(_0513_),
    .A1(_0024_),
    .A2(net33));
 sg13g2_o21ai_1 _2155_ (.B1(_0513_),
    .Y(_0514_),
    .A1(net49),
    .A2(_0512_));
 sg13g2_nand2_1 _2156_ (.Y(_0515_),
    .A(_0514_),
    .B(net36));
 sg13g2_a21oi_1 _2157_ (.A1(net25),
    .A2(net33),
    .Y(_0516_),
    .B1(_0327_));
 sg13g2_o21ai_1 _2158_ (.B1(_0516_),
    .Y(_0517_),
    .A1(_1978_),
    .A2(_0397_));
 sg13g2_nand3_1 _2159_ (.B(net42),
    .C(_0517_),
    .A(_0515_),
    .Y(_0518_));
 sg13g2_a21oi_1 _2160_ (.A1(_1985_),
    .A2(net35),
    .Y(_0519_),
    .B1(net30));
 sg13g2_a21oi_1 _2161_ (.A1(_0518_),
    .A2(_0519_),
    .Y(_0520_),
    .B1(_0221_));
 sg13g2_inv_1 _2162_ (.Y(_0521_),
    .A(_0243_));
 sg13g2_nor2_1 _2163_ (.A(_0521_),
    .B(_0299_),
    .Y(_0522_));
 sg13g2_inv_1 _2164_ (.Y(_0523_),
    .A(_0522_));
 sg13g2_a21oi_1 _2165_ (.A1(_0051_),
    .A2(_1624_),
    .Y(_0524_),
    .B1(_0523_));
 sg13g2_o21ai_1 _2166_ (.B1(_0524_),
    .Y(_0525_),
    .A1(net56),
    .A2(_0520_));
 sg13g2_nor2b_1 _2167_ (.A(_0248_),
    .B_N(_0525_),
    .Y(_0526_));
 sg13g2_inv_1 _2168_ (.Y(_0527_),
    .A(net51));
 sg13g2_nand2_1 _2169_ (.Y(_0528_),
    .A(_0408_),
    .B(_0527_));
 sg13g2_nand2_1 _2170_ (.Y(_0529_),
    .A(net22),
    .B(_0528_));
 sg13g2_nand2_1 _2171_ (.Y(_0530_),
    .A(_0526_),
    .B(_0529_));
 sg13g2_nand2_1 _2172_ (.Y(_0531_),
    .A(_0530_),
    .B(_0455_));
 sg13g2_nor2_1 _2173_ (.A(net22),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_nor2_1 _2174_ (.A(_0503_),
    .B(_0532_),
    .Y(_0533_));
 sg13g2_nand2_2 _2175_ (.Y(_0534_),
    .A(_0500_),
    .B(_0533_));
 sg13g2_nand3_1 _2176_ (.B(net22),
    .C(_0529_),
    .A(_0526_),
    .Y(_0535_));
 sg13g2_buf_2 _2177_ (.A(_0535_),
    .X(_0536_));
 sg13g2_nand2_2 _2178_ (.Y(_0537_),
    .A(_0534_),
    .B(_0536_));
 sg13g2_nand2_1 _2179_ (.Y(_0538_),
    .A(_0537_),
    .B(_0463_));
 sg13g2_inv_1 _2180_ (.Y(_0539_),
    .A(_0463_));
 sg13g2_nand3_1 _2181_ (.B(_0539_),
    .C(_0536_),
    .A(_0534_),
    .Y(_0540_));
 sg13g2_nand2_1 _2182_ (.Y(_0541_),
    .A(_0538_),
    .B(_0540_));
 sg13g2_nor2_2 _2183_ (.A(_0454_),
    .B(_0453_),
    .Y(_0542_));
 sg13g2_nor2_1 _2184_ (.A(_0542_),
    .B(_0463_),
    .Y(_0543_));
 sg13g2_xnor2_1 _2185_ (.Y(_0544_),
    .A(_0501_),
    .B(_0543_));
 sg13g2_nand2_1 _2186_ (.Y(_0545_),
    .A(_0537_),
    .B(_0544_));
 sg13g2_nand3_1 _2187_ (.B(_0536_),
    .C(_0497_),
    .A(_0534_),
    .Y(_0546_));
 sg13g2_nand2_2 _2188_ (.Y(_0547_),
    .A(_0545_),
    .B(_0546_));
 sg13g2_inv_4 _2189_ (.A(_0547_),
    .Y(_0548_));
 sg13g2_nor2_1 _2190_ (.A(_0502_),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_xnor2_1 _2191_ (.Y(_0550_),
    .A(_0542_),
    .B(_0463_));
 sg13g2_nand2_1 _2192_ (.Y(_0551_),
    .A(_0537_),
    .B(_0550_));
 sg13g2_nand3_1 _2193_ (.B(_0536_),
    .C(_0542_),
    .A(_0534_),
    .Y(_0552_));
 sg13g2_nand2_2 _2194_ (.Y(_0553_),
    .A(_0551_),
    .B(_0552_));
 sg13g2_nand2_1 _2195_ (.Y(_0554_),
    .A(_0448_),
    .B(_0455_));
 sg13g2_nand2_1 _2196_ (.Y(_0555_),
    .A(_0553_),
    .B(_0554_));
 sg13g2_nor2_1 _2197_ (.A(_0454_),
    .B(_0413_),
    .Y(_0556_));
 sg13g2_inv_1 _2198_ (.Y(_0557_),
    .A(_0556_));
 sg13g2_nand3_1 _2199_ (.B(_0540_),
    .C(_0557_),
    .A(_0538_),
    .Y(_0558_));
 sg13g2_buf_2 _2200_ (.A(_0558_),
    .X(_0559_));
 sg13g2_nor2_1 _2201_ (.A(_0554_),
    .B(_0553_),
    .Y(_0560_));
 sg13g2_a21oi_1 _2202_ (.A1(_0555_),
    .A2(_0559_),
    .Y(_0561_),
    .B1(_0560_));
 sg13g2_nand2b_1 _2203_ (.Y(_0562_),
    .B(_0561_),
    .A_N(_0549_));
 sg13g2_nand2_1 _2204_ (.Y(_0563_),
    .A(_0548_),
    .B(_0502_));
 sg13g2_nor3_1 _2205_ (.A(_0542_),
    .B(_0463_),
    .C(_0501_),
    .Y(_0564_));
 sg13g2_xnor2_1 _2206_ (.Y(_0565_),
    .A(net22),
    .B(_0564_));
 sg13g2_nand2_1 _2207_ (.Y(_0566_),
    .A(_0537_),
    .B(_0565_));
 sg13g2_nand3_1 _2208_ (.B(_0459_),
    .C(_0536_),
    .A(_0534_),
    .Y(_0567_));
 sg13g2_nand2_1 _2209_ (.Y(_0568_),
    .A(_0566_),
    .B(_0567_));
 sg13g2_nor2_1 _2210_ (.A(_0459_),
    .B(_0531_),
    .Y(_0569_));
 sg13g2_a21oi_2 _2211_ (.B1(_0569_),
    .Y(_0570_),
    .A2(_0531_),
    .A1(_0568_));
 sg13g2_nand3_1 _2212_ (.B(_0563_),
    .C(_0570_),
    .A(_0562_),
    .Y(_0571_));
 sg13g2_xnor2_1 _2213_ (.Y(_0572_),
    .A(_0502_),
    .B(_0547_));
 sg13g2_nand2b_1 _2214_ (.Y(_0573_),
    .B(_0553_),
    .A_N(_0554_));
 sg13g2_nand3_1 _2215_ (.B(_0552_),
    .C(_0554_),
    .A(_0551_),
    .Y(_0574_));
 sg13g2_nand2_1 _2216_ (.Y(_0575_),
    .A(_0573_),
    .B(_0574_));
 sg13g2_nand3_1 _2217_ (.B(_0575_),
    .C(_0559_),
    .A(_0572_),
    .Y(_0576_));
 sg13g2_a21oi_1 _2218_ (.A1(_0563_),
    .A2(_0560_),
    .Y(_0577_),
    .B1(_0549_));
 sg13g2_inv_1 _2219_ (.Y(_0578_),
    .A(_0570_));
 sg13g2_nand3_1 _2220_ (.B(_0577_),
    .C(_0578_),
    .A(_0576_),
    .Y(_0579_));
 sg13g2_nand2_1 _2221_ (.Y(_0580_),
    .A(_0571_),
    .B(_0579_));
 sg13g2_inv_2 _2222_ (.Y(_0581_),
    .A(_1698_));
 sg13g2_nand2_1 _2223_ (.Y(_0582_),
    .A(_0580_),
    .B(_0581_));
 sg13g2_nand3_1 _2224_ (.B(_0579_),
    .C(_1698_),
    .A(_0571_),
    .Y(_0583_));
 sg13g2_nand2_1 _2225_ (.Y(_0584_),
    .A(_0582_),
    .B(_0583_));
 sg13g2_inv_1 _2226_ (.Y(_0585_),
    .A(_0561_));
 sg13g2_xor2_1 _2227_ (.B(_0547_),
    .A(_0502_),
    .X(_0586_));
 sg13g2_nor2_1 _2228_ (.A(_0570_),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_nand2_1 _2229_ (.Y(_0588_),
    .A(_0585_),
    .B(_0587_));
 sg13g2_a21oi_1 _2230_ (.A1(_0503_),
    .A2(_0536_),
    .Y(_0589_),
    .B1(_0532_));
 sg13g2_nand2_1 _2231_ (.Y(_0590_),
    .A(_0588_),
    .B(_0589_));
 sg13g2_nand2_1 _2232_ (.Y(_0591_),
    .A(_0590_),
    .B(_0537_));
 sg13g2_nand2_1 _2233_ (.Y(_0592_),
    .A(_0591_),
    .B(_1670_));
 sg13g2_nand3_1 _2234_ (.B(_1706_),
    .C(_0537_),
    .A(_0590_),
    .Y(_0593_));
 sg13g2_nand2_1 _2235_ (.Y(_0594_),
    .A(_0592_),
    .B(_0593_));
 sg13g2_xnor2_1 _2236_ (.Y(_0595_),
    .A(_0559_),
    .B(_0575_));
 sg13g2_xnor2_1 _2237_ (.Y(_0596_),
    .A(_1661_),
    .B(_0595_));
 sg13g2_xnor2_1 _2238_ (.Y(_0597_),
    .A(_0572_),
    .B(_0561_));
 sg13g2_xnor2_1 _2239_ (.Y(_0598_),
    .A(_1664_),
    .B(_0597_));
 sg13g2_nor2_1 _2240_ (.A(_0596_),
    .B(_0598_),
    .Y(_0599_));
 sg13g2_nand3_1 _2241_ (.B(_0594_),
    .C(_0599_),
    .A(_0584_),
    .Y(_0600_));
 sg13g2_inv_1 _2242_ (.Y(_0601_),
    .A(_0559_));
 sg13g2_inv_2 _2243_ (.Y(_0602_),
    .A(_0541_));
 sg13g2_nor2_1 _2244_ (.A(_0557_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_o21ai_1 _2245_ (.B1(_0029_),
    .Y(_0604_),
    .A1(_0601_),
    .A2(_0603_));
 sg13g2_nor2b_1 _2246_ (.A(_0600_),
    .B_N(_0604_),
    .Y(_0605_));
 sg13g2_xnor2_1 _2247_ (.Y(_0606_),
    .A(_1706_),
    .B(_0591_));
 sg13g2_nand3_1 _2248_ (.B(_0579_),
    .C(_0581_),
    .A(_0571_),
    .Y(_0607_));
 sg13g2_nand3_1 _2249_ (.B(_0563_),
    .C(_0578_),
    .A(_0562_),
    .Y(_0608_));
 sg13g2_nand3_1 _2250_ (.B(_0577_),
    .C(_0570_),
    .A(_0576_),
    .Y(_0609_));
 sg13g2_nand3_1 _2251_ (.B(_0609_),
    .C(_1698_),
    .A(_0608_),
    .Y(_0610_));
 sg13g2_nand2_1 _2252_ (.Y(_0611_),
    .A(_0607_),
    .B(_0610_));
 sg13g2_nor2_1 _2253_ (.A(_0606_),
    .B(_0611_),
    .Y(_0612_));
 sg13g2_nand2_1 _2254_ (.Y(_0613_),
    .A(_0595_),
    .B(_1661_));
 sg13g2_nand2b_1 _2255_ (.Y(_0614_),
    .B(_1658_),
    .A_N(_0597_));
 sg13g2_o21ai_1 _2256_ (.B1(_0614_),
    .Y(_0615_),
    .A1(_0613_),
    .A2(_0598_));
 sg13g2_nand2_1 _2257_ (.Y(_0616_),
    .A(_0612_),
    .B(_0615_));
 sg13g2_nor2_1 _2258_ (.A(_1694_),
    .B(_0580_),
    .Y(_0617_));
 sg13g2_a22oi_1 _2259_ (.Y(_0618_),
    .B1(_0617_),
    .B2(_0594_),
    .A2(_0591_),
    .A1(\dither_threshold[4] ));
 sg13g2_nand2_1 _2260_ (.Y(_0619_),
    .A(_0616_),
    .B(_0618_));
 sg13g2_nor2_2 _2261_ (.A(_0605_),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_xnor2_1 _2262_ (.Y(net8),
    .A(_0541_),
    .B(_0620_));
 sg13g2_a21oi_1 _2263_ (.A1(_0620_),
    .A2(_0602_),
    .Y(_0621_),
    .B1(_0553_));
 sg13g2_nand3_1 _2264_ (.B(_0602_),
    .C(_0553_),
    .A(_0620_),
    .Y(_0622_));
 sg13g2_nor2b_1 _2265_ (.A(_0621_),
    .B_N(_0622_),
    .Y(net9));
 sg13g2_nand2_1 _2266_ (.Y(_0623_),
    .A(_0622_),
    .B(_0548_));
 sg13g2_nand4_1 _2267_ (.B(_0602_),
    .C(_0547_),
    .A(_0620_),
    .Y(_0624_),
    .D(_0553_));
 sg13g2_nand2_1 _2268_ (.Y(net10),
    .A(_0623_),
    .B(_0624_));
 sg13g2_a21oi_1 _2269_ (.A1(_0551_),
    .A2(_0552_),
    .Y(_0625_),
    .B1(_0547_));
 sg13g2_nand3_1 _2270_ (.B(_0602_),
    .C(_0625_),
    .A(_0620_),
    .Y(_0626_));
 sg13g2_inv_1 _2271_ (.Y(_0627_),
    .A(_0568_));
 sg13g2_nand2_1 _2272_ (.Y(_0628_),
    .A(_0626_),
    .B(_0627_));
 sg13g2_nand4_1 _2273_ (.B(_0602_),
    .C(_0568_),
    .A(_0620_),
    .Y(_0629_),
    .D(_0625_));
 sg13g2_nand2_1 _2274_ (.Y(net11),
    .A(_0628_),
    .B(_0629_));
 sg13g2_xnor2_1 _2275_ (.Y(_0630_),
    .A(_1867_),
    .B(_0199_));
 sg13g2_nand2_1 _2276_ (.Y(_0631_),
    .A(net34),
    .B(_0039_));
 sg13g2_nor2_1 _2277_ (.A(_1994_),
    .B(_1916_),
    .Y(_0632_));
 sg13g2_nor2_1 _2278_ (.A(_0039_),
    .B(net34),
    .Y(_0633_));
 sg13g2_a21oi_1 _2279_ (.A1(_0631_),
    .A2(_0632_),
    .Y(_0634_),
    .B1(_0633_));
 sg13g2_xnor2_1 _2280_ (.Y(_0635_),
    .A(_1840_),
    .B(net32));
 sg13g2_nand2b_1 _2281_ (.Y(_0636_),
    .B(net26),
    .A_N(_0037_));
 sg13g2_nand3_1 _2282_ (.B(_0212_),
    .C(_0037_),
    .A(_0211_),
    .Y(_0637_));
 sg13g2_nand2_1 _2283_ (.Y(_0638_),
    .A(_0636_),
    .B(_0637_));
 sg13g2_nand2b_1 _2284_ (.Y(_0639_),
    .B(_0638_),
    .A_N(_0635_));
 sg13g2_nor2_1 _2285_ (.A(_0634_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_nor2_1 _2286_ (.A(_0037_),
    .B(net26),
    .Y(_0641_));
 sg13g2_inv_1 _2287_ (.Y(_0642_),
    .A(_0038_));
 sg13g2_nand2_1 _2288_ (.Y(_0643_),
    .A(_0146_),
    .B(_0642_));
 sg13g2_a21oi_1 _2289_ (.A1(_0037_),
    .A2(net26),
    .Y(_0644_),
    .B1(_0643_));
 sg13g2_nor2_1 _2290_ (.A(_0641_),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_nor2b_1 _2291_ (.A(_0640_),
    .B_N(_0645_),
    .Y(_0646_));
 sg13g2_xnor2_1 _2292_ (.Y(_0647_),
    .A(_1994_),
    .B(_1909_));
 sg13g2_inv_2 _2293_ (.Y(_0648_),
    .A(_0647_));
 sg13g2_xnor2_1 _2294_ (.Y(_0649_),
    .A(_1861_),
    .B(_1935_));
 sg13g2_nor2_1 _2295_ (.A(_0648_),
    .B(_0649_),
    .Y(_0650_));
 sg13g2_nor2b_1 _2296_ (.A(_0639_),
    .B_N(_0650_),
    .Y(_0651_));
 sg13g2_nor2_1 _2297_ (.A(_1936_),
    .B(net33),
    .Y(_0652_));
 sg13g2_xnor2_1 _2298_ (.Y(_0653_),
    .A(net73),
    .B(net38));
 sg13g2_nand2_1 _2299_ (.Y(_0654_),
    .A(_1958_),
    .B(_0043_));
 sg13g2_nor2_1 _2300_ (.A(_1844_),
    .B(_1963_),
    .Y(_0655_));
 sg13g2_nor2_1 _2301_ (.A(_0043_),
    .B(_1958_),
    .Y(_0656_));
 sg13g2_a21oi_1 _2302_ (.A1(_0654_),
    .A2(_0655_),
    .Y(_0657_),
    .B1(_0656_));
 sg13g2_inv_1 _2303_ (.Y(_0658_),
    .A(_0657_));
 sg13g2_nand2_1 _2304_ (.Y(_0659_),
    .A(_0653_),
    .B(_0658_));
 sg13g2_nand2_1 _2305_ (.Y(_0660_),
    .A(_1982_),
    .B(_1911_));
 sg13g2_nand2_1 _2306_ (.Y(_0661_),
    .A(_0659_),
    .B(_0660_));
 sg13g2_xnor2_1 _2307_ (.Y(_0662_),
    .A(net60),
    .B(_1977_));
 sg13g2_nand2_1 _2308_ (.Y(_0663_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_nand2b_2 _2309_ (.Y(_0664_),
    .B(_0663_),
    .A_N(_0652_));
 sg13g2_nand2_1 _2310_ (.Y(_0665_),
    .A(_0651_),
    .B(_0664_));
 sg13g2_nand2_1 _2311_ (.Y(_0666_),
    .A(_0646_),
    .B(_0665_));
 sg13g2_nand2b_1 _2312_ (.Y(_0667_),
    .B(_0666_),
    .A_N(_0630_));
 sg13g2_nand3_1 _2313_ (.B(_0665_),
    .C(_0630_),
    .A(_0646_),
    .Y(_0668_));
 sg13g2_nand2_1 _2314_ (.Y(_0669_),
    .A(_0667_),
    .B(_0668_));
 sg13g2_xor2_1 _2315_ (.B(\i_project.controller_0.t[11] ),
    .A(_1529_),
    .X(_0670_));
 sg13g2_nand2_1 _2316_ (.Y(_0671_),
    .A(net68),
    .B(_1841_));
 sg13g2_xnor2_1 _2317_ (.Y(_0672_),
    .A(net65),
    .B(_1856_));
 sg13g2_nand2_1 _2318_ (.Y(_0673_),
    .A(net65),
    .B(net60));
 sg13g2_o21ai_1 _2319_ (.B1(_0673_),
    .Y(_0674_),
    .A1(_0671_),
    .A2(_0672_));
 sg13g2_xor2_1 _2320_ (.B(_1861_),
    .A(_1526_),
    .X(_0675_));
 sg13g2_inv_1 _2321_ (.Y(_0676_),
    .A(_0675_));
 sg13g2_xor2_1 _2322_ (.B(net70),
    .A(net67),
    .X(_0677_));
 sg13g2_nor2b_1 _2323_ (.A(_0676_),
    .B_N(_0677_),
    .Y(_0678_));
 sg13g2_nand2_1 _2324_ (.Y(_0679_),
    .A(net67),
    .B(net70));
 sg13g2_nand2_1 _2325_ (.Y(_0680_),
    .A(net64),
    .B(_1861_));
 sg13g2_o21ai_1 _2326_ (.B1(_0680_),
    .Y(_0681_),
    .A1(_0679_),
    .A2(_0676_));
 sg13g2_a21oi_1 _2327_ (.A1(_0674_),
    .A2(_0678_),
    .Y(_0682_),
    .B1(_0681_));
 sg13g2_nand2_1 _2328_ (.Y(_0683_),
    .A(net80),
    .B(net72));
 sg13g2_xnor2_1 _2329_ (.Y(_0684_),
    .A(\i_project.controller_0.h[1] ),
    .B(_1852_));
 sg13g2_nand2_1 _2330_ (.Y(_0685_),
    .A(net79),
    .B(net61));
 sg13g2_o21ai_1 _2331_ (.B1(_0685_),
    .Y(_0686_),
    .A1(_0683_),
    .A2(_0684_));
 sg13g2_buf_1 _2332_ (.A(_0686_),
    .X(_0687_));
 sg13g2_xor2_1 _2333_ (.B(\i_project.controller_0.mode_ramp_base[5] ),
    .A(_1520_),
    .X(_0688_));
 sg13g2_inv_1 _2334_ (.Y(_0689_),
    .A(_0688_));
 sg13g2_nor2_1 _2335_ (.A(_0672_),
    .B(_0689_),
    .Y(_0690_));
 sg13g2_nand3_1 _2336_ (.B(_0690_),
    .C(_0678_),
    .A(_0687_),
    .Y(_0691_));
 sg13g2_nand2_1 _2337_ (.Y(_0692_),
    .A(_0682_),
    .B(_0691_));
 sg13g2_xor2_1 _2338_ (.B(_1839_),
    .A(_1532_),
    .X(_0693_));
 sg13g2_nand2_1 _2339_ (.Y(_0694_),
    .A(_0692_),
    .B(_0693_));
 sg13g2_nand2_1 _2340_ (.Y(_0695_),
    .A(net66),
    .B(_1839_));
 sg13g2_nand2_1 _2341_ (.Y(_0696_),
    .A(_0694_),
    .B(_0695_));
 sg13g2_inv_1 _2342_ (.Y(_0697_),
    .A(_0696_));
 sg13g2_nand2_1 _2343_ (.Y(_0698_),
    .A(net78),
    .B(\i_project.controller_0.t[10] ));
 sg13g2_nor2_1 _2344_ (.A(net78),
    .B(\i_project.controller_0.t[10] ),
    .Y(_0699_));
 sg13g2_a21oi_1 _2345_ (.A1(_0697_),
    .A2(_0698_),
    .Y(_0700_),
    .B1(_0699_));
 sg13g2_xnor2_1 _2346_ (.Y(_0701_),
    .A(_0670_),
    .B(_0700_));
 sg13g2_nand2_1 _2347_ (.Y(_0702_),
    .A(_0669_),
    .B(_0701_));
 sg13g2_inv_1 _2348_ (.Y(_0703_),
    .A(_0701_));
 sg13g2_nand3_1 _2349_ (.B(_0668_),
    .C(_0703_),
    .A(_0667_),
    .Y(_0704_));
 sg13g2_nand3_1 _2350_ (.B(_0704_),
    .C(_0315_),
    .A(_0702_),
    .Y(_0705_));
 sg13g2_a21oi_1 _2351_ (.A1(_0199_),
    .A2(_1530_),
    .Y(_0706_),
    .B1(net48));
 sg13g2_o21ai_1 _2352_ (.B1(_0706_),
    .Y(_0707_),
    .A1(_1530_),
    .A2(_0199_));
 sg13g2_a21oi_1 _2353_ (.A1(_0284_),
    .A2(net57),
    .Y(_0708_),
    .B1(net52));
 sg13g2_nand3_1 _2354_ (.B(_0707_),
    .C(_0708_),
    .A(_0705_),
    .Y(_0709_));
 sg13g2_xnor2_1 _2355_ (.Y(_0710_),
    .A(_0283_),
    .B(_0167_));
 sg13g2_a21oi_1 _2356_ (.A1(_0710_),
    .A2(net45),
    .Y(_0711_),
    .B1(net46));
 sg13g2_nand2_1 _2357_ (.Y(_0712_),
    .A(_0709_),
    .B(_0711_));
 sg13g2_a21oi_1 _2358_ (.A1(_0283_),
    .A2(net46),
    .Y(_0713_),
    .B1(net37));
 sg13g2_nand2_1 _2359_ (.Y(_0714_),
    .A(_0712_),
    .B(_0713_));
 sg13g2_nand2_1 _2360_ (.Y(_0715_),
    .A(_0714_),
    .B(_0220_));
 sg13g2_a21oi_1 _2361_ (.A1(_0715_),
    .A2(_0225_),
    .Y(_0716_),
    .B1(_0301_));
 sg13g2_buf_2 _2362_ (.A(_0716_),
    .X(_0717_));
 sg13g2_nand2_1 _2363_ (.Y(_0718_),
    .A(_0717_),
    .B(net51));
 sg13g2_nand2_1 _2364_ (.Y(_0719_),
    .A(_0717_),
    .B(_0245_));
 sg13g2_xor2_1 _2365_ (.B(_0692_),
    .A(_0693_),
    .X(_0720_));
 sg13g2_xnor2_1 _2366_ (.Y(_0721_),
    .A(_0038_),
    .B(net32));
 sg13g2_xnor2_1 _2367_ (.Y(_0722_),
    .A(_0720_),
    .B(_0721_));
 sg13g2_nand3b_1 _2368_ (.B(_0664_),
    .C(_0647_),
    .Y(_0723_),
    .A_N(_0649_));
 sg13g2_nand2_1 _2369_ (.Y(_0724_),
    .A(_0723_),
    .B(_0634_));
 sg13g2_nand2b_1 _2370_ (.Y(_0725_),
    .B(_0724_),
    .A_N(_0722_));
 sg13g2_nand3_1 _2371_ (.B(_0722_),
    .C(_0634_),
    .A(_0723_),
    .Y(_0726_));
 sg13g2_nand3_1 _2372_ (.B(_0726_),
    .C(_0315_),
    .A(_0725_),
    .Y(_0727_));
 sg13g2_nand2_1 _2373_ (.Y(_0728_),
    .A(_0727_),
    .B(_2054_));
 sg13g2_a21oi_1 _2374_ (.A1(_0354_),
    .A2(net57),
    .Y(_0729_),
    .B1(net52));
 sg13g2_nand2_1 _2375_ (.Y(_0730_),
    .A(_0728_),
    .B(_0729_));
 sg13g2_nor2b_1 _2376_ (.A(_0167_),
    .B_N(_0359_),
    .Y(_0731_));
 sg13g2_nor2_1 _2377_ (.A(_0359_),
    .B(_0168_),
    .Y(_0732_));
 sg13g2_nor3_1 _2378_ (.A(_0326_),
    .B(_0731_),
    .C(_0732_),
    .Y(_0733_));
 sg13g2_nor2_1 _2379_ (.A(_0333_),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_nand2_1 _2380_ (.Y(_0735_),
    .A(_0730_),
    .B(_0734_));
 sg13g2_a21oi_1 _2381_ (.A1(_0359_),
    .A2(_0333_),
    .Y(_0736_),
    .B1(net37));
 sg13g2_nand2_1 _2382_ (.Y(_0737_),
    .A(_0735_),
    .B(_0736_));
 sg13g2_nand2_1 _2383_ (.Y(_0738_),
    .A(_0737_),
    .B(_0223_));
 sg13g2_nand2_1 _2384_ (.Y(_0739_),
    .A(_0738_),
    .B(_0374_));
 sg13g2_nand2_1 _2385_ (.Y(_0740_),
    .A(_0739_),
    .B(_0237_));
 sg13g2_a21oi_1 _2386_ (.A1(_1889_),
    .A2(_0408_),
    .Y(_0741_),
    .B1(_0740_));
 sg13g2_a21oi_1 _2387_ (.A1(_0522_),
    .A2(_0739_),
    .Y(_0742_),
    .B1(_0741_));
 sg13g2_nand3_1 _2388_ (.B(_0719_),
    .C(_0742_),
    .A(_0718_),
    .Y(_0743_));
 sg13g2_buf_2 _2389_ (.A(_0743_),
    .X(_0744_));
 sg13g2_inv_2 _2390_ (.Y(_0745_),
    .A(_0744_));
 sg13g2_nand2_1 _2391_ (.Y(_0746_),
    .A(_0717_),
    .B(_1888_));
 sg13g2_o21ai_1 _2392_ (.B1(net43),
    .Y(_0747_),
    .A1(_0310_),
    .A2(_0379_));
 sg13g2_inv_1 _2393_ (.Y(_0748_),
    .A(_0633_));
 sg13g2_nand2_1 _2394_ (.Y(_0749_),
    .A(_0748_),
    .B(_0631_));
 sg13g2_a21o_1 _2395_ (.A2(_0690_),
    .A1(_0687_),
    .B1(_0674_),
    .X(_0750_));
 sg13g2_nand2_1 _2396_ (.Y(_0751_),
    .A(_0750_),
    .B(_0677_));
 sg13g2_nand2_1 _2397_ (.Y(_0752_),
    .A(_0751_),
    .B(_0679_));
 sg13g2_xnor2_1 _2398_ (.Y(_0753_),
    .A(_0675_),
    .B(_0752_));
 sg13g2_xnor2_1 _2399_ (.Y(_0754_),
    .A(_0749_),
    .B(_0753_));
 sg13g2_a21oi_1 _2400_ (.A1(_0664_),
    .A2(_0647_),
    .Y(_0755_),
    .B1(_0632_));
 sg13g2_xnor2_1 _2401_ (.Y(_0756_),
    .A(_0754_),
    .B(_0755_));
 sg13g2_a21oi_1 _2402_ (.A1(_0756_),
    .A2(_0388_),
    .Y(_0757_),
    .B1(_0355_));
 sg13g2_nor2b_1 _2403_ (.A(net29),
    .B_N(_0386_),
    .Y(_0758_));
 sg13g2_nor2_1 _2404_ (.A(_0386_),
    .B(_0169_),
    .Y(_0759_));
 sg13g2_nor3_1 _2405_ (.A(net43),
    .B(_0758_),
    .C(_0759_),
    .Y(_0760_));
 sg13g2_nor2_1 _2406_ (.A(net46),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_o21ai_1 _2407_ (.B1(_0761_),
    .Y(_0762_),
    .A1(_0747_),
    .A2(_0757_));
 sg13g2_a21oi_1 _2408_ (.A1(_0386_),
    .A2(net41),
    .Y(_0763_),
    .B1(net37));
 sg13g2_a21oi_1 _2409_ (.A1(_0762_),
    .A2(_0763_),
    .Y(_0764_),
    .B1(_0404_));
 sg13g2_nand2b_1 _2410_ (.Y(_0765_),
    .B(_0406_),
    .A_N(_0764_));
 sg13g2_nor2_1 _2411_ (.A(_0649_),
    .B(_0635_),
    .Y(_0766_));
 sg13g2_nand2_1 _2412_ (.Y(_0767_),
    .A(_0647_),
    .B(_0652_));
 sg13g2_nand2b_1 _2413_ (.Y(_0768_),
    .B(_0767_),
    .A_N(_0632_));
 sg13g2_nor2_1 _2414_ (.A(_0642_),
    .B(_0146_),
    .Y(_0769_));
 sg13g2_a21oi_1 _2415_ (.A1(_0748_),
    .A2(_0643_),
    .Y(_0770_),
    .B1(_0769_));
 sg13g2_a21oi_1 _2416_ (.A1(_0766_),
    .A2(_0768_),
    .Y(_0771_),
    .B1(_0770_));
 sg13g2_nor2b_1 _2417_ (.A(_0648_),
    .B_N(_0662_),
    .Y(_0772_));
 sg13g2_nand3_1 _2418_ (.B(_0661_),
    .C(_0772_),
    .A(_0766_),
    .Y(_0773_));
 sg13g2_nand2_1 _2419_ (.Y(_0774_),
    .A(_0771_),
    .B(_0773_));
 sg13g2_nor2b_1 _2420_ (.A(_0699_),
    .B_N(_0698_),
    .Y(_0775_));
 sg13g2_nand2_1 _2421_ (.Y(_0776_),
    .A(_0638_),
    .B(_0775_));
 sg13g2_inv_1 _2422_ (.Y(_0777_),
    .A(_0775_));
 sg13g2_nand3_1 _2423_ (.B(_0637_),
    .C(_0777_),
    .A(_0636_),
    .Y(_0778_));
 sg13g2_nand2_1 _2424_ (.Y(_0779_),
    .A(_0776_),
    .B(_0778_));
 sg13g2_xnor2_1 _2425_ (.Y(_0780_),
    .A(_0696_),
    .B(_0779_));
 sg13g2_nand2b_1 _2426_ (.Y(_0781_),
    .B(_0780_),
    .A_N(_0774_));
 sg13g2_xnor2_1 _2427_ (.Y(_0782_),
    .A(_0697_),
    .B(_0779_));
 sg13g2_nand2_1 _2428_ (.Y(_0783_),
    .A(_0782_),
    .B(_0774_));
 sg13g2_nand3_1 _2429_ (.B(_0783_),
    .C(_2038_),
    .A(_0781_),
    .Y(_0784_));
 sg13g2_nand2_1 _2430_ (.Y(_0785_),
    .A(_0784_),
    .B(_0285_));
 sg13g2_a21oi_1 _2431_ (.A1(_2053_),
    .A2(_2041_),
    .Y(_0786_),
    .B1(_0150_));
 sg13g2_nand2_1 _2432_ (.Y(_0787_),
    .A(_0785_),
    .B(_0786_));
 sg13g2_nor2b_1 _2433_ (.A(_0167_),
    .B_N(_2052_),
    .Y(_0788_));
 sg13g2_nor2_1 _2434_ (.A(_2052_),
    .B(_0168_),
    .Y(_0789_));
 sg13g2_nor3_1 _2435_ (.A(_0170_),
    .B(_0788_),
    .C(_0789_),
    .Y(_0790_));
 sg13g2_nor2_1 _2436_ (.A(_0154_),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_nand2_1 _2437_ (.Y(_0792_),
    .A(_0787_),
    .B(_0791_));
 sg13g2_a21oi_1 _2438_ (.A1(_2052_),
    .A2(_0154_),
    .Y(_0793_),
    .B1(_0176_));
 sg13g2_nand2_1 _2439_ (.Y(_0794_),
    .A(_0792_),
    .B(_0793_));
 sg13g2_nand2_1 _2440_ (.Y(_0795_),
    .A(_0794_),
    .B(_0223_));
 sg13g2_a21oi_1 _2441_ (.A1(_0795_),
    .A2(_0227_),
    .Y(_0796_),
    .B1(_0299_));
 sg13g2_a22oi_1 _2442_ (.Y(_0797_),
    .B1(net51),
    .B2(_0796_),
    .A2(_0765_),
    .A1(_0450_));
 sg13g2_nand3_1 _2443_ (.B(_0719_),
    .C(_0797_),
    .A(_0746_),
    .Y(_0798_));
 sg13g2_buf_8 _2444_ (.A(_0798_),
    .X(_0799_));
 sg13g2_inv_1 _2445_ (.Y(_0800_),
    .A(_0304_));
 sg13g2_nand2_1 _2446_ (.Y(_0801_),
    .A(_0715_),
    .B(_0225_));
 sg13g2_nand2_1 _2447_ (.Y(_0802_),
    .A(_0801_),
    .B(_0300_));
 sg13g2_a21oi_1 _2448_ (.A1(_0800_),
    .A2(_0247_),
    .Y(_0803_),
    .B1(_0802_));
 sg13g2_nand2_1 _2449_ (.Y(_0804_),
    .A(_0795_),
    .B(_0227_));
 sg13g2_nand2_1 _2450_ (.Y(_0805_),
    .A(_0804_),
    .B(_0237_));
 sg13g2_inv_1 _2451_ (.Y(_0806_),
    .A(_0343_));
 sg13g2_nor2_1 _2452_ (.A(_0806_),
    .B(_0740_),
    .Y(_0807_));
 sg13g2_nand2_1 _2453_ (.Y(_0808_),
    .A(_0765_),
    .B(_0410_));
 sg13g2_o21ai_1 _2454_ (.B1(_0326_),
    .Y(_0809_),
    .A1(net50),
    .A2(_0321_));
 sg13g2_xor2_1 _2455_ (.B(_0684_),
    .A(_0683_),
    .X(_0810_));
 sg13g2_nor2b_1 _2456_ (.A(_0656_),
    .B_N(_0654_),
    .Y(_0811_));
 sg13g2_xor2_1 _2457_ (.B(_0811_),
    .A(_0655_),
    .X(_0812_));
 sg13g2_xnor2_1 _2458_ (.Y(_0813_),
    .A(_0810_),
    .B(_0812_));
 sg13g2_a21oi_1 _2459_ (.A1(_0813_),
    .A2(net40),
    .Y(_0814_),
    .B1(_0425_));
 sg13g2_xnor2_1 _2460_ (.Y(_0815_),
    .A(_0163_),
    .B(net29));
 sg13g2_a21oi_1 _2461_ (.A1(_0815_),
    .A2(_0399_),
    .Y(_0816_),
    .B1(net41));
 sg13g2_o21ai_1 _2462_ (.B1(_0816_),
    .Y(_0817_),
    .A1(_0809_),
    .A2(_0814_));
 sg13g2_o21ai_1 _2463_ (.B1(_0817_),
    .Y(_0818_),
    .A1(_0329_),
    .A2(_0164_));
 sg13g2_o21ai_1 _2464_ (.B1(_0341_),
    .Y(_0819_),
    .A1(_0402_),
    .A2(_0818_));
 sg13g2_nand2_1 _2465_ (.Y(_0820_),
    .A(_0808_),
    .B(_0819_));
 sg13g2_nor2_1 _2466_ (.A(_0807_),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_o21ai_1 _2467_ (.B1(_0821_),
    .Y(_0822_),
    .A1(_0416_),
    .A2(_0805_));
 sg13g2_nor2_1 _2468_ (.A(_0803_),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_nand2_1 _2469_ (.Y(_0824_),
    .A(_0799_),
    .B(_0823_));
 sg13g2_nor2_1 _2470_ (.A(_0745_),
    .B(_0824_),
    .Y(_0825_));
 sg13g2_xor2_1 _2471_ (.B(_0750_),
    .A(_0677_),
    .X(_0826_));
 sg13g2_xnor2_1 _2472_ (.Y(_0827_),
    .A(_0647_),
    .B(_0664_));
 sg13g2_xnor2_1 _2473_ (.Y(_0828_),
    .A(_0826_),
    .B(_0827_));
 sg13g2_inv_1 _2474_ (.Y(_0829_),
    .A(_0381_));
 sg13g2_o21ai_1 _2475_ (.B1(_0829_),
    .Y(_0830_),
    .A1(_0316_),
    .A2(_0828_));
 sg13g2_a21oi_1 _2476_ (.A1(_0504_),
    .A2(net49),
    .Y(_0831_),
    .B1(net45));
 sg13g2_nand2_1 _2477_ (.Y(_0832_),
    .A(_0830_),
    .B(_0831_));
 sg13g2_nand2_1 _2478_ (.Y(_0833_),
    .A(_0169_),
    .B(_0507_));
 sg13g2_nand2b_1 _2479_ (.Y(_0834_),
    .B(net29),
    .A_N(_0507_));
 sg13g2_nand3_1 _2480_ (.B(net39),
    .C(_0834_),
    .A(_0833_),
    .Y(_0835_));
 sg13g2_nand3_1 _2481_ (.B(_0155_),
    .C(_0835_),
    .A(_0832_),
    .Y(_0836_));
 sg13g2_a21oi_1 _2482_ (.A1(_0507_),
    .A2(_0334_),
    .Y(_0837_),
    .B1(_0402_));
 sg13g2_a21oi_1 _2483_ (.A1(_0836_),
    .A2(_0837_),
    .Y(_0838_),
    .B1(_0221_));
 sg13g2_nor2_1 _2484_ (.A(net56),
    .B(_0838_),
    .Y(_0839_));
 sg13g2_nor2b_1 _2485_ (.A(_0839_),
    .B_N(_0524_),
    .Y(_0840_));
 sg13g2_a21oi_1 _2486_ (.A1(_0796_),
    .A2(net54),
    .Y(_0841_),
    .B1(_0840_));
 sg13g2_nor2_1 _2487_ (.A(_0528_),
    .B(_0245_),
    .Y(_0842_));
 sg13g2_nand3_1 _2488_ (.B(_0717_),
    .C(_0842_),
    .A(_0841_),
    .Y(_0843_));
 sg13g2_nand2b_1 _2489_ (.Y(_0844_),
    .B(_0802_),
    .A_N(_0841_));
 sg13g2_nand2_1 _2490_ (.Y(_0845_),
    .A(_0843_),
    .B(_0844_));
 sg13g2_nand3_1 _2491_ (.B(_0414_),
    .C(net51),
    .A(_0804_),
    .Y(_0846_));
 sg13g2_nand2_1 _2492_ (.Y(_0847_),
    .A(_0846_),
    .B(net31));
 sg13g2_nand2_1 _2493_ (.Y(_0848_),
    .A(_0804_),
    .B(net23));
 sg13g2_nand3_1 _2494_ (.B(_0414_),
    .C(net54),
    .A(_0739_),
    .Y(_0849_));
 sg13g2_nand2_1 _2495_ (.Y(_0850_),
    .A(_0687_),
    .B(_0688_));
 sg13g2_nand2_1 _2496_ (.Y(_0851_),
    .A(_0850_),
    .B(_0671_));
 sg13g2_xnor2_1 _2497_ (.Y(_0852_),
    .A(_0672_),
    .B(_0851_));
 sg13g2_xnor2_1 _2498_ (.Y(_0853_),
    .A(_0662_),
    .B(_0661_));
 sg13g2_xnor2_1 _2499_ (.Y(_0854_),
    .A(_0852_),
    .B(_0853_));
 sg13g2_inv_1 _2500_ (.Y(_0855_),
    .A(_0505_));
 sg13g2_o21ai_1 _2501_ (.B1(_0855_),
    .Y(_0856_),
    .A1(_0316_),
    .A2(_0854_));
 sg13g2_a21oi_1 _2502_ (.A1(_0470_),
    .A2(net49),
    .Y(_0857_),
    .B1(net45));
 sg13g2_nand2_1 _2503_ (.Y(_0858_),
    .A(_0856_),
    .B(_0857_));
 sg13g2_nand2_1 _2504_ (.Y(_0859_),
    .A(net27),
    .B(_0473_));
 sg13g2_nand2b_1 _2505_ (.Y(_0860_),
    .B(net29),
    .A_N(_0473_));
 sg13g2_nand3_1 _2506_ (.B(net39),
    .C(_0860_),
    .A(_0859_),
    .Y(_0861_));
 sg13g2_nand3_1 _2507_ (.B(net42),
    .C(_0861_),
    .A(_0858_),
    .Y(_0862_));
 sg13g2_a21oi_1 _2508_ (.A1(_0473_),
    .A2(net35),
    .Y(_0863_),
    .B1(net30));
 sg13g2_a21oi_1 _2509_ (.A1(_0862_),
    .A2(_0863_),
    .Y(_0864_),
    .B1(_0221_));
 sg13g2_o21ai_1 _2510_ (.B1(_0486_),
    .Y(_0865_),
    .A1(net56),
    .A2(_0864_));
 sg13g2_nand3_1 _2511_ (.B(_0849_),
    .C(_0865_),
    .A(_0848_),
    .Y(_0866_));
 sg13g2_nor2_1 _2512_ (.A(_0847_),
    .B(_0866_),
    .Y(_0867_));
 sg13g2_nand2_1 _2513_ (.Y(_0868_),
    .A(_0717_),
    .B(_0343_));
 sg13g2_nand2_1 _2514_ (.Y(_0869_),
    .A(_0867_),
    .B(_0868_));
 sg13g2_nand2_1 _2515_ (.Y(_0870_),
    .A(_0848_),
    .B(_0246_));
 sg13g2_nor2_1 _2516_ (.A(_0420_),
    .B(_0805_),
    .Y(_0871_));
 sg13g2_nor2_1 _2517_ (.A(_0870_),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_o21ai_1 _2518_ (.B1(_0796_),
    .Y(_0873_),
    .A1(_0343_),
    .A2(_0417_));
 sg13g2_nand2_1 _2519_ (.Y(_0874_),
    .A(_0872_),
    .B(_0873_));
 sg13g2_nand2_1 _2520_ (.Y(_0875_),
    .A(_0802_),
    .B(_0245_));
 sg13g2_nand2_1 _2521_ (.Y(_0876_),
    .A(_0874_),
    .B(_0875_));
 sg13g2_nor2_1 _2522_ (.A(_0869_),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_nor2_1 _2523_ (.A(_0845_),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_nand3_1 _2524_ (.B(_0869_),
    .C(_0875_),
    .A(_0876_),
    .Y(_0879_));
 sg13g2_nand2_1 _2525_ (.Y(_0880_),
    .A(_0878_),
    .B(_0879_));
 sg13g2_nor2_1 _2526_ (.A(_0825_),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_nand2_1 _2527_ (.Y(_0882_),
    .A(_0824_),
    .B(_0745_));
 sg13g2_nor2_1 _2528_ (.A(_0806_),
    .B(_0805_),
    .Y(_0883_));
 sg13g2_a21oi_1 _2529_ (.A1(_0739_),
    .A2(_0410_),
    .Y(_0884_),
    .B1(_0245_));
 sg13g2_o21ai_1 _2530_ (.B1(net36),
    .Y(_0885_),
    .A1(net50),
    .A2(_0423_));
 sg13g2_xnor2_1 _2531_ (.Y(_0886_),
    .A(_0689_),
    .B(_0687_));
 sg13g2_xnor2_1 _2532_ (.Y(_0887_),
    .A(_0657_),
    .B(_0653_));
 sg13g2_xnor2_1 _2533_ (.Y(_0888_),
    .A(_0886_),
    .B(_0887_));
 sg13g2_a21oi_1 _2534_ (.A1(_0888_),
    .A2(net40),
    .Y(_0889_),
    .B1(_0471_));
 sg13g2_xnor2_1 _2535_ (.Y(_0890_),
    .A(_0432_),
    .B(net25));
 sg13g2_a21oi_1 _2536_ (.A1(_0890_),
    .A2(net39),
    .Y(_0891_),
    .B1(net35));
 sg13g2_o21ai_1 _2537_ (.B1(_0891_),
    .Y(_0892_),
    .A1(_0885_),
    .A2(_0889_));
 sg13g2_o21ai_1 _2538_ (.B1(_0892_),
    .Y(_0893_),
    .A1(net42),
    .A2(_0431_));
 sg13g2_o21ai_1 _2539_ (.B1(_0422_),
    .Y(_0894_),
    .A1(net30),
    .A2(_0893_));
 sg13g2_nand3b_1 _2540_ (.B(_0884_),
    .C(_0894_),
    .Y(_0895_),
    .A_N(_0883_));
 sg13g2_a22oi_1 _2541_ (.Y(_0896_),
    .B1(_0875_),
    .B2(_0895_),
    .A2(_0717_),
    .A1(_0417_));
 sg13g2_buf_1 _2542_ (.A(_0896_),
    .X(_0897_));
 sg13g2_nand2_1 _2543_ (.Y(_0898_),
    .A(_0882_),
    .B(_0897_));
 sg13g2_nand2_1 _2544_ (.Y(_0899_),
    .A(_0881_),
    .B(_0898_));
 sg13g2_buf_8 _2545_ (.A(_0899_),
    .X(_0900_));
 sg13g2_inv_1 _2546_ (.Y(_0901_),
    .A(_0844_));
 sg13g2_nor2_1 _2547_ (.A(_0845_),
    .B(_0879_),
    .Y(_0902_));
 sg13g2_nor2_1 _2548_ (.A(_0901_),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_buf_2 _2549_ (.A(_0903_),
    .X(_0904_));
 sg13g2_nand2_1 _2550_ (.Y(_0905_),
    .A(_0900_),
    .B(_0904_));
 sg13g2_inv_1 _2551_ (.Y(_0906_),
    .A(_0799_));
 sg13g2_nand2_1 _2552_ (.Y(_0907_),
    .A(_0905_),
    .B(_0906_));
 sg13g2_nand3_1 _2553_ (.B(_0799_),
    .C(_0904_),
    .A(_0900_),
    .Y(_0908_));
 sg13g2_nand2_1 _2554_ (.Y(_0909_),
    .A(_0907_),
    .B(_0908_));
 sg13g2_nand2b_1 _2555_ (.Y(_0910_),
    .B(_0909_),
    .A_N(_0823_));
 sg13g2_nand3_1 _2556_ (.B(_0908_),
    .C(_0823_),
    .A(_0907_),
    .Y(_0911_));
 sg13g2_buf_1 _2557_ (.A(_0911_),
    .X(_0912_));
 sg13g2_inv_1 _2558_ (.Y(_0913_),
    .A(_0029_));
 sg13g2_a21oi_1 _2559_ (.A1(_0910_),
    .A2(_0912_),
    .Y(_0914_),
    .B1(_0913_));
 sg13g2_nand2_1 _2560_ (.Y(_0915_),
    .A(_0905_),
    .B(_0744_));
 sg13g2_xnor2_1 _2561_ (.Y(_0916_),
    .A(_0799_),
    .B(_0744_));
 sg13g2_nand3_1 _2562_ (.B(_0904_),
    .C(_0916_),
    .A(_0900_),
    .Y(_0917_));
 sg13g2_nand2_2 _2563_ (.Y(_0918_),
    .A(_0915_),
    .B(_0917_));
 sg13g2_nand2_1 _2564_ (.Y(_0919_),
    .A(_0918_),
    .B(_0897_));
 sg13g2_nor2_1 _2565_ (.A(_0897_),
    .B(_0918_),
    .Y(_0920_));
 sg13g2_a21oi_2 _2566_ (.B1(_0920_),
    .Y(_0921_),
    .A2(_0912_),
    .A1(_0919_));
 sg13g2_nand2_1 _2567_ (.Y(_0922_),
    .A(_0869_),
    .B(_0875_));
 sg13g2_nand2_1 _2568_ (.Y(_0923_),
    .A(_0905_),
    .B(_0876_));
 sg13g2_inv_1 _2569_ (.Y(_0924_),
    .A(_0876_));
 sg13g2_nor2_1 _2570_ (.A(_0799_),
    .B(_0744_),
    .Y(_0925_));
 sg13g2_xnor2_1 _2571_ (.Y(_0926_),
    .A(_0924_),
    .B(_0925_));
 sg13g2_nand3_1 _2572_ (.B(_0904_),
    .C(_0926_),
    .A(_0900_),
    .Y(_0927_));
 sg13g2_nand2_1 _2573_ (.Y(_0928_),
    .A(_0923_),
    .B(_0927_));
 sg13g2_xnor2_1 _2574_ (.Y(_0929_),
    .A(_0922_),
    .B(_0928_));
 sg13g2_nand2_1 _2575_ (.Y(_0930_),
    .A(_0905_),
    .B(_0717_));
 sg13g2_nor2_1 _2576_ (.A(_0924_),
    .B(_0744_),
    .Y(_0931_));
 sg13g2_nand2_1 _2577_ (.Y(_0932_),
    .A(_0931_),
    .B(_0906_));
 sg13g2_xnor2_1 _2578_ (.Y(_0933_),
    .A(_0717_),
    .B(_0932_));
 sg13g2_nand3_1 _2579_ (.B(_0933_),
    .C(_0904_),
    .A(_0900_),
    .Y(_0934_));
 sg13g2_nand2_1 _2580_ (.Y(_0935_),
    .A(_0930_),
    .B(_0934_));
 sg13g2_o21ai_1 _2581_ (.B1(_0841_),
    .Y(_0936_),
    .A1(_0842_),
    .A2(_0802_));
 sg13g2_inv_1 _2582_ (.Y(_0937_),
    .A(_0936_));
 sg13g2_a21oi_1 _2583_ (.A1(_0935_),
    .A2(_0937_),
    .Y(_0938_),
    .B1(_0901_));
 sg13g2_nand2_1 _2584_ (.Y(_0939_),
    .A(_0929_),
    .B(_0938_));
 sg13g2_nor2_1 _2585_ (.A(_0921_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_nand3_1 _2586_ (.B(_0900_),
    .C(_0904_),
    .A(_0940_),
    .Y(_0941_));
 sg13g2_nand2_1 _2587_ (.Y(_0942_),
    .A(_0941_),
    .B(_1706_));
 sg13g2_nand4_1 _2588_ (.B(_1670_),
    .C(_0900_),
    .A(_0940_),
    .Y(_0943_),
    .D(_0904_));
 sg13g2_nand2_1 _2589_ (.Y(_0944_),
    .A(_0942_),
    .B(_0943_));
 sg13g2_nand2b_1 _2590_ (.Y(_0945_),
    .B(_0918_),
    .A_N(_0897_));
 sg13g2_nand3_1 _2591_ (.B(_0917_),
    .C(_0897_),
    .A(_0915_),
    .Y(_0946_));
 sg13g2_nand2_1 _2592_ (.Y(_0947_),
    .A(_0945_),
    .B(_0946_));
 sg13g2_xnor2_1 _2593_ (.Y(_0948_),
    .A(_0912_),
    .B(_0947_));
 sg13g2_xnor2_1 _2594_ (.Y(_0949_),
    .A(_0018_),
    .B(_0948_));
 sg13g2_xor2_1 _2595_ (.B(_0921_),
    .A(_0929_),
    .X(_0950_));
 sg13g2_nand2_1 _2596_ (.Y(_0951_),
    .A(_0950_),
    .B(_1665_));
 sg13g2_xnor2_1 _2597_ (.Y(_0952_),
    .A(_0929_),
    .B(_0921_));
 sg13g2_nand2_1 _2598_ (.Y(_0953_),
    .A(_0952_),
    .B(_1664_));
 sg13g2_nand3_1 _2599_ (.B(_0951_),
    .C(_0953_),
    .A(_0949_),
    .Y(_0954_));
 sg13g2_nand3_1 _2600_ (.B(_0947_),
    .C(_0912_),
    .A(_0929_),
    .Y(_0955_));
 sg13g2_inv_1 _2601_ (.Y(_0956_),
    .A(_0928_));
 sg13g2_nand2_1 _2602_ (.Y(_0957_),
    .A(_0956_),
    .B(_0922_));
 sg13g2_nor2_1 _2603_ (.A(_0922_),
    .B(_0956_),
    .Y(_0958_));
 sg13g2_a21oi_1 _2604_ (.A1(_0957_),
    .A2(_0920_),
    .Y(_0959_),
    .B1(_0958_));
 sg13g2_nand2_1 _2605_ (.Y(_0960_),
    .A(_0955_),
    .B(_0959_));
 sg13g2_nand2_1 _2606_ (.Y(_0961_),
    .A(_0960_),
    .B(_0938_));
 sg13g2_inv_1 _2607_ (.Y(_0962_),
    .A(_0938_));
 sg13g2_nand3_1 _2608_ (.B(_0959_),
    .C(_0962_),
    .A(_0955_),
    .Y(_0963_));
 sg13g2_nand2_1 _2609_ (.Y(_0964_),
    .A(_0961_),
    .B(_0963_));
 sg13g2_nand2_1 _2610_ (.Y(_0965_),
    .A(_0964_),
    .B(_0581_));
 sg13g2_nand3_1 _2611_ (.B(_0963_),
    .C(_1698_),
    .A(_0961_),
    .Y(_0966_));
 sg13g2_nand2_1 _2612_ (.Y(_0967_),
    .A(_0965_),
    .B(_0966_));
 sg13g2_nor4_1 _2613_ (.A(_0914_),
    .B(_0944_),
    .C(_0954_),
    .D(_0967_),
    .Y(_0968_));
 sg13g2_nor2_1 _2614_ (.A(_0944_),
    .B(_0967_),
    .Y(_0969_));
 sg13g2_inv_1 _2615_ (.Y(_0970_),
    .A(_0948_));
 sg13g2_nor2_1 _2616_ (.A(_0018_),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_nand3_1 _2617_ (.B(_0953_),
    .C(_0971_),
    .A(_0951_),
    .Y(_0972_));
 sg13g2_nand2_1 _2618_ (.Y(_0973_),
    .A(_0950_),
    .B(_1658_));
 sg13g2_nand2_1 _2619_ (.Y(_0974_),
    .A(_0972_),
    .B(_0973_));
 sg13g2_nand2_1 _2620_ (.Y(_0975_),
    .A(_0969_),
    .B(_0974_));
 sg13g2_nand2_1 _2621_ (.Y(_0976_),
    .A(_0964_),
    .B(_1657_));
 sg13g2_nor2_1 _2622_ (.A(_0976_),
    .B(_0944_),
    .Y(_0977_));
 sg13g2_a21oi_1 _2623_ (.A1(\dither_threshold[4] ),
    .A2(_0941_),
    .Y(_0978_),
    .B1(_0977_));
 sg13g2_nand2_1 _2624_ (.Y(_0979_),
    .A(_0975_),
    .B(_0978_));
 sg13g2_nor2_2 _2625_ (.A(_0968_),
    .B(_0979_),
    .Y(_0980_));
 sg13g2_xnor2_1 _2626_ (.Y(net14),
    .A(_0909_),
    .B(_0980_));
 sg13g2_inv_1 _2627_ (.Y(_0981_),
    .A(_0909_));
 sg13g2_a21oi_1 _2628_ (.A1(_0980_),
    .A2(_0981_),
    .Y(_0982_),
    .B1(_0918_));
 sg13g2_nand3_1 _2629_ (.B(_0981_),
    .C(_0918_),
    .A(_0980_),
    .Y(_0983_));
 sg13g2_nor2b_1 _2630_ (.A(_0982_),
    .B_N(_0983_),
    .Y(net15));
 sg13g2_nand2_1 _2631_ (.Y(_0984_),
    .A(_0983_),
    .B(_0956_));
 sg13g2_nand4_1 _2632_ (.B(_0981_),
    .C(_0928_),
    .A(_0980_),
    .Y(_0985_),
    .D(_0918_));
 sg13g2_nand2_1 _2633_ (.Y(net16),
    .A(_0984_),
    .B(_0985_));
 sg13g2_a21oi_1 _2634_ (.A1(_0917_),
    .A2(_0915_),
    .Y(_0986_),
    .B1(_0928_));
 sg13g2_nand3_1 _2635_ (.B(_0981_),
    .C(_0986_),
    .A(_0980_),
    .Y(_0987_));
 sg13g2_nand2_1 _2636_ (.Y(_0988_),
    .A(_0987_),
    .B(_0935_));
 sg13g2_inv_1 _2637_ (.Y(_0989_),
    .A(_0935_));
 sg13g2_nand4_1 _2638_ (.B(_0981_),
    .C(_0989_),
    .A(_0980_),
    .Y(_0990_),
    .D(_0986_));
 sg13g2_nand2_1 _2639_ (.Y(net17),
    .A(_0988_),
    .B(_0990_));
 sg13g2_nand2_1 _2640_ (.Y(_0991_),
    .A(_1519_),
    .B(_1844_));
 sg13g2_nand2_1 _2641_ (.Y(_0992_),
    .A(_1518_),
    .B(net72));
 sg13g2_nand2_1 _2642_ (.Y(_0993_),
    .A(_0991_),
    .B(_0992_));
 sg13g2_inv_1 _2643_ (.Y(_0994_),
    .A(_0993_));
 sg13g2_nand2_1 _2644_ (.Y(_0995_),
    .A(_1977_),
    .B(_0994_));
 sg13g2_nand3_1 _2645_ (.B(_1976_),
    .C(_0993_),
    .A(_1975_),
    .Y(_0996_));
 sg13g2_xor2_1 _2646_ (.B(net71),
    .A(_1520_),
    .X(_0997_));
 sg13g2_nand2_1 _2647_ (.Y(_0998_),
    .A(net38),
    .B(_0997_));
 sg13g2_nand2_1 _2648_ (.Y(_0999_),
    .A(net68),
    .B(net71));
 sg13g2_nand2_1 _2649_ (.Y(_1000_),
    .A(_0998_),
    .B(_0999_));
 sg13g2_nand3_1 _2650_ (.B(_0996_),
    .C(_1000_),
    .A(_0995_),
    .Y(_1001_));
 sg13g2_inv_1 _2651_ (.Y(_1002_),
    .A(_1001_));
 sg13g2_nand2_1 _2652_ (.Y(_1003_),
    .A(_1556_),
    .B(_1970_));
 sg13g2_nand2_1 _2653_ (.Y(_1004_),
    .A(_1524_),
    .B(_1853_));
 sg13g2_nand2_1 _2654_ (.Y(_1005_),
    .A(_1003_),
    .B(_1004_));
 sg13g2_inv_1 _2655_ (.Y(_1006_),
    .A(_1005_));
 sg13g2_nand2_1 _2656_ (.Y(_1007_),
    .A(_1916_),
    .B(_1006_));
 sg13g2_nand2_1 _2657_ (.Y(_1008_),
    .A(_1909_),
    .B(_1005_));
 sg13g2_nand2_1 _2658_ (.Y(_1009_),
    .A(_1007_),
    .B(_1008_));
 sg13g2_nand2_1 _2659_ (.Y(_1010_),
    .A(_0995_),
    .B(_0992_));
 sg13g2_inv_1 _2660_ (.Y(_1011_),
    .A(_1010_));
 sg13g2_nor2_1 _2661_ (.A(_1009_),
    .B(_1011_),
    .Y(_1012_));
 sg13g2_nand2_1 _2662_ (.Y(_1013_),
    .A(_1011_),
    .B(_1009_));
 sg13g2_o21ai_1 _2663_ (.B1(_1013_),
    .Y(_1014_),
    .A1(_1002_),
    .A2(_1012_));
 sg13g2_xor2_1 _2664_ (.B(_1857_),
    .A(_1532_),
    .X(_1015_));
 sg13g2_inv_1 _2665_ (.Y(_1016_),
    .A(_1015_));
 sg13g2_xnor2_1 _2666_ (.Y(_1017_),
    .A(_1016_),
    .B(net32));
 sg13g2_nand2_1 _2667_ (.Y(_1018_),
    .A(_1527_),
    .B(_1842_));
 sg13g2_nand2_1 _2668_ (.Y(_1019_),
    .A(net64),
    .B(net73));
 sg13g2_inv_1 _2669_ (.Y(_1020_),
    .A(_1019_));
 sg13g2_a21oi_1 _2670_ (.A1(net34),
    .A2(_1018_),
    .Y(_1021_),
    .B1(_1020_));
 sg13g2_nand2_1 _2671_ (.Y(_1022_),
    .A(_1017_),
    .B(_1021_));
 sg13g2_nand2_1 _2672_ (.Y(_1023_),
    .A(_2007_),
    .B(_1015_));
 sg13g2_nand3_1 _2673_ (.B(_2005_),
    .C(_1016_),
    .A(_2004_),
    .Y(_1024_));
 sg13g2_nand2_1 _2674_ (.Y(_1025_),
    .A(_1023_),
    .B(_1024_));
 sg13g2_nand2_1 _2675_ (.Y(_1026_),
    .A(_1018_),
    .B(_1019_));
 sg13g2_nand2b_1 _2676_ (.Y(_1027_),
    .B(net34),
    .A_N(_1026_));
 sg13g2_nand2_1 _2677_ (.Y(_1028_),
    .A(_1027_),
    .B(_1019_));
 sg13g2_nand2_1 _2678_ (.Y(_1029_),
    .A(_1025_),
    .B(_1028_));
 sg13g2_nand2_1 _2679_ (.Y(_1030_),
    .A(_1022_),
    .B(_1029_));
 sg13g2_nand3_1 _2680_ (.B(_1940_),
    .C(_1026_),
    .A(_1939_),
    .Y(_1031_));
 sg13g2_nand2_1 _2681_ (.Y(_1032_),
    .A(_1027_),
    .B(_1031_));
 sg13g2_nand2_1 _2682_ (.Y(_1033_),
    .A(_1007_),
    .B(_1004_));
 sg13g2_nand2_1 _2683_ (.Y(_1034_),
    .A(_1032_),
    .B(_1033_));
 sg13g2_inv_1 _2684_ (.Y(_1035_),
    .A(_1004_));
 sg13g2_a21oi_1 _2685_ (.A1(_1916_),
    .A2(_1003_),
    .Y(_1036_),
    .B1(_1035_));
 sg13g2_nand3_1 _2686_ (.B(_1036_),
    .C(_1031_),
    .A(_1027_),
    .Y(_1037_));
 sg13g2_nand2_1 _2687_ (.Y(_1038_),
    .A(_1034_),
    .B(_1037_));
 sg13g2_nand2_1 _2688_ (.Y(_1039_),
    .A(_1030_),
    .B(_1038_));
 sg13g2_nor2_1 _2689_ (.A(_1014_),
    .B(_1039_),
    .Y(_1040_));
 sg13g2_nand3_1 _2690_ (.B(_1031_),
    .C(_1033_),
    .A(_1027_),
    .Y(_1041_));
 sg13g2_inv_1 _2691_ (.Y(_1042_),
    .A(_1041_));
 sg13g2_nand2_1 _2692_ (.Y(_1043_),
    .A(_1025_),
    .B(_1021_));
 sg13g2_nor2_1 _2693_ (.A(_1021_),
    .B(_1025_),
    .Y(_1044_));
 sg13g2_a21oi_1 _2694_ (.A1(_1042_),
    .A2(_1043_),
    .Y(_1045_),
    .B1(_1044_));
 sg13g2_nor2b_1 _2695_ (.A(_1040_),
    .B_N(_1045_),
    .Y(_1046_));
 sg13g2_xor2_1 _2696_ (.B(_1845_),
    .A(net79),
    .X(_1047_));
 sg13g2_nand2_1 _2697_ (.Y(_1048_),
    .A(net44),
    .B(_1047_));
 sg13g2_o21ai_1 _2698_ (.B1(_1048_),
    .Y(_1049_),
    .A1(_1516_),
    .A2(_1846_));
 sg13g2_xor2_1 _2699_ (.B(net38),
    .A(_0997_),
    .X(_1050_));
 sg13g2_nor2_1 _2700_ (.A(_1049_),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_xnor2_1 _2701_ (.Y(_1052_),
    .A(_1047_),
    .B(net44));
 sg13g2_nor2_1 _2702_ (.A(_1836_),
    .B(_1963_),
    .Y(_1053_));
 sg13g2_nand2_1 _2703_ (.Y(_1054_),
    .A(_1052_),
    .B(_1053_));
 sg13g2_xnor2_1 _2704_ (.Y(_1055_),
    .A(_1847_),
    .B(_1963_));
 sg13g2_nor2_1 _2705_ (.A(_0193_),
    .B(_1055_),
    .Y(_1056_));
 sg13g2_nor2_1 _2706_ (.A(_1053_),
    .B(_1052_),
    .Y(_1057_));
 sg13g2_a21oi_2 _2707_ (.B1(_1057_),
    .Y(_1058_),
    .A2(_1056_),
    .A1(_1054_));
 sg13g2_nand2_1 _2708_ (.Y(_1059_),
    .A(_1050_),
    .B(_1049_));
 sg13g2_o21ai_1 _2709_ (.B1(_1059_),
    .Y(_1060_),
    .A1(_1051_),
    .A2(_1058_));
 sg13g2_xnor2_1 _2710_ (.Y(_1061_),
    .A(_1006_),
    .B(_1909_));
 sg13g2_nand2_1 _2711_ (.Y(_1062_),
    .A(_1061_),
    .B(_1011_));
 sg13g2_nand2_1 _2712_ (.Y(_1063_),
    .A(_1009_),
    .B(_1010_));
 sg13g2_nand2_2 _2713_ (.Y(_1064_),
    .A(_1062_),
    .B(_1063_));
 sg13g2_nand2_1 _2714_ (.Y(_1065_),
    .A(_0995_),
    .B(_0996_));
 sg13g2_xnor2_1 _2715_ (.Y(_1066_),
    .A(_1000_),
    .B(_1065_));
 sg13g2_nand3_1 _2716_ (.B(_1064_),
    .C(_1066_),
    .A(_1060_),
    .Y(_1067_));
 sg13g2_or2_1 _2717_ (.X(_1068_),
    .B(_1039_),
    .A(_1067_));
 sg13g2_nand2_1 _2718_ (.Y(_1069_),
    .A(_1046_),
    .B(_1068_));
 sg13g2_o21ai_1 _2719_ (.B1(_1023_),
    .Y(_1070_),
    .A1(_1548_),
    .A2(_0253_));
 sg13g2_xor2_1 _2720_ (.B(net70),
    .A(_1534_),
    .X(_1071_));
 sg13g2_xnor2_1 _2721_ (.Y(_1072_),
    .A(_1071_),
    .B(net26));
 sg13g2_xnor2_1 _2722_ (.Y(_1073_),
    .A(_1070_),
    .B(_1072_));
 sg13g2_nand2_1 _2723_ (.Y(_1074_),
    .A(_1069_),
    .B(_1073_));
 sg13g2_inv_1 _2724_ (.Y(_1075_),
    .A(_1073_));
 sg13g2_nand3_1 _2725_ (.B(_1068_),
    .C(_1075_),
    .A(_1046_),
    .Y(_1076_));
 sg13g2_nand3_1 _2726_ (.B(_1076_),
    .C(_2041_),
    .A(_1074_),
    .Y(_1077_));
 sg13g2_xor2_1 _2727_ (.B(_1859_),
    .A(net66),
    .X(_1078_));
 sg13g2_nand2_1 _2728_ (.Y(_1079_),
    .A(net68),
    .B(net72));
 sg13g2_xnor2_1 _2729_ (.Y(_1080_),
    .A(net65),
    .B(net61));
 sg13g2_nand2_1 _2730_ (.Y(_1081_),
    .A(net65),
    .B(net61));
 sg13g2_o21ai_1 _2731_ (.B1(_1081_),
    .Y(_1082_),
    .A1(_1079_),
    .A2(_1080_));
 sg13g2_xnor2_1 _2732_ (.Y(_1083_),
    .A(net67),
    .B(net73));
 sg13g2_xnor2_1 _2733_ (.Y(_1084_),
    .A(net64),
    .B(net60));
 sg13g2_nor2_1 _2734_ (.A(_1083_),
    .B(_1084_),
    .Y(_1085_));
 sg13g2_nand2_1 _2735_ (.Y(_1086_),
    .A(net67),
    .B(net73));
 sg13g2_nand2_1 _2736_ (.Y(_1087_),
    .A(net64),
    .B(net60));
 sg13g2_o21ai_1 _2737_ (.B1(_1087_),
    .Y(_1088_),
    .A1(_1086_),
    .A2(_1084_));
 sg13g2_a21oi_1 _2738_ (.A1(_1082_),
    .A2(_1085_),
    .Y(_1089_),
    .B1(_1088_));
 sg13g2_nand2_1 _2739_ (.Y(_1090_),
    .A(net80),
    .B(_1845_));
 sg13g2_xnor2_1 _2740_ (.Y(_1091_),
    .A(net79),
    .B(net71));
 sg13g2_nand2_1 _2741_ (.Y(_1092_),
    .A(net79),
    .B(_1849_));
 sg13g2_o21ai_1 _2742_ (.B1(_1092_),
    .Y(_1093_),
    .A1(_1090_),
    .A2(_1091_));
 sg13g2_buf_1 _2743_ (.A(_1093_),
    .X(_1094_));
 sg13g2_xor2_1 _2744_ (.B(net72),
    .A(net68),
    .X(_1095_));
 sg13g2_nor2b_1 _2745_ (.A(_1080_),
    .B_N(_1095_),
    .Y(_1096_));
 sg13g2_nand3_1 _2746_ (.B(_1096_),
    .C(_1085_),
    .A(_1094_),
    .Y(_1097_));
 sg13g2_nand2_1 _2747_ (.Y(_1098_),
    .A(_1089_),
    .B(_1097_));
 sg13g2_xnor2_1 _2748_ (.Y(_1099_),
    .A(_1078_),
    .B(_1098_));
 sg13g2_xnor2_1 _2749_ (.Y(_1100_),
    .A(_0264_),
    .B(net32));
 sg13g2_xnor2_1 _2750_ (.Y(_1101_),
    .A(_1099_),
    .B(_1100_));
 sg13g2_xnor2_1 _2751_ (.Y(_1102_),
    .A(_1936_),
    .B(_1909_));
 sg13g2_inv_1 _2752_ (.Y(_1103_),
    .A(_1102_));
 sg13g2_nand2_1 _2753_ (.Y(_1104_),
    .A(net33),
    .B(_1910_));
 sg13g2_nor2_1 _2754_ (.A(_0043_),
    .B(net38),
    .Y(_1105_));
 sg13g2_nor2_1 _2755_ (.A(_1910_),
    .B(net33),
    .Y(_1106_));
 sg13g2_a21oi_1 _2756_ (.A1(_1104_),
    .A2(_1105_),
    .Y(_1107_),
    .B1(_1106_));
 sg13g2_nand2_1 _2757_ (.Y(_1108_),
    .A(net34),
    .B(_1994_));
 sg13g2_nand2_1 _2758_ (.Y(_1109_),
    .A(_1935_),
    .B(_0256_));
 sg13g2_nand2_1 _2759_ (.Y(_1110_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_nor3_1 _2760_ (.A(_1103_),
    .B(_1107_),
    .C(_1110_),
    .Y(_1111_));
 sg13g2_nor2_1 _2761_ (.A(_1936_),
    .B(_1916_),
    .Y(_1112_));
 sg13g2_inv_1 _2762_ (.Y(_1113_),
    .A(_1109_));
 sg13g2_a21oi_1 _2763_ (.A1(_1108_),
    .A2(_1112_),
    .Y(_1114_),
    .B1(_1113_));
 sg13g2_nor2b_1 _2764_ (.A(_1111_),
    .B_N(_1114_),
    .Y(_1115_));
 sg13g2_nor2_1 _2765_ (.A(_1103_),
    .B(_1110_),
    .Y(_1116_));
 sg13g2_xnor2_1 _2766_ (.Y(_1117_),
    .A(net72),
    .B(net44));
 sg13g2_nor2_1 _2767_ (.A(_0312_),
    .B(_1963_),
    .Y(_1118_));
 sg13g2_nand2_1 _2768_ (.Y(_1119_),
    .A(_1117_),
    .B(_1118_));
 sg13g2_nand2_1 _2769_ (.Y(_1120_),
    .A(_1966_),
    .B(_1983_));
 sg13g2_nand2_2 _2770_ (.Y(_1121_),
    .A(_1119_),
    .B(_1120_));
 sg13g2_nand2_1 _2771_ (.Y(_1122_),
    .A(net33),
    .B(_1911_));
 sg13g2_nand3_1 _2772_ (.B(_1976_),
    .C(_1910_),
    .A(_1975_),
    .Y(_1123_));
 sg13g2_nand2_1 _2773_ (.Y(_1124_),
    .A(_1122_),
    .B(_1123_));
 sg13g2_inv_1 _2774_ (.Y(_1125_),
    .A(_1124_));
 sg13g2_xnor2_1 _2775_ (.Y(_1126_),
    .A(_1853_),
    .B(net38));
 sg13g2_nor2b_1 _2776_ (.A(_1125_),
    .B_N(_1126_),
    .Y(_1127_));
 sg13g2_nand3_1 _2777_ (.B(_1121_),
    .C(_1127_),
    .A(_1116_),
    .Y(_1128_));
 sg13g2_nand2_1 _2778_ (.Y(_1129_),
    .A(_1115_),
    .B(_1128_));
 sg13g2_nand2b_1 _2779_ (.Y(_1130_),
    .B(_1129_),
    .A_N(_1101_));
 sg13g2_nand3_1 _2780_ (.B(_1128_),
    .C(_1101_),
    .A(_1115_),
    .Y(_1131_));
 sg13g2_nand3_1 _2781_ (.B(_1131_),
    .C(_2038_),
    .A(_1130_),
    .Y(_1132_));
 sg13g2_a21oi_1 _2782_ (.A1(_1132_),
    .A2(_2054_),
    .Y(_1133_),
    .B1(net52));
 sg13g2_nand2_1 _2783_ (.Y(_1134_),
    .A(_1077_),
    .B(_1133_));
 sg13g2_xnor2_1 _2784_ (.Y(_1135_),
    .A(net70),
    .B(_0167_));
 sg13g2_a21oi_1 _2785_ (.A1(_1135_),
    .A2(_0367_),
    .Y(_1136_),
    .B1(net46));
 sg13g2_nand2_1 _2786_ (.Y(_1137_),
    .A(_1134_),
    .B(_1136_));
 sg13g2_a21oi_1 _2787_ (.A1(_0256_),
    .A2(net46),
    .Y(_1138_),
    .B1(net37));
 sg13g2_nand2_1 _2788_ (.Y(_1139_),
    .A(_1137_),
    .B(_1138_));
 sg13g2_nand2_1 _2789_ (.Y(_1140_),
    .A(_1139_),
    .B(_0220_));
 sg13g2_nand2_1 _2790_ (.Y(_1141_),
    .A(_1140_),
    .B(_0225_));
 sg13g2_nand3_1 _2791_ (.B(_0300_),
    .C(net51),
    .A(_1141_),
    .Y(_1142_));
 sg13g2_inv_1 _2792_ (.Y(_1143_),
    .A(_1142_));
 sg13g2_inv_1 _2793_ (.Y(_1144_),
    .A(_1064_));
 sg13g2_nand2b_1 _2794_ (.Y(_1145_),
    .B(_1065_),
    .A_N(_1000_));
 sg13g2_inv_1 _2795_ (.Y(_1146_),
    .A(_1059_));
 sg13g2_a21oi_1 _2796_ (.A1(_1145_),
    .A2(_1146_),
    .Y(_1147_),
    .B1(_1002_));
 sg13g2_nand2_1 _2797_ (.Y(_1148_),
    .A(_1032_),
    .B(_1036_));
 sg13g2_nand2_1 _2798_ (.Y(_1149_),
    .A(_1148_),
    .B(_1041_));
 sg13g2_nor3_1 _2799_ (.A(_1144_),
    .B(_1147_),
    .C(_1149_),
    .Y(_1150_));
 sg13g2_a21oi_1 _2800_ (.A1(_1148_),
    .A2(_1012_),
    .Y(_1151_),
    .B1(_1042_));
 sg13g2_nor2b_1 _2801_ (.A(_1150_),
    .B_N(_1151_),
    .Y(_1152_));
 sg13g2_nand2b_1 _2802_ (.Y(_1153_),
    .B(_1059_),
    .A_N(_1051_));
 sg13g2_nand2_1 _2803_ (.Y(_1154_),
    .A(_1145_),
    .B(_1001_));
 sg13g2_nor2_1 _2804_ (.A(_1153_),
    .B(_1154_),
    .Y(_1155_));
 sg13g2_inv_1 _2805_ (.Y(_1156_),
    .A(_1058_));
 sg13g2_nand4_1 _2806_ (.B(_1155_),
    .C(_1156_),
    .A(_1038_),
    .Y(_1157_),
    .D(_1064_));
 sg13g2_nand2_1 _2807_ (.Y(_1158_),
    .A(_1152_),
    .B(_1157_));
 sg13g2_nand2_1 _2808_ (.Y(_1159_),
    .A(_1158_),
    .B(_1030_));
 sg13g2_inv_1 _2809_ (.Y(_1160_),
    .A(_1030_));
 sg13g2_nand3_1 _2810_ (.B(_1160_),
    .C(_1157_),
    .A(_1152_),
    .Y(_1161_));
 sg13g2_nand3_1 _2811_ (.B(_1161_),
    .C(net57),
    .A(_1159_),
    .Y(_1162_));
 sg13g2_a21oi_1 _2812_ (.A1(_1094_),
    .A2(_1096_),
    .Y(_1163_),
    .B1(_1082_));
 sg13g2_o21ai_1 _2813_ (.B1(_1086_),
    .Y(_1164_),
    .A1(_1083_),
    .A2(_1163_));
 sg13g2_xnor2_1 _2814_ (.Y(_1165_),
    .A(_1084_),
    .B(_1164_));
 sg13g2_xnor2_1 _2815_ (.Y(_1166_),
    .A(_1110_),
    .B(_1165_));
 sg13g2_nand3_1 _2816_ (.B(_1121_),
    .C(_1126_),
    .A(_1124_),
    .Y(_1167_));
 sg13g2_nand2_1 _2817_ (.Y(_1168_),
    .A(_1167_),
    .B(_1107_));
 sg13g2_nand2_1 _2818_ (.Y(_1169_),
    .A(_1168_),
    .B(_1102_));
 sg13g2_inv_1 _2819_ (.Y(_1170_),
    .A(_1112_));
 sg13g2_nand2_1 _2820_ (.Y(_1171_),
    .A(_1169_),
    .B(_1170_));
 sg13g2_xnor2_1 _2821_ (.Y(_1172_),
    .A(_1166_),
    .B(_1171_));
 sg13g2_a21oi_1 _2822_ (.A1(_1172_),
    .A2(net47),
    .Y(_1173_),
    .B1(_0355_));
 sg13g2_nor2_1 _2823_ (.A(net45),
    .B(_1173_),
    .Y(_1174_));
 sg13g2_nand2_1 _2824_ (.Y(_1175_),
    .A(_1162_),
    .B(_1174_));
 sg13g2_xnor2_1 _2825_ (.Y(_1176_),
    .A(net60),
    .B(_0396_));
 sg13g2_a21oi_1 _2826_ (.A1(_1176_),
    .A2(net45),
    .Y(_1177_),
    .B1(net46));
 sg13g2_nand2_1 _2827_ (.Y(_1178_),
    .A(_1175_),
    .B(_1177_));
 sg13g2_a21oi_1 _2828_ (.A1(_1937_),
    .A2(_0334_),
    .Y(_1179_),
    .B1(net37));
 sg13g2_nand2_1 _2829_ (.Y(_1180_),
    .A(_1178_),
    .B(_1179_));
 sg13g2_nand2_1 _2830_ (.Y(_1181_),
    .A(_1180_),
    .B(_0223_));
 sg13g2_nand2_2 _2831_ (.Y(_1182_),
    .A(_1181_),
    .B(_0227_));
 sg13g2_nand3_1 _2832_ (.B(net24),
    .C(net54),
    .A(_1182_),
    .Y(_1183_));
 sg13g2_nand2_1 _2833_ (.Y(_1184_),
    .A(_1183_),
    .B(net31));
 sg13g2_nor2_1 _2834_ (.A(_1143_),
    .B(_1184_),
    .Y(_1185_));
 sg13g2_a21oi_1 _2835_ (.A1(_1140_),
    .A2(_0225_),
    .Y(_1186_),
    .B1(_0301_));
 sg13g2_buf_8 _2836_ (.A(_1186_),
    .X(_1187_));
 sg13g2_xnor2_1 _2837_ (.Y(_1188_),
    .A(_1066_),
    .B(_1060_));
 sg13g2_xnor2_1 _2838_ (.Y(_1189_),
    .A(_1095_),
    .B(_1094_));
 sg13g2_xnor2_1 _2839_ (.Y(_1190_),
    .A(_1126_),
    .B(_1121_));
 sg13g2_xnor2_1 _2840_ (.Y(_1191_),
    .A(_1189_),
    .B(_1190_));
 sg13g2_a21oi_1 _2841_ (.A1(_1191_),
    .A2(net40),
    .Y(_1192_),
    .B1(_0471_));
 sg13g2_nor2_1 _2842_ (.A(net39),
    .B(_1192_),
    .Y(_1193_));
 sg13g2_o21ai_1 _2843_ (.B1(_1193_),
    .Y(_1194_),
    .A1(net50),
    .A2(_1188_));
 sg13g2_a21oi_1 _2844_ (.A1(_0397_),
    .A2(_1844_),
    .Y(_1195_),
    .B1(net43));
 sg13g2_o21ai_1 _2845_ (.B1(_1195_),
    .Y(_1196_),
    .A1(_1844_),
    .A2(net25));
 sg13g2_nand3_1 _2846_ (.B(net42),
    .C(_1196_),
    .A(_1194_),
    .Y(_1197_));
 sg13g2_nand2_1 _2847_ (.Y(_1198_),
    .A(net35),
    .B(_1983_));
 sg13g2_nand3_1 _2848_ (.B(_0174_),
    .C(_1198_),
    .A(_1197_),
    .Y(_1199_));
 sg13g2_a21oi_1 _2849_ (.A1(_1199_),
    .A2(_0220_),
    .Y(_1200_),
    .B1(net56));
 sg13g2_nor2b_1 _2850_ (.A(_1200_),
    .B_N(_0524_),
    .Y(_1201_));
 sg13g2_a21oi_1 _2851_ (.A1(_1187_),
    .A2(_0242_),
    .Y(_1202_),
    .B1(_1201_));
 sg13g2_nand2_1 _2852_ (.Y(_1203_),
    .A(_1185_),
    .B(_1202_));
 sg13g2_nand2_1 _2853_ (.Y(_1204_),
    .A(_1141_),
    .B(_0300_));
 sg13g2_nand3_1 _2854_ (.B(_0247_),
    .C(_1204_),
    .A(_1203_),
    .Y(_1205_));
 sg13g2_nand3_1 _2855_ (.B(_1187_),
    .C(_1202_),
    .A(_1185_),
    .Y(_1206_));
 sg13g2_nand2_1 _2856_ (.Y(_1207_),
    .A(_1205_),
    .B(_1206_));
 sg13g2_nand3_1 _2857_ (.B(_1103_),
    .C(_1107_),
    .A(_1167_),
    .Y(_1208_));
 sg13g2_nand2_1 _2858_ (.Y(_1209_),
    .A(_1169_),
    .B(_1208_));
 sg13g2_xor2_1 _2859_ (.B(_1163_),
    .A(_1083_),
    .X(_1210_));
 sg13g2_nand2_1 _2860_ (.Y(_1211_),
    .A(_1209_),
    .B(_1210_));
 sg13g2_inv_1 _2861_ (.Y(_1212_),
    .A(_1210_));
 sg13g2_nand3_1 _2862_ (.B(_1208_),
    .C(_1212_),
    .A(_1169_),
    .Y(_1213_));
 sg13g2_nand3_1 _2863_ (.B(_1213_),
    .C(net40),
    .A(_1211_),
    .Y(_1214_));
 sg13g2_nand2_1 _2864_ (.Y(_1215_),
    .A(_1214_),
    .B(_0829_));
 sg13g2_nand2_1 _2865_ (.Y(_1216_),
    .A(_1067_),
    .B(_1014_));
 sg13g2_nand2_1 _2866_ (.Y(_1217_),
    .A(_1216_),
    .B(_1038_));
 sg13g2_nand3_1 _2867_ (.B(_1014_),
    .C(_1149_),
    .A(_1067_),
    .Y(_1218_));
 sg13g2_nand3_1 _2868_ (.B(_1218_),
    .C(net57),
    .A(_1217_),
    .Y(_1219_));
 sg13g2_nand3_1 _2869_ (.B(net43),
    .C(_1219_),
    .A(_1215_),
    .Y(_1220_));
 sg13g2_xnor2_1 _2870_ (.Y(_1221_),
    .A(_1841_),
    .B(net29));
 sg13g2_a21oi_1 _2871_ (.A1(_1221_),
    .A2(net45),
    .Y(_1222_),
    .B1(net41));
 sg13g2_nand2_1 _2872_ (.Y(_1223_),
    .A(_1220_),
    .B(_1222_));
 sg13g2_a21oi_1 _2873_ (.A1(_1911_),
    .A2(net41),
    .Y(_1224_),
    .B1(net30));
 sg13g2_nand2_1 _2874_ (.Y(_1225_),
    .A(_1223_),
    .B(_1224_));
 sg13g2_nand2_1 _2875_ (.Y(_1226_),
    .A(_1225_),
    .B(_0223_));
 sg13g2_nand2_2 _2876_ (.Y(_1227_),
    .A(_1226_),
    .B(_0374_));
 sg13g2_nand3_1 _2877_ (.B(net24),
    .C(net54),
    .A(_1227_),
    .Y(_1228_));
 sg13g2_xor2_1 _2878_ (.B(_1091_),
    .A(_1090_),
    .X(_1229_));
 sg13g2_xor2_1 _2879_ (.B(_1117_),
    .A(_1118_),
    .X(_1230_));
 sg13g2_xnor2_1 _2880_ (.Y(_1231_),
    .A(_1229_),
    .B(_1230_));
 sg13g2_a21oi_1 _2881_ (.A1(_1231_),
    .A2(net40),
    .Y(_1232_),
    .B1(_0425_));
 sg13g2_o21ai_1 _2882_ (.B1(net57),
    .Y(_1233_),
    .A1(_1058_),
    .A2(_1153_));
 sg13g2_a21oi_1 _2883_ (.A1(_1153_),
    .A2(_1058_),
    .Y(_1234_),
    .B1(_1233_));
 sg13g2_nor3_1 _2884_ (.A(net39),
    .B(_1232_),
    .C(_1234_),
    .Y(_1235_));
 sg13g2_a21oi_1 _2885_ (.A1(net29),
    .A2(_0312_),
    .Y(_1236_),
    .B1(net43));
 sg13g2_o21ai_1 _2886_ (.B1(_1236_),
    .Y(_1237_),
    .A1(_0312_),
    .A2(net25));
 sg13g2_nand3b_1 _2887_ (.B(net42),
    .C(_1237_),
    .Y(_1238_),
    .A_N(_1235_));
 sg13g2_nand2_1 _2888_ (.Y(_1239_),
    .A(net35),
    .B(_1967_));
 sg13g2_nand3_1 _2889_ (.B(_0174_),
    .C(_1239_),
    .A(_1238_),
    .Y(_1240_));
 sg13g2_a21oi_1 _2890_ (.A1(_1240_),
    .A2(_0220_),
    .Y(_1241_),
    .B1(net56));
 sg13g2_nand2b_1 _2891_ (.Y(_1242_),
    .B(_0486_),
    .A_N(_1241_));
 sg13g2_nand2_1 _2892_ (.Y(_1243_),
    .A(_1228_),
    .B(_1242_));
 sg13g2_nand3_1 _2893_ (.B(net24),
    .C(net51),
    .A(_1182_),
    .Y(_1244_));
 sg13g2_nand2_1 _2894_ (.Y(_1245_),
    .A(_1244_),
    .B(net31));
 sg13g2_nor2_1 _2895_ (.A(_1243_),
    .B(_1245_),
    .Y(_1246_));
 sg13g2_a22oi_1 _2896_ (.Y(_1247_),
    .B1(_0343_),
    .B2(_1187_),
    .A2(_1182_),
    .A1(net23));
 sg13g2_nand2_1 _2897_ (.Y(_1248_),
    .A(_1246_),
    .B(_1247_));
 sg13g2_nor2_2 _2898_ (.A(net31),
    .B(_1187_),
    .Y(_1249_));
 sg13g2_inv_8 _2899_ (.Y(_1250_),
    .A(_1249_));
 sg13g2_nand2_1 _2900_ (.Y(_1251_),
    .A(_0420_),
    .B(_0806_));
 sg13g2_inv_1 _2901_ (.Y(_1252_),
    .A(_1251_));
 sg13g2_nand2_1 _2902_ (.Y(_1253_),
    .A(_1182_),
    .B(net24));
 sg13g2_a21oi_1 _2903_ (.A1(_0408_),
    .A2(_1252_),
    .Y(_1254_),
    .B1(_1253_));
 sg13g2_nand3_1 _2904_ (.B(net24),
    .C(_0417_),
    .A(_1182_),
    .Y(_1255_));
 sg13g2_nand2_1 _2905_ (.Y(_1256_),
    .A(_1255_),
    .B(net31));
 sg13g2_nor2_1 _2906_ (.A(_1254_),
    .B(_1256_),
    .Y(_1257_));
 sg13g2_nand3_1 _2907_ (.B(_1250_),
    .C(_1257_),
    .A(_1248_),
    .Y(_1258_));
 sg13g2_nor2_1 _2908_ (.A(_1249_),
    .B(_1257_),
    .Y(_1259_));
 sg13g2_nand2b_1 _2909_ (.Y(_1260_),
    .B(_1259_),
    .A_N(_1248_));
 sg13g2_nand2_1 _2910_ (.Y(_1261_),
    .A(_1258_),
    .B(_1260_));
 sg13g2_nor2_1 _2911_ (.A(_1207_),
    .B(_1261_),
    .Y(_1262_));
 sg13g2_nand3_1 _2912_ (.B(net24),
    .C(_0493_),
    .A(_1227_),
    .Y(_1263_));
 sg13g2_nand2_1 _2913_ (.Y(_1264_),
    .A(_1227_),
    .B(net23));
 sg13g2_nand3_1 _2914_ (.B(net31),
    .C(_1264_),
    .A(_1263_),
    .Y(_1265_));
 sg13g2_nor2b_1 _2915_ (.A(_1265_),
    .B_N(_1142_),
    .Y(_1266_));
 sg13g2_nor2b_1 _2916_ (.A(_1266_),
    .B_N(_1250_),
    .Y(_1267_));
 sg13g2_nor2_1 _2917_ (.A(_0800_),
    .B(_1204_),
    .Y(_1268_));
 sg13g2_nor2_1 _2918_ (.A(_0056_),
    .B(net42),
    .Y(_1269_));
 sg13g2_a21oi_1 _2919_ (.A1(_1055_),
    .A2(_0053_),
    .Y(_1270_),
    .B1(net50));
 sg13g2_o21ai_1 _2920_ (.B1(_1270_),
    .Y(_1271_),
    .A1(_0053_),
    .A2(_1055_));
 sg13g2_nand2_1 _2921_ (.Y(_1272_),
    .A(net25),
    .B(_1847_));
 sg13g2_a21oi_1 _2922_ (.A1(net27),
    .A2(\i_project.controller_0.mode_ramp_base[0] ),
    .Y(_1273_),
    .B1(net36));
 sg13g2_a22oi_1 _2923_ (.Y(_1274_),
    .B1(_1272_),
    .B2(_1273_),
    .A2(_1271_),
    .A1(net36));
 sg13g2_nor2_1 _2924_ (.A(_1269_),
    .B(_1274_),
    .Y(_1275_));
 sg13g2_nand2_1 _2925_ (.Y(_1276_),
    .A(_1275_),
    .B(_0174_));
 sg13g2_nand2_1 _2926_ (.Y(_1277_),
    .A(_1094_),
    .B(_1095_));
 sg13g2_nand2_1 _2927_ (.Y(_1278_),
    .A(_1277_),
    .B(_1079_));
 sg13g2_xnor2_1 _2928_ (.Y(_1279_),
    .A(_1080_),
    .B(_1278_));
 sg13g2_a21oi_1 _2929_ (.A1(_1121_),
    .A2(_1126_),
    .Y(_1280_),
    .B1(_1105_));
 sg13g2_xnor2_1 _2930_ (.Y(_1281_),
    .A(_1124_),
    .B(_1280_));
 sg13g2_xor2_1 _2931_ (.B(_1281_),
    .A(_1279_),
    .X(_1282_));
 sg13g2_o21ai_1 _2932_ (.B1(_0855_),
    .Y(_1283_),
    .A1(_0316_),
    .A2(_1282_));
 sg13g2_a21oi_1 _2933_ (.A1(_1060_),
    .A2(_1145_),
    .Y(_1284_),
    .B1(_1002_));
 sg13g2_xnor2_1 _2934_ (.Y(_1285_),
    .A(_1064_),
    .B(_1284_));
 sg13g2_nand2_1 _2935_ (.Y(_1286_),
    .A(_1285_),
    .B(net49));
 sg13g2_nand3_1 _2936_ (.B(_1286_),
    .C(net43),
    .A(_1283_),
    .Y(_1287_));
 sg13g2_xnor2_1 _2937_ (.Y(_1288_),
    .A(net61),
    .B(net29));
 sg13g2_a21oi_1 _2938_ (.A1(_1288_),
    .A2(net39),
    .Y(_1289_),
    .B1(net41));
 sg13g2_nand2_1 _2939_ (.Y(_1290_),
    .A(_1287_),
    .B(_1289_));
 sg13g2_a21oi_1 _2940_ (.A1(_1986_),
    .A2(net41),
    .Y(_1291_),
    .B1(net30));
 sg13g2_nand2_1 _2941_ (.Y(_1292_),
    .A(_1290_),
    .B(_1291_));
 sg13g2_nand2_1 _2942_ (.Y(_1293_),
    .A(_1292_),
    .B(_0223_));
 sg13g2_nand2_1 _2943_ (.Y(_1294_),
    .A(_1293_),
    .B(_0406_));
 sg13g2_a22oi_1 _2944_ (.Y(_1295_),
    .B1(net23),
    .B2(_1294_),
    .A2(_1276_),
    .A1(_0341_));
 sg13g2_nand3_1 _2945_ (.B(net24),
    .C(_0343_),
    .A(_1227_),
    .Y(_1296_));
 sg13g2_nand2_1 _2946_ (.Y(_1297_),
    .A(_1295_),
    .B(_1296_));
 sg13g2_nor3_1 _2947_ (.A(_1268_),
    .B(_1297_),
    .C(_1256_),
    .Y(_1298_));
 sg13g2_and2_1 _2948_ (.A(_1294_),
    .B(_0450_),
    .X(_1299_));
 sg13g2_a21oi_1 _2949_ (.A1(_1187_),
    .A2(net54),
    .Y(_1300_),
    .B1(_1299_));
 sg13g2_inv_2 _2950_ (.Y(_1301_),
    .A(_1245_));
 sg13g2_nand2_1 _2951_ (.Y(_1302_),
    .A(_1300_),
    .B(_1301_));
 sg13g2_nand3_1 _2952_ (.B(_1298_),
    .C(_1302_),
    .A(_1267_),
    .Y(_1303_));
 sg13g2_nor2_1 _2953_ (.A(_0806_),
    .B(_1253_),
    .Y(_1304_));
 sg13g2_a21oi_1 _2954_ (.A1(_1227_),
    .A2(net23),
    .Y(_1305_),
    .B1(_0245_));
 sg13g2_o21ai_1 _2955_ (.B1(net39),
    .Y(_1306_),
    .A1(_1845_),
    .A2(net27));
 sg13g2_a21oi_1 _2956_ (.A1(_1845_),
    .A2(net27),
    .Y(_1307_),
    .B1(_1306_));
 sg13g2_nor2b_1 _2957_ (.A(_1057_),
    .B_N(_1054_),
    .Y(_1308_));
 sg13g2_xnor2_1 _2958_ (.Y(_1309_),
    .A(_1056_),
    .B(_1308_));
 sg13g2_nand2_1 _2959_ (.Y(_1310_),
    .A(_1309_),
    .B(net49));
 sg13g2_a21oi_1 _2960_ (.A1(_1310_),
    .A2(_0324_),
    .Y(_1311_),
    .B1(net39));
 sg13g2_nor3_1 _2961_ (.A(net35),
    .B(_1307_),
    .C(_1311_),
    .Y(_1312_));
 sg13g2_o21ai_1 _2962_ (.B1(_0174_),
    .Y(_1313_),
    .A1(_0021_),
    .A2(net42));
 sg13g2_o21ai_1 _2963_ (.B1(_0422_),
    .Y(_1314_),
    .A1(_1312_),
    .A2(_1313_));
 sg13g2_nand2_1 _2964_ (.Y(_1315_),
    .A(_1305_),
    .B(_1314_));
 sg13g2_o21ai_1 _2965_ (.B1(_1250_),
    .Y(_1316_),
    .A1(_1304_),
    .A2(_1315_));
 sg13g2_o21ai_1 _2966_ (.B1(_1316_),
    .Y(_1317_),
    .A1(_0416_),
    .A2(_1204_));
 sg13g2_nand2_1 _2967_ (.Y(_1318_),
    .A(_1303_),
    .B(_1317_));
 sg13g2_a21oi_2 _2968_ (.B1(_1249_),
    .Y(_1319_),
    .A2(_1301_),
    .A1(_1300_));
 sg13g2_nand2_1 _2969_ (.Y(_1320_),
    .A(_1319_),
    .B(_1298_));
 sg13g2_inv_1 _2970_ (.Y(_1321_),
    .A(_1267_));
 sg13g2_nand2_1 _2971_ (.Y(_1322_),
    .A(_1320_),
    .B(_1321_));
 sg13g2_nand2_1 _2972_ (.Y(_1323_),
    .A(_1318_),
    .B(_1322_));
 sg13g2_nand2_2 _2973_ (.Y(_1324_),
    .A(_1262_),
    .B(_1323_));
 sg13g2_inv_1 _2974_ (.Y(_1325_),
    .A(_1258_));
 sg13g2_inv_1 _2975_ (.Y(_1326_),
    .A(_1205_));
 sg13g2_a21oi_2 _2976_ (.B1(_1326_),
    .Y(_1327_),
    .A2(_1206_),
    .A1(_1325_));
 sg13g2_nand2_1 _2977_ (.Y(_1328_),
    .A(_1324_),
    .B(_1327_));
 sg13g2_inv_2 _2978_ (.Y(_1329_),
    .A(_1319_));
 sg13g2_nand2_1 _2979_ (.Y(_1330_),
    .A(_1328_),
    .B(_1329_));
 sg13g2_nand3_1 _2980_ (.B(_1319_),
    .C(_1327_),
    .A(_1324_),
    .Y(_1331_));
 sg13g2_nand2_1 _2981_ (.Y(_1332_),
    .A(_1330_),
    .B(_1331_));
 sg13g2_inv_1 _2982_ (.Y(_1333_),
    .A(_1259_));
 sg13g2_nand2_1 _2983_ (.Y(_1334_),
    .A(_1328_),
    .B(_1333_));
 sg13g2_nand2_1 _2984_ (.Y(_1335_),
    .A(_1329_),
    .B(_1321_));
 sg13g2_xnor2_1 _2985_ (.Y(_1336_),
    .A(_1333_),
    .B(_1335_));
 sg13g2_nand3_1 _2986_ (.B(_1327_),
    .C(_1336_),
    .A(_1324_),
    .Y(_1337_));
 sg13g2_nand2_1 _2987_ (.Y(_1338_),
    .A(_1334_),
    .B(_1337_));
 sg13g2_nand2_1 _2988_ (.Y(_1339_),
    .A(_1248_),
    .B(_1250_));
 sg13g2_nand2_1 _2989_ (.Y(_1340_),
    .A(_1338_),
    .B(_1339_));
 sg13g2_inv_1 _2990_ (.Y(_1341_),
    .A(_1339_));
 sg13g2_nand3_1 _2991_ (.B(_1337_),
    .C(_1341_),
    .A(_1334_),
    .Y(_1342_));
 sg13g2_nand2_1 _2992_ (.Y(_1343_),
    .A(_1340_),
    .B(_1342_));
 sg13g2_nand2_1 _2993_ (.Y(_1344_),
    .A(_1328_),
    .B(_1267_));
 sg13g2_o21ai_1 _2994_ (.B1(_1335_),
    .Y(_1345_),
    .A1(_1329_),
    .A2(_1266_));
 sg13g2_nand3_1 _2995_ (.B(_1327_),
    .C(_1345_),
    .A(_1324_),
    .Y(_1346_));
 sg13g2_nand2_1 _2996_ (.Y(_1347_),
    .A(_1344_),
    .B(_1346_));
 sg13g2_buf_8 _2997_ (.A(_1347_),
    .X(_1348_));
 sg13g2_nand2_1 _2998_ (.Y(_1349_),
    .A(_1348_),
    .B(_1317_));
 sg13g2_inv_1 _2999_ (.Y(_1350_),
    .A(_1317_));
 sg13g2_nand3_1 _3000_ (.B(_1346_),
    .C(_1350_),
    .A(_1344_),
    .Y(_1351_));
 sg13g2_nand2_1 _3001_ (.Y(_1352_),
    .A(_1349_),
    .B(_1351_));
 sg13g2_nor2_1 _3002_ (.A(_1249_),
    .B(_1298_),
    .Y(_1353_));
 sg13g2_inv_1 _3003_ (.Y(_1354_),
    .A(_1353_));
 sg13g2_nand3_1 _3004_ (.B(_1331_),
    .C(_1354_),
    .A(_1330_),
    .Y(_1355_));
 sg13g2_buf_2 _3005_ (.A(_1355_),
    .X(_1356_));
 sg13g2_nand3_1 _3006_ (.B(_1352_),
    .C(_1356_),
    .A(_1343_),
    .Y(_1357_));
 sg13g2_inv_2 _3007_ (.Y(_1358_),
    .A(_1338_));
 sg13g2_nand2_1 _3008_ (.Y(_1359_),
    .A(_1358_),
    .B(_1339_));
 sg13g2_nor2_1 _3009_ (.A(_1350_),
    .B(_1348_),
    .Y(_1360_));
 sg13g2_nor2_1 _3010_ (.A(_1339_),
    .B(_1358_),
    .Y(_1361_));
 sg13g2_a21oi_1 _3011_ (.A1(_1359_),
    .A2(_1360_),
    .Y(_1362_),
    .B1(_1361_));
 sg13g2_nand2_1 _3012_ (.Y(_1363_),
    .A(_1357_),
    .B(_1362_));
 sg13g2_nand2_1 _3013_ (.Y(_1364_),
    .A(_1328_),
    .B(_1187_));
 sg13g2_nor2_1 _3014_ (.A(_1259_),
    .B(_1267_),
    .Y(_1365_));
 sg13g2_nand2_1 _3015_ (.Y(_1366_),
    .A(_1365_),
    .B(_1329_));
 sg13g2_xnor2_1 _3016_ (.Y(_1367_),
    .A(_1187_),
    .B(_1366_));
 sg13g2_nand3_1 _3017_ (.B(_1327_),
    .C(_1367_),
    .A(_1324_),
    .Y(_1368_));
 sg13g2_nand2_1 _3018_ (.Y(_1369_),
    .A(_1203_),
    .B(_1250_));
 sg13g2_nand3_1 _3019_ (.B(_1368_),
    .C(_1369_),
    .A(_1364_),
    .Y(_1370_));
 sg13g2_nand3_1 _3020_ (.B(_1187_),
    .C(_1250_),
    .A(_1203_),
    .Y(_1371_));
 sg13g2_nand2_1 _3021_ (.Y(_1372_),
    .A(_1370_),
    .B(_1371_));
 sg13g2_inv_1 _3022_ (.Y(_1373_),
    .A(_1372_));
 sg13g2_nand2_1 _3023_ (.Y(_1374_),
    .A(_1363_),
    .B(_1373_));
 sg13g2_nand3_1 _3024_ (.B(_1362_),
    .C(_1372_),
    .A(_1357_),
    .Y(_1375_));
 sg13g2_nand3_1 _3025_ (.B(_1375_),
    .C(_1698_),
    .A(_1374_),
    .Y(_1376_));
 sg13g2_nand2_1 _3026_ (.Y(_1377_),
    .A(_1363_),
    .B(_1372_));
 sg13g2_nand3_1 _3027_ (.B(_1362_),
    .C(_1373_),
    .A(_1357_),
    .Y(_1378_));
 sg13g2_nand3_1 _3028_ (.B(_1378_),
    .C(_0581_),
    .A(_1377_),
    .Y(_1379_));
 sg13g2_nand2_1 _3029_ (.Y(_1380_),
    .A(_1376_),
    .B(_1379_));
 sg13g2_nand2_1 _3030_ (.Y(_1381_),
    .A(_1343_),
    .B(_1372_));
 sg13g2_nand2_1 _3031_ (.Y(_1382_),
    .A(_1348_),
    .B(_1350_));
 sg13g2_a21oi_1 _3032_ (.A1(_1382_),
    .A2(_1356_),
    .Y(_1383_),
    .B1(_1360_));
 sg13g2_nor2_1 _3033_ (.A(_1381_),
    .B(_1383_),
    .Y(_1384_));
 sg13g2_nand3_1 _3034_ (.B(_1324_),
    .C(_1327_),
    .A(_1384_),
    .Y(_1385_));
 sg13g2_xnor2_1 _3035_ (.Y(_1386_),
    .A(_1667_),
    .B(_1385_));
 sg13g2_nand3b_1 _3036_ (.B(_1349_),
    .C(_1351_),
    .Y(_1387_),
    .A_N(_1356_));
 sg13g2_nand2_1 _3037_ (.Y(_1388_),
    .A(_1352_),
    .B(_1356_));
 sg13g2_nand2_1 _3038_ (.Y(_1389_),
    .A(_1387_),
    .B(_1388_));
 sg13g2_nand2b_1 _3039_ (.Y(_1390_),
    .B(_1389_),
    .A_N(_0018_));
 sg13g2_nand3_1 _3040_ (.B(_1388_),
    .C(_0018_),
    .A(_1387_),
    .Y(_1391_));
 sg13g2_nand2_1 _3041_ (.Y(_1392_),
    .A(_1332_),
    .B(_1353_));
 sg13g2_nand3_1 _3042_ (.B(_1356_),
    .C(_1668_),
    .A(_1392_),
    .Y(_1393_));
 sg13g2_nand3_1 _3043_ (.B(_1391_),
    .C(_1393_),
    .A(_1390_),
    .Y(_1394_));
 sg13g2_inv_1 _3044_ (.Y(_1395_),
    .A(_1343_));
 sg13g2_xnor2_1 _3045_ (.Y(_1396_),
    .A(_1395_),
    .B(_1383_));
 sg13g2_xnor2_1 _3046_ (.Y(_1397_),
    .A(_1665_),
    .B(_1396_));
 sg13g2_nor2_1 _3047_ (.A(_1394_),
    .B(_1397_),
    .Y(_1398_));
 sg13g2_nand3_1 _3048_ (.B(_1386_),
    .C(_1398_),
    .A(_1380_),
    .Y(_1399_));
 sg13g2_a21oi_1 _3049_ (.A1(_1374_),
    .A2(_1375_),
    .Y(_1400_),
    .B1(_1657_));
 sg13g2_nor2_1 _3050_ (.A(\dither_threshold[4] ),
    .B(_1385_),
    .Y(_1401_));
 sg13g2_a21oi_1 _3051_ (.A1(_1386_),
    .A2(_1400_),
    .Y(_1402_),
    .B1(_1401_));
 sg13g2_nand2_1 _3052_ (.Y(_1403_),
    .A(_1399_),
    .B(_1402_));
 sg13g2_nand3_1 _3053_ (.B(_1375_),
    .C(_0581_),
    .A(_1374_),
    .Y(_1404_));
 sg13g2_nand3_1 _3054_ (.B(_1378_),
    .C(_1698_),
    .A(_1377_),
    .Y(_1405_));
 sg13g2_nand2_1 _3055_ (.Y(_1406_),
    .A(_1404_),
    .B(_1405_));
 sg13g2_nor2b_1 _3056_ (.A(_1406_),
    .B_N(_1386_),
    .Y(_1407_));
 sg13g2_xnor2_1 _3057_ (.Y(_1408_),
    .A(_1664_),
    .B(_1396_));
 sg13g2_nor2_1 _3058_ (.A(_1661_),
    .B(_1389_),
    .Y(_1409_));
 sg13g2_nand2_1 _3059_ (.Y(_1410_),
    .A(_1408_),
    .B(_1409_));
 sg13g2_nand2b_1 _3060_ (.Y(_1411_),
    .B(_1695_),
    .A_N(_1396_));
 sg13g2_nand2_1 _3061_ (.Y(_1412_),
    .A(_1410_),
    .B(_1411_));
 sg13g2_nand2_1 _3062_ (.Y(_1413_),
    .A(_1407_),
    .B(_1412_));
 sg13g2_nor2b_1 _3063_ (.A(_1403_),
    .B_N(_1413_),
    .Y(_1414_));
 sg13g2_a21o_1 _3064_ (.A2(_1356_),
    .A1(_1392_),
    .B1(_1668_),
    .X(_1415_));
 sg13g2_nand3_1 _3065_ (.B(_1398_),
    .C(_1415_),
    .A(_1407_),
    .Y(_1416_));
 sg13g2_nor2b_1 _3066_ (.A(_1414_),
    .B_N(_1416_),
    .Y(_1417_));
 sg13g2_xnor2_1 _3067_ (.Y(net18),
    .A(_1332_),
    .B(_1417_));
 sg13g2_inv_1 _3068_ (.Y(_1418_),
    .A(_1332_));
 sg13g2_nand2_1 _3069_ (.Y(_1419_),
    .A(_1417_),
    .B(_1418_));
 sg13g2_xnor2_1 _3070_ (.Y(net19),
    .A(_1348_),
    .B(_1419_));
 sg13g2_nand4_1 _3071_ (.B(_1418_),
    .C(_1338_),
    .A(_1417_),
    .Y(_1420_),
    .D(_1348_));
 sg13g2_nand3_1 _3072_ (.B(_1399_),
    .C(_1402_),
    .A(_1413_),
    .Y(_1421_));
 sg13g2_nand4_1 _3073_ (.B(_1418_),
    .C(_1348_),
    .A(_1421_),
    .Y(_1422_),
    .D(_1416_));
 sg13g2_nand2_1 _3074_ (.Y(_1423_),
    .A(_1422_),
    .B(_1358_));
 sg13g2_nand2_1 _3075_ (.Y(net20),
    .A(_1420_),
    .B(_1423_));
 sg13g2_nand2_1 _3076_ (.Y(_1424_),
    .A(_1364_),
    .B(_1368_));
 sg13g2_nand4_1 _3077_ (.B(_1418_),
    .C(_1358_),
    .A(_1417_),
    .Y(_1425_),
    .D(_1348_));
 sg13g2_nand2b_1 _3078_ (.Y(net21),
    .B(_1425_),
    .A_N(_1424_));
 sg13g2_nor4_1 _3079_ (.A(\counter[21] ),
    .B(\counter[20] ),
    .C(\counter[23] ),
    .D(\counter[22] ),
    .Y(_1426_));
 sg13g2_nor4_1 _3080_ (.A(\counter[17] ),
    .B(\counter[16] ),
    .C(\counter[19] ),
    .D(\counter[18] ),
    .Y(_1427_));
 sg13g2_nor3_1 _3081_ (.A(\counter[25] ),
    .B(\counter[24] ),
    .C(\counter[26] ),
    .Y(_1428_));
 sg13g2_and3_1 _3082_ (.X(_1429_),
    .A(_1426_),
    .B(_1427_),
    .C(_1428_));
 sg13g2_inv_1 _3083_ (.Y(_1430_),
    .A(\counter[4] ));
 sg13g2_inv_1 _3084_ (.Y(_1431_),
    .A(\counter[7] ));
 sg13g2_nand2_1 _3085_ (.Y(_1432_),
    .A(_1430_),
    .B(_1431_));
 sg13g2_nor2_1 _3086_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .Y(_1433_));
 sg13g2_inv_1 _3087_ (.Y(_1434_),
    .A(\counter[2] ));
 sg13g2_nand3b_1 _3088_ (.B(_1433_),
    .C(_1434_),
    .Y(_1435_),
    .A_N(\counter[3] ));
 sg13g2_nor4_1 _3089_ (.A(\counter[5] ),
    .B(\counter[6] ),
    .C(_1432_),
    .D(_1435_),
    .Y(_1436_));
 sg13g2_nor4_1 _3090_ (.A(\counter[13] ),
    .B(\counter[12] ),
    .C(\counter[15] ),
    .D(\counter[14] ),
    .Y(_1437_));
 sg13g2_nor4_1 _3091_ (.A(\counter[9] ),
    .B(\counter[8] ),
    .C(\counter[11] ),
    .D(\counter[10] ),
    .Y(_1438_));
 sg13g2_nand4_1 _3092_ (.B(_1436_),
    .C(_1437_),
    .A(_1429_),
    .Y(_0008_),
    .D(_1438_));
 sg13g2_inv_1 _3093_ (.Y(_1439_),
    .A(\counter[21] ));
 sg13g2_inv_1 _3094_ (.Y(_1440_),
    .A(\counter[19] ));
 sg13g2_nand2_1 _3095_ (.Y(_1441_),
    .A(\counter[17] ),
    .B(\counter[18] ));
 sg13g2_inv_1 _3096_ (.Y(_1442_),
    .A(\counter[11] ));
 sg13g2_inv_1 _3097_ (.Y(_1443_),
    .A(\counter[10] ));
 sg13g2_inv_1 _3098_ (.Y(_1444_),
    .A(\counter[9] ));
 sg13g2_inv_1 _3099_ (.Y(_1445_),
    .A(\counter[8] ));
 sg13g2_nand2_1 _3100_ (.Y(_1446_),
    .A(\counter[1] ),
    .B(\counter[0] ));
 sg13g2_nor2_1 _3101_ (.A(_1434_),
    .B(_1446_),
    .Y(_1447_));
 sg13g2_nand2_1 _3102_ (.Y(_1448_),
    .A(_1447_),
    .B(\counter[3] ));
 sg13g2_inv_1 _3103_ (.Y(_1449_),
    .A(_1448_));
 sg13g2_inv_1 _3104_ (.Y(_1450_),
    .A(\counter[6] ));
 sg13g2_nand2_1 _3105_ (.Y(_1451_),
    .A(\counter[5] ),
    .B(\counter[4] ));
 sg13g2_nor3_1 _3106_ (.A(_1431_),
    .B(_1450_),
    .C(_1451_),
    .Y(_1452_));
 sg13g2_nand2_1 _3107_ (.Y(_1453_),
    .A(_1449_),
    .B(_1452_));
 sg13g2_nor2_1 _3108_ (.A(_1445_),
    .B(_1453_),
    .Y(_1454_));
 sg13g2_inv_1 _3109_ (.Y(_1455_),
    .A(_1454_));
 sg13g2_nor2_1 _3110_ (.A(_1444_),
    .B(_1455_),
    .Y(_1456_));
 sg13g2_inv_1 _3111_ (.Y(_1457_),
    .A(_1456_));
 sg13g2_nor3_1 _3112_ (.A(_1442_),
    .B(_1443_),
    .C(_1457_),
    .Y(_1458_));
 sg13g2_nand2_1 _3113_ (.Y(_1459_),
    .A(_1458_),
    .B(\counter[12] ));
 sg13g2_nor2b_1 _3114_ (.A(_1459_),
    .B_N(\counter[13] ),
    .Y(_1460_));
 sg13g2_nand2_1 _3115_ (.Y(_1461_),
    .A(_1460_),
    .B(\counter[14] ));
 sg13g2_nor2b_1 _3116_ (.A(_1461_),
    .B_N(\counter[15] ),
    .Y(_1462_));
 sg13g2_nand2_1 _3117_ (.Y(_1463_),
    .A(_1462_),
    .B(\counter[16] ));
 sg13g2_nor3_1 _3118_ (.A(_1440_),
    .B(_1441_),
    .C(_1463_),
    .Y(_1464_));
 sg13g2_nand2_1 _3119_ (.Y(_1465_),
    .A(_1464_),
    .B(\counter[20] ));
 sg13g2_nor2_2 _3120_ (.A(_1439_),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_inv_1 _3121_ (.Y(_1467_),
    .A(\counter[25] ));
 sg13g2_inv_1 _3122_ (.Y(_1468_),
    .A(\counter[24] ));
 sg13g2_nand2_1 _3123_ (.Y(_1469_),
    .A(\counter[23] ),
    .B(\counter[22] ));
 sg13g2_nor3_1 _3124_ (.A(_1467_),
    .B(_1468_),
    .C(_1469_),
    .Y(_1470_));
 sg13g2_and3_1 _3125_ (.X(_1471_),
    .A(_1466_),
    .B(\counter[26] ),
    .C(_1470_));
 sg13g2_buf_1 _3126_ (.A(_1471_),
    .X(_1472_));
 sg13g2_nand2_1 _3127_ (.Y(_1473_),
    .A(\counter[27] ),
    .B(\counter[28] ));
 sg13g2_inv_1 _3128_ (.Y(_1474_),
    .A(_1473_));
 sg13g2_nand2_1 _3129_ (.Y(_1475_),
    .A(_1472_),
    .B(\counter[27] ));
 sg13g2_inv_1 _3130_ (.Y(_1476_),
    .A(\counter[28] ));
 sg13g2_buf_1 _3131_ (.A(rst_n),
    .X(_1477_));
 sg13g2_inv_1 _3132_ (.Y(_1478_),
    .A(_1477_));
 sg13g2_a221oi_1 _3133_ (.B2(_1476_),
    .C1(net82),
    .B1(_1475_),
    .A1(_1472_),
    .Y(_1479_),
    .A2(_1474_));
 sg13g2_buf_1 _3134_ (.A(_1479_),
    .X(_0078_));
 sg13g2_inv_2 _3135_ (.Y(_1480_),
    .A(_1463_));
 sg13g2_inv_1 _3136_ (.Y(_1481_),
    .A(\counter[23] ));
 sg13g2_inv_1 _3137_ (.Y(_1482_),
    .A(\counter[26] ));
 sg13g2_nor4_1 _3138_ (.A(_1481_),
    .B(_1467_),
    .C(_1468_),
    .D(_1482_),
    .Y(_1483_));
 sg13g2_inv_1 _3139_ (.Y(_1484_),
    .A(\counter[22] ));
 sg13g2_nand2_1 _3140_ (.Y(_1485_),
    .A(\counter[21] ),
    .B(\counter[20] ));
 sg13g2_nor4_2 _3141_ (.A(_1440_),
    .B(_1484_),
    .C(_1441_),
    .Y(_1486_),
    .D(_1485_));
 sg13g2_and3_1 _3142_ (.X(_1487_),
    .A(_1480_),
    .B(_1483_),
    .C(_1486_));
 sg13g2_nor2_1 _3143_ (.A(\counter[27] ),
    .B(_1487_),
    .Y(_1488_));
 sg13g2_inv_1 _3144_ (.Y(_1489_),
    .A(_1487_));
 sg13g2_nor2b_1 _3145_ (.A(_1489_),
    .B_N(\counter[27] ),
    .Y(_1490_));
 sg13g2_nor3_1 _3146_ (.A(net82),
    .B(_1488_),
    .C(_1490_),
    .Y(_0077_));
 sg13g2_inv_1 _3147_ (.Y(_1491_),
    .A(_0077_));
 sg13g2_nand2_1 _3148_ (.Y(_1492_),
    .A(_0078_),
    .B(_1491_));
 sg13g2_inv_1 _3149_ (.Y(_1493_),
    .A(\counter[29] ));
 sg13g2_nor3_1 _3150_ (.A(_1493_),
    .B(_1473_),
    .C(_1489_),
    .Y(_1494_));
 sg13g2_a21oi_1 _3151_ (.A1(_1490_),
    .A2(\counter[28] ),
    .Y(_1495_),
    .B1(\counter[29] ));
 sg13g2_nor3_2 _3152_ (.A(net82),
    .B(_1494_),
    .C(_1495_),
    .Y(_0079_));
 sg13g2_nor2_1 _3153_ (.A(_1491_),
    .B(_0078_),
    .Y(_1496_));
 sg13g2_a21oi_1 _3154_ (.A1(_1492_),
    .A2(_0079_),
    .Y(_0000_),
    .B1(_1496_));
 sg13g2_inv_1 _3155_ (.Y(_1497_),
    .A(_0079_));
 sg13g2_o21ai_1 _3156_ (.B1(_1492_),
    .Y(_0001_),
    .A1(_1497_),
    .A2(_1496_));
 sg13g2_a21o_1 _3157_ (.A2(_0079_),
    .A1(_0078_),
    .B1(_0077_),
    .X(_0002_));
 sg13g2_buf_1 _3158_ (.A(\i_project.controller_0.rst_n ),
    .X(_1498_));
 sg13g2_buf_1 _3159_ (.A(_1498_),
    .X(_1499_));
 sg13g2_buf_2 _3160_ (.A(\i_project.controller_0.divider[0] ),
    .X(_1500_));
 sg13g2_inv_1 _3161_ (.Y(_1501_),
    .A(_1500_));
 sg13g2_nor2_1 _3162_ (.A(_1498_),
    .B(\i_project.controller_0.grey_pass[10] ),
    .Y(_1502_));
 sg13g2_a21oi_1 _3163_ (.A1(net69),
    .A2(_1501_),
    .Y(_0003_),
    .B1(_1502_));
 sg13g2_buf_1 _3164_ (.A(\i_project.controller_0.divider[1] ),
    .X(_1503_));
 sg13g2_inv_1 _3165_ (.Y(_1504_),
    .A(_1503_));
 sg13g2_nor2_1 _3166_ (.A(net69),
    .B(\i_project.controller_0.grey_pass[11] ),
    .Y(_1505_));
 sg13g2_a21oi_1 _3167_ (.A1(net69),
    .A2(_1504_),
    .Y(_0004_),
    .B1(_1505_));
 sg13g2_buf_1 _3168_ (.A(ui_in[7]),
    .X(_1506_));
 sg13g2_mux2_1 _3169_ (.A0(_0012_),
    .A1(net1),
    .S(net83),
    .X(_0009_));
 sg13g2_mux2_1 _3170_ (.A0(_0013_),
    .A1(net2),
    .S(net83),
    .X(_0010_));
 sg13g2_mux2_1 _3171_ (.A0(_0014_),
    .A1(net3),
    .S(net83),
    .X(_0011_));
 sg13g2_nand2_1 _3172_ (.Y(_1507_),
    .A(net83),
    .B(net5));
 sg13g2_o21ai_1 _3173_ (.B1(_1507_),
    .Y(_0005_),
    .A1(net83),
    .A2(_1468_));
 sg13g2_nand2_1 _3174_ (.Y(_1508_),
    .A(_1506_),
    .B(net6));
 sg13g2_o21ai_1 _3175_ (.B1(_1508_),
    .Y(_0006_),
    .A1(net83),
    .A2(_1467_));
 sg13g2_nand2_1 _3176_ (.Y(_1509_),
    .A(_1506_),
    .B(net7));
 sg13g2_o21ai_1 _3177_ (.B1(_1509_),
    .Y(_0007_),
    .A1(net83),
    .A2(_1482_));
 sg13g2_buf_2 _3178_ (.A(\i_project.controller_0.vga_sync.mode ),
    .X(_1510_));
 sg13g2_inv_2 _3179_ (.Y(_1511_),
    .A(_1510_));
 sg13g2_nor2_1 _3180_ (.A(_1498_),
    .B(_1477_),
    .Y(_1512_));
 sg13g2_buf_2 _3181_ (.A(_1512_),
    .X(_1513_));
 sg13g2_buf_1 _3182_ (.A(\i_project.controller_0.h[0] ),
    .X(_1514_));
 sg13g2_buf_1 _3183_ (.A(\i_project.controller_0.h[1] ),
    .X(_1515_));
 sg13g2_inv_1 _3184_ (.Y(_1516_),
    .A(net79));
 sg13g2_nor2_1 _3185_ (.A(net80),
    .B(_1516_),
    .Y(_1517_));
 sg13g2_buf_1 _3186_ (.A(\i_project.controller_0.h[3] ),
    .X(_1518_));
 sg13g2_inv_1 _3187_ (.Y(_1519_),
    .A(_1518_));
 sg13g2_buf_2 _3188_ (.A(\i_project.controller_0.h[2] ),
    .X(_1520_));
 sg13g2_buf_1 _3189_ (.A(_1520_),
    .X(_1521_));
 sg13g2_inv_1 _3190_ (.Y(_1522_),
    .A(net68));
 sg13g2_nand3_1 _3191_ (.B(_1519_),
    .C(_1522_),
    .A(_1517_),
    .Y(_1523_));
 sg13g2_buf_1 _3192_ (.A(\i_project.controller_0.h[4] ),
    .X(_1524_));
 sg13g2_buf_1 _3193_ (.A(_1524_),
    .X(_1525_));
 sg13g2_buf_1 _3194_ (.A(\i_project.controller_0.h[5] ),
    .X(_1526_));
 sg13g2_inv_1 _3195_ (.Y(_1527_),
    .A(_1526_));
 sg13g2_nor2_1 _3196_ (.A(net67),
    .B(_1527_),
    .Y(_1528_));
 sg13g2_buf_2 _3197_ (.A(\i_project.controller_0.h[8] ),
    .X(_1529_));
 sg13g2_inv_1 _3198_ (.Y(_1530_),
    .A(_1529_));
 sg13g2_nor2_1 _3199_ (.A(\i_project.controller_0.h[9] ),
    .B(_1530_),
    .Y(_1531_));
 sg13g2_buf_2 _3200_ (.A(\i_project.controller_0.h[6] ),
    .X(_1532_));
 sg13g2_buf_1 _3201_ (.A(_1532_),
    .X(_1533_));
 sg13g2_buf_2 _3202_ (.A(\i_project.controller_0.h[7] ),
    .X(_1534_));
 sg13g2_inv_1 _3203_ (.Y(_1535_),
    .A(net78));
 sg13g2_nor2_1 _3204_ (.A(net66),
    .B(_1535_),
    .Y(_1536_));
 sg13g2_nand3_1 _3205_ (.B(_1531_),
    .C(_1536_),
    .A(_1528_),
    .Y(_1537_));
 sg13g2_nor2_1 _3206_ (.A(_1523_),
    .B(_1537_),
    .Y(_1538_));
 sg13g2_nor3_1 _3207_ (.A(_1511_),
    .B(_1513_),
    .C(_1538_),
    .Y(_1539_));
 sg13g2_buf_1 _3208_ (.A(_1518_),
    .X(_1540_));
 sg13g2_nor2_2 _3209_ (.A(_1515_),
    .B(net80),
    .Y(_1541_));
 sg13g2_inv_1 _3210_ (.Y(_1542_),
    .A(_1541_));
 sg13g2_nor3_1 _3211_ (.A(net65),
    .B(net68),
    .C(_1542_),
    .Y(_1543_));
 sg13g2_inv_2 _3212_ (.Y(_1544_),
    .A(\i_project.controller_0.h[9] ));
 sg13g2_nor2_1 _3213_ (.A(_1529_),
    .B(_1544_),
    .Y(_1545_));
 sg13g2_nand2_1 _3214_ (.Y(_1546_),
    .A(_1543_),
    .B(_1545_));
 sg13g2_inv_1 _3215_ (.Y(_1547_),
    .A(_1546_));
 sg13g2_inv_1 _3216_ (.Y(_1548_),
    .A(net66));
 sg13g2_buf_1 _3217_ (.A(_1526_),
    .X(_1549_));
 sg13g2_nand2_1 _3218_ (.Y(_1550_),
    .A(net67),
    .B(net64));
 sg13g2_nor3_1 _3219_ (.A(_1548_),
    .B(_1535_),
    .C(_1550_),
    .Y(_1551_));
 sg13g2_inv_1 _3220_ (.Y(_1552_),
    .A(_1513_));
 sg13g2_nand2_1 _3221_ (.Y(_1553_),
    .A(_1552_),
    .B(_0022_));
 sg13g2_a21oi_1 _3222_ (.A1(_1547_),
    .A2(_1551_),
    .Y(_1554_),
    .B1(_1553_));
 sg13g2_nor2_1 _3223_ (.A(_1539_),
    .B(_1554_),
    .Y(_1555_));
 sg13g2_inv_1 _3224_ (.Y(_1556_),
    .A(_1524_));
 sg13g2_nor2_1 _3225_ (.A(net64),
    .B(_1556_),
    .Y(_1557_));
 sg13g2_nand2_1 _3226_ (.Y(_1558_),
    .A(_1536_),
    .B(_1557_));
 sg13g2_o21ai_1 _3227_ (.B1(_1554_),
    .Y(_1559_),
    .A1(_1546_),
    .A2(_1558_));
 sg13g2_nor3_1 _3228_ (.A(_1548_),
    .B(net78),
    .C(_1550_),
    .Y(_1560_));
 sg13g2_nand2_1 _3229_ (.Y(_1561_),
    .A(_1540_),
    .B(net68));
 sg13g2_inv_1 _3230_ (.Y(_1562_),
    .A(_1561_));
 sg13g2_nand4_1 _3231_ (.B(_1531_),
    .C(_1541_),
    .A(_1560_),
    .Y(_1563_),
    .D(_1562_));
 sg13g2_nand2_1 _3232_ (.Y(_1564_),
    .A(_1539_),
    .B(_1563_));
 sg13g2_a21oi_1 _3233_ (.A1(_1559_),
    .A2(_1564_),
    .Y(_1565_),
    .B1(\i_project.controller_0.vga_sync.hsync ));
 sg13g2_nor2_1 _3234_ (.A(_1555_),
    .B(_1565_),
    .Y(_0123_));
 sg13g2_nor2_1 _3235_ (.A(\i_project.controller_0.vga_sync.vsync ),
    .B(_1511_),
    .Y(_1566_));
 sg13g2_buf_1 _3236_ (.A(\i_project.controller_0.v[7] ),
    .X(_1567_));
 sg13g2_inv_1 _3237_ (.Y(_1568_),
    .A(_1567_));
 sg13g2_buf_8 _3238_ (.A(\i_project.controller_0.v[4] ),
    .X(_1569_));
 sg13g2_buf_2 _3239_ (.A(\i_project.controller_0.v[6] ),
    .X(_1570_));
 sg13g2_nor2_1 _3240_ (.A(_1569_),
    .B(_1570_),
    .Y(_1571_));
 sg13g2_buf_8 _3241_ (.A(\i_project.controller_0.v[5] ),
    .X(_1572_));
 sg13g2_inv_1 _3242_ (.Y(_1573_),
    .A(_1572_));
 sg13g2_nand2_1 _3243_ (.Y(_1574_),
    .A(_1571_),
    .B(_1573_));
 sg13g2_nor2_1 _3244_ (.A(_1568_),
    .B(_1574_),
    .Y(_1575_));
 sg13g2_buf_8 _3245_ (.A(\i_project.controller_0.v[0] ),
    .X(_1576_));
 sg13g2_inv_2 _3246_ (.Y(_1577_),
    .A(_1576_));
 sg13g2_buf_8 _3247_ (.A(\i_project.controller_0.v[1] ),
    .X(_1578_));
 sg13g2_buf_2 _3248_ (.A(\i_project.controller_0.v[8] ),
    .X(_1579_));
 sg13g2_buf_1 _3249_ (.A(\i_project.controller_0.v[9] ),
    .X(_1580_));
 sg13g2_nand2_1 _3250_ (.Y(_1581_),
    .A(_1579_),
    .B(_1580_));
 sg13g2_nor3_1 _3251_ (.A(_1577_),
    .B(net77),
    .C(_1581_),
    .Y(_1582_));
 sg13g2_buf_1 _3252_ (.A(\i_project.controller_0.v[2] ),
    .X(_1583_));
 sg13g2_buf_1 _3253_ (.A(\i_project.controller_0.v[3] ),
    .X(_1584_));
 sg13g2_inv_1 _3254_ (.Y(_1585_),
    .A(net75));
 sg13g2_nand4_1 _3255_ (.B(_1582_),
    .C(net76),
    .A(_1575_),
    .Y(_1586_),
    .D(_1585_));
 sg13g2_inv_1 _3256_ (.Y(_1587_),
    .A(net76));
 sg13g2_nand4_1 _3257_ (.B(_1587_),
    .C(net77),
    .A(_1577_),
    .Y(_1588_),
    .D(net75));
 sg13g2_nand2_1 _3258_ (.Y(_1589_),
    .A(_1567_),
    .B(_1579_));
 sg13g2_inv_1 _3259_ (.Y(_1590_),
    .A(_1589_));
 sg13g2_nor2_1 _3260_ (.A(_1569_),
    .B(_1580_),
    .Y(_1591_));
 sg13g2_nand4_1 _3261_ (.B(_1591_),
    .C(_1572_),
    .A(_1590_),
    .Y(_1592_),
    .D(_1570_));
 sg13g2_nor2_1 _3262_ (.A(_1588_),
    .B(_1592_),
    .Y(_1593_));
 sg13g2_nor4_1 _3263_ (.A(_1576_),
    .B(net77),
    .C(_1587_),
    .D(_1585_),
    .Y(_1594_));
 sg13g2_nand2b_1 _3264_ (.Y(_1595_),
    .B(_1594_),
    .A_N(_1592_));
 sg13g2_o21ai_1 _3265_ (.B1(_1595_),
    .Y(_1596_),
    .A1(\i_project.controller_0.vga_sync.vsync ),
    .A2(_1593_));
 sg13g2_nor2_1 _3266_ (.A(_1576_),
    .B(net77),
    .Y(_1597_));
 sg13g2_nand3_1 _3267_ (.B(_1587_),
    .C(net75),
    .A(_1597_),
    .Y(_1598_));
 sg13g2_nor2_1 _3268_ (.A(_1574_),
    .B(_1598_),
    .Y(_1599_));
 sg13g2_nor3_1 _3269_ (.A(_1511_),
    .B(_1568_),
    .C(_1581_),
    .Y(_1600_));
 sg13g2_a21o_1 _3270_ (.A2(_1600_),
    .A1(_1599_),
    .B1(_1513_),
    .X(_1601_));
 sg13g2_a221oi_1 _3271_ (.B2(_1511_),
    .C1(_1601_),
    .B1(_1596_),
    .A1(_1566_),
    .Y(_0134_),
    .A2(_1586_));
 sg13g2_inv_1 _3272_ (.Y(_1602_),
    .A(\i_project.controller_0.voffset[0] ));
 sg13g2_nand3_1 _3273_ (.B(net66),
    .C(_1535_),
    .A(_1531_),
    .Y(_1603_));
 sg13g2_nor2_1 _3274_ (.A(_1521_),
    .B(_1519_),
    .Y(_1604_));
 sg13g2_nand3_1 _3275_ (.B(_1604_),
    .C(_1541_),
    .A(_1528_),
    .Y(_1605_));
 sg13g2_a21oi_1 _3276_ (.A1(_1556_),
    .A2(_0024_),
    .Y(_1606_),
    .B1(_1527_));
 sg13g2_nor2_1 _3277_ (.A(net66),
    .B(net78),
    .Y(_1607_));
 sg13g2_o21ai_1 _3278_ (.B1(_1544_),
    .Y(_1608_),
    .A1(_1530_),
    .A2(_1607_));
 sg13g2_o21ai_1 _3279_ (.B1(_1608_),
    .Y(_1609_),
    .A1(_1606_),
    .A2(_1603_));
 sg13g2_o21ai_1 _3280_ (.B1(_1609_),
    .Y(_1610_),
    .A1(_1603_),
    .A2(_1605_));
 sg13g2_nor2_1 _3281_ (.A(_1510_),
    .B(_1544_),
    .Y(_1611_));
 sg13g2_nand4_1 _3282_ (.B(_1556_),
    .C(_1527_),
    .A(_1543_),
    .Y(_1612_),
    .D(_1536_));
 sg13g2_nand3_1 _3283_ (.B(_1530_),
    .C(_0023_),
    .A(_1612_),
    .Y(_1613_));
 sg13g2_a22oi_1 _3284_ (.Y(_1614_),
    .B1(_1611_),
    .B2(_1613_),
    .A2(_1610_),
    .A1(_1510_));
 sg13g2_xor2_1 _3285_ (.B(\i_project.controller_0.mode[2] ),
    .A(\i_project.controller_0.grey_pass[14] ),
    .X(_1615_));
 sg13g2_buf_2 _3286_ (.A(\i_project.controller_0.mode[1] ),
    .X(_1616_));
 sg13g2_xor2_1 _3287_ (.B(\i_project.controller_0.grey_pass[13] ),
    .A(_1616_),
    .X(_1617_));
 sg13g2_nor2_1 _3288_ (.A(_1615_),
    .B(_1617_),
    .Y(_1618_));
 sg13g2_buf_2 _3289_ (.A(\i_project.controller_0.mode[0] ),
    .X(_1619_));
 sg13g2_xnor2_1 _3290_ (.Y(_1620_),
    .A(_1619_),
    .B(\i_project.controller_0.grey_pass[12] ));
 sg13g2_inv_1 _3291_ (.Y(_1621_),
    .A(_0025_));
 sg13g2_nor3_1 _3292_ (.A(_1616_),
    .B(_1619_),
    .C(_1621_),
    .Y(_1622_));
 sg13g2_buf_2 _3293_ (.A(_1622_),
    .X(_1623_));
 sg13g2_buf_1 _3294_ (.A(_1623_),
    .X(_1624_));
 sg13g2_a21oi_1 _3295_ (.A1(_1618_),
    .A2(_1620_),
    .Y(_1625_),
    .B1(net56));
 sg13g2_nand2b_1 _3296_ (.Y(_1626_),
    .B(_1625_),
    .A_N(_1614_));
 sg13g2_nand2_2 _3297_ (.Y(_1627_),
    .A(_1626_),
    .B(_1498_));
 sg13g2_inv_2 _3298_ (.Y(_1628_),
    .A(_1627_));
 sg13g2_nand2b_1 _3299_ (.Y(_1629_),
    .B(net69),
    .A_N(_1620_));
 sg13g2_inv_1 _3300_ (.Y(_1630_),
    .A(\i_project.controller_0.mode[2] ));
 sg13g2_nor3_1 _3301_ (.A(_1616_),
    .B(_1498_),
    .C(_1630_),
    .Y(_1631_));
 sg13g2_nand2_1 _3302_ (.Y(_1632_),
    .A(_1631_),
    .B(_0016_));
 sg13g2_nor2b_2 _3303_ (.A(_1628_),
    .B_N(_1632_),
    .Y(_1633_));
 sg13g2_a22oi_1 _3304_ (.Y(_0135_),
    .B1(_1629_),
    .B2(_1633_),
    .A2(_1628_),
    .A1(_1602_));
 sg13g2_a22oi_1 _3305_ (.Y(_1634_),
    .B1(net69),
    .B2(_1617_),
    .A2(_0015_),
    .A1(_1631_));
 sg13g2_buf_8 _3306_ (.A(\i_project.controller_0.voffset[1] ),
    .X(_1635_));
 sg13g2_nor2_1 _3307_ (.A(_1635_),
    .B(_1627_),
    .Y(_1636_));
 sg13g2_a21oi_1 _3308_ (.A1(_1627_),
    .A2(_1634_),
    .Y(_0136_),
    .B1(_1636_));
 sg13g2_buf_2 _3309_ (.A(\i_project.controller_0.voffset[2] ),
    .X(_1637_));
 sg13g2_inv_1 _3310_ (.Y(_1638_),
    .A(_1637_));
 sg13g2_nand2_1 _3311_ (.Y(_1639_),
    .A(_1615_),
    .B(net69));
 sg13g2_a22oi_1 _3312_ (.Y(_0137_),
    .B1(_1639_),
    .B2(_1633_),
    .A2(_1628_),
    .A1(_1638_));
 sg13g2_inv_1 _3313_ (.Y(_1640_),
    .A(\i_project.controller_0.voffset[3] ));
 sg13g2_nand2_1 _3314_ (.Y(_1641_),
    .A(_1631_),
    .B(_0145_));
 sg13g2_o21ai_1 _3315_ (.B1(_1641_),
    .Y(_0138_),
    .A1(_1640_),
    .A2(_1627_));
 sg13g2_inv_1 _3316_ (.Y(_1642_),
    .A(\i_project.controller_0.voffset[4] ));
 sg13g2_o21ai_1 _3317_ (.B1(_1632_),
    .Y(_0139_),
    .A1(_1642_),
    .A2(_1627_));
 sg13g2_inv_1 _3318_ (.Y(_1643_),
    .A(\i_project.controller_0.voffset[5] ));
 sg13g2_buf_1 _3319_ (.A(_1499_),
    .X(_1644_));
 sg13g2_nand2_1 _3320_ (.Y(_1645_),
    .A(net58),
    .B(\i_project.controller_0.grey_pass[10] ));
 sg13g2_a22oi_1 _3321_ (.Y(_0140_),
    .B1(_1645_),
    .B2(_1633_),
    .A2(_1628_),
    .A1(_1643_));
 sg13g2_inv_1 _3322_ (.Y(_1646_),
    .A(\i_project.controller_0.voffset[6] ));
 sg13g2_nand2_1 _3323_ (.Y(_1647_),
    .A(net58),
    .B(\i_project.controller_0.grey_pass[11] ));
 sg13g2_a22oi_1 _3324_ (.Y(_0141_),
    .B1(_1647_),
    .B2(_1633_),
    .A2(_1628_),
    .A1(_1646_));
 sg13g2_inv_1 _3325_ (.Y(_1648_),
    .A(net69));
 sg13g2_inv_1 _3326_ (.Y(_1649_),
    .A(\i_project.controller_0.grey_pass[15] ));
 sg13g2_nor3_1 _3327_ (.A(_1648_),
    .B(_1649_),
    .C(_1626_),
    .Y(_1650_));
 sg13g2_a21o_1 _3328_ (.A2(_1628_),
    .A1(\i_project.controller_0.voffset[7] ),
    .B1(_1650_),
    .X(_0142_));
 sg13g2_inv_1 _3329_ (.Y(_1651_),
    .A(_1619_));
 sg13g2_nor2_1 _3330_ (.A(\i_project.controller_0.grey_pass[12] ),
    .B(net58),
    .Y(_1652_));
 sg13g2_a21oi_1 _3331_ (.A1(_1651_),
    .A2(net58),
    .Y(_0097_),
    .B1(_1652_));
 sg13g2_inv_1 _3332_ (.Y(_1653_),
    .A(_1616_));
 sg13g2_nor2_1 _3333_ (.A(\i_project.controller_0.grey_pass[13] ),
    .B(net58),
    .Y(_1654_));
 sg13g2_a21oi_1 _3334_ (.A1(_1653_),
    .A2(net58),
    .Y(_0098_),
    .B1(_1654_));
 sg13g2_nor2_1 _3335_ (.A(\i_project.controller_0.grey_pass[14] ),
    .B(_1644_),
    .Y(_1655_));
 sg13g2_a21oi_1 _3336_ (.A1(_1630_),
    .A2(_1644_),
    .Y(_0099_),
    .B1(_1655_));
 sg13g2_nand2_1 _3337_ (.Y(_1656_),
    .A(_1510_),
    .B(net58));
 sg13g2_o21ai_1 _3338_ (.B1(_1656_),
    .Y(_0100_),
    .A1(net58),
    .A2(_1649_));
 sg13g2_buf_2 _3339_ (.A(\dither_threshold[3] ),
    .X(_1657_));
 sg13g2_buf_1 _3340_ (.A(\dither_threshold[2] ),
    .X(_1658_));
 sg13g2_nand2_1 _3341_ (.Y(_1659_),
    .A(_1657_),
    .B(_1658_));
 sg13g2_inv_1 _3342_ (.Y(_1660_),
    .A(_1659_));
 sg13g2_buf_2 _3343_ (.A(\dither_threshold[1] ),
    .X(_1661_));
 sg13g2_inv_1 _3344_ (.Y(_1662_),
    .A(_1661_));
 sg13g2_nand3_1 _3345_ (.B(_1662_),
    .C(_0029_),
    .A(_1660_),
    .Y(_1663_));
 sg13g2_buf_2 _3346_ (.A(_0028_),
    .X(_1664_));
 sg13g2_inv_1 _3347_ (.Y(_1665_),
    .A(_1664_));
 sg13g2_nand3_1 _3348_ (.B(_1657_),
    .C(_1665_),
    .A(_1663_),
    .Y(_1666_));
 sg13g2_inv_1 _3349_ (.Y(_1667_),
    .A(\dither_threshold[4] ));
 sg13g2_buf_1 _3350_ (.A(\dither_threshold[0] ),
    .X(_1668_));
 sg13g2_inv_1 _3351_ (.Y(_1669_),
    .A(_1668_));
 sg13g2_buf_1 _3352_ (.A(_0027_),
    .X(_1670_));
 sg13g2_nand4_1 _3353_ (.B(_1662_),
    .C(_1669_),
    .A(_1660_),
    .Y(_1671_),
    .D(_1670_));
 sg13g2_nand3_1 _3354_ (.B(_1667_),
    .C(_1671_),
    .A(_1666_),
    .Y(_1672_));
 sg13g2_buf_1 _3355_ (.A(_1672_),
    .X(_1673_));
 sg13g2_inv_1 _3356_ (.Y(_1674_),
    .A(_1673_));
 sg13g2_nand2_1 _3357_ (.Y(_1675_),
    .A(_1674_),
    .B(_1669_));
 sg13g2_nand2_1 _3358_ (.Y(_1676_),
    .A(_1673_),
    .B(_1668_));
 sg13g2_inv_1 _3359_ (.Y(_1677_),
    .A(\frame_counter[1] ));
 sg13g2_inv_1 _3360_ (.Y(_1678_),
    .A(\frame_counter[0] ));
 sg13g2_nand2_1 _3361_ (.Y(_1679_),
    .A(_1677_),
    .B(_1678_));
 sg13g2_nand2_1 _3362_ (.Y(_1680_),
    .A(_1649_),
    .B(prev_vsync));
 sg13g2_xnor2_1 _3363_ (.Y(\i_project.controller_0.vga_sync.o_vsync ),
    .A(_1510_),
    .B(\i_project.controller_0.vga_sync.vsync ));
 sg13g2_nor2_1 _3364_ (.A(_1680_),
    .B(\i_project.controller_0.vga_sync.o_vsync ),
    .Y(_1681_));
 sg13g2_nand3b_1 _3365_ (.B(\i_project.controller_0.vga_sync.o_vsync ),
    .C(\i_project.controller_0.grey_pass[15] ),
    .Y(_1682_),
    .A_N(prev_vsync));
 sg13g2_nand2b_1 _3366_ (.Y(_1683_),
    .B(_1682_),
    .A_N(_1681_));
 sg13g2_inv_1 _3367_ (.Y(_1684_),
    .A(_1683_));
 sg13g2_buf_1 _3368_ (.A(_1477_),
    .X(_1685_));
 sg13g2_o21ai_1 _3369_ (.B1(_1685_),
    .Y(_1686_),
    .A1(_1679_),
    .A2(_1684_));
 sg13g2_buf_1 _3370_ (.A(_1686_),
    .X(_1687_));
 sg13g2_a21oi_1 _3371_ (.A1(_1675_),
    .A2(_1676_),
    .Y(_0090_),
    .B1(_1687_));
 sg13g2_nor2_1 _3372_ (.A(_1661_),
    .B(_1674_),
    .Y(_1688_));
 sg13g2_nand2_1 _3373_ (.Y(_1689_),
    .A(_1662_),
    .B(_1669_));
 sg13g2_nand2_1 _3374_ (.Y(_1690_),
    .A(_1661_),
    .B(_1668_));
 sg13g2_a21oi_1 _3375_ (.A1(_1689_),
    .A2(_1690_),
    .Y(_1691_),
    .B1(_1673_));
 sg13g2_nor3_1 _3376_ (.A(_1687_),
    .B(_1688_),
    .C(_1691_),
    .Y(_0091_));
 sg13g2_nor2_1 _3377_ (.A(_1690_),
    .B(_1673_),
    .Y(_1692_));
 sg13g2_xnor2_1 _3378_ (.Y(_1693_),
    .A(_1664_),
    .B(_1692_));
 sg13g2_nor2_1 _3379_ (.A(_1687_),
    .B(_1693_),
    .Y(_0092_));
 sg13g2_inv_1 _3380_ (.Y(_1694_),
    .A(_1657_));
 sg13g2_inv_1 _3381_ (.Y(_1695_),
    .A(_1658_));
 sg13g2_nand2_1 _3382_ (.Y(_1696_),
    .A(_1694_),
    .B(_1695_));
 sg13g2_nand3_1 _3383_ (.B(_1659_),
    .C(_1696_),
    .A(_1673_),
    .Y(_1697_));
 sg13g2_buf_2 _3384_ (.A(_0033_),
    .X(_1698_));
 sg13g2_o21ai_1 _3385_ (.B1(_1664_),
    .Y(_1699_),
    .A1(_1658_),
    .A2(_1690_));
 sg13g2_xnor2_1 _3386_ (.Y(_1700_),
    .A(_1698_),
    .B(_1699_));
 sg13g2_nand2_1 _3387_ (.Y(_1701_),
    .A(_1674_),
    .B(_1700_));
 sg13g2_a21oi_1 _3388_ (.A1(_1697_),
    .A2(_1701_),
    .Y(_0093_),
    .B1(_1687_));
 sg13g2_a21oi_1 _3389_ (.A1(_1690_),
    .A2(_1695_),
    .Y(_1702_),
    .B1(_1694_));
 sg13g2_nor2_1 _3390_ (.A(_1660_),
    .B(_1674_),
    .Y(_1703_));
 sg13g2_a21oi_1 _3391_ (.A1(_1674_),
    .A2(_1702_),
    .Y(_1704_),
    .B1(_1703_));
 sg13g2_nor2_1 _3392_ (.A(_1670_),
    .B(_1704_),
    .Y(_1705_));
 sg13g2_inv_1 _3393_ (.Y(_1706_),
    .A(_1670_));
 sg13g2_nor2b_1 _3394_ (.A(_1706_),
    .B_N(_1704_),
    .Y(_1707_));
 sg13g2_nor3_1 _3395_ (.A(_1687_),
    .B(_1705_),
    .C(_1707_),
    .Y(_0094_));
 sg13g2_inv_1 _3396_ (.Y(_1708_),
    .A(_0053_));
 sg13g2_nand4_1 _3397_ (.B(net66),
    .C(net78),
    .A(_1544_),
    .Y(_1709_),
    .D(_1510_));
 sg13g2_nand2_1 _3398_ (.Y(_1710_),
    .A(net79),
    .B(_1514_));
 sg13g2_inv_1 _3399_ (.Y(_1711_),
    .A(_1710_));
 sg13g2_inv_1 _3400_ (.Y(_1712_),
    .A(_0024_));
 sg13g2_inv_1 _3401_ (.Y(_1713_),
    .A(_0026_));
 sg13g2_nand4_1 _3402_ (.B(_1557_),
    .C(_1712_),
    .A(_1711_),
    .Y(_1714_),
    .D(_1713_));
 sg13g2_a21oi_1 _3403_ (.A1(_1522_),
    .A2(_1709_),
    .Y(_1715_),
    .B1(_1714_));
 sg13g2_a21o_1 _3404_ (.A2(_1607_),
    .A1(_1611_),
    .B1(_1522_),
    .X(_1716_));
 sg13g2_nand2_2 _3405_ (.Y(_1717_),
    .A(_1715_),
    .B(_1716_));
 sg13g2_inv_1 _3406_ (.Y(_1718_),
    .A(_1717_));
 sg13g2_nor2_1 _3407_ (.A(_1513_),
    .B(_1718_),
    .Y(_1719_));
 sg13g2_inv_1 _3408_ (.Y(_1720_),
    .A(_1719_));
 sg13g2_buf_1 _3409_ (.A(_1720_),
    .X(_1721_));
 sg13g2_nor2_1 _3410_ (.A(_1708_),
    .B(net28),
    .Y(_0113_));
 sg13g2_nor3_1 _3411_ (.A(_1541_),
    .B(_1711_),
    .C(_1721_),
    .Y(_0114_));
 sg13g2_nor2_1 _3412_ (.A(_1521_),
    .B(_1711_),
    .Y(_1722_));
 sg13g2_nor2_1 _3413_ (.A(_1522_),
    .B(_1710_),
    .Y(_1723_));
 sg13g2_nor3_1 _3414_ (.A(_1722_),
    .B(_1723_),
    .C(net28),
    .Y(_0115_));
 sg13g2_nor2_1 _3415_ (.A(net65),
    .B(_1723_),
    .Y(_1724_));
 sg13g2_nor2_1 _3416_ (.A(_1561_),
    .B(_1710_),
    .Y(_1725_));
 sg13g2_nor3_1 _3417_ (.A(_1724_),
    .B(_1725_),
    .C(net28),
    .Y(_0116_));
 sg13g2_nor2_1 _3418_ (.A(net67),
    .B(_1725_),
    .Y(_1726_));
 sg13g2_nand2_1 _3419_ (.Y(_1727_),
    .A(_1725_),
    .B(_1525_));
 sg13g2_inv_1 _3420_ (.Y(_1728_),
    .A(_1727_));
 sg13g2_nor3_1 _3421_ (.A(_1726_),
    .B(_1728_),
    .C(net28),
    .Y(_0117_));
 sg13g2_nor2_1 _3422_ (.A(_1549_),
    .B(_1728_),
    .Y(_1729_));
 sg13g2_nor2_1 _3423_ (.A(_1527_),
    .B(_1727_),
    .Y(_1730_));
 sg13g2_nor3_1 _3424_ (.A(_1729_),
    .B(_1730_),
    .C(net28),
    .Y(_0118_));
 sg13g2_nor2_1 _3425_ (.A(_1533_),
    .B(_1730_),
    .Y(_1731_));
 sg13g2_nand2_1 _3426_ (.Y(_1732_),
    .A(_1730_),
    .B(_1533_));
 sg13g2_inv_1 _3427_ (.Y(_1733_),
    .A(_1732_));
 sg13g2_nor3_1 _3428_ (.A(_1731_),
    .B(_1733_),
    .C(net28),
    .Y(_0119_));
 sg13g2_nor2_1 _3429_ (.A(net78),
    .B(_1733_),
    .Y(_1734_));
 sg13g2_nor2_1 _3430_ (.A(_1535_),
    .B(_1732_),
    .Y(_1735_));
 sg13g2_nor3_1 _3431_ (.A(_1734_),
    .B(_1735_),
    .C(net28),
    .Y(_0120_));
 sg13g2_nor2_1 _3432_ (.A(_1529_),
    .B(_1735_),
    .Y(_1736_));
 sg13g2_nand2_1 _3433_ (.Y(_1737_),
    .A(_1735_),
    .B(_1529_));
 sg13g2_inv_1 _3434_ (.Y(_1738_),
    .A(_1737_));
 sg13g2_nor3_1 _3435_ (.A(_1736_),
    .B(_1738_),
    .C(net28),
    .Y(_0121_));
 sg13g2_o21ai_1 _3436_ (.B1(_1719_),
    .Y(_1739_),
    .A1(_1544_),
    .A2(_1737_));
 sg13g2_a21oi_1 _3437_ (.A1(_1544_),
    .A2(_1737_),
    .Y(_0122_),
    .B1(_1739_));
 sg13g2_nor2_1 _3438_ (.A(_1567_),
    .B(_1574_),
    .Y(_1740_));
 sg13g2_inv_1 _3439_ (.Y(_1741_),
    .A(_1579_));
 sg13g2_nand4_1 _3440_ (.B(_1511_),
    .C(_1740_),
    .A(_1594_),
    .Y(_1742_),
    .D(_1741_));
 sg13g2_nor3_1 _3441_ (.A(_1511_),
    .B(_1573_),
    .C(_1589_),
    .Y(_1743_));
 sg13g2_nor2_1 _3442_ (.A(net76),
    .B(net75),
    .Y(_1744_));
 sg13g2_nand2_1 _3443_ (.Y(_1745_),
    .A(_1576_),
    .B(net77));
 sg13g2_inv_1 _3444_ (.Y(_1746_),
    .A(_1745_));
 sg13g2_nand4_1 _3445_ (.B(_1571_),
    .C(_1744_),
    .A(_1743_),
    .Y(_1747_),
    .D(_1746_));
 sg13g2_a21o_1 _3446_ (.A2(_1747_),
    .A1(_1742_),
    .B1(_0030_),
    .X(_1748_));
 sg13g2_nand2_1 _3447_ (.Y(_1749_),
    .A(_1748_),
    .B(_1718_));
 sg13g2_nor2_1 _3448_ (.A(_1577_),
    .B(_1717_),
    .Y(_1750_));
 sg13g2_a221oi_1 _3449_ (.B2(_1577_),
    .C1(_1750_),
    .B1(_1749_),
    .A1(_1648_),
    .Y(_0124_),
    .A2(net82));
 sg13g2_nor2_1 _3450_ (.A(_1578_),
    .B(_1750_),
    .Y(_1751_));
 sg13g2_inv_1 _3451_ (.Y(_1752_),
    .A(_1578_));
 sg13g2_inv_1 _3452_ (.Y(_1753_),
    .A(_1750_));
 sg13g2_nor2_1 _3453_ (.A(_1752_),
    .B(_1753_),
    .Y(_1754_));
 sg13g2_nor3_1 _3454_ (.A(_1513_),
    .B(_1751_),
    .C(_1754_),
    .Y(_0125_));
 sg13g2_nor3_1 _3455_ (.A(_1752_),
    .B(_1587_),
    .C(_1753_),
    .Y(_1755_));
 sg13g2_nor2_1 _3456_ (.A(net76),
    .B(_1754_),
    .Y(_1756_));
 sg13g2_nor2_2 _3457_ (.A(_1717_),
    .B(_1748_),
    .Y(_1757_));
 sg13g2_inv_1 _3458_ (.Y(_1758_),
    .A(_1757_));
 sg13g2_nand2_1 _3459_ (.Y(_1759_),
    .A(_1758_),
    .B(_1552_));
 sg13g2_nor3_1 _3460_ (.A(_1755_),
    .B(_1756_),
    .C(_1759_),
    .Y(_0126_));
 sg13g2_nand3_1 _3461_ (.B(_1583_),
    .C(net75),
    .A(_1746_),
    .Y(_1760_));
 sg13g2_nor2_1 _3462_ (.A(_1760_),
    .B(_1717_),
    .Y(_1761_));
 sg13g2_nor2_1 _3463_ (.A(_1584_),
    .B(_1755_),
    .Y(_1762_));
 sg13g2_nor3_1 _3464_ (.A(_1761_),
    .B(_1762_),
    .C(_1759_),
    .Y(_0127_));
 sg13g2_inv_1 _3465_ (.Y(_1763_),
    .A(_1569_));
 sg13g2_nor3_1 _3466_ (.A(_1763_),
    .B(_1760_),
    .C(_1717_),
    .Y(_1764_));
 sg13g2_nor2_1 _3467_ (.A(_1569_),
    .B(_1761_),
    .Y(_1765_));
 sg13g2_nor3_1 _3468_ (.A(_1513_),
    .B(_1764_),
    .C(_1765_),
    .Y(_0128_));
 sg13g2_nor2_1 _3469_ (.A(_1513_),
    .B(_1749_),
    .Y(_1766_));
 sg13g2_nor2_1 _3470_ (.A(_1763_),
    .B(_1760_),
    .Y(_1767_));
 sg13g2_xnor2_1 _3471_ (.Y(_1768_),
    .A(_0031_),
    .B(_1767_));
 sg13g2_nand2_1 _3472_ (.Y(_1769_),
    .A(_1766_),
    .B(_1768_));
 sg13g2_o21ai_1 _3473_ (.B1(_1769_),
    .Y(_0129_),
    .A1(_1573_),
    .A2(_1721_));
 sg13g2_a21oi_1 _3474_ (.A1(_1764_),
    .A2(_1572_),
    .Y(_1770_),
    .B1(_1570_));
 sg13g2_nand3_1 _3475_ (.B(_1572_),
    .C(_1570_),
    .A(_1764_),
    .Y(_1771_));
 sg13g2_nand2b_1 _3476_ (.Y(_1772_),
    .B(_1771_),
    .A_N(_1770_));
 sg13g2_nor2_1 _3477_ (.A(_1759_),
    .B(_1772_),
    .Y(_0130_));
 sg13g2_nand3_1 _3478_ (.B(_1572_),
    .C(_1570_),
    .A(_1767_),
    .Y(_1773_));
 sg13g2_nor2_1 _3479_ (.A(_1568_),
    .B(_1773_),
    .Y(_1774_));
 sg13g2_a221oi_1 _3480_ (.B2(_1568_),
    .C1(_1759_),
    .B1(_1771_),
    .A1(_1718_),
    .Y(_0131_),
    .A2(_1774_));
 sg13g2_xnor2_1 _3481_ (.Y(_1775_),
    .A(_0032_),
    .B(_1774_));
 sg13g2_nand2_1 _3482_ (.Y(_1776_),
    .A(_1766_),
    .B(_1775_));
 sg13g2_o21ai_1 _3483_ (.B1(_1776_),
    .Y(_0132_),
    .A1(_1741_),
    .A2(_1720_));
 sg13g2_inv_1 _3484_ (.Y(_1777_),
    .A(_1580_));
 sg13g2_nor2_1 _3485_ (.A(_1589_),
    .B(_1773_),
    .Y(_1778_));
 sg13g2_xnor2_1 _3486_ (.Y(_1779_),
    .A(_0030_),
    .B(_1778_));
 sg13g2_nand2_1 _3487_ (.Y(_1780_),
    .A(_1766_),
    .B(_1779_));
 sg13g2_o21ai_1 _3488_ (.B1(_1780_),
    .Y(_0133_),
    .A1(_1777_),
    .A2(_1720_));
 sg13g2_and2_1 _3489_ (.A(_0004_),
    .B(_0003_),
    .X(_0057_));
 sg13g2_nand2_1 _3490_ (.Y(_1781_),
    .A(net74),
    .B(_0055_));
 sg13g2_inv_1 _3491_ (.Y(_0058_),
    .A(_1781_));
 sg13g2_o21ai_1 _3492_ (.B1(net74),
    .Y(_1782_),
    .A1(_1443_),
    .A2(_1457_));
 sg13g2_a21oi_1 _3493_ (.A1(_1443_),
    .A2(_1457_),
    .Y(_0059_),
    .B1(_1782_));
 sg13g2_buf_1 _3494_ (.A(net82),
    .X(_1783_));
 sg13g2_nor3_1 _3495_ (.A(_1444_),
    .B(_1443_),
    .C(_1455_),
    .Y(_1784_));
 sg13g2_nor2_1 _3496_ (.A(\counter[11] ),
    .B(_1784_),
    .Y(_1785_));
 sg13g2_nor3_1 _3497_ (.A(net63),
    .B(_1785_),
    .C(_1458_),
    .Y(_0060_));
 sg13g2_nor2_1 _3498_ (.A(\counter[12] ),
    .B(_1458_),
    .Y(_1786_));
 sg13g2_inv_1 _3499_ (.Y(_1787_),
    .A(_1459_));
 sg13g2_nor3_1 _3500_ (.A(net63),
    .B(_1786_),
    .C(_1787_),
    .Y(_0061_));
 sg13g2_nor2_1 _3501_ (.A(\counter[13] ),
    .B(_1787_),
    .Y(_1788_));
 sg13g2_nor3_1 _3502_ (.A(net63),
    .B(_1460_),
    .C(_1788_),
    .Y(_0062_));
 sg13g2_nor2_1 _3503_ (.A(\counter[14] ),
    .B(_1460_),
    .Y(_1789_));
 sg13g2_inv_1 _3504_ (.Y(_1790_),
    .A(_1461_));
 sg13g2_nor3_1 _3505_ (.A(net63),
    .B(_1789_),
    .C(_1790_),
    .Y(_0063_));
 sg13g2_nand3_1 _3506_ (.B(\counter[11] ),
    .C(\counter[12] ),
    .A(_1784_),
    .Y(_1791_));
 sg13g2_nand3b_1 _3507_ (.B(\counter[13] ),
    .C(\counter[14] ),
    .Y(_1792_),
    .A_N(_1791_));
 sg13g2_inv_1 _3508_ (.Y(_1793_),
    .A(_1792_));
 sg13g2_nor2_1 _3509_ (.A(\counter[15] ),
    .B(_1793_),
    .Y(_1794_));
 sg13g2_nor3_1 _3510_ (.A(_1783_),
    .B(_1462_),
    .C(_1794_),
    .Y(_0064_));
 sg13g2_buf_1 _3511_ (.A(_1478_),
    .X(_1795_));
 sg13g2_nor2_1 _3512_ (.A(\counter[16] ),
    .B(_1462_),
    .Y(_1796_));
 sg13g2_nor3_1 _3513_ (.A(net62),
    .B(_1796_),
    .C(_1480_),
    .Y(_0065_));
 sg13g2_inv_1 _3514_ (.Y(_1797_),
    .A(\counter[17] ));
 sg13g2_nand2_1 _3515_ (.Y(_1798_),
    .A(_1480_),
    .B(\counter[17] ));
 sg13g2_nand2_1 _3516_ (.Y(_1799_),
    .A(_1798_),
    .B(net74));
 sg13g2_a21oi_1 _3517_ (.A1(_1797_),
    .A2(_1463_),
    .Y(_0066_),
    .B1(_1799_));
 sg13g2_inv_1 _3518_ (.Y(_1800_),
    .A(_1441_));
 sg13g2_inv_1 _3519_ (.Y(_1801_),
    .A(\counter[18] ));
 sg13g2_a221oi_1 _3520_ (.B2(_1801_),
    .C1(_1783_),
    .B1(_1798_),
    .A1(_1480_),
    .Y(_0067_),
    .A2(_1800_));
 sg13g2_a21oi_1 _3521_ (.A1(_1480_),
    .A2(_1800_),
    .Y(_1802_),
    .B1(\counter[19] ));
 sg13g2_nor3_1 _3522_ (.A(net62),
    .B(_1464_),
    .C(_1802_),
    .Y(_0068_));
 sg13g2_inv_1 _3523_ (.Y(_1803_),
    .A(_1446_));
 sg13g2_nor3_1 _3524_ (.A(net62),
    .B(_1433_),
    .C(_1803_),
    .Y(_0069_));
 sg13g2_nor2_1 _3525_ (.A(\counter[20] ),
    .B(_1464_),
    .Y(_1804_));
 sg13g2_inv_1 _3526_ (.Y(_1805_),
    .A(_1465_));
 sg13g2_nor3_1 _3527_ (.A(net62),
    .B(_1804_),
    .C(_1805_),
    .Y(_0070_));
 sg13g2_nor2_1 _3528_ (.A(\counter[21] ),
    .B(_1805_),
    .Y(_1806_));
 sg13g2_nor3_1 _3529_ (.A(_1795_),
    .B(_1466_),
    .C(_1806_),
    .Y(_0071_));
 sg13g2_inv_1 _3530_ (.Y(_1807_),
    .A(_1466_));
 sg13g2_a221oi_1 _3531_ (.B2(_1484_),
    .C1(net63),
    .B1(_1807_),
    .A1(_1480_),
    .Y(_0072_),
    .A2(_1486_));
 sg13g2_nand2_1 _3532_ (.Y(_1808_),
    .A(_1480_),
    .B(_1486_));
 sg13g2_nand3_1 _3533_ (.B(\counter[23] ),
    .C(_1486_),
    .A(_1480_),
    .Y(_1809_));
 sg13g2_nand2_1 _3534_ (.Y(_1810_),
    .A(_1809_),
    .B(net74));
 sg13g2_a21oi_1 _3535_ (.A1(_1481_),
    .A2(_1808_),
    .Y(_0073_),
    .B1(_1810_));
 sg13g2_o21ai_1 _3536_ (.B1(_1468_),
    .Y(_1811_),
    .A1(_1469_),
    .A2(_1807_));
 sg13g2_nor3_1 _3537_ (.A(_1468_),
    .B(_1469_),
    .C(_1807_),
    .Y(_1812_));
 sg13g2_inv_1 _3538_ (.Y(_1813_),
    .A(_1812_));
 sg13g2_and3_1 _3539_ (.X(_0074_),
    .A(_1811_),
    .B(_1813_),
    .C(_1685_));
 sg13g2_a221oi_1 _3540_ (.B2(_1467_),
    .C1(net63),
    .B1(_1813_),
    .A1(_1470_),
    .Y(_0075_),
    .A2(_1466_));
 sg13g2_a21oi_1 _3541_ (.A1(_1466_),
    .A2(_1470_),
    .Y(_1814_),
    .B1(\counter[26] ));
 sg13g2_nor3_1 _3542_ (.A(_1795_),
    .B(_1814_),
    .C(_1472_),
    .Y(_0076_));
 sg13g2_nor2_1 _3543_ (.A(\counter[2] ),
    .B(_1803_),
    .Y(_1815_));
 sg13g2_nor3_1 _3544_ (.A(net62),
    .B(_1447_),
    .C(_1815_),
    .Y(_0080_));
 sg13g2_inv_1 _3545_ (.Y(_1816_),
    .A(\counter[30] ));
 sg13g2_nor3_1 _3546_ (.A(_1493_),
    .B(_1816_),
    .C(_1473_),
    .Y(_1817_));
 sg13g2_nand3_1 _3547_ (.B(\counter[29] ),
    .C(_1474_),
    .A(_1472_),
    .Y(_1818_));
 sg13g2_a221oi_1 _3548_ (.B2(_1816_),
    .C1(net63),
    .B1(_1818_),
    .A1(_1472_),
    .Y(_0081_),
    .A2(_1817_));
 sg13g2_inv_1 _3549_ (.Y(_1819_),
    .A(\counter[31] ));
 sg13g2_nand2_1 _3550_ (.Y(_1820_),
    .A(_1494_),
    .B(\counter[30] ));
 sg13g2_o21ai_1 _3551_ (.B1(net74),
    .Y(_1821_),
    .A1(_1819_),
    .A2(_1820_));
 sg13g2_a21oi_1 _3552_ (.A1(_1819_),
    .A2(_1820_),
    .Y(_0082_),
    .B1(_1821_));
 sg13g2_nor2_1 _3553_ (.A(\counter[3] ),
    .B(_1447_),
    .Y(_1822_));
 sg13g2_nor3_1 _3554_ (.A(net62),
    .B(_1822_),
    .C(_1449_),
    .Y(_0083_));
 sg13g2_nor2_1 _3555_ (.A(_1430_),
    .B(_1448_),
    .Y(_1823_));
 sg13g2_nor2_1 _3556_ (.A(\counter[4] ),
    .B(_1449_),
    .Y(_1824_));
 sg13g2_nor3_1 _3557_ (.A(net62),
    .B(_1823_),
    .C(_1824_),
    .Y(_0084_));
 sg13g2_nor2_1 _3558_ (.A(_1451_),
    .B(_1448_),
    .Y(_1825_));
 sg13g2_nor2_1 _3559_ (.A(\counter[5] ),
    .B(_1823_),
    .Y(_1826_));
 sg13g2_nor3_1 _3560_ (.A(net62),
    .B(_1825_),
    .C(_1826_),
    .Y(_0085_));
 sg13g2_nor3_1 _3561_ (.A(_1450_),
    .B(_1451_),
    .C(_1448_),
    .Y(_1827_));
 sg13g2_nor2_1 _3562_ (.A(\counter[6] ),
    .B(_1825_),
    .Y(_1828_));
 sg13g2_nor3_1 _3563_ (.A(net82),
    .B(_1827_),
    .C(_1828_),
    .Y(_0086_));
 sg13g2_o21ai_1 _3564_ (.B1(net74),
    .Y(_1829_),
    .A1(\counter[7] ),
    .A2(_1827_));
 sg13g2_nor2b_1 _3565_ (.A(_1829_),
    .B_N(_1453_),
    .Y(_0087_));
 sg13g2_nand2_1 _3566_ (.Y(_1830_),
    .A(_1455_),
    .B(net74));
 sg13g2_a21oi_1 _3567_ (.A1(_1445_),
    .A2(_1453_),
    .Y(_0088_),
    .B1(_1830_));
 sg13g2_nor2_1 _3568_ (.A(\counter[9] ),
    .B(_1454_),
    .Y(_1831_));
 sg13g2_nor3_1 _3569_ (.A(net82),
    .B(_1831_),
    .C(_1456_),
    .Y(_0089_));
 sg13g2_inv_1 _3570_ (.Y(_1832_),
    .A(_0054_));
 sg13g2_o21ai_1 _3571_ (.B1(net74),
    .Y(_1833_),
    .A1(\frame_counter[0] ),
    .A2(_1683_));
 sg13g2_a21oi_1 _3572_ (.A1(_1832_),
    .A2(_1683_),
    .Y(_0095_),
    .B1(_1833_));
 sg13g2_a21oi_1 _3573_ (.A1(_1683_),
    .A2(\frame_counter[0] ),
    .Y(_1834_),
    .B1(\frame_counter[1] ));
 sg13g2_nor3_1 _3574_ (.A(_1677_),
    .B(_1678_),
    .C(_1684_),
    .Y(_1835_));
 sg13g2_nor3_1 _3575_ (.A(net82),
    .B(_1834_),
    .C(_1835_),
    .Y(_0096_));
 sg13g2_inv_1 _3576_ (.Y(_1836_),
    .A(_0056_));
 sg13g2_o21ai_1 _3577_ (.B1(_1499_),
    .Y(_1837_),
    .A1(\i_project.controller_0.mode_ramp_base[0] ),
    .A2(_1757_));
 sg13g2_a21oi_1 _3578_ (.A1(_1836_),
    .A2(_1757_),
    .Y(_0101_),
    .B1(_1837_));
 sg13g2_buf_1 _3579_ (.A(_1648_),
    .X(_1838_));
 sg13g2_buf_1 _3580_ (.A(\i_project.controller_0.t[9] ),
    .X(_1839_));
 sg13g2_inv_1 _3581_ (.Y(_1840_),
    .A(_1839_));
 sg13g2_buf_8 _3582_ (.A(\i_project.controller_0.mode_ramp_base[5] ),
    .X(_1841_));
 sg13g2_inv_1 _3583_ (.Y(_1842_),
    .A(net73));
 sg13g2_buf_1 _3584_ (.A(\i_project.controller_0.mode_ramp_base[3] ),
    .X(_1843_));
 sg13g2_inv_1 _3585_ (.Y(_1844_),
    .A(_1843_));
 sg13g2_buf_2 _3586_ (.A(\i_project.controller_0.mode_ramp_base[1] ),
    .X(_1845_));
 sg13g2_inv_1 _3587_ (.Y(_1846_),
    .A(_1845_));
 sg13g2_inv_1 _3588_ (.Y(_1847_),
    .A(\i_project.controller_0.mode_ramp_base[0] ));
 sg13g2_nor3_1 _3589_ (.A(_1846_),
    .B(_1847_),
    .C(_1758_),
    .Y(_1848_));
 sg13g2_buf_1 _3590_ (.A(\i_project.controller_0.mode_ramp_base[2] ),
    .X(_1849_));
 sg13g2_nand2_1 _3591_ (.Y(_1850_),
    .A(_1848_),
    .B(net71));
 sg13g2_nor2_1 _3592_ (.A(_1844_),
    .B(_1850_),
    .Y(_1851_));
 sg13g2_buf_1 _3593_ (.A(\i_project.controller_0.mode_ramp_base[4] ),
    .X(_1852_));
 sg13g2_buf_1 _3594_ (.A(_1852_),
    .X(_1853_));
 sg13g2_nand2_1 _3595_ (.Y(_1854_),
    .A(_1851_),
    .B(net61));
 sg13g2_nor2_1 _3596_ (.A(_1842_),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_buf_1 _3597_ (.A(\i_project.controller_0.mode_ramp_base[6] ),
    .X(_1856_));
 sg13g2_buf_8 _3598_ (.A(_1856_),
    .X(_1857_));
 sg13g2_nand2_1 _3599_ (.Y(_1858_),
    .A(_1855_),
    .B(net60));
 sg13g2_buf_1 _3600_ (.A(\i_project.controller_0.mode_ramp_base[7] ),
    .X(_1859_));
 sg13g2_nor2b_1 _3601_ (.A(_1858_),
    .B_N(net70),
    .Y(_1860_));
 sg13g2_buf_2 _3602_ (.A(\i_project.controller_0.t[8] ),
    .X(_1861_));
 sg13g2_nand2_1 _3603_ (.Y(_1862_),
    .A(_1860_),
    .B(_1861_));
 sg13g2_nor2_1 _3604_ (.A(_1840_),
    .B(_1862_),
    .Y(_1863_));
 sg13g2_nor2_1 _3605_ (.A(\i_project.controller_0.t[10] ),
    .B(_1863_),
    .Y(_1864_));
 sg13g2_nand2_1 _3606_ (.Y(_1865_),
    .A(_1863_),
    .B(\i_project.controller_0.t[10] ));
 sg13g2_inv_1 _3607_ (.Y(_1866_),
    .A(_1865_));
 sg13g2_nor3_1 _3608_ (.A(net55),
    .B(_1864_),
    .C(_1866_),
    .Y(_0102_));
 sg13g2_inv_1 _3609_ (.Y(_1867_),
    .A(\i_project.controller_0.t[11] ));
 sg13g2_o21ai_1 _3610_ (.B1(net69),
    .Y(_1868_),
    .A1(_1867_),
    .A2(_1865_));
 sg13g2_a21oi_1 _3611_ (.A1(_1867_),
    .A2(_1865_),
    .Y(_0103_),
    .B1(_1868_));
 sg13g2_a21oi_1 _3612_ (.A1(_1757_),
    .A2(\i_project.controller_0.mode_ramp_base[0] ),
    .Y(_1869_),
    .B1(_1845_));
 sg13g2_nor3_1 _3613_ (.A(net55),
    .B(_1869_),
    .C(_1848_),
    .Y(_0104_));
 sg13g2_nor2_1 _3614_ (.A(net71),
    .B(_1848_),
    .Y(_1870_));
 sg13g2_inv_1 _3615_ (.Y(_1871_),
    .A(_1850_));
 sg13g2_nor3_1 _3616_ (.A(net55),
    .B(_1870_),
    .C(_1871_),
    .Y(_0105_));
 sg13g2_nor2_1 _3617_ (.A(_1843_),
    .B(_1871_),
    .Y(_1872_));
 sg13g2_nor3_1 _3618_ (.A(net55),
    .B(_1851_),
    .C(_1872_),
    .Y(_0106_));
 sg13g2_nor2_1 _3619_ (.A(net61),
    .B(_1851_),
    .Y(_1873_));
 sg13g2_inv_1 _3620_ (.Y(_1874_),
    .A(_1854_));
 sg13g2_nor3_1 _3621_ (.A(net55),
    .B(_1873_),
    .C(_1874_),
    .Y(_0107_));
 sg13g2_nor2_1 _3622_ (.A(net73),
    .B(_1874_),
    .Y(_1875_));
 sg13g2_nor3_1 _3623_ (.A(net55),
    .B(_1855_),
    .C(_1875_),
    .Y(_0108_));
 sg13g2_nor2_1 _3624_ (.A(net60),
    .B(_1855_),
    .Y(_1876_));
 sg13g2_inv_1 _3625_ (.Y(_1877_),
    .A(_1858_));
 sg13g2_nor3_1 _3626_ (.A(net55),
    .B(_1876_),
    .C(_1877_),
    .Y(_0109_));
 sg13g2_nor2_1 _3627_ (.A(net70),
    .B(_1877_),
    .Y(_1878_));
 sg13g2_nor3_1 _3628_ (.A(net55),
    .B(_1860_),
    .C(_1878_),
    .Y(_0110_));
 sg13g2_nor2_1 _3629_ (.A(_1861_),
    .B(_1860_),
    .Y(_1879_));
 sg13g2_inv_1 _3630_ (.Y(_1880_),
    .A(_1862_));
 sg13g2_nor3_1 _3631_ (.A(_1838_),
    .B(_1879_),
    .C(_1880_),
    .Y(_0111_));
 sg13g2_nor2_1 _3632_ (.A(_1839_),
    .B(_1880_),
    .Y(_1881_));
 sg13g2_nor3_1 _3633_ (.A(_1838_),
    .B(_1863_),
    .C(_1881_),
    .Y(_0112_));
 sg13g2_nor2b_1 _3634_ (.A(net63),
    .B_N(\i_project.controller_0.vga_sync.o_vsync ),
    .Y(_0143_));
 sg13g2_nand2_1 _3635_ (.Y(_1882_),
    .A(net83),
    .B(net4));
 sg13g2_inv_1 _3636_ (.Y(_0144_),
    .A(_1882_));
 sg13g2_buf_1 _3637_ (.A(\depth[0] ),
    .X(_1883_));
 sg13g2_buf_1 _3638_ (.A(\depth[1] ),
    .X(_1884_));
 sg13g2_inv_1 _3639_ (.Y(_1885_),
    .A(_1884_));
 sg13g2_inv_1 _3640_ (.Y(_1886_),
    .A(_0044_));
 sg13g2_nor3_1 _3641_ (.A(_1883_),
    .B(_1885_),
    .C(_1886_),
    .Y(_1887_));
 sg13g2_buf_1 _3642_ (.A(_1887_),
    .X(_1888_));
 sg13g2_inv_1 _3643_ (.Y(_1889_),
    .A(_1888_));
 sg13g2_nand2_2 _3644_ (.Y(_1890_),
    .A(_1576_),
    .B(\i_project.controller_0.voffset[0] ));
 sg13g2_nor2_1 _3645_ (.A(net77),
    .B(_1635_),
    .Y(_1891_));
 sg13g2_nand2_1 _3646_ (.Y(_1892_),
    .A(\i_project.controller_0.v[1] ),
    .B(_1635_));
 sg13g2_o21ai_1 _3647_ (.B1(_1892_),
    .Y(_1893_),
    .A1(_1890_),
    .A2(_1891_));
 sg13g2_xnor2_1 _3648_ (.Y(_1894_),
    .A(net76),
    .B(_1637_));
 sg13g2_xnor2_1 _3649_ (.Y(_1895_),
    .A(net75),
    .B(\i_project.controller_0.voffset[3] ));
 sg13g2_nor2_1 _3650_ (.A(_1894_),
    .B(_1895_),
    .Y(_1896_));
 sg13g2_nand2_1 _3651_ (.Y(_1897_),
    .A(_1893_),
    .B(_1896_));
 sg13g2_nand2_1 _3652_ (.Y(_1898_),
    .A(net76),
    .B(_1637_));
 sg13g2_nor2_1 _3653_ (.A(net75),
    .B(\i_project.controller_0.voffset[3] ),
    .Y(_1899_));
 sg13g2_nand2_1 _3654_ (.Y(_1900_),
    .A(net75),
    .B(\i_project.controller_0.voffset[3] ));
 sg13g2_o21ai_1 _3655_ (.B1(_1900_),
    .Y(_1901_),
    .A1(_1898_),
    .A2(_1899_));
 sg13g2_inv_1 _3656_ (.Y(_1902_),
    .A(_1901_));
 sg13g2_nand2_1 _3657_ (.Y(_1903_),
    .A(_1897_),
    .B(_1902_));
 sg13g2_xnor2_1 _3658_ (.Y(_1904_),
    .A(_1569_),
    .B(\i_project.controller_0.voffset[4] ));
 sg13g2_nand2_1 _3659_ (.Y(_1905_),
    .A(_1903_),
    .B(_1904_));
 sg13g2_inv_1 _3660_ (.Y(_1906_),
    .A(_1904_));
 sg13g2_nand3_1 _3661_ (.B(_1902_),
    .C(_1906_),
    .A(_1897_),
    .Y(_1907_));
 sg13g2_nand2_1 _3662_ (.Y(_1908_),
    .A(_1905_),
    .B(_1907_));
 sg13g2_buf_8 _3663_ (.A(_1908_),
    .X(_1909_));
 sg13g2_buf_2 _3664_ (.A(_0042_),
    .X(_1910_));
 sg13g2_inv_1 _3665_ (.Y(_1911_),
    .A(_1910_));
 sg13g2_nand2_1 _3666_ (.Y(_1912_),
    .A(_1909_),
    .B(_1911_));
 sg13g2_nand2_1 _3667_ (.Y(_1913_),
    .A(_1903_),
    .B(_1906_));
 sg13g2_nand3_1 _3668_ (.B(_1902_),
    .C(_1904_),
    .A(_1897_),
    .Y(_1914_));
 sg13g2_nand2_1 _3669_ (.Y(_1915_),
    .A(_1913_),
    .B(_1914_));
 sg13g2_buf_2 _3670_ (.A(_1915_),
    .X(_1916_));
 sg13g2_nand2_1 _3671_ (.Y(_1917_),
    .A(_1916_),
    .B(_1910_));
 sg13g2_nand2_2 _3672_ (.Y(_1918_),
    .A(_1912_),
    .B(_1917_));
 sg13g2_nor2_1 _3673_ (.A(net76),
    .B(_1637_),
    .Y(_1919_));
 sg13g2_o21ai_1 _3674_ (.B1(_1898_),
    .Y(_1920_),
    .A1(_1892_),
    .A2(_1919_));
 sg13g2_nor2_1 _3675_ (.A(_1895_),
    .B(_1904_),
    .Y(_1921_));
 sg13g2_nand2_1 _3676_ (.Y(_1922_),
    .A(_1569_),
    .B(\i_project.controller_0.voffset[4] ));
 sg13g2_nor2_1 _3677_ (.A(_1569_),
    .B(\i_project.controller_0.voffset[4] ),
    .Y(_1923_));
 sg13g2_a21oi_1 _3678_ (.A1(_1922_),
    .A2(_1900_),
    .Y(_1924_),
    .B1(_1923_));
 sg13g2_a21oi_1 _3679_ (.A1(_1920_),
    .A2(_1921_),
    .Y(_1925_),
    .B1(_1924_));
 sg13g2_xnor2_1 _3680_ (.Y(_1926_),
    .A(net77),
    .B(_1635_));
 sg13g2_nor2_1 _3681_ (.A(_1926_),
    .B(_1894_),
    .Y(_1927_));
 sg13g2_inv_2 _3682_ (.Y(_1928_),
    .A(_1890_));
 sg13g2_nand3_1 _3683_ (.B(_1921_),
    .C(_1928_),
    .A(_1927_),
    .Y(_1929_));
 sg13g2_nand2_1 _3684_ (.Y(_1930_),
    .A(_1925_),
    .B(_1929_));
 sg13g2_xnor2_1 _3685_ (.Y(_1931_),
    .A(_1572_),
    .B(\i_project.controller_0.voffset[5] ));
 sg13g2_nand2_1 _3686_ (.Y(_1932_),
    .A(_1930_),
    .B(_1931_));
 sg13g2_inv_2 _3687_ (.Y(_1933_),
    .A(_1931_));
 sg13g2_nand3_1 _3688_ (.B(_1929_),
    .C(_1933_),
    .A(_1925_),
    .Y(_1934_));
 sg13g2_nand2_2 _3689_ (.Y(_1935_),
    .A(_1932_),
    .B(_1934_));
 sg13g2_buf_1 _3690_ (.A(_0041_),
    .X(_1936_));
 sg13g2_inv_1 _3691_ (.Y(_1937_),
    .A(_1936_));
 sg13g2_nand2_1 _3692_ (.Y(_1938_),
    .A(_1935_),
    .B(_1937_));
 sg13g2_nand2_1 _3693_ (.Y(_1939_),
    .A(_1930_),
    .B(_1933_));
 sg13g2_nand3_1 _3694_ (.B(_1929_),
    .C(_1931_),
    .A(_1925_),
    .Y(_1940_));
 sg13g2_nand2_1 _3695_ (.Y(_1941_),
    .A(_1939_),
    .B(_1940_));
 sg13g2_buf_8 _3696_ (.A(_1941_),
    .X(_1942_));
 sg13g2_nand2_1 _3697_ (.Y(_1943_),
    .A(net34),
    .B(_1936_));
 sg13g2_nand2_1 _3698_ (.Y(_1944_),
    .A(_1938_),
    .B(_1943_));
 sg13g2_nor2_1 _3699_ (.A(_1918_),
    .B(_1944_),
    .Y(_1945_));
 sg13g2_inv_1 _3700_ (.Y(_1946_),
    .A(_1891_));
 sg13g2_inv_1 _3701_ (.Y(_1947_),
    .A(_1892_));
 sg13g2_a21oi_1 _3702_ (.A1(_1946_),
    .A2(_1928_),
    .Y(_1948_),
    .B1(_1947_));
 sg13g2_nand2_1 _3703_ (.Y(_1949_),
    .A(_1948_),
    .B(_1894_));
 sg13g2_xor2_1 _3704_ (.B(_1637_),
    .A(net76),
    .X(_1950_));
 sg13g2_nand2_1 _3705_ (.Y(_1951_),
    .A(_1893_),
    .B(_1950_));
 sg13g2_nand2_1 _3706_ (.Y(_1952_),
    .A(_1949_),
    .B(_1951_));
 sg13g2_buf_8 _3707_ (.A(_1952_),
    .X(_1953_));
 sg13g2_xnor2_1 _3708_ (.Y(_1954_),
    .A(net72),
    .B(net38));
 sg13g2_xor2_1 _3709_ (.B(_1635_),
    .A(net77),
    .X(_1955_));
 sg13g2_nand2_1 _3710_ (.Y(_1956_),
    .A(_1955_),
    .B(_1928_));
 sg13g2_nand2_1 _3711_ (.Y(_1957_),
    .A(_1926_),
    .B(_1890_));
 sg13g2_nand2_1 _3712_ (.Y(_1958_),
    .A(_1956_),
    .B(_1957_));
 sg13g2_buf_1 _3713_ (.A(_1958_),
    .X(_1959_));
 sg13g2_xnor2_1 _3714_ (.Y(_1960_),
    .A(net71),
    .B(net44));
 sg13g2_nand2_1 _3715_ (.Y(_1961_),
    .A(_1577_),
    .B(_1602_));
 sg13g2_nand2_1 _3716_ (.Y(_1962_),
    .A(_1961_),
    .B(_1890_));
 sg13g2_buf_2 _3717_ (.A(_1962_),
    .X(_1963_));
 sg13g2_nor2_1 _3718_ (.A(_1846_),
    .B(_1963_),
    .Y(_1964_));
 sg13g2_nand2_1 _3719_ (.Y(_1965_),
    .A(_1960_),
    .B(_1964_));
 sg13g2_inv_1 _3720_ (.Y(_1966_),
    .A(net44));
 sg13g2_inv_1 _3721_ (.Y(_1967_),
    .A(_0020_));
 sg13g2_nand2_1 _3722_ (.Y(_1968_),
    .A(_1966_),
    .B(_1967_));
 sg13g2_nand2_1 _3723_ (.Y(_1969_),
    .A(_1965_),
    .B(_1968_));
 sg13g2_inv_1 _3724_ (.Y(_1970_),
    .A(_1852_));
 sg13g2_nand3_1 _3725_ (.B(_1950_),
    .C(_1928_),
    .A(_1955_),
    .Y(_1971_));
 sg13g2_inv_1 _3726_ (.Y(_1972_),
    .A(_1920_));
 sg13g2_nand2_1 _3727_ (.Y(_1973_),
    .A(_1971_),
    .B(_1972_));
 sg13g2_inv_1 _3728_ (.Y(_1974_),
    .A(_1895_));
 sg13g2_nand2_1 _3729_ (.Y(_1975_),
    .A(_1973_),
    .B(_1974_));
 sg13g2_nand3_1 _3730_ (.B(_1972_),
    .C(_1895_),
    .A(_1971_),
    .Y(_1976_));
 sg13g2_nand2_2 _3731_ (.Y(_1977_),
    .A(_1975_),
    .B(_1976_));
 sg13g2_buf_8 _3732_ (.A(_1977_),
    .X(_1978_));
 sg13g2_xnor2_1 _3733_ (.Y(_1979_),
    .A(_1970_),
    .B(_1978_));
 sg13g2_inv_1 _3734_ (.Y(_1980_),
    .A(_1979_));
 sg13g2_nand4_1 _3735_ (.B(_1954_),
    .C(_1969_),
    .A(_1945_),
    .Y(_1981_),
    .D(_1980_));
 sg13g2_inv_1 _3736_ (.Y(_1982_),
    .A(net38));
 sg13g2_inv_1 _3737_ (.Y(_1983_),
    .A(_0019_));
 sg13g2_nand2_1 _3738_ (.Y(_1984_),
    .A(_1982_),
    .B(_1983_));
 sg13g2_inv_1 _3739_ (.Y(_1985_),
    .A(net33));
 sg13g2_inv_1 _3740_ (.Y(_1986_),
    .A(_0043_));
 sg13g2_nand2_1 _3741_ (.Y(_1987_),
    .A(_1985_),
    .B(_1986_));
 sg13g2_o21ai_1 _3742_ (.B1(_1987_),
    .Y(_1988_),
    .A1(_1984_),
    .A2(_1979_));
 sg13g2_inv_1 _3743_ (.Y(_1989_),
    .A(_1912_));
 sg13g2_inv_1 _3744_ (.Y(_1990_),
    .A(_1938_));
 sg13g2_a21oi_1 _3745_ (.A1(_1943_),
    .A2(_1989_),
    .Y(_1991_),
    .B1(_1990_));
 sg13g2_inv_1 _3746_ (.Y(_1992_),
    .A(_1991_));
 sg13g2_a21oi_1 _3747_ (.A1(_1988_),
    .A2(_1945_),
    .Y(_1993_),
    .B1(_1992_));
 sg13g2_buf_2 _3748_ (.A(_0040_),
    .X(_1994_));
 sg13g2_nor2_1 _3749_ (.A(_1931_),
    .B(_1904_),
    .Y(_1995_));
 sg13g2_nor2_1 _3750_ (.A(_1572_),
    .B(\i_project.controller_0.voffset[5] ),
    .Y(_1996_));
 sg13g2_nand2_1 _3751_ (.Y(_1997_),
    .A(_1572_),
    .B(\i_project.controller_0.voffset[5] ));
 sg13g2_o21ai_1 _3752_ (.B1(_1997_),
    .Y(_1998_),
    .A1(_1922_),
    .A2(_1996_));
 sg13g2_a21oi_1 _3753_ (.A1(_1901_),
    .A2(_1995_),
    .Y(_1999_),
    .B1(_1998_));
 sg13g2_nand3_1 _3754_ (.B(_1896_),
    .C(_1995_),
    .A(_1893_),
    .Y(_2000_));
 sg13g2_nand2_1 _3755_ (.Y(_2001_),
    .A(_1999_),
    .B(_2000_));
 sg13g2_xnor2_1 _3756_ (.Y(_2002_),
    .A(_1570_),
    .B(\i_project.controller_0.voffset[6] ));
 sg13g2_inv_1 _3757_ (.Y(_2003_),
    .A(_2002_));
 sg13g2_nand2_1 _3758_ (.Y(_2004_),
    .A(_2001_),
    .B(_2003_));
 sg13g2_nand3_1 _3759_ (.B(_2000_),
    .C(_2002_),
    .A(_1999_),
    .Y(_2005_));
 sg13g2_nand2_1 _3760_ (.Y(_2006_),
    .A(_2004_),
    .B(_2005_));
 sg13g2_buf_1 _3761_ (.A(_2006_),
    .X(_2007_));
 sg13g2_xnor2_1 _3762_ (.Y(_2008_),
    .A(_1994_),
    .B(net32));
 sg13g2_nor2_1 _3763_ (.A(_1532_),
    .B(_1861_),
    .Y(_2009_));
 sg13g2_nand2_1 _3764_ (.Y(_2010_),
    .A(_1532_),
    .B(_1861_));
 sg13g2_nand2b_1 _3765_ (.Y(_2011_),
    .B(_2010_),
    .A_N(_2009_));
 sg13g2_xnor2_1 _3766_ (.Y(_2012_),
    .A(net64),
    .B(net70));
 sg13g2_nand2_1 _3767_ (.Y(_2013_),
    .A(net79),
    .B(net72));
 sg13g2_xnor2_1 _3768_ (.Y(_2014_),
    .A(_1520_),
    .B(net61));
 sg13g2_nand2_1 _3769_ (.Y(_2015_),
    .A(net68),
    .B(net61));
 sg13g2_o21ai_1 _3770_ (.B1(_2015_),
    .Y(_2016_),
    .A1(_2013_),
    .A2(_2014_));
 sg13g2_xnor2_1 _3771_ (.Y(_2017_),
    .A(_1524_),
    .B(_1856_));
 sg13g2_xnor2_1 _3772_ (.Y(_2018_),
    .A(net65),
    .B(net73));
 sg13g2_nor2_1 _3773_ (.A(_2017_),
    .B(_2018_),
    .Y(_2019_));
 sg13g2_nand2_1 _3774_ (.Y(_2020_),
    .A(net65),
    .B(net73));
 sg13g2_nand2_1 _3775_ (.Y(_2021_),
    .A(net67),
    .B(net60));
 sg13g2_o21ai_1 _3776_ (.B1(_2021_),
    .Y(_2022_),
    .A1(_2020_),
    .A2(_2017_));
 sg13g2_a21oi_1 _3777_ (.A1(_2016_),
    .A2(_2019_),
    .Y(_2023_),
    .B1(_2022_));
 sg13g2_xnor2_1 _3778_ (.Y(_2024_),
    .A(net79),
    .B(net72));
 sg13g2_nor2_1 _3779_ (.A(_2014_),
    .B(_2024_),
    .Y(_2025_));
 sg13g2_nand2_1 _3780_ (.Y(_2026_),
    .A(net80),
    .B(net71));
 sg13g2_inv_1 _3781_ (.Y(_2027_),
    .A(_2026_));
 sg13g2_nand3_1 _3782_ (.B(_2019_),
    .C(_2027_),
    .A(_2025_),
    .Y(_2028_));
 sg13g2_nand2_1 _3783_ (.Y(_2029_),
    .A(_2023_),
    .B(_2028_));
 sg13g2_nand2b_1 _3784_ (.Y(_2030_),
    .B(_2029_),
    .A_N(_2012_));
 sg13g2_nand2_1 _3785_ (.Y(_2031_),
    .A(net64),
    .B(net70));
 sg13g2_nand2_1 _3786_ (.Y(_2032_),
    .A(_2030_),
    .B(_2031_));
 sg13g2_xnor2_1 _3787_ (.Y(_2033_),
    .A(_2011_),
    .B(_2032_));
 sg13g2_xnor2_1 _3788_ (.Y(_2034_),
    .A(_2008_),
    .B(_2033_));
 sg13g2_a21oi_1 _3789_ (.A1(_1981_),
    .A2(_1993_),
    .Y(_2035_),
    .B1(_2034_));
 sg13g2_nand3_1 _3790_ (.B(_1993_),
    .C(_2034_),
    .A(_1981_),
    .Y(_2036_));
 sg13g2_nor3_1 _3791_ (.A(_1616_),
    .B(_1651_),
    .C(_1630_),
    .Y(_2037_));
 sg13g2_buf_2 _3792_ (.A(_2037_),
    .X(_2038_));
 sg13g2_nand2_1 _3793_ (.Y(_2039_),
    .A(_2036_),
    .B(_2038_));
 sg13g2_nor3_2 _3794_ (.A(_1616_),
    .B(_1619_),
    .C(_1630_),
    .Y(_2040_));
 sg13g2_buf_8 _3795_ (.A(_2040_),
    .X(_2041_));
 sg13g2_nor3_1 _3796_ (.A(_1619_),
    .B(_0025_),
    .C(_1653_),
    .Y(_2042_));
 sg13g2_buf_1 _3797_ (.A(_2042_),
    .X(_2043_));
 sg13g2_inv_1 _3798_ (.Y(_2044_),
    .A(_2043_));
 sg13g2_a21oi_1 _3799_ (.A1(_1713_),
    .A2(_1501_),
    .Y(_2045_),
    .B1(_1504_));
 sg13g2_buf_1 _3800_ (.A(_1500_),
    .X(_2046_));
 sg13g2_nand2b_1 _3801_ (.Y(_2047_),
    .B(net59),
    .A_N(_0050_));
 sg13g2_nor2b_1 _3802_ (.A(_2046_),
    .B_N(_0048_),
    .Y(_2048_));
 sg13g2_a21oi_1 _3803_ (.A1(_0023_),
    .A2(_2046_),
    .Y(_2049_),
    .B1(_2048_));
 sg13g2_inv_1 _3804_ (.Y(_2050_),
    .A(_2049_));
 sg13g2_a22oi_1 _3805_ (.Y(_2051_),
    .B1(_1504_),
    .B2(_2050_),
    .A2(_2047_),
    .A1(_2045_));
 sg13g2_buf_1 _3806_ (.A(_2051_),
    .X(_2052_));
 sg13g2_xnor2_1 _3807_ (.Y(_2053_),
    .A(net66),
    .B(net32));
 sg13g2_a21o_1 _3808_ (.A2(net53),
    .A1(_2053_),
    .B1(_2038_),
    .X(_2054_));
 sg13g2_a21oi_1 _3809_ (.A1(net48),
    .A2(_2052_),
    .Y(_2055_),
    .B1(_2054_));
 sg13g2_nor2_1 _3810_ (.A(net57),
    .B(_2055_),
    .Y(_2056_));
 sg13g2_o21ai_1 _3811_ (.B1(_2056_),
    .Y(_2057_),
    .A1(_2035_),
    .A2(_2039_));
 sg13g2_inv_2 _3812_ (.Y(_0146_),
    .A(net32));
 sg13g2_inv_1 _3813_ (.Y(_0147_),
    .A(_2040_));
 sg13g2_nor2_1 _3814_ (.A(_0048_),
    .B(_0147_),
    .Y(_0148_));
 sg13g2_nor3_1 _3815_ (.A(_1619_),
    .B(_1653_),
    .C(_1621_),
    .Y(_0149_));
 sg13g2_buf_8 _3816_ (.A(_0149_),
    .X(_0150_));
 sg13g2_a21oi_1 _3817_ (.A1(_0146_),
    .A2(_0148_),
    .Y(_0151_),
    .B1(net52));
 sg13g2_nand2_1 _3818_ (.Y(_0152_),
    .A(_2057_),
    .B(_0151_));
 sg13g2_nor3_1 _3819_ (.A(_1616_),
    .B(_1651_),
    .C(_1621_),
    .Y(_0153_));
 sg13g2_buf_2 _3820_ (.A(_0153_),
    .X(_0154_));
 sg13g2_inv_1 _3821_ (.Y(_0155_),
    .A(_0154_));
 sg13g2_nor2_1 _3822_ (.A(_1579_),
    .B(_1580_),
    .Y(_0156_));
 sg13g2_inv_1 _3823_ (.Y(_0157_),
    .A(_0156_));
 sg13g2_nand2_1 _3824_ (.Y(_0158_),
    .A(_1712_),
    .B(_1500_));
 sg13g2_o21ai_1 _3825_ (.B1(_0158_),
    .Y(_0159_),
    .A1(_1500_),
    .A2(_0035_));
 sg13g2_nand2_1 _3826_ (.Y(_0160_),
    .A(_0159_),
    .B(net81));
 sg13g2_a21oi_1 _3827_ (.A1(_1500_),
    .A2(_0036_),
    .Y(_0161_),
    .B1(\i_project.controller_0.divider[1] ));
 sg13g2_o21ai_1 _3828_ (.B1(_0161_),
    .Y(_0162_),
    .A1(_1500_),
    .A2(_1708_));
 sg13g2_nand2_1 _3829_ (.Y(_0163_),
    .A(_0160_),
    .B(_0162_));
 sg13g2_inv_1 _3830_ (.Y(_0164_),
    .A(_0163_));
 sg13g2_nand2_1 _3831_ (.Y(_0165_),
    .A(_0157_),
    .B(_1708_));
 sg13g2_o21ai_1 _3832_ (.B1(_0165_),
    .Y(_0166_),
    .A1(_0157_),
    .A2(_0164_));
 sg13g2_buf_2 _3833_ (.A(_0166_),
    .X(_0167_));
 sg13g2_inv_1 _3834_ (.Y(_0168_),
    .A(_0167_));
 sg13g2_buf_1 _3835_ (.A(_0168_),
    .X(_0169_));
 sg13g2_inv_1 _3836_ (.Y(_0170_),
    .A(net52));
 sg13g2_a21oi_1 _3837_ (.A1(_0146_),
    .A2(_0168_),
    .Y(_0171_),
    .B1(_0170_));
 sg13g2_o21ai_1 _3838_ (.B1(_0171_),
    .Y(_0172_),
    .A1(_0146_),
    .A2(net27));
 sg13g2_nand3_1 _3839_ (.B(_0155_),
    .C(_0172_),
    .A(_0152_),
    .Y(_0173_));
 sg13g2_nand2_2 _3840_ (.Y(_0174_),
    .A(_1560_),
    .B(_1545_));
 sg13g2_inv_1 _3841_ (.Y(_0175_),
    .A(_0174_));
 sg13g2_buf_8 _3842_ (.A(_0175_),
    .X(_0176_));
 sg13g2_a21oi_1 _3843_ (.A1(_0146_),
    .A2(_0154_),
    .Y(_0177_),
    .B1(net37));
 sg13g2_nand2_1 _3844_ (.Y(_0178_),
    .A(_0173_),
    .B(_0177_));
 sg13g2_nand2_1 _3845_ (.Y(_0179_),
    .A(_1567_),
    .B(\i_project.controller_0.voffset[7] ));
 sg13g2_nand2_1 _3846_ (.Y(_0180_),
    .A(_1933_),
    .B(_2003_));
 sg13g2_nor2b_1 _3847_ (.A(_0180_),
    .B_N(_1921_),
    .Y(_0181_));
 sg13g2_nand2_1 _3848_ (.Y(_0182_),
    .A(_1973_),
    .B(_0181_));
 sg13g2_nand2_1 _3849_ (.Y(_0183_),
    .A(_1570_),
    .B(\i_project.controller_0.voffset[6] ));
 sg13g2_o21ai_1 _3850_ (.B1(_0183_),
    .Y(_0184_),
    .A1(_1997_),
    .A2(_2002_));
 sg13g2_nor2b_1 _3851_ (.A(_0180_),
    .B_N(_1924_),
    .Y(_0185_));
 sg13g2_nor2_1 _3852_ (.A(_0184_),
    .B(_0185_),
    .Y(_0186_));
 sg13g2_nand2_1 _3853_ (.Y(_0187_),
    .A(_0182_),
    .B(_0186_));
 sg13g2_nor2_1 _3854_ (.A(_1567_),
    .B(\i_project.controller_0.voffset[7] ),
    .Y(_0188_));
 sg13g2_nor2b_1 _3855_ (.A(_0188_),
    .B_N(_0179_),
    .Y(_0189_));
 sg13g2_nand3_1 _3856_ (.B(_1579_),
    .C(_0189_),
    .A(_0187_),
    .Y(_0190_));
 sg13g2_o21ai_1 _3857_ (.B1(_0190_),
    .Y(_0191_),
    .A1(_0032_),
    .A2(_0179_));
 sg13g2_nand2b_1 _3858_ (.Y(_0192_),
    .B(_1580_),
    .A_N(_0191_));
 sg13g2_inv_1 _3859_ (.Y(_0193_),
    .A(net80));
 sg13g2_nand2_1 _3860_ (.Y(_0194_),
    .A(_0191_),
    .B(_1777_));
 sg13g2_nand3_1 _3861_ (.B(_0193_),
    .C(_0194_),
    .A(_0192_),
    .Y(_0195_));
 sg13g2_nand2_1 _3862_ (.Y(_0196_),
    .A(_0183_),
    .B(_0179_));
 sg13g2_inv_1 _3863_ (.Y(_0197_),
    .A(_0196_));
 sg13g2_a21oi_1 _3864_ (.A1(_2004_),
    .A2(_0197_),
    .Y(_0198_),
    .B1(_0188_));
 sg13g2_xnor2_1 _3865_ (.Y(_0199_),
    .A(_1579_),
    .B(_0198_));
 sg13g2_nand2_1 _3866_ (.Y(_0200_),
    .A(_0199_),
    .B(net80));
 sg13g2_nor2_1 _3867_ (.A(_0036_),
    .B(_0035_),
    .Y(_0201_));
 sg13g2_nand3_1 _3868_ (.B(_0200_),
    .C(_0201_),
    .A(_0195_),
    .Y(_0202_));
 sg13g2_nand2_1 _3869_ (.Y(_0203_),
    .A(_0202_),
    .B(_1519_));
 sg13g2_nor2_1 _3870_ (.A(_1515_),
    .B(_0193_),
    .Y(_0204_));
 sg13g2_inv_2 _3871_ (.Y(_0205_),
    .A(_1963_));
 sg13g2_nor2_1 _3872_ (.A(_1710_),
    .B(_0205_),
    .Y(_0206_));
 sg13g2_a221oi_1 _3873_ (.B2(_0204_),
    .C1(_0206_),
    .B1(_1953_),
    .A1(_1517_),
    .Y(_0207_),
    .A2(_1959_));
 sg13g2_o21ai_1 _3874_ (.B1(_0207_),
    .Y(_0208_),
    .A1(_1542_),
    .A2(_1985_));
 sg13g2_a22oi_1 _3875_ (.Y(_0209_),
    .B1(_1517_),
    .B2(_1942_),
    .A2(_1916_),
    .A1(_1711_));
 sg13g2_nand2_1 _3876_ (.Y(_0210_),
    .A(net32),
    .B(_0204_));
 sg13g2_nand3b_1 _3877_ (.B(_0182_),
    .C(_0186_),
    .Y(_0211_),
    .A_N(_0189_));
 sg13g2_nand2_1 _3878_ (.Y(_0212_),
    .A(_0187_),
    .B(_0189_));
 sg13g2_nand2_1 _3879_ (.Y(_0213_),
    .A(_0211_),
    .B(_0212_));
 sg13g2_buf_8 _3880_ (.A(_0213_),
    .X(_0214_));
 sg13g2_nand2_1 _3881_ (.Y(_0215_),
    .A(net26),
    .B(_1541_));
 sg13g2_nand3_1 _3882_ (.B(_0210_),
    .C(_0215_),
    .A(_0209_),
    .Y(_0216_));
 sg13g2_a22oi_1 _3883_ (.Y(_0217_),
    .B1(_1604_),
    .B2(_0216_),
    .A2(_0208_),
    .A1(_1562_));
 sg13g2_nand2_1 _3884_ (.Y(_0218_),
    .A(_0203_),
    .B(_0217_));
 sg13g2_nand2_1 _3885_ (.Y(_0219_),
    .A(_0218_),
    .B(_0175_));
 sg13g2_buf_8 _3886_ (.A(_0219_),
    .X(_0220_));
 sg13g2_inv_4 _3887_ (.A(_0220_),
    .Y(_0221_));
 sg13g2_nor2_1 _3888_ (.A(_1623_),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_buf_8 _3889_ (.A(_0222_),
    .X(_0223_));
 sg13g2_nand2_1 _3890_ (.Y(_0224_),
    .A(_0178_),
    .B(_0223_));
 sg13g2_inv_4 _3891_ (.A(_1623_),
    .Y(_0225_));
 sg13g2_nor2_1 _3892_ (.A(_0049_),
    .B(_0225_),
    .Y(_0226_));
 sg13g2_inv_2 _3893_ (.Y(_0227_),
    .A(_0226_));
 sg13g2_nand2_1 _3894_ (.Y(_0228_),
    .A(_0224_),
    .B(_0227_));
 sg13g2_nand3_1 _3895_ (.B(_1744_),
    .C(_1573_),
    .A(_1571_),
    .Y(_0229_));
 sg13g2_nand2_1 _3896_ (.Y(_0230_),
    .A(_1597_),
    .B(_1744_));
 sg13g2_nor2b_1 _3897_ (.A(_0031_),
    .B_N(_1570_),
    .Y(_0231_));
 sg13g2_a21oi_1 _3898_ (.A1(_0231_),
    .A2(_1590_),
    .Y(_0232_),
    .B1(_1580_));
 sg13g2_o21ai_1 _3899_ (.B1(_0232_),
    .Y(_0233_),
    .A1(_0230_),
    .A2(_1592_));
 sg13g2_a22oi_1 _3900_ (.Y(_0234_),
    .B1(_1511_),
    .B2(_0233_),
    .A2(_0229_),
    .A1(_1600_));
 sg13g2_nand2_1 _3901_ (.Y(_0235_),
    .A(_1614_),
    .B(_0234_));
 sg13g2_nand2_1 _3902_ (.Y(_0236_),
    .A(_0235_),
    .B(_0225_));
 sg13g2_buf_2 _3903_ (.A(_0236_),
    .X(_0237_));
 sg13g2_nand2_1 _3904_ (.Y(_0238_),
    .A(_0228_),
    .B(_0237_));
 sg13g2_inv_1 _3905_ (.Y(_0239_),
    .A(_1883_));
 sg13g2_a21oi_1 _3906_ (.A1(_1885_),
    .A2(_0239_),
    .Y(_0240_),
    .B1(_1886_));
 sg13g2_a21oi_1 _3907_ (.A1(_1884_),
    .A2(_1883_),
    .Y(_0241_),
    .B1(\depth[2] ));
 sg13g2_nor3_2 _3908_ (.A(_1885_),
    .B(_0239_),
    .C(_1886_),
    .Y(_0242_));
 sg13g2_nor2_1 _3909_ (.A(_0241_),
    .B(_0242_),
    .Y(_0243_));
 sg13g2_nor2_1 _3910_ (.A(_0240_),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_buf_2 _3911_ (.A(_0244_),
    .X(_0245_));
 sg13g2_inv_1 _3912_ (.Y(_0246_),
    .A(_0245_));
 sg13g2_buf_1 _3913_ (.A(_0246_),
    .X(_0247_));
 sg13g2_o21ai_1 _3914_ (.B1(net31),
    .Y(_0248_),
    .A1(_1889_),
    .A2(_0238_));
 sg13g2_inv_1 _3915_ (.Y(_0249_),
    .A(\depth[2] ));
 sg13g2_nor3_1 _3916_ (.A(_1884_),
    .B(_0239_),
    .C(_0249_),
    .Y(_0250_));
 sg13g2_inv_1 _3917_ (.Y(_0251_),
    .A(_0250_));
 sg13g2_o21ai_1 _3918_ (.B1(_1912_),
    .Y(_0252_),
    .A1(_1987_),
    .A2(_1918_));
 sg13g2_inv_1 _3919_ (.Y(_0253_),
    .A(_1857_));
 sg13g2_xnor2_1 _3920_ (.Y(_0254_),
    .A(_0253_),
    .B(net34));
 sg13g2_nor2_1 _3921_ (.A(_0254_),
    .B(_2008_),
    .Y(_0255_));
 sg13g2_inv_1 _3922_ (.Y(_0256_),
    .A(_1994_));
 sg13g2_nand2_1 _3923_ (.Y(_0257_),
    .A(_0146_),
    .B(_0256_));
 sg13g2_o21ai_1 _3924_ (.B1(_0257_),
    .Y(_0258_),
    .A1(_1938_),
    .A2(_2008_));
 sg13g2_a21oi_1 _3925_ (.A1(_0252_),
    .A2(_0255_),
    .Y(_0259_),
    .B1(_0258_));
 sg13g2_nand2_1 _3926_ (.Y(_0260_),
    .A(_1969_),
    .B(_1954_));
 sg13g2_nand2_1 _3927_ (.Y(_0261_),
    .A(_0260_),
    .B(_1984_));
 sg13g2_nor2_1 _3928_ (.A(_1979_),
    .B(_1918_),
    .Y(_0262_));
 sg13g2_nand3_1 _3929_ (.B(_0261_),
    .C(_0262_),
    .A(_0255_),
    .Y(_0263_));
 sg13g2_inv_1 _3930_ (.Y(_0264_),
    .A(_0039_));
 sg13g2_xnor2_1 _3931_ (.Y(_0265_),
    .A(_0264_),
    .B(net26));
 sg13g2_xor2_1 _3932_ (.B(_1839_),
    .A(net78),
    .X(_0266_));
 sg13g2_a21o_1 _3933_ (.A2(_2025_),
    .A1(_2027_),
    .B1(_2016_),
    .X(_0267_));
 sg13g2_nor2_1 _3934_ (.A(_2012_),
    .B(_2011_),
    .Y(_0268_));
 sg13g2_nand3_1 _3935_ (.B(_2019_),
    .C(_0268_),
    .A(_0267_),
    .Y(_0269_));
 sg13g2_o21ai_1 _3936_ (.B1(_2010_),
    .Y(_0270_),
    .A1(_2031_),
    .A2(_2009_));
 sg13g2_a21oi_1 _3937_ (.A1(_2022_),
    .A2(_0268_),
    .Y(_0271_),
    .B1(_0270_));
 sg13g2_nand2_1 _3938_ (.Y(_0272_),
    .A(_0269_),
    .B(_0271_));
 sg13g2_xnor2_1 _3939_ (.Y(_0273_),
    .A(_0266_),
    .B(_0272_));
 sg13g2_xnor2_1 _3940_ (.Y(_0274_),
    .A(_0265_),
    .B(_0273_));
 sg13g2_a21oi_1 _3941_ (.A1(_0259_),
    .A2(_0263_),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_nand3_1 _3942_ (.B(_0263_),
    .C(_0274_),
    .A(_0259_),
    .Y(_0276_));
 sg13g2_nand2_1 _3943_ (.Y(_0277_),
    .A(_0276_),
    .B(_2038_));
 sg13g2_nand2_1 _3944_ (.Y(_0278_),
    .A(_0026_),
    .B(_1500_));
 sg13g2_inv_1 _3945_ (.Y(_0279_),
    .A(_0278_));
 sg13g2_a21oi_1 _3946_ (.A1(_0023_),
    .A2(_1501_),
    .Y(_0280_),
    .B1(_0279_));
 sg13g2_o21ai_1 _3947_ (.B1(net81),
    .Y(_0281_),
    .A1(net59),
    .A2(_1544_));
 sg13g2_o21ai_1 _3948_ (.B1(_0281_),
    .Y(_0282_),
    .A1(net81),
    .A2(_0280_));
 sg13g2_inv_1 _3949_ (.Y(_0283_),
    .A(_0282_));
 sg13g2_xnor2_1 _3950_ (.Y(_0284_),
    .A(_1534_),
    .B(net26));
 sg13g2_a21o_1 _3951_ (.A2(net53),
    .A1(_0284_),
    .B1(_2038_),
    .X(_0285_));
 sg13g2_a21oi_1 _3952_ (.A1(net48),
    .A2(_0283_),
    .Y(_0286_),
    .B1(_0285_));
 sg13g2_nor2_1 _3953_ (.A(net57),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_o21ai_1 _3954_ (.B1(_0287_),
    .Y(_0288_),
    .A1(_0275_),
    .A2(_0277_));
 sg13g2_inv_1 _3955_ (.Y(_0289_),
    .A(net26));
 sg13g2_nor2_1 _3956_ (.A(_0023_),
    .B(_0147_),
    .Y(_0290_));
 sg13g2_a21oi_1 _3957_ (.A1(_0289_),
    .A2(_0290_),
    .Y(_0291_),
    .B1(net52));
 sg13g2_nand2_1 _3958_ (.Y(_0292_),
    .A(_0288_),
    .B(_0291_));
 sg13g2_xnor2_1 _3959_ (.Y(_0293_),
    .A(_0168_),
    .B(_0214_));
 sg13g2_a21oi_1 _3960_ (.A1(_0293_),
    .A2(_0150_),
    .Y(_0294_),
    .B1(_0154_));
 sg13g2_nand2_1 _3961_ (.Y(_0295_),
    .A(_0292_),
    .B(_0294_));
 sg13g2_a21oi_1 _3962_ (.A1(_0289_),
    .A2(_0154_),
    .Y(_0296_),
    .B1(_0176_));
 sg13g2_nand2_1 _3963_ (.Y(_0297_),
    .A(_0295_),
    .B(_0296_));
 sg13g2_nand2_1 _3964_ (.Y(_0298_),
    .A(_0297_),
    .B(_0220_));
 sg13g2_inv_2 _3965_ (.Y(_0299_),
    .A(_0237_));
 sg13g2_a21oi_2 _3966_ (.B1(_0299_),
    .Y(_0300_),
    .A2(_1623_),
    .A1(_0034_));
 sg13g2_inv_1 _3967_ (.Y(_0301_),
    .A(_0300_));
 sg13g2_a21oi_1 _3968_ (.A1(_0298_),
    .A2(_0225_),
    .Y(_0302_),
    .B1(_0301_));
 sg13g2_buf_8 _3969_ (.A(_0302_),
    .X(_0303_));
 sg13g2_nor3_1 _3970_ (.A(_1883_),
    .B(_1885_),
    .C(_0249_),
    .Y(_0304_));
 sg13g2_nand2_1 _3971_ (.Y(_0305_),
    .A(net22),
    .B(_0304_));
 sg13g2_o21ai_1 _3972_ (.B1(_0305_),
    .Y(_0306_),
    .A1(_0251_),
    .A2(_0238_));
 sg13g2_nor3_1 _3973_ (.A(_1884_),
    .B(_0239_),
    .C(_1886_),
    .Y(_0307_));
 sg13g2_buf_1 _3974_ (.A(_0307_),
    .X(_0308_));
 sg13g2_nand3_1 _3975_ (.B(_0237_),
    .C(net51),
    .A(_0228_),
    .Y(_0309_));
 sg13g2_buf_1 _3976_ (.A(_0147_),
    .X(_0310_));
 sg13g2_a21oi_1 _3977_ (.A1(_0205_),
    .A2(_1708_),
    .Y(_0311_),
    .B1(net50));
 sg13g2_inv_1 _3978_ (.Y(_0312_),
    .A(net71));
 sg13g2_xnor2_1 _3979_ (.Y(_0313_),
    .A(net80),
    .B(_1845_));
 sg13g2_xnor2_1 _3980_ (.Y(_0314_),
    .A(_0312_),
    .B(_0313_));
 sg13g2_buf_1 _3981_ (.A(_2038_),
    .X(_0315_));
 sg13g2_inv_1 _3982_ (.Y(_0316_),
    .A(net47));
 sg13g2_a21oi_1 _3983_ (.A1(_0314_),
    .A2(_0205_),
    .Y(_0317_),
    .B1(_0316_));
 sg13g2_o21ai_1 _3984_ (.B1(_0317_),
    .Y(_0318_),
    .A1(_0205_),
    .A2(_0314_));
 sg13g2_nor2_1 _3985_ (.A(net53),
    .B(_0164_),
    .Y(_0319_));
 sg13g2_xnor2_1 _3986_ (.Y(_0320_),
    .A(_1514_),
    .B(_1963_));
 sg13g2_inv_1 _3987_ (.Y(_0321_),
    .A(_0320_));
 sg13g2_o21ai_1 _3988_ (.B1(_0316_),
    .Y(_0322_),
    .A1(net48),
    .A2(_0321_));
 sg13g2_buf_1 _3989_ (.A(net57),
    .X(_0323_));
 sg13g2_a21o_1 _3990_ (.A2(_0322_),
    .A1(_0318_),
    .B1(net49),
    .X(_0324_));
 sg13g2_a21oi_1 _3991_ (.A1(_0318_),
    .A2(_0319_),
    .Y(_0325_),
    .B1(_0324_));
 sg13g2_buf_1 _3992_ (.A(_0170_),
    .X(_0326_));
 sg13g2_buf_1 _3993_ (.A(net43),
    .X(_0327_));
 sg13g2_o21ai_1 _3994_ (.B1(net36),
    .Y(_0328_),
    .A1(_0311_),
    .A2(_0325_));
 sg13g2_buf_1 _3995_ (.A(_0155_),
    .X(_0329_));
 sg13g2_a21oi_1 _3996_ (.A1(net27),
    .A2(_0205_),
    .Y(_0330_),
    .B1(_0327_));
 sg13g2_o21ai_1 _3997_ (.B1(_0330_),
    .Y(_0331_),
    .A1(_0205_),
    .A2(net27));
 sg13g2_nand3_1 _3998_ (.B(_0329_),
    .C(_0331_),
    .A(_0328_),
    .Y(_0332_));
 sg13g2_buf_8 _3999_ (.A(_0154_),
    .X(_0333_));
 sg13g2_buf_1 _4000_ (.A(net46),
    .X(_0334_));
 sg13g2_buf_1 _4001_ (.A(net41),
    .X(_0335_));
 sg13g2_nand2_1 _4002_ (.Y(_0336_),
    .A(_0205_),
    .B(_0335_));
 sg13g2_nand3_1 _4003_ (.B(_0174_),
    .C(_0336_),
    .A(_0332_),
    .Y(_0337_));
 sg13g2_nor2_1 _4004_ (.A(_1623_),
    .B(_0235_),
    .Y(_0338_));
 sg13g2_nor3_1 _4005_ (.A(_0044_),
    .B(_1885_),
    .C(_0239_),
    .Y(_0339_));
 sg13g2_nand3_1 _4006_ (.B(_0338_),
    .C(_0339_),
    .A(_0220_),
    .Y(_0340_));
 sg13g2_inv_1 _4007_ (.Y(_0341_),
    .A(_0340_));
 sg13g2_nor3_1 _4008_ (.A(_1884_),
    .B(_1883_),
    .C(_0249_),
    .Y(_0342_));
 sg13g2_buf_2 _4009_ (.A(_0342_),
    .X(_0343_));
 sg13g2_xor2_1 _4010_ (.B(_2029_),
    .A(_2012_),
    .X(_0344_));
 sg13g2_xnor2_1 _4011_ (.Y(_0345_),
    .A(_0344_),
    .B(_1944_));
 sg13g2_inv_1 _4012_ (.Y(_0346_),
    .A(_1954_));
 sg13g2_o21ai_1 _4013_ (.B1(_1984_),
    .Y(_0347_),
    .A1(_1968_),
    .A2(_0346_));
 sg13g2_a21oi_1 _4014_ (.A1(_0347_),
    .A2(_0262_),
    .Y(_0348_),
    .B1(_0252_));
 sg13g2_nand4_1 _4015_ (.B(_1954_),
    .C(_1964_),
    .A(_0262_),
    .Y(_0349_),
    .D(_1960_));
 sg13g2_nand3b_1 _4016_ (.B(_0348_),
    .C(_0349_),
    .Y(_0350_),
    .A_N(_0345_));
 sg13g2_nand2_1 _4017_ (.Y(_0351_),
    .A(_0348_),
    .B(_0349_));
 sg13g2_nand2_1 _4018_ (.Y(_0352_),
    .A(_0351_),
    .B(_0345_));
 sg13g2_nand3_1 _4019_ (.B(_0352_),
    .C(net47),
    .A(_0350_),
    .Y(_0353_));
 sg13g2_xnor2_1 _4020_ (.Y(_0354_),
    .A(_1549_),
    .B(net34));
 sg13g2_a21oi_1 _4021_ (.A1(_0354_),
    .A2(net53),
    .Y(_0355_),
    .B1(_2038_));
 sg13g2_nor2b_1 _4022_ (.A(net59),
    .B_N(_0047_),
    .Y(_0356_));
 sg13g2_a21oi_1 _4023_ (.A1(net59),
    .A2(_0048_),
    .Y(_0357_),
    .B1(_0356_));
 sg13g2_mux2_1 _4024_ (.A0(_0357_),
    .A1(_0280_),
    .S(net81),
    .X(_0358_));
 sg13g2_buf_1 _4025_ (.A(_0358_),
    .X(_0359_));
 sg13g2_nand3_1 _4026_ (.B(_0147_),
    .C(_2044_),
    .A(_0359_),
    .Y(_0360_));
 sg13g2_nand2_1 _4027_ (.Y(_0361_),
    .A(_0355_),
    .B(_0360_));
 sg13g2_nand2_1 _4028_ (.Y(_0362_),
    .A(_0353_),
    .B(_0361_));
 sg13g2_nor2_1 _4029_ (.A(_0047_),
    .B(net50),
    .Y(_0363_));
 sg13g2_a21oi_1 _4030_ (.A1(_1935_),
    .A2(_0363_),
    .Y(_0364_),
    .B1(net52));
 sg13g2_nand2_1 _4031_ (.Y(_0365_),
    .A(_0362_),
    .B(_0364_));
 sg13g2_xnor2_1 _4032_ (.Y(_0366_),
    .A(net27),
    .B(_1942_));
 sg13g2_buf_1 _4033_ (.A(net52),
    .X(_0367_));
 sg13g2_a21oi_1 _4034_ (.A1(_0366_),
    .A2(_0367_),
    .Y(_0368_),
    .B1(_0154_));
 sg13g2_nand2_1 _4035_ (.Y(_0369_),
    .A(_0365_),
    .B(_0368_));
 sg13g2_a21oi_1 _4036_ (.A1(_1935_),
    .A2(net46),
    .Y(_0370_),
    .B1(net37));
 sg13g2_nand2_1 _4037_ (.Y(_0371_),
    .A(_0369_),
    .B(_0370_));
 sg13g2_nand2_1 _4038_ (.Y(_0372_),
    .A(_0371_),
    .B(_0223_));
 sg13g2_nand2b_1 _4039_ (.Y(_0373_),
    .B(_1623_),
    .A_N(_0017_));
 sg13g2_buf_1 _4040_ (.A(_0373_),
    .X(_0374_));
 sg13g2_a21oi_1 _4041_ (.A1(_0372_),
    .A2(_0374_),
    .Y(_0375_),
    .B1(_0299_));
 sg13g2_a22oi_1 _4042_ (.Y(_0376_),
    .B1(_0343_),
    .B2(_0375_),
    .A2(_0341_),
    .A1(_0337_));
 sg13g2_nand2b_1 _4043_ (.Y(_0377_),
    .B(_0323_),
    .A_N(_0046_));
 sg13g2_o21ai_1 _4044_ (.B1(net36),
    .Y(_0378_),
    .A1(_0377_),
    .A2(_1916_));
 sg13g2_xnor2_1 _4045_ (.Y(_0379_),
    .A(_1525_),
    .B(_1909_));
 sg13g2_inv_1 _4046_ (.Y(_0380_),
    .A(_0379_));
 sg13g2_a21oi_1 _4047_ (.A1(_0380_),
    .A2(net53),
    .Y(_0381_),
    .B1(net47));
 sg13g2_nand2_1 _4048_ (.Y(_0382_),
    .A(net59),
    .B(_0047_));
 sg13g2_inv_1 _4049_ (.Y(_0383_),
    .A(_0382_));
 sg13g2_a21oi_1 _4050_ (.A1(_1501_),
    .A2(_0046_),
    .Y(_0384_),
    .B1(_0383_));
 sg13g2_nor2_1 _4051_ (.A(net81),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_a21oi_2 _4052_ (.B1(_0385_),
    .Y(_0386_),
    .A2(_2050_),
    .A1(_1503_));
 sg13g2_nand3_1 _4053_ (.B(_0310_),
    .C(net48),
    .A(_0386_),
    .Y(_0387_));
 sg13g2_buf_1 _4054_ (.A(net47),
    .X(_0388_));
 sg13g2_nand2b_1 _4055_ (.Y(_0389_),
    .B(_0267_),
    .A_N(_2018_));
 sg13g2_nand2_1 _4056_ (.Y(_0390_),
    .A(_0389_),
    .B(_2020_));
 sg13g2_xnor2_1 _4057_ (.Y(_0391_),
    .A(_2017_),
    .B(_0390_));
 sg13g2_a22oi_1 _4058_ (.Y(_0392_),
    .B1(_1980_),
    .B2(_0261_),
    .A2(_1985_),
    .A1(_1986_));
 sg13g2_xor2_1 _4059_ (.B(_0392_),
    .A(_1918_),
    .X(_0393_));
 sg13g2_xnor2_1 _4060_ (.Y(_0394_),
    .A(_0391_),
    .B(_0393_));
 sg13g2_a22oi_1 _4061_ (.Y(_0395_),
    .B1(_0388_),
    .B2(_0394_),
    .A2(_0387_),
    .A1(_0381_));
 sg13g2_buf_1 _4062_ (.A(_0167_),
    .X(_0396_));
 sg13g2_buf_1 _4063_ (.A(net29),
    .X(_0397_));
 sg13g2_xnor2_1 _4064_ (.Y(_0398_),
    .A(_1909_),
    .B(net25));
 sg13g2_buf_1 _4065_ (.A(net45),
    .X(_0399_));
 sg13g2_a21oi_1 _4066_ (.A1(_0398_),
    .A2(_0399_),
    .Y(_0400_),
    .B1(net35));
 sg13g2_o21ai_1 _4067_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_0378_),
    .A2(_0395_));
 sg13g2_buf_1 _4068_ (.A(net37),
    .X(_0402_));
 sg13g2_a21oi_1 _4069_ (.A1(_1909_),
    .A2(_0335_),
    .Y(_0403_),
    .B1(net30));
 sg13g2_inv_2 _4070_ (.Y(_0404_),
    .A(_0223_));
 sg13g2_a21oi_1 _4071_ (.A1(_0401_),
    .A2(_0403_),
    .Y(_0405_),
    .B1(_0404_));
 sg13g2_nand2b_1 _4072_ (.Y(_0406_),
    .B(_1624_),
    .A_N(_0045_));
 sg13g2_nand2b_1 _4073_ (.Y(_0407_),
    .B(_0406_),
    .A_N(_0405_));
 sg13g2_inv_1 _4074_ (.Y(_0408_),
    .A(_0242_));
 sg13g2_nor2_1 _4075_ (.A(_0408_),
    .B(_0299_),
    .Y(_0409_));
 sg13g2_buf_1 _4076_ (.A(_0409_),
    .X(_0410_));
 sg13g2_nand2_1 _4077_ (.Y(_0411_),
    .A(_0407_),
    .B(net23));
 sg13g2_nand3_1 _4078_ (.B(_0376_),
    .C(_0411_),
    .A(_0309_),
    .Y(_0412_));
 sg13g2_nor3_1 _4079_ (.A(_0248_),
    .B(_0306_),
    .C(_0412_),
    .Y(_0413_));
 sg13g2_buf_1 _4080_ (.A(_0237_),
    .X(_0414_));
 sg13g2_nand3_1 _4081_ (.B(net24),
    .C(_0343_),
    .A(_0228_),
    .Y(_0415_));
 sg13g2_nor3_1 _4082_ (.A(_0308_),
    .B(net54),
    .C(_0250_),
    .Y(_0416_));
 sg13g2_inv_1 _4083_ (.Y(_0417_),
    .A(_0416_));
 sg13g2_nand2_1 _4084_ (.Y(_0418_),
    .A(net22),
    .B(_0417_));
 sg13g2_nand2_1 _4085_ (.Y(_0419_),
    .A(_0372_),
    .B(_0374_));
 sg13g2_nor2_1 _4086_ (.A(_0339_),
    .B(_0304_),
    .Y(_0420_));
 sg13g2_nor2_1 _4087_ (.A(_0420_),
    .B(_0299_),
    .Y(_0421_));
 sg13g2_nor2b_1 _4088_ (.A(_0404_),
    .B_N(_0421_),
    .Y(_0422_));
 sg13g2_xnor2_1 _4089_ (.Y(_0423_),
    .A(_1516_),
    .B(net44));
 sg13g2_inv_1 _4090_ (.Y(_0424_),
    .A(_0423_));
 sg13g2_a21oi_1 _4091_ (.A1(_0424_),
    .A2(net53),
    .Y(_0425_),
    .B1(net47));
 sg13g2_nand2_1 _4092_ (.Y(_0426_),
    .A(_1501_),
    .B(_0036_));
 sg13g2_a21oi_1 _4093_ (.A1(net59),
    .A2(_0035_),
    .Y(_0427_),
    .B1(net81));
 sg13g2_nand2_1 _4094_ (.Y(_0428_),
    .A(net59),
    .B(_0046_));
 sg13g2_o21ai_1 _4095_ (.B1(_0428_),
    .Y(_0429_),
    .A1(net59),
    .A2(_1712_));
 sg13g2_inv_1 _4096_ (.Y(_0430_),
    .A(_0429_));
 sg13g2_a22oi_1 _4097_ (.Y(_0431_),
    .B1(net81),
    .B2(_0430_),
    .A2(_0427_),
    .A1(_0426_));
 sg13g2_inv_1 _4098_ (.Y(_0432_),
    .A(_0431_));
 sg13g2_nand2_1 _4099_ (.Y(_0433_),
    .A(_0432_),
    .B(net48));
 sg13g2_xnor2_1 _4100_ (.Y(_0434_),
    .A(_2027_),
    .B(_2024_));
 sg13g2_xor2_1 _4101_ (.B(_1960_),
    .A(_1964_),
    .X(_0435_));
 sg13g2_xnor2_1 _4102_ (.Y(_0436_),
    .A(_0434_),
    .B(_0435_));
 sg13g2_a22oi_1 _4103_ (.Y(_0437_),
    .B1(net40),
    .B2(_0436_),
    .A2(_0433_),
    .A1(_0425_));
 sg13g2_o21ai_1 _4104_ (.B1(net49),
    .Y(_0438_),
    .A1(_0036_),
    .A2(net44));
 sg13g2_o21ai_1 _4105_ (.B1(_0438_),
    .Y(_0439_),
    .A1(net49),
    .A2(_0437_));
 sg13g2_nand2_1 _4106_ (.Y(_0440_),
    .A(_0439_),
    .B(net36));
 sg13g2_a21oi_1 _4107_ (.A1(net25),
    .A2(_1959_),
    .Y(_0441_),
    .B1(net36));
 sg13g2_o21ai_1 _4108_ (.B1(_0441_),
    .Y(_0442_),
    .A1(net44),
    .A2(net25));
 sg13g2_nand3_1 _4109_ (.B(net42),
    .C(_0442_),
    .A(_0440_),
    .Y(_0443_));
 sg13g2_a21oi_1 _4110_ (.A1(_1966_),
    .A2(net35),
    .Y(_0444_),
    .B1(net30));
 sg13g2_nand2_1 _4111_ (.Y(_0445_),
    .A(_0443_),
    .B(_0444_));
 sg13g2_a21o_1 _4112_ (.A2(_0445_),
    .A1(_0422_),
    .B1(_0245_),
    .X(_0446_));
 sg13g2_a21oi_1 _4113_ (.A1(_0419_),
    .A2(net23),
    .Y(_0447_),
    .B1(_0446_));
 sg13g2_nand3_1 _4114_ (.B(_0418_),
    .C(_0447_),
    .A(_0415_),
    .Y(_0448_));
 sg13g2_nand3_1 _4115_ (.B(_0237_),
    .C(net54),
    .A(_0419_),
    .Y(_0449_));
 sg13g2_a21oi_2 _4116_ (.B1(_0299_),
    .Y(_0450_),
    .A2(_0241_),
    .A1(_0408_));
 sg13g2_nand2_1 _4117_ (.Y(_0451_),
    .A(_0419_),
    .B(_0450_));
 sg13g2_nand3_1 _4118_ (.B(net31),
    .C(_0451_),
    .A(_0449_),
    .Y(_0452_));
 sg13g2_a21oi_2 _4119_ (.B1(_0452_),
    .Y(_0453_),
    .A2(net51),
    .A1(_0303_));
 sg13g2_nor2_2 _4120_ (.A(_0246_),
    .B(net22),
    .Y(_0454_));
 sg13g2_inv_2 _4121_ (.Y(_0455_),
    .A(_0454_));
 sg13g2_nand3_1 _4122_ (.B(_0453_),
    .C(_0455_),
    .A(_0448_),
    .Y(_0456_));
 sg13g2_nand2_1 _4123_ (.Y(_0457_),
    .A(_0309_),
    .B(_0246_));
 sg13g2_nand2_1 _4124_ (.Y(_0458_),
    .A(_0298_),
    .B(_0225_));
 sg13g2_nand2_1 _4125_ (.Y(_0459_),
    .A(_0458_),
    .B(_0300_));
 sg13g2_nand2_1 _4126_ (.Y(_0460_),
    .A(_0407_),
    .B(_0450_));
 sg13g2_o21ai_1 _4127_ (.B1(_0460_),
    .Y(_0461_),
    .A1(_0459_),
    .A2(_1889_));
 sg13g2_nor2_1 _4128_ (.A(_0457_),
    .B(_0461_),
    .Y(_0462_));
 sg13g2_nor2_2 _4129_ (.A(_0454_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_nand3_1 _4130_ (.B(_0456_),
    .C(_0463_),
    .A(_0413_),
    .Y(_0464_));
 sg13g2_nor3_1 _4131_ (.A(_0454_),
    .B(_0453_),
    .C(_0448_),
    .Y(_0465_));
 sg13g2_inv_4 _4132_ (.A(_0457_),
    .Y(_0466_));
 sg13g2_xnor2_1 _4133_ (.Y(_0467_),
    .A(_1953_),
    .B(_0396_));
 sg13g2_o21ai_1 _4134_ (.B1(_0155_),
    .Y(_0468_),
    .A1(net43),
    .A2(_0467_));
 sg13g2_xnor2_1 _4135_ (.Y(_0469_),
    .A(_1522_),
    .B(net38));
 sg13g2_inv_1 _4136_ (.Y(_0470_),
    .A(_0469_));
 sg13g2_a21oi_1 _4137_ (.A1(_0470_),
    .A2(net53),
    .Y(_0471_),
    .B1(net47));
 sg13g2_mux2_1 _4138_ (.A0(_0159_),
    .A1(_0384_),
    .S(net81),
    .X(_0472_));
 sg13g2_buf_1 _4139_ (.A(_0472_),
    .X(_0473_));
 sg13g2_nand3_1 _4140_ (.B(net50),
    .C(net48),
    .A(_0473_),
    .Y(_0474_));
 sg13g2_o21ai_1 _4141_ (.B1(_2013_),
    .Y(_0475_),
    .A1(_2026_),
    .A2(_2024_));
 sg13g2_xnor2_1 _4142_ (.Y(_0476_),
    .A(_2014_),
    .B(_0475_));
 sg13g2_xnor2_1 _4143_ (.Y(_0477_),
    .A(_0346_),
    .B(_1969_));
 sg13g2_xnor2_1 _4144_ (.Y(_0478_),
    .A(_0476_),
    .B(_0477_));
 sg13g2_a22oi_1 _4145_ (.Y(_0479_),
    .B1(net40),
    .B2(_0478_),
    .A2(_0474_),
    .A1(_0471_));
 sg13g2_nor2_1 _4146_ (.A(_0035_),
    .B(net50),
    .Y(_0480_));
 sg13g2_a21oi_1 _4147_ (.A1(_1982_),
    .A2(_0480_),
    .Y(_0481_),
    .B1(net45));
 sg13g2_dfrbp_1 _4148_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net86),
    .D(_0000_),
    .Q_N(_2113_),
    .Q(_0012_));
 sg13g2_dfrbp_1 _4149_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net87),
    .D(_0001_),
    .Q_N(_2114_),
    .Q(_0013_));
 sg13g2_dfrbp_1 _4150_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net88),
    .D(_0002_),
    .Q_N(_2112_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _4151_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net89),
    .D(_0057_),
    .Q_N(_2115_),
    .Q(_0016_));
 sg13g2_dfrbp_1 _4152_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net90),
    .D(_0003_),
    .Q_N(_2111_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _4153_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net91),
    .D(_0004_),
    .Q_N(_2110_),
    .Q(_0145_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _4148__86 (.L_HI(net86));
 sg13g2_buf_1 _4156_ (.A(net92),
    .X(uio_oe[0]));
 sg13g2_buf_1 _4157_ (.A(net93),
    .X(uio_oe[1]));
 sg13g2_buf_1 _4158_ (.A(net94),
    .X(uio_oe[2]));
 sg13g2_buf_1 _4159_ (.A(net95),
    .X(uio_oe[3]));
 sg13g2_buf_1 _4160_ (.A(net96),
    .X(uio_oe[4]));
 sg13g2_buf_1 _4161_ (.A(net97),
    .X(uio_oe[5]));
 sg13g2_buf_1 _4162_ (.A(net98),
    .X(uio_oe[6]));
 sg13g2_buf_1 _4163_ (.A(net99),
    .X(uio_oe[7]));
 sg13g2_buf_1 _4164_ (.A(hsync),
    .X(net12));
 sg13g2_buf_1 _4165_ (.A(\i_project.controller_0.vga_sync.o_vsync ),
    .X(net13));
 sg13g2_buf_1 _4166_ (.A(net84),
    .X(uio_out[6]));
 sg13g2_buf_1 _4167_ (.A(net85),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \counter[0]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net100),
    .D(_0058_),
    .Q_N(_0055_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 \counter[10]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net101),
    .D(_0059_),
    .Q_N(_2109_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 \counter[11]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net102),
    .D(_0060_),
    .Q_N(_2108_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 \counter[12]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net103),
    .D(_0061_),
    .Q_N(_2107_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 \counter[13]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net104),
    .D(_0062_),
    .Q_N(_2106_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 \counter[14]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net105),
    .D(_0063_),
    .Q_N(_2105_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 \counter[15]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net106),
    .D(_0064_),
    .Q_N(_2104_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 \counter[16]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net107),
    .D(_0065_),
    .Q_N(_2103_),
    .Q(\counter[16] ));
 sg13g2_dfrbp_1 \counter[17]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net108),
    .D(_0066_),
    .Q_N(_2102_),
    .Q(\counter[17] ));
 sg13g2_dfrbp_1 \counter[18]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net109),
    .D(_0067_),
    .Q_N(_2101_),
    .Q(\counter[18] ));
 sg13g2_dfrbp_1 \counter[19]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net110),
    .D(_0068_),
    .Q_N(_2100_),
    .Q(\counter[19] ));
 sg13g2_dfrbp_1 \counter[1]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net111),
    .D(_0069_),
    .Q_N(_2099_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 \counter[20]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net112),
    .D(_0070_),
    .Q_N(_2098_),
    .Q(\counter[20] ));
 sg13g2_dfrbp_1 \counter[21]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net113),
    .D(_0071_),
    .Q_N(_2097_),
    .Q(\counter[21] ));
 sg13g2_dfrbp_1 \counter[22]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net114),
    .D(_0072_),
    .Q_N(_2096_),
    .Q(\counter[22] ));
 sg13g2_dfrbp_1 \counter[23]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net115),
    .D(_0073_),
    .Q_N(_2095_),
    .Q(\counter[23] ));
 sg13g2_dfrbp_1 \counter[24]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net116),
    .D(_0074_),
    .Q_N(_2094_),
    .Q(\counter[24] ));
 sg13g2_dfrbp_1 \counter[25]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net117),
    .D(_0075_),
    .Q_N(_2093_),
    .Q(\counter[25] ));
 sg13g2_dfrbp_1 \counter[26]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net118),
    .D(_0076_),
    .Q_N(_2092_),
    .Q(\counter[26] ));
 sg13g2_dfrbp_1 \counter[27]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net119),
    .D(_0077_),
    .Q_N(_2091_),
    .Q(\counter[27] ));
 sg13g2_dfrbp_1 \counter[28]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net120),
    .D(_0078_),
    .Q_N(_2090_),
    .Q(\counter[28] ));
 sg13g2_dfrbp_1 \counter[29]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net121),
    .D(_0079_),
    .Q_N(_2089_),
    .Q(\counter[29] ));
 sg13g2_dfrbp_1 \counter[2]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net122),
    .D(_0080_),
    .Q_N(_2088_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 \counter[30]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net123),
    .D(_0081_),
    .Q_N(_2087_),
    .Q(\counter[30] ));
 sg13g2_dfrbp_1 \counter[31]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net124),
    .D(_0082_),
    .Q_N(_2086_),
    .Q(\counter[31] ));
 sg13g2_dfrbp_1 \counter[3]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net125),
    .D(_0083_),
    .Q_N(_2085_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 \counter[4]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net126),
    .D(_0084_),
    .Q_N(_2084_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 \counter[5]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net127),
    .D(_0085_),
    .Q_N(_2083_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 \counter[6]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net128),
    .D(_0086_),
    .Q_N(_2082_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 \counter[7]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(_0087_),
    .Q_N(_2081_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 \counter[8]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net130),
    .D(_0088_),
    .Q_N(_2080_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 \counter[9]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net131),
    .D(_0089_),
    .Q_N(_2116_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 \depth[0]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net132),
    .D(_0005_),
    .Q_N(_2117_),
    .Q(\depth[0] ));
 sg13g2_dfrbp_1 \depth[1]$_DFF_P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net133),
    .D(_0006_),
    .Q_N(_2118_),
    .Q(\depth[1] ));
 sg13g2_dfrbp_1 \depth[2]$_DFF_P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net134),
    .D(_0007_),
    .Q_N(_0044_),
    .Q(\depth[2] ));
 sg13g2_dfrbp_1 \dither_threshold[0]$_SDFFE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net135),
    .D(_0090_),
    .Q_N(_0029_),
    .Q(\dither_threshold[0] ));
 sg13g2_dfrbp_1 \dither_threshold[1]$_SDFFE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net136),
    .D(_0091_),
    .Q_N(_0018_),
    .Q(\dither_threshold[1] ));
 sg13g2_dfrbp_1 \dither_threshold[2]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net137),
    .D(_0092_),
    .Q_N(_0028_),
    .Q(\dither_threshold[2] ));
 sg13g2_dfrbp_1 \dither_threshold[3]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net138),
    .D(_0093_),
    .Q_N(_0033_),
    .Q(\dither_threshold[3] ));
 sg13g2_dfrbp_1 \dither_threshold[4]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net139),
    .D(_0094_),
    .Q_N(_0027_),
    .Q(\dither_threshold[4] ));
 sg13g2_dfrbp_1 \frame_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net140),
    .D(_0095_),
    .Q_N(_0054_),
    .Q(\frame_counter[0] ));
 sg13g2_dfrbp_1 \frame_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net141),
    .D(_0096_),
    .Q_N(_2079_),
    .Q(\frame_counter[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[2]$_DFFE_PN_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net142),
    .D(_0003_),
    .Q_N(_2078_),
    .Q(\i_project.controller_0.divider[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[3]$_DFFE_PN_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net143),
    .D(_0004_),
    .Q_N(_2077_),
    .Q(\i_project.controller_0.divider[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[4]$_DFFE_PN_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net144),
    .D(_0097_),
    .Q_N(_2076_),
    .Q(\i_project.controller_0.mode[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[5]$_DFFE_PN_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net145),
    .D(_0098_),
    .Q_N(_2075_),
    .Q(\i_project.controller_0.mode[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[6]$_DFFE_PN_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net146),
    .D(_0099_),
    .Q_N(_0025_),
    .Q(\i_project.controller_0.mode[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[7]$_DFFE_PN_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net147),
    .D(_0100_),
    .Q_N(_0022_),
    .Q(\i_project.controller_0.vga_sync.mode ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[0]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net148),
    .D(_0101_),
    .Q_N(_0056_),
    .Q(\i_project.controller_0.mode_ramp_base[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[10]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net149),
    .D(_0102_),
    .Q_N(_0037_),
    .Q(\i_project.controller_0.t[10] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[11]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net150),
    .D(_0103_),
    .Q_N(_2074_),
    .Q(\i_project.controller_0.t[11] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[1]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net151),
    .D(_0104_),
    .Q_N(_0021_),
    .Q(\i_project.controller_0.mode_ramp_base[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[2]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net152),
    .D(_0105_),
    .Q_N(_0020_),
    .Q(\i_project.controller_0.mode_ramp_base[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[3]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net153),
    .D(_0106_),
    .Q_N(_0019_),
    .Q(\i_project.controller_0.mode_ramp_base[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[4]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net154),
    .D(_0107_),
    .Q_N(_0043_),
    .Q(\i_project.controller_0.mode_ramp_base[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[5]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net155),
    .D(_0108_),
    .Q_N(_0042_),
    .Q(\i_project.controller_0.mode_ramp_base[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[6]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net156),
    .D(_0109_),
    .Q_N(_0041_),
    .Q(\i_project.controller_0.mode_ramp_base[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[7]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net157),
    .D(_0110_),
    .Q_N(_0040_),
    .Q(\i_project.controller_0.mode_ramp_base[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[8]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net158),
    .D(_0111_),
    .Q_N(_0039_),
    .Q(\i_project.controller_0.t[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[9]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net159),
    .D(_0112_),
    .Q_N(_0038_),
    .Q(\i_project.controller_0.t[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[0]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net160),
    .D(_0113_),
    .Q_N(_0053_),
    .Q(\i_project.controller_0.h[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[1]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net161),
    .D(_0114_),
    .Q_N(_0036_),
    .Q(\i_project.controller_0.h[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[2]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net162),
    .D(_0115_),
    .Q_N(_0035_),
    .Q(\i_project.controller_0.h[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[3]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net163),
    .D(_0116_),
    .Q_N(_0024_),
    .Q(\i_project.controller_0.h[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[4]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net164),
    .D(_0117_),
    .Q_N(_0046_),
    .Q(\i_project.controller_0.h[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[5]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net165),
    .D(_0118_),
    .Q_N(_0047_),
    .Q(\i_project.controller_0.h[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[6]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net166),
    .D(_0119_),
    .Q_N(_0048_),
    .Q(\i_project.controller_0.h[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[7]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net167),
    .D(_0120_),
    .Q_N(_0023_),
    .Q(\i_project.controller_0.h[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[8]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net168),
    .D(_0121_),
    .Q_N(_0026_),
    .Q(\i_project.controller_0.h[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[9]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net169),
    .D(_0122_),
    .Q_N(_0050_),
    .Q(\i_project.controller_0.h[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hsync$_DFFE_PP_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net170),
    .D(_0123_),
    .Q_N(hsync),
    .Q(\i_project.controller_0.vga_sync.hsync ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[0]$_SDFFE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net171),
    .D(_0124_),
    .Q_N(_2073_),
    .Q(\i_project.controller_0.v[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[1]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net172),
    .D(_0125_),
    .Q_N(_2072_),
    .Q(\i_project.controller_0.v[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[2]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net173),
    .D(_0126_),
    .Q_N(_2071_),
    .Q(\i_project.controller_0.v[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[3]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net174),
    .D(_0127_),
    .Q_N(_2070_),
    .Q(\i_project.controller_0.v[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[4]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net175),
    .D(_0128_),
    .Q_N(_2069_),
    .Q(\i_project.controller_0.v[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[5]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net176),
    .D(_0129_),
    .Q_N(_0031_),
    .Q(\i_project.controller_0.v[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[6]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net177),
    .D(_0130_),
    .Q_N(_2068_),
    .Q(\i_project.controller_0.v[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[7]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net178),
    .D(_0131_),
    .Q_N(_2067_),
    .Q(\i_project.controller_0.v[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[8]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net179),
    .D(_0132_),
    .Q_N(_0032_),
    .Q(\i_project.controller_0.v[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[9]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net180),
    .D(_0133_),
    .Q_N(_0030_),
    .Q(\i_project.controller_0.v[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vsync$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net181),
    .D(_0134_),
    .Q_N(_2066_),
    .Q(\i_project.controller_0.vga_sync.vsync ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[0]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net182),
    .D(_0135_),
    .Q_N(_2065_),
    .Q(\i_project.controller_0.voffset[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[1]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net183),
    .D(_0136_),
    .Q_N(_2064_),
    .Q(\i_project.controller_0.voffset[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[2]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net184),
    .D(_0137_),
    .Q_N(_2063_),
    .Q(\i_project.controller_0.voffset[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[3]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net185),
    .D(_0138_),
    .Q_N(_2062_),
    .Q(\i_project.controller_0.voffset[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[4]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net186),
    .D(_0139_),
    .Q_N(_2061_),
    .Q(\i_project.controller_0.voffset[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[5]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net187),
    .D(_0140_),
    .Q_N(_2060_),
    .Q(\i_project.controller_0.voffset[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[6]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net188),
    .D(_0141_),
    .Q_N(_2059_),
    .Q(\i_project.controller_0.voffset[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[7]$_SDFFCE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net189),
    .D(_0142_),
    .Q_N(_2058_),
    .Q(\i_project.controller_0.voffset[7] ));
 sg13g2_dfrbp_1 \prev_vsync$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net190),
    .D(_0143_),
    .Q_N(_2119_),
    .Q(prev_vsync));
 sg13g2_dfrbp_1 \project_rst_n$_DFF_P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net191),
    .D(_0008_),
    .Q_N(_2120_),
    .Q(\i_project.controller_0.rst_n ));
 sg13g2_dfrbp_1 \project_ui_in[2]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net192),
    .D(\counter[30] ),
    .Q_N(_0052_),
    .Q(\i_project.controller_0.grey_pass[10] ));
 sg13g2_dfrbp_1 \project_ui_in[3]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net193),
    .D(\counter[31] ),
    .Q_N(_0051_),
    .Q(\i_project.controller_0.grey_pass[11] ));
 sg13g2_dfrbp_1 \project_ui_in[4]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net194),
    .D(_0009_),
    .Q_N(_0045_),
    .Q(\i_project.controller_0.grey_pass[12] ));
 sg13g2_dfrbp_1 \project_ui_in[5]$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net195),
    .D(_0010_),
    .Q_N(_0017_),
    .Q(\i_project.controller_0.grey_pass[13] ));
 sg13g2_dfrbp_1 \project_ui_in[6]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net196),
    .D(_0011_),
    .Q_N(_0049_),
    .Q(\i_project.controller_0.grey_pass[14] ));
 sg13g2_dfrbp_1 \project_ui_in[7]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net197),
    .D(_0144_),
    .Q_N(_0034_),
    .Q(\i_project.controller_0.grey_pass[15] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[3]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[4]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[2]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[3]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[4]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[5]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[6]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout22 (.A(_0303_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0410_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0414_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0397_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0214_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0169_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1721_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0396_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0402_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0247_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_2007_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1978_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1942_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0335_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0327_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0176_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1953_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0399_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0388_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0334_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0329_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0326_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1959_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0367_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0333_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0315_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2044_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0323_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0310_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0308_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0150_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2043_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1888_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1838_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1624_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2041_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1644_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_2046_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1857_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1853_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1795_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1783_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1549_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1540_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1533_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1525_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1521_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1499_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1859_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1849_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_1843_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1841_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1685_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1584_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1583_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1578_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1534_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1515_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1514_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1503_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1478_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1506_),
    .X(net83));
 sg13g2_tielo _4166__84 (.L_LO(net84));
 sg13g2_tielo _4167__85 (.L_LO(net85));
 sg13g2_tiehi _4149__87 (.L_HI(net87));
 sg13g2_tiehi _4150__88 (.L_HI(net88));
 sg13g2_tiehi _4151__89 (.L_HI(net89));
 sg13g2_tiehi _4152__90 (.L_HI(net90));
 sg13g2_tiehi _4153__91 (.L_HI(net91));
 sg13g2_tiehi _4156__92 (.L_HI(net92));
 sg13g2_tiehi _4157__93 (.L_HI(net93));
 sg13g2_tiehi _4158__94 (.L_HI(net94));
 sg13g2_tiehi _4159__95 (.L_HI(net95));
 sg13g2_tiehi _4160__96 (.L_HI(net96));
 sg13g2_tiehi _4161__97 (.L_HI(net97));
 sg13g2_tiehi _4162__98 (.L_HI(net98));
 sg13g2_tiehi _4163__99 (.L_HI(net99));
 sg13g2_tiehi \counter[0]$_SDFF_PN0__100  (.L_HI(net100));
 sg13g2_tiehi \counter[10]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_tiehi \counter[11]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \counter[12]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_tiehi \counter[13]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_tiehi \counter[14]$_SDFF_PN0__105  (.L_HI(net105));
 sg13g2_tiehi \counter[15]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_tiehi \counter[16]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_tiehi \counter[17]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \counter[18]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_tiehi \counter[19]$_SDFF_PN0__110  (.L_HI(net110));
 sg13g2_tiehi \counter[1]$_SDFF_PN0__111  (.L_HI(net111));
 sg13g2_tiehi \counter[20]$_SDFF_PN0__112  (.L_HI(net112));
 sg13g2_tiehi \counter[21]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_tiehi \counter[22]$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_tiehi \counter[23]$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \counter[24]$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \counter[25]$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_tiehi \counter[26]$_SDFF_PN0__118  (.L_HI(net118));
 sg13g2_tiehi \counter[27]$_SDFF_PN0__119  (.L_HI(net119));
 sg13g2_tiehi \counter[28]$_SDFF_PN0__120  (.L_HI(net120));
 sg13g2_tiehi \counter[29]$_SDFF_PN0__121  (.L_HI(net121));
 sg13g2_tiehi \counter[2]$_SDFF_PN0__122  (.L_HI(net122));
 sg13g2_tiehi \counter[30]$_SDFF_PN0__123  (.L_HI(net123));
 sg13g2_tiehi \counter[31]$_SDFF_PN0__124  (.L_HI(net124));
 sg13g2_tiehi \counter[3]$_SDFF_PN0__125  (.L_HI(net125));
 sg13g2_tiehi \counter[4]$_SDFF_PN0__126  (.L_HI(net126));
 sg13g2_tiehi \counter[5]$_SDFF_PN0__127  (.L_HI(net127));
 sg13g2_tiehi \counter[6]$_SDFF_PN0__128  (.L_HI(net128));
 sg13g2_tiehi \counter[7]$_SDFF_PN0__129  (.L_HI(net129));
 sg13g2_tiehi \counter[8]$_SDFF_PN0__130  (.L_HI(net130));
 sg13g2_tiehi \counter[9]$_SDFF_PN0__131  (.L_HI(net131));
 sg13g2_tiehi \depth[0]$_DFF_P__132  (.L_HI(net132));
 sg13g2_tiehi \depth[1]$_DFF_P__133  (.L_HI(net133));
 sg13g2_tiehi \depth[2]$_DFF_P__134  (.L_HI(net134));
 sg13g2_tiehi \dither_threshold[0]$_SDFFE_PP0P__135  (.L_HI(net135));
 sg13g2_tiehi \dither_threshold[1]$_SDFFE_PP0P__136  (.L_HI(net136));
 sg13g2_tiehi \dither_threshold[2]$_SDFF_PP0__137  (.L_HI(net137));
 sg13g2_tiehi \dither_threshold[3]$_SDFF_PP0__138  (.L_HI(net138));
 sg13g2_tiehi \dither_threshold[4]$_SDFF_PP0__139  (.L_HI(net139));
 sg13g2_tiehi \frame_counter[0]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \frame_counter[1]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \i_project.controller_0.mode_params[2]$_DFFE_PN__142  (.L_HI(net142));
 sg13g2_tiehi \i_project.controller_0.mode_params[3]$_DFFE_PN__143  (.L_HI(net143));
 sg13g2_tiehi \i_project.controller_0.mode_params[4]$_DFFE_PN__144  (.L_HI(net144));
 sg13g2_tiehi \i_project.controller_0.mode_params[5]$_DFFE_PN__145  (.L_HI(net145));
 sg13g2_tiehi \i_project.controller_0.mode_params[6]$_DFFE_PN__146  (.L_HI(net146));
 sg13g2_tiehi \i_project.controller_0.mode_params[7]$_DFFE_PN__147  (.L_HI(net147));
 sg13g2_tiehi \i_project.controller_0.t[0]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \i_project.controller_0.t[10]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \i_project.controller_0.t[11]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \i_project.controller_0.t[1]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \i_project.controller_0.t[2]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \i_project.controller_0.t[3]$_SDFFE_PN0P__153  (.L_HI(net153));
 sg13g2_tiehi \i_project.controller_0.t[4]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \i_project.controller_0.t[5]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \i_project.controller_0.t[6]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \i_project.controller_0.t[7]$_SDFFE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \i_project.controller_0.t[8]$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \i_project.controller_0.t[9]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[0]$_SDFF_PP0__160  (.L_HI(net160));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[1]$_SDFF_PP0__161  (.L_HI(net161));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[2]$_SDFF_PP0__162  (.L_HI(net162));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[3]$_SDFF_PP0__163  (.L_HI(net163));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[4]$_SDFF_PP0__164  (.L_HI(net164));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[5]$_SDFF_PP0__165  (.L_HI(net165));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[6]$_SDFF_PP0__166  (.L_HI(net166));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[7]$_SDFF_PP0__167  (.L_HI(net167));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[8]$_SDFF_PP0__168  (.L_HI(net168));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[9]$_SDFF_PP0__169  (.L_HI(net169));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hsync$_DFFE_PP__170  (.L_HI(net170));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[0]$_SDFFE_PP0P__171  (.L_HI(net171));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[1]$_SDFFE_PP0P__172  (.L_HI(net172));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[2]$_SDFFE_PP0P__173  (.L_HI(net173));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[3]$_SDFFE_PP0P__174  (.L_HI(net174));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[4]$_SDFFE_PP0P__175  (.L_HI(net175));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[5]$_SDFFE_PP0P__176  (.L_HI(net176));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[6]$_SDFFE_PP0P__177  (.L_HI(net177));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[7]$_SDFFE_PP0P__178  (.L_HI(net178));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[8]$_SDFFE_PP0P__179  (.L_HI(net179));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[9]$_SDFFE_PP0P__180  (.L_HI(net180));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vsync$_DFFE_PP__181  (.L_HI(net181));
 sg13g2_tiehi \i_project.controller_0.voffset[0]$_DFFE_PP__182  (.L_HI(net182));
 sg13g2_tiehi \i_project.controller_0.voffset[1]$_DFFE_PP__183  (.L_HI(net183));
 sg13g2_tiehi \i_project.controller_0.voffset[2]$_DFFE_PP__184  (.L_HI(net184));
 sg13g2_tiehi \i_project.controller_0.voffset[3]$_SDFFCE_PP0P__185  (.L_HI(net185));
 sg13g2_tiehi \i_project.controller_0.voffset[4]$_SDFFCE_PP0P__186  (.L_HI(net186));
 sg13g2_tiehi \i_project.controller_0.voffset[5]$_DFFE_PP__187  (.L_HI(net187));
 sg13g2_tiehi \i_project.controller_0.voffset[6]$_DFFE_PP__188  (.L_HI(net188));
 sg13g2_tiehi \i_project.controller_0.voffset[7]$_SDFFCE_PN0P__189  (.L_HI(net189));
 sg13g2_tiehi \prev_vsync$_SDFF_PN0__190  (.L_HI(net190));
 sg13g2_tiehi \project_rst_n$_DFF_P__191  (.L_HI(net191));
 sg13g2_tiehi \project_ui_in[2]$_DFF_P__192  (.L_HI(net192));
 sg13g2_tiehi \project_ui_in[3]$_DFF_P__193  (.L_HI(net193));
 sg13g2_tiehi \project_ui_in[4]$_DFF_P__194  (.L_HI(net194));
 sg13g2_tiehi \project_ui_in[5]$_DFF_P__195  (.L_HI(net195));
 sg13g2_tiehi \project_ui_in[6]$_DFF_P__196  (.L_HI(net196));
 sg13g2_tiehi \project_ui_in[7]$_SDFF_PN0__197  (.L_HI(net197));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_fill_2 FILLER_0_67 ();
 sg13g2_fill_1 FILLER_0_74 ();
 sg13g2_decap_4 FILLER_0_101 ();
 sg13g2_fill_1 FILLER_0_110 ();
 sg13g2_fill_1 FILLER_0_119 ();
 sg13g2_decap_4 FILLER_0_133 ();
 sg13g2_decap_4 FILLER_0_145 ();
 sg13g2_fill_1 FILLER_0_149 ();
 sg13g2_fill_2 FILLER_0_190 ();
 sg13g2_fill_1 FILLER_0_192 ();
 sg13g2_decap_4 FILLER_0_240 ();
 sg13g2_fill_2 FILLER_0_244 ();
 sg13g2_fill_1 FILLER_0_251 ();
 sg13g2_fill_1 FILLER_0_260 ();
 sg13g2_decap_4 FILLER_0_278 ();
 sg13g2_decap_4 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_4 FILLER_0_425 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_4 FILLER_1_49 ();
 sg13g2_fill_1 FILLER_1_110 ();
 sg13g2_fill_1 FILLER_1_114 ();
 sg13g2_fill_1 FILLER_1_119 ();
 sg13g2_fill_2 FILLER_1_128 ();
 sg13g2_fill_2 FILLER_1_138 ();
 sg13g2_fill_2 FILLER_1_148 ();
 sg13g2_fill_1 FILLER_1_150 ();
 sg13g2_decap_4 FILLER_1_159 ();
 sg13g2_fill_2 FILLER_1_167 ();
 sg13g2_fill_1 FILLER_1_169 ();
 sg13g2_fill_1 FILLER_1_174 ();
 sg13g2_fill_1 FILLER_1_186 ();
 sg13g2_fill_1 FILLER_1_194 ();
 sg13g2_fill_1 FILLER_1_200 ();
 sg13g2_fill_2 FILLER_1_220 ();
 sg13g2_fill_2 FILLER_1_233 ();
 sg13g2_fill_1 FILLER_1_253 ();
 sg13g2_fill_2 FILLER_1_264 ();
 sg13g2_fill_1 FILLER_1_287 ();
 sg13g2_fill_1 FILLER_1_292 ();
 sg13g2_fill_1 FILLER_1_296 ();
 sg13g2_fill_1 FILLER_1_302 ();
 sg13g2_fill_1 FILLER_1_308 ();
 sg13g2_fill_2 FILLER_1_313 ();
 sg13g2_fill_1 FILLER_1_320 ();
 sg13g2_fill_2 FILLER_1_325 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_fill_2 FILLER_1_350 ();
 sg13g2_fill_1 FILLER_1_352 ();
 sg13g2_fill_2 FILLER_1_384 ();
 sg13g2_fill_1 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_8 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_1_412 ();
 sg13g2_decap_8 FILLER_1_419 ();
 sg13g2_decap_4 FILLER_1_426 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_75 ();
 sg13g2_fill_2 FILLER_2_90 ();
 sg13g2_fill_1 FILLER_2_92 ();
 sg13g2_fill_1 FILLER_2_118 ();
 sg13g2_fill_1 FILLER_2_123 ();
 sg13g2_fill_1 FILLER_2_132 ();
 sg13g2_fill_2 FILLER_2_137 ();
 sg13g2_fill_1 FILLER_2_147 ();
 sg13g2_fill_1 FILLER_2_152 ();
 sg13g2_fill_2 FILLER_2_161 ();
 sg13g2_fill_2 FILLER_2_168 ();
 sg13g2_fill_2 FILLER_2_175 ();
 sg13g2_fill_1 FILLER_2_208 ();
 sg13g2_fill_1 FILLER_2_247 ();
 sg13g2_decap_4 FILLER_2_270 ();
 sg13g2_fill_1 FILLER_2_274 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_fill_1 FILLER_2_329 ();
 sg13g2_fill_1 FILLER_2_334 ();
 sg13g2_fill_2 FILLER_2_345 ();
 sg13g2_fill_1 FILLER_2_347 ();
 sg13g2_decap_4 FILLER_2_351 ();
 sg13g2_fill_2 FILLER_2_355 ();
 sg13g2_fill_2 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_4 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_38 ();
 sg13g2_fill_2 FILLER_3_45 ();
 sg13g2_decap_4 FILLER_3_69 ();
 sg13g2_fill_1 FILLER_3_73 ();
 sg13g2_decap_4 FILLER_3_79 ();
 sg13g2_fill_1 FILLER_3_100 ();
 sg13g2_fill_2 FILLER_3_114 ();
 sg13g2_fill_2 FILLER_3_124 ();
 sg13g2_fill_2 FILLER_3_134 ();
 sg13g2_fill_1 FILLER_3_136 ();
 sg13g2_fill_1 FILLER_3_149 ();
 sg13g2_decap_4 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_174 ();
 sg13g2_fill_1 FILLER_3_185 ();
 sg13g2_fill_1 FILLER_3_189 ();
 sg13g2_fill_2 FILLER_3_195 ();
 sg13g2_decap_8 FILLER_3_205 ();
 sg13g2_fill_1 FILLER_3_217 ();
 sg13g2_decap_4 FILLER_3_222 ();
 sg13g2_fill_2 FILLER_3_249 ();
 sg13g2_decap_4 FILLER_3_255 ();
 sg13g2_fill_2 FILLER_3_271 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_fill_1 FILLER_3_288 ();
 sg13g2_decap_4 FILLER_3_297 ();
 sg13g2_fill_2 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_311 ();
 sg13g2_decap_4 FILLER_3_318 ();
 sg13g2_fill_1 FILLER_3_352 ();
 sg13g2_fill_2 FILLER_3_388 ();
 sg13g2_fill_1 FILLER_3_390 ();
 sg13g2_decap_4 FILLER_3_395 ();
 sg13g2_fill_1 FILLER_3_403 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_13 ();
 sg13g2_fill_1 FILLER_4_20 ();
 sg13g2_fill_2 FILLER_4_33 ();
 sg13g2_fill_1 FILLER_4_35 ();
 sg13g2_fill_2 FILLER_4_70 ();
 sg13g2_fill_1 FILLER_4_83 ();
 sg13g2_fill_1 FILLER_4_92 ();
 sg13g2_fill_1 FILLER_4_101 ();
 sg13g2_decap_8 FILLER_4_115 ();
 sg13g2_fill_2 FILLER_4_137 ();
 sg13g2_fill_1 FILLER_4_149 ();
 sg13g2_fill_1 FILLER_4_162 ();
 sg13g2_fill_2 FILLER_4_167 ();
 sg13g2_fill_1 FILLER_4_177 ();
 sg13g2_fill_1 FILLER_4_186 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_fill_2 FILLER_4_205 ();
 sg13g2_decap_8 FILLER_4_215 ();
 sg13g2_decap_4 FILLER_4_222 ();
 sg13g2_fill_1 FILLER_4_226 ();
 sg13g2_decap_4 FILLER_4_240 ();
 sg13g2_decap_8 FILLER_4_249 ();
 sg13g2_decap_4 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_fill_1 FILLER_4_289 ();
 sg13g2_fill_2 FILLER_4_295 ();
 sg13g2_fill_1 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_320 ();
 sg13g2_fill_1 FILLER_4_327 ();
 sg13g2_decap_4 FILLER_4_335 ();
 sg13g2_fill_1 FILLER_4_339 ();
 sg13g2_fill_2 FILLER_4_344 ();
 sg13g2_fill_2 FILLER_4_358 ();
 sg13g2_fill_1 FILLER_4_360 ();
 sg13g2_fill_1 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_27 ();
 sg13g2_fill_1 FILLER_5_48 ();
 sg13g2_fill_2 FILLER_5_72 ();
 sg13g2_fill_2 FILLER_5_82 ();
 sg13g2_fill_1 FILLER_5_84 ();
 sg13g2_fill_2 FILLER_5_89 ();
 sg13g2_fill_1 FILLER_5_91 ();
 sg13g2_fill_2 FILLER_5_100 ();
 sg13g2_fill_1 FILLER_5_102 ();
 sg13g2_fill_2 FILLER_5_108 ();
 sg13g2_fill_2 FILLER_5_123 ();
 sg13g2_fill_1 FILLER_5_134 ();
 sg13g2_fill_1 FILLER_5_140 ();
 sg13g2_fill_1 FILLER_5_146 ();
 sg13g2_fill_1 FILLER_5_155 ();
 sg13g2_decap_4 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_fill_2 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_fill_2 FILLER_5_193 ();
 sg13g2_fill_1 FILLER_5_195 ();
 sg13g2_fill_2 FILLER_5_212 ();
 sg13g2_fill_2 FILLER_5_218 ();
 sg13g2_fill_1 FILLER_5_220 ();
 sg13g2_fill_2 FILLER_5_229 ();
 sg13g2_fill_1 FILLER_5_231 ();
 sg13g2_fill_1 FILLER_5_235 ();
 sg13g2_fill_2 FILLER_5_245 ();
 sg13g2_fill_1 FILLER_5_251 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_4 FILLER_5_293 ();
 sg13g2_fill_1 FILLER_5_297 ();
 sg13g2_fill_1 FILLER_5_301 ();
 sg13g2_fill_2 FILLER_5_307 ();
 sg13g2_fill_1 FILLER_5_309 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_fill_1 FILLER_5_316 ();
 sg13g2_fill_1 FILLER_5_320 ();
 sg13g2_decap_4 FILLER_5_337 ();
 sg13g2_fill_1 FILLER_5_341 ();
 sg13g2_fill_2 FILLER_5_355 ();
 sg13g2_fill_1 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_fill_1 FILLER_5_368 ();
 sg13g2_fill_1 FILLER_5_413 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_fill_1 FILLER_6_20 ();
 sg13g2_fill_2 FILLER_6_25 ();
 sg13g2_fill_2 FILLER_6_67 ();
 sg13g2_fill_1 FILLER_6_77 ();
 sg13g2_fill_1 FILLER_6_86 ();
 sg13g2_fill_1 FILLER_6_91 ();
 sg13g2_fill_2 FILLER_6_125 ();
 sg13g2_fill_1 FILLER_6_140 ();
 sg13g2_fill_2 FILLER_6_146 ();
 sg13g2_decap_4 FILLER_6_152 ();
 sg13g2_fill_2 FILLER_6_173 ();
 sg13g2_fill_1 FILLER_6_186 ();
 sg13g2_fill_2 FILLER_6_195 ();
 sg13g2_fill_1 FILLER_6_205 ();
 sg13g2_fill_2 FILLER_6_209 ();
 sg13g2_fill_2 FILLER_6_215 ();
 sg13g2_decap_8 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_281 ();
 sg13g2_fill_2 FILLER_6_295 ();
 sg13g2_fill_1 FILLER_6_302 ();
 sg13g2_fill_2 FILLER_6_308 ();
 sg13g2_fill_2 FILLER_6_341 ();
 sg13g2_decap_4 FILLER_6_360 ();
 sg13g2_fill_2 FILLER_6_364 ();
 sg13g2_decap_4 FILLER_6_373 ();
 sg13g2_fill_2 FILLER_6_412 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_27 ();
 sg13g2_decap_4 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_43 ();
 sg13g2_fill_1 FILLER_7_56 ();
 sg13g2_fill_2 FILLER_7_65 ();
 sg13g2_fill_2 FILLER_7_80 ();
 sg13g2_fill_1 FILLER_7_82 ();
 sg13g2_fill_1 FILLER_7_88 ();
 sg13g2_fill_1 FILLER_7_94 ();
 sg13g2_fill_2 FILLER_7_104 ();
 sg13g2_fill_1 FILLER_7_122 ();
 sg13g2_fill_1 FILLER_7_130 ();
 sg13g2_fill_1 FILLER_7_135 ();
 sg13g2_fill_2 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_151 ();
 sg13g2_decap_4 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_fill_1 FILLER_7_191 ();
 sg13g2_decap_8 FILLER_7_198 ();
 sg13g2_decap_4 FILLER_7_205 ();
 sg13g2_fill_1 FILLER_7_209 ();
 sg13g2_decap_4 FILLER_7_238 ();
 sg13g2_fill_2 FILLER_7_242 ();
 sg13g2_fill_2 FILLER_7_260 ();
 sg13g2_decap_4 FILLER_7_276 ();
 sg13g2_fill_2 FILLER_7_283 ();
 sg13g2_fill_2 FILLER_7_289 ();
 sg13g2_fill_2 FILLER_7_297 ();
 sg13g2_fill_1 FILLER_7_299 ();
 sg13g2_fill_2 FILLER_7_317 ();
 sg13g2_fill_2 FILLER_7_336 ();
 sg13g2_fill_1 FILLER_7_350 ();
 sg13g2_fill_1 FILLER_7_356 ();
 sg13g2_fill_1 FILLER_7_361 ();
 sg13g2_fill_1 FILLER_7_366 ();
 sg13g2_fill_1 FILLER_7_373 ();
 sg13g2_fill_1 FILLER_7_381 ();
 sg13g2_fill_1 FILLER_7_403 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_12 ();
 sg13g2_fill_1 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_27 ();
 sg13g2_fill_1 FILLER_8_29 ();
 sg13g2_fill_1 FILLER_8_39 ();
 sg13g2_fill_2 FILLER_8_68 ();
 sg13g2_fill_1 FILLER_8_70 ();
 sg13g2_fill_2 FILLER_8_75 ();
 sg13g2_decap_4 FILLER_8_85 ();
 sg13g2_fill_1 FILLER_8_89 ();
 sg13g2_fill_1 FILLER_8_94 ();
 sg13g2_fill_1 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_137 ();
 sg13g2_fill_2 FILLER_8_143 ();
 sg13g2_fill_1 FILLER_8_145 ();
 sg13g2_fill_1 FILLER_8_150 ();
 sg13g2_decap_4 FILLER_8_163 ();
 sg13g2_fill_1 FILLER_8_180 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_210 ();
 sg13g2_fill_2 FILLER_8_247 ();
 sg13g2_fill_1 FILLER_8_256 ();
 sg13g2_fill_1 FILLER_8_262 ();
 sg13g2_fill_1 FILLER_8_267 ();
 sg13g2_fill_1 FILLER_8_272 ();
 sg13g2_fill_1 FILLER_8_278 ();
 sg13g2_fill_1 FILLER_8_283 ();
 sg13g2_decap_4 FILLER_8_306 ();
 sg13g2_fill_1 FILLER_8_310 ();
 sg13g2_fill_1 FILLER_8_322 ();
 sg13g2_fill_1 FILLER_8_336 ();
 sg13g2_fill_2 FILLER_8_341 ();
 sg13g2_fill_1 FILLER_8_343 ();
 sg13g2_fill_1 FILLER_8_357 ();
 sg13g2_fill_1 FILLER_8_367 ();
 sg13g2_fill_1 FILLER_8_376 ();
 sg13g2_fill_2 FILLER_8_385 ();
 sg13g2_fill_1 FILLER_8_414 ();
 sg13g2_decap_8 FILLER_8_419 ();
 sg13g2_decap_4 FILLER_8_426 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_14 ();
 sg13g2_fill_1 FILLER_9_18 ();
 sg13g2_fill_1 FILLER_9_40 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_fill_2 FILLER_9_57 ();
 sg13g2_fill_1 FILLER_9_59 ();
 sg13g2_fill_2 FILLER_9_68 ();
 sg13g2_fill_2 FILLER_9_86 ();
 sg13g2_fill_1 FILLER_9_102 ();
 sg13g2_decap_4 FILLER_9_111 ();
 sg13g2_fill_2 FILLER_9_115 ();
 sg13g2_decap_4 FILLER_9_145 ();
 sg13g2_fill_1 FILLER_9_158 ();
 sg13g2_fill_1 FILLER_9_163 ();
 sg13g2_fill_1 FILLER_9_168 ();
 sg13g2_fill_2 FILLER_9_173 ();
 sg13g2_decap_4 FILLER_9_184 ();
 sg13g2_fill_1 FILLER_9_188 ();
 sg13g2_fill_2 FILLER_9_213 ();
 sg13g2_fill_2 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_220 ();
 sg13g2_decap_4 FILLER_9_225 ();
 sg13g2_decap_4 FILLER_9_233 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_fill_1 FILLER_9_244 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_4 FILLER_9_315 ();
 sg13g2_fill_2 FILLER_9_319 ();
 sg13g2_fill_2 FILLER_9_326 ();
 sg13g2_fill_2 FILLER_9_332 ();
 sg13g2_fill_1 FILLER_9_334 ();
 sg13g2_fill_2 FILLER_9_338 ();
 sg13g2_fill_1 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_4 FILLER_9_365 ();
 sg13g2_fill_2 FILLER_9_369 ();
 sg13g2_fill_1 FILLER_9_375 ();
 sg13g2_fill_2 FILLER_9_414 ();
 sg13g2_fill_1 FILLER_9_416 ();
 sg13g2_decap_8 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_9 ();
 sg13g2_fill_1 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_52 ();
 sg13g2_decap_4 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_65 ();
 sg13g2_decap_4 FILLER_10_72 ();
 sg13g2_fill_1 FILLER_10_76 ();
 sg13g2_fill_2 FILLER_10_108 ();
 sg13g2_fill_2 FILLER_10_119 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_fill_2 FILLER_10_146 ();
 sg13g2_fill_1 FILLER_10_152 ();
 sg13g2_fill_1 FILLER_10_158 ();
 sg13g2_fill_2 FILLER_10_168 ();
 sg13g2_fill_2 FILLER_10_175 ();
 sg13g2_fill_2 FILLER_10_186 ();
 sg13g2_fill_1 FILLER_10_188 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_259 ();
 sg13g2_fill_2 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_272 ();
 sg13g2_fill_2 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_10_299 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_fill_2 FILLER_10_313 ();
 sg13g2_fill_1 FILLER_10_315 ();
 sg13g2_fill_1 FILLER_10_324 ();
 sg13g2_fill_1 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_fill_2 FILLER_10_364 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_32 ();
 sg13g2_fill_2 FILLER_11_53 ();
 sg13g2_fill_1 FILLER_11_71 ();
 sg13g2_decap_8 FILLER_11_85 ();
 sg13g2_fill_2 FILLER_11_97 ();
 sg13g2_decap_4 FILLER_11_106 ();
 sg13g2_decap_4 FILLER_11_121 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_139 ();
 sg13g2_fill_2 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_fill_2 FILLER_11_243 ();
 sg13g2_fill_1 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_277 ();
 sg13g2_fill_1 FILLER_11_283 ();
 sg13g2_decap_8 FILLER_11_356 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_11 ();
 sg13g2_fill_1 FILLER_12_20 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_fill_2 FILLER_12_82 ();
 sg13g2_fill_1 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_fill_1 FILLER_12_122 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_fill_1 FILLER_12_129 ();
 sg13g2_fill_2 FILLER_12_156 ();
 sg13g2_fill_2 FILLER_12_162 ();
 sg13g2_decap_8 FILLER_12_177 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_196 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_fill_1 FILLER_12_217 ();
 sg13g2_fill_1 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_235 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_269 ();
 sg13g2_fill_2 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_290 ();
 sg13g2_fill_2 FILLER_12_312 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_fill_2 FILLER_12_335 ();
 sg13g2_fill_1 FILLER_12_337 ();
 sg13g2_decap_4 FILLER_12_342 ();
 sg13g2_fill_1 FILLER_12_346 ();
 sg13g2_decap_4 FILLER_12_392 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_36 ();
 sg13g2_fill_1 FILLER_13_53 ();
 sg13g2_fill_1 FILLER_13_62 ();
 sg13g2_fill_2 FILLER_13_66 ();
 sg13g2_fill_1 FILLER_13_73 ();
 sg13g2_fill_2 FILLER_13_82 ();
 sg13g2_fill_1 FILLER_13_109 ();
 sg13g2_fill_1 FILLER_13_114 ();
 sg13g2_fill_2 FILLER_13_120 ();
 sg13g2_decap_4 FILLER_13_130 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_fill_2 FILLER_13_148 ();
 sg13g2_fill_1 FILLER_13_150 ();
 sg13g2_fill_1 FILLER_13_169 ();
 sg13g2_decap_4 FILLER_13_195 ();
 sg13g2_fill_1 FILLER_13_233 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_258 ();
 sg13g2_fill_2 FILLER_13_314 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_1 FILLER_13_358 ();
 sg13g2_fill_2 FILLER_13_368 ();
 sg13g2_fill_1 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_8 FILLER_13_419 ();
 sg13g2_decap_4 FILLER_13_426 ();
 sg13g2_fill_2 FILLER_14_30 ();
 sg13g2_fill_1 FILLER_14_32 ();
 sg13g2_fill_2 FILLER_14_41 ();
 sg13g2_fill_1 FILLER_14_60 ();
 sg13g2_decap_4 FILLER_14_66 ();
 sg13g2_fill_1 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_117 ();
 sg13g2_fill_1 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_128 ();
 sg13g2_fill_2 FILLER_14_144 ();
 sg13g2_fill_1 FILLER_14_146 ();
 sg13g2_fill_1 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_181 ();
 sg13g2_fill_2 FILLER_14_222 ();
 sg13g2_decap_4 FILLER_14_231 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_278 ();
 sg13g2_fill_2 FILLER_14_285 ();
 sg13g2_fill_2 FILLER_14_313 ();
 sg13g2_fill_1 FILLER_14_320 ();
 sg13g2_fill_1 FILLER_14_329 ();
 sg13g2_fill_2 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_fill_2 FILLER_14_354 ();
 sg13g2_fill_2 FILLER_14_377 ();
 sg13g2_fill_1 FILLER_14_379 ();
 sg13g2_fill_1 FILLER_14_390 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_fill_2 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_16 ();
 sg13g2_fill_2 FILLER_15_55 ();
 sg13g2_decap_4 FILLER_15_64 ();
 sg13g2_fill_1 FILLER_15_68 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_fill_2 FILLER_15_97 ();
 sg13g2_decap_4 FILLER_15_104 ();
 sg13g2_fill_1 FILLER_15_118 ();
 sg13g2_fill_1 FILLER_15_122 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_4 FILLER_15_151 ();
 sg13g2_fill_2 FILLER_15_160 ();
 sg13g2_fill_2 FILLER_15_166 ();
 sg13g2_fill_1 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_174 ();
 sg13g2_decap_4 FILLER_15_198 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_2 FILLER_15_209 ();
 sg13g2_fill_2 FILLER_15_226 ();
 sg13g2_fill_2 FILLER_15_254 ();
 sg13g2_fill_1 FILLER_15_267 ();
 sg13g2_decap_4 FILLER_15_271 ();
 sg13g2_fill_1 FILLER_15_275 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_fill_1 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_299 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_fill_2 FILLER_15_330 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_decap_4 FILLER_15_362 ();
 sg13g2_fill_1 FILLER_15_366 ();
 sg13g2_fill_2 FILLER_15_402 ();
 sg13g2_fill_1 FILLER_15_404 ();
 sg13g2_decap_8 FILLER_15_418 ();
 sg13g2_decap_4 FILLER_15_425 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_26 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_45 ();
 sg13g2_fill_1 FILLER_16_50 ();
 sg13g2_fill_1 FILLER_16_56 ();
 sg13g2_fill_2 FILLER_16_80 ();
 sg13g2_fill_1 FILLER_16_87 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_132 ();
 sg13g2_decap_4 FILLER_16_155 ();
 sg13g2_fill_1 FILLER_16_159 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_204 ();
 sg13g2_fill_1 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_215 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_decap_4 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_229 ();
 sg13g2_fill_1 FILLER_16_244 ();
 sg13g2_fill_1 FILLER_16_250 ();
 sg13g2_fill_1 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_265 ();
 sg13g2_fill_1 FILLER_16_271 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_288 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_299 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_fill_2 FILLER_16_315 ();
 sg13g2_fill_2 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_386 ();
 sg13g2_fill_2 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_26 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_1 FILLER_17_40 ();
 sg13g2_fill_1 FILLER_17_45 ();
 sg13g2_fill_1 FILLER_17_51 ();
 sg13g2_fill_1 FILLER_17_60 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_93 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_decap_4 FILLER_17_135 ();
 sg13g2_fill_1 FILLER_17_163 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_179 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_208 ();
 sg13g2_fill_1 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_fill_1 FILLER_17_237 ();
 sg13g2_fill_2 FILLER_17_245 ();
 sg13g2_decap_4 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_285 ();
 sg13g2_fill_1 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_325 ();
 sg13g2_fill_1 FILLER_17_327 ();
 sg13g2_fill_1 FILLER_17_352 ();
 sg13g2_fill_2 FILLER_17_357 ();
 sg13g2_fill_1 FILLER_17_365 ();
 sg13g2_fill_2 FILLER_17_392 ();
 sg13g2_fill_2 FILLER_17_402 ();
 sg13g2_fill_2 FILLER_18_38 ();
 sg13g2_fill_1 FILLER_18_40 ();
 sg13g2_fill_2 FILLER_18_44 ();
 sg13g2_fill_1 FILLER_18_57 ();
 sg13g2_fill_2 FILLER_18_62 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_fill_1 FILLER_18_81 ();
 sg13g2_fill_1 FILLER_18_86 ();
 sg13g2_fill_2 FILLER_18_92 ();
 sg13g2_fill_1 FILLER_18_98 ();
 sg13g2_fill_2 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_129 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_1 FILLER_18_137 ();
 sg13g2_decap_4 FILLER_18_155 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_fill_1 FILLER_18_195 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_fill_2 FILLER_18_255 ();
 sg13g2_fill_1 FILLER_18_281 ();
 sg13g2_fill_1 FILLER_18_286 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_1 FILLER_18_302 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_fill_2 FILLER_18_316 ();
 sg13g2_fill_2 FILLER_18_331 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_fill_1 FILLER_18_339 ();
 sg13g2_decap_4 FILLER_18_392 ();
 sg13g2_fill_1 FILLER_18_396 ();
 sg13g2_fill_1 FILLER_18_407 ();
 sg13g2_fill_2 FILLER_18_412 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_1 FILLER_19_5 ();
 sg13g2_fill_2 FILLER_19_10 ();
 sg13g2_fill_2 FILLER_19_16 ();
 sg13g2_fill_2 FILLER_19_22 ();
 sg13g2_fill_1 FILLER_19_24 ();
 sg13g2_fill_2 FILLER_19_30 ();
 sg13g2_fill_1 FILLER_19_32 ();
 sg13g2_fill_2 FILLER_19_37 ();
 sg13g2_decap_4 FILLER_19_52 ();
 sg13g2_decap_4 FILLER_19_71 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_121 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_fill_1 FILLER_19_208 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_232 ();
 sg13g2_fill_1 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_decap_4 FILLER_19_364 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_14 ();
 sg13g2_decap_4 FILLER_20_19 ();
 sg13g2_fill_1 FILLER_20_46 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_127 ();
 sg13g2_fill_1 FILLER_20_150 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_157 ();
 sg13g2_fill_2 FILLER_20_178 ();
 sg13g2_decap_4 FILLER_20_203 ();
 sg13g2_fill_2 FILLER_20_207 ();
 sg13g2_fill_1 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_236 ();
 sg13g2_fill_2 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_fill_2 FILLER_20_262 ();
 sg13g2_fill_1 FILLER_20_269 ();
 sg13g2_decap_4 FILLER_20_274 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_decap_4 FILLER_20_297 ();
 sg13g2_fill_2 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_fill_2 FILLER_20_394 ();
 sg13g2_fill_1 FILLER_20_396 ();
 sg13g2_fill_1 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_410 ();
 sg13g2_fill_1 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_fill_2 FILLER_20_427 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_12 ();
 sg13g2_fill_2 FILLER_21_17 ();
 sg13g2_fill_2 FILLER_21_24 ();
 sg13g2_fill_2 FILLER_21_30 ();
 sg13g2_decap_4 FILLER_21_37 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_fill_2 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_83 ();
 sg13g2_fill_2 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_104 ();
 sg13g2_fill_1 FILLER_21_110 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_137 ();
 sg13g2_fill_1 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_159 ();
 sg13g2_fill_2 FILLER_21_169 ();
 sg13g2_fill_1 FILLER_21_171 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_fill_1 FILLER_21_188 ();
 sg13g2_fill_2 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_fill_2 FILLER_21_207 ();
 sg13g2_fill_1 FILLER_21_213 ();
 sg13g2_decap_4 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_fill_1 FILLER_21_335 ();
 sg13g2_fill_1 FILLER_21_375 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_fill_1 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_5 ();
 sg13g2_fill_1 FILLER_22_32 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_fill_2 FILLER_22_51 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_fill_1 FILLER_22_86 ();
 sg13g2_decap_4 FILLER_22_92 ();
 sg13g2_decap_8 FILLER_22_100 ();
 sg13g2_fill_1 FILLER_22_107 ();
 sg13g2_fill_2 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_125 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_fill_1 FILLER_22_136 ();
 sg13g2_fill_2 FILLER_22_142 ();
 sg13g2_fill_2 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_fill_2 FILLER_22_187 ();
 sg13g2_decap_4 FILLER_22_195 ();
 sg13g2_fill_1 FILLER_22_199 ();
 sg13g2_decap_4 FILLER_22_217 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_decap_4 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_299 ();
 sg13g2_fill_2 FILLER_22_309 ();
 sg13g2_fill_2 FILLER_22_319 ();
 sg13g2_fill_2 FILLER_22_365 ();
 sg13g2_fill_2 FILLER_22_402 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_27 ();
 sg13g2_fill_1 FILLER_23_55 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_fill_1 FILLER_23_65 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_77 ();
 sg13g2_decap_4 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_87 ();
 sg13g2_fill_2 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_decap_4 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_decap_4 FILLER_23_132 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_decap_4 FILLER_23_152 ();
 sg13g2_fill_2 FILLER_23_156 ();
 sg13g2_fill_1 FILLER_23_166 ();
 sg13g2_decap_4 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_decap_8 FILLER_23_197 ();
 sg13g2_decap_4 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_234 ();
 sg13g2_decap_4 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_250 ();
 sg13g2_decap_8 FILLER_23_257 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_fill_1 FILLER_23_421 ();
 sg13g2_decap_4 FILLER_23_426 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_6 ();
 sg13g2_fill_1 FILLER_24_8 ();
 sg13g2_fill_1 FILLER_24_13 ();
 sg13g2_fill_2 FILLER_24_19 ();
 sg13g2_decap_8 FILLER_24_26 ();
 sg13g2_decap_4 FILLER_24_33 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_fill_1 FILLER_24_47 ();
 sg13g2_decap_4 FILLER_24_51 ();
 sg13g2_decap_8 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_fill_1 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_86 ();
 sg13g2_fill_1 FILLER_24_92 ();
 sg13g2_fill_2 FILLER_24_113 ();
 sg13g2_fill_1 FILLER_24_115 ();
 sg13g2_fill_2 FILLER_24_139 ();
 sg13g2_decap_4 FILLER_24_166 ();
 sg13g2_fill_2 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_216 ();
 sg13g2_decap_4 FILLER_24_233 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_263 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_fill_1 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_fill_2 FILLER_24_346 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_fill_2 FILLER_24_397 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_13 ();
 sg13g2_fill_1 FILLER_25_15 ();
 sg13g2_fill_1 FILLER_25_20 ();
 sg13g2_fill_1 FILLER_25_29 ();
 sg13g2_fill_1 FILLER_25_34 ();
 sg13g2_fill_1 FILLER_25_45 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_99 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_fill_2 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_123 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_decap_4 FILLER_25_188 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_2 FILLER_25_208 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_fill_2 FILLER_25_221 ();
 sg13g2_fill_2 FILLER_25_231 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_decap_4 FILLER_25_239 ();
 sg13g2_decap_8 FILLER_25_255 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_decap_4 FILLER_25_336 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_fill_1 FILLER_25_374 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_398 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_13 ();
 sg13g2_fill_2 FILLER_26_17 ();
 sg13g2_fill_2 FILLER_26_34 ();
 sg13g2_fill_1 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_66 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_83 ();
 sg13g2_fill_1 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_108 ();
 sg13g2_fill_1 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_128 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_215 ();
 sg13g2_fill_2 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_234 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_decap_4 FILLER_26_253 ();
 sg13g2_fill_1 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_269 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_4 FILLER_26_323 ();
 sg13g2_fill_2 FILLER_26_327 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_fill_2 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_394 ();
 sg13g2_fill_1 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_decap_8 FILLER_27_32 ();
 sg13g2_decap_4 FILLER_27_53 ();
 sg13g2_fill_2 FILLER_27_57 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_101 ();
 sg13g2_fill_1 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_fill_2 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_162 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_213 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_decap_4 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_276 ();
 sg13g2_decap_4 FILLER_27_282 ();
 sg13g2_decap_4 FILLER_27_290 ();
 sg13g2_fill_1 FILLER_27_305 ();
 sg13g2_fill_2 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_fill_2 FILLER_27_395 ();
 sg13g2_fill_1 FILLER_27_414 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_30 ();
 sg13g2_fill_2 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_54 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_69 ();
 sg13g2_decap_8 FILLER_28_76 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_94 ();
 sg13g2_fill_2 FILLER_28_103 ();
 sg13g2_fill_1 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_115 ();
 sg13g2_fill_2 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_128 ();
 sg13g2_fill_2 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_decap_4 FILLER_28_208 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_decap_4 FILLER_28_240 ();
 sg13g2_fill_2 FILLER_28_244 ();
 sg13g2_decap_4 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_decap_4 FILLER_28_274 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_fill_2 FILLER_28_318 ();
 sg13g2_fill_1 FILLER_28_325 ();
 sg13g2_fill_1 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_342 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_1 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_396 ();
 sg13g2_fill_1 FILLER_28_402 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_19 ();
 sg13g2_fill_2 FILLER_29_23 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_82 ();
 sg13g2_decap_4 FILLER_29_88 ();
 sg13g2_fill_2 FILLER_29_120 ();
 sg13g2_decap_4 FILLER_29_132 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_decap_4 FILLER_29_168 ();
 sg13g2_fill_1 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_fill_2 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_196 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_2 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_decap_4 FILLER_29_221 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_decap_4 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_fill_2 FILLER_29_373 ();
 sg13g2_fill_1 FILLER_29_379 ();
 sg13g2_fill_1 FILLER_29_385 ();
 sg13g2_fill_1 FILLER_29_395 ();
 sg13g2_fill_2 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_30 ();
 sg13g2_decap_4 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_71 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_decap_4 FILLER_30_92 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_fill_1 FILLER_30_118 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_145 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_156 ();
 sg13g2_decap_8 FILLER_30_173 ();
 sg13g2_decap_8 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_2 FILLER_30_314 ();
 sg13g2_fill_1 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_347 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_24 ();
 sg13g2_fill_1 FILLER_31_34 ();
 sg13g2_fill_1 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_54 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_121 ();
 sg13g2_fill_1 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_4 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_2 FILLER_31_396 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_26 ();
 sg13g2_decap_4 FILLER_32_45 ();
 sg13g2_decap_4 FILLER_32_54 ();
 sg13g2_decap_4 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_71 ();
 sg13g2_decap_8 FILLER_32_78 ();
 sg13g2_decap_8 FILLER_32_85 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_fill_2 FILLER_32_135 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_decap_8 FILLER_32_148 ();
 sg13g2_fill_2 FILLER_32_155 ();
 sg13g2_decap_8 FILLER_32_177 ();
 sg13g2_decap_8 FILLER_32_184 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_decap_4 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_239 ();
 sg13g2_decap_4 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_decap_4 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_fill_2 FILLER_32_335 ();
 sg13g2_decap_4 FILLER_32_380 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_fill_2 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_9 ();
 sg13g2_fill_2 FILLER_33_25 ();
 sg13g2_fill_1 FILLER_33_40 ();
 sg13g2_fill_1 FILLER_33_53 ();
 sg13g2_decap_4 FILLER_33_64 ();
 sg13g2_fill_2 FILLER_33_68 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_decap_8 FILLER_33_80 ();
 sg13g2_decap_4 FILLER_33_87 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_107 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_decap_4 FILLER_33_152 ();
 sg13g2_fill_1 FILLER_33_156 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_185 ();
 sg13g2_decap_8 FILLER_33_192 ();
 sg13g2_decap_8 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_227 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_261 ();
 sg13g2_decap_4 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_323 ();
 sg13g2_decap_4 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_fill_2 FILLER_33_384 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_423 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_fill_2 FILLER_34_15 ();
 sg13g2_fill_1 FILLER_34_17 ();
 sg13g2_fill_1 FILLER_34_22 ();
 sg13g2_decap_4 FILLER_34_31 ();
 sg13g2_fill_1 FILLER_34_45 ();
 sg13g2_fill_1 FILLER_34_50 ();
 sg13g2_fill_1 FILLER_34_59 ();
 sg13g2_fill_2 FILLER_34_93 ();
 sg13g2_fill_2 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_decap_8 FILLER_34_152 ();
 sg13g2_decap_4 FILLER_34_159 ();
 sg13g2_fill_2 FILLER_34_163 ();
 sg13g2_decap_8 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_200 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_decap_4 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_decap_4 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_35_38 ();
 sg13g2_fill_1 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_fill_1 FILLER_35_59 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_fill_1 FILLER_35_92 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_134 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_decap_4 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_229 ();
 sg13g2_decap_4 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_258 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_315 ();
 sg13g2_fill_1 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_fill_1 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_13 ();
 sg13g2_fill_1 FILLER_36_20 ();
 sg13g2_fill_2 FILLER_36_25 ();
 sg13g2_fill_2 FILLER_36_37 ();
 sg13g2_fill_1 FILLER_36_39 ();
 sg13g2_fill_2 FILLER_36_79 ();
 sg13g2_decap_8 FILLER_36_90 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_fill_2 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_fill_2 FILLER_36_137 ();
 sg13g2_fill_2 FILLER_36_162 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_fill_1 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_fill_2 FILLER_36_194 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_fill_2 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_238 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_decap_4 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_fill_2 FILLER_36_312 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_371 ();
 sg13g2_fill_2 FILLER_36_396 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_fill_1 FILLER_36_416 ();
 sg13g2_fill_1 FILLER_36_421 ();
 sg13g2_decap_4 FILLER_36_426 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_11 ();
 sg13g2_fill_1 FILLER_37_16 ();
 sg13g2_fill_2 FILLER_37_25 ();
 sg13g2_fill_1 FILLER_37_31 ();
 sg13g2_fill_2 FILLER_37_37 ();
 sg13g2_fill_2 FILLER_37_48 ();
 sg13g2_fill_1 FILLER_37_54 ();
 sg13g2_fill_1 FILLER_37_65 ();
 sg13g2_decap_4 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_106 ();
 sg13g2_fill_2 FILLER_37_136 ();
 sg13g2_decap_4 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_fill_1 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_179 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_339 ();
 sg13g2_fill_1 FILLER_37_386 ();
 sg13g2_fill_1 FILLER_37_391 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_fill_1 FILLER_38_26 ();
 sg13g2_fill_1 FILLER_38_31 ();
 sg13g2_fill_1 FILLER_38_40 ();
 sg13g2_fill_1 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_129 ();
 sg13g2_fill_1 FILLER_38_134 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_fill_2 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_223 ();
 sg13g2_decap_4 FILLER_38_231 ();
 sg13g2_fill_2 FILLER_38_279 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_291 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_fill_1 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_323 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_358 ();
 sg13g2_fill_2 FILLER_38_363 ();
 sg13g2_fill_1 FILLER_38_365 ();
 sg13g2_fill_2 FILLER_38_370 ();
 sg13g2_fill_1 FILLER_38_372 ();
 sg13g2_fill_1 FILLER_38_403 ();
endmodule
