module tt_um_urish_silife_max (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire clknet_leaf_0_clk;
 wire net1214;
 wire demo_mode;
 wire \demo_row_select[0] ;
 wire \demo_row_select[1] ;
 wire \demo_row_select[2] ;
 wire \demo_row_select[3] ;
 wire \demo_row_select[4] ;
 wire demo_step;
 wire demo_wr_en;
 wire \grid.cell_0_0.e ;
 wire \grid.cell_0_0.n ;
 wire \grid.cell_0_0.ne ;
 wire \grid.cell_0_0.nw ;
 wire \grid.cell_0_0.out ;
 wire \grid.cell_0_0.s ;
 wire \grid.cell_0_0.se ;
 wire \grid.cell_0_0.sw ;
 wire \grid.cell_0_0.w ;
 wire \grid.cell_0_1.e ;
 wire \grid.cell_0_1.ne ;
 wire \grid.cell_0_1.se ;
 wire \grid.cell_0_2.e ;
 wire \grid.cell_0_2.ne ;
 wire \grid.cell_0_2.se ;
 wire \grid.cell_0_3.e ;
 wire \grid.cell_0_3.ne ;
 wire \grid.cell_0_3.se ;
 wire \grid.cell_0_4.e ;
 wire \grid.cell_0_4.ne ;
 wire \grid.cell_0_4.se ;
 wire \grid.cell_0_5.e ;
 wire \grid.cell_0_5.ne ;
 wire \grid.cell_0_5.se ;
 wire \grid.cell_10_0.e ;
 wire \grid.cell_10_0.n ;
 wire \grid.cell_10_0.ne ;
 wire \grid.cell_10_0.nw ;
 wire \grid.cell_10_0.out ;
 wire \grid.cell_10_0.s ;
 wire \grid.cell_10_0.se ;
 wire \grid.cell_10_0.sw ;
 wire \grid.cell_10_0.w ;
 wire \grid.cell_10_1.e ;
 wire \grid.cell_10_1.ne ;
 wire \grid.cell_10_1.se ;
 wire \grid.cell_10_2.e ;
 wire \grid.cell_10_2.ne ;
 wire \grid.cell_10_2.se ;
 wire \grid.cell_10_3.e ;
 wire \grid.cell_10_3.ne ;
 wire \grid.cell_10_3.se ;
 wire \grid.cell_10_4.e ;
 wire \grid.cell_10_4.ne ;
 wire \grid.cell_10_4.se ;
 wire \grid.cell_10_5.e ;
 wire \grid.cell_10_5.ne ;
 wire \grid.cell_10_5.se ;
 wire \grid.cell_11_0.s ;
 wire \grid.cell_11_0.se ;
 wire \grid.cell_11_0.sw ;
 wire \grid.cell_11_1.se ;
 wire \grid.cell_11_2.se ;
 wire \grid.cell_11_3.se ;
 wire \grid.cell_11_4.se ;
 wire \grid.cell_11_5.se ;
 wire \grid.cell_12_0.s ;
 wire \grid.cell_12_0.se ;
 wire \grid.cell_12_0.sw ;
 wire \grid.cell_12_1.se ;
 wire \grid.cell_12_2.se ;
 wire \grid.cell_12_3.se ;
 wire \grid.cell_12_4.se ;
 wire \grid.cell_12_5.se ;
 wire \grid.cell_13_0.s ;
 wire \grid.cell_13_0.se ;
 wire \grid.cell_13_0.sw ;
 wire \grid.cell_13_1.se ;
 wire \grid.cell_13_2.se ;
 wire \grid.cell_13_3.se ;
 wire \grid.cell_13_4.se ;
 wire \grid.cell_13_5.se ;
 wire \grid.cell_14_0.s ;
 wire \grid.cell_14_0.se ;
 wire \grid.cell_14_0.sw ;
 wire \grid.cell_14_1.se ;
 wire \grid.cell_14_2.se ;
 wire \grid.cell_14_3.se ;
 wire \grid.cell_14_4.se ;
 wire \grid.cell_14_5.se ;
 wire \grid.cell_15_0.s ;
 wire \grid.cell_15_0.se ;
 wire \grid.cell_15_0.sw ;
 wire \grid.cell_15_1.se ;
 wire \grid.cell_15_2.se ;
 wire \grid.cell_15_3.se ;
 wire \grid.cell_15_4.se ;
 wire \grid.cell_15_5.se ;
 wire \grid.cell_16_0.s ;
 wire \grid.cell_16_0.se ;
 wire \grid.cell_16_0.sw ;
 wire \grid.cell_16_1.se ;
 wire \grid.cell_16_2.se ;
 wire \grid.cell_16_3.se ;
 wire \grid.cell_16_4.se ;
 wire \grid.cell_16_5.se ;
 wire \grid.cell_17_0.s ;
 wire \grid.cell_17_0.se ;
 wire \grid.cell_17_0.sw ;
 wire \grid.cell_17_1.se ;
 wire \grid.cell_17_2.se ;
 wire \grid.cell_17_3.se ;
 wire \grid.cell_17_4.se ;
 wire \grid.cell_17_5.se ;
 wire \grid.cell_18_0.s ;
 wire \grid.cell_18_0.se ;
 wire \grid.cell_18_0.sw ;
 wire \grid.cell_18_1.se ;
 wire \grid.cell_18_2.se ;
 wire \grid.cell_18_3.se ;
 wire \grid.cell_18_4.se ;
 wire \grid.cell_18_5.se ;
 wire \grid.cell_19_0.s ;
 wire \grid.cell_19_0.se ;
 wire \grid.cell_19_0.sw ;
 wire \grid.cell_19_1.se ;
 wire \grid.cell_19_2.se ;
 wire \grid.cell_19_3.se ;
 wire \grid.cell_19_4.se ;
 wire \grid.cell_19_5.se ;
 wire \grid.cell_1_0.s ;
 wire \grid.cell_1_0.se ;
 wire \grid.cell_1_0.sw ;
 wire \grid.cell_1_1.se ;
 wire \grid.cell_1_2.se ;
 wire \grid.cell_1_3.se ;
 wire \grid.cell_1_4.se ;
 wire \grid.cell_1_5.se ;
 wire \grid.cell_20_0.s ;
 wire \grid.cell_20_0.se ;
 wire \grid.cell_20_0.sw ;
 wire \grid.cell_20_1.se ;
 wire \grid.cell_20_2.se ;
 wire \grid.cell_20_3.se ;
 wire \grid.cell_20_4.se ;
 wire \grid.cell_20_5.se ;
 wire \grid.cell_21_0.s ;
 wire \grid.cell_21_0.se ;
 wire \grid.cell_21_0.sw ;
 wire \grid.cell_21_1.se ;
 wire \grid.cell_21_2.se ;
 wire \grid.cell_21_3.se ;
 wire \grid.cell_21_4.se ;
 wire \grid.cell_21_5.se ;
 wire \grid.cell_22_0.s ;
 wire \grid.cell_22_0.se ;
 wire \grid.cell_22_0.sw ;
 wire \grid.cell_22_1.se ;
 wire \grid.cell_22_2.se ;
 wire \grid.cell_22_3.se ;
 wire \grid.cell_22_4.se ;
 wire \grid.cell_22_5.se ;
 wire \grid.cell_23_0.s ;
 wire \grid.cell_23_0.se ;
 wire \grid.cell_23_0.sw ;
 wire \grid.cell_23_1.se ;
 wire \grid.cell_23_2.se ;
 wire \grid.cell_23_3.se ;
 wire \grid.cell_23_4.se ;
 wire \grid.cell_23_5.se ;
 wire \grid.cell_24_0.s ;
 wire \grid.cell_24_0.se ;
 wire \grid.cell_24_0.sw ;
 wire \grid.cell_24_1.se ;
 wire \grid.cell_24_2.se ;
 wire \grid.cell_24_3.se ;
 wire \grid.cell_24_4.se ;
 wire \grid.cell_24_5.se ;
 wire \grid.cell_25_0.s ;
 wire \grid.cell_25_0.se ;
 wire \grid.cell_25_0.sw ;
 wire \grid.cell_25_1.se ;
 wire \grid.cell_25_2.se ;
 wire \grid.cell_25_3.se ;
 wire \grid.cell_25_4.se ;
 wire \grid.cell_25_5.se ;
 wire \grid.cell_26_0.s ;
 wire \grid.cell_26_0.se ;
 wire \grid.cell_26_0.sw ;
 wire \grid.cell_26_1.se ;
 wire \grid.cell_26_2.se ;
 wire \grid.cell_26_3.se ;
 wire \grid.cell_26_4.se ;
 wire \grid.cell_26_5.se ;
 wire \grid.cell_27_0.s ;
 wire \grid.cell_27_0.se ;
 wire \grid.cell_27_0.sw ;
 wire \grid.cell_27_1.se ;
 wire \grid.cell_27_2.se ;
 wire \grid.cell_27_3.se ;
 wire \grid.cell_27_4.se ;
 wire \grid.cell_27_5.se ;
 wire \grid.cell_28_0.s ;
 wire \grid.cell_28_0.se ;
 wire \grid.cell_28_0.sw ;
 wire \grid.cell_28_1.se ;
 wire \grid.cell_28_2.se ;
 wire \grid.cell_28_3.se ;
 wire \grid.cell_28_4.se ;
 wire \grid.cell_28_5.se ;
 wire \grid.cell_29_0.s ;
 wire \grid.cell_29_0.se ;
 wire \grid.cell_29_0.sw ;
 wire \grid.cell_29_1.se ;
 wire \grid.cell_29_2.se ;
 wire \grid.cell_29_3.se ;
 wire \grid.cell_29_4.se ;
 wire \grid.cell_29_5.se ;
 wire \grid.cell_2_0.s ;
 wire \grid.cell_2_0.se ;
 wire \grid.cell_2_0.sw ;
 wire \grid.cell_2_1.se ;
 wire \grid.cell_2_2.se ;
 wire \grid.cell_2_3.se ;
 wire \grid.cell_2_4.se ;
 wire \grid.cell_2_5.se ;
 wire \grid.cell_3_0.s ;
 wire \grid.cell_3_0.se ;
 wire \grid.cell_3_0.sw ;
 wire \grid.cell_3_1.se ;
 wire \grid.cell_3_2.se ;
 wire \grid.cell_3_3.se ;
 wire \grid.cell_3_4.se ;
 wire \grid.cell_3_5.se ;
 wire \grid.cell_4_0.s ;
 wire \grid.cell_4_0.se ;
 wire \grid.cell_4_0.sw ;
 wire \grid.cell_4_1.se ;
 wire \grid.cell_4_2.se ;
 wire \grid.cell_4_3.se ;
 wire \grid.cell_4_4.se ;
 wire \grid.cell_4_5.se ;
 wire \grid.cell_5_0.s ;
 wire \grid.cell_5_0.se ;
 wire \grid.cell_5_0.sw ;
 wire \grid.cell_5_1.se ;
 wire \grid.cell_5_2.se ;
 wire \grid.cell_5_3.se ;
 wire \grid.cell_5_4.se ;
 wire \grid.cell_5_5.se ;
 wire \grid.cell_6_0.s ;
 wire \grid.cell_6_0.se ;
 wire \grid.cell_6_0.sw ;
 wire \grid.cell_6_1.se ;
 wire \grid.cell_6_2.se ;
 wire \grid.cell_6_3.se ;
 wire \grid.cell_6_4.se ;
 wire \grid.cell_6_5.se ;
 wire \grid.cell_7_0.s ;
 wire \grid.cell_7_0.se ;
 wire \grid.cell_7_0.sw ;
 wire \grid.cell_7_1.se ;
 wire \grid.cell_7_2.se ;
 wire \grid.cell_7_3.se ;
 wire \grid.cell_7_4.se ;
 wire \grid.cell_7_5.se ;
 wire \grid.row_select2[0] ;
 wire \grid.row_select2[1] ;
 wire \grid.row_select2[2] ;
 wire \grid.row_select2[3] ;
 wire \grid.row_select2[4] ;
 wire \max7219.init_index[0] ;
 wire \max7219.init_index[1] ;
 wire \max7219.load_row ;
 wire \max7219.max7219_enabled ;
 wire \max7219.max7219_row[0] ;
 wire \max7219.max7219_row[1] ;
 wire \max7219.max7219_row[2] ;
 wire \max7219.o_cs ;
 wire \max7219.o_mosi ;
 wire \max7219.o_sck ;
 wire \max7219.row_data[0] ;
 wire \max7219.row_data[1] ;
 wire \max7219.row_data[2] ;
 wire \max7219.row_data[3] ;
 wire \max7219.row_data[4] ;
 wire \max7219.row_data[5] ;
 wire \max7219.row_data[6] ;
 wire \max7219.row_data[7] ;
 wire \max7219.spi_busy ;
 wire \max7219.spi_start ;
 wire \max7219.spim.bit_index[0] ;
 wire \max7219.spim.bit_index[1] ;
 wire \max7219.spim.bit_index[2] ;
 wire \max7219.spim.bit_index[3] ;
 wire \max7219.spim.clk_count[0] ;
 wire \max7219.spim.clk_count[1] ;
 wire \max7219.spim.finish ;
 wire \max7219.state[0] ;
 wire \max7219.state[1] ;
 wire \max7219.state[2] ;
 wire \max7219.state[3] ;
 wire prev_rst_n;
 wire \silife_demo_inst.counter[0] ;
 wire \silife_demo_inst.counter[10] ;
 wire \silife_demo_inst.counter[11] ;
 wire \silife_demo_inst.counter[12] ;
 wire \silife_demo_inst.counter[13] ;
 wire \silife_demo_inst.counter[14] ;
 wire \silife_demo_inst.counter[15] ;
 wire \silife_demo_inst.counter[16] ;
 wire \silife_demo_inst.counter[17] ;
 wire \silife_demo_inst.counter[18] ;
 wire \silife_demo_inst.counter[19] ;
 wire \silife_demo_inst.counter[1] ;
 wire \silife_demo_inst.counter[20] ;
 wire \silife_demo_inst.counter[21] ;
 wire \silife_demo_inst.counter[22] ;
 wire \silife_demo_inst.counter[23] ;
 wire \silife_demo_inst.counter[24] ;
 wire \silife_demo_inst.counter[25] ;
 wire \silife_demo_inst.counter[26] ;
 wire \silife_demo_inst.counter[27] ;
 wire \silife_demo_inst.counter[28] ;
 wire \silife_demo_inst.counter[29] ;
 wire \silife_demo_inst.counter[2] ;
 wire \silife_demo_inst.counter[30] ;
 wire \silife_demo_inst.counter[31] ;
 wire \silife_demo_inst.counter[3] ;
 wire \silife_demo_inst.counter[4] ;
 wire \silife_demo_inst.counter[5] ;
 wire \silife_demo_inst.counter[6] ;
 wire \silife_demo_inst.counter[7] ;
 wire \silife_demo_inst.counter[8] ;
 wire \silife_demo_inst.counter[9] ;
 wire \silife_demo_inst.init_done ;
 wire wr_available;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net1549;

 sg13g2_buf_2 _13376_ (.A(net1),
    .X(_12956_));
 sg13g2_buf_2 _13377_ (.A(_12956_),
    .X(_12967_));
 sg13g2_buf_1 _13378_ (.A(net1197),
    .X(_12977_));
 sg13g2_buf_1 _13379_ (.A(net1060),
    .X(_12988_));
 sg13g2_buf_1 _13380_ (.A(_12988_),
    .X(_12999_));
 sg13g2_buf_2 _13381_ (.A(ui_in[5]),
    .X(_13010_));
 sg13g2_buf_2 _13382_ (.A(\max7219.spi_busy ),
    .X(_13020_));
 sg13g2_nor2_1 _13383_ (.A(\max7219.spi_start ),
    .B(_13020_),
    .Y(_13031_));
 sg13g2_and2_1 _13384_ (.A(_13010_),
    .B(_13031_),
    .X(_13042_));
 sg13g2_buf_1 _13385_ (.A(_13042_),
    .X(_13053_));
 sg13g2_buf_1 _13386_ (.A(\max7219.state[0] ),
    .X(_13063_));
 sg13g2_buf_1 _13387_ (.A(net1197),
    .X(_13074_));
 sg13g2_nand2_1 _13388_ (.Y(_13085_),
    .A(net1059),
    .B(_13010_));
 sg13g2_nor2_1 _13389_ (.A(_13063_),
    .B(_13085_),
    .Y(_13096_));
 sg13g2_a21oi_1 _13390_ (.A1(net378),
    .A2(net377),
    .Y(_00000_),
    .B1(_13096_));
 sg13g2_buf_1 _13391_ (.A(\max7219.o_cs ),
    .X(_13116_));
 sg13g2_buf_1 _13392_ (.A(\grid.row_select2[3] ),
    .X(_13127_));
 sg13g2_buf_1 _13393_ (.A(\grid.row_select2[4] ),
    .X(_13138_));
 sg13g2_nand2_1 _13394_ (.Y(_13149_),
    .A(net1196),
    .B(_13138_));
 sg13g2_buf_2 _13395_ (.A(_13149_),
    .X(_13159_));
 sg13g2_nor3_2 _13396_ (.A(\max7219.spi_start ),
    .B(_13020_),
    .C(_13159_),
    .Y(_13170_));
 sg13g2_nand2_1 _13397_ (.Y(_13181_),
    .A(_13116_),
    .B(_13170_));
 sg13g2_buf_1 _13398_ (.A(\max7219.state[1] ),
    .X(_13191_));
 sg13g2_buf_1 _13399_ (.A(_13191_),
    .X(_13202_));
 sg13g2_buf_1 _13400_ (.A(\max7219.max7219_row[2] ),
    .X(_13213_));
 sg13g2_inv_1 _13401_ (.Y(_13224_),
    .A(_13213_));
 sg13g2_buf_1 _13402_ (.A(\max7219.max7219_row[1] ),
    .X(_13235_));
 sg13g2_buf_1 _13403_ (.A(\max7219.max7219_row[0] ),
    .X(_13246_));
 sg13g2_nand2_1 _13404_ (.Y(_13256_),
    .A(_13235_),
    .B(net1195));
 sg13g2_nor3_1 _13405_ (.A(_13224_),
    .B(\max7219.max7219_enabled ),
    .C(_13256_),
    .Y(_13267_));
 sg13g2_nand4_1 _13406_ (.B(_13010_),
    .C(net1058),
    .A(net716),
    .Y(_13278_),
    .D(_13267_));
 sg13g2_buf_1 _13407_ (.A(\max7219.state[3] ),
    .X(_13289_));
 sg13g2_nor2_2 _13408_ (.A(_13116_),
    .B(_13159_),
    .Y(_13300_));
 sg13g2_nand3_1 _13409_ (.B(net377),
    .C(_13300_),
    .A(net1059),
    .Y(_00606_));
 sg13g2_o21ai_1 _13410_ (.B1(_00606_),
    .Y(_00616_),
    .A1(_13085_),
    .A2(_13170_));
 sg13g2_nand2_1 _13411_ (.Y(_00627_),
    .A(_13289_),
    .B(_00616_));
 sg13g2_o21ai_1 _13412_ (.B1(_00627_),
    .Y(_00003_),
    .A1(_13181_),
    .A2(_13278_));
 sg13g2_inv_2 _13413_ (.Y(_00648_),
    .A(_12956_));
 sg13g2_buf_1 _13414_ (.A(_00648_),
    .X(_00659_));
 sg13g2_buf_1 _13415_ (.A(net1057),
    .X(_00669_));
 sg13g2_nand2b_1 _13416_ (.Y(_00680_),
    .B(net377),
    .A_N(_00024_));
 sg13g2_buf_1 _13417_ (.A(_00025_),
    .X(_00691_));
 sg13g2_nand2b_1 _13418_ (.Y(_00702_),
    .B(_13170_),
    .A_N(_00691_));
 sg13g2_inv_1 _13419_ (.Y(_00712_),
    .A(_13116_));
 sg13g2_buf_2 _13420_ (.A(\max7219.init_index[0] ),
    .X(_00723_));
 sg13g2_buf_1 _13421_ (.A(\max7219.init_index[1] ),
    .X(_00734_));
 sg13g2_and2_1 _13422_ (.A(_00723_),
    .B(_00734_),
    .X(_00745_));
 sg13g2_buf_1 _13423_ (.A(_00745_),
    .X(_00755_));
 sg13g2_nor2_1 _13424_ (.A(_00712_),
    .B(_00755_),
    .Y(_00766_));
 sg13g2_buf_1 _13425_ (.A(_12956_),
    .X(_00777_));
 sg13g2_buf_1 _13426_ (.A(net1194),
    .X(_00788_));
 sg13g2_buf_1 _13427_ (.A(\max7219.state[2] ),
    .X(_00798_));
 sg13g2_and3_1 _13428_ (.X(_00809_),
    .A(net1056),
    .B(_13010_),
    .C(_00798_));
 sg13g2_o21ai_1 _13429_ (.B1(_00809_),
    .Y(_00820_),
    .A1(_00702_),
    .A2(_00766_));
 sg13g2_o21ai_1 _13430_ (.B1(_00820_),
    .Y(_00002_),
    .A1(net715),
    .A2(_00680_));
 sg13g2_and3_1 _13431_ (.X(_00840_),
    .A(net1193),
    .B(_00723_),
    .C(_00734_));
 sg13g2_nor2_1 _13432_ (.A(_13289_),
    .B(_00840_),
    .Y(_00851_));
 sg13g2_or2_1 _13433_ (.X(_00862_),
    .B(_00851_),
    .A(_13181_));
 sg13g2_nand3b_1 _13434_ (.B(_13170_),
    .C(_13267_),
    .Y(_00872_),
    .A_N(_00691_));
 sg13g2_nand2_1 _13435_ (.Y(_00883_),
    .A(net1058),
    .B(_00872_));
 sg13g2_a21oi_1 _13436_ (.A1(_00862_),
    .A2(_00883_),
    .Y(_00001_),
    .B1(_13085_));
 sg13g2_buf_1 _13437_ (.A(\max7219.spim.clk_count[1] ),
    .X(_00904_));
 sg13g2_nand2b_1 _13438_ (.Y(_00915_),
    .B(net1194),
    .A_N(\max7219.spim.finish ));
 sg13g2_buf_1 _13439_ (.A(_00915_),
    .X(_00926_));
 sg13g2_buf_2 _13440_ (.A(\max7219.spim.bit_index[2] ),
    .X(_00936_));
 sg13g2_buf_1 _13441_ (.A(\max7219.spim.bit_index[3] ),
    .X(_00947_));
 sg13g2_nand3_1 _13442_ (.B(_00947_),
    .C(\max7219.o_sck ),
    .A(_00936_),
    .Y(_00958_));
 sg13g2_buf_1 _13443_ (.A(\max7219.spim.clk_count[0] ),
    .X(_00969_));
 sg13g2_buf_1 _13444_ (.A(\max7219.spim.bit_index[0] ),
    .X(_00979_));
 sg13g2_buf_1 _13445_ (.A(_00979_),
    .X(_00990_));
 sg13g2_buf_1 _13446_ (.A(\max7219.spim.bit_index[1] ),
    .X(_01001_));
 sg13g2_nand4_1 _13447_ (.B(_00969_),
    .C(net1055),
    .A(_13020_),
    .Y(_01012_),
    .D(net1192));
 sg13g2_nor4_1 _13448_ (.A(_00904_),
    .B(_00926_),
    .C(_00958_),
    .D(_01012_),
    .Y(_01022_));
 sg13g2_a21o_1 _13449_ (.A2(\max7219.spim.finish ),
    .A1(net715),
    .B1(_01022_),
    .X(_00561_));
 sg13g2_buf_2 _13450_ (.A(demo_mode),
    .X(_01043_));
 sg13g2_buf_1 _13451_ (.A(net1197),
    .X(_01053_));
 sg13g2_buf_1 _13452_ (.A(_01053_),
    .X(_01064_));
 sg13g2_nand2_1 _13453_ (.Y(_01075_),
    .A(net1191),
    .B(net714));
 sg13g2_buf_1 _13454_ (.A(\silife_demo_inst.counter[19] ),
    .X(_01086_));
 sg13g2_buf_1 _13455_ (.A(\silife_demo_inst.counter[18] ),
    .X(_01096_));
 sg13g2_and4_1 _13456_ (.A(_01086_),
    .B(_01096_),
    .C(\silife_demo_inst.counter[21] ),
    .D(\silife_demo_inst.counter[20] ),
    .X(_01107_));
 sg13g2_buf_1 _13457_ (.A(\silife_demo_inst.counter[10] ),
    .X(_01118_));
 sg13g2_buf_1 _13458_ (.A(\silife_demo_inst.counter[24] ),
    .X(_01129_));
 sg13g2_buf_1 _13459_ (.A(\silife_demo_inst.counter[27] ),
    .X(_01139_));
 sg13g2_nor4_1 _13460_ (.A(\silife_demo_inst.counter[8] ),
    .B(_01118_),
    .C(_01129_),
    .D(_01139_),
    .Y(_01150_));
 sg13g2_buf_1 _13461_ (.A(\silife_demo_inst.counter[26] ),
    .X(_01161_));
 sg13g2_buf_2 _13462_ (.A(\silife_demo_inst.counter[29] ),
    .X(_01172_));
 sg13g2_nor4_1 _13463_ (.A(_01161_),
    .B(_01172_),
    .C(\silife_demo_inst.counter[28] ),
    .D(\silife_demo_inst.counter[31] ),
    .Y(_01182_));
 sg13g2_nand2_1 _13464_ (.Y(_01193_),
    .A(_01150_),
    .B(_01182_));
 sg13g2_buf_1 _13465_ (.A(\silife_demo_inst.counter[1] ),
    .X(_01204_));
 sg13g2_buf_1 _13466_ (.A(\silife_demo_inst.counter[6] ),
    .X(_01215_));
 sg13g2_nand2_1 _13467_ (.Y(_01225_),
    .A(_01204_),
    .B(_01215_));
 sg13g2_nor4_1 _13468_ (.A(\silife_demo_inst.counter[9] ),
    .B(\silife_demo_inst.counter[30] ),
    .C(_01193_),
    .D(_01225_),
    .Y(_01236_));
 sg13g2_buf_1 _13469_ (.A(\silife_demo_inst.counter[23] ),
    .X(_01247_));
 sg13g2_buf_1 _13470_ (.A(\silife_demo_inst.counter[17] ),
    .X(_01258_));
 sg13g2_buf_1 _13471_ (.A(\silife_demo_inst.counter[16] ),
    .X(_01268_));
 sg13g2_nand2b_1 _13472_ (.Y(_01279_),
    .B(_01268_),
    .A_N(_01258_));
 sg13g2_inv_1 _13473_ (.Y(_01290_),
    .A(\silife_demo_inst.counter[11] ));
 sg13g2_buf_1 _13474_ (.A(\silife_demo_inst.counter[13] ),
    .X(_01301_));
 sg13g2_buf_1 _13475_ (.A(\silife_demo_inst.counter[12] ),
    .X(_01312_));
 sg13g2_or4_1 _13476_ (.A(_01290_),
    .B(_01301_),
    .C(_01312_),
    .D(\silife_demo_inst.counter[15] ),
    .X(_01322_));
 sg13g2_nor4_1 _13477_ (.A(_01247_),
    .B(\silife_demo_inst.counter[25] ),
    .C(_01279_),
    .D(_01322_),
    .Y(_01333_));
 sg13g2_buf_1 _13478_ (.A(\silife_demo_inst.counter[14] ),
    .X(_01344_));
 sg13g2_buf_1 _13479_ (.A(\silife_demo_inst.counter[22] ),
    .X(_01354_));
 sg13g2_buf_2 _13480_ (.A(\silife_demo_inst.counter[5] ),
    .X(_01365_));
 sg13g2_and2_1 _13481_ (.A(\silife_demo_inst.counter[3] ),
    .B(\silife_demo_inst.counter[4] ),
    .X(_01376_));
 sg13g2_buf_1 _13482_ (.A(_01376_),
    .X(_01386_));
 sg13g2_nand3_1 _13483_ (.B(\silife_demo_inst.counter[7] ),
    .C(_01386_),
    .A(_01365_),
    .Y(_01397_));
 sg13g2_buf_8 _13484_ (.A(\silife_demo_inst.counter[0] ),
    .X(_01408_));
 sg13g2_nand2_1 _13485_ (.Y(_01418_),
    .A(_01408_),
    .B(\silife_demo_inst.counter[2] ));
 sg13g2_nor4_1 _13486_ (.A(_01344_),
    .B(_01354_),
    .C(_01397_),
    .D(_01418_),
    .Y(_01429_));
 sg13g2_nand4_1 _13487_ (.B(_01236_),
    .C(_01333_),
    .A(_01107_),
    .Y(_01440_),
    .D(_01429_));
 sg13g2_nand2_1 _13488_ (.Y(_01451_),
    .A(demo_step),
    .B(_01075_));
 sg13g2_o21ai_1 _13489_ (.B1(_01451_),
    .Y(_00603_),
    .A1(_01075_),
    .A2(_01440_));
 sg13g2_buf_2 _13490_ (.A(demo_wr_en),
    .X(_01471_));
 sg13g2_buf_8 _13491_ (.A(_01471_),
    .X(_01482_));
 sg13g2_buf_1 _13492_ (.A(net1053),
    .X(_01492_));
 sg13g2_buf_1 _13493_ (.A(_01492_),
    .X(_01503_));
 sg13g2_buf_1 _13494_ (.A(\demo_row_select[3] ),
    .X(_01514_));
 sg13g2_buf_1 _13495_ (.A(net1190),
    .X(_01525_));
 sg13g2_buf_2 _13496_ (.A(\demo_row_select[4] ),
    .X(_01536_));
 sg13g2_inv_1 _13497_ (.Y(_01547_),
    .A(_01536_));
 sg13g2_nor2_1 _13498_ (.A(net1052),
    .B(_01547_),
    .Y(_01557_));
 sg13g2_buf_2 _13499_ (.A(ui_in[0]),
    .X(_01568_));
 sg13g2_buf_1 _13500_ (.A(_01568_),
    .X(_01579_));
 sg13g2_buf_1 _13501_ (.A(net1189),
    .X(_01590_));
 sg13g2_buf_1 _13502_ (.A(\demo_row_select[0] ),
    .X(_01601_));
 sg13g2_buf_1 _13503_ (.A(_01601_),
    .X(_01612_));
 sg13g2_buf_2 _13504_ (.A(\demo_row_select[2] ),
    .X(_01622_));
 sg13g2_buf_1 _13505_ (.A(_00020_),
    .X(_01633_));
 sg13g2_nor2_1 _13506_ (.A(_01622_),
    .B(_01633_),
    .Y(_01644_));
 sg13g2_buf_2 _13507_ (.A(_01644_),
    .X(_01655_));
 sg13g2_buf_1 _13508_ (.A(_01622_),
    .X(_01666_));
 sg13g2_buf_1 _13509_ (.A(net1049),
    .X(_01676_));
 sg13g2_nand3_1 _13510_ (.B(net712),
    .C(_01633_),
    .A(net1189),
    .Y(_01687_));
 sg13g2_nor2b_1 _13511_ (.A(_01655_),
    .B_N(_01687_),
    .Y(_01698_));
 sg13g2_a21oi_1 _13512_ (.A1(_01590_),
    .A2(net1050),
    .Y(_01709_),
    .B1(_01698_));
 sg13g2_buf_1 _13513_ (.A(\demo_row_select[1] ),
    .X(_01720_));
 sg13g2_xor2_1 _13514_ (.B(net1187),
    .A(net1188),
    .X(_01731_));
 sg13g2_buf_1 _13515_ (.A(_01536_),
    .X(_01742_));
 sg13g2_buf_1 _13516_ (.A(_00021_),
    .X(_01752_));
 sg13g2_nor4_1 _13517_ (.A(net1051),
    .B(net1048),
    .C(_01752_),
    .D(_00019_),
    .Y(_01763_));
 sg13g2_a22oi_1 _13518_ (.Y(_01774_),
    .B1(_01731_),
    .B2(_01763_),
    .A2(_01709_),
    .A1(_01557_));
 sg13g2_nor2_1 _13519_ (.A(net713),
    .B(net8),
    .Y(_01784_));
 sg13g2_a21oi_1 _13520_ (.A1(net376),
    .A2(_01774_),
    .Y(_01795_),
    .B1(_01784_));
 sg13g2_buf_2 _13521_ (.A(_01795_),
    .X(_01806_));
 sg13g2_inv_1 _13522_ (.Y(_01817_),
    .A(_01806_));
 sg13g2_nor2_1 _13523_ (.A(_01622_),
    .B(net1190),
    .Y(_01827_));
 sg13g2_nor2_1 _13524_ (.A(net1053),
    .B(net3),
    .Y(_01838_));
 sg13g2_inv_1 _13525_ (.Y(_01849_),
    .A(net4));
 sg13g2_a22oi_1 _13526_ (.Y(_01860_),
    .B1(_01838_),
    .B2(_01849_),
    .A2(_01827_),
    .A1(net1053));
 sg13g2_buf_1 _13527_ (.A(_01860_),
    .X(_01870_));
 sg13g2_nand2_1 _13528_ (.Y(_01881_),
    .A(_01471_),
    .B(_00017_));
 sg13g2_o21ai_1 _13529_ (.B1(_01881_),
    .Y(_01892_),
    .A1(net1053),
    .A2(net5));
 sg13g2_buf_1 _13530_ (.A(_01892_),
    .X(_01903_));
 sg13g2_buf_1 _13531_ (.A(_01903_),
    .X(_01913_));
 sg13g2_mux2_1 _13532_ (.A0(_01568_),
    .A1(\demo_row_select[0] ),
    .S(_01482_),
    .X(_01924_));
 sg13g2_buf_2 _13533_ (.A(_01924_),
    .X(_01935_));
 sg13g2_mux2_1 _13534_ (.A0(net2),
    .A1(\demo_row_select[1] ),
    .S(_01471_),
    .X(_01946_));
 sg13g2_buf_1 _13535_ (.A(_01946_),
    .X(_01956_));
 sg13g2_nor2_1 _13536_ (.A(_01935_),
    .B(_01956_),
    .Y(_01967_));
 sg13g2_nand2_1 _13537_ (.Y(_01978_),
    .A(net177),
    .B(_01967_));
 sg13g2_buf_2 _13538_ (.A(_01978_),
    .X(_01989_));
 sg13g2_nand2_1 _13539_ (.Y(_02000_),
    .A(wr_available),
    .B(net7));
 sg13g2_and2_1 _13540_ (.A(_00018_),
    .B(_02000_),
    .X(_02011_));
 sg13g2_buf_2 _13541_ (.A(_02011_),
    .X(_02021_));
 sg13g2_buf_1 _13542_ (.A(_02021_),
    .X(_02032_));
 sg13g2_buf_2 _13543_ (.A(net375),
    .X(_02043_));
 sg13g2_nor3_2 _13544_ (.A(_01870_),
    .B(_01989_),
    .C(net176),
    .Y(_02054_));
 sg13g2_nand2_2 _13545_ (.Y(_02065_),
    .A(net714),
    .B(_02054_));
 sg13g2_buf_2 _13546_ (.A(\grid.cell_0_0.se ),
    .X(_02076_));
 sg13g2_inv_2 _13547_ (.Y(_02087_),
    .A(_02076_));
 sg13g2_buf_1 _13548_ (.A(_00217_),
    .X(_02097_));
 sg13g2_buf_1 _13549_ (.A(_02097_),
    .X(_02108_));
 sg13g2_buf_1 _13550_ (.A(\grid.cell_0_0.e ),
    .X(_02119_));
 sg13g2_buf_1 _13551_ (.A(net1186),
    .X(_02130_));
 sg13g2_o21ai_1 _13552_ (.B1(net1046),
    .Y(_02140_),
    .A1(_02087_),
    .A2(net1047));
 sg13g2_buf_1 _13553_ (.A(_02076_),
    .X(_02151_));
 sg13g2_buf_1 _13554_ (.A(net1045),
    .X(_02162_));
 sg13g2_buf_1 _13555_ (.A(\grid.cell_0_0.s ),
    .X(_02173_));
 sg13g2_inv_2 _13556_ (.Y(_02183_),
    .A(net1185));
 sg13g2_buf_1 _13557_ (.A(\grid.cell_0_0.ne ),
    .X(_02194_));
 sg13g2_buf_2 _13558_ (.A(\grid.cell_0_0.nw ),
    .X(_02205_));
 sg13g2_xor2_1 _13559_ (.B(_02205_),
    .A(_02194_),
    .X(_02216_));
 sg13g2_buf_2 _13560_ (.A(_02216_),
    .X(_02226_));
 sg13g2_buf_1 _13561_ (.A(\grid.cell_0_0.w ),
    .X(_02237_));
 sg13g2_buf_1 _13562_ (.A(\grid.cell_0_0.sw ),
    .X(_02248_));
 sg13g2_xnor2_1 _13563_ (.Y(_02259_),
    .A(_02237_),
    .B(_02248_));
 sg13g2_xnor2_1 _13564_ (.Y(_02269_),
    .A(_02226_),
    .B(_02259_));
 sg13g2_xnor2_1 _13565_ (.Y(_02280_),
    .A(_02183_),
    .B(_02269_));
 sg13g2_o21ai_1 _13566_ (.B1(_02280_),
    .Y(_02291_),
    .A1(net1046),
    .A2(net1047));
 sg13g2_inv_1 _13567_ (.Y(_02302_),
    .A(_02097_));
 sg13g2_nor2_1 _13568_ (.A(net1045),
    .B(net1044),
    .Y(_02312_));
 sg13g2_a22oi_1 _13569_ (.Y(_02323_),
    .B1(_02312_),
    .B2(_02280_),
    .A2(_02291_),
    .A1(net711));
 sg13g2_buf_1 _13570_ (.A(_00250_),
    .X(_02334_));
 sg13g2_buf_1 _13571_ (.A(_02334_),
    .X(_02345_));
 sg13g2_a21o_1 _13572_ (.A2(_02323_),
    .A1(_02140_),
    .B1(net1043),
    .X(_02356_));
 sg13g2_buf_1 _13573_ (.A(_02119_),
    .X(_02366_));
 sg13g2_buf_1 _13574_ (.A(net1042),
    .X(_02377_));
 sg13g2_xnor2_1 _13575_ (.Y(_02388_),
    .A(_02087_),
    .B(_02280_));
 sg13g2_and2_1 _13576_ (.A(net1044),
    .B(_02280_),
    .X(_02399_));
 sg13g2_buf_2 _13577_ (.A(_00161_),
    .X(_02410_));
 sg13g2_buf_1 _13578_ (.A(_02248_),
    .X(_02421_));
 sg13g2_buf_1 _13579_ (.A(net1041),
    .X(_02432_));
 sg13g2_buf_1 _13580_ (.A(_02432_),
    .X(_02442_));
 sg13g2_xnor2_1 _13581_ (.Y(_02453_),
    .A(net374),
    .B(_02226_));
 sg13g2_buf_2 _13582_ (.A(net1185),
    .X(_02464_));
 sg13g2_buf_1 _13583_ (.A(net1040),
    .X(_02475_));
 sg13g2_nand2_1 _13584_ (.Y(_02486_),
    .A(net708),
    .B(_02269_));
 sg13g2_o21ai_1 _13585_ (.B1(_02486_),
    .Y(_02496_),
    .A1(_02410_),
    .A2(_02453_));
 sg13g2_a221oi_1 _13586_ (.B2(net1043),
    .C1(_02496_),
    .B1(_02399_),
    .A1(net710),
    .Y(_02507_),
    .A2(_02388_));
 sg13g2_inv_2 _13587_ (.Y(_02518_),
    .A(_02334_));
 sg13g2_a21oi_1 _13588_ (.A1(net710),
    .A2(_02518_),
    .Y(_02529_),
    .B1(_02399_));
 sg13g2_o21ai_1 _13589_ (.B1(_02388_),
    .Y(_02540_),
    .A1(net710),
    .A2(_02518_));
 sg13g2_nand2_1 _13590_ (.Y(_02550_),
    .A(_02529_),
    .B(_02540_));
 sg13g2_inv_1 _13591_ (.Y(_02561_),
    .A(net1041));
 sg13g2_buf_1 _13592_ (.A(_02561_),
    .X(_02572_));
 sg13g2_buf_1 _13593_ (.A(_02205_),
    .X(_02583_));
 sg13g2_buf_1 _13594_ (.A(net1039),
    .X(_02593_));
 sg13g2_inv_1 _13595_ (.Y(_02604_),
    .A(net707));
 sg13g2_buf_1 _13596_ (.A(_02604_),
    .X(_02615_));
 sg13g2_buf_1 _13597_ (.A(net374),
    .X(_02626_));
 sg13g2_buf_1 _13598_ (.A(net707),
    .X(_02636_));
 sg13g2_buf_1 _13599_ (.A(net372),
    .X(_02647_));
 sg13g2_buf_2 _13600_ (.A(_02194_),
    .X(_02658_));
 sg13g2_buf_1 _13601_ (.A(net1038),
    .X(_02669_));
 sg13g2_buf_2 _13602_ (.A(net706),
    .X(_02679_));
 sg13g2_a21oi_1 _13603_ (.A1(net174),
    .A2(net173),
    .Y(_02690_),
    .B1(net371));
 sg13g2_a21oi_1 _13604_ (.A1(net373),
    .A2(net175),
    .Y(_02701_),
    .B1(_02690_));
 sg13g2_a221oi_1 _13605_ (.B2(_02496_),
    .C1(_02701_),
    .B1(_02550_),
    .A1(_02356_),
    .Y(_02712_),
    .A2(_02507_));
 sg13g2_nand2b_1 _13606_ (.Y(_02722_),
    .B(_02701_),
    .A_N(_02496_));
 sg13g2_nand2b_1 _13607_ (.Y(_02733_),
    .B(net1191),
    .A_N(demo_step));
 sg13g2_and2_1 _13608_ (.A(net6),
    .B(_02733_),
    .X(_02744_));
 sg13g2_buf_2 _13609_ (.A(_02744_),
    .X(_02755_));
 sg13g2_buf_2 _13610_ (.A(_02755_),
    .X(_02765_));
 sg13g2_buf_2 _13611_ (.A(net172),
    .X(_02776_));
 sg13g2_buf_2 _13612_ (.A(net127),
    .X(_02787_));
 sg13g2_o21ai_1 _13613_ (.B1(net85),
    .Y(_02798_),
    .A1(_02550_),
    .A2(_02722_));
 sg13g2_buf_1 _13614_ (.A(_02755_),
    .X(_02809_));
 sg13g2_buf_1 _13615_ (.A(net171),
    .X(_02820_));
 sg13g2_buf_1 _13616_ (.A(\grid.cell_0_0.n ),
    .X(_02830_));
 sg13g2_xnor2_1 _13617_ (.Y(_02841_),
    .A(net1184),
    .B(net1186));
 sg13g2_xnor2_1 _13618_ (.Y(_02852_),
    .A(_02388_),
    .B(_02841_));
 sg13g2_buf_1 _13619_ (.A(\grid.cell_0_0.out ),
    .X(_02863_));
 sg13g2_buf_1 _13620_ (.A(net1183),
    .X(_02874_));
 sg13g2_a21oi_1 _13621_ (.A1(net126),
    .A2(_02852_),
    .Y(_02884_),
    .B1(net1037));
 sg13g2_or3_1 _13622_ (.A(_01870_),
    .B(_01989_),
    .C(_02021_),
    .X(_02895_));
 sg13g2_buf_2 _13623_ (.A(_02895_),
    .X(_02906_));
 sg13g2_nand2_1 _13624_ (.Y(_02917_),
    .A(net1197),
    .B(_02906_));
 sg13g2_buf_1 _13625_ (.A(_02917_),
    .X(_02928_));
 sg13g2_nor2_1 _13626_ (.A(_02884_),
    .B(_02928_),
    .Y(_02938_));
 sg13g2_o21ai_1 _13627_ (.B1(_02938_),
    .Y(_02949_),
    .A1(_02712_),
    .A2(_02798_));
 sg13g2_o21ai_1 _13628_ (.B1(_02949_),
    .Y(_00277_),
    .A1(net50),
    .A2(_02065_));
 sg13g2_buf_1 _13629_ (.A(net715),
    .X(_02970_));
 sg13g2_nand3_1 _13630_ (.B(net1050),
    .C(_01655_),
    .A(net1189),
    .Y(_02980_));
 sg13g2_and2_1 _13631_ (.A(_01557_),
    .B(_02980_),
    .X(_02991_));
 sg13g2_inv_2 _13632_ (.Y(_03002_),
    .A(_01601_));
 sg13g2_nor2b_1 _13633_ (.A(net1187),
    .B_N(_01666_),
    .Y(_03013_));
 sg13g2_buf_1 _13634_ (.A(_03013_),
    .X(_03023_));
 sg13g2_nand2_1 _13635_ (.Y(_03034_),
    .A(_03002_),
    .B(_03023_));
 sg13g2_inv_1 _13636_ (.Y(_03045_),
    .A(net1187));
 sg13g2_nand2_1 _13637_ (.Y(_03056_),
    .A(net1189),
    .B(_03045_));
 sg13g2_o21ai_1 _13638_ (.B1(_01525_),
    .Y(_03066_),
    .A1(_01752_),
    .A2(_03056_));
 sg13g2_nand3b_1 _13639_ (.B(net1049),
    .C(_01633_),
    .Y(_03077_),
    .A_N(net1188));
 sg13g2_buf_1 _13640_ (.A(_03077_),
    .X(_03088_));
 sg13g2_nand2b_1 _13641_ (.Y(_03099_),
    .B(net1190),
    .A_N(net1189));
 sg13g2_nor3_1 _13642_ (.A(net1048),
    .B(_03088_),
    .C(_03099_),
    .Y(_03109_));
 sg13g2_a21oi_1 _13643_ (.A1(net1048),
    .A2(_03066_),
    .Y(_03120_),
    .B1(_03109_));
 sg13g2_a21oi_1 _13644_ (.A1(_02991_),
    .A2(_03034_),
    .Y(_03131_),
    .B1(_03120_));
 sg13g2_mux2_1 _13645_ (.A0(net9),
    .A1(_03131_),
    .S(net376),
    .X(_03142_));
 sg13g2_buf_1 _13646_ (.A(_03142_),
    .X(_03153_));
 sg13g2_buf_1 _13647_ (.A(_03153_),
    .X(_03164_));
 sg13g2_buf_2 _13648_ (.A(\grid.cell_0_1.e ),
    .X(_03174_));
 sg13g2_buf_2 _13649_ (.A(\grid.cell_0_1.se ),
    .X(_03185_));
 sg13g2_xnor2_1 _13650_ (.Y(_03196_),
    .A(_03174_),
    .B(_03185_));
 sg13g2_buf_2 _13651_ (.A(_03196_),
    .X(_03207_));
 sg13g2_buf_1 _13652_ (.A(\grid.cell_0_1.ne ),
    .X(_03218_));
 sg13g2_buf_1 _13653_ (.A(_03218_),
    .X(_03229_));
 sg13g2_xnor2_1 _13654_ (.Y(_03240_),
    .A(_02194_),
    .B(net1036));
 sg13g2_xnor2_1 _13655_ (.Y(_03250_),
    .A(_03207_),
    .B(_03240_));
 sg13g2_xnor2_1 _13656_ (.Y(_03261_),
    .A(net1185),
    .B(_03250_));
 sg13g2_buf_1 _13657_ (.A(net1184),
    .X(_03272_));
 sg13g2_xor2_1 _13658_ (.B(_02076_),
    .A(net1183),
    .X(_03283_));
 sg13g2_xnor2_1 _13659_ (.Y(_03294_),
    .A(net1035),
    .B(_03283_));
 sg13g2_xnor2_1 _13660_ (.Y(_03304_),
    .A(_03261_),
    .B(_03294_));
 sg13g2_inv_1 _13661_ (.Y(_03315_),
    .A(net1036));
 sg13g2_buf_1 _13662_ (.A(_03174_),
    .X(_03326_));
 sg13g2_buf_1 _13663_ (.A(_03185_),
    .X(_03337_));
 sg13g2_nand2_1 _13664_ (.Y(_03347_),
    .A(net1034),
    .B(net1033));
 sg13g2_mux2_1 _13665_ (.A0(_03347_),
    .A1(_03207_),
    .S(net706),
    .X(_03358_));
 sg13g2_buf_1 _13666_ (.A(net1034),
    .X(_03369_));
 sg13g2_buf_1 _13667_ (.A(net1033),
    .X(_03380_));
 sg13g2_nand4_1 _13668_ (.B(net705),
    .C(net704),
    .A(net706),
    .Y(_03390_),
    .D(_03315_));
 sg13g2_o21ai_1 _13669_ (.B1(_03390_),
    .Y(_03401_),
    .A1(_03315_),
    .A2(_03358_));
 sg13g2_nor3_1 _13670_ (.A(net1047),
    .B(_02345_),
    .C(_03283_),
    .Y(_03412_));
 sg13g2_nand2_1 _13671_ (.Y(_03423_),
    .A(net371),
    .B(net704));
 sg13g2_buf_1 _13672_ (.A(_00216_),
    .X(_03433_));
 sg13g2_nand2b_1 _13673_ (.Y(_03444_),
    .B(_03229_),
    .A_N(net1182));
 sg13g2_o21ai_1 _13674_ (.B1(_02755_),
    .Y(_03455_),
    .A1(_03423_),
    .A2(_03444_));
 sg13g2_a221oi_1 _13675_ (.B2(_03412_),
    .C1(_03455_),
    .B1(_03261_),
    .A1(net708),
    .Y(_03466_),
    .A2(_03401_));
 sg13g2_o21ai_1 _13676_ (.B1(_03466_),
    .Y(_03477_),
    .A1(net710),
    .A2(_03304_));
 sg13g2_nor2_1 _13677_ (.A(net1183),
    .B(_02518_),
    .Y(_03487_));
 sg13g2_xnor2_1 _13678_ (.Y(_03498_),
    .A(net1045),
    .B(_03261_));
 sg13g2_a22oi_1 _13679_ (.Y(_03509_),
    .B1(_03261_),
    .B2(net1044),
    .A2(_02518_),
    .A1(net1037));
 sg13g2_o21ai_1 _13680_ (.B1(_03509_),
    .Y(_03519_),
    .A1(_03487_),
    .A2(_03498_));
 sg13g2_inv_2 _13681_ (.Y(_03530_),
    .A(net1034));
 sg13g2_buf_1 _13682_ (.A(net1036),
    .X(_03541_));
 sg13g2_nor3_1 _13683_ (.A(net706),
    .B(net704),
    .C(net703),
    .Y(_03552_));
 sg13g2_nand4_1 _13684_ (.B(net706),
    .C(net704),
    .A(net1040),
    .Y(_03563_),
    .D(net703));
 sg13g2_nand2b_1 _13685_ (.Y(_03573_),
    .B(_03563_),
    .A_N(_03552_));
 sg13g2_nand2_1 _13686_ (.Y(_03584_),
    .A(net1185),
    .B(net1034));
 sg13g2_o21ai_1 _13687_ (.B1(_03444_),
    .Y(_03595_),
    .A1(net703),
    .A2(_03584_));
 sg13g2_buf_1 _13688_ (.A(net1036),
    .X(_03606_));
 sg13g2_nor2_1 _13689_ (.A(net702),
    .B(net1182),
    .Y(_03617_));
 sg13g2_nor3_1 _13690_ (.A(net1033),
    .B(_03584_),
    .C(_03617_),
    .Y(_03628_));
 sg13g2_a21oi_1 _13691_ (.A1(net704),
    .A2(_03595_),
    .Y(_03638_),
    .B1(_03628_));
 sg13g2_nand2_1 _13692_ (.Y(_03649_),
    .A(_02679_),
    .B(_03638_));
 sg13g2_nand2_1 _13693_ (.Y(_03660_),
    .A(_03315_),
    .B(net1182));
 sg13g2_inv_1 _13694_ (.Y(_03671_),
    .A(_03185_));
 sg13g2_buf_1 _13695_ (.A(_03671_),
    .X(_03682_));
 sg13g2_nand2_1 _13696_ (.Y(_03692_),
    .A(net701),
    .B(_03444_));
 sg13g2_a21oi_1 _13697_ (.A1(_03660_),
    .A2(_03692_),
    .Y(_03703_),
    .B1(net1040));
 sg13g2_nand2_1 _13698_ (.Y(_03714_),
    .A(net702),
    .B(net1182));
 sg13g2_o21ai_1 _13699_ (.B1(net1033),
    .Y(_03724_),
    .A1(net702),
    .A2(net1182));
 sg13g2_a21oi_1 _13700_ (.A1(_03714_),
    .A2(_03724_),
    .Y(_03735_),
    .B1(_03584_));
 sg13g2_or3_1 _13701_ (.A(_02669_),
    .B(_03703_),
    .C(_03735_),
    .X(_03746_));
 sg13g2_buf_1 _13702_ (.A(net704),
    .X(_03756_));
 sg13g2_nor3_1 _13703_ (.A(net708),
    .B(net369),
    .C(_03660_),
    .Y(_03767_));
 sg13g2_a221oi_1 _13704_ (.B2(_03746_),
    .C1(_03767_),
    .B1(_03649_),
    .A1(_03530_),
    .Y(_03778_),
    .A2(_03573_));
 sg13g2_xnor2_1 _13705_ (.Y(_03789_),
    .A(_03519_),
    .B(_03778_));
 sg13g2_nand2_1 _13706_ (.Y(_03799_),
    .A(net6),
    .B(_02733_));
 sg13g2_buf_2 _13707_ (.A(_03799_),
    .X(_03810_));
 sg13g2_buf_2 _13708_ (.A(net368),
    .X(_03821_));
 sg13g2_buf_1 _13709_ (.A(net170),
    .X(_03831_));
 sg13g2_a21oi_1 _13710_ (.A1(net710),
    .A2(net125),
    .Y(_03842_),
    .B1(_02054_));
 sg13g2_o21ai_1 _13711_ (.B1(_03842_),
    .Y(_03853_),
    .A1(_03477_),
    .A2(_03789_));
 sg13g2_o21ai_1 _13712_ (.B1(_03853_),
    .Y(_03864_),
    .A1(_02906_),
    .A2(net49));
 sg13g2_nor2_1 _13713_ (.A(net370),
    .B(_03864_),
    .Y(_00278_));
 sg13g2_nand2b_1 _13714_ (.Y(_03884_),
    .B(net10),
    .A_N(net713));
 sg13g2_buf_1 _13715_ (.A(net1187),
    .X(_03895_));
 sg13g2_nor3_1 _13716_ (.A(net1051),
    .B(net1050),
    .C(net1032),
    .Y(_03906_));
 sg13g2_a21oi_1 _13717_ (.A1(net1051),
    .A2(_01731_),
    .Y(_03916_),
    .B1(_03906_));
 sg13g2_inv_1 _13718_ (.Y(_03927_),
    .A(net1190));
 sg13g2_nor2_1 _13719_ (.A(_03927_),
    .B(_01547_),
    .Y(_03938_));
 sg13g2_o21ai_1 _13720_ (.B1(_03938_),
    .Y(_03949_),
    .A1(_01752_),
    .A2(_03916_));
 sg13g2_nand2b_1 _13721_ (.Y(_03960_),
    .B(net1049),
    .A_N(_01568_));
 sg13g2_nand2_1 _13722_ (.Y(_03970_),
    .A(_01612_),
    .B(_03895_));
 sg13g2_nand2b_1 _13723_ (.Y(_03981_),
    .B(_03970_),
    .A_N(_03960_));
 sg13g2_nor4_1 _13724_ (.A(net1188),
    .B(_03895_),
    .C(_01525_),
    .D(_01752_),
    .Y(_03992_));
 sg13g2_nand2b_1 _13725_ (.Y(_04003_),
    .B(net1187),
    .A_N(net1049));
 sg13g2_a21oi_1 _13726_ (.A1(_03088_),
    .A2(_04003_),
    .Y(_04013_),
    .B1(_03099_));
 sg13g2_nor3_1 _13727_ (.A(_01536_),
    .B(_03992_),
    .C(_04013_),
    .Y(_04024_));
 sg13g2_a21oi_1 _13728_ (.A1(_02991_),
    .A2(_03981_),
    .Y(_04035_),
    .B1(_04024_));
 sg13g2_nand3_1 _13729_ (.B(_03949_),
    .C(_04035_),
    .A(net713),
    .Y(_04046_));
 sg13g2_and2_1 _13730_ (.A(_03884_),
    .B(_04046_),
    .X(_04056_));
 sg13g2_buf_2 _13731_ (.A(_04056_),
    .X(_04067_));
 sg13g2_buf_2 _13732_ (.A(_04067_),
    .X(_04077_));
 sg13g2_buf_1 _13733_ (.A(net35),
    .X(_04088_));
 sg13g2_buf_1 _13734_ (.A(net702),
    .X(_04099_));
 sg13g2_buf_1 _13735_ (.A(net367),
    .X(_04109_));
 sg13g2_buf_1 _13736_ (.A(_00033_),
    .X(_04120_));
 sg13g2_buf_2 _13737_ (.A(\grid.cell_0_2.e ),
    .X(_04131_));
 sg13g2_buf_2 _13738_ (.A(_04131_),
    .X(_04142_));
 sg13g2_inv_1 _13739_ (.Y(_04152_),
    .A(net1031));
 sg13g2_buf_2 _13740_ (.A(\grid.cell_0_2.ne ),
    .X(_04163_));
 sg13g2_buf_1 _13741_ (.A(_04163_),
    .X(_04174_));
 sg13g2_inv_1 _13742_ (.Y(_04185_),
    .A(net1030));
 sg13g2_buf_1 _13743_ (.A(\grid.cell_0_2.se ),
    .X(_04195_));
 sg13g2_buf_1 _13744_ (.A(_04195_),
    .X(_04206_));
 sg13g2_buf_1 _13745_ (.A(_04206_),
    .X(_04217_));
 sg13g2_nor2_1 _13746_ (.A(_02087_),
    .B(net699),
    .Y(_04228_));
 sg13g2_inv_2 _13747_ (.Y(_04236_),
    .A(net1029));
 sg13g2_nor2_1 _13748_ (.A(_04236_),
    .B(_04185_),
    .Y(_04244_));
 sg13g2_a221oi_1 _13749_ (.B2(_04228_),
    .C1(_04244_),
    .B1(_04185_),
    .A1(_02076_),
    .Y(_04254_),
    .A2(net700));
 sg13g2_buf_1 _13750_ (.A(net1030),
    .X(_04264_));
 sg13g2_nor2_1 _13751_ (.A(net699),
    .B(net698),
    .Y(_04274_));
 sg13g2_buf_1 _13752_ (.A(net1031),
    .X(_04283_));
 sg13g2_nand2_1 _13753_ (.Y(_04294_),
    .A(net1045),
    .B(net697));
 sg13g2_a22oi_1 _13754_ (.Y(_04303_),
    .B1(_04274_),
    .B2(_04294_),
    .A2(_04254_),
    .A1(net1181));
 sg13g2_nand2_1 _13755_ (.Y(_04313_),
    .A(_03606_),
    .B(net1031));
 sg13g2_nand2_1 _13756_ (.Y(_04322_),
    .A(net1045),
    .B(_04313_));
 sg13g2_nand3_1 _13757_ (.B(_04274_),
    .C(_04322_),
    .A(net1181),
    .Y(_04332_));
 sg13g2_o21ai_1 _13758_ (.B1(_04332_),
    .Y(_04341_),
    .A1(net169),
    .A2(_04303_));
 sg13g2_inv_2 _13759_ (.Y(_04352_),
    .A(net1186));
 sg13g2_buf_1 _13760_ (.A(_00252_),
    .X(_04363_));
 sg13g2_nand2_1 _13761_ (.Y(_04374_),
    .A(_04352_),
    .B(_04363_));
 sg13g2_xor2_1 _13762_ (.B(_04131_),
    .A(net1029),
    .X(_04385_));
 sg13g2_xnor2_1 _13763_ (.Y(_04396_),
    .A(_03229_),
    .B(_04163_));
 sg13g2_xnor2_1 _13764_ (.Y(_04407_),
    .A(_04385_),
    .B(_04396_));
 sg13g2_xnor2_1 _13765_ (.Y(_04418_),
    .A(_02076_),
    .B(_04407_));
 sg13g2_xnor2_1 _13766_ (.Y(_04429_),
    .A(net704),
    .B(_04418_));
 sg13g2_buf_1 _13767_ (.A(_00214_),
    .X(_04440_));
 sg13g2_nand2b_1 _13768_ (.Y(_04451_),
    .B(net1046),
    .A_N(_04363_));
 sg13g2_o21ai_1 _13769_ (.B1(_04451_),
    .Y(_04462_),
    .A1(_04440_),
    .A2(_04418_));
 sg13g2_a21oi_1 _13770_ (.A1(_04374_),
    .A2(_04429_),
    .Y(_04473_),
    .B1(_04462_));
 sg13g2_xor2_1 _13771_ (.B(_04473_),
    .A(_04341_),
    .X(_04484_));
 sg13g2_buf_2 _13772_ (.A(net699),
    .X(_04495_));
 sg13g2_xor2_1 _13773_ (.B(_04163_),
    .A(_04131_),
    .X(_04506_));
 sg13g2_nand2_1 _13774_ (.Y(_04516_),
    .A(net1031),
    .B(_04174_));
 sg13g2_nor2_1 _13775_ (.A(net699),
    .B(_04516_),
    .Y(_04526_));
 sg13g2_a21oi_1 _13776_ (.A1(net366),
    .A2(_04506_),
    .Y(_04536_),
    .B1(_04526_));
 sg13g2_buf_1 _13777_ (.A(net698),
    .X(_04545_));
 sg13g2_nand4_1 _13778_ (.B(net366),
    .C(net697),
    .A(_03315_),
    .Y(_04554_),
    .D(net365));
 sg13g2_o21ai_1 _13779_ (.B1(_04554_),
    .Y(_04563_),
    .A1(_03315_),
    .A2(_04536_));
 sg13g2_nor2b_1 _13780_ (.A(net1181),
    .B_N(net169),
    .Y(_04573_));
 sg13g2_xor2_1 _13781_ (.B(net704),
    .A(net1046),
    .X(_04583_));
 sg13g2_nor4_1 _13782_ (.A(_04440_),
    .B(_04363_),
    .C(_04418_),
    .D(_04583_),
    .Y(_04592_));
 sg13g2_a221oi_1 _13783_ (.B2(_04244_),
    .C1(_04592_),
    .B1(_04573_),
    .A1(net711),
    .Y(_04603_),
    .A2(_04563_));
 sg13g2_buf_1 _13784_ (.A(net368),
    .X(_04614_));
 sg13g2_buf_1 _13785_ (.A(net168),
    .X(_04624_));
 sg13g2_a21oi_1 _13786_ (.A1(_04484_),
    .A2(_04603_),
    .Y(_04634_),
    .B1(net124));
 sg13g2_buf_1 _13787_ (.A(net172),
    .X(_04642_));
 sg13g2_buf_1 _13788_ (.A(net123),
    .X(_04650_));
 sg13g2_xor2_1 _13789_ (.B(_04583_),
    .A(_02679_),
    .X(_04658_));
 sg13g2_xnor2_1 _13790_ (.Y(_04666_),
    .A(_04418_),
    .B(_04658_));
 sg13g2_buf_1 _13791_ (.A(net705),
    .X(_04674_));
 sg13g2_a21oi_1 _13792_ (.A1(net84),
    .A2(_04666_),
    .Y(_04682_),
    .B1(net364));
 sg13g2_or3_1 _13793_ (.A(_02928_),
    .B(_04634_),
    .C(_04682_),
    .X(_04691_));
 sg13g2_o21ai_1 _13794_ (.B1(_04691_),
    .Y(_00279_),
    .A1(_02065_),
    .A2(net27));
 sg13g2_buf_2 _13795_ (.A(\grid.cell_0_3.se ),
    .X(_04705_));
 sg13g2_inv_2 _13796_ (.Y(_04712_),
    .A(_04705_));
 sg13g2_buf_1 _13797_ (.A(_04712_),
    .X(_04721_));
 sg13g2_buf_1 _13798_ (.A(\grid.cell_0_3.e ),
    .X(_04729_));
 sg13g2_buf_1 _13799_ (.A(\grid.cell_0_3.ne ),
    .X(_04737_));
 sg13g2_xnor2_1 _13800_ (.Y(_04748_),
    .A(net1180),
    .B(_04737_));
 sg13g2_buf_1 _13801_ (.A(net1180),
    .X(_04758_));
 sg13g2_buf_1 _13802_ (.A(net1028),
    .X(_04768_));
 sg13g2_buf_2 _13803_ (.A(_04737_),
    .X(_04779_));
 sg13g2_buf_1 _13804_ (.A(net1027),
    .X(_04789_));
 sg13g2_buf_1 _13805_ (.A(net694),
    .X(_04800_));
 sg13g2_nand3_1 _13806_ (.B(net695),
    .C(net363),
    .A(net696),
    .Y(_04810_));
 sg13g2_o21ai_1 _13807_ (.B1(_04810_),
    .Y(_04820_),
    .A1(net696),
    .A2(_04748_));
 sg13g2_inv_2 _13808_ (.Y(_04830_),
    .A(net1180));
 sg13g2_inv_1 _13809_ (.Y(_04841_),
    .A(net1027));
 sg13g2_nor4_1 _13810_ (.A(net696),
    .B(_04830_),
    .C(_04841_),
    .D(net365),
    .Y(_04851_));
 sg13g2_a21oi_1 _13811_ (.A1(net365),
    .A2(_04820_),
    .Y(_04855_),
    .B1(_04851_));
 sg13g2_nor2_1 _13812_ (.A(net701),
    .B(_04855_),
    .Y(_04856_));
 sg13g2_buf_2 _13813_ (.A(_00065_),
    .X(_04857_));
 sg13g2_nor4_1 _13814_ (.A(_04857_),
    .B(net696),
    .C(_04841_),
    .D(_04185_),
    .Y(_04858_));
 sg13g2_buf_1 _13815_ (.A(_02755_),
    .X(_04859_));
 sg13g2_buf_1 _13816_ (.A(net167),
    .X(_04860_));
 sg13g2_xor2_1 _13817_ (.B(_04163_),
    .A(_04737_),
    .X(_04861_));
 sg13g2_xnor2_1 _13818_ (.Y(_04862_),
    .A(_04705_),
    .B(net1180));
 sg13g2_xor2_1 _13819_ (.B(_04862_),
    .A(_04861_),
    .X(_04863_));
 sg13g2_xnor2_1 _13820_ (.Y(_04864_),
    .A(net1029),
    .B(_04863_));
 sg13g2_xor2_1 _13821_ (.B(_03207_),
    .A(net367),
    .X(_04865_));
 sg13g2_xnor2_1 _13822_ (.Y(_04866_),
    .A(_04864_),
    .B(_04865_));
 sg13g2_a21oi_1 _13823_ (.A1(net122),
    .A2(_04866_),
    .Y(_04867_),
    .B1(net697));
 sg13g2_nor4_1 _13824_ (.A(_02928_),
    .B(_04856_),
    .C(_04858_),
    .D(_04867_),
    .Y(_04868_));
 sg13g2_xnor2_1 _13825_ (.Y(_04869_),
    .A(net701),
    .B(_04864_));
 sg13g2_buf_2 _13826_ (.A(_00032_),
    .X(_04870_));
 sg13g2_xnor2_1 _13827_ (.Y(_04871_),
    .A(net701),
    .B(_04863_));
 sg13g2_nor2_1 _13828_ (.A(_04870_),
    .B(_04871_),
    .Y(_04872_));
 sg13g2_nor2_1 _13829_ (.A(_00251_),
    .B(_04872_),
    .Y(_04873_));
 sg13g2_nand2_1 _13830_ (.Y(_04874_),
    .A(_04869_),
    .B(_04873_));
 sg13g2_inv_1 _13831_ (.Y(_04875_),
    .A(_00251_));
 sg13g2_o21ai_1 _13832_ (.B1(_04875_),
    .Y(_04876_),
    .A1(net364),
    .A2(_04869_));
 sg13g2_nand2_1 _13833_ (.Y(_04877_),
    .A(_04872_),
    .B(_04876_));
 sg13g2_o21ai_1 _13834_ (.B1(net364),
    .Y(_04878_),
    .A1(_04869_),
    .A2(_04873_));
 sg13g2_nand3_1 _13835_ (.B(_04877_),
    .C(_04878_),
    .A(_04874_),
    .Y(_04879_));
 sg13g2_a21o_1 _13836_ (.A2(_04869_),
    .A1(_04875_),
    .B1(net364),
    .X(_04880_));
 sg13g2_or2_1 _13837_ (.X(_04881_),
    .B(_04869_),
    .A(_04875_));
 sg13g2_a21oi_1 _13838_ (.A1(_04880_),
    .A2(_04881_),
    .Y(_04882_),
    .B1(_04872_));
 sg13g2_nand2_1 _13839_ (.Y(_04883_),
    .A(net369),
    .B(net695));
 sg13g2_buf_1 _13840_ (.A(_04705_),
    .X(_04884_));
 sg13g2_buf_1 _13841_ (.A(net1026),
    .X(_04885_));
 sg13g2_nor3_1 _13842_ (.A(net693),
    .B(net363),
    .C(net365),
    .Y(_04886_));
 sg13g2_nand2_1 _13843_ (.Y(_04887_),
    .A(_04800_),
    .B(net365));
 sg13g2_a22oi_1 _13844_ (.Y(_04888_),
    .B1(_04887_),
    .B2(net701),
    .A2(_04861_),
    .A1(net695));
 sg13g2_a21oi_1 _13845_ (.A1(net1026),
    .A2(net1028),
    .Y(_04889_),
    .B1(net701));
 sg13g2_or3_1 _13846_ (.A(_04800_),
    .B(_04545_),
    .C(_04889_),
    .X(_04890_));
 sg13g2_o21ai_1 _13847_ (.B1(_04890_),
    .Y(_04891_),
    .A1(net693),
    .A2(_04888_));
 sg13g2_a22oi_1 _13848_ (.Y(_04892_),
    .B1(_04891_),
    .B2(_04857_),
    .A2(_04886_),
    .A1(_04883_));
 sg13g2_mux2_1 _13849_ (.A0(_04879_),
    .A1(_04882_),
    .S(_04892_),
    .X(_04893_));
 sg13g2_inv_1 _13850_ (.Y(_04894_),
    .A(_01579_));
 sg13g2_a21oi_1 _13851_ (.A1(net1188),
    .A2(_01655_),
    .Y(_04895_),
    .B1(_03023_));
 sg13g2_nand2b_1 _13852_ (.Y(_04896_),
    .B(_01666_),
    .A_N(_01633_));
 sg13g2_nand2b_1 _13853_ (.Y(_04897_),
    .B(_01720_),
    .A_N(net1190));
 sg13g2_or2_1 _13854_ (.X(_04898_),
    .B(net1049),
    .A(_01720_));
 sg13g2_nand4_1 _13855_ (.B(_04896_),
    .C(_04897_),
    .A(_03002_),
    .Y(_04899_),
    .D(_04898_));
 sg13g2_o21ai_1 _13856_ (.B1(_04899_),
    .Y(_04900_),
    .A1(net1052),
    .A2(_04895_));
 sg13g2_a21oi_1 _13857_ (.A1(_01579_),
    .A2(_01655_),
    .Y(_04901_),
    .B1(_03023_));
 sg13g2_nor3_1 _13858_ (.A(net1050),
    .B(net1052),
    .C(_04901_),
    .Y(_04902_));
 sg13g2_a21oi_1 _13859_ (.A1(_04894_),
    .A2(_04900_),
    .Y(_04903_),
    .B1(_04902_));
 sg13g2_nor2_1 _13860_ (.A(_03099_),
    .B(_04895_),
    .Y(_04904_));
 sg13g2_nor2_1 _13861_ (.A(net1189),
    .B(_01752_),
    .Y(_04905_));
 sg13g2_and2_1 _13862_ (.A(_01622_),
    .B(net1190),
    .X(_04906_));
 sg13g2_buf_1 _13863_ (.A(_04906_),
    .X(_04907_));
 sg13g2_a22oi_1 _13864_ (.Y(_04908_),
    .B1(_04907_),
    .B2(_03045_),
    .A2(_04905_),
    .A1(_03927_));
 sg13g2_nor2_1 _13865_ (.A(net1050),
    .B(_04908_),
    .Y(_04909_));
 sg13g2_o21ai_1 _13866_ (.B1(net1048),
    .Y(_04910_),
    .A1(_04904_),
    .A2(_04909_));
 sg13g2_o21ai_1 _13867_ (.B1(_04910_),
    .Y(_04911_),
    .A1(net1048),
    .A2(_04903_));
 sg13g2_nor2b_1 _13868_ (.A(net713),
    .B_N(net11),
    .Y(_04912_));
 sg13g2_a21oi_1 _13869_ (.A1(net376),
    .A2(_04911_),
    .Y(_04913_),
    .B1(_04912_));
 sg13g2_buf_1 _13870_ (.A(_04913_),
    .X(_04914_));
 sg13g2_buf_1 _13871_ (.A(net368),
    .X(_04915_));
 sg13g2_nand3_1 _13872_ (.B(_02906_),
    .C(net166),
    .A(net697),
    .Y(_04916_));
 sg13g2_o21ai_1 _13873_ (.B1(_04916_),
    .Y(_04917_),
    .A1(_02906_),
    .A2(net48));
 sg13g2_and2_1 _13874_ (.A(net716),
    .B(_04917_),
    .X(_04918_));
 sg13g2_a21o_1 _13875_ (.A2(_04893_),
    .A1(_04868_),
    .B1(_04918_),
    .X(_00280_));
 sg13g2_a21oi_1 _13876_ (.A1(_04894_),
    .A2(_03023_),
    .Y(_04919_),
    .B1(_01655_));
 sg13g2_nand2_1 _13877_ (.Y(_04920_),
    .A(_03002_),
    .B(net712));
 sg13g2_nand3_1 _13878_ (.B(_04003_),
    .C(_04920_),
    .A(_01590_),
    .Y(_04921_));
 sg13g2_o21ai_1 _13879_ (.B1(_04921_),
    .Y(_04922_),
    .A1(net1050),
    .A2(_04919_));
 sg13g2_nand2_1 _13880_ (.Y(_04923_),
    .A(net1049),
    .B(_01536_));
 sg13g2_nor2_1 _13881_ (.A(net1032),
    .B(_04923_),
    .Y(_04924_));
 sg13g2_o21ai_1 _13882_ (.B1(net1050),
    .Y(_04925_),
    .A1(_01655_),
    .A2(_04924_));
 sg13g2_nor2_1 _13883_ (.A(net1188),
    .B(_03045_),
    .Y(_04926_));
 sg13g2_nand3_1 _13884_ (.B(net1048),
    .C(_04926_),
    .A(_01676_),
    .Y(_04927_));
 sg13g2_a21oi_1 _13885_ (.A1(_04925_),
    .A2(_04927_),
    .Y(_04928_),
    .B1(net1051));
 sg13g2_a21oi_1 _13886_ (.A1(_01547_),
    .A2(_04922_),
    .Y(_04929_),
    .B1(_04928_));
 sg13g2_nor2b_1 _13887_ (.A(_01536_),
    .B_N(net712),
    .Y(_04930_));
 sg13g2_a22oi_1 _13888_ (.Y(_04931_),
    .B1(_04930_),
    .B2(_03045_),
    .A2(_04905_),
    .A1(_01536_));
 sg13g2_nor2_1 _13889_ (.A(net1050),
    .B(_04931_),
    .Y(_04932_));
 sg13g2_inv_1 _13890_ (.Y(_04933_),
    .A(_01752_));
 sg13g2_a21oi_1 _13891_ (.A1(_01536_),
    .A2(_04933_),
    .Y(_04934_),
    .B1(_04930_));
 sg13g2_nor3_1 _13892_ (.A(net1051),
    .B(net1032),
    .C(_04934_),
    .Y(_04935_));
 sg13g2_nor3_1 _13893_ (.A(net712),
    .B(net1048),
    .C(_03970_),
    .Y(_04936_));
 sg13g2_nor4_1 _13894_ (.A(net1052),
    .B(_04932_),
    .C(_04935_),
    .D(_04936_),
    .Y(_04937_));
 sg13g2_a21oi_1 _13895_ (.A1(net1052),
    .A2(_04929_),
    .Y(_04938_),
    .B1(_04937_));
 sg13g2_nor2b_1 _13896_ (.A(net376),
    .B_N(net12),
    .Y(_04939_));
 sg13g2_a21oi_1 _13897_ (.A1(net376),
    .A2(_04938_),
    .Y(_04940_),
    .B1(_04939_));
 sg13g2_buf_2 _13898_ (.A(_04940_),
    .X(_04941_));
 sg13g2_buf_2 _13899_ (.A(net47),
    .X(_04942_));
 sg13g2_buf_2 _13900_ (.A(\grid.cell_0_4.se ),
    .X(_04943_));
 sg13g2_buf_1 _13901_ (.A(_04943_),
    .X(_04944_));
 sg13g2_buf_1 _13902_ (.A(net1025),
    .X(_04945_));
 sg13g2_buf_2 _13903_ (.A(_00097_),
    .X(_04946_));
 sg13g2_buf_2 _13904_ (.A(\grid.cell_0_4.ne ),
    .X(_04947_));
 sg13g2_buf_1 _13905_ (.A(_04947_),
    .X(_04948_));
 sg13g2_nand2_2 _13906_ (.Y(_04949_),
    .A(net1024),
    .B(_04779_));
 sg13g2_buf_1 _13907_ (.A(\grid.cell_0_4.e ),
    .X(_04950_));
 sg13g2_buf_1 _13908_ (.A(net1179),
    .X(_04951_));
 sg13g2_xor2_1 _13909_ (.B(_04737_),
    .A(_04947_),
    .X(_04952_));
 sg13g2_nand2_1 _13910_ (.Y(_04953_),
    .A(net1023),
    .B(_04952_));
 sg13g2_o21ai_1 _13911_ (.B1(_04953_),
    .Y(_04954_),
    .A1(net1023),
    .A2(_04949_));
 sg13g2_nand2_1 _13912_ (.Y(_04955_),
    .A(net366),
    .B(_04954_));
 sg13g2_o21ai_1 _13913_ (.B1(_04955_),
    .Y(_04956_),
    .A1(_04946_),
    .A2(_04949_));
 sg13g2_inv_1 _13914_ (.Y(_04957_),
    .A(_04943_));
 sg13g2_buf_1 _13915_ (.A(_04957_),
    .X(_04958_));
 sg13g2_nand2_1 _13916_ (.Y(_04959_),
    .A(net691),
    .B(net1023));
 sg13g2_nor2_1 _13917_ (.A(_04949_),
    .B(_04959_),
    .Y(_04960_));
 sg13g2_a22oi_1 _13918_ (.Y(_04961_),
    .B1(_04960_),
    .B2(net366),
    .A2(_04956_),
    .A1(net692));
 sg13g2_buf_1 _13919_ (.A(_00062_),
    .X(_04962_));
 sg13g2_xnor2_1 _13920_ (.Y(_04963_),
    .A(_04943_),
    .B(net1179));
 sg13g2_xor2_1 _13921_ (.B(_04963_),
    .A(_04952_),
    .X(_04964_));
 sg13g2_xnor2_1 _13922_ (.Y(_04965_),
    .A(_04195_),
    .B(_04131_));
 sg13g2_xnor2_1 _13923_ (.Y(_04966_),
    .A(_04712_),
    .B(_04965_));
 sg13g2_xnor2_1 _13924_ (.Y(_04967_),
    .A(_04964_),
    .B(_04966_));
 sg13g2_or2_1 _13925_ (.X(_04968_),
    .B(_04967_),
    .A(_04962_));
 sg13g2_nor2_1 _13926_ (.A(_04712_),
    .B(net700),
    .Y(_04969_));
 sg13g2_buf_2 _13927_ (.A(_00064_),
    .X(_04970_));
 sg13g2_o21ai_1 _13928_ (.B1(_04970_),
    .Y(_04971_),
    .A1(net1026),
    .A2(net700));
 sg13g2_xnor2_1 _13929_ (.Y(_04972_),
    .A(_04217_),
    .B(_04964_));
 sg13g2_mux2_1 _13930_ (.A0(_04969_),
    .A1(_04971_),
    .S(_04972_),
    .X(_04973_));
 sg13g2_a22oi_1 _13931_ (.Y(_04974_),
    .B1(_04949_),
    .B2(_04236_),
    .A2(_04952_),
    .A1(net1179));
 sg13g2_nand2_1 _13932_ (.Y(_04975_),
    .A(_04943_),
    .B(_04950_));
 sg13g2_or2_1 _13933_ (.X(_04976_),
    .B(net1027),
    .A(net1024));
 sg13g2_buf_1 _13934_ (.A(_04976_),
    .X(_04977_));
 sg13g2_a21o_1 _13935_ (.A2(_04975_),
    .A1(net1029),
    .B1(_04977_),
    .X(_04978_));
 sg13g2_o21ai_1 _13936_ (.B1(_04978_),
    .Y(_04979_),
    .A1(net1025),
    .A2(_04974_));
 sg13g2_a21oi_1 _13937_ (.A1(net1023),
    .A2(net699),
    .Y(_04980_),
    .B1(_04977_));
 sg13g2_a22oi_1 _13938_ (.Y(_04981_),
    .B1(_04980_),
    .B2(net691),
    .A2(_04979_),
    .A1(_04946_));
 sg13g2_xor2_1 _13939_ (.B(_04981_),
    .A(_04973_),
    .X(_04982_));
 sg13g2_nor3_1 _13940_ (.A(_04973_),
    .B(_04981_),
    .C(_04968_),
    .Y(_04983_));
 sg13g2_a21o_1 _13941_ (.A2(_04982_),
    .A1(_04968_),
    .B1(_04983_),
    .X(_04984_));
 sg13g2_a21oi_1 _13942_ (.A1(_04961_),
    .A2(_04984_),
    .Y(_04985_),
    .B1(net124));
 sg13g2_xnor2_1 _13943_ (.Y(_04986_),
    .A(_04545_),
    .B(_04967_));
 sg13g2_a21oi_1 _13944_ (.A1(net84),
    .A2(_04986_),
    .Y(_04987_),
    .B1(net695));
 sg13g2_or3_1 _13945_ (.A(_02928_),
    .B(_04985_),
    .C(_04987_),
    .X(_04988_));
 sg13g2_o21ai_1 _13946_ (.B1(_04988_),
    .Y(_00281_),
    .A1(_02065_),
    .A2(net34));
 sg13g2_a21oi_1 _13947_ (.A1(net1032),
    .A2(_01547_),
    .Y(_04989_),
    .B1(_03960_));
 sg13g2_nand2b_1 _13948_ (.Y(_04990_),
    .B(_01568_),
    .A_N(net1049));
 sg13g2_a21oi_1 _13949_ (.A1(_01633_),
    .A2(_01547_),
    .Y(_04991_),
    .B1(_04990_));
 sg13g2_or2_1 _13950_ (.X(_04992_),
    .B(_04991_),
    .A(_04989_));
 sg13g2_nor3_1 _13951_ (.A(net1032),
    .B(net712),
    .C(_01547_),
    .Y(_04993_));
 sg13g2_a21o_1 _13952_ (.A2(_04930_),
    .A1(net1032),
    .B1(_04993_),
    .X(_04994_));
 sg13g2_nor3_1 _13953_ (.A(net1051),
    .B(net1032),
    .C(_04923_),
    .Y(_04995_));
 sg13g2_a221oi_1 _13954_ (.B2(net1051),
    .C1(_04995_),
    .B1(_04994_),
    .A1(_03002_),
    .Y(_04996_),
    .A2(_04992_));
 sg13g2_nor2_1 _13955_ (.A(net1051),
    .B(_03088_),
    .Y(_04997_));
 sg13g2_nor2_1 _13956_ (.A(net1052),
    .B(_04997_),
    .Y(_04998_));
 sg13g2_a21oi_1 _13957_ (.A1(net1052),
    .A2(_04996_),
    .Y(_04999_),
    .B1(_04998_));
 sg13g2_nor2b_1 _13958_ (.A(net376),
    .B_N(net13),
    .Y(_05000_));
 sg13g2_a21oi_1 _13959_ (.A1(net376),
    .A2(_04999_),
    .Y(_05001_),
    .B1(_05000_));
 sg13g2_buf_2 _13960_ (.A(_05001_),
    .X(_05002_));
 sg13g2_buf_1 _13961_ (.A(_05002_),
    .X(_05003_));
 sg13g2_buf_1 _13962_ (.A(\grid.cell_0_5.se ),
    .X(_05004_));
 sg13g2_buf_2 _13963_ (.A(_05004_),
    .X(_05005_));
 sg13g2_buf_1 _13964_ (.A(net1022),
    .X(_05006_));
 sg13g2_buf_1 _13965_ (.A(net690),
    .X(_05007_));
 sg13g2_buf_1 _13966_ (.A(_00129_),
    .X(_05008_));
 sg13g2_buf_1 _13967_ (.A(net1178),
    .X(_05009_));
 sg13g2_buf_1 _13968_ (.A(net1021),
    .X(_05010_));
 sg13g2_buf_1 _13969_ (.A(\grid.cell_0_5.ne ),
    .X(_05011_));
 sg13g2_buf_1 _13970_ (.A(_05011_),
    .X(_05012_));
 sg13g2_buf_1 _13971_ (.A(net1020),
    .X(_05013_));
 sg13g2_buf_1 _13972_ (.A(_04948_),
    .X(_05014_));
 sg13g2_nand2_1 _13973_ (.Y(_05015_),
    .A(net688),
    .B(net687));
 sg13g2_buf_2 _13974_ (.A(\grid.cell_0_5.e ),
    .X(_05016_));
 sg13g2_buf_1 _13975_ (.A(_05016_),
    .X(_05017_));
 sg13g2_buf_1 _13976_ (.A(net1019),
    .X(_05018_));
 sg13g2_xor2_1 _13977_ (.B(_04947_),
    .A(_05011_),
    .X(_05019_));
 sg13g2_nand2_1 _13978_ (.Y(_05020_),
    .A(net1019),
    .B(_05019_));
 sg13g2_o21ai_1 _13979_ (.B1(_05020_),
    .Y(_05021_),
    .A1(net686),
    .A2(_05015_));
 sg13g2_nand2_1 _13980_ (.Y(_05022_),
    .A(net693),
    .B(_05021_));
 sg13g2_o21ai_1 _13981_ (.B1(_05022_),
    .Y(_05023_),
    .A1(net689),
    .A2(_05015_));
 sg13g2_buf_1 _13982_ (.A(_00096_),
    .X(_05024_));
 sg13g2_inv_1 _13983_ (.Y(_05025_),
    .A(_05024_));
 sg13g2_xnor2_1 _13984_ (.Y(_05026_),
    .A(_05004_),
    .B(_05016_));
 sg13g2_xor2_1 _13985_ (.B(_05026_),
    .A(_05019_),
    .X(_05027_));
 sg13g2_xnor2_1 _13986_ (.Y(_05028_),
    .A(net1026),
    .B(_05027_));
 sg13g2_and2_1 _13987_ (.A(_05025_),
    .B(_05028_),
    .X(_05029_));
 sg13g2_buf_2 _13988_ (.A(_00094_),
    .X(_05030_));
 sg13g2_xor2_1 _13989_ (.B(net695),
    .A(net692),
    .X(_05031_));
 sg13g2_nor2_1 _13990_ (.A(_05030_),
    .B(_05031_),
    .Y(_05032_));
 sg13g2_nand2_1 _13991_ (.Y(_05033_),
    .A(net686),
    .B(net693));
 sg13g2_nor3_1 _13992_ (.A(net362),
    .B(_05015_),
    .C(_05033_),
    .Y(_05034_));
 sg13g2_a221oi_1 _13993_ (.B2(_05032_),
    .C1(_05034_),
    .B1(_05029_),
    .A1(net362),
    .Y(_05035_),
    .A2(_05023_));
 sg13g2_xnor2_1 _13994_ (.Y(_05036_),
    .A(net691),
    .B(_05028_));
 sg13g2_nand2_1 _13995_ (.Y(_05037_),
    .A(_05030_),
    .B(_04830_));
 sg13g2_nor2_1 _13996_ (.A(_05030_),
    .B(_04830_),
    .Y(_05038_));
 sg13g2_a221oi_1 _13997_ (.B2(_05037_),
    .C1(_05038_),
    .B1(_05036_),
    .A1(_05025_),
    .Y(_05039_),
    .A2(_05028_));
 sg13g2_a22oi_1 _13998_ (.Y(_05040_),
    .B1(_05015_),
    .B2(net696),
    .A2(_05019_),
    .A1(_05017_));
 sg13g2_nand2_1 _13999_ (.Y(_05041_),
    .A(net1022),
    .B(net1019));
 sg13g2_or2_1 _14000_ (.X(_05042_),
    .B(net1024),
    .A(_05013_));
 sg13g2_buf_1 _14001_ (.A(_05042_),
    .X(_05043_));
 sg13g2_a21o_1 _14002_ (.A2(_05041_),
    .A1(net1026),
    .B1(_05043_),
    .X(_05044_));
 sg13g2_o21ai_1 _14003_ (.B1(_05044_),
    .Y(_05045_),
    .A1(net690),
    .A2(_05040_));
 sg13g2_nor2_1 _14004_ (.A(net362),
    .B(_05043_),
    .Y(_05046_));
 sg13g2_a22oi_1 _14005_ (.Y(_05047_),
    .B1(_05046_),
    .B2(_05033_),
    .A2(_05045_),
    .A1(net689));
 sg13g2_xnor2_1 _14006_ (.Y(_05048_),
    .A(_05039_),
    .B(_05047_));
 sg13g2_a21oi_1 _14007_ (.A1(_05035_),
    .A2(_05048_),
    .Y(_05049_),
    .B1(net124));
 sg13g2_xnor2_1 _14008_ (.Y(_05050_),
    .A(_04748_),
    .B(_05036_));
 sg13g2_buf_1 _14009_ (.A(_04951_),
    .X(_05051_));
 sg13g2_a21oi_1 _14010_ (.A1(net84),
    .A2(_05050_),
    .Y(_05052_),
    .B1(net685));
 sg13g2_or3_1 _14011_ (.A(_02928_),
    .B(_05049_),
    .C(_05052_),
    .X(_05053_));
 sg13g2_o21ai_1 _14012_ (.B1(_05053_),
    .Y(_00282_),
    .A1(_02065_),
    .A2(net46));
 sg13g2_inv_1 _14013_ (.Y(_05054_),
    .A(_02410_));
 sg13g2_and2_1 _14014_ (.A(net1020),
    .B(_02205_),
    .X(_05055_));
 sg13g2_buf_1 _14015_ (.A(_05055_),
    .X(_05056_));
 sg13g2_buf_1 _14016_ (.A(_05056_),
    .X(_05057_));
 sg13g2_xor2_1 _14017_ (.B(net1039),
    .A(net1020),
    .X(_05058_));
 sg13g2_buf_1 _14018_ (.A(_02237_),
    .X(_05059_));
 sg13g2_buf_1 _14019_ (.A(net1018),
    .X(_05060_));
 sg13g2_mux2_1 _14020_ (.A0(net165),
    .A1(_05058_),
    .S(net684),
    .X(_05061_));
 sg13g2_a22oi_1 _14021_ (.Y(_05062_),
    .B1(_05061_),
    .B2(net692),
    .A2(net165),
    .A1(_05054_));
 sg13g2_nor2_1 _14022_ (.A(net373),
    .B(_05062_),
    .Y(_05063_));
 sg13g2_buf_1 _14023_ (.A(net687),
    .X(_05064_));
 sg13g2_xnor2_1 _14024_ (.Y(_05065_),
    .A(_05011_),
    .B(_02205_));
 sg13g2_xnor2_1 _14025_ (.Y(_05066_),
    .A(net1041),
    .B(_05065_));
 sg13g2_xnor2_1 _14026_ (.Y(_05067_),
    .A(net1018),
    .B(_05066_));
 sg13g2_xnor2_1 _14027_ (.Y(_05068_),
    .A(net1022),
    .B(_04963_));
 sg13g2_xnor2_1 _14028_ (.Y(_05069_),
    .A(_05067_),
    .B(_05068_));
 sg13g2_xor2_1 _14029_ (.B(_05069_),
    .A(net361),
    .X(_05070_));
 sg13g2_buf_1 _14030_ (.A(_05018_),
    .X(_05071_));
 sg13g2_a21oi_1 _14031_ (.A1(net123),
    .A2(_05070_),
    .Y(_05072_),
    .B1(net360));
 sg13g2_buf_1 _14032_ (.A(net684),
    .X(_05073_));
 sg13g2_buf_2 _14033_ (.A(net688),
    .X(_05074_));
 sg13g2_buf_1 _14034_ (.A(net358),
    .X(_05075_));
 sg13g2_nand4_1 _14035_ (.B(net692),
    .C(_05075_),
    .A(net359),
    .Y(_05076_),
    .D(net173));
 sg13g2_o21ai_1 _14036_ (.B1(_02906_),
    .Y(_05077_),
    .A1(net174),
    .A2(_05076_));
 sg13g2_nor3_1 _14037_ (.A(_05063_),
    .B(_05072_),
    .C(_05077_),
    .Y(_05078_));
 sg13g2_or2_1 _14038_ (.X(_05079_),
    .B(_02205_),
    .A(net1020));
 sg13g2_buf_1 _14039_ (.A(_05079_),
    .X(_05080_));
 sg13g2_nand2b_1 _14040_ (.Y(_05081_),
    .B(_02561_),
    .A_N(_05080_));
 sg13g2_a21oi_1 _14041_ (.A1(net1041),
    .A2(_05080_),
    .Y(_05082_),
    .B1(_05056_));
 sg13g2_nand2_1 _14042_ (.Y(_05083_),
    .A(_02410_),
    .B(_05082_));
 sg13g2_a21oi_1 _14043_ (.A1(_05081_),
    .A2(_05083_),
    .Y(_05084_),
    .B1(net1025));
 sg13g2_nand2_1 _14044_ (.Y(_05085_),
    .A(net709),
    .B(net165));
 sg13g2_nor2_1 _14045_ (.A(_02410_),
    .B(_05085_),
    .Y(_05086_));
 sg13g2_nor3_1 _14046_ (.A(_05054_),
    .B(_02561_),
    .C(net165),
    .Y(_05087_));
 sg13g2_a21oi_1 _14047_ (.A1(_05054_),
    .A2(net165),
    .Y(_05088_),
    .B1(_05087_));
 sg13g2_xor2_1 _14048_ (.B(net1041),
    .A(_02410_),
    .X(_05089_));
 sg13g2_nand2_1 _14049_ (.Y(_05090_),
    .A(_05080_),
    .B(_05089_));
 sg13g2_nand2_1 _14050_ (.Y(_05091_),
    .A(_05059_),
    .B(net1025));
 sg13g2_a21oi_1 _14051_ (.A1(_05088_),
    .A2(_05090_),
    .Y(_05092_),
    .B1(_05091_));
 sg13g2_nand3_1 _14052_ (.B(net1025),
    .C(net165),
    .A(net709),
    .Y(_05093_));
 sg13g2_a21oi_1 _14053_ (.A1(_05081_),
    .A2(_05093_),
    .Y(_05094_),
    .B1(net684));
 sg13g2_nor4_2 _14054_ (.A(_05084_),
    .B(_05086_),
    .C(_05092_),
    .Y(_05095_),
    .D(_05094_));
 sg13g2_buf_1 _14055_ (.A(_00126_),
    .X(_05096_));
 sg13g2_nor2b_1 _14056_ (.A(_05096_),
    .B_N(_05069_),
    .Y(_05097_));
 sg13g2_nor2_1 _14057_ (.A(_05095_),
    .B(_05097_),
    .Y(_05098_));
 sg13g2_xor2_1 _14058_ (.B(_05097_),
    .A(_05095_),
    .X(_05099_));
 sg13g2_xnor2_1 _14059_ (.Y(_05100_),
    .A(net691),
    .B(_05067_));
 sg13g2_inv_2 _14060_ (.Y(_05101_),
    .A(net1179));
 sg13g2_buf_1 _14061_ (.A(_00128_),
    .X(_05102_));
 sg13g2_o21ai_1 _14062_ (.B1(net1177),
    .Y(_05103_),
    .A1(net362),
    .A2(_05101_));
 sg13g2_inv_1 _14063_ (.Y(_05104_),
    .A(net1022));
 sg13g2_buf_1 _14064_ (.A(_05104_),
    .X(_05105_));
 sg13g2_o21ai_1 _14065_ (.B1(_05100_),
    .Y(_05106_),
    .A1(net357),
    .A2(_05101_));
 sg13g2_o21ai_1 _14066_ (.B1(_05106_),
    .Y(_05107_),
    .A1(_05100_),
    .A2(_05103_));
 sg13g2_mux2_1 _14067_ (.A0(_05098_),
    .A1(_05099_),
    .S(_05107_),
    .X(_05108_));
 sg13g2_a22oi_1 _14068_ (.Y(_05109_),
    .B1(_03023_),
    .B2(_01514_),
    .A2(_01827_),
    .A1(net1187));
 sg13g2_and2_1 _14069_ (.A(net1189),
    .B(_01655_),
    .X(_05110_));
 sg13g2_nand3_1 _14070_ (.B(_01514_),
    .C(_05110_),
    .A(_03002_),
    .Y(_05111_));
 sg13g2_o21ai_1 _14071_ (.B1(_05111_),
    .Y(_05112_),
    .A1(net1189),
    .A2(_05109_));
 sg13g2_a21oi_1 _14072_ (.A1(_03960_),
    .A2(_04990_),
    .Y(_05113_),
    .B1(net1187));
 sg13g2_a22oi_1 _14073_ (.Y(_05114_),
    .B1(_05113_),
    .B2(net1188),
    .A2(_04926_),
    .A1(net712));
 sg13g2_nor3_1 _14074_ (.A(_01536_),
    .B(_00019_),
    .C(_05114_),
    .Y(_05115_));
 sg13g2_a21o_1 _14075_ (.A2(_05112_),
    .A1(net1048),
    .B1(_05115_),
    .X(_05116_));
 sg13g2_mux2_1 _14076_ (.A0(net14),
    .A1(_05116_),
    .S(net713),
    .X(_05117_));
 sg13g2_buf_1 _14077_ (.A(_05117_),
    .X(_05118_));
 sg13g2_buf_1 _14078_ (.A(_05118_),
    .X(_05119_));
 sg13g2_inv_1 _14079_ (.Y(_05120_),
    .A(_05016_));
 sg13g2_buf_1 _14080_ (.A(_05120_),
    .X(_05121_));
 sg13g2_nor3_1 _14081_ (.A(_05121_),
    .B(_02054_),
    .C(net85),
    .Y(_05122_));
 sg13g2_a221oi_1 _14082_ (.B2(_02054_),
    .C1(_05122_),
    .B1(net45),
    .A1(_05078_),
    .Y(_05123_),
    .A2(_05108_));
 sg13g2_nor2_1 _14083_ (.A(net370),
    .B(_05123_),
    .Y(_00283_));
 sg13g2_buf_1 _14084_ (.A(net714),
    .X(_05124_));
 sg13g2_or2_1 _14085_ (.X(_05125_),
    .B(_00019_),
    .A(_00017_));
 sg13g2_nor4_1 _14086_ (.A(_03002_),
    .B(net712),
    .C(_03056_),
    .D(_05125_),
    .Y(_05126_));
 sg13g2_nor2b_1 _14087_ (.A(net713),
    .B_N(net15),
    .Y(_05127_));
 sg13g2_a21oi_1 _14088_ (.A1(net713),
    .A2(_05126_),
    .Y(_05128_),
    .B1(_05127_));
 sg13g2_buf_1 _14089_ (.A(_05128_),
    .X(_05129_));
 sg13g2_buf_2 _14090_ (.A(net368),
    .X(_05130_));
 sg13g2_buf_2 _14091_ (.A(net163),
    .X(_05131_));
 sg13g2_nand3_1 _14092_ (.B(_02906_),
    .C(net120),
    .A(net359),
    .Y(_05132_));
 sg13g2_o21ai_1 _14093_ (.B1(_05132_),
    .Y(_05133_),
    .A1(_02906_),
    .A2(net121));
 sg13g2_nand2_1 _14094_ (.Y(_05134_),
    .A(net174),
    .B(net358));
 sg13g2_nor3_1 _14095_ (.A(net689),
    .B(net175),
    .C(_05134_),
    .Y(_05135_));
 sg13g2_buf_1 _14096_ (.A(net172),
    .X(_05136_));
 sg13g2_xnor2_1 _14097_ (.Y(_05137_),
    .A(net1183),
    .B(net1185));
 sg13g2_xor2_1 _14098_ (.B(_05137_),
    .A(_05026_),
    .X(_05138_));
 sg13g2_xnor2_1 _14099_ (.Y(_05139_),
    .A(_05066_),
    .B(_05138_));
 sg13g2_xnor2_1 _14100_ (.Y(_05140_),
    .A(_03272_),
    .B(_05139_));
 sg13g2_a21oi_1 _14101_ (.A1(net119),
    .A2(_05140_),
    .Y(_05141_),
    .B1(net359));
 sg13g2_nor2_1 _14102_ (.A(net360),
    .B(_05134_),
    .Y(_05142_));
 sg13g2_xnor2_1 _14103_ (.Y(_05143_),
    .A(net374),
    .B(_05074_));
 sg13g2_nor2_1 _14104_ (.A(net683),
    .B(_05143_),
    .Y(_05144_));
 sg13g2_o21ai_1 _14105_ (.B1(_02647_),
    .Y(_05145_),
    .A1(_05142_),
    .A2(_05144_));
 sg13g2_nand4_1 _14106_ (.B(net174),
    .C(_05075_),
    .A(net360),
    .Y(_05146_),
    .D(_02615_));
 sg13g2_a21oi_1 _14107_ (.A1(_05145_),
    .A2(_05146_),
    .Y(_05147_),
    .B1(_02183_));
 sg13g2_nor4_1 _14108_ (.A(_02928_),
    .B(_05135_),
    .C(_05141_),
    .D(_05147_),
    .Y(_05148_));
 sg13g2_nor2_1 _14109_ (.A(_02345_),
    .B(_05139_),
    .Y(_05149_));
 sg13g2_inv_1 _14110_ (.Y(_05150_),
    .A(net1177));
 sg13g2_xnor2_1 _14111_ (.Y(_05151_),
    .A(net1185),
    .B(net1019));
 sg13g2_xnor2_1 _14112_ (.Y(_05152_),
    .A(_05066_),
    .B(_05151_));
 sg13g2_xnor2_1 _14113_ (.Y(_05153_),
    .A(net357),
    .B(_05152_));
 sg13g2_a22oi_1 _14114_ (.Y(_05154_),
    .B1(_05153_),
    .B2(_02874_),
    .A2(_05152_),
    .A1(_05150_));
 sg13g2_nor3_1 _14115_ (.A(net1040),
    .B(net374),
    .C(_05080_),
    .Y(_05155_));
 sg13g2_nand3_1 _14116_ (.B(net709),
    .C(_05057_),
    .A(net1040),
    .Y(_05156_));
 sg13g2_a21oi_1 _14117_ (.A1(_05081_),
    .A2(_05156_),
    .Y(_05157_),
    .B1(net686));
 sg13g2_nor2_1 _14118_ (.A(_05155_),
    .B(_05157_),
    .Y(_05158_));
 sg13g2_nand4_1 _14119_ (.B(net1019),
    .C(_02561_),
    .A(net1040),
    .Y(_05159_),
    .D(_05080_));
 sg13g2_o21ai_1 _14120_ (.B1(_05159_),
    .Y(_05160_),
    .A1(net1040),
    .A2(_05080_));
 sg13g2_nand2_1 _14121_ (.Y(_05161_),
    .A(net1185),
    .B(_05017_));
 sg13g2_mux2_1 _14122_ (.A0(net1185),
    .A1(_05161_),
    .S(net709),
    .X(_05162_));
 sg13g2_nor2_1 _14123_ (.A(_05057_),
    .B(_05162_),
    .Y(_05163_));
 sg13g2_o21ai_1 _14124_ (.B1(_05010_),
    .Y(_05164_),
    .A1(_05160_),
    .A2(_05163_));
 sg13g2_o21ai_1 _14125_ (.B1(_05085_),
    .Y(_05165_),
    .A1(_05082_),
    .A2(_05161_));
 sg13g2_nand2b_1 _14126_ (.Y(_05166_),
    .B(_05165_),
    .A_N(net1021));
 sg13g2_nand3_1 _14127_ (.B(_05164_),
    .C(_05166_),
    .A(_05158_),
    .Y(_05167_));
 sg13g2_xnor2_1 _14128_ (.Y(_05168_),
    .A(_05154_),
    .B(_05167_));
 sg13g2_nand3_1 _14129_ (.B(_05167_),
    .C(_05149_),
    .A(_05154_),
    .Y(_05169_));
 sg13g2_o21ai_1 _14130_ (.B1(_05169_),
    .Y(_05170_),
    .A1(_05149_),
    .A2(_05168_));
 sg13g2_a22oi_1 _14131_ (.Y(_05171_),
    .B1(_05148_),
    .B2(_05170_),
    .A2(_05133_),
    .A1(net356));
 sg13g2_inv_1 _14132_ (.Y(_00284_),
    .A(_05171_));
 sg13g2_buf_2 _14133_ (.A(\grid.cell_10_0.out ),
    .X(_05172_));
 sg13g2_buf_1 _14134_ (.A(_05172_),
    .X(_05173_));
 sg13g2_nand2_1 _14135_ (.Y(_05174_),
    .A(_00018_),
    .B(_02000_));
 sg13g2_buf_1 _14136_ (.A(_05174_),
    .X(_05175_));
 sg13g2_mux2_1 _14137_ (.A0(net3),
    .A1(_01622_),
    .S(_01471_),
    .X(_05176_));
 sg13g2_buf_4 _14138_ (.X(_05177_),
    .A(_05176_));
 sg13g2_mux2_1 _14139_ (.A0(net4),
    .A1(net1190),
    .S(_01471_),
    .X(_05178_));
 sg13g2_buf_4 _14140_ (.X(_05179_),
    .A(_05178_));
 sg13g2_nor2b_2 _14141_ (.A(_05177_),
    .B_N(_05179_),
    .Y(_05180_));
 sg13g2_nand2_1 _14142_ (.Y(_05181_),
    .A(_05175_),
    .B(_05180_));
 sg13g2_buf_2 _14143_ (.A(_05181_),
    .X(_05182_));
 sg13g2_nor2b_2 _14144_ (.A(_01935_),
    .B_N(_01956_),
    .Y(_05183_));
 sg13g2_nand2_1 _14145_ (.Y(_05184_),
    .A(net177),
    .B(_05183_));
 sg13g2_buf_2 _14146_ (.A(_05184_),
    .X(_05185_));
 sg13g2_or2_1 _14147_ (.X(_05186_),
    .B(_05185_),
    .A(_05182_));
 sg13g2_buf_2 _14148_ (.A(_05186_),
    .X(_05187_));
 sg13g2_buf_1 _14149_ (.A(\grid.cell_10_0.ne ),
    .X(_05188_));
 sg13g2_buf_2 _14150_ (.A(_05188_),
    .X(_05189_));
 sg13g2_buf_1 _14151_ (.A(net1016),
    .X(_05190_));
 sg13g2_buf_1 _14152_ (.A(\grid.cell_10_0.sw ),
    .X(_05191_));
 sg13g2_buf_1 _14153_ (.A(_05191_),
    .X(_05192_));
 sg13g2_buf_1 _14154_ (.A(net1015),
    .X(_05193_));
 sg13g2_buf_1 _14155_ (.A(net681),
    .X(_05194_));
 sg13g2_buf_2 _14156_ (.A(\grid.cell_10_0.w ),
    .X(_05195_));
 sg13g2_buf_1 _14157_ (.A(_05195_),
    .X(_05196_));
 sg13g2_buf_1 _14158_ (.A(net1014),
    .X(_05197_));
 sg13g2_xnor2_1 _14159_ (.Y(_05198_),
    .A(_05194_),
    .B(net680));
 sg13g2_inv_1 _14160_ (.Y(_05199_),
    .A(net1015));
 sg13g2_inv_1 _14161_ (.Y(_05200_),
    .A(net1014));
 sg13g2_nor2_1 _14162_ (.A(net679),
    .B(net678),
    .Y(_05201_));
 sg13g2_buf_2 _14163_ (.A(\grid.cell_10_0.nw ),
    .X(_05202_));
 sg13g2_buf_1 _14164_ (.A(_05202_),
    .X(_05203_));
 sg13g2_buf_1 _14165_ (.A(net1013),
    .X(_05204_));
 sg13g2_buf_1 _14166_ (.A(_05204_),
    .X(_05205_));
 sg13g2_o21ai_1 _14167_ (.B1(net354),
    .Y(_05206_),
    .A1(net682),
    .A2(_05201_));
 sg13g2_a21oi_1 _14168_ (.A1(net682),
    .A2(_05198_),
    .Y(_05207_),
    .B1(_05206_));
 sg13g2_nand2_1 _14169_ (.Y(_05208_),
    .A(net355),
    .B(net680));
 sg13g2_buf_1 _14170_ (.A(_05203_),
    .X(_05209_));
 sg13g2_buf_1 _14171_ (.A(net1016),
    .X(_05210_));
 sg13g2_nand2b_1 _14172_ (.Y(_05211_),
    .B(net675),
    .A_N(net676));
 sg13g2_nor2_1 _14173_ (.A(_05208_),
    .B(_05211_),
    .Y(_05212_));
 sg13g2_buf_1 _14174_ (.A(\grid.cell_10_0.s ),
    .X(_05213_));
 sg13g2_buf_1 _14175_ (.A(_05213_),
    .X(_05214_));
 sg13g2_buf_1 _14176_ (.A(net1012),
    .X(_05215_));
 sg13g2_buf_1 _14177_ (.A(_05215_),
    .X(_05216_));
 sg13g2_o21ai_1 _14178_ (.B1(_05216_),
    .Y(_05217_),
    .A1(_05207_),
    .A2(_05212_));
 sg13g2_buf_1 _14179_ (.A(_00243_),
    .X(_05218_));
 sg13g2_buf_1 _14180_ (.A(_05218_),
    .X(_05219_));
 sg13g2_buf_1 _14181_ (.A(_00247_),
    .X(_05220_));
 sg13g2_buf_1 _14182_ (.A(_05220_),
    .X(_05221_));
 sg13g2_xnor2_1 _14183_ (.Y(_05222_),
    .A(_05195_),
    .B(_05202_));
 sg13g2_xnor2_1 _14184_ (.Y(_05223_),
    .A(net1015),
    .B(_05222_));
 sg13g2_xor2_1 _14185_ (.B(_05188_),
    .A(_05213_),
    .X(_05224_));
 sg13g2_xnor2_1 _14186_ (.Y(_05225_),
    .A(_05223_),
    .B(_05224_));
 sg13g2_buf_2 _14187_ (.A(\grid.cell_10_0.e ),
    .X(_05226_));
 sg13g2_buf_1 _14188_ (.A(_05226_),
    .X(_05227_));
 sg13g2_buf_2 _14189_ (.A(\grid.cell_10_0.se ),
    .X(_05228_));
 sg13g2_buf_1 _14190_ (.A(_05228_),
    .X(_05229_));
 sg13g2_xor2_1 _14191_ (.B(net1008),
    .A(net1009),
    .X(_05230_));
 sg13g2_nor4_1 _14192_ (.A(net1011),
    .B(net1010),
    .C(_05225_),
    .D(_05230_),
    .Y(_05231_));
 sg13g2_buf_1 _14193_ (.A(_00171_),
    .X(_05232_));
 sg13g2_buf_1 _14194_ (.A(_05232_),
    .X(_05233_));
 sg13g2_nand3_1 _14195_ (.B(_05193_),
    .C(net676),
    .A(net675),
    .Y(_05234_));
 sg13g2_nor2_1 _14196_ (.A(_05233_),
    .B(_05234_),
    .Y(_05235_));
 sg13g2_nor3_1 _14197_ (.A(net368),
    .B(_05231_),
    .C(_05235_),
    .Y(_05236_));
 sg13g2_nand2_1 _14198_ (.Y(_05237_),
    .A(_05217_),
    .B(_05236_));
 sg13g2_inv_1 _14199_ (.Y(_05238_),
    .A(net1009));
 sg13g2_buf_1 _14200_ (.A(_05238_),
    .X(_05239_));
 sg13g2_nand2_1 _14201_ (.Y(_05240_),
    .A(net352),
    .B(net1010));
 sg13g2_buf_1 _14202_ (.A(net1008),
    .X(_05241_));
 sg13g2_xnor2_1 _14203_ (.Y(_05242_),
    .A(net673),
    .B(_05225_));
 sg13g2_inv_2 _14204_ (.Y(_05243_),
    .A(_05220_));
 sg13g2_nand2_1 _14205_ (.Y(_05244_),
    .A(_05227_),
    .B(_05243_));
 sg13g2_o21ai_1 _14206_ (.B1(_05244_),
    .Y(_05245_),
    .A1(net1011),
    .A2(_05225_));
 sg13g2_a21oi_1 _14207_ (.A1(_05240_),
    .A2(_05242_),
    .Y(_05246_),
    .B1(_05245_));
 sg13g2_inv_2 _14208_ (.Y(_05247_),
    .A(_05213_));
 sg13g2_or2_1 _14209_ (.X(_05248_),
    .B(_05234_),
    .A(_05247_));
 sg13g2_inv_2 _14210_ (.Y(_05249_),
    .A(_05189_));
 sg13g2_buf_1 _14211_ (.A(_05249_),
    .X(_05250_));
 sg13g2_nor2_1 _14212_ (.A(_05193_),
    .B(net1013),
    .Y(_05251_));
 sg13g2_nand2_1 _14213_ (.Y(_05252_),
    .A(_05250_),
    .B(_05251_));
 sg13g2_a21oi_1 _14214_ (.A1(_05248_),
    .A2(_05252_),
    .Y(_05253_),
    .B1(net680));
 sg13g2_xor2_1 _14215_ (.B(net1007),
    .A(net1016),
    .X(_05254_));
 sg13g2_nand2b_1 _14216_ (.Y(_05255_),
    .B(_05254_),
    .A_N(_05251_));
 sg13g2_nand2_1 _14217_ (.Y(_05256_),
    .A(_05192_),
    .B(net1013));
 sg13g2_nand2b_1 _14218_ (.Y(_05257_),
    .B(_05249_),
    .A_N(_05256_));
 sg13g2_nand3_1 _14219_ (.B(net1007),
    .C(_05256_),
    .A(net682),
    .Y(_05258_));
 sg13g2_nand3_1 _14220_ (.B(_05257_),
    .C(_05258_),
    .A(_05255_),
    .Y(_05259_));
 sg13g2_and3_1 _14221_ (.X(_05260_),
    .A(net674),
    .B(_05197_),
    .C(_05259_));
 sg13g2_a21oi_1 _14222_ (.A1(net1007),
    .A2(_05256_),
    .Y(_05261_),
    .B1(_05251_));
 sg13g2_nand2_1 _14223_ (.Y(_05262_),
    .A(net1007),
    .B(_05251_));
 sg13g2_o21ai_1 _14224_ (.B1(_05262_),
    .Y(_05263_),
    .A1(net682),
    .A2(_05261_));
 sg13g2_and2_1 _14225_ (.A(_05247_),
    .B(_05263_),
    .X(_05264_));
 sg13g2_nor4_1 _14226_ (.A(_05235_),
    .B(_05253_),
    .C(_05260_),
    .D(_05264_),
    .Y(_05265_));
 sg13g2_xor2_1 _14227_ (.B(_05265_),
    .A(_05246_),
    .X(_05266_));
 sg13g2_buf_2 _14228_ (.A(net172),
    .X(_05267_));
 sg13g2_buf_1 _14229_ (.A(net118),
    .X(_05268_));
 sg13g2_o21ai_1 _14230_ (.B1(_05268_),
    .Y(_05269_),
    .A1(_05237_),
    .A2(_05266_));
 sg13g2_nand3_1 _14231_ (.B(_05187_),
    .C(_05269_),
    .A(net1017),
    .Y(_05270_));
 sg13g2_nor2_2 _14232_ (.A(_05182_),
    .B(_05185_),
    .Y(_05271_));
 sg13g2_nor2_1 _14233_ (.A(_05237_),
    .B(_05266_),
    .Y(_05272_));
 sg13g2_buf_1 _14234_ (.A(\grid.cell_10_0.n ),
    .X(_05273_));
 sg13g2_buf_1 _14235_ (.A(_05273_),
    .X(_05274_));
 sg13g2_buf_1 _14236_ (.A(_05274_),
    .X(_05275_));
 sg13g2_xor2_1 _14237_ (.B(_05226_),
    .A(_05210_),
    .X(_05276_));
 sg13g2_xnor2_1 _14238_ (.Y(_05277_),
    .A(net1012),
    .B(net1008));
 sg13g2_xor2_1 _14239_ (.B(_05277_),
    .A(_05276_),
    .X(_05278_));
 sg13g2_xnor2_1 _14240_ (.Y(_05279_),
    .A(_05223_),
    .B(_05278_));
 sg13g2_xnor2_1 _14241_ (.Y(_05280_),
    .A(net672),
    .B(_05279_));
 sg13g2_nor2_1 _14242_ (.A(_05271_),
    .B(_05280_),
    .Y(_05281_));
 sg13g2_a22oi_1 _14243_ (.Y(_05282_),
    .B1(_05272_),
    .B2(_05281_),
    .A2(_05271_),
    .A1(_01806_));
 sg13g2_buf_1 _14244_ (.A(net715),
    .X(_05283_));
 sg13g2_a21oi_1 _14245_ (.A1(_05270_),
    .A2(_05282_),
    .Y(_00285_),
    .B1(net350));
 sg13g2_buf_2 _14246_ (.A(\grid.cell_10_1.e ),
    .X(_05284_));
 sg13g2_buf_2 _14247_ (.A(\grid.cell_10_1.se ),
    .X(_05285_));
 sg13g2_xnor2_1 _14248_ (.Y(_05286_),
    .A(_05284_),
    .B(_05285_));
 sg13g2_buf_2 _14249_ (.A(\grid.cell_10_1.ne ),
    .X(_05287_));
 sg13g2_xnor2_1 _14250_ (.Y(_05288_),
    .A(_05228_),
    .B(_05287_));
 sg13g2_xor2_1 _14251_ (.B(_05288_),
    .A(_05286_),
    .X(_05289_));
 sg13g2_xnor2_1 _14252_ (.Y(_05290_),
    .A(_05224_),
    .B(_05289_));
 sg13g2_buf_1 _14253_ (.A(_05290_),
    .X(_05291_));
 sg13g2_nor2_1 _14254_ (.A(net1010),
    .B(_05291_),
    .Y(_05292_));
 sg13g2_inv_1 _14255_ (.Y(_05293_),
    .A(_05172_));
 sg13g2_buf_1 _14256_ (.A(_05293_),
    .X(_05294_));
 sg13g2_a21o_1 _14257_ (.A2(_05291_),
    .A1(_05294_),
    .B1(net1010),
    .X(_05295_));
 sg13g2_inv_1 _14258_ (.Y(_05296_),
    .A(_05285_));
 sg13g2_buf_1 _14259_ (.A(_05296_),
    .X(_05297_));
 sg13g2_xnor2_1 _14260_ (.Y(_05298_),
    .A(_05287_),
    .B(_05284_));
 sg13g2_xor2_1 _14261_ (.B(_05298_),
    .A(_05224_),
    .X(_05299_));
 sg13g2_xnor2_1 _14262_ (.Y(_05300_),
    .A(net670),
    .B(_05299_));
 sg13g2_nor2_1 _14263_ (.A(_05219_),
    .B(_05300_),
    .Y(_05301_));
 sg13g2_mux2_1 _14264_ (.A0(_05292_),
    .A1(_05295_),
    .S(_05301_),
    .X(_05302_));
 sg13g2_nand2_1 _14265_ (.Y(_05303_),
    .A(_05287_),
    .B(_05284_));
 sg13g2_mux2_1 _14266_ (.A0(_05298_),
    .A1(_05303_),
    .S(_05249_),
    .X(_05304_));
 sg13g2_buf_1 _14267_ (.A(_05287_),
    .X(_05305_));
 sg13g2_buf_1 _14268_ (.A(net1005),
    .X(_05306_));
 sg13g2_buf_1 _14269_ (.A(_05284_),
    .X(_05307_));
 sg13g2_nand4_1 _14270_ (.B(net669),
    .C(net1004),
    .A(net675),
    .Y(_05308_),
    .D(_05296_));
 sg13g2_o21ai_1 _14271_ (.B1(_05308_),
    .Y(_05309_),
    .A1(_05297_),
    .A2(_05304_));
 sg13g2_buf_1 _14272_ (.A(_00245_),
    .X(_05310_));
 sg13g2_buf_1 _14273_ (.A(_05285_),
    .X(_05311_));
 sg13g2_nand2b_1 _14274_ (.Y(_05312_),
    .B(_05311_),
    .A_N(net1176));
 sg13g2_nand2_1 _14275_ (.Y(_05313_),
    .A(net675),
    .B(net669));
 sg13g2_o21ai_1 _14276_ (.B1(_02755_),
    .Y(_05314_),
    .A1(_05312_),
    .A2(_05313_));
 sg13g2_a21o_1 _14277_ (.A2(_05309_),
    .A1(net674),
    .B1(_05314_),
    .X(_05315_));
 sg13g2_buf_1 _14278_ (.A(_05315_),
    .X(_05316_));
 sg13g2_nand3b_1 _14279_ (.B(net1004),
    .C(net1012),
    .Y(_05317_),
    .A_N(net1003));
 sg13g2_inv_1 _14280_ (.Y(_05318_),
    .A(net1005));
 sg13g2_buf_1 _14281_ (.A(_05318_),
    .X(_05319_));
 sg13g2_a21oi_1 _14282_ (.A1(_05312_),
    .A2(_05317_),
    .Y(_05320_),
    .B1(net349));
 sg13g2_inv_2 _14283_ (.Y(_05321_),
    .A(net1004));
 sg13g2_nor2_1 _14284_ (.A(_05285_),
    .B(net1176),
    .Y(_05322_));
 sg13g2_nor4_1 _14285_ (.A(_05247_),
    .B(net669),
    .C(_05321_),
    .D(_05322_),
    .Y(_05323_));
 sg13g2_nor3_1 _14286_ (.A(net351),
    .B(_05320_),
    .C(_05323_),
    .Y(_05324_));
 sg13g2_nor2_1 _14287_ (.A(_05247_),
    .B(_05321_),
    .Y(_05325_));
 sg13g2_nand2_1 _14288_ (.Y(_05326_),
    .A(net1003),
    .B(net1176));
 sg13g2_o21ai_1 _14289_ (.B1(_05326_),
    .Y(_05327_),
    .A1(_05318_),
    .A2(_05322_));
 sg13g2_nor2b_1 _14290_ (.A(net1003),
    .B_N(net1176),
    .Y(_05328_));
 sg13g2_a21o_1 _14291_ (.A2(_05312_),
    .A1(_05318_),
    .B1(_05328_),
    .X(_05329_));
 sg13g2_a221oi_1 _14292_ (.B2(_05247_),
    .C1(net682),
    .B1(_05329_),
    .A1(_05325_),
    .Y(_05330_),
    .A2(_05327_));
 sg13g2_or2_1 _14293_ (.X(_05331_),
    .B(net1003),
    .A(net1005));
 sg13g2_nand4_1 _14294_ (.B(net1016),
    .C(net1005),
    .A(net1012),
    .Y(_05332_),
    .D(net1003));
 sg13g2_o21ai_1 _14295_ (.B1(_05332_),
    .Y(_05333_),
    .A1(net675),
    .A2(_05331_));
 sg13g2_inv_1 _14296_ (.Y(_05334_),
    .A(net1176));
 sg13g2_nor3_1 _14297_ (.A(net1012),
    .B(_05334_),
    .C(_05331_),
    .Y(_05335_));
 sg13g2_a21oi_1 _14298_ (.A1(_05321_),
    .A2(_05333_),
    .Y(_05336_),
    .B1(_05335_));
 sg13g2_o21ai_1 _14299_ (.B1(_05336_),
    .Y(_05337_),
    .A1(_05324_),
    .A2(_05330_));
 sg13g2_nor2b_1 _14300_ (.A(_05316_),
    .B_N(_05337_),
    .Y(_05338_));
 sg13g2_nor3_1 _14301_ (.A(_05316_),
    .B(_05337_),
    .C(_05301_),
    .Y(_05339_));
 sg13g2_nand2_1 _14302_ (.Y(_05340_),
    .A(net1010),
    .B(_05291_));
 sg13g2_o21ai_1 _14303_ (.B1(_05340_),
    .Y(_05341_),
    .A1(net1017),
    .A2(_05292_));
 sg13g2_or2_1 _14304_ (.X(_05342_),
    .B(_05330_),
    .A(_05324_));
 sg13g2_nor2_1 _14305_ (.A(net671),
    .B(net1010),
    .Y(_05343_));
 sg13g2_o21ai_1 _14306_ (.B1(_05343_),
    .Y(_05344_),
    .A1(_05219_),
    .A2(_05300_));
 sg13g2_or2_1 _14307_ (.X(_05345_),
    .B(_05291_),
    .A(_05294_));
 sg13g2_a221oi_1 _14308_ (.B2(_05345_),
    .C1(_05316_),
    .B1(_05344_),
    .A1(_05336_),
    .Y(_05346_),
    .A2(_05342_));
 sg13g2_a221oi_1 _14309_ (.B2(_05341_),
    .C1(_05346_),
    .B1(_05339_),
    .A1(_05302_),
    .Y(_05347_),
    .A2(_05338_));
 sg13g2_a21oi_1 _14310_ (.A1(net85),
    .A2(_05347_),
    .Y(_05348_),
    .B1(_05239_));
 sg13g2_xnor2_1 _14311_ (.Y(_05349_),
    .A(_05273_),
    .B(_05172_));
 sg13g2_xnor2_1 _14312_ (.Y(_05350_),
    .A(_05291_),
    .B(_05349_));
 sg13g2_o21ai_1 _14313_ (.B1(_05187_),
    .Y(_05351_),
    .A1(_05347_),
    .A2(_05350_));
 sg13g2_nor2_1 _14314_ (.A(_05348_),
    .B(_05351_),
    .Y(_05352_));
 sg13g2_o21ai_1 _14315_ (.B1(_05124_),
    .Y(_05353_),
    .A1(net49),
    .A2(_05187_));
 sg13g2_nor2_1 _14316_ (.A(_05352_),
    .B(_05353_),
    .Y(_00286_));
 sg13g2_buf_1 _14317_ (.A(net1194),
    .X(_05354_));
 sg13g2_buf_2 _14318_ (.A(net1002),
    .X(_05355_));
 sg13g2_nand2_1 _14319_ (.Y(_05356_),
    .A(net668),
    .B(_05271_));
 sg13g2_buf_1 _14320_ (.A(net669),
    .X(_05357_));
 sg13g2_buf_2 _14321_ (.A(\grid.cell_10_2.se ),
    .X(_05358_));
 sg13g2_buf_1 _14322_ (.A(_05358_),
    .X(_05359_));
 sg13g2_buf_1 _14323_ (.A(net1001),
    .X(_05360_));
 sg13g2_buf_2 _14324_ (.A(\grid.cell_10_2.e ),
    .X(_05361_));
 sg13g2_buf_1 _14325_ (.A(_05361_),
    .X(_05362_));
 sg13g2_buf_1 _14326_ (.A(net1000),
    .X(_05363_));
 sg13g2_buf_1 _14327_ (.A(\grid.cell_10_2.ne ),
    .X(_05364_));
 sg13g2_buf_1 _14328_ (.A(_05364_),
    .X(_05365_));
 sg13g2_buf_1 _14329_ (.A(net999),
    .X(_05366_));
 sg13g2_buf_1 _14330_ (.A(net665),
    .X(_05367_));
 sg13g2_nand3_1 _14331_ (.B(net666),
    .C(net347),
    .A(net667),
    .Y(_05368_));
 sg13g2_xor2_1 _14332_ (.B(_05364_),
    .A(_05361_),
    .X(_05369_));
 sg13g2_and2_1 _14333_ (.A(net1001),
    .B(_05369_),
    .X(_05370_));
 sg13g2_nand2_1 _14334_ (.Y(_05371_),
    .A(net1000),
    .B(net665));
 sg13g2_nor2_1 _14335_ (.A(net667),
    .B(_05371_),
    .Y(_05372_));
 sg13g2_o21ai_1 _14336_ (.B1(net348),
    .Y(_05373_),
    .A1(_05370_),
    .A2(_05372_));
 sg13g2_o21ai_1 _14337_ (.B1(_05373_),
    .Y(_05374_),
    .A1(net348),
    .A2(_05368_));
 sg13g2_inv_1 _14338_ (.Y(_05375_),
    .A(_05358_));
 sg13g2_buf_1 _14339_ (.A(_05375_),
    .X(_05376_));
 sg13g2_inv_2 _14340_ (.Y(_05377_),
    .A(net999));
 sg13g2_nor2_1 _14341_ (.A(net664),
    .B(_05377_),
    .Y(_05378_));
 sg13g2_buf_2 _14342_ (.A(_00043_),
    .X(_05379_));
 sg13g2_nor2_1 _14343_ (.A(net349),
    .B(_05379_),
    .Y(_05380_));
 sg13g2_inv_1 _14344_ (.Y(_05381_),
    .A(_00242_));
 sg13g2_inv_1 _14345_ (.Y(_05382_),
    .A(_00249_));
 sg13g2_xnor2_1 _14346_ (.Y(_05383_),
    .A(_05358_),
    .B(_05361_));
 sg13g2_xnor2_1 _14347_ (.Y(_05384_),
    .A(_05288_),
    .B(_05383_));
 sg13g2_xnor2_1 _14348_ (.Y(_05385_),
    .A(net665),
    .B(_05384_));
 sg13g2_buf_1 _14349_ (.A(net1003),
    .X(_05386_));
 sg13g2_buf_1 _14350_ (.A(net663),
    .X(_05387_));
 sg13g2_xnor2_1 _14351_ (.Y(_05388_),
    .A(net1009),
    .B(_05387_));
 sg13g2_and4_1 _14352_ (.A(_05381_),
    .B(_05382_),
    .C(_05385_),
    .D(_05388_),
    .X(_05389_));
 sg13g2_a221oi_1 _14353_ (.B2(_05380_),
    .C1(_05389_),
    .B1(_05378_),
    .A1(net673),
    .Y(_05390_),
    .A2(_05374_));
 sg13g2_inv_2 _14354_ (.Y(_05391_),
    .A(net1000));
 sg13g2_inv_1 _14355_ (.Y(_05392_),
    .A(net1008));
 sg13g2_nor2_1 _14356_ (.A(_05392_),
    .B(net1001),
    .Y(_05393_));
 sg13g2_a221oi_1 _14357_ (.B2(_05393_),
    .C1(_05378_),
    .B1(_05377_),
    .A1(_05229_),
    .Y(_05394_),
    .A2(_05391_));
 sg13g2_nor2_1 _14358_ (.A(net1001),
    .B(net665),
    .Y(_05395_));
 sg13g2_nand2_1 _14359_ (.Y(_05396_),
    .A(_05229_),
    .B(net666));
 sg13g2_a22oi_1 _14360_ (.Y(_05397_),
    .B1(_05395_),
    .B2(_05396_),
    .A2(_05394_),
    .A1(_05379_));
 sg13g2_o21ai_1 _14361_ (.B1(net673),
    .Y(_05398_),
    .A1(net349),
    .A2(_05391_));
 sg13g2_nand3_1 _14362_ (.B(_05395_),
    .C(_05398_),
    .A(_05379_),
    .Y(_05399_));
 sg13g2_o21ai_1 _14363_ (.B1(_05399_),
    .Y(_05400_),
    .A1(net348),
    .A2(_05397_));
 sg13g2_buf_1 _14364_ (.A(net1009),
    .X(_05401_));
 sg13g2_xnor2_1 _14365_ (.Y(_05402_),
    .A(_05285_),
    .B(_05364_));
 sg13g2_xnor2_1 _14366_ (.Y(_05403_),
    .A(_05384_),
    .B(_05402_));
 sg13g2_a21oi_1 _14367_ (.A1(net352),
    .A2(_00249_),
    .Y(_05404_),
    .B1(_05403_));
 sg13g2_a221oi_1 _14368_ (.B2(_05381_),
    .C1(_05404_),
    .B1(_05385_),
    .A1(_05401_),
    .Y(_05405_),
    .A2(_05382_));
 sg13g2_xor2_1 _14369_ (.B(_05405_),
    .A(_05400_),
    .X(_05406_));
 sg13g2_buf_2 _14370_ (.A(net368),
    .X(_05407_));
 sg13g2_buf_1 _14371_ (.A(_05407_),
    .X(_05408_));
 sg13g2_a21oi_1 _14372_ (.A1(_05390_),
    .A2(_05406_),
    .Y(_05409_),
    .B1(net117));
 sg13g2_xnor2_1 _14373_ (.Y(_05410_),
    .A(_05276_),
    .B(_05403_));
 sg13g2_buf_1 _14374_ (.A(net1004),
    .X(_05411_));
 sg13g2_a21oi_1 _14375_ (.A1(net122),
    .A2(_05410_),
    .Y(_05412_),
    .B1(net661));
 sg13g2_nand2_2 _14376_ (.Y(_05413_),
    .A(net1054),
    .B(_05187_));
 sg13g2_or3_1 _14377_ (.A(_05409_),
    .B(_05412_),
    .C(_05413_),
    .X(_05414_));
 sg13g2_o21ai_1 _14378_ (.B1(_05414_),
    .Y(_00287_),
    .A1(net27),
    .A2(_05356_));
 sg13g2_buf_1 _14379_ (.A(net171),
    .X(_05415_));
 sg13g2_buf_2 _14380_ (.A(net116),
    .X(_05416_));
 sg13g2_inv_1 _14381_ (.Y(_05417_),
    .A(_00042_));
 sg13g2_buf_2 _14382_ (.A(\grid.cell_10_3.ne ),
    .X(_05418_));
 sg13g2_buf_1 _14383_ (.A(\grid.cell_10_3.se ),
    .X(_05419_));
 sg13g2_buf_1 _14384_ (.A(\grid.cell_10_3.e ),
    .X(_05420_));
 sg13g2_xnor2_1 _14385_ (.Y(_05421_),
    .A(net1175),
    .B(_05420_));
 sg13g2_xnor2_1 _14386_ (.Y(_05422_),
    .A(_05402_),
    .B(_05421_));
 sg13g2_xnor2_1 _14387_ (.Y(_05423_),
    .A(_05418_),
    .B(_05422_));
 sg13g2_and2_1 _14388_ (.A(_05417_),
    .B(_05423_),
    .X(_05424_));
 sg13g2_buf_1 _14389_ (.A(_05424_),
    .X(_05425_));
 sg13g2_buf_1 _14390_ (.A(_05321_),
    .X(_05426_));
 sg13g2_xnor2_1 _14391_ (.Y(_05427_),
    .A(net1001),
    .B(_05423_));
 sg13g2_buf_1 _14392_ (.A(_05427_),
    .X(_05428_));
 sg13g2_buf_2 _14393_ (.A(_00248_),
    .X(_05429_));
 sg13g2_a21o_1 _14394_ (.A2(_05428_),
    .A1(net345),
    .B1(_05429_),
    .X(_05430_));
 sg13g2_o21ai_1 _14395_ (.B1(_05428_),
    .Y(_05431_),
    .A1(_05429_),
    .A2(_05425_));
 sg13g2_nor3_1 _14396_ (.A(_05429_),
    .B(_05425_),
    .C(_05428_),
    .Y(_05432_));
 sg13g2_a221oi_1 _14397_ (.B2(net661),
    .C1(_05432_),
    .B1(_05431_),
    .A1(_05425_),
    .Y(_05433_),
    .A2(_05430_));
 sg13g2_buf_2 _14398_ (.A(_00075_),
    .X(_05434_));
 sg13g2_buf_1 _14399_ (.A(net1175),
    .X(_05435_));
 sg13g2_buf_1 _14400_ (.A(_05435_),
    .X(_05436_));
 sg13g2_nand2_1 _14401_ (.Y(_05437_),
    .A(_05418_),
    .B(net999));
 sg13g2_buf_1 _14402_ (.A(_05420_),
    .X(_05438_));
 sg13g2_xor2_1 _14403_ (.B(_05364_),
    .A(_05418_),
    .X(_05439_));
 sg13g2_and2_1 _14404_ (.A(net997),
    .B(_05439_),
    .X(_05440_));
 sg13g2_a21oi_1 _14405_ (.A1(net670),
    .A2(_05437_),
    .Y(_05441_),
    .B1(_05440_));
 sg13g2_buf_2 _14406_ (.A(_05418_),
    .X(_05442_));
 sg13g2_inv_1 _14407_ (.Y(_05443_),
    .A(net1175));
 sg13g2_buf_1 _14408_ (.A(_05443_),
    .X(_05444_));
 sg13g2_inv_2 _14409_ (.Y(_05445_),
    .A(net997));
 sg13g2_o21ai_1 _14410_ (.B1(net663),
    .Y(_05446_),
    .A1(_05444_),
    .A2(_05445_));
 sg13g2_nand3b_1 _14411_ (.B(_05377_),
    .C(_05446_),
    .Y(_05447_),
    .A_N(net996));
 sg13g2_o21ai_1 _14412_ (.B1(_05447_),
    .Y(_05448_),
    .A1(net660),
    .A2(_05441_));
 sg13g2_buf_1 _14413_ (.A(net997),
    .X(_05449_));
 sg13g2_nand2_1 _14414_ (.Y(_05450_),
    .A(net346),
    .B(net658));
 sg13g2_buf_1 _14415_ (.A(net996),
    .X(_05451_));
 sg13g2_nor3_1 _14416_ (.A(net660),
    .B(net657),
    .C(net347),
    .Y(_05452_));
 sg13g2_a22oi_1 _14417_ (.Y(_05453_),
    .B1(_05450_),
    .B2(_05452_),
    .A2(_05448_),
    .A1(_05434_));
 sg13g2_or2_1 _14418_ (.X(_05454_),
    .B(_05453_),
    .A(_05433_));
 sg13g2_nand2_1 _14419_ (.Y(_05455_),
    .A(_05429_),
    .B(_05428_));
 sg13g2_o21ai_1 _14420_ (.B1(net345),
    .Y(_05456_),
    .A1(_05429_),
    .A2(_05428_));
 sg13g2_nand2_1 _14421_ (.Y(_05457_),
    .A(net659),
    .B(net997));
 sg13g2_nor2_1 _14422_ (.A(net997),
    .B(_05437_),
    .Y(_05458_));
 sg13g2_o21ai_1 _14423_ (.B1(net998),
    .Y(_05459_),
    .A1(_05440_),
    .A2(_05458_));
 sg13g2_o21ai_1 _14424_ (.B1(_05459_),
    .Y(_05460_),
    .A1(_05437_),
    .A2(_05457_));
 sg13g2_nor3_1 _14425_ (.A(_05434_),
    .B(net659),
    .C(_05437_),
    .Y(_05461_));
 sg13g2_a21oi_1 _14426_ (.A1(net346),
    .A2(_05460_),
    .Y(_05462_),
    .B1(_05461_));
 sg13g2_nand3b_1 _14427_ (.B(_05453_),
    .C(_05462_),
    .Y(_05463_),
    .A_N(_05425_));
 sg13g2_a21o_1 _14428_ (.A2(_05456_),
    .A1(_05455_),
    .B1(_05463_),
    .X(_05464_));
 sg13g2_and3_1 _14429_ (.X(_05465_),
    .A(net82),
    .B(_05454_),
    .C(_05464_));
 sg13g2_xor2_1 _14430_ (.B(_05428_),
    .A(_05298_),
    .X(_05466_));
 sg13g2_a21oi_1 _14431_ (.A1(net122),
    .A2(_05466_),
    .Y(_05467_),
    .B1(net666));
 sg13g2_or2_1 _14432_ (.X(_05468_),
    .B(_05467_),
    .A(_05413_));
 sg13g2_nand2b_1 _14433_ (.Y(_05469_),
    .B(net1054),
    .A_N(net48));
 sg13g2_or2_1 _14434_ (.X(_05470_),
    .B(_05469_),
    .A(_05187_));
 sg13g2_o21ai_1 _14435_ (.B1(_05470_),
    .Y(_00288_),
    .A1(_05465_),
    .A2(_05468_));
 sg13g2_buf_1 _14436_ (.A(_05407_),
    .X(_05471_));
 sg13g2_buf_1 _14437_ (.A(net115),
    .X(_05472_));
 sg13g2_buf_2 _14438_ (.A(_00040_),
    .X(_05473_));
 sg13g2_nand2_1 _14439_ (.Y(_05474_),
    .A(_05473_),
    .B(_05391_));
 sg13g2_buf_1 _14440_ (.A(\grid.cell_10_4.se ),
    .X(_05475_));
 sg13g2_buf_1 _14441_ (.A(_05475_),
    .X(_05476_));
 sg13g2_buf_1 _14442_ (.A(\grid.cell_10_4.e ),
    .X(_05477_));
 sg13g2_buf_2 _14443_ (.A(\grid.cell_10_4.ne ),
    .X(_05478_));
 sg13g2_xor2_1 _14444_ (.B(_05478_),
    .A(_05477_),
    .X(_05479_));
 sg13g2_xnor2_1 _14445_ (.Y(_05480_),
    .A(_05358_),
    .B(_05418_));
 sg13g2_xnor2_1 _14446_ (.Y(_05481_),
    .A(_05479_),
    .B(_05480_));
 sg13g2_xnor2_1 _14447_ (.Y(_05482_),
    .A(net995),
    .B(_05481_));
 sg13g2_xnor2_1 _14448_ (.Y(_05483_),
    .A(net660),
    .B(_05482_));
 sg13g2_buf_1 _14449_ (.A(_00074_),
    .X(_05484_));
 sg13g2_nand2b_1 _14450_ (.Y(_05485_),
    .B(net666),
    .A_N(_05473_));
 sg13g2_o21ai_1 _14451_ (.B1(_05485_),
    .Y(_05486_),
    .A1(_05484_),
    .A2(_05482_));
 sg13g2_a21oi_1 _14452_ (.A1(_05474_),
    .A2(_05483_),
    .Y(_05487_),
    .B1(_05486_));
 sg13g2_buf_2 _14453_ (.A(_00107_),
    .X(_05488_));
 sg13g2_buf_1 _14454_ (.A(net995),
    .X(_05489_));
 sg13g2_buf_1 _14455_ (.A(net656),
    .X(_05490_));
 sg13g2_buf_1 _14456_ (.A(_05477_),
    .X(_05491_));
 sg13g2_buf_1 _14457_ (.A(net994),
    .X(_05492_));
 sg13g2_buf_1 _14458_ (.A(_05478_),
    .X(_05493_));
 sg13g2_xor2_1 _14459_ (.B(net996),
    .A(net993),
    .X(_05494_));
 sg13g2_nand2_1 _14460_ (.Y(_05495_),
    .A(net993),
    .B(net996));
 sg13g2_a22oi_1 _14461_ (.Y(_05496_),
    .B1(_05495_),
    .B2(net664),
    .A2(_05494_),
    .A1(net655));
 sg13g2_buf_1 _14462_ (.A(net993),
    .X(_05497_));
 sg13g2_a21oi_1 _14463_ (.A1(net995),
    .A2(net994),
    .Y(_05498_),
    .B1(net664));
 sg13g2_or3_1 _14464_ (.A(net654),
    .B(net996),
    .C(_05498_),
    .X(_05499_));
 sg13g2_o21ai_1 _14465_ (.B1(_05499_),
    .Y(_05500_),
    .A1(net344),
    .A2(_05496_));
 sg13g2_nand2_1 _14466_ (.Y(_05501_),
    .A(net667),
    .B(_05492_));
 sg13g2_buf_1 _14467_ (.A(net654),
    .X(_05502_));
 sg13g2_nor3_1 _14468_ (.A(net344),
    .B(net343),
    .C(net657),
    .Y(_05503_));
 sg13g2_a22oi_1 _14469_ (.Y(_05504_),
    .B1(_05501_),
    .B2(_05503_),
    .A2(_05500_),
    .A1(_05488_));
 sg13g2_xor2_1 _14470_ (.B(_05504_),
    .A(_05487_),
    .X(_05505_));
 sg13g2_inv_2 _14471_ (.Y(_05506_),
    .A(_05475_));
 sg13g2_buf_1 _14472_ (.A(net655),
    .X(_05507_));
 sg13g2_nand2_1 _14473_ (.Y(_05508_),
    .A(net655),
    .B(_05494_));
 sg13g2_o21ai_1 _14474_ (.B1(_05508_),
    .Y(_05509_),
    .A1(net342),
    .A2(_05495_));
 sg13g2_nor2_1 _14475_ (.A(_05488_),
    .B(_05495_),
    .Y(_05510_));
 sg13g2_a21oi_1 _14476_ (.A1(net667),
    .A2(_05509_),
    .Y(_05511_),
    .B1(_05510_));
 sg13g2_nor2_1 _14477_ (.A(_05506_),
    .B(_05511_),
    .Y(_05512_));
 sg13g2_nor3_1 _14478_ (.A(net344),
    .B(_05495_),
    .C(_05501_),
    .Y(_05513_));
 sg13g2_xor2_1 _14479_ (.B(net1000),
    .A(net1175),
    .X(_05514_));
 sg13g2_nor4_1 _14480_ (.A(_05473_),
    .B(_05484_),
    .C(_05482_),
    .D(_05514_),
    .Y(_05515_));
 sg13g2_nor4_1 _14481_ (.A(_05505_),
    .B(_05512_),
    .C(_05513_),
    .D(_05515_),
    .Y(_05516_));
 sg13g2_buf_1 _14482_ (.A(net171),
    .X(_05517_));
 sg13g2_xnor2_1 _14483_ (.Y(_05518_),
    .A(_05377_),
    .B(_05514_));
 sg13g2_xnor2_1 _14484_ (.Y(_05519_),
    .A(_05482_),
    .B(_05518_));
 sg13g2_a21oi_1 _14485_ (.A1(net114),
    .A2(_05519_),
    .Y(_05520_),
    .B1(net658));
 sg13g2_nor2_1 _14486_ (.A(_05413_),
    .B(_05520_),
    .Y(_05521_));
 sg13g2_o21ai_1 _14487_ (.B1(_05521_),
    .Y(_05522_),
    .A1(net81),
    .A2(_05516_));
 sg13g2_o21ai_1 _14488_ (.B1(_05522_),
    .Y(_00289_),
    .A1(net34),
    .A2(_05356_));
 sg13g2_buf_2 _14489_ (.A(\grid.cell_10_5.se ),
    .X(_05523_));
 sg13g2_buf_1 _14490_ (.A(_05523_),
    .X(_05524_));
 sg13g2_buf_1 _14491_ (.A(net992),
    .X(_05525_));
 sg13g2_buf_1 _14492_ (.A(net653),
    .X(_05526_));
 sg13g2_buf_1 _14493_ (.A(net341),
    .X(_05527_));
 sg13g2_buf_1 _14494_ (.A(_00139_),
    .X(_05528_));
 sg13g2_buf_1 _14495_ (.A(_05528_),
    .X(_05529_));
 sg13g2_buf_1 _14496_ (.A(net991),
    .X(_05530_));
 sg13g2_buf_1 _14497_ (.A(\grid.cell_10_5.ne ),
    .X(_05531_));
 sg13g2_buf_1 _14498_ (.A(_05531_),
    .X(_05532_));
 sg13g2_nand2_1 _14499_ (.Y(_05533_),
    .A(net990),
    .B(net993));
 sg13g2_buf_1 _14500_ (.A(\grid.cell_10_5.e ),
    .X(_05534_));
 sg13g2_buf_8 _14501_ (.A(_05534_),
    .X(_05535_));
 sg13g2_buf_1 _14502_ (.A(net989),
    .X(_05536_));
 sg13g2_buf_1 _14503_ (.A(net651),
    .X(_05537_));
 sg13g2_xor2_1 _14504_ (.B(_05478_),
    .A(_05531_),
    .X(_05538_));
 sg13g2_nand2_1 _14505_ (.Y(_05539_),
    .A(net651),
    .B(_05538_));
 sg13g2_o21ai_1 _14506_ (.B1(_05539_),
    .Y(_05540_),
    .A1(net340),
    .A2(_05533_));
 sg13g2_nand2_1 _14507_ (.Y(_05541_),
    .A(_05436_),
    .B(_05540_));
 sg13g2_o21ai_1 _14508_ (.B1(_05541_),
    .Y(_05542_),
    .A1(net652),
    .A2(_05533_));
 sg13g2_nand2_1 _14509_ (.Y(_05543_),
    .A(_05435_),
    .B(net651));
 sg13g2_nor3_1 _14510_ (.A(net162),
    .B(_05533_),
    .C(_05543_),
    .Y(_05544_));
 sg13g2_a21oi_1 _14511_ (.A1(net162),
    .A2(_05542_),
    .Y(_05545_),
    .B1(_05544_));
 sg13g2_buf_1 _14512_ (.A(_00072_),
    .X(_05546_));
 sg13g2_xnor2_1 _14513_ (.Y(_05547_),
    .A(_05523_),
    .B(_05534_));
 sg13g2_xor2_1 _14514_ (.B(_05547_),
    .A(_05538_),
    .X(_05548_));
 sg13g2_xnor2_1 _14515_ (.Y(_05549_),
    .A(_05506_),
    .B(_05421_));
 sg13g2_xnor2_1 _14516_ (.Y(_05550_),
    .A(_05548_),
    .B(_05549_));
 sg13g2_or2_1 _14517_ (.X(_05551_),
    .B(_05550_),
    .A(_05546_));
 sg13g2_nor2_1 _14518_ (.A(_05506_),
    .B(_05445_),
    .Y(_05552_));
 sg13g2_buf_1 _14519_ (.A(_00106_),
    .X(_05553_));
 sg13g2_o21ai_1 _14520_ (.B1(_05553_),
    .Y(_05554_),
    .A1(net995),
    .A2(_05445_));
 sg13g2_xnor2_1 _14521_ (.Y(_05555_),
    .A(_05419_),
    .B(_05548_));
 sg13g2_mux2_1 _14522_ (.A0(_05552_),
    .A1(_05554_),
    .S(_05555_),
    .X(_05556_));
 sg13g2_a22oi_1 _14523_ (.Y(_05557_),
    .B1(_05533_),
    .B2(_05443_),
    .A2(_05538_),
    .A1(net989));
 sg13g2_nand2_1 _14524_ (.Y(_05558_),
    .A(_05523_),
    .B(net989));
 sg13g2_or2_1 _14525_ (.X(_05559_),
    .B(net993),
    .A(net990));
 sg13g2_a21o_1 _14526_ (.A2(_05558_),
    .A1(net1175),
    .B1(_05559_),
    .X(_05560_));
 sg13g2_o21ai_1 _14527_ (.B1(_05560_),
    .Y(_05561_),
    .A1(_05524_),
    .A2(_05557_));
 sg13g2_nor2_1 _14528_ (.A(net653),
    .B(_05559_),
    .Y(_05562_));
 sg13g2_a22oi_1 _14529_ (.Y(_05563_),
    .B1(_05562_),
    .B2(_05543_),
    .A2(_05561_),
    .A1(net991));
 sg13g2_xor2_1 _14530_ (.B(_05563_),
    .A(_05556_),
    .X(_05564_));
 sg13g2_nor3_1 _14531_ (.A(_05556_),
    .B(_05563_),
    .C(_05551_),
    .Y(_05565_));
 sg13g2_a21o_1 _14532_ (.A2(_05564_),
    .A1(_05551_),
    .B1(_05565_),
    .X(_05566_));
 sg13g2_a21oi_1 _14533_ (.A1(_05545_),
    .A2(_05566_),
    .Y(_05567_),
    .B1(net124));
 sg13g2_buf_1 _14534_ (.A(net657),
    .X(_05568_));
 sg13g2_xnor2_1 _14535_ (.Y(_05569_),
    .A(_05568_),
    .B(_05550_));
 sg13g2_a21oi_1 _14536_ (.A1(net84),
    .A2(_05569_),
    .Y(_05570_),
    .B1(net342));
 sg13g2_or3_1 _14537_ (.A(_05413_),
    .B(_05567_),
    .C(_05570_),
    .X(_05571_));
 sg13g2_o21ai_1 _14538_ (.B1(_05571_),
    .Y(_00290_),
    .A1(net46),
    .A2(_05356_));
 sg13g2_xor2_1 _14539_ (.B(net990),
    .A(net995),
    .X(_05572_));
 sg13g2_xnor2_1 _14540_ (.Y(_05573_),
    .A(_05223_),
    .B(_05572_));
 sg13g2_buf_1 _14541_ (.A(_05573_),
    .X(_05574_));
 sg13g2_buf_1 _14542_ (.A(_00104_),
    .X(_05575_));
 sg13g2_inv_1 _14543_ (.Y(_05576_),
    .A(_05575_));
 sg13g2_or2_1 _14544_ (.X(_05577_),
    .B(_05202_),
    .A(net990));
 sg13g2_buf_1 _14545_ (.A(_05577_),
    .X(_05578_));
 sg13g2_and2_1 _14546_ (.A(_05532_),
    .B(_05203_),
    .X(_05579_));
 sg13g2_buf_1 _14547_ (.A(_05579_),
    .X(_05580_));
 sg13g2_a21oi_1 _14548_ (.A1(net681),
    .A2(_05578_),
    .Y(_05581_),
    .B1(_05580_));
 sg13g2_nor3_1 _14549_ (.A(net1015),
    .B(net990),
    .C(net1013),
    .Y(_05582_));
 sg13g2_a21oi_1 _14550_ (.A1(net1007),
    .A2(_05581_),
    .Y(_05583_),
    .B1(_05582_));
 sg13g2_nand2_1 _14551_ (.Y(_05584_),
    .A(net1007),
    .B(net681));
 sg13g2_nand2_1 _14552_ (.Y(_05585_),
    .A(net990),
    .B(net1013));
 sg13g2_mux2_1 _14553_ (.A0(net1007),
    .A1(_05584_),
    .S(_05585_),
    .X(_05586_));
 sg13g2_xor2_1 _14554_ (.B(net681),
    .A(_05232_),
    .X(_05587_));
 sg13g2_nand2_1 _14555_ (.Y(_05588_),
    .A(_05578_),
    .B(_05587_));
 sg13g2_nand2_1 _14556_ (.Y(_05589_),
    .A(_05476_),
    .B(net1014));
 sg13g2_a21oi_1 _14557_ (.A1(_05586_),
    .A2(_05588_),
    .Y(_05590_),
    .B1(_05589_));
 sg13g2_and3_1 _14558_ (.X(_05591_),
    .A(net1015),
    .B(net990),
    .C(_05202_));
 sg13g2_buf_1 _14559_ (.A(_05591_),
    .X(_05592_));
 sg13g2_a21oi_1 _14560_ (.A1(_05476_),
    .A2(_05592_),
    .Y(_05593_),
    .B1(_05582_));
 sg13g2_inv_1 _14561_ (.Y(_05594_),
    .A(net1007));
 sg13g2_nand2_1 _14562_ (.Y(_05595_),
    .A(_05594_),
    .B(_05592_));
 sg13g2_o21ai_1 _14563_ (.B1(_05595_),
    .Y(_05596_),
    .A1(net1014),
    .A2(_05593_));
 sg13g2_nor2_1 _14564_ (.A(_05590_),
    .B(_05596_),
    .Y(_05597_));
 sg13g2_o21ai_1 _14565_ (.B1(_05597_),
    .Y(_05598_),
    .A1(_05489_),
    .A2(_05583_));
 sg13g2_buf_1 _14566_ (.A(_05598_),
    .X(_05599_));
 sg13g2_buf_1 _14567_ (.A(_00138_),
    .X(_05600_));
 sg13g2_buf_1 _14568_ (.A(_05600_),
    .X(_05601_));
 sg13g2_nand3b_1 _14569_ (.B(net162),
    .C(net342),
    .Y(_05602_),
    .A_N(net988));
 sg13g2_o21ai_1 _14570_ (.B1(_05602_),
    .Y(_05603_),
    .A1(net162),
    .A2(_05599_));
 sg13g2_inv_2 _14571_ (.Y(_05604_),
    .A(net994));
 sg13g2_o21ai_1 _14572_ (.B1(net988),
    .Y(_05605_),
    .A1(net162),
    .A2(_05604_));
 sg13g2_nor2b_1 _14573_ (.A(_05599_),
    .B_N(_05605_),
    .Y(_05606_));
 sg13g2_a21oi_1 _14574_ (.A1(_05576_),
    .A2(_05603_),
    .Y(_05607_),
    .B1(_05606_));
 sg13g2_or2_1 _14575_ (.X(_05608_),
    .B(_05607_),
    .A(_05574_));
 sg13g2_nor3_1 _14576_ (.A(_05575_),
    .B(net988),
    .C(net341),
    .Y(_05609_));
 sg13g2_o21ai_1 _14577_ (.B1(_05575_),
    .Y(_05610_),
    .A1(net988),
    .A2(_05574_));
 sg13g2_nand2b_1 _14578_ (.Y(_05611_),
    .B(_05610_),
    .A_N(_05609_));
 sg13g2_a21oi_1 _14579_ (.A1(net988),
    .A2(net341),
    .Y(_05612_),
    .B1(_05574_));
 sg13g2_a221oi_1 _14580_ (.B2(net162),
    .C1(_05612_),
    .B1(_05574_),
    .A1(_05576_),
    .Y(_05613_),
    .A2(net342));
 sg13g2_a21oi_1 _14581_ (.A1(_05604_),
    .A2(_05611_),
    .Y(_05614_),
    .B1(_05613_));
 sg13g2_and2_1 _14582_ (.A(_05527_),
    .B(_05574_),
    .X(_05615_));
 sg13g2_o21ai_1 _14583_ (.B1(_05576_),
    .Y(_05616_),
    .A1(net342),
    .A2(_05615_));
 sg13g2_a21oi_1 _14584_ (.A1(_05507_),
    .A2(_05615_),
    .Y(_05617_),
    .B1(_05599_));
 sg13g2_a22oi_1 _14585_ (.Y(_05618_),
    .B1(_05616_),
    .B2(_05617_),
    .A2(_05614_),
    .A1(_05599_));
 sg13g2_buf_1 _14586_ (.A(net167),
    .X(_05619_));
 sg13g2_xor2_1 _14587_ (.B(_05479_),
    .A(_05527_),
    .X(_05620_));
 sg13g2_xnor2_1 _14588_ (.Y(_05621_),
    .A(_05574_),
    .B(_05620_));
 sg13g2_a21oi_1 _14589_ (.A1(net113),
    .A2(_05621_),
    .Y(_05622_),
    .B1(_05537_));
 sg13g2_or2_1 _14590_ (.X(_05623_),
    .B(_05589_),
    .A(_05585_));
 sg13g2_buf_1 _14591_ (.A(net680),
    .X(_05624_));
 sg13g2_buf_1 _14592_ (.A(_05532_),
    .X(_05625_));
 sg13g2_buf_1 _14593_ (.A(net650),
    .X(_05626_));
 sg13g2_buf_1 _14594_ (.A(_05204_),
    .X(_05627_));
 sg13g2_xor2_1 _14595_ (.B(net336),
    .A(_05626_),
    .X(_05628_));
 sg13g2_nand2_1 _14596_ (.Y(_05629_),
    .A(net338),
    .B(_05628_));
 sg13g2_o21ai_1 _14597_ (.B1(_05629_),
    .Y(_05630_),
    .A1(net338),
    .A2(_05585_));
 sg13g2_a221oi_1 _14598_ (.B2(_05490_),
    .C1(net679),
    .B1(_05630_),
    .A1(_05594_),
    .Y(_05631_),
    .A2(_05580_));
 sg13g2_a21oi_1 _14599_ (.A1(net679),
    .A2(_05623_),
    .Y(_05632_),
    .B1(_05631_));
 sg13g2_nor4_1 _14600_ (.A(_05413_),
    .B(_05618_),
    .C(_05622_),
    .D(_05632_),
    .Y(_05633_));
 sg13g2_inv_1 _14601_ (.Y(_05634_),
    .A(net989));
 sg13g2_nor3_1 _14602_ (.A(net649),
    .B(_05136_),
    .C(_05271_),
    .Y(_05635_));
 sg13g2_a21oi_1 _14603_ (.A1(_05119_),
    .A2(_05271_),
    .Y(_05636_),
    .B1(_05635_));
 sg13g2_nor2_1 _14604_ (.A(net715),
    .B(_05636_),
    .Y(_05637_));
 sg13g2_a21o_1 _14605_ (.A2(_05633_),
    .A1(_05608_),
    .B1(_05637_),
    .X(_00291_));
 sg13g2_xor2_1 _14606_ (.B(_05531_),
    .A(net989),
    .X(_05638_));
 sg13g2_xnor2_1 _14607_ (.Y(_05639_),
    .A(_05191_),
    .B(_05202_));
 sg13g2_xnor2_1 _14608_ (.Y(_05640_),
    .A(_05638_),
    .B(_05639_));
 sg13g2_xnor2_1 _14609_ (.Y(_05641_),
    .A(net1012),
    .B(_05640_));
 sg13g2_xor2_1 _14610_ (.B(net341),
    .A(net1017),
    .X(_05642_));
 sg13g2_nor4_1 _14611_ (.A(net988),
    .B(net1010),
    .C(_05641_),
    .D(_05642_),
    .Y(_05643_));
 sg13g2_inv_1 _14612_ (.Y(_05644_),
    .A(_05528_));
 sg13g2_nand3_1 _14613_ (.B(_05536_),
    .C(_05626_),
    .A(_05194_),
    .Y(_05645_));
 sg13g2_buf_1 _14614_ (.A(net681),
    .X(_05646_));
 sg13g2_and2_1 _14615_ (.A(net335),
    .B(_05638_),
    .X(_05647_));
 sg13g2_inv_1 _14616_ (.Y(_05648_),
    .A(net650));
 sg13g2_nor3_1 _14617_ (.A(net335),
    .B(net649),
    .C(_05648_),
    .Y(_05649_));
 sg13g2_o21ai_1 _14618_ (.B1(net336),
    .Y(_05650_),
    .A1(_05647_),
    .A2(_05649_));
 sg13g2_o21ai_1 _14619_ (.B1(_05650_),
    .Y(_05651_),
    .A1(net354),
    .A2(_05645_));
 sg13g2_a221oi_1 _14620_ (.B2(_05216_),
    .C1(_03810_),
    .B1(_05651_),
    .A1(net987),
    .Y(_05652_),
    .A2(_05592_));
 sg13g2_nand2b_1 _14621_ (.Y(_05653_),
    .B(_05652_),
    .A_N(_05643_));
 sg13g2_nand2_1 _14622_ (.Y(_05654_),
    .A(net671),
    .B(net1010));
 sg13g2_xnor2_1 _14623_ (.Y(_05655_),
    .A(_05525_),
    .B(_05641_));
 sg13g2_nand2_1 _14624_ (.Y(_05656_),
    .A(net1017),
    .B(_05243_));
 sg13g2_o21ai_1 _14625_ (.B1(_05656_),
    .Y(_05657_),
    .A1(_05601_),
    .A2(_05641_));
 sg13g2_a21oi_1 _14626_ (.A1(_05654_),
    .A2(_05655_),
    .Y(_05658_),
    .B1(_05657_));
 sg13g2_nand3_1 _14627_ (.B(net335),
    .C(net651),
    .A(_05214_),
    .Y(_05659_));
 sg13g2_o21ai_1 _14628_ (.B1(_05659_),
    .Y(_05660_),
    .A1(net674),
    .A2(_05646_));
 sg13g2_nand4_1 _14629_ (.B(_05199_),
    .C(net651),
    .A(net674),
    .Y(_05661_),
    .D(_05578_));
 sg13g2_o21ai_1 _14630_ (.B1(_05661_),
    .Y(_05662_),
    .A1(net674),
    .A2(_05578_));
 sg13g2_a21oi_1 _14631_ (.A1(_05585_),
    .A2(_05660_),
    .Y(_05663_),
    .B1(_05662_));
 sg13g2_nand2_1 _14632_ (.Y(_05664_),
    .A(net1012),
    .B(_05535_));
 sg13g2_nand2_1 _14633_ (.Y(_05665_),
    .A(_05646_),
    .B(_05580_));
 sg13g2_o21ai_1 _14634_ (.B1(_05665_),
    .Y(_05666_),
    .A1(_05581_),
    .A2(_05664_));
 sg13g2_a21oi_1 _14635_ (.A1(net674),
    .A2(_05592_),
    .Y(_05667_),
    .B1(_05582_));
 sg13g2_nor2b_1 _14636_ (.A(_05667_),
    .B_N(_05664_),
    .Y(_05668_));
 sg13g2_a21oi_1 _14637_ (.A1(net987),
    .A2(_05666_),
    .Y(_05669_),
    .B1(_05668_));
 sg13g2_o21ai_1 _14638_ (.B1(_05669_),
    .Y(_05670_),
    .A1(_05644_),
    .A2(_05663_));
 sg13g2_xnor2_1 _14639_ (.Y(_05671_),
    .A(_05658_),
    .B(_05670_));
 sg13g2_xor2_1 _14640_ (.B(_05655_),
    .A(_05349_),
    .X(_05672_));
 sg13g2_nor3_1 _14641_ (.A(_05653_),
    .B(_05671_),
    .C(_05672_),
    .Y(_05673_));
 sg13g2_o21ai_1 _14642_ (.B1(net85),
    .Y(_05674_),
    .A1(_05653_),
    .A2(_05671_));
 sg13g2_o21ai_1 _14643_ (.B1(_05674_),
    .Y(_05675_),
    .A1(net338),
    .A2(_05673_));
 sg13g2_a21o_1 _14644_ (.A2(_05126_),
    .A1(net713),
    .B1(_05127_),
    .X(_05676_));
 sg13g2_buf_1 _14645_ (.A(_05676_),
    .X(_05677_));
 sg13g2_buf_2 _14646_ (.A(_05677_),
    .X(_05678_));
 sg13g2_buf_1 _14647_ (.A(_01064_),
    .X(_05679_));
 sg13g2_o21ai_1 _14648_ (.B1(net334),
    .Y(_05680_),
    .A1(net80),
    .A2(_05187_));
 sg13g2_a21oi_1 _14649_ (.A1(_05187_),
    .A2(_05675_),
    .Y(_00292_),
    .B1(_05680_));
 sg13g2_buf_1 _14650_ (.A(_00241_),
    .X(_05681_));
 sg13g2_inv_1 _14651_ (.Y(_05682_),
    .A(_05681_));
 sg13g2_nor2_1 _14652_ (.A(net1017),
    .B(_05682_),
    .Y(_05683_));
 sg13g2_buf_1 _14653_ (.A(\grid.cell_11_0.se ),
    .X(_05684_));
 sg13g2_buf_1 _14654_ (.A(_05684_),
    .X(_05685_));
 sg13g2_xor2_1 _14655_ (.B(net986),
    .A(_05226_),
    .X(_05686_));
 sg13g2_buf_2 _14656_ (.A(\grid.cell_11_0.sw ),
    .X(_05687_));
 sg13g2_xnor2_1 _14657_ (.Y(_05688_),
    .A(_05687_),
    .B(_05191_));
 sg13g2_xnor2_1 _14658_ (.Y(_05689_),
    .A(_05195_),
    .B(_05688_));
 sg13g2_xor2_1 _14659_ (.B(_05689_),
    .A(_05686_),
    .X(_05690_));
 sg13g2_xnor2_1 _14660_ (.Y(_05691_),
    .A(_05241_),
    .B(_05690_));
 sg13g2_nor2b_1 _14661_ (.A(net1011),
    .B_N(_05690_),
    .Y(_05692_));
 sg13g2_buf_1 _14662_ (.A(_05681_),
    .X(_05693_));
 sg13g2_nor2_1 _14663_ (.A(net671),
    .B(_05693_),
    .Y(_05694_));
 sg13g2_nor2_1 _14664_ (.A(_05692_),
    .B(_05694_),
    .Y(_05695_));
 sg13g2_o21ai_1 _14665_ (.B1(_05695_),
    .Y(_05696_),
    .A1(_05683_),
    .A2(_05691_));
 sg13g2_buf_1 _14666_ (.A(_05685_),
    .X(_05697_));
 sg13g2_buf_1 _14667_ (.A(_05697_),
    .X(_05698_));
 sg13g2_buf_1 _14668_ (.A(_05687_),
    .X(_05699_));
 sg13g2_buf_1 _14669_ (.A(net984),
    .X(_05700_));
 sg13g2_nor2_1 _14670_ (.A(net647),
    .B(net681),
    .Y(_05701_));
 sg13g2_nand2_1 _14671_ (.Y(_05702_),
    .A(net680),
    .B(_05701_));
 sg13g2_buf_1 _14672_ (.A(_00246_),
    .X(_05703_));
 sg13g2_buf_1 _14673_ (.A(_05703_),
    .X(_05704_));
 sg13g2_and2_1 _14674_ (.A(net984),
    .B(net1015),
    .X(_05705_));
 sg13g2_buf_1 _14675_ (.A(_05705_),
    .X(_05706_));
 sg13g2_nand3_1 _14676_ (.B(net983),
    .C(_05706_),
    .A(net648),
    .Y(_05707_));
 sg13g2_o21ai_1 _14677_ (.B1(_05707_),
    .Y(_05708_),
    .A1(net333),
    .A2(_05702_));
 sg13g2_buf_1 _14678_ (.A(net647),
    .X(_05709_));
 sg13g2_buf_1 _14679_ (.A(net332),
    .X(_05710_));
 sg13g2_inv_2 _14680_ (.Y(_05711_),
    .A(_05703_));
 sg13g2_nand2_1 _14681_ (.Y(_05712_),
    .A(net335),
    .B(_05711_));
 sg13g2_nor2_1 _14682_ (.A(net332),
    .B(net679),
    .Y(_05713_));
 sg13g2_a21oi_1 _14683_ (.A1(net161),
    .A2(_05712_),
    .Y(_05714_),
    .B1(_05713_));
 sg13g2_inv_2 _14684_ (.Y(_05715_),
    .A(net647));
 sg13g2_mux2_1 _14685_ (.A0(net679),
    .A1(net680),
    .S(_05715_),
    .X(_05716_));
 sg13g2_a22oi_1 _14686_ (.Y(_05717_),
    .B1(_05716_),
    .B2(net352),
    .A2(_05701_),
    .A1(_05711_));
 sg13g2_o21ai_1 _14687_ (.B1(_05717_),
    .Y(_05718_),
    .A1(net338),
    .A2(_05714_));
 sg13g2_mux2_1 _14688_ (.A0(net678),
    .A1(_05711_),
    .S(net679),
    .X(_05719_));
 sg13g2_nand2b_1 _14689_ (.Y(_05720_),
    .B(net1014),
    .A_N(_05226_));
 sg13g2_or2_1 _14690_ (.X(_05721_),
    .B(_05720_),
    .A(_05701_));
 sg13g2_o21ai_1 _14691_ (.B1(_05721_),
    .Y(_05722_),
    .A1(net161),
    .A2(_05712_));
 sg13g2_a21oi_1 _14692_ (.A1(_05710_),
    .A2(_05719_),
    .Y(_05723_),
    .B1(_05722_));
 sg13g2_nor2_1 _14693_ (.A(net333),
    .B(_05723_),
    .Y(_05724_));
 sg13g2_a221oi_1 _14694_ (.B2(net333),
    .C1(_05724_),
    .B1(_05718_),
    .A1(net662),
    .Y(_05725_),
    .A2(_05708_));
 sg13g2_xnor2_1 _14695_ (.Y(_05726_),
    .A(_05696_),
    .B(_05725_));
 sg13g2_nor2_1 _14696_ (.A(net352),
    .B(_05688_),
    .Y(_05727_));
 sg13g2_nand2_1 _14697_ (.Y(_05728_),
    .A(net647),
    .B(net681));
 sg13g2_nor2_1 _14698_ (.A(net662),
    .B(_05728_),
    .Y(_05729_));
 sg13g2_o21ai_1 _14699_ (.B1(net338),
    .Y(_05730_),
    .A1(_05727_),
    .A2(_05729_));
 sg13g2_o21ai_1 _14700_ (.B1(_05730_),
    .Y(_05731_),
    .A1(_05715_),
    .A2(_05712_));
 sg13g2_xor2_1 _14701_ (.B(net1008),
    .A(_05172_),
    .X(_05732_));
 sg13g2_nor2_1 _14702_ (.A(_05693_),
    .B(_05732_),
    .Y(_05733_));
 sg13g2_nand2b_1 _14703_ (.Y(_05734_),
    .B(_05699_),
    .A_N(net986));
 sg13g2_nor3_1 _14704_ (.A(net352),
    .B(_05208_),
    .C(_05734_),
    .Y(_05735_));
 sg13g2_a221oi_1 _14705_ (.B2(_05692_),
    .C1(_05735_),
    .B1(_05733_),
    .A1(net333),
    .Y(_05736_),
    .A2(_05731_));
 sg13g2_buf_1 _14706_ (.A(net115),
    .X(_05737_));
 sg13g2_a21oi_1 _14707_ (.A1(_05726_),
    .A2(_05736_),
    .Y(_05738_),
    .B1(net79));
 sg13g2_buf_1 _14708_ (.A(net167),
    .X(_05739_));
 sg13g2_buf_1 _14709_ (.A(\grid.cell_11_0.s ),
    .X(_05740_));
 sg13g2_buf_1 _14710_ (.A(net1174),
    .X(_05741_));
 sg13g2_xnor2_1 _14711_ (.Y(_05742_),
    .A(net982),
    .B(_05732_));
 sg13g2_xnor2_1 _14712_ (.Y(_05743_),
    .A(_05690_),
    .B(_05742_));
 sg13g2_a21oi_1 _14713_ (.A1(net112),
    .A2(_05743_),
    .Y(_05744_),
    .B1(net353));
 sg13g2_nor2b_1 _14714_ (.A(_01482_),
    .B_N(_01568_),
    .Y(_05745_));
 sg13g2_and3_1 _14715_ (.X(_05746_),
    .A(net1188),
    .B(net1053),
    .C(net1187));
 sg13g2_a21o_1 _14716_ (.A2(_05745_),
    .A1(net2),
    .B1(_05746_),
    .X(_05747_));
 sg13g2_buf_2 _14717_ (.A(_05747_),
    .X(_05748_));
 sg13g2_nand2_1 _14718_ (.Y(_05749_),
    .A(net177),
    .B(_05748_));
 sg13g2_buf_2 _14719_ (.A(_05749_),
    .X(_05750_));
 sg13g2_o21ai_1 _14720_ (.B1(net1194),
    .Y(_05751_),
    .A1(_05182_),
    .A2(_05750_));
 sg13g2_buf_1 _14721_ (.A(_05751_),
    .X(_05752_));
 sg13g2_or2_1 _14722_ (.X(_05753_),
    .B(_05752_),
    .A(_05744_));
 sg13g2_nor2_1 _14723_ (.A(_05182_),
    .B(_05750_),
    .Y(_05754_));
 sg13g2_buf_2 _14724_ (.A(_05754_),
    .X(_05755_));
 sg13g2_nand2_2 _14725_ (.Y(_05756_),
    .A(net1060),
    .B(_05755_));
 sg13g2_buf_1 _14726_ (.A(_01806_),
    .X(_05757_));
 sg13g2_nand2b_1 _14727_ (.Y(_05758_),
    .B(net44),
    .A_N(_05756_));
 sg13g2_o21ai_1 _14728_ (.B1(_05758_),
    .Y(_00293_),
    .A1(_05738_),
    .A2(_05753_));
 sg13g2_buf_1 _14729_ (.A(\grid.cell_11_1.se ),
    .X(_05759_));
 sg13g2_buf_1 _14730_ (.A(_05759_),
    .X(_05760_));
 sg13g2_nor2_1 _14731_ (.A(net663),
    .B(net981),
    .Y(_05761_));
 sg13g2_nand2b_1 _14732_ (.Y(_05762_),
    .B(_05761_),
    .A_N(net648));
 sg13g2_buf_1 _14733_ (.A(net981),
    .X(_05763_));
 sg13g2_buf_1 _14734_ (.A(net646),
    .X(_05764_));
 sg13g2_nand4_1 _14735_ (.B(net661),
    .C(net346),
    .A(net648),
    .Y(_05765_),
    .D(net331));
 sg13g2_a21oi_1 _14736_ (.A1(_05762_),
    .A2(_05765_),
    .Y(_05766_),
    .B1(net662));
 sg13g2_buf_1 _14737_ (.A(net331),
    .X(_05767_));
 sg13g2_nor4_1 _14738_ (.A(net661),
    .B(_05387_),
    .C(_05767_),
    .D(_05711_),
    .Y(_05768_));
 sg13g2_nand2b_1 _14739_ (.Y(_05769_),
    .B(net646),
    .A_N(_05703_));
 sg13g2_nor2_1 _14740_ (.A(net646),
    .B(_05711_),
    .Y(_05770_));
 sg13g2_a21o_1 _14741_ (.A2(_05769_),
    .A1(_05297_),
    .B1(_05770_),
    .X(_05771_));
 sg13g2_nand2_1 _14742_ (.Y(_05772_),
    .A(net646),
    .B(net983));
 sg13g2_o21ai_1 _14743_ (.B1(net663),
    .Y(_05773_),
    .A1(net646),
    .A2(net983));
 sg13g2_nand2_1 _14744_ (.Y(_05774_),
    .A(_05226_),
    .B(net1004));
 sg13g2_a21oi_1 _14745_ (.A1(_05772_),
    .A2(_05773_),
    .Y(_05775_),
    .B1(_05774_));
 sg13g2_a21oi_1 _14746_ (.A1(net345),
    .A2(_05771_),
    .Y(_05776_),
    .B1(_05775_));
 sg13g2_o21ai_1 _14747_ (.B1(_05769_),
    .Y(_05777_),
    .A1(_05763_),
    .A2(_05774_));
 sg13g2_nor2_1 _14748_ (.A(_05763_),
    .B(net983),
    .Y(_05778_));
 sg13g2_nor3_1 _14749_ (.A(net663),
    .B(_05774_),
    .C(_05778_),
    .Y(_05779_));
 sg13g2_a21oi_1 _14750_ (.A1(_05386_),
    .A2(_05777_),
    .Y(_05780_),
    .B1(_05779_));
 sg13g2_buf_1 _14751_ (.A(_05697_),
    .X(_05781_));
 sg13g2_nand2b_1 _14752_ (.Y(_05782_),
    .B(_05781_),
    .A_N(_05780_));
 sg13g2_o21ai_1 _14753_ (.B1(_05782_),
    .Y(_05783_),
    .A1(_05698_),
    .A2(_05776_));
 sg13g2_nor3_1 _14754_ (.A(_05766_),
    .B(_05768_),
    .C(_05783_),
    .Y(_05784_));
 sg13g2_xnor2_1 _14755_ (.Y(_05785_),
    .A(net981),
    .B(_05286_));
 sg13g2_xor2_1 _14756_ (.B(_05785_),
    .A(_05686_),
    .X(_05786_));
 sg13g2_xnor2_1 _14757_ (.Y(_05787_),
    .A(net353),
    .B(_05786_));
 sg13g2_inv_1 _14758_ (.Y(_05788_),
    .A(_00244_));
 sg13g2_and2_1 _14759_ (.A(_05788_),
    .B(_05786_),
    .X(_05789_));
 sg13g2_nor2_1 _14760_ (.A(_05694_),
    .B(_05789_),
    .Y(_05790_));
 sg13g2_o21ai_1 _14761_ (.B1(_05790_),
    .Y(_05791_),
    .A1(_05683_),
    .A2(_05787_));
 sg13g2_xnor2_1 _14762_ (.Y(_05792_),
    .A(_05784_),
    .B(_05791_));
 sg13g2_xnor2_1 _14763_ (.Y(_05793_),
    .A(_05172_),
    .B(net1012));
 sg13g2_xnor2_1 _14764_ (.Y(_05794_),
    .A(net1174),
    .B(_05793_));
 sg13g2_xor2_1 _14765_ (.B(_05794_),
    .A(_05786_),
    .X(_05795_));
 sg13g2_nand2_1 _14766_ (.Y(_05796_),
    .A(_05386_),
    .B(net331));
 sg13g2_xnor2_1 _14767_ (.Y(_05797_),
    .A(_05285_),
    .B(_05759_));
 sg13g2_nor2_1 _14768_ (.A(_05238_),
    .B(_05797_),
    .Y(_05798_));
 sg13g2_nor2_1 _14769_ (.A(net1009),
    .B(_05796_),
    .Y(_05799_));
 sg13g2_o21ai_1 _14770_ (.B1(net661),
    .Y(_05800_),
    .A1(_05798_),
    .A2(_05799_));
 sg13g2_o21ai_1 _14771_ (.B1(_05800_),
    .Y(_05801_),
    .A1(net983),
    .A2(_05796_));
 sg13g2_and2_1 _14772_ (.A(_05682_),
    .B(_05793_),
    .X(_05802_));
 sg13g2_nor3_1 _14773_ (.A(_05781_),
    .B(_05796_),
    .C(_05774_),
    .Y(_05803_));
 sg13g2_nand2b_1 _14774_ (.Y(_05804_),
    .B(net171),
    .A_N(_05803_));
 sg13g2_a221oi_1 _14775_ (.B2(_05789_),
    .C1(_05804_),
    .B1(_05802_),
    .A1(net333),
    .Y(_05805_),
    .A2(_05801_));
 sg13g2_o21ai_1 _14776_ (.B1(_05805_),
    .Y(_05806_),
    .A1(_05241_),
    .A2(_05795_));
 sg13g2_a21oi_1 _14777_ (.A1(net673),
    .A2(net115),
    .Y(_05807_),
    .B1(_05755_));
 sg13g2_o21ai_1 _14778_ (.B1(_05807_),
    .Y(_05808_),
    .A1(_05792_),
    .A2(_05806_));
 sg13g2_nand2b_1 _14779_ (.Y(_05809_),
    .B(_05755_),
    .A_N(_03153_));
 sg13g2_and3_1 _14780_ (.X(_00294_),
    .A(_12999_),
    .B(_05808_),
    .C(_05809_));
 sg13g2_nand2_1 _14781_ (.Y(_05810_),
    .A(_03884_),
    .B(_04046_));
 sg13g2_buf_2 _14782_ (.A(_05810_),
    .X(_05811_));
 sg13g2_buf_1 _14783_ (.A(_05811_),
    .X(_05812_));
 sg13g2_nand2_1 _14784_ (.Y(_05813_),
    .A(net33),
    .B(_05755_));
 sg13g2_buf_1 _14785_ (.A(net167),
    .X(_05814_));
 sg13g2_buf_1 _14786_ (.A(_05814_),
    .X(_05815_));
 sg13g2_xnor2_1 _14787_ (.Y(_05816_),
    .A(_05284_),
    .B(_05759_));
 sg13g2_buf_2 _14788_ (.A(\grid.cell_11_2.se ),
    .X(_05817_));
 sg13g2_xnor2_1 _14789_ (.Y(_05818_),
    .A(_05817_),
    .B(_05358_));
 sg13g2_buf_1 _14790_ (.A(_05818_),
    .X(_05819_));
 sg13g2_xnor2_1 _14791_ (.Y(_05820_),
    .A(_05361_),
    .B(_05819_));
 sg13g2_xnor2_1 _14792_ (.Y(_05821_),
    .A(_05816_),
    .B(_05820_));
 sg13g2_nand2b_1 _14793_ (.Y(_05822_),
    .B(_05821_),
    .A_N(net1011));
 sg13g2_buf_1 _14794_ (.A(_00240_),
    .X(_05823_));
 sg13g2_xnor2_1 _14795_ (.Y(_05824_),
    .A(_05228_),
    .B(_05817_));
 sg13g2_xnor2_1 _14796_ (.Y(_05825_),
    .A(_05816_),
    .B(_05824_));
 sg13g2_xnor2_1 _14797_ (.Y(_05826_),
    .A(_05383_),
    .B(_05825_));
 sg13g2_buf_1 _14798_ (.A(_05826_),
    .X(_05827_));
 sg13g2_nor2_1 _14799_ (.A(_05823_),
    .B(_05827_),
    .Y(_05828_));
 sg13g2_buf_1 _14800_ (.A(_05823_),
    .X(_05829_));
 sg13g2_nor2b_1 _14801_ (.A(net1011),
    .B_N(_05821_),
    .Y(_05830_));
 sg13g2_o21ai_1 _14802_ (.B1(_05827_),
    .Y(_05831_),
    .A1(_05829_),
    .A2(_05830_));
 sg13g2_a21oi_1 _14803_ (.A1(net352),
    .A2(_05827_),
    .Y(_05832_),
    .B1(_05829_));
 sg13g2_nor2_1 _14804_ (.A(_05822_),
    .B(_05832_),
    .Y(_05833_));
 sg13g2_a221oi_1 _14805_ (.B2(net662),
    .C1(_05833_),
    .B1(_05831_),
    .A1(_05822_),
    .Y(_05834_),
    .A2(_05828_));
 sg13g2_nor2_1 _14806_ (.A(_05321_),
    .B(_05819_),
    .Y(_05835_));
 sg13g2_buf_1 _14807_ (.A(_05817_),
    .X(_05836_));
 sg13g2_nand2_1 _14808_ (.Y(_05837_),
    .A(net979),
    .B(_05359_));
 sg13g2_nor2_1 _14809_ (.A(net1004),
    .B(_05837_),
    .Y(_05838_));
 sg13g2_or2_1 _14810_ (.X(_05839_),
    .B(_05838_),
    .A(_05835_));
 sg13g2_nor2_1 _14811_ (.A(net1176),
    .B(_05837_),
    .Y(_05840_));
 sg13g2_a21oi_1 _14812_ (.A1(net666),
    .A2(_05839_),
    .Y(_05841_),
    .B1(_05840_));
 sg13g2_nand2_1 _14813_ (.Y(_05842_),
    .A(_05307_),
    .B(net1000));
 sg13g2_or2_1 _14814_ (.X(_05843_),
    .B(_05837_),
    .A(_05842_));
 sg13g2_inv_2 _14815_ (.Y(_05844_),
    .A(_05759_));
 sg13g2_mux2_1 _14816_ (.A0(_05841_),
    .A1(_05843_),
    .S(_05844_),
    .X(_05845_));
 sg13g2_nand2_1 _14817_ (.Y(_05846_),
    .A(net980),
    .B(_05827_));
 sg13g2_o21ai_1 _14818_ (.B1(_05846_),
    .Y(_05847_),
    .A1(net662),
    .A2(_05828_));
 sg13g2_nand3_1 _14819_ (.B(_05845_),
    .C(_05847_),
    .A(_05822_),
    .Y(_05848_));
 sg13g2_buf_1 _14820_ (.A(net979),
    .X(_05849_));
 sg13g2_a21oi_1 _14821_ (.A1(net661),
    .A2(net331),
    .Y(_05850_),
    .B1(_05391_));
 sg13g2_nor4_1 _14822_ (.A(_05849_),
    .B(_05360_),
    .C(_05334_),
    .D(_05850_),
    .Y(_05851_));
 sg13g2_nor2_1 _14823_ (.A(net645),
    .B(net1001),
    .Y(_05852_));
 sg13g2_nand2_1 _14824_ (.Y(_05853_),
    .A(_05852_),
    .B(_05842_));
 sg13g2_a21oi_1 _14825_ (.A1(_05849_),
    .A2(_05359_),
    .Y(_05854_),
    .B1(net1000));
 sg13g2_o21ai_1 _14826_ (.B1(net1176),
    .Y(_05855_),
    .A1(_05835_),
    .A2(_05854_));
 sg13g2_a21oi_1 _14827_ (.A1(_05853_),
    .A2(_05855_),
    .Y(_05856_),
    .B1(_05767_));
 sg13g2_nor2_1 _14828_ (.A(_05851_),
    .B(_05856_),
    .Y(_05857_));
 sg13g2_mux2_1 _14829_ (.A0(_05834_),
    .A1(_05848_),
    .S(_05857_),
    .X(_05858_));
 sg13g2_xnor2_1 _14830_ (.Y(_05859_),
    .A(_05686_),
    .B(_05827_));
 sg13g2_a21oi_1 _14831_ (.A1(net167),
    .A2(_05859_),
    .Y(_05860_),
    .B1(net346));
 sg13g2_or2_1 _14832_ (.X(_05861_),
    .B(_05860_),
    .A(_05755_));
 sg13g2_a21o_1 _14833_ (.A2(_05858_),
    .A1(net78),
    .B1(_05861_),
    .X(_05862_));
 sg13g2_a21oi_1 _14834_ (.A1(_05813_),
    .A2(_05862_),
    .Y(_00295_),
    .B1(_05283_));
 sg13g2_buf_1 _14835_ (.A(net48),
    .X(_05863_));
 sg13g2_buf_1 _14836_ (.A(\grid.cell_11_3.se ),
    .X(_05864_));
 sg13g2_buf_1 _14837_ (.A(net1172),
    .X(_05865_));
 sg13g2_buf_1 _14838_ (.A(net978),
    .X(_05866_));
 sg13g2_nand2_1 _14839_ (.Y(_05867_),
    .A(net979),
    .B(net998));
 sg13g2_nand2_1 _14840_ (.Y(_05868_),
    .A(net998),
    .B(net1000));
 sg13g2_nand2_1 _14841_ (.Y(_05869_),
    .A(net979),
    .B(_05514_));
 sg13g2_o21ai_1 _14842_ (.B1(_05869_),
    .Y(_05870_),
    .A1(net645),
    .A2(_05868_));
 sg13g2_nand2_1 _14843_ (.Y(_05871_),
    .A(net658),
    .B(_05870_));
 sg13g2_o21ai_1 _14844_ (.B1(_05871_),
    .Y(_05872_),
    .A1(_05379_),
    .A2(_05867_));
 sg13g2_xnor2_1 _14845_ (.Y(_05873_),
    .A(net1172),
    .B(_05421_));
 sg13g2_xnor2_1 _14846_ (.Y(_05874_),
    .A(_05817_),
    .B(_05361_));
 sg13g2_xnor2_1 _14847_ (.Y(_05875_),
    .A(_05873_),
    .B(_05874_));
 sg13g2_and2_1 _14848_ (.A(_05381_),
    .B(_05875_),
    .X(_05876_));
 sg13g2_buf_1 _14849_ (.A(_00239_),
    .X(_05877_));
 sg13g2_nor2b_1 _14850_ (.A(_05877_),
    .B_N(_05286_),
    .Y(_05878_));
 sg13g2_nand2_1 _14851_ (.Y(_05879_),
    .A(net658),
    .B(net666));
 sg13g2_nor3_1 _14852_ (.A(_05866_),
    .B(_05867_),
    .C(_05879_),
    .Y(_05880_));
 sg13g2_a221oi_1 _14853_ (.B2(_05878_),
    .C1(_05880_),
    .B1(_05876_),
    .A1(net644),
    .Y(_05881_),
    .A2(_05872_));
 sg13g2_nor3_1 _14854_ (.A(net978),
    .B(net645),
    .C(net660),
    .Y(_05882_));
 sg13g2_buf_1 _14855_ (.A(net1172),
    .X(_05883_));
 sg13g2_nor3_1 _14856_ (.A(net977),
    .B(_05836_),
    .C(_05457_),
    .Y(_05884_));
 sg13g2_o21ai_1 _14857_ (.B1(_05867_),
    .Y(_05885_),
    .A1(_05445_),
    .A2(net1000));
 sg13g2_nand2_1 _14858_ (.Y(_05886_),
    .A(_05864_),
    .B(net998));
 sg13g2_nand2_1 _14859_ (.Y(_05887_),
    .A(net977),
    .B(_05836_));
 sg13g2_nand3_1 _14860_ (.B(_05886_),
    .C(_05887_),
    .A(_05379_),
    .Y(_05888_));
 sg13g2_nor3_1 _14861_ (.A(_05884_),
    .B(_05885_),
    .C(_05888_),
    .Y(_05889_));
 sg13g2_a21o_1 _14862_ (.A2(_05882_),
    .A1(_05879_),
    .B1(_05889_),
    .X(_05890_));
 sg13g2_nand2_1 _14863_ (.Y(_05891_),
    .A(net345),
    .B(_05877_));
 sg13g2_xnor2_1 _14864_ (.Y(_05892_),
    .A(net670),
    .B(_05875_));
 sg13g2_nor2_1 _14865_ (.A(net345),
    .B(_05877_),
    .Y(_05893_));
 sg13g2_a221oi_1 _14866_ (.B2(_05892_),
    .C1(_05893_),
    .B1(_05891_),
    .A1(_05381_),
    .Y(_05894_),
    .A2(_05875_));
 sg13g2_xor2_1 _14867_ (.B(_05894_),
    .A(_05890_),
    .X(_05895_));
 sg13g2_a21oi_1 _14868_ (.A1(_05881_),
    .A2(_05895_),
    .Y(_05896_),
    .B1(net124));
 sg13g2_buf_1 _14869_ (.A(net123),
    .X(_05897_));
 sg13g2_xor2_1 _14870_ (.B(_05875_),
    .A(_05785_),
    .X(_05898_));
 sg13g2_a21oi_1 _14871_ (.A1(net77),
    .A2(_05898_),
    .Y(_05899_),
    .B1(net667));
 sg13g2_or3_1 _14872_ (.A(_05752_),
    .B(_05896_),
    .C(_05899_),
    .X(_05900_));
 sg13g2_o21ai_1 _14873_ (.B1(_05900_),
    .Y(_00296_),
    .A1(_05863_),
    .A2(_05756_));
 sg13g2_buf_2 _14874_ (.A(\grid.cell_11_4.se ),
    .X(_05901_));
 sg13g2_buf_1 _14875_ (.A(_05901_),
    .X(_05902_));
 sg13g2_buf_1 _14876_ (.A(net976),
    .X(_05903_));
 sg13g2_buf_1 _14877_ (.A(net643),
    .X(_05904_));
 sg13g2_nand2_1 _14878_ (.Y(_05905_),
    .A(net977),
    .B(net656));
 sg13g2_nor2_1 _14879_ (.A(_05434_),
    .B(_05905_),
    .Y(_05906_));
 sg13g2_xnor2_1 _14880_ (.Y(_05907_),
    .A(net656),
    .B(net997));
 sg13g2_o21ai_1 _14881_ (.B1(net655),
    .Y(_05908_),
    .A1(net977),
    .A2(_05552_));
 sg13g2_a21oi_1 _14882_ (.A1(net978),
    .A2(_05907_),
    .Y(_05909_),
    .B1(_05908_));
 sg13g2_or2_1 _14883_ (.X(_05910_),
    .B(_05909_),
    .A(_05906_));
 sg13g2_xnor2_1 _14884_ (.Y(_05911_),
    .A(_05901_),
    .B(_05475_));
 sg13g2_xnor2_1 _14885_ (.Y(_05912_),
    .A(net994),
    .B(_05911_));
 sg13g2_xnor2_1 _14886_ (.Y(_05913_),
    .A(net1172),
    .B(_05420_));
 sg13g2_xnor2_1 _14887_ (.Y(_05914_),
    .A(_05912_),
    .B(_05913_));
 sg13g2_and2_1 _14888_ (.A(_05417_),
    .B(_05914_),
    .X(_05915_));
 sg13g2_buf_2 _14889_ (.A(_00045_),
    .X(_05916_));
 sg13g2_nor2b_1 _14890_ (.A(_05916_),
    .B_N(_05383_),
    .Y(_05917_));
 sg13g2_nand2_1 _14891_ (.Y(_05918_),
    .A(net655),
    .B(net658));
 sg13g2_nor3_1 _14892_ (.A(net329),
    .B(_05905_),
    .C(_05918_),
    .Y(_05919_));
 sg13g2_a221oi_1 _14893_ (.B2(_05917_),
    .C1(_05919_),
    .B1(_05915_),
    .A1(net329),
    .Y(_05920_),
    .A2(_05910_));
 sg13g2_nor4_1 _14894_ (.A(net976),
    .B(net977),
    .C(net656),
    .D(_05604_),
    .Y(_05921_));
 sg13g2_a221oi_1 _14895_ (.B2(_05445_),
    .C1(_05921_),
    .B1(net655),
    .A1(net978),
    .Y(_05922_),
    .A2(net656));
 sg13g2_o21ai_1 _14896_ (.B1(_05903_),
    .Y(_05923_),
    .A1(_05883_),
    .A2(net656));
 sg13g2_and2_1 _14897_ (.A(_05434_),
    .B(_05923_),
    .X(_05924_));
 sg13g2_nor3_1 _14898_ (.A(_05904_),
    .B(net978),
    .C(net344),
    .Y(_05925_));
 sg13g2_a22oi_1 _14899_ (.Y(_05926_),
    .B1(_05925_),
    .B2(_05918_),
    .A2(_05924_),
    .A1(_05922_));
 sg13g2_nand2_1 _14900_ (.Y(_05927_),
    .A(_05916_),
    .B(_05391_));
 sg13g2_xnor2_1 _14901_ (.Y(_05928_),
    .A(net664),
    .B(_05914_));
 sg13g2_nor2_1 _14902_ (.A(_05916_),
    .B(_05391_),
    .Y(_05929_));
 sg13g2_a221oi_1 _14903_ (.B2(_05928_),
    .C1(_05929_),
    .B1(_05927_),
    .A1(_05417_),
    .Y(_05930_),
    .A2(_05914_));
 sg13g2_xnor2_1 _14904_ (.Y(_05931_),
    .A(_05926_),
    .B(_05930_));
 sg13g2_a21oi_1 _14905_ (.A1(_05920_),
    .A2(_05931_),
    .Y(_05932_),
    .B1(net124));
 sg13g2_xor2_1 _14906_ (.B(_05914_),
    .A(_05820_),
    .X(_05933_));
 sg13g2_a21oi_1 _14907_ (.A1(_05897_),
    .A2(_05933_),
    .Y(_05934_),
    .B1(_05436_));
 sg13g2_or3_1 _14908_ (.A(_05752_),
    .B(_05932_),
    .C(_05934_),
    .X(_05935_));
 sg13g2_o21ai_1 _14909_ (.B1(_05935_),
    .Y(_00297_),
    .A1(net34),
    .A2(_05756_));
 sg13g2_buf_1 _14910_ (.A(\grid.cell_11_5.se ),
    .X(_05936_));
 sg13g2_buf_1 _14911_ (.A(net1171),
    .X(_05937_));
 sg13g2_buf_1 _14912_ (.A(net975),
    .X(_05938_));
 sg13g2_buf_1 _14913_ (.A(net642),
    .X(_05939_));
 sg13g2_nand2_1 _14914_ (.Y(_05940_),
    .A(net976),
    .B(net992));
 sg13g2_xnor2_1 _14915_ (.Y(_05941_),
    .A(net992),
    .B(net994));
 sg13g2_a21oi_1 _14916_ (.A1(net653),
    .A2(net994),
    .Y(_05942_),
    .B1(_05902_));
 sg13g2_a21oi_1 _14917_ (.A1(_05903_),
    .A2(_05941_),
    .Y(_05943_),
    .B1(_05942_));
 sg13g2_nand2_1 _14918_ (.Y(_05944_),
    .A(net340),
    .B(_05943_));
 sg13g2_o21ai_1 _14919_ (.B1(_05944_),
    .Y(_05945_),
    .A1(_05488_),
    .A2(_05940_));
 sg13g2_inv_1 _14920_ (.Y(_05946_),
    .A(_05484_));
 sg13g2_xnor2_1 _14921_ (.Y(_05947_),
    .A(net1171),
    .B(_05901_));
 sg13g2_xnor2_1 _14922_ (.Y(_05948_),
    .A(_05547_),
    .B(_05947_));
 sg13g2_xnor2_1 _14923_ (.Y(_05949_),
    .A(net994),
    .B(_05948_));
 sg13g2_and2_1 _14924_ (.A(_05946_),
    .B(_05949_),
    .X(_05950_));
 sg13g2_buf_1 _14925_ (.A(_00077_),
    .X(_05951_));
 sg13g2_inv_2 _14926_ (.Y(_05952_),
    .A(_05951_));
 sg13g2_and2_1 _14927_ (.A(_05952_),
    .B(_05421_),
    .X(_05953_));
 sg13g2_nand2_1 _14928_ (.Y(_05954_),
    .A(net340),
    .B(net655));
 sg13g2_nor3_1 _14929_ (.A(_05939_),
    .B(_05940_),
    .C(_05954_),
    .Y(_05955_));
 sg13g2_a221oi_1 _14930_ (.B2(_05953_),
    .C1(_05955_),
    .B1(_05950_),
    .A1(net328),
    .Y(_05956_),
    .A2(_05945_));
 sg13g2_buf_1 _14931_ (.A(net975),
    .X(_05957_));
 sg13g2_nor4_1 _14932_ (.A(net641),
    .B(_05902_),
    .C(net653),
    .D(net649),
    .Y(_05958_));
 sg13g2_nand2_1 _14933_ (.Y(_05959_),
    .A(net641),
    .B(net992));
 sg13g2_nand2_1 _14934_ (.Y(_05960_),
    .A(_05940_),
    .B(_05959_));
 sg13g2_nand2_1 _14935_ (.Y(_05961_),
    .A(net641),
    .B(net976));
 sg13g2_o21ai_1 _14936_ (.B1(_05961_),
    .Y(_05962_),
    .A1(net649),
    .A2(net655));
 sg13g2_nor3_1 _14937_ (.A(_05958_),
    .B(_05960_),
    .C(_05962_),
    .Y(_05963_));
 sg13g2_nor3_1 _14938_ (.A(_05938_),
    .B(_05904_),
    .C(net341),
    .Y(_05964_));
 sg13g2_a22oi_1 _14939_ (.Y(_05965_),
    .B1(_05964_),
    .B2(_05954_),
    .A2(_05963_),
    .A1(_05488_));
 sg13g2_nor2_1 _14940_ (.A(_05952_),
    .B(_05449_),
    .Y(_05966_));
 sg13g2_xnor2_1 _14941_ (.Y(_05967_),
    .A(net660),
    .B(_05949_));
 sg13g2_a22oi_1 _14942_ (.Y(_05968_),
    .B1(_05949_),
    .B2(_05946_),
    .A2(_05449_),
    .A1(_05952_));
 sg13g2_o21ai_1 _14943_ (.B1(_05968_),
    .Y(_05969_),
    .A1(_05966_),
    .A2(_05967_));
 sg13g2_xor2_1 _14944_ (.B(_05969_),
    .A(_05965_),
    .X(_05970_));
 sg13g2_a21oi_1 _14945_ (.A1(_05956_),
    .A2(_05970_),
    .Y(_05971_),
    .B1(_04624_));
 sg13g2_xor2_1 _14946_ (.B(_05949_),
    .A(_05873_),
    .X(_05972_));
 sg13g2_a21oi_1 _14947_ (.A1(_05897_),
    .A2(_05972_),
    .Y(_05973_),
    .B1(net344));
 sg13g2_or3_1 _14948_ (.A(_05752_),
    .B(_05971_),
    .C(_05973_),
    .X(_05974_));
 sg13g2_o21ai_1 _14949_ (.B1(_05974_),
    .Y(_00298_),
    .A1(net46),
    .A2(_05756_));
 sg13g2_xnor2_1 _14950_ (.Y(_05975_),
    .A(net355),
    .B(net651));
 sg13g2_a21oi_1 _14951_ (.A1(net355),
    .A2(net651),
    .Y(_05976_),
    .B1(net161));
 sg13g2_a21oi_1 _14952_ (.A1(net161),
    .A2(_05975_),
    .Y(_05977_),
    .B1(_05976_));
 sg13g2_nand2_1 _14953_ (.Y(_05978_),
    .A(net338),
    .B(_05977_));
 sg13g2_o21ai_1 _14954_ (.B1(_05978_),
    .Y(_05979_),
    .A1(net652),
    .A2(_05728_));
 sg13g2_inv_1 _14955_ (.Y(_05980_),
    .A(_05553_));
 sg13g2_xnor2_1 _14956_ (.Y(_05981_),
    .A(_05936_),
    .B(net989));
 sg13g2_xnor2_1 _14957_ (.Y(_05982_),
    .A(_05689_),
    .B(_05981_));
 sg13g2_and2_1 _14958_ (.A(_05980_),
    .B(_05982_),
    .X(_05983_));
 sg13g2_buf_1 _14959_ (.A(_00109_),
    .X(_05984_));
 sg13g2_buf_1 _14960_ (.A(_05984_),
    .X(_05985_));
 sg13g2_xor2_1 _14961_ (.B(_05507_),
    .A(net344),
    .X(_05986_));
 sg13g2_nor2_1 _14962_ (.A(net974),
    .B(_05986_),
    .Y(_05987_));
 sg13g2_nand2_1 _14963_ (.Y(_05988_),
    .A(net989),
    .B(_05195_));
 sg13g2_buf_2 _14964_ (.A(_05988_),
    .X(_05989_));
 sg13g2_nor3_1 _14965_ (.A(net328),
    .B(_05728_),
    .C(_05989_),
    .Y(_05990_));
 sg13g2_a221oi_1 _14966_ (.B2(_05987_),
    .C1(_05990_),
    .B1(_05983_),
    .A1(net328),
    .Y(_05991_),
    .A2(_05979_));
 sg13g2_nor3_1 _14967_ (.A(net641),
    .B(net332),
    .C(net335),
    .Y(_05992_));
 sg13g2_nor2_1 _14968_ (.A(net642),
    .B(_05706_),
    .Y(_05993_));
 sg13g2_o21ai_1 _14969_ (.B1(net652),
    .Y(_05994_),
    .A1(_05701_),
    .A2(_05993_));
 sg13g2_nor2b_1 _14970_ (.A(_05992_),
    .B_N(_05994_),
    .Y(_05995_));
 sg13g2_nor3_1 _14971_ (.A(_05528_),
    .B(net647),
    .C(net681),
    .Y(_05996_));
 sg13g2_nor3_1 _14972_ (.A(_05706_),
    .B(_05989_),
    .C(_05996_),
    .Y(_05997_));
 sg13g2_a21o_1 _14973_ (.A2(_05706_),
    .A1(net987),
    .B1(_05997_),
    .X(_05998_));
 sg13g2_nand2_1 _14974_ (.Y(_05999_),
    .A(net987),
    .B(_05709_));
 sg13g2_nor2_1 _14975_ (.A(_05715_),
    .B(net678),
    .Y(_06000_));
 sg13g2_nor2_1 _14976_ (.A(net987),
    .B(_05957_),
    .Y(_06001_));
 sg13g2_o21ai_1 _14977_ (.B1(_06001_),
    .Y(_06002_),
    .A1(_05713_),
    .A2(_06000_));
 sg13g2_o21ai_1 _14978_ (.B1(_06002_),
    .Y(_06003_),
    .A1(_05208_),
    .A2(_05999_));
 sg13g2_and2_1 _14979_ (.A(net975),
    .B(_05700_),
    .X(_06004_));
 sg13g2_buf_1 _14980_ (.A(_06004_),
    .X(_06005_));
 sg13g2_a21oi_1 _14981_ (.A1(_05201_),
    .A2(_06005_),
    .Y(_06006_),
    .B1(_05992_));
 sg13g2_nor2_1 _14982_ (.A(net340),
    .B(_06006_),
    .Y(_06007_));
 sg13g2_a221oi_1 _14983_ (.B2(net340),
    .C1(_06007_),
    .B1(_06003_),
    .A1(net328),
    .Y(_06008_),
    .A2(_05998_));
 sg13g2_o21ai_1 _14984_ (.B1(_06008_),
    .Y(_06009_),
    .A1(net338),
    .A2(_05995_));
 sg13g2_xnor2_1 _14985_ (.Y(_06010_),
    .A(net344),
    .B(_05982_));
 sg13g2_a21oi_1 _14986_ (.A1(net974),
    .A2(_05604_),
    .Y(_06011_),
    .B1(_06010_));
 sg13g2_nor2_1 _14987_ (.A(net974),
    .B(_05604_),
    .Y(_06012_));
 sg13g2_nor3_1 _14988_ (.A(_05983_),
    .B(_06011_),
    .C(_06012_),
    .Y(_06013_));
 sg13g2_xor2_1 _14989_ (.B(_06013_),
    .A(_06009_),
    .X(_06014_));
 sg13g2_a21oi_1 _14990_ (.A1(_05991_),
    .A2(_06014_),
    .Y(_06015_),
    .B1(net79));
 sg13g2_xor2_1 _14991_ (.B(_05982_),
    .A(_05912_),
    .X(_06016_));
 sg13g2_a21oi_1 _14992_ (.A1(_04860_),
    .A2(_06016_),
    .Y(_06017_),
    .B1(net162));
 sg13g2_or2_1 _14993_ (.X(_06018_),
    .B(_06017_),
    .A(_05752_));
 sg13g2_buf_2 _14994_ (.A(net45),
    .X(_06019_));
 sg13g2_nand2b_1 _14995_ (.Y(_06020_),
    .B(_06019_),
    .A_N(_05756_));
 sg13g2_o21ai_1 _14996_ (.B1(_06020_),
    .Y(_00299_),
    .A1(_06015_),
    .A2(_06018_));
 sg13g2_nand2_1 _14997_ (.Y(_06021_),
    .A(net80),
    .B(_05755_));
 sg13g2_nand4_1 _14998_ (.B(net332),
    .C(net653),
    .A(net987),
    .Y(_06022_),
    .D(net680));
 sg13g2_nor2b_1 _14999_ (.A(net332),
    .B_N(net653),
    .Y(_06023_));
 sg13g2_o21ai_1 _15000_ (.B1(_06001_),
    .Y(_06024_),
    .A1(_06000_),
    .A2(_06023_));
 sg13g2_nand3_1 _15001_ (.B(_06022_),
    .C(_06024_),
    .A(net340),
    .Y(_06025_));
 sg13g2_nor2_1 _15002_ (.A(net332),
    .B(net992),
    .Y(_06026_));
 sg13g2_nand2b_1 _15003_ (.Y(_06027_),
    .B(_06026_),
    .A_N(net642));
 sg13g2_nand3_1 _15004_ (.B(net680),
    .C(_06005_),
    .A(_05526_),
    .Y(_06028_));
 sg13g2_nand3_1 _15005_ (.B(_06027_),
    .C(_06028_),
    .A(_05634_),
    .Y(_06029_));
 sg13g2_and2_1 _15006_ (.A(net984),
    .B(_05523_),
    .X(_06030_));
 sg13g2_buf_1 _15007_ (.A(_06030_),
    .X(_06031_));
 sg13g2_nor3_1 _15008_ (.A(net991),
    .B(net332),
    .C(net653),
    .Y(_06032_));
 sg13g2_nor3_1 _15009_ (.A(_05989_),
    .B(_06031_),
    .C(_06032_),
    .Y(_06033_));
 sg13g2_a21o_1 _15010_ (.A2(_06031_),
    .A1(net987),
    .B1(_06033_),
    .X(_06034_));
 sg13g2_nor2_1 _15011_ (.A(net642),
    .B(_06031_),
    .Y(_06035_));
 sg13g2_o21ai_1 _15012_ (.B1(net652),
    .Y(_06036_),
    .A1(_06026_),
    .A2(_06035_));
 sg13g2_a21oi_1 _15013_ (.A1(_06027_),
    .A2(_06036_),
    .Y(_06037_),
    .B1(net338));
 sg13g2_a221oi_1 _15014_ (.B2(_05939_),
    .C1(_06037_),
    .B1(_06034_),
    .A1(_06025_),
    .Y(_06038_),
    .A2(_06029_));
 sg13g2_xnor2_1 _15015_ (.Y(_06039_),
    .A(net1171),
    .B(_05687_));
 sg13g2_xnor2_1 _15016_ (.Y(_06040_),
    .A(_05547_),
    .B(_06039_));
 sg13g2_xnor2_1 _15017_ (.Y(_06041_),
    .A(_05195_),
    .B(_06040_));
 sg13g2_xnor2_1 _15018_ (.Y(_06042_),
    .A(_05247_),
    .B(_06041_));
 sg13g2_a22oi_1 _15019_ (.Y(_06043_),
    .B1(_06042_),
    .B2(net1017),
    .A2(_06041_),
    .A1(_05788_));
 sg13g2_xnor2_1 _15020_ (.Y(_06044_),
    .A(_05793_),
    .B(_06041_));
 sg13g2_nand2_1 _15021_ (.Y(_06045_),
    .A(_05682_),
    .B(_06044_));
 sg13g2_and2_1 _15022_ (.A(_06043_),
    .B(_06045_),
    .X(_06046_));
 sg13g2_xor2_1 _15023_ (.B(_06045_),
    .A(_06043_),
    .X(_06047_));
 sg13g2_inv_1 _15024_ (.Y(_06048_),
    .A(_05989_));
 sg13g2_nor4_1 _15025_ (.A(_05957_),
    .B(_05709_),
    .C(_05525_),
    .D(net678),
    .Y(_06049_));
 sg13g2_nor2_1 _15026_ (.A(net651),
    .B(net678),
    .Y(_06050_));
 sg13g2_nor3_1 _15027_ (.A(_06049_),
    .B(_06031_),
    .C(_06050_),
    .Y(_06051_));
 sg13g2_o21ai_1 _15028_ (.B1(_05938_),
    .Y(_06052_),
    .A1(net161),
    .A2(_05526_));
 sg13g2_nand3_1 _15029_ (.B(_06051_),
    .C(_06052_),
    .A(net652),
    .Y(_06053_));
 sg13g2_o21ai_1 _15030_ (.B1(_06053_),
    .Y(_06054_),
    .A1(_06048_),
    .A2(_06027_));
 sg13g2_buf_2 _15031_ (.A(net163),
    .X(_06055_));
 sg13g2_a221oi_1 _15032_ (.B2(_06054_),
    .C1(_06055_),
    .B1(_06047_),
    .A1(_06038_),
    .Y(_06056_),
    .A2(_06046_));
 sg13g2_buf_1 _15033_ (.A(net167),
    .X(_06057_));
 sg13g2_xor2_1 _15034_ (.B(_06041_),
    .A(_05794_),
    .X(_06058_));
 sg13g2_a21oi_1 _15035_ (.A1(net109),
    .A2(_06058_),
    .Y(_06059_),
    .B1(net355));
 sg13g2_or3_1 _15036_ (.A(_05755_),
    .B(_06056_),
    .C(_06059_),
    .X(_06060_));
 sg13g2_a21oi_1 _15037_ (.A1(_06021_),
    .A2(_06060_),
    .Y(_00300_),
    .B1(net350));
 sg13g2_nor2b_1 _15038_ (.A(net1053),
    .B_N(net3),
    .Y(_06061_));
 sg13g2_a22oi_1 _15039_ (.Y(_06062_),
    .B1(_06061_),
    .B2(net4),
    .A2(_04907_),
    .A1(net1053));
 sg13g2_buf_1 _15040_ (.A(_06062_),
    .X(_06063_));
 sg13g2_nor3_1 _15041_ (.A(_01989_),
    .B(_02021_),
    .C(net159),
    .Y(_06064_));
 sg13g2_buf_1 _15042_ (.A(_06064_),
    .X(_06065_));
 sg13g2_buf_1 _15043_ (.A(\grid.cell_12_0.se ),
    .X(_06066_));
 sg13g2_buf_1 _15044_ (.A(\grid.cell_12_0.sw ),
    .X(_06067_));
 sg13g2_xnor2_1 _15045_ (.Y(_06068_),
    .A(_06066_),
    .B(net1170));
 sg13g2_xnor2_1 _15046_ (.Y(_06069_),
    .A(_05715_),
    .B(_06068_));
 sg13g2_nand2_1 _15047_ (.Y(_06070_),
    .A(net1008),
    .B(net355));
 sg13g2_o21ai_1 _15048_ (.B1(net1011),
    .Y(_06071_),
    .A1(net1008),
    .A2(net679));
 sg13g2_nor2_1 _15049_ (.A(_06071_),
    .B(_06069_),
    .Y(_06072_));
 sg13g2_a21oi_1 _15050_ (.A1(_06069_),
    .A2(_06070_),
    .Y(_06073_),
    .B1(_06072_));
 sg13g2_buf_1 _15051_ (.A(_06066_),
    .X(_06074_));
 sg13g2_buf_1 _15052_ (.A(_06074_),
    .X(_06075_));
 sg13g2_buf_1 _15053_ (.A(_06067_),
    .X(_06076_));
 sg13g2_buf_1 _15054_ (.A(net972),
    .X(_06077_));
 sg13g2_or2_1 _15055_ (.X(_06078_),
    .B(net647),
    .A(net639));
 sg13g2_and2_1 _15056_ (.A(net1170),
    .B(_05687_),
    .X(_06079_));
 sg13g2_buf_1 _15057_ (.A(_06079_),
    .X(_06080_));
 sg13g2_a21oi_1 _15058_ (.A1(net640),
    .A2(_06078_),
    .Y(_06081_),
    .B1(_06080_));
 sg13g2_nor2b_1 _15059_ (.A(_06073_),
    .B_N(_06081_),
    .Y(_06082_));
 sg13g2_xnor2_1 _15060_ (.Y(_06083_),
    .A(_06073_),
    .B(_06081_));
 sg13g2_inv_1 _15061_ (.Y(_06084_),
    .A(net1173));
 sg13g2_xnor2_1 _15062_ (.Y(_06085_),
    .A(net639),
    .B(_05688_));
 sg13g2_xnor2_1 _15063_ (.Y(_06086_),
    .A(_05228_),
    .B(net973));
 sg13g2_xnor2_1 _15064_ (.Y(_06087_),
    .A(_06085_),
    .B(_06086_));
 sg13g2_xnor2_1 _15065_ (.Y(_06088_),
    .A(net986),
    .B(_06086_));
 sg13g2_xor2_1 _15066_ (.B(_06088_),
    .A(_06085_),
    .X(_06089_));
 sg13g2_a22oi_1 _15067_ (.Y(_06090_),
    .B1(_06089_),
    .B2(net353),
    .A2(_06087_),
    .A1(_06084_));
 sg13g2_mux2_1 _15068_ (.A0(_06082_),
    .A1(_06083_),
    .S(_06090_),
    .X(_06091_));
 sg13g2_xnor2_1 _15069_ (.Y(_06092_),
    .A(_05684_),
    .B(_06066_));
 sg13g2_xnor2_1 _15070_ (.Y(_06093_),
    .A(_05277_),
    .B(_06092_));
 sg13g2_xnor2_1 _15071_ (.Y(_06094_),
    .A(_06085_),
    .B(_06093_));
 sg13g2_buf_2 _15072_ (.A(\grid.cell_12_0.s ),
    .X(_06095_));
 sg13g2_buf_1 _15073_ (.A(_06095_),
    .X(_06096_));
 sg13g2_inv_1 _15074_ (.Y(_06097_),
    .A(net971));
 sg13g2_buf_1 _15075_ (.A(_00238_),
    .X(_06098_));
 sg13g2_buf_1 _15076_ (.A(_06098_),
    .X(_06099_));
 sg13g2_o21ai_1 _15077_ (.B1(net970),
    .Y(_06100_),
    .A1(net982),
    .A2(_06097_));
 sg13g2_o21ai_1 _15078_ (.B1(net127),
    .Y(_06101_),
    .A1(net971),
    .A2(_06094_));
 sg13g2_inv_1 _15079_ (.Y(_06102_),
    .A(net1174));
 sg13g2_a22oi_1 _15080_ (.Y(_06103_),
    .B1(_06101_),
    .B2(_06102_),
    .A2(_06100_),
    .A1(_06094_));
 sg13g2_nand2_1 _15081_ (.Y(_06104_),
    .A(_06091_),
    .B(_06103_));
 sg13g2_inv_1 _15082_ (.Y(_06105_),
    .A(_06098_));
 sg13g2_nand4_1 _15083_ (.B(_06090_),
    .C(_06082_),
    .A(_06105_),
    .Y(_06106_),
    .D(_06094_));
 sg13g2_a21oi_1 _15084_ (.A1(_06097_),
    .A2(_05267_),
    .Y(_06107_),
    .B1(net982));
 sg13g2_a21oi_1 _15085_ (.A1(net84),
    .A2(_06106_),
    .Y(_06108_),
    .B1(_06107_));
 sg13g2_nor2_1 _15086_ (.A(net61),
    .B(_06108_),
    .Y(_06109_));
 sg13g2_buf_2 _15087_ (.A(_00648_),
    .X(_06110_));
 sg13g2_buf_2 _15088_ (.A(_06110_),
    .X(_06111_));
 sg13g2_a221oi_1 _15089_ (.B2(_06109_),
    .C1(_06111_),
    .B1(_06104_),
    .A1(net50),
    .Y(_00301_),
    .A2(net61));
 sg13g2_buf_1 _15090_ (.A(_05175_),
    .X(_06112_));
 sg13g2_buf_2 _15091_ (.A(_06112_),
    .X(_06113_));
 sg13g2_buf_1 _15092_ (.A(_06113_),
    .X(_06114_));
 sg13g2_nor2_2 _15093_ (.A(_01989_),
    .B(net159),
    .Y(_06115_));
 sg13g2_nand2_2 _15094_ (.Y(_06116_),
    .A(net108),
    .B(_06115_));
 sg13g2_nand4_1 _15095_ (.B(net333),
    .C(net79),
    .A(net668),
    .Y(_06117_),
    .D(_06116_));
 sg13g2_buf_1 _15096_ (.A(net1056),
    .X(_06118_));
 sg13g2_nand3_1 _15097_ (.B(net49),
    .C(net61),
    .A(net637),
    .Y(_06119_));
 sg13g2_nor3_1 _15098_ (.A(net982),
    .B(net970),
    .C(net985),
    .Y(_06120_));
 sg13g2_buf_2 _15099_ (.A(\grid.cell_12_1.se ),
    .X(_06121_));
 sg13g2_buf_1 _15100_ (.A(_06121_),
    .X(_06122_));
 sg13g2_nand2_1 _15101_ (.Y(_06123_),
    .A(_05228_),
    .B(_05285_));
 sg13g2_nand2b_1 _15102_ (.Y(_06124_),
    .B(_06121_),
    .A_N(_05218_));
 sg13g2_o21ai_1 _15103_ (.B1(_06124_),
    .Y(_06125_),
    .A1(net969),
    .A2(_06123_));
 sg13g2_or2_1 _15104_ (.X(_06126_),
    .B(_05218_),
    .A(_06121_));
 sg13g2_nor2_1 _15105_ (.A(net981),
    .B(_06123_),
    .Y(_06127_));
 sg13g2_inv_2 _15106_ (.Y(_06128_),
    .A(_06074_));
 sg13g2_a221oi_1 _15107_ (.B2(_06127_),
    .C1(_06128_),
    .B1(_06126_),
    .A1(_05760_),
    .Y(_06129_),
    .A2(_06125_));
 sg13g2_nor2b_1 _15108_ (.A(_06121_),
    .B_N(_05218_),
    .Y(_06130_));
 sg13g2_a21o_1 _15109_ (.A2(_06124_),
    .A1(_05844_),
    .B1(_06130_),
    .X(_06131_));
 sg13g2_and2_1 _15110_ (.A(_06121_),
    .B(net1011),
    .X(_06132_));
 sg13g2_a21o_1 _15111_ (.A2(_06126_),
    .A1(net981),
    .B1(_06132_),
    .X(_06133_));
 sg13g2_inv_1 _15112_ (.Y(_06134_),
    .A(_06123_));
 sg13g2_a221oi_1 _15113_ (.B2(_06134_),
    .C1(net973),
    .B1(_06133_),
    .A1(_05296_),
    .Y(_06135_),
    .A2(_06131_));
 sg13g2_nor3_1 _15114_ (.A(net973),
    .B(_05760_),
    .C(_06121_),
    .Y(_06136_));
 sg13g2_nand4_1 _15115_ (.B(net1003),
    .C(net981),
    .A(net973),
    .Y(_06137_),
    .D(net969));
 sg13g2_nand2b_1 _15116_ (.Y(_06138_),
    .B(_06137_),
    .A_N(_06136_));
 sg13g2_a22oi_1 _15117_ (.Y(_06139_),
    .B1(_06130_),
    .B2(_05761_),
    .A2(_06138_),
    .A1(_05392_));
 sg13g2_o21ai_1 _15118_ (.B1(_06139_),
    .Y(_06140_),
    .A1(_06129_),
    .A2(_06135_));
 sg13g2_buf_1 _15119_ (.A(_06140_),
    .X(_06141_));
 sg13g2_and3_1 _15120_ (.X(_06142_),
    .A(net982),
    .B(net985),
    .C(_06141_));
 sg13g2_o21ai_1 _15121_ (.B1(_05247_),
    .Y(_06143_),
    .A1(_06120_),
    .A2(_06142_));
 sg13g2_nor2_1 _15122_ (.A(net674),
    .B(_06105_),
    .Y(_06144_));
 sg13g2_o21ai_1 _15123_ (.B1(net985),
    .Y(_06145_),
    .A1(_05741_),
    .A2(_06144_));
 sg13g2_nand3_1 _15124_ (.B(net970),
    .C(net985),
    .A(net982),
    .Y(_06146_));
 sg13g2_nand2_1 _15125_ (.Y(_06147_),
    .A(_06141_),
    .B(_06146_));
 sg13g2_o21ai_1 _15126_ (.B1(_06147_),
    .Y(_06148_),
    .A1(_06141_),
    .A2(_06145_));
 sg13g2_xnor2_1 _15127_ (.Y(_06149_),
    .A(_06122_),
    .B(_05797_));
 sg13g2_xor2_1 _15128_ (.B(_06149_),
    .A(_06086_),
    .X(_06150_));
 sg13g2_buf_1 _15129_ (.A(_06150_),
    .X(_06151_));
 sg13g2_a21oi_1 _15130_ (.A1(_06143_),
    .A2(_06148_),
    .Y(_06152_),
    .B1(_06151_));
 sg13g2_a21oi_1 _15131_ (.A1(net982),
    .A2(_06151_),
    .Y(_06153_),
    .B1(_06105_));
 sg13g2_nor2_1 _15132_ (.A(_06102_),
    .B(_06098_),
    .Y(_06154_));
 sg13g2_a21oi_1 _15133_ (.A1(_06151_),
    .A2(_06154_),
    .Y(_06155_),
    .B1(net353));
 sg13g2_nor3_1 _15134_ (.A(_06141_),
    .B(_06153_),
    .C(_06155_),
    .Y(_06156_));
 sg13g2_nand3_1 _15135_ (.B(net970),
    .C(net985),
    .A(_05247_),
    .Y(_06157_));
 sg13g2_nand2_1 _15136_ (.Y(_06158_),
    .A(_06102_),
    .B(_06098_));
 sg13g2_o21ai_1 _15137_ (.B1(_06158_),
    .Y(_06159_),
    .A1(net353),
    .A2(_06154_));
 sg13g2_nand2_1 _15138_ (.Y(_06160_),
    .A(_06151_),
    .B(_06159_));
 sg13g2_nand2_1 _15139_ (.Y(_06161_),
    .A(_06157_),
    .B(_06160_));
 sg13g2_and2_1 _15140_ (.A(_06141_),
    .B(_06161_),
    .X(_06162_));
 sg13g2_xnor2_1 _15141_ (.Y(_06163_),
    .A(net1174),
    .B(_06095_));
 sg13g2_xnor2_1 _15142_ (.Y(_06164_),
    .A(net674),
    .B(_06163_));
 sg13g2_xnor2_1 _15143_ (.Y(_06165_),
    .A(_06151_),
    .B(_06164_));
 sg13g2_a21oi_1 _15144_ (.A1(_04859_),
    .A2(_06165_),
    .Y(_06166_),
    .B1(net333));
 sg13g2_inv_1 _15145_ (.Y(_06167_),
    .A(net969));
 sg13g2_buf_1 _15146_ (.A(_06167_),
    .X(_06168_));
 sg13g2_nor2_1 _15147_ (.A(net326),
    .B(net1011),
    .Y(_06169_));
 sg13g2_buf_1 _15148_ (.A(net969),
    .X(_06170_));
 sg13g2_xnor2_1 _15149_ (.Y(_06171_),
    .A(net646),
    .B(net636));
 sg13g2_a21oi_1 _15150_ (.A1(net331),
    .A2(net636),
    .Y(_06172_),
    .B1(net1008));
 sg13g2_a21oi_1 _15151_ (.A1(net673),
    .A2(_06171_),
    .Y(_06173_),
    .B1(_06172_));
 sg13g2_a22oi_1 _15152_ (.Y(_06174_),
    .B1(_06173_),
    .B2(net346),
    .A2(_06169_),
    .A1(_05764_));
 sg13g2_nor2_1 _15153_ (.A(_06128_),
    .B(_06174_),
    .Y(_06175_));
 sg13g2_nand2_1 _15154_ (.Y(_06176_),
    .A(net353),
    .B(net1174));
 sg13g2_nor4_1 _15155_ (.A(_06099_),
    .B(net985),
    .C(_06151_),
    .D(_06176_),
    .Y(_06177_));
 sg13g2_buf_1 _15156_ (.A(net636),
    .X(_06178_));
 sg13g2_buf_1 _15157_ (.A(net325),
    .X(_06179_));
 sg13g2_nand3_1 _15158_ (.B(net157),
    .C(_06134_),
    .A(_05764_),
    .Y(_06180_));
 sg13g2_o21ai_1 _15159_ (.B1(_12967_),
    .Y(_06181_),
    .A1(_06075_),
    .A2(_06180_));
 sg13g2_nor4_1 _15160_ (.A(net61),
    .B(_06175_),
    .C(_06177_),
    .D(_06181_),
    .Y(_06182_));
 sg13g2_nand2b_1 _15161_ (.Y(_06183_),
    .B(_06182_),
    .A_N(_06166_));
 sg13g2_or4_1 _15162_ (.A(_06152_),
    .B(_06156_),
    .C(_06162_),
    .D(_06183_),
    .X(_06184_));
 sg13g2_nand3_1 _15163_ (.B(_06119_),
    .C(_06184_),
    .A(_06117_),
    .Y(_00302_));
 sg13g2_buf_1 _15164_ (.A(\grid.cell_12_2.se ),
    .X(_06185_));
 sg13g2_buf_1 _15165_ (.A(_06185_),
    .X(_06186_));
 sg13g2_inv_1 _15166_ (.Y(_06187_),
    .A(net968));
 sg13g2_inv_2 _15167_ (.Y(_06188_),
    .A(_05817_));
 sg13g2_nor2_2 _15168_ (.A(_06187_),
    .B(_06188_),
    .Y(_06189_));
 sg13g2_xnor2_1 _15169_ (.Y(_06190_),
    .A(_06185_),
    .B(_05817_));
 sg13g2_nor2_1 _15170_ (.A(net670),
    .B(_06190_),
    .Y(_06191_));
 sg13g2_a21o_1 _15171_ (.A2(_06189_),
    .A1(net670),
    .B1(_06191_),
    .X(_06192_));
 sg13g2_a22oi_1 _15172_ (.Y(_06193_),
    .B1(_06192_),
    .B2(net667),
    .A2(_06189_),
    .A1(_05381_));
 sg13g2_buf_1 _15173_ (.A(net968),
    .X(_06194_));
 sg13g2_buf_1 _15174_ (.A(_06194_),
    .X(_06195_));
 sg13g2_nor2_1 _15175_ (.A(net670),
    .B(net325),
    .Y(_06196_));
 sg13g2_nand4_1 _15176_ (.B(net645),
    .C(_05360_),
    .A(net324),
    .Y(_06197_),
    .D(_06196_));
 sg13g2_o21ai_1 _15177_ (.B1(_06197_),
    .Y(_06198_),
    .A1(net326),
    .A2(_06193_));
 sg13g2_buf_2 _15178_ (.A(_00237_),
    .X(_06199_));
 sg13g2_buf_1 _15179_ (.A(_06199_),
    .X(_06200_));
 sg13g2_nor2b_1 _15180_ (.A(net967),
    .B_N(net986),
    .Y(_06201_));
 sg13g2_nor2_1 _15181_ (.A(_05392_),
    .B(net980),
    .Y(_06202_));
 sg13g2_xor2_1 _15182_ (.B(net968),
    .A(net636),
    .X(_06203_));
 sg13g2_nand3_1 _15183_ (.B(_06170_),
    .C(_06187_),
    .A(net663),
    .Y(_06204_));
 sg13g2_o21ai_1 _15184_ (.B1(_06204_),
    .Y(_06205_),
    .A1(net346),
    .A2(_06203_));
 sg13g2_xor2_1 _15185_ (.B(net969),
    .A(net1003),
    .X(_06206_));
 sg13g2_xnor2_1 _15186_ (.Y(_06207_),
    .A(net635),
    .B(_06206_));
 sg13g2_nor2_1 _15187_ (.A(_05819_),
    .B(_06207_),
    .Y(_06208_));
 sg13g2_a21oi_1 _15188_ (.A1(_05819_),
    .A2(_06205_),
    .Y(_06209_),
    .B1(_06208_));
 sg13g2_nand3_1 _15189_ (.B(_05852_),
    .C(_06196_),
    .A(net324),
    .Y(_06210_));
 sg13g2_nand4_1 _15190_ (.B(_06202_),
    .C(_06209_),
    .A(_06201_),
    .Y(_06211_),
    .D(_06210_));
 sg13g2_nand2b_1 _15191_ (.Y(_06212_),
    .B(_06211_),
    .A_N(_06198_));
 sg13g2_nor2_1 _15192_ (.A(net636),
    .B(_06189_),
    .Y(_06213_));
 sg13g2_nor2_1 _15193_ (.A(net968),
    .B(_05817_),
    .Y(_06214_));
 sg13g2_o21ai_1 _15194_ (.B1(_00242_),
    .Y(_06215_),
    .A1(net663),
    .A2(net664));
 sg13g2_o21ai_1 _15195_ (.B1(_06214_),
    .Y(_06216_),
    .A1(net670),
    .A2(_05376_));
 sg13g2_o21ai_1 _15196_ (.B1(_06216_),
    .Y(_06217_),
    .A1(_06214_),
    .A2(_06215_));
 sg13g2_a21oi_1 _15197_ (.A1(net663),
    .A2(_06122_),
    .Y(_06218_),
    .B1(_05376_));
 sg13g2_nor4_1 _15198_ (.A(_06186_),
    .B(net979),
    .C(_05381_),
    .D(_06218_),
    .Y(_06219_));
 sg13g2_a21oi_2 _15199_ (.B1(_06219_),
    .Y(_06220_),
    .A2(_06217_),
    .A1(_06213_));
 sg13g2_xnor2_1 _15200_ (.Y(_06221_),
    .A(_05358_),
    .B(_06190_));
 sg13g2_xnor2_1 _15201_ (.Y(_06222_),
    .A(_06206_),
    .B(_06221_));
 sg13g2_buf_1 _15202_ (.A(_06222_),
    .X(_06223_));
 sg13g2_inv_2 _15203_ (.Y(_06224_),
    .A(_06200_));
 sg13g2_a21oi_1 _15204_ (.A1(net330),
    .A2(_06223_),
    .Y(_06225_),
    .B1(_06224_));
 sg13g2_a21oi_1 _15205_ (.A1(_06223_),
    .A2(_06201_),
    .Y(_06226_),
    .B1(net673));
 sg13g2_nor2_1 _15206_ (.A(_06225_),
    .B(_06226_),
    .Y(_06227_));
 sg13g2_nand2b_1 _15207_ (.Y(_06228_),
    .B(net967),
    .A_N(net648));
 sg13g2_o21ai_1 _15208_ (.B1(_06228_),
    .Y(_06229_),
    .A1(net673),
    .A2(_06201_));
 sg13g2_nand2_1 _15209_ (.Y(_06230_),
    .A(_06223_),
    .B(_06229_));
 sg13g2_nand3_1 _15210_ (.B(net967),
    .C(net980),
    .A(_05392_),
    .Y(_06231_));
 sg13g2_a21oi_1 _15211_ (.A1(_06230_),
    .A2(_06231_),
    .Y(_06232_),
    .B1(_06220_));
 sg13g2_a21o_1 _15212_ (.A2(_06227_),
    .A1(_06220_),
    .B1(_06232_),
    .X(_06233_));
 sg13g2_o21ai_1 _15213_ (.B1(_05268_),
    .Y(_06234_),
    .A1(_06212_),
    .A2(_06233_));
 sg13g2_nand2_1 _15214_ (.Y(_06235_),
    .A(net330),
    .B(net980));
 sg13g2_or3_1 _15215_ (.A(net648),
    .B(net967),
    .C(net980),
    .X(_06236_));
 sg13g2_o21ai_1 _15216_ (.B1(_06236_),
    .Y(_06237_),
    .A1(_06220_),
    .A2(_06235_));
 sg13g2_a21o_1 _15217_ (.A2(net967),
    .A1(_05392_),
    .B1(net330),
    .X(_06238_));
 sg13g2_nand3_1 _15218_ (.B(_06220_),
    .C(_06238_),
    .A(net980),
    .Y(_06239_));
 sg13g2_nand3_1 _15219_ (.B(_06200_),
    .C(net980),
    .A(net330),
    .Y(_06240_));
 sg13g2_nand2b_1 _15220_ (.Y(_06241_),
    .B(_06240_),
    .A_N(_06220_));
 sg13g2_a22oi_1 _15221_ (.Y(_06242_),
    .B1(_06239_),
    .B2(_06241_),
    .A2(_06237_),
    .A1(_05392_));
 sg13g2_or3_1 _15222_ (.A(net125),
    .B(_06223_),
    .C(_06242_),
    .X(_06243_));
 sg13g2_buf_1 _15223_ (.A(_05407_),
    .X(_06244_));
 sg13g2_xor2_1 _15224_ (.B(_06223_),
    .A(_06088_),
    .X(_06245_));
 sg13g2_o21ai_1 _15225_ (.B1(_05844_),
    .Y(_06246_),
    .A1(net107),
    .A2(_06245_));
 sg13g2_nand4_1 _15226_ (.B(_06234_),
    .C(_06243_),
    .A(_06116_),
    .Y(_06247_),
    .D(_06246_));
 sg13g2_nand2_1 _15227_ (.Y(_06248_),
    .A(net33),
    .B(net61));
 sg13g2_a21oi_1 _15228_ (.A1(_06247_),
    .A2(_06248_),
    .Y(_00303_),
    .B1(_05283_));
 sg13g2_buf_1 _15229_ (.A(_05469_),
    .X(_06249_));
 sg13g2_buf_1 _15230_ (.A(\grid.cell_12_3.se ),
    .X(_06250_));
 sg13g2_buf_1 _15231_ (.A(net1169),
    .X(_06251_));
 sg13g2_nor4_1 _15232_ (.A(net966),
    .B(net635),
    .C(net977),
    .D(net659),
    .Y(_06252_));
 sg13g2_inv_1 _15233_ (.Y(_06253_),
    .A(net1169));
 sg13g2_buf_1 _15234_ (.A(_06253_),
    .X(_06254_));
 sg13g2_inv_2 _15235_ (.Y(_06255_),
    .A(net1172));
 sg13g2_a21oi_1 _15236_ (.A1(_06254_),
    .A2(_06187_),
    .Y(_06256_),
    .B1(_06255_));
 sg13g2_nand2_1 _15237_ (.Y(_06257_),
    .A(net1169),
    .B(net968));
 sg13g2_o21ai_1 _15238_ (.B1(_06257_),
    .Y(_06258_),
    .A1(net659),
    .A2(net1001));
 sg13g2_nor3_1 _15239_ (.A(_06252_),
    .B(_06256_),
    .C(_06258_),
    .Y(_06259_));
 sg13g2_nand2_1 _15240_ (.Y(_06260_),
    .A(net660),
    .B(net667));
 sg13g2_nor3_1 _15241_ (.A(net966),
    .B(net324),
    .C(net978),
    .Y(_06261_));
 sg13g2_a22oi_1 _15242_ (.Y(_06262_),
    .B1(_06260_),
    .B2(_06261_),
    .A2(_06259_),
    .A1(_00042_));
 sg13g2_buf_1 _15243_ (.A(_00236_),
    .X(_06263_));
 sg13g2_nand2_1 _15244_ (.Y(_06264_),
    .A(net670),
    .B(_06263_));
 sg13g2_xnor2_1 _15245_ (.Y(_06265_),
    .A(net1169),
    .B(net1172));
 sg13g2_xnor2_1 _15246_ (.Y(_06266_),
    .A(net1175),
    .B(_06265_));
 sg13g2_xor2_1 _15247_ (.B(_05358_),
    .A(_06186_),
    .X(_06267_));
 sg13g2_xnor2_1 _15248_ (.Y(_06268_),
    .A(_06266_),
    .B(_06267_));
 sg13g2_xnor2_1 _15249_ (.Y(_06269_),
    .A(net331),
    .B(_06268_));
 sg13g2_inv_2 _15250_ (.Y(_06270_),
    .A(_06263_));
 sg13g2_nand2_1 _15251_ (.Y(_06271_),
    .A(net346),
    .B(_06270_));
 sg13g2_o21ai_1 _15252_ (.B1(_06271_),
    .Y(_06272_),
    .A1(_05877_),
    .A2(_06268_));
 sg13g2_a21oi_1 _15253_ (.A1(_06264_),
    .A2(_06269_),
    .Y(_06273_),
    .B1(_06272_));
 sg13g2_xnor2_1 _15254_ (.Y(_06274_),
    .A(_06262_),
    .B(_06273_));
 sg13g2_nor2_1 _15255_ (.A(_05877_),
    .B(_06268_),
    .Y(_06275_));
 sg13g2_and2_1 _15256_ (.A(_06270_),
    .B(_05797_),
    .X(_06276_));
 sg13g2_xor2_1 _15257_ (.B(net1001),
    .A(net977),
    .X(_06277_));
 sg13g2_nor3_1 _15258_ (.A(_06194_),
    .B(_06255_),
    .C(net664),
    .Y(_06278_));
 sg13g2_a21oi_1 _15259_ (.A1(_06195_),
    .A2(_06277_),
    .Y(_06279_),
    .B1(_06278_));
 sg13g2_nand3_1 _15260_ (.B(_06195_),
    .C(net644),
    .A(_05417_),
    .Y(_06280_));
 sg13g2_o21ai_1 _15261_ (.B1(_06280_),
    .Y(_06281_),
    .A1(net659),
    .A2(_06279_));
 sg13g2_buf_1 _15262_ (.A(net966),
    .X(_06282_));
 sg13g2_nor4_1 _15263_ (.A(net633),
    .B(_06187_),
    .C(net664),
    .D(_05886_),
    .Y(_06283_));
 sg13g2_a221oi_1 _15264_ (.B2(net633),
    .C1(_06283_),
    .B1(_06281_),
    .A1(_06275_),
    .Y(_06284_),
    .A2(_06276_));
 sg13g2_buf_1 _15265_ (.A(_05407_),
    .X(_06285_));
 sg13g2_a21oi_1 _15266_ (.A1(_06274_),
    .A2(_06284_),
    .Y(_06286_),
    .B1(net106));
 sg13g2_xnor2_1 _15267_ (.Y(_06287_),
    .A(_06149_),
    .B(_06268_));
 sg13g2_a21oi_1 _15268_ (.A1(net112),
    .A2(_06287_),
    .Y(_06288_),
    .B1(net645));
 sg13g2_or4_1 _15269_ (.A(_06110_),
    .B(net61),
    .C(_06286_),
    .D(_06288_),
    .X(_06289_));
 sg13g2_o21ai_1 _15270_ (.B1(_06289_),
    .Y(_00304_),
    .A1(net26),
    .A2(_06116_));
 sg13g2_nand2_1 _15271_ (.Y(_06290_),
    .A(net637),
    .B(_06065_));
 sg13g2_buf_1 _15272_ (.A(\grid.cell_12_4.se ),
    .X(_06291_));
 sg13g2_buf_1 _15273_ (.A(_06291_),
    .X(_06292_));
 sg13g2_buf_1 _15274_ (.A(_06292_),
    .X(_06293_));
 sg13g2_nor4_1 _15275_ (.A(net632),
    .B(net966),
    .C(net976),
    .D(_05506_),
    .Y(_06294_));
 sg13g2_inv_2 _15276_ (.Y(_06295_),
    .A(net965));
 sg13g2_inv_1 _15277_ (.Y(_06296_),
    .A(net976));
 sg13g2_a21oi_1 _15278_ (.A1(_06295_),
    .A2(net634),
    .Y(_06297_),
    .B1(_06296_));
 sg13g2_nand2_1 _15279_ (.Y(_06298_),
    .A(net632),
    .B(net1169));
 sg13g2_o21ai_1 _15280_ (.B1(_06298_),
    .Y(_06299_),
    .A1(_05506_),
    .A2(net998));
 sg13g2_nor3_1 _15281_ (.A(_06294_),
    .B(_06297_),
    .C(_06299_),
    .Y(_06300_));
 sg13g2_nand2_1 _15282_ (.Y(_06301_),
    .A(net656),
    .B(net660));
 sg13g2_nor3_1 _15283_ (.A(net632),
    .B(net633),
    .C(net329),
    .Y(_06302_));
 sg13g2_a22oi_1 _15284_ (.Y(_06303_),
    .B1(_06301_),
    .B2(_06302_),
    .A2(_06300_),
    .A1(_05484_));
 sg13g2_buf_1 _15285_ (.A(_00044_),
    .X(_06304_));
 sg13g2_nand2_1 _15286_ (.Y(_06305_),
    .A(_06304_),
    .B(net664));
 sg13g2_xnor2_1 _15287_ (.Y(_06306_),
    .A(net965),
    .B(_05911_));
 sg13g2_xor2_1 _15288_ (.B(net1175),
    .A(net1169),
    .X(_06307_));
 sg13g2_xnor2_1 _15289_ (.Y(_06308_),
    .A(_06306_),
    .B(_06307_));
 sg13g2_xnor2_1 _15290_ (.Y(_06309_),
    .A(net645),
    .B(_06308_));
 sg13g2_inv_1 _15291_ (.Y(_06310_),
    .A(_06304_));
 sg13g2_nand2_1 _15292_ (.Y(_06311_),
    .A(_06310_),
    .B(net667));
 sg13g2_o21ai_1 _15293_ (.B1(_06311_),
    .Y(_06312_),
    .A1(_05916_),
    .A2(_06308_));
 sg13g2_a21oi_1 _15294_ (.A1(_06305_),
    .A2(_06309_),
    .Y(_06313_),
    .B1(_06312_));
 sg13g2_xnor2_1 _15295_ (.Y(_06314_),
    .A(_06303_),
    .B(_06313_));
 sg13g2_nor2_1 _15296_ (.A(_05916_),
    .B(_06308_),
    .Y(_06315_));
 sg13g2_and2_1 _15297_ (.A(_06310_),
    .B(_05819_),
    .X(_06316_));
 sg13g2_nand2_1 _15298_ (.Y(_06317_),
    .A(net966),
    .B(net643));
 sg13g2_xnor2_1 _15299_ (.Y(_06318_),
    .A(net976),
    .B(net998));
 sg13g2_nor2_1 _15300_ (.A(net634),
    .B(_06318_),
    .Y(_06319_));
 sg13g2_nor3_1 _15301_ (.A(_06251_),
    .B(_06296_),
    .C(net659),
    .Y(_06320_));
 sg13g2_o21ai_1 _15302_ (.B1(net344),
    .Y(_06321_),
    .A1(_06319_),
    .A2(_06320_));
 sg13g2_o21ai_1 _15303_ (.B1(_06321_),
    .Y(_06322_),
    .A1(_05484_),
    .A2(_06317_));
 sg13g2_buf_1 _15304_ (.A(_06293_),
    .X(_06323_));
 sg13g2_nor3_1 _15305_ (.A(net323),
    .B(_06317_),
    .C(_06301_),
    .Y(_06324_));
 sg13g2_a221oi_1 _15306_ (.B2(_06323_),
    .C1(_06324_),
    .B1(_06322_),
    .A1(_06315_),
    .Y(_06325_),
    .A2(_06316_));
 sg13g2_a21oi_1 _15307_ (.A1(_06314_),
    .A2(_06325_),
    .Y(_06326_),
    .B1(net106));
 sg13g2_xnor2_1 _15308_ (.Y(_06327_),
    .A(_06221_),
    .B(_06308_));
 sg13g2_a21oi_1 _15309_ (.A1(net112),
    .A2(_06327_),
    .Y(_06328_),
    .B1(net644));
 sg13g2_or4_1 _15310_ (.A(_00659_),
    .B(_06065_),
    .C(_06326_),
    .D(_06328_),
    .X(_06329_));
 sg13g2_o21ai_1 _15311_ (.B1(_06329_),
    .Y(_00305_),
    .A1(_04942_),
    .A2(_06290_));
 sg13g2_inv_2 _15312_ (.Y(_06330_),
    .A(_05002_));
 sg13g2_buf_1 _15313_ (.A(_05407_),
    .X(_06331_));
 sg13g2_buf_1 _15314_ (.A(_00076_),
    .X(_06332_));
 sg13g2_a22oi_1 _15315_ (.Y(_06333_),
    .B1(_06255_),
    .B2(net660),
    .A2(net1168),
    .A1(_05952_));
 sg13g2_nand3_1 _15316_ (.B(_05865_),
    .C(net659),
    .A(_05952_),
    .Y(_06334_));
 sg13g2_nor2b_1 _15317_ (.A(net1171),
    .B_N(_05523_),
    .Y(_06335_));
 sg13g2_buf_2 _15318_ (.A(\grid.cell_12_5.se ),
    .X(_06336_));
 sg13g2_nor2_1 _15319_ (.A(_06336_),
    .B(net965),
    .Y(_06337_));
 sg13g2_and2_1 _15320_ (.A(net965),
    .B(net1171),
    .X(_06338_));
 sg13g2_a221oi_1 _15321_ (.B2(_06337_),
    .C1(_06338_),
    .B1(_06335_),
    .A1(_05523_),
    .Y(_06339_),
    .A2(_05506_));
 sg13g2_buf_1 _15322_ (.A(_06336_),
    .X(_06340_));
 sg13g2_o21ai_1 _15323_ (.B1(net964),
    .Y(_06341_),
    .A1(net965),
    .A2(net1171));
 sg13g2_and2_1 _15324_ (.A(_05553_),
    .B(_06341_),
    .X(_06342_));
 sg13g2_nand2_1 _15325_ (.Y(_06343_),
    .A(net992),
    .B(net995));
 sg13g2_nor3_1 _15326_ (.A(net964),
    .B(net965),
    .C(net975),
    .Y(_06344_));
 sg13g2_a22oi_1 _15327_ (.Y(_06345_),
    .B1(_06343_),
    .B2(_06344_),
    .A2(_06342_),
    .A1(_06339_));
 sg13g2_buf_1 _15328_ (.A(_06345_),
    .X(_06346_));
 sg13g2_a21oi_1 _15329_ (.A1(_06333_),
    .A2(_06334_),
    .Y(_06347_),
    .B1(_06346_));
 sg13g2_nand2b_1 _15330_ (.Y(_06348_),
    .B(net998),
    .A_N(_00076_));
 sg13g2_and4_1 _15331_ (.A(_05951_),
    .B(_05865_),
    .C(_06346_),
    .D(_06348_),
    .X(_06349_));
 sg13g2_xor2_1 _15332_ (.B(_05523_),
    .A(net1171),
    .X(_06350_));
 sg13g2_xnor2_1 _15333_ (.Y(_06351_),
    .A(_06336_),
    .B(_06292_));
 sg13g2_xor2_1 _15334_ (.B(_06351_),
    .A(_06350_),
    .X(_06352_));
 sg13g2_xnor2_1 _15335_ (.Y(_06353_),
    .A(net995),
    .B(_06352_));
 sg13g2_buf_1 _15336_ (.A(_06353_),
    .X(_06354_));
 sg13g2_o21ai_1 _15337_ (.B1(_06354_),
    .Y(_06355_),
    .A1(_06347_),
    .A2(_06349_));
 sg13g2_nor2_1 _15338_ (.A(_05883_),
    .B(net998),
    .Y(_06356_));
 sg13g2_a21oi_1 _15339_ (.A1(net1168),
    .A2(_05886_),
    .Y(_06357_),
    .B1(_06356_));
 sg13g2_nand3_1 _15340_ (.B(net1168),
    .C(net659),
    .A(_05951_),
    .Y(_06358_));
 sg13g2_o21ai_1 _15341_ (.B1(_06358_),
    .Y(_06359_),
    .A1(_06354_),
    .A2(_06357_));
 sg13g2_nor3_1 _15342_ (.A(_05886_),
    .B(_06354_),
    .C(_06346_),
    .Y(_06360_));
 sg13g2_a21oi_1 _15343_ (.A1(_06346_),
    .A2(_06359_),
    .Y(_06361_),
    .B1(_06360_));
 sg13g2_inv_1 _15344_ (.Y(_06362_),
    .A(net964));
 sg13g2_xnor2_1 _15345_ (.Y(_06363_),
    .A(net641),
    .B(net995));
 sg13g2_a21oi_1 _15346_ (.A1(net642),
    .A2(net656),
    .Y(_06364_),
    .B1(net632));
 sg13g2_a21oi_1 _15347_ (.A1(_06293_),
    .A2(_06363_),
    .Y(_06365_),
    .B1(_06364_));
 sg13g2_a22oi_1 _15348_ (.Y(_06366_),
    .B1(_06365_),
    .B2(net162),
    .A2(_06338_),
    .A1(_05980_));
 sg13g2_buf_1 _15349_ (.A(_06340_),
    .X(_06367_));
 sg13g2_buf_1 _15350_ (.A(net630),
    .X(_06368_));
 sg13g2_nor2_1 _15351_ (.A(net322),
    .B(_05959_),
    .Y(_06369_));
 sg13g2_nand3_1 _15352_ (.B(_05490_),
    .C(_06369_),
    .A(_06323_),
    .Y(_06370_));
 sg13g2_o21ai_1 _15353_ (.B1(_06370_),
    .Y(_06371_),
    .A1(net631),
    .A2(_06366_));
 sg13g2_a21oi_1 _15354_ (.A1(_06355_),
    .A2(_06361_),
    .Y(_06372_),
    .B1(_06371_));
 sg13g2_a21oi_1 _15355_ (.A1(_05866_),
    .A2(_05444_),
    .Y(_06373_),
    .B1(_05952_));
 sg13g2_nor2_1 _15356_ (.A(_06354_),
    .B(_06356_),
    .Y(_06374_));
 sg13g2_a21oi_1 _15357_ (.A1(_06354_),
    .A2(_06373_),
    .Y(_06375_),
    .B1(_06374_));
 sg13g2_nor3_1 _15358_ (.A(net1168),
    .B(_06346_),
    .C(_06375_),
    .Y(_06376_));
 sg13g2_or3_1 _15359_ (.A(net105),
    .B(_06372_),
    .C(_06376_),
    .X(_06377_));
 sg13g2_xor2_1 _15360_ (.B(_06354_),
    .A(_06266_),
    .X(_06378_));
 sg13g2_a21oi_1 _15361_ (.A1(net113),
    .A2(_06378_),
    .Y(_06379_),
    .B1(net329));
 sg13g2_nor2_1 _15362_ (.A(net61),
    .B(_06379_),
    .Y(_06380_));
 sg13g2_a22oi_1 _15363_ (.Y(_06381_),
    .B1(_06377_),
    .B2(_06380_),
    .A2(net61),
    .A1(_06330_));
 sg13g2_nor2_1 _15364_ (.A(net370),
    .B(_06381_),
    .Y(_00306_));
 sg13g2_nor2b_1 _15365_ (.A(_05600_),
    .B_N(_06080_),
    .Y(_06382_));
 sg13g2_buf_1 _15366_ (.A(net972),
    .X(_06383_));
 sg13g2_xnor2_1 _15367_ (.Y(_06384_),
    .A(net332),
    .B(net992));
 sg13g2_o21ai_1 _15368_ (.B1(net335),
    .Y(_06385_),
    .A1(net629),
    .A2(_06031_));
 sg13g2_a21oi_1 _15369_ (.A1(net629),
    .A2(_06384_),
    .Y(_06386_),
    .B1(_06385_));
 sg13g2_nor2_1 _15370_ (.A(_06382_),
    .B(_06386_),
    .Y(_06387_));
 sg13g2_and2_1 _15371_ (.A(net1170),
    .B(net1015),
    .X(_06388_));
 sg13g2_buf_1 _15372_ (.A(_06388_),
    .X(_06389_));
 sg13g2_a21oi_1 _15373_ (.A1(_06031_),
    .A2(_06389_),
    .Y(_06390_),
    .B1(net322));
 sg13g2_a21oi_1 _15374_ (.A1(_06368_),
    .A2(_06387_),
    .Y(_06391_),
    .B1(_06390_));
 sg13g2_buf_2 _15375_ (.A(_00108_),
    .X(_06392_));
 sg13g2_inv_1 _15376_ (.Y(_06393_),
    .A(_05911_));
 sg13g2_xnor2_1 _15377_ (.Y(_06394_),
    .A(_06336_),
    .B(net1170));
 sg13g2_xor2_1 _15378_ (.B(_06394_),
    .A(_05688_),
    .X(_06395_));
 sg13g2_xnor2_1 _15379_ (.Y(_06396_),
    .A(net992),
    .B(_06395_));
 sg13g2_nor4_1 _15380_ (.A(_05985_),
    .B(_06392_),
    .C(_06393_),
    .D(_06396_),
    .Y(_06397_));
 sg13g2_nor3_1 _15381_ (.A(net170),
    .B(_06391_),
    .C(_06397_),
    .Y(_06398_));
 sg13g2_nand2_1 _15382_ (.Y(_06399_),
    .A(_06392_),
    .B(_05506_));
 sg13g2_xnor2_1 _15383_ (.Y(_06400_),
    .A(net643),
    .B(_06396_));
 sg13g2_nand2b_1 _15384_ (.Y(_06401_),
    .B(_05489_),
    .A_N(_06392_));
 sg13g2_o21ai_1 _15385_ (.B1(_06401_),
    .Y(_06402_),
    .A1(_05985_),
    .A2(_06396_));
 sg13g2_a21oi_1 _15386_ (.A1(_06399_),
    .A2(_06400_),
    .Y(_06403_),
    .B1(_06402_));
 sg13g2_o21ai_1 _15387_ (.B1(_06078_),
    .Y(_06404_),
    .A1(net630),
    .A2(_06080_));
 sg13g2_nor3_1 _15388_ (.A(net964),
    .B(net639),
    .C(_05700_),
    .Y(_06405_));
 sg13g2_a21oi_1 _15389_ (.A1(net988),
    .A2(_06404_),
    .Y(_06406_),
    .B1(_06405_));
 sg13g2_nand2_1 _15390_ (.Y(_06407_),
    .A(_05523_),
    .B(net1015));
 sg13g2_nor3_1 _15391_ (.A(_05600_),
    .B(_06076_),
    .C(net984),
    .Y(_06408_));
 sg13g2_nor3_1 _15392_ (.A(_06080_),
    .B(_06407_),
    .C(_06408_),
    .Y(_06409_));
 sg13g2_or2_1 _15393_ (.X(_06410_),
    .B(_06409_),
    .A(_06382_));
 sg13g2_nand2b_1 _15394_ (.Y(_06411_),
    .B(net639),
    .A_N(_05600_));
 sg13g2_nor2b_1 _15395_ (.A(net639),
    .B_N(_05699_),
    .Y(_06412_));
 sg13g2_nor2b_1 _15396_ (.A(net964),
    .B_N(_05600_),
    .Y(_06413_));
 sg13g2_o21ai_1 _15397_ (.B1(_06413_),
    .Y(_06414_),
    .A1(_06412_),
    .A2(_06389_));
 sg13g2_o21ai_1 _15398_ (.B1(_06414_),
    .Y(_06415_),
    .A1(_05728_),
    .A2(_06411_));
 sg13g2_and2_1 _15399_ (.A(_06340_),
    .B(net972),
    .X(_06416_));
 sg13g2_buf_2 _15400_ (.A(_06416_),
    .X(_06417_));
 sg13g2_a21oi_1 _15401_ (.A1(_05706_),
    .A2(_06417_),
    .Y(_06418_),
    .B1(_06405_));
 sg13g2_nor2_1 _15402_ (.A(net653),
    .B(_06418_),
    .Y(_06419_));
 sg13g2_a221oi_1 _15403_ (.B2(net341),
    .C1(_06419_),
    .B1(_06415_),
    .A1(_06367_),
    .Y(_06420_),
    .A2(_06410_));
 sg13g2_o21ai_1 _15404_ (.B1(_06420_),
    .Y(_06421_),
    .A1(net355),
    .A2(_06406_));
 sg13g2_xor2_1 _15405_ (.B(_06421_),
    .A(_06403_),
    .X(_06422_));
 sg13g2_xnor2_1 _15406_ (.Y(_06423_),
    .A(_06306_),
    .B(_06396_));
 sg13g2_and3_1 _15407_ (.X(_06424_),
    .A(_06398_),
    .B(_06422_),
    .C(_06423_));
 sg13g2_buf_1 _15408_ (.A(net168),
    .X(_06425_));
 sg13g2_a21o_1 _15409_ (.A2(_06422_),
    .A1(_06398_),
    .B1(net104),
    .X(_06426_));
 sg13g2_o21ai_1 _15410_ (.B1(_06426_),
    .Y(_06427_),
    .A1(net328),
    .A2(_06424_));
 sg13g2_o21ai_1 _15411_ (.B1(net334),
    .Y(_06428_),
    .A1(net31),
    .A2(_06116_));
 sg13g2_a21oi_1 _15412_ (.A1(_06116_),
    .A2(_06427_),
    .Y(_00307_),
    .B1(_06428_));
 sg13g2_nor2_1 _15413_ (.A(_06077_),
    .B(_05937_),
    .Y(_06429_));
 sg13g2_nand2_1 _15414_ (.Y(_06430_),
    .A(net631),
    .B(_06429_));
 sg13g2_and2_1 _15415_ (.A(_06076_),
    .B(net1171),
    .X(_06431_));
 sg13g2_buf_1 _15416_ (.A(_06431_),
    .X(_06432_));
 sg13g2_nor2_1 _15417_ (.A(_06367_),
    .B(_06432_),
    .Y(_06433_));
 sg13g2_o21ai_1 _15418_ (.B1(net988),
    .Y(_06434_),
    .A1(_06429_),
    .A2(_06433_));
 sg13g2_a21oi_1 _15419_ (.A1(_06430_),
    .A2(_06434_),
    .Y(_06435_),
    .B1(net355));
 sg13g2_nor2b_1 _15420_ (.A(_05600_),
    .B_N(_06432_),
    .Y(_06436_));
 sg13g2_nor3_1 _15421_ (.A(_05600_),
    .B(_06383_),
    .C(net641),
    .Y(_06437_));
 sg13g2_nor3_1 _15422_ (.A(_06407_),
    .B(_06432_),
    .C(_06437_),
    .Y(_06438_));
 sg13g2_o21ai_1 _15423_ (.B1(_06368_),
    .Y(_06439_),
    .A1(_06436_),
    .A2(_06438_));
 sg13g2_nand2_1 _15424_ (.Y(_06440_),
    .A(net641),
    .B(net335));
 sg13g2_nor2b_1 _15425_ (.A(_06077_),
    .B_N(net975),
    .Y(_06441_));
 sg13g2_o21ai_1 _15426_ (.B1(_06413_),
    .Y(_06442_),
    .A1(_06389_),
    .A2(_06441_));
 sg13g2_o21ai_1 _15427_ (.B1(_06442_),
    .Y(_06443_),
    .A1(_06411_),
    .A2(_06440_));
 sg13g2_nand3_1 _15428_ (.B(net335),
    .C(_06417_),
    .A(net641),
    .Y(_06444_));
 sg13g2_a21oi_1 _15429_ (.A1(_06430_),
    .A2(_06444_),
    .Y(_06445_),
    .B1(net341));
 sg13g2_a21oi_1 _15430_ (.A1(net341),
    .A2(_06443_),
    .Y(_06446_),
    .B1(_06445_));
 sg13g2_nand3b_1 _15431_ (.B(_06439_),
    .C(_06446_),
    .Y(_06447_),
    .A_N(_06435_));
 sg13g2_xor2_1 _15432_ (.B(_06394_),
    .A(_06350_),
    .X(_06448_));
 sg13g2_xnor2_1 _15433_ (.Y(_06449_),
    .A(net679),
    .B(_06448_));
 sg13g2_xnor2_1 _15434_ (.Y(_06450_),
    .A(_06102_),
    .B(_06449_));
 sg13g2_nor2_1 _15435_ (.A(net985),
    .B(_06449_),
    .Y(_06451_));
 sg13g2_a21oi_1 _15436_ (.A1(net353),
    .A2(_06105_),
    .Y(_06452_),
    .B1(_06451_));
 sg13g2_o21ai_1 _15437_ (.B1(_06452_),
    .Y(_06453_),
    .A1(_06144_),
    .A2(_06450_));
 sg13g2_xor2_1 _15438_ (.B(_06453_),
    .A(_06447_),
    .X(_06454_));
 sg13g2_xor2_1 _15439_ (.B(_05741_),
    .A(net353),
    .X(_06455_));
 sg13g2_nor4_1 _15440_ (.A(_06099_),
    .B(net985),
    .C(_06449_),
    .D(_06455_),
    .Y(_06456_));
 sg13g2_buf_1 _15441_ (.A(_06383_),
    .X(_06457_));
 sg13g2_nand2_1 _15442_ (.Y(_06458_),
    .A(net321),
    .B(_06350_));
 sg13g2_o21ai_1 _15443_ (.B1(_06458_),
    .Y(_06459_),
    .A1(_06457_),
    .A2(_05959_));
 sg13g2_a21oi_1 _15444_ (.A1(net355),
    .A2(_06459_),
    .Y(_06460_),
    .B1(_06436_));
 sg13g2_a21oi_1 _15445_ (.A1(_06369_),
    .A2(_06389_),
    .Y(_06461_),
    .B1(net163));
 sg13g2_o21ai_1 _15446_ (.B1(_06461_),
    .Y(_06462_),
    .A1(_06362_),
    .A2(_06460_));
 sg13g2_xnor2_1 _15447_ (.Y(_06463_),
    .A(_06164_),
    .B(_06449_));
 sg13g2_nor2_1 _15448_ (.A(_05710_),
    .B(_06463_),
    .Y(_06464_));
 sg13g2_or4_1 _15449_ (.A(_06454_),
    .B(_06456_),
    .C(_06462_),
    .D(_06464_),
    .X(_06465_));
 sg13g2_buf_1 _15450_ (.A(net168),
    .X(_06466_));
 sg13g2_nor2_1 _15451_ (.A(net176),
    .B(_05128_),
    .Y(_06467_));
 sg13g2_buf_2 _15452_ (.A(_06467_),
    .X(_06468_));
 sg13g2_a22oi_1 _15453_ (.Y(_06469_),
    .B1(_06115_),
    .B2(net76),
    .A2(net103),
    .A1(net161));
 sg13g2_nor2_1 _15454_ (.A(net176),
    .B(net80),
    .Y(_06470_));
 sg13g2_buf_2 _15455_ (.A(_06470_),
    .X(_06471_));
 sg13g2_a221oi_1 _15456_ (.B2(_06115_),
    .C1(net638),
    .B1(_06471_),
    .A1(_06465_),
    .Y(_00308_),
    .A2(_06469_));
 sg13g2_buf_1 _15457_ (.A(_01956_),
    .X(_06472_));
 sg13g2_nand3b_1 _15458_ (.B(_01935_),
    .C(net177),
    .Y(_06473_),
    .A_N(net320));
 sg13g2_buf_2 _15459_ (.A(_06473_),
    .X(_06474_));
 sg13g2_nor3_1 _15460_ (.A(net375),
    .B(net159),
    .C(_06474_),
    .Y(_06475_));
 sg13g2_buf_1 _15461_ (.A(_06475_),
    .X(_06476_));
 sg13g2_nand2_1 _15462_ (.Y(_06477_),
    .A(_05757_),
    .B(net60));
 sg13g2_buf_2 _15463_ (.A(\grid.cell_13_0.se ),
    .X(_06478_));
 sg13g2_buf_2 _15464_ (.A(\grid.cell_13_0.sw ),
    .X(_06479_));
 sg13g2_xnor2_1 _15465_ (.Y(_06480_),
    .A(_06479_),
    .B(net1170));
 sg13g2_xnor2_1 _15466_ (.Y(_06481_),
    .A(_06478_),
    .B(_06480_));
 sg13g2_buf_2 _15467_ (.A(_06481_),
    .X(_06482_));
 sg13g2_xor2_1 _15468_ (.B(_06482_),
    .A(net648),
    .X(_06483_));
 sg13g2_a22oi_1 _15469_ (.Y(_06484_),
    .B1(_06483_),
    .B2(net161),
    .A2(_06482_),
    .A1(_06084_));
 sg13g2_or2_1 _15470_ (.X(_06485_),
    .B(net1170),
    .A(_06479_));
 sg13g2_buf_1 _15471_ (.A(_06485_),
    .X(_06486_));
 sg13g2_inv_1 _15472_ (.Y(_06487_),
    .A(_06478_));
 sg13g2_buf_1 _15473_ (.A(_06487_),
    .X(_06488_));
 sg13g2_nand2_1 _15474_ (.Y(_06489_),
    .A(net628),
    .B(net647));
 sg13g2_and2_1 _15475_ (.A(_06479_),
    .B(net1170),
    .X(_06490_));
 sg13g2_buf_2 _15476_ (.A(_06490_),
    .X(_06491_));
 sg13g2_nand3_1 _15477_ (.B(net1173),
    .C(_06491_),
    .A(_06478_),
    .Y(_06492_));
 sg13g2_o21ai_1 _15478_ (.B1(_06492_),
    .Y(_06493_),
    .A1(_06486_),
    .A2(_06489_));
 sg13g2_and2_1 _15479_ (.A(net648),
    .B(_06493_),
    .X(_06494_));
 sg13g2_buf_1 _15480_ (.A(_06478_),
    .X(_06495_));
 sg13g2_buf_1 _15481_ (.A(_06479_),
    .X(_06496_));
 sg13g2_nor2_1 _15482_ (.A(net962),
    .B(net972),
    .Y(_06497_));
 sg13g2_nand2b_1 _15483_ (.Y(_06498_),
    .B(net1170),
    .A_N(net1173));
 sg13g2_mux2_1 _15484_ (.A0(net972),
    .A1(_06498_),
    .S(net962),
    .X(_06499_));
 sg13g2_nand2b_1 _15485_ (.Y(_06500_),
    .B(net962),
    .A_N(net972));
 sg13g2_nand2b_1 _15486_ (.Y(_06501_),
    .B(net984),
    .A_N(net962));
 sg13g2_a21oi_1 _15487_ (.A1(_06500_),
    .A2(_06501_),
    .Y(_06502_),
    .B1(net986));
 sg13g2_a221oi_1 _15488_ (.B2(_05715_),
    .C1(_06502_),
    .B1(_06499_),
    .A1(_06084_),
    .Y(_06503_),
    .A2(_06497_));
 sg13g2_nor2_1 _15489_ (.A(_05734_),
    .B(_06497_),
    .Y(_06504_));
 sg13g2_mux2_1 _15490_ (.A0(net1173),
    .A1(net984),
    .S(net972),
    .X(_06505_));
 sg13g2_nor2b_1 _15491_ (.A(_06505_),
    .B_N(_06496_),
    .Y(_06506_));
 sg13g2_buf_1 _15492_ (.A(_06496_),
    .X(_06507_));
 sg13g2_nor2_1 _15493_ (.A(net627),
    .B(_06498_),
    .Y(_06508_));
 sg13g2_nor4_1 _15494_ (.A(net963),
    .B(_06504_),
    .C(_06506_),
    .D(_06508_),
    .Y(_06509_));
 sg13g2_a21oi_1 _15495_ (.A1(net963),
    .A2(_06503_),
    .Y(_06510_),
    .B1(_06509_));
 sg13g2_buf_1 _15496_ (.A(_00235_),
    .X(_06511_));
 sg13g2_inv_1 _15497_ (.Y(_06512_),
    .A(_06511_));
 sg13g2_xnor2_1 _15498_ (.Y(_06513_),
    .A(net1174),
    .B(_05687_));
 sg13g2_xnor2_1 _15499_ (.Y(_06514_),
    .A(_06092_),
    .B(_06513_));
 sg13g2_xnor2_1 _15500_ (.Y(_06515_),
    .A(_06482_),
    .B(_06514_));
 sg13g2_and2_1 _15501_ (.A(_06512_),
    .B(_06515_),
    .X(_06516_));
 sg13g2_o21ai_1 _15502_ (.B1(_06516_),
    .Y(_06517_),
    .A1(_06494_),
    .A2(_06510_));
 sg13g2_or3_1 _15503_ (.A(_06516_),
    .B(_06494_),
    .C(_06510_),
    .X(_06518_));
 sg13g2_xnor2_1 _15504_ (.Y(_06519_),
    .A(_05685_),
    .B(net984));
 sg13g2_xnor2_1 _15505_ (.Y(_06520_),
    .A(_06482_),
    .B(_06519_));
 sg13g2_nand2_1 _15506_ (.Y(_06521_),
    .A(_06224_),
    .B(_06520_));
 sg13g2_xnor2_1 _15507_ (.Y(_06522_),
    .A(_06128_),
    .B(_06520_));
 sg13g2_nand2_1 _15508_ (.Y(_06523_),
    .A(net982),
    .B(_06522_));
 sg13g2_and4_1 _15509_ (.A(_06517_),
    .B(_06518_),
    .C(_06521_),
    .D(_06523_),
    .X(_06524_));
 sg13g2_a21oi_1 _15510_ (.A1(_06495_),
    .A2(_06486_),
    .Y(_06525_),
    .B1(_06491_));
 sg13g2_nand2_1 _15511_ (.Y(_06526_),
    .A(_06484_),
    .B(_06525_));
 sg13g2_a221oi_1 _15512_ (.B2(_06523_),
    .C1(_06526_),
    .B1(_06521_),
    .A1(_06517_),
    .Y(_06527_),
    .A2(_06518_));
 sg13g2_a21oi_1 _15513_ (.A1(_06484_),
    .A2(_06524_),
    .Y(_06528_),
    .B1(_06527_));
 sg13g2_a21oi_1 _15514_ (.A1(_06524_),
    .A2(_06525_),
    .Y(_06529_),
    .B1(net117));
 sg13g2_nor2_2 _15515_ (.A(net159),
    .B(_06474_),
    .Y(_06530_));
 sg13g2_nand2_2 _15516_ (.Y(_06531_),
    .A(net108),
    .B(_06530_));
 sg13g2_buf_1 _15517_ (.A(\grid.cell_13_0.s ),
    .X(_06532_));
 sg13g2_buf_1 _15518_ (.A(_06532_),
    .X(_06533_));
 sg13g2_xnor2_1 _15519_ (.Y(_06534_),
    .A(_06533_),
    .B(_06515_));
 sg13g2_o21ai_1 _15520_ (.B1(_06097_),
    .Y(_06535_),
    .A1(_04915_),
    .A2(_06534_));
 sg13g2_nand2_1 _15521_ (.Y(_06536_),
    .A(_06531_),
    .B(_06535_));
 sg13g2_a21o_1 _15522_ (.A2(_06529_),
    .A1(_06528_),
    .B1(_06536_),
    .X(_06537_));
 sg13g2_a21oi_1 _15523_ (.A1(_06477_),
    .A2(_06537_),
    .Y(_00309_),
    .B1(net350));
 sg13g2_buf_1 _15524_ (.A(net105),
    .X(_06538_));
 sg13g2_buf_2 _15525_ (.A(\grid.cell_13_1.se ),
    .X(_06539_));
 sg13g2_buf_1 _15526_ (.A(_06539_),
    .X(_06540_));
 sg13g2_inv_1 _15527_ (.Y(_06541_),
    .A(net960));
 sg13g2_buf_1 _15528_ (.A(_06541_),
    .X(_06542_));
 sg13g2_nand3_1 _15529_ (.B(_06168_),
    .C(_06542_),
    .A(net628),
    .Y(_06543_));
 sg13g2_buf_1 _15530_ (.A(net960),
    .X(_06544_));
 sg13g2_nand4_1 _15531_ (.B(net331),
    .C(_06178_),
    .A(_06495_),
    .Y(_06545_),
    .D(net626));
 sg13g2_a21oi_1 _15532_ (.A1(_06543_),
    .A2(_06545_),
    .Y(_06546_),
    .B1(net333));
 sg13g2_nor4_1 _15533_ (.A(net160),
    .B(net157),
    .C(_06544_),
    .D(_06084_),
    .Y(_06547_));
 sg13g2_buf_1 _15534_ (.A(net960),
    .X(_06548_));
 sg13g2_nand2_1 _15535_ (.Y(_06549_),
    .A(net986),
    .B(net646));
 sg13g2_nand2b_1 _15536_ (.Y(_06550_),
    .B(net960),
    .A_N(net1173));
 sg13g2_o21ai_1 _15537_ (.B1(_06550_),
    .Y(_06551_),
    .A1(net625),
    .A2(_06549_));
 sg13g2_nor2_1 _15538_ (.A(net625),
    .B(net1173),
    .Y(_06552_));
 sg13g2_nor3_1 _15539_ (.A(_06178_),
    .B(_06549_),
    .C(_06552_),
    .Y(_06553_));
 sg13g2_a21oi_1 _15540_ (.A1(net157),
    .A2(_06551_),
    .Y(_06554_),
    .B1(_06553_));
 sg13g2_nor2_1 _15541_ (.A(net628),
    .B(_06554_),
    .Y(_06555_));
 sg13g2_buf_1 _15542_ (.A(net963),
    .X(_06556_));
 sg13g2_nand2_1 _15543_ (.Y(_06557_),
    .A(_06168_),
    .B(_06550_));
 sg13g2_o21ai_1 _15544_ (.B1(_06557_),
    .Y(_06558_),
    .A1(net625),
    .A2(_06084_));
 sg13g2_nand2_1 _15545_ (.Y(_06559_),
    .A(net625),
    .B(net1173));
 sg13g2_o21ai_1 _15546_ (.B1(_06170_),
    .Y(_06560_),
    .A1(_06540_),
    .A2(net1173));
 sg13g2_a21oi_1 _15547_ (.A1(_06559_),
    .A2(_06560_),
    .Y(_06561_),
    .B1(_06549_));
 sg13g2_a21oi_1 _15548_ (.A1(_05844_),
    .A2(_06558_),
    .Y(_06562_),
    .B1(_06561_));
 sg13g2_nor2_1 _15549_ (.A(_06556_),
    .B(_06562_),
    .Y(_06563_));
 sg13g2_nor4_1 _15550_ (.A(_06546_),
    .B(_06547_),
    .C(_06555_),
    .D(_06563_),
    .Y(_06564_));
 sg13g2_nand2_1 _15551_ (.Y(_06565_),
    .A(_06102_),
    .B(_06511_));
 sg13g2_xnor2_1 _15552_ (.Y(_06566_),
    .A(_06121_),
    .B(_06539_));
 sg13g2_xnor2_1 _15553_ (.Y(_06567_),
    .A(net646),
    .B(_06566_));
 sg13g2_xor2_1 _15554_ (.B(_06478_),
    .A(net986),
    .X(_06568_));
 sg13g2_xnor2_1 _15555_ (.Y(_06569_),
    .A(_06567_),
    .B(_06568_));
 sg13g2_xnor2_1 _15556_ (.Y(_06570_),
    .A(net971),
    .B(_06569_));
 sg13g2_nand2_1 _15557_ (.Y(_06571_),
    .A(_05740_),
    .B(_06512_));
 sg13g2_o21ai_1 _15558_ (.B1(_06571_),
    .Y(_06572_),
    .A1(net970),
    .A2(_06569_));
 sg13g2_a21oi_1 _15559_ (.A1(_06565_),
    .A2(_06570_),
    .Y(_06573_),
    .B1(_06572_));
 sg13g2_xnor2_1 _15560_ (.Y(_06574_),
    .A(_06564_),
    .B(_06573_));
 sg13g2_nor2_1 _15561_ (.A(net319),
    .B(net980),
    .Y(_06575_));
 sg13g2_a21oi_1 _15562_ (.A1(net325),
    .A2(net626),
    .Y(_06576_),
    .B1(net648));
 sg13g2_a21oi_1 _15563_ (.A1(net330),
    .A2(_06566_),
    .Y(_06577_),
    .B1(_06576_));
 sg13g2_a22oi_1 _15564_ (.Y(_06578_),
    .B1(_06577_),
    .B2(net160),
    .A2(_06575_),
    .A1(_06179_));
 sg13g2_nand4_1 _15565_ (.B(net160),
    .C(_06179_),
    .A(net330),
    .Y(_06579_),
    .D(_06544_));
 sg13g2_nand2b_1 _15566_ (.Y(_06580_),
    .B(_06488_),
    .A_N(_06579_));
 sg13g2_o21ai_1 _15567_ (.B1(_06580_),
    .Y(_06581_),
    .A1(_06488_),
    .A2(_06578_));
 sg13g2_xor2_1 _15568_ (.B(_06095_),
    .A(_05740_),
    .X(_06582_));
 sg13g2_nor4_1 _15569_ (.A(_06511_),
    .B(net970),
    .C(_06582_),
    .D(_06569_),
    .Y(_06583_));
 sg13g2_xnor2_1 _15570_ (.Y(_06584_),
    .A(_06532_),
    .B(_06163_));
 sg13g2_xnor2_1 _15571_ (.Y(_06585_),
    .A(_06569_),
    .B(_06584_));
 sg13g2_nor2_1 _15572_ (.A(net640),
    .B(_06585_),
    .Y(_06586_));
 sg13g2_nor4_1 _15573_ (.A(net107),
    .B(_06581_),
    .C(_06583_),
    .D(_06586_),
    .Y(_06587_));
 sg13g2_a22oi_1 _15574_ (.Y(_06588_),
    .B1(_06574_),
    .B2(_06587_),
    .A2(net75),
    .A1(net640));
 sg13g2_o21ai_1 _15575_ (.B1(_05679_),
    .Y(_06589_),
    .A1(net49),
    .A2(_06531_));
 sg13g2_a21oi_1 _15576_ (.A1(_06531_),
    .A2(_06588_),
    .Y(_00310_),
    .B1(_06589_));
 sg13g2_nor2_1 _15577_ (.A(_05844_),
    .B(_06188_),
    .Y(_06590_));
 sg13g2_o21ai_1 _15578_ (.B1(_05877_),
    .Y(_06591_),
    .A1(net331),
    .A2(_06188_));
 sg13g2_buf_1 _15579_ (.A(\grid.cell_13_2.se ),
    .X(_06592_));
 sg13g2_xnor2_1 _15580_ (.Y(_06593_),
    .A(_06592_),
    .B(_06185_));
 sg13g2_xnor2_1 _15581_ (.Y(_06594_),
    .A(_06539_),
    .B(_06593_));
 sg13g2_mux2_1 _15582_ (.A0(_06590_),
    .A1(_06591_),
    .S(_06594_),
    .X(_06595_));
 sg13g2_buf_1 _15583_ (.A(_06592_),
    .X(_06596_));
 sg13g2_buf_1 _15584_ (.A(net959),
    .X(_06597_));
 sg13g2_nand2_1 _15585_ (.Y(_06598_),
    .A(net623),
    .B(net635));
 sg13g2_o21ai_1 _15586_ (.B1(net625),
    .Y(_06599_),
    .A1(net623),
    .A2(net635));
 sg13g2_nand2_1 _15587_ (.Y(_06600_),
    .A(_06598_),
    .B(_06599_));
 sg13g2_xnor2_1 _15588_ (.Y(_06601_),
    .A(_06595_),
    .B(_06600_));
 sg13g2_xnor2_1 _15589_ (.Y(_06602_),
    .A(net981),
    .B(_05817_));
 sg13g2_xnor2_1 _15590_ (.Y(_06603_),
    .A(_06594_),
    .B(_06602_));
 sg13g2_nand2_1 _15591_ (.Y(_06604_),
    .A(_06224_),
    .B(_06603_));
 sg13g2_buf_1 _15592_ (.A(_00234_),
    .X(_06605_));
 sg13g2_inv_2 _15593_ (.Y(_06606_),
    .A(_06605_));
 sg13g2_nand2_1 _15594_ (.Y(_06607_),
    .A(_06606_),
    .B(_06092_));
 sg13g2_nor2_1 _15595_ (.A(_06595_),
    .B(_06600_),
    .Y(_06608_));
 sg13g2_o21ai_1 _15596_ (.B1(_06608_),
    .Y(_06609_),
    .A1(_06604_),
    .A2(_06607_));
 sg13g2_nor2_1 _15597_ (.A(net330),
    .B(_06606_),
    .Y(_06610_));
 sg13g2_xnor2_1 _15598_ (.Y(_06611_),
    .A(_06075_),
    .B(_06603_));
 sg13g2_a22oi_1 _15599_ (.Y(_06612_),
    .B1(_06224_),
    .B2(_06603_),
    .A2(_06606_),
    .A1(net330));
 sg13g2_o21ai_1 _15600_ (.B1(_06612_),
    .Y(_06613_),
    .A1(_06610_),
    .A2(_06611_));
 sg13g2_mux2_1 _15601_ (.A0(_06601_),
    .A1(_06609_),
    .S(_06613_),
    .X(_06614_));
 sg13g2_nand2_1 _15602_ (.Y(_06615_),
    .A(net82),
    .B(_06614_));
 sg13g2_xnor2_1 _15603_ (.Y(_06616_),
    .A(net628),
    .B(_06092_));
 sg13g2_xnor2_1 _15604_ (.Y(_06617_),
    .A(_06603_),
    .B(_06616_));
 sg13g2_a21oi_1 _15605_ (.A1(net113),
    .A2(_06617_),
    .Y(_06618_),
    .B1(net157));
 sg13g2_nor2_1 _15606_ (.A(net60),
    .B(_06618_),
    .Y(_06619_));
 sg13g2_a22oi_1 _15607_ (.Y(_06620_),
    .B1(_06615_),
    .B2(_06619_),
    .A2(_06476_),
    .A1(net33));
 sg13g2_nor2_1 _15608_ (.A(net370),
    .B(_06620_),
    .Y(_00311_));
 sg13g2_inv_2 _15609_ (.Y(_06621_),
    .A(net48));
 sg13g2_nand2_1 _15610_ (.Y(_06622_),
    .A(_06621_),
    .B(net60));
 sg13g2_nor2_1 _15611_ (.A(_06251_),
    .B(_06255_),
    .Y(_06623_));
 sg13g2_buf_1 _15612_ (.A(\grid.cell_13_3.se ),
    .X(_06624_));
 sg13g2_buf_1 _15613_ (.A(net1166),
    .X(_06625_));
 sg13g2_nor2_1 _15614_ (.A(net958),
    .B(_06597_),
    .Y(_06626_));
 sg13g2_nand2_1 _15615_ (.Y(_06627_),
    .A(_06596_),
    .B(_06250_));
 sg13g2_o21ai_1 _15616_ (.B1(_06627_),
    .Y(_06628_),
    .A1(_06255_),
    .A2(net645));
 sg13g2_a21oi_1 _15617_ (.A1(_06623_),
    .A2(_06626_),
    .Y(_06629_),
    .B1(_06628_));
 sg13g2_o21ai_1 _15618_ (.B1(net958),
    .Y(_06630_),
    .A1(_06597_),
    .A2(net966));
 sg13g2_and2_1 _15619_ (.A(_05916_),
    .B(_06630_),
    .X(_06631_));
 sg13g2_buf_1 _15620_ (.A(net958),
    .X(_06632_));
 sg13g2_buf_1 _15621_ (.A(net623),
    .X(_06633_));
 sg13g2_nor3_1 _15622_ (.A(net622),
    .B(_06633_),
    .C(net633),
    .Y(_06634_));
 sg13g2_a22oi_1 _15623_ (.Y(_06635_),
    .B1(_06634_),
    .B2(_05887_),
    .A2(_06631_),
    .A1(_06629_));
 sg13g2_buf_1 _15624_ (.A(_00233_),
    .X(_06636_));
 sg13g2_nand2_1 _15625_ (.Y(_06637_),
    .A(net325),
    .B(_06270_));
 sg13g2_xnor2_1 _15626_ (.Y(_06638_),
    .A(net1166),
    .B(_06596_));
 sg13g2_xnor2_1 _15627_ (.Y(_06639_),
    .A(_06265_),
    .B(_06638_));
 sg13g2_xnor2_1 _15628_ (.Y(_06640_),
    .A(net979),
    .B(_06639_));
 sg13g2_buf_2 _15629_ (.A(_06640_),
    .X(_06641_));
 sg13g2_nor2_1 _15630_ (.A(net325),
    .B(_06270_),
    .Y(_06642_));
 sg13g2_nand2_1 _15631_ (.Y(_06643_),
    .A(_05844_),
    .B(_06270_));
 sg13g2_a21oi_1 _15632_ (.A1(_06641_),
    .A2(_06643_),
    .Y(_06644_),
    .B1(net326));
 sg13g2_a221oi_1 _15633_ (.B2(_06642_),
    .C1(_06644_),
    .B1(_06641_),
    .A1(net160),
    .Y(_06645_),
    .A2(_06637_));
 sg13g2_and2_1 _15634_ (.A(_06270_),
    .B(_06641_),
    .X(_06646_));
 sg13g2_xnor2_1 _15635_ (.Y(_06647_),
    .A(net326),
    .B(_06641_));
 sg13g2_a22oi_1 _15636_ (.Y(_06648_),
    .B1(_06647_),
    .B2(net160),
    .A2(_06646_),
    .A1(_06636_));
 sg13g2_o21ai_1 _15637_ (.B1(_06648_),
    .Y(_06649_),
    .A1(_06636_),
    .A2(_06645_));
 sg13g2_nor3_1 _15638_ (.A(net166),
    .B(_06635_),
    .C(_06649_),
    .Y(_06650_));
 sg13g2_xor2_1 _15639_ (.B(_06641_),
    .A(_06567_),
    .X(_06651_));
 sg13g2_a21oi_1 _15640_ (.A1(net116),
    .A2(_06651_),
    .Y(_06652_),
    .B1(net324));
 sg13g2_inv_2 _15641_ (.Y(_06653_),
    .A(_06636_));
 sg13g2_o21ai_1 _15642_ (.B1(_06647_),
    .Y(_06654_),
    .A1(net160),
    .A2(_06653_));
 sg13g2_xor2_1 _15643_ (.B(_06250_),
    .A(net959),
    .X(_06655_));
 sg13g2_nand2_1 _15644_ (.Y(_06656_),
    .A(net979),
    .B(_06655_));
 sg13g2_o21ai_1 _15645_ (.B1(_06656_),
    .Y(_06657_),
    .A1(net645),
    .A2(_06627_));
 sg13g2_nor2_1 _15646_ (.A(_05916_),
    .B(_06627_),
    .Y(_06658_));
 sg13g2_a21oi_1 _15647_ (.A1(net978),
    .A2(_06657_),
    .Y(_06659_),
    .B1(_06658_));
 sg13g2_nand2b_1 _15648_ (.Y(_06660_),
    .B(net622),
    .A_N(_06659_));
 sg13g2_nor3_1 _15649_ (.A(net958),
    .B(_05887_),
    .C(_06627_),
    .Y(_06661_));
 sg13g2_a221oi_1 _15650_ (.B2(_06641_),
    .C1(_06661_),
    .B1(_06270_),
    .A1(net160),
    .Y(_06662_),
    .A2(_06653_));
 sg13g2_and2_1 _15651_ (.A(_06660_),
    .B(_06662_),
    .X(_06663_));
 sg13g2_nand2_1 _15652_ (.Y(_06664_),
    .A(net118),
    .B(_06635_));
 sg13g2_a21oi_1 _15653_ (.A1(_06654_),
    .A2(_06663_),
    .Y(_06665_),
    .B1(_06664_));
 sg13g2_or4_1 _15654_ (.A(net60),
    .B(_06650_),
    .C(_06652_),
    .D(_06665_),
    .X(_06666_));
 sg13g2_a21oi_1 _15655_ (.A1(_06622_),
    .A2(_06666_),
    .Y(_00312_),
    .B1(net350));
 sg13g2_buf_1 _15656_ (.A(net716),
    .X(_06667_));
 sg13g2_nand3_1 _15657_ (.B(_06425_),
    .C(_06531_),
    .A(net633),
    .Y(_06668_));
 sg13g2_o21ai_1 _15658_ (.B1(_06668_),
    .Y(_06669_),
    .A1(net47),
    .A2(_06531_));
 sg13g2_buf_2 _15659_ (.A(\grid.cell_13_4.se ),
    .X(_06670_));
 sg13g2_buf_1 _15660_ (.A(_06670_),
    .X(_06671_));
 sg13g2_buf_1 _15661_ (.A(net957),
    .X(_06672_));
 sg13g2_buf_1 _15662_ (.A(net621),
    .X(_06673_));
 sg13g2_nand2_1 _15663_ (.Y(_06674_),
    .A(net643),
    .B(net977));
 sg13g2_nor2_1 _15664_ (.A(net1166),
    .B(net965),
    .Y(_06675_));
 sg13g2_nand2_1 _15665_ (.Y(_06676_),
    .A(_06674_),
    .B(_06675_));
 sg13g2_inv_2 _15666_ (.Y(_06677_),
    .A(net957));
 sg13g2_nand3_1 _15667_ (.B(net643),
    .C(_06675_),
    .A(_06677_),
    .Y(_06678_));
 sg13g2_o21ai_1 _15668_ (.B1(net632),
    .Y(_06679_),
    .A1(_06672_),
    .A2(_06625_));
 sg13g2_and2_1 _15669_ (.A(net957),
    .B(net1166),
    .X(_06680_));
 sg13g2_buf_1 _15670_ (.A(_06680_),
    .X(_06681_));
 sg13g2_a21oi_1 _15671_ (.A1(net643),
    .A2(_06255_),
    .Y(_06682_),
    .B1(_06681_));
 sg13g2_nand4_1 _15672_ (.B(_06678_),
    .C(_06679_),
    .A(_05951_),
    .Y(_06683_),
    .D(_06682_));
 sg13g2_o21ai_1 _15673_ (.B1(_06683_),
    .Y(_06684_),
    .A1(net316),
    .A2(_06676_));
 sg13g2_o21ai_1 _15674_ (.B1(_06304_),
    .Y(_06685_),
    .A1(net635),
    .A2(_06188_));
 sg13g2_xnor2_1 _15675_ (.Y(_06686_),
    .A(_06670_),
    .B(_06291_));
 sg13g2_xnor2_1 _15676_ (.Y(_06687_),
    .A(_05901_),
    .B(_06686_));
 sg13g2_xnor2_1 _15677_ (.Y(_06688_),
    .A(net1172),
    .B(_06687_));
 sg13g2_xnor2_1 _15678_ (.Y(_06689_),
    .A(_06625_),
    .B(_06688_));
 sg13g2_mux2_1 _15679_ (.A0(_06189_),
    .A1(_06685_),
    .S(_06689_),
    .X(_06690_));
 sg13g2_buf_1 _15680_ (.A(_00047_),
    .X(_06691_));
 sg13g2_xnor2_1 _15681_ (.Y(_06692_),
    .A(_06624_),
    .B(net968));
 sg13g2_xnor2_1 _15682_ (.Y(_06693_),
    .A(_06188_),
    .B(_06692_));
 sg13g2_xnor2_1 _15683_ (.Y(_06694_),
    .A(_06688_),
    .B(_06693_));
 sg13g2_nor2_1 _15684_ (.A(_06691_),
    .B(_06694_),
    .Y(_06695_));
 sg13g2_xor2_1 _15685_ (.B(_06695_),
    .A(_06690_),
    .X(_06696_));
 sg13g2_nor3_1 _15686_ (.A(_06684_),
    .B(_06690_),
    .C(_06695_),
    .Y(_06697_));
 sg13g2_a21oi_1 _15687_ (.A1(_06684_),
    .A2(_06696_),
    .Y(_06698_),
    .B1(_06697_));
 sg13g2_inv_1 _15688_ (.Y(_06699_),
    .A(net1166));
 sg13g2_buf_1 _15689_ (.A(_06699_),
    .X(_06700_));
 sg13g2_nor2_1 _15690_ (.A(net620),
    .B(_06295_),
    .Y(_06701_));
 sg13g2_nand2b_1 _15691_ (.Y(_06702_),
    .B(_06701_),
    .A_N(_06674_));
 sg13g2_o21ai_1 _15692_ (.B1(net1002),
    .Y(_06703_),
    .A1(net316),
    .A2(_06702_));
 sg13g2_xnor2_1 _15693_ (.Y(_06704_),
    .A(net323),
    .B(net644));
 sg13g2_a21oi_1 _15694_ (.A1(net323),
    .A2(net644),
    .Y(_06705_),
    .B1(net622));
 sg13g2_a21oi_1 _15695_ (.A1(_06632_),
    .A2(_06704_),
    .Y(_06706_),
    .B1(_06705_));
 sg13g2_a22oi_1 _15696_ (.Y(_06707_),
    .B1(_06706_),
    .B2(net329),
    .A2(_06701_),
    .A1(_05952_));
 sg13g2_xnor2_1 _15697_ (.Y(_06708_),
    .A(_06190_),
    .B(_06638_));
 sg13g2_xnor2_1 _15698_ (.Y(_06709_),
    .A(_06688_),
    .B(_06708_));
 sg13g2_o21ai_1 _15699_ (.B1(_06254_),
    .Y(_06710_),
    .A1(_04614_),
    .A2(_06709_));
 sg13g2_o21ai_1 _15700_ (.B1(_06710_),
    .Y(_06711_),
    .A1(_06677_),
    .A2(_06707_));
 sg13g2_nor4_1 _15701_ (.A(net60),
    .B(_06698_),
    .C(_06703_),
    .D(_06711_),
    .Y(_06712_));
 sg13g2_a21o_1 _15702_ (.A2(_06669_),
    .A1(net317),
    .B1(_06712_),
    .X(_00313_));
 sg13g2_buf_1 _15703_ (.A(\grid.cell_13_5.se ),
    .X(_06713_));
 sg13g2_buf_1 _15704_ (.A(_06713_),
    .X(_06714_));
 sg13g2_xor2_1 _15705_ (.B(_06336_),
    .A(net957),
    .X(_06715_));
 sg13g2_xnor2_1 _15706_ (.Y(_06716_),
    .A(_05947_),
    .B(_06715_));
 sg13g2_xnor2_1 _15707_ (.Y(_06717_),
    .A(net956),
    .B(_06716_));
 sg13g2_buf_1 _15708_ (.A(_06717_),
    .X(_06718_));
 sg13g2_xnor2_1 _15709_ (.Y(_06719_),
    .A(net633),
    .B(_06718_));
 sg13g2_nor2_1 _15710_ (.A(_06332_),
    .B(_06718_),
    .Y(_06720_));
 sg13g2_buf_2 _15711_ (.A(_00079_),
    .X(_06721_));
 sg13g2_o21ai_1 _15712_ (.B1(_06255_),
    .Y(_06722_),
    .A1(_06282_),
    .A2(_06718_));
 sg13g2_nor2_1 _15713_ (.A(net1168),
    .B(net978),
    .Y(_06723_));
 sg13g2_or2_1 _15714_ (.X(_06724_),
    .B(_06723_),
    .A(_06718_));
 sg13g2_a221oi_1 _15715_ (.B2(_06282_),
    .C1(_06623_),
    .B1(_06724_),
    .A1(_06332_),
    .Y(_06725_),
    .A2(_06722_));
 sg13g2_nor2_1 _15716_ (.A(_06721_),
    .B(_06725_),
    .Y(_06726_));
 sg13g2_a221oi_1 _15717_ (.B2(_06721_),
    .C1(_06726_),
    .B1(_06720_),
    .A1(net644),
    .Y(_06727_),
    .A2(_06719_));
 sg13g2_buf_1 _15718_ (.A(_06714_),
    .X(_06728_));
 sg13g2_buf_1 _15719_ (.A(net619),
    .X(_06729_));
 sg13g2_nand2_1 _15720_ (.Y(_06730_),
    .A(_06677_),
    .B(net631));
 sg13g2_inv_1 _15721_ (.Y(_06731_),
    .A(_06713_));
 sg13g2_buf_1 _15722_ (.A(_06731_),
    .X(_06732_));
 sg13g2_nand2_1 _15723_ (.Y(_06733_),
    .A(net618),
    .B(net328));
 sg13g2_o21ai_1 _15724_ (.B1(net322),
    .Y(_06734_),
    .A1(net315),
    .A2(_06673_));
 sg13g2_o21ai_1 _15725_ (.B1(_06734_),
    .Y(_06735_),
    .A1(_06730_),
    .A2(_06733_));
 sg13g2_a221oi_1 _15726_ (.B2(_06296_),
    .C1(_06735_),
    .B1(net328),
    .A1(net315),
    .Y(_06736_),
    .A2(_06673_));
 sg13g2_nor2_1 _15727_ (.A(net619),
    .B(_06730_),
    .Y(_06737_));
 sg13g2_a22oi_1 _15728_ (.Y(_06738_),
    .B1(_06737_),
    .B2(_05961_),
    .A2(_06736_),
    .A1(net974));
 sg13g2_mux2_1 _15729_ (.A0(net630),
    .A1(net975),
    .S(net957),
    .X(_06739_));
 sg13g2_nand3_1 _15730_ (.B(net643),
    .C(_06739_),
    .A(net974),
    .Y(_06740_));
 sg13g2_o21ai_1 _15731_ (.B1(_06740_),
    .Y(_06741_),
    .A1(net643),
    .A2(_06730_));
 sg13g2_nand2_1 _15732_ (.Y(_06742_),
    .A(net618),
    .B(_06741_));
 sg13g2_inv_1 _15733_ (.Y(_06743_),
    .A(_06721_));
 sg13g2_and2_1 _15734_ (.A(net957),
    .B(net964),
    .X(_06744_));
 sg13g2_buf_1 _15735_ (.A(_06744_),
    .X(_06745_));
 sg13g2_nor3_1 _15736_ (.A(_05984_),
    .B(_06671_),
    .C(net630),
    .Y(_06746_));
 sg13g2_a22oi_1 _15737_ (.Y(_06747_),
    .B1(_05937_),
    .B2(net976),
    .A2(net630),
    .A1(_06671_));
 sg13g2_or2_1 _15738_ (.X(_06748_),
    .B(_06747_),
    .A(_06746_));
 sg13g2_a21oi_1 _15739_ (.A1(net974),
    .A2(_06745_),
    .Y(_06749_),
    .B1(_06748_));
 sg13g2_mux2_1 _15740_ (.A0(_05984_),
    .A1(_06731_),
    .S(_06296_),
    .X(_06750_));
 sg13g2_nand2_1 _15741_ (.Y(_06751_),
    .A(net642),
    .B(_06745_));
 sg13g2_nor2_1 _15742_ (.A(_06750_),
    .B(_06751_),
    .Y(_06752_));
 sg13g2_a221oi_1 _15743_ (.B2(net315),
    .C1(_06752_),
    .B1(_06749_),
    .A1(_06743_),
    .Y(_06753_),
    .A2(net644));
 sg13g2_nand2_1 _15744_ (.Y(_06754_),
    .A(_06742_),
    .B(_06753_));
 sg13g2_o21ai_1 _15745_ (.B1(_06730_),
    .Y(_06755_),
    .A1(_06728_),
    .A2(_06745_));
 sg13g2_a21oi_1 _15746_ (.A1(net974),
    .A2(_06755_),
    .Y(_06756_),
    .B1(_06737_));
 sg13g2_nor2_1 _15747_ (.A(net328),
    .B(_06756_),
    .Y(_06757_));
 sg13g2_nor3_1 _15748_ (.A(_06720_),
    .B(_06754_),
    .C(_06757_),
    .Y(_06758_));
 sg13g2_o21ai_1 _15749_ (.B1(_06719_),
    .Y(_06759_),
    .A1(_06743_),
    .A2(net644));
 sg13g2_a221oi_1 _15750_ (.B2(_06759_),
    .C1(net115),
    .B1(_06758_),
    .A1(net108),
    .Y(_06760_),
    .A2(_06530_));
 sg13g2_o21ai_1 _15751_ (.B1(_06760_),
    .Y(_06761_),
    .A1(_06727_),
    .A2(_06738_));
 sg13g2_buf_1 _15752_ (.A(_05002_),
    .X(_06762_));
 sg13g2_xnor2_1 _15753_ (.Y(_06763_),
    .A(_06632_),
    .B(_06265_));
 sg13g2_xnor2_1 _15754_ (.Y(_06764_),
    .A(_06718_),
    .B(_06763_));
 sg13g2_a221oi_1 _15755_ (.B2(net111),
    .C1(net323),
    .B1(_06764_),
    .A1(net108),
    .Y(_06765_),
    .A2(_06530_));
 sg13g2_a21oi_1 _15756_ (.A1(net43),
    .A2(net60),
    .Y(_06766_),
    .B1(_06765_));
 sg13g2_and3_1 _15757_ (.X(_00314_),
    .A(net317),
    .B(_06761_),
    .C(_06766_));
 sg13g2_buf_2 _15758_ (.A(_00141_),
    .X(_06767_));
 sg13g2_o21ai_1 _15759_ (.B1(_06005_),
    .Y(_06768_),
    .A1(_06767_),
    .A2(_06486_));
 sg13g2_nand2b_1 _15760_ (.Y(_06769_),
    .B(_06491_),
    .A_N(_06767_));
 sg13g2_o21ai_1 _15761_ (.B1(_06769_),
    .Y(_06770_),
    .A1(_06491_),
    .A2(_06768_));
 sg13g2_o21ai_1 _15762_ (.B1(_06486_),
    .Y(_06771_),
    .A1(net619),
    .A2(_06491_));
 sg13g2_nor2_1 _15763_ (.A(net956),
    .B(_06486_),
    .Y(_06772_));
 sg13g2_a21oi_1 _15764_ (.A1(_06767_),
    .A2(_06771_),
    .Y(_06773_),
    .B1(_06772_));
 sg13g2_and2_1 _15765_ (.A(net956),
    .B(net627),
    .X(_06774_));
 sg13g2_a21oi_1 _15766_ (.A1(_06080_),
    .A2(_06774_),
    .Y(_06775_),
    .B1(_06772_));
 sg13g2_nor2b_1 _15767_ (.A(_06767_),
    .B_N(net627),
    .Y(_06776_));
 sg13g2_nand2b_1 _15768_ (.Y(_06777_),
    .B(net639),
    .A_N(net962));
 sg13g2_nand2_1 _15769_ (.Y(_06778_),
    .A(_06507_),
    .B(net647));
 sg13g2_a21oi_1 _15770_ (.A1(_06777_),
    .A2(_06778_),
    .Y(_06779_),
    .B1(_06714_));
 sg13g2_a22oi_1 _15771_ (.Y(_06780_),
    .B1(_06779_),
    .B2(_06767_),
    .A2(_06776_),
    .A1(_06080_));
 sg13g2_mux2_1 _15772_ (.A0(_06775_),
    .A1(_06780_),
    .S(net642),
    .X(_06781_));
 sg13g2_o21ai_1 _15773_ (.B1(_06781_),
    .Y(_06782_),
    .A1(net161),
    .A2(_06773_));
 sg13g2_a21oi_1 _15774_ (.A1(net315),
    .A2(_06770_),
    .Y(_06783_),
    .B1(_06782_));
 sg13g2_buf_1 _15775_ (.A(_00111_),
    .X(_06784_));
 sg13g2_inv_1 _15776_ (.Y(_06785_),
    .A(_06784_));
 sg13g2_xnor2_1 _15777_ (.Y(_06786_),
    .A(_06713_),
    .B(_06479_));
 sg13g2_xnor2_1 _15778_ (.Y(_06787_),
    .A(_06039_),
    .B(_06786_));
 sg13g2_xnor2_1 _15779_ (.Y(_06788_),
    .A(net629),
    .B(_06787_));
 sg13g2_xnor2_1 _15780_ (.Y(_06789_),
    .A(_06295_),
    .B(_06788_));
 sg13g2_o21ai_1 _15781_ (.B1(_06789_),
    .Y(_06790_),
    .A1(_06785_),
    .A2(net329));
 sg13g2_nor2b_1 _15782_ (.A(_06392_),
    .B_N(_06788_),
    .Y(_06791_));
 sg13g2_a21oi_1 _15783_ (.A1(_06785_),
    .A2(net329),
    .Y(_06792_),
    .B1(_06791_));
 sg13g2_nand2_1 _15784_ (.Y(_06793_),
    .A(_06790_),
    .B(_06792_));
 sg13g2_xnor2_1 _15785_ (.Y(_06794_),
    .A(_06783_),
    .B(_06793_));
 sg13g2_xor2_1 _15786_ (.B(_06788_),
    .A(_06687_),
    .X(_06795_));
 sg13g2_buf_1 _15787_ (.A(net627),
    .X(_06796_));
 sg13g2_buf_1 _15788_ (.A(_06796_),
    .X(_06797_));
 sg13g2_nand2b_1 _15789_ (.Y(_06798_),
    .B(net629),
    .A_N(net975));
 sg13g2_nand3b_1 _15790_ (.B(_06798_),
    .C(net314),
    .Y(_06799_),
    .A_N(_06441_));
 sg13g2_o21ai_1 _15791_ (.B1(_06799_),
    .Y(_06800_),
    .A1(_06797_),
    .A2(_06432_));
 sg13g2_o21ai_1 _15792_ (.B1(_06769_),
    .Y(_06801_),
    .A1(_05715_),
    .A2(_06800_));
 sg13g2_xor2_1 _15793_ (.B(net329),
    .A(net632),
    .X(_06802_));
 sg13g2_nor2_1 _15794_ (.A(_06784_),
    .B(_06802_),
    .Y(_06803_));
 sg13g2_nand3_1 _15795_ (.B(_06005_),
    .C(_06491_),
    .A(_06732_),
    .Y(_06804_));
 sg13g2_nand2_1 _15796_ (.Y(_06805_),
    .A(_02765_),
    .B(_06804_));
 sg13g2_a221oi_1 _15797_ (.B2(_06791_),
    .C1(_06805_),
    .B1(_06803_),
    .A1(_06729_),
    .Y(_06806_),
    .A2(_06801_));
 sg13g2_o21ai_1 _15798_ (.B1(_06806_),
    .Y(_06807_),
    .A1(net322),
    .A2(_06795_));
 sg13g2_or2_1 _15799_ (.X(_06808_),
    .B(_06807_),
    .A(_06794_));
 sg13g2_and2_1 _15800_ (.A(net158),
    .B(_05118_),
    .X(_06809_));
 sg13g2_buf_2 _15801_ (.A(_06809_),
    .X(_06810_));
 sg13g2_a22oi_1 _15802_ (.Y(_06811_),
    .B1(_06530_),
    .B2(_06810_),
    .A2(net103),
    .A1(net322));
 sg13g2_nor2_1 _15803_ (.A(net176),
    .B(_05119_),
    .Y(_06812_));
 sg13g2_buf_2 _15804_ (.A(_06812_),
    .X(_06813_));
 sg13g2_buf_1 _15805_ (.A(_06813_),
    .X(_06814_));
 sg13g2_buf_1 _15806_ (.A(_06110_),
    .X(_06815_));
 sg13g2_a221oi_1 _15807_ (.B2(_06530_),
    .C1(_06815_),
    .B1(net24),
    .A1(_06808_),
    .Y(_00315_),
    .A2(_06811_));
 sg13g2_nand2_1 _15808_ (.Y(_06816_),
    .A(net80),
    .B(net60));
 sg13g2_buf_1 _15809_ (.A(net105),
    .X(_06817_));
 sg13g2_xnor2_1 _15810_ (.Y(_06818_),
    .A(net964),
    .B(_06786_));
 sg13g2_xor2_1 _15811_ (.B(_06818_),
    .A(_06039_),
    .X(_06819_));
 sg13g2_xnor2_1 _15812_ (.Y(_06820_),
    .A(net971),
    .B(_06819_));
 sg13g2_o21ai_1 _15813_ (.B1(_06571_),
    .Y(_06821_),
    .A1(net970),
    .A2(_06819_));
 sg13g2_a21oi_1 _15814_ (.A1(_06565_),
    .A2(_06820_),
    .Y(_06822_),
    .B1(_06821_));
 sg13g2_nand2_1 _15815_ (.Y(_06823_),
    .A(net314),
    .B(net630));
 sg13g2_o21ai_1 _15816_ (.B1(net315),
    .Y(_06824_),
    .A1(net314),
    .A2(net630));
 sg13g2_nand2_1 _15817_ (.Y(_06825_),
    .A(_06823_),
    .B(_06824_));
 sg13g2_o21ai_1 _15818_ (.B1(_06767_),
    .Y(_06826_),
    .A1(net642),
    .A2(_05715_));
 sg13g2_mux2_1 _15819_ (.A0(_06005_),
    .A1(_06826_),
    .S(_06818_),
    .X(_06827_));
 sg13g2_xnor2_1 _15820_ (.Y(_06828_),
    .A(_06825_),
    .B(_06827_));
 sg13g2_nor4_1 _15821_ (.A(_06511_),
    .B(net970),
    .C(_06582_),
    .D(_06819_),
    .Y(_06829_));
 sg13g2_nor3_1 _15822_ (.A(_06825_),
    .B(_06829_),
    .C(_06827_),
    .Y(_06830_));
 sg13g2_nor2_1 _15823_ (.A(_06822_),
    .B(_06830_),
    .Y(_06831_));
 sg13g2_a21oi_1 _15824_ (.A1(_06822_),
    .A2(_06828_),
    .Y(_06832_),
    .B1(_06831_));
 sg13g2_xnor2_1 _15825_ (.Y(_06833_),
    .A(_06584_),
    .B(_06819_));
 sg13g2_a21oi_1 _15826_ (.A1(net116),
    .A2(_06833_),
    .Y(_06834_),
    .B1(_06457_));
 sg13g2_nor2_1 _15827_ (.A(net60),
    .B(_06834_),
    .Y(_06835_));
 sg13g2_o21ai_1 _15828_ (.B1(_06835_),
    .Y(_06836_),
    .A1(net74),
    .A2(_06832_));
 sg13g2_a21oi_1 _15829_ (.A1(_06816_),
    .A2(_06836_),
    .Y(_00316_),
    .B1(net350));
 sg13g2_buf_1 _15830_ (.A(\grid.cell_14_0.se ),
    .X(_06837_));
 sg13g2_inv_1 _15831_ (.Y(_06838_),
    .A(net1165));
 sg13g2_buf_1 _15832_ (.A(_06838_),
    .X(_06839_));
 sg13g2_buf_1 _15833_ (.A(\grid.cell_14_0.sw ),
    .X(_06840_));
 sg13g2_buf_1 _15834_ (.A(_06840_),
    .X(_06841_));
 sg13g2_and2_1 _15835_ (.A(_06841_),
    .B(_06479_),
    .X(_06842_));
 sg13g2_buf_1 _15836_ (.A(_06842_),
    .X(_06843_));
 sg13g2_buf_1 _15837_ (.A(_06843_),
    .X(_06844_));
 sg13g2_xnor2_1 _15838_ (.Y(_06845_),
    .A(net955),
    .B(_06479_));
 sg13g2_nor2_1 _15839_ (.A(_06128_),
    .B(_06845_),
    .Y(_06846_));
 sg13g2_a21o_1 _15840_ (.A2(net155),
    .A1(_06128_),
    .B1(_06846_),
    .X(_06847_));
 sg13g2_a22oi_1 _15841_ (.Y(_06848_),
    .B1(_06847_),
    .B2(net321),
    .A2(net155),
    .A1(_06224_));
 sg13g2_buf_1 _15842_ (.A(net1165),
    .X(_06849_));
 sg13g2_nor2_1 _15843_ (.A(_06128_),
    .B(_06849_),
    .Y(_06850_));
 sg13g2_nand3_1 _15844_ (.B(net155),
    .C(_06850_),
    .A(net321),
    .Y(_06851_));
 sg13g2_o21ai_1 _15845_ (.B1(_06851_),
    .Y(_06852_),
    .A1(net616),
    .A2(_06848_));
 sg13g2_nor2_1 _15846_ (.A(_05185_),
    .B(net159),
    .Y(_06853_));
 sg13g2_nand2_2 _15847_ (.Y(_06854_),
    .A(net158),
    .B(_06853_));
 sg13g2_nand2_1 _15848_ (.Y(_06855_),
    .A(net1054),
    .B(_06854_));
 sg13g2_buf_2 _15849_ (.A(\grid.cell_14_0.s ),
    .X(_06856_));
 sg13g2_buf_1 _15850_ (.A(_06856_),
    .X(_06857_));
 sg13g2_xor2_1 _15851_ (.B(net1165),
    .A(_06066_),
    .X(_06858_));
 sg13g2_buf_1 _15852_ (.A(net955),
    .X(_06859_));
 sg13g2_xnor2_1 _15853_ (.Y(_06860_),
    .A(_06095_),
    .B(net615));
 sg13g2_xnor2_1 _15854_ (.Y(_06861_),
    .A(_06858_),
    .B(_06860_));
 sg13g2_xnor2_1 _15855_ (.Y(_06862_),
    .A(_06482_),
    .B(_06861_));
 sg13g2_xnor2_1 _15856_ (.Y(_06863_),
    .A(net953),
    .B(_06862_));
 sg13g2_a21oi_1 _15857_ (.A1(net126),
    .A2(_06863_),
    .Y(_06864_),
    .B1(_06533_));
 sg13g2_nor3_1 _15858_ (.A(_06852_),
    .B(_06855_),
    .C(_06864_),
    .Y(_06865_));
 sg13g2_xnor2_1 _15859_ (.Y(_06866_),
    .A(_06068_),
    .B(_06845_));
 sg13g2_xnor2_1 _15860_ (.Y(_06867_),
    .A(_06837_),
    .B(_06866_));
 sg13g2_xnor2_1 _15861_ (.Y(_06868_),
    .A(net628),
    .B(_06867_));
 sg13g2_a22oi_1 _15862_ (.Y(_06869_),
    .B1(_06868_),
    .B2(_06096_),
    .A2(_06867_),
    .A1(_06606_));
 sg13g2_buf_1 _15863_ (.A(net955),
    .X(_06870_));
 sg13g2_nand2b_1 _15864_ (.Y(_06871_),
    .B(net627),
    .A_N(net614));
 sg13g2_nand2b_1 _15865_ (.Y(_06872_),
    .B(net962),
    .A_N(_06199_));
 sg13g2_nand2_1 _15866_ (.Y(_06873_),
    .A(net615),
    .B(_06872_));
 sg13g2_a21oi_1 _15867_ (.A1(_06871_),
    .A2(_06873_),
    .Y(_06874_),
    .B1(net629));
 sg13g2_nand2b_1 _15868_ (.Y(_06875_),
    .B(net614),
    .A_N(net627));
 sg13g2_nand2b_1 _15869_ (.Y(_06876_),
    .B(net629),
    .A_N(net614));
 sg13g2_a21oi_1 _15870_ (.A1(_06875_),
    .A2(_06876_),
    .Y(_06877_),
    .B1(net973));
 sg13g2_or2_1 _15871_ (.X(_06878_),
    .B(net962),
    .A(_06841_));
 sg13g2_buf_1 _15872_ (.A(_06878_),
    .X(_06879_));
 sg13g2_nor2_1 _15873_ (.A(net967),
    .B(_06879_),
    .Y(_06880_));
 sg13g2_nor4_1 _15874_ (.A(net616),
    .B(_06874_),
    .C(_06877_),
    .D(_06880_),
    .Y(_06881_));
 sg13g2_nor2b_1 _15875_ (.A(net973),
    .B_N(net639),
    .Y(_06882_));
 sg13g2_o21ai_1 _15876_ (.B1(_06500_),
    .Y(_06883_),
    .A1(_06507_),
    .A2(_06199_));
 sg13g2_nor2_1 _15877_ (.A(net615),
    .B(_06872_),
    .Y(_06884_));
 sg13g2_a221oi_1 _15878_ (.B2(net615),
    .C1(_06884_),
    .B1(_06883_),
    .A1(_06882_),
    .Y(_06885_),
    .A2(_06879_));
 sg13g2_and2_1 _15879_ (.A(net616),
    .B(_06885_),
    .X(_06886_));
 sg13g2_and3_1 _15880_ (.X(_06887_),
    .A(net1165),
    .B(net967),
    .C(_06843_));
 sg13g2_buf_1 _15881_ (.A(net614),
    .X(_06888_));
 sg13g2_nor3_1 _15882_ (.A(net954),
    .B(net313),
    .C(_06777_),
    .Y(_06889_));
 sg13g2_o21ai_1 _15883_ (.B1(net640),
    .Y(_06890_),
    .A1(_06887_),
    .A2(_06889_));
 sg13g2_o21ai_1 _15884_ (.B1(_06890_),
    .Y(_06891_),
    .A1(_06881_),
    .A2(_06886_));
 sg13g2_xnor2_1 _15885_ (.Y(_06892_),
    .A(_06869_),
    .B(_06891_));
 sg13g2_a221oi_1 _15886_ (.B2(_06096_),
    .C1(_06891_),
    .B1(_06868_),
    .A1(_06606_),
    .Y(_06893_),
    .A2(_06867_));
 sg13g2_buf_1 _15887_ (.A(_00232_),
    .X(_06894_));
 sg13g2_nor2_1 _15888_ (.A(_06894_),
    .B(_06862_),
    .Y(_06895_));
 sg13g2_mux2_1 _15889_ (.A0(_06892_),
    .A1(_06893_),
    .S(_06895_),
    .X(_06896_));
 sg13g2_buf_1 _15890_ (.A(_05407_),
    .X(_06897_));
 sg13g2_nand3_1 _15891_ (.B(net102),
    .C(_06854_),
    .A(net961),
    .Y(_06898_));
 sg13g2_o21ai_1 _15892_ (.B1(_06898_),
    .Y(_06899_),
    .A1(net50),
    .A2(_06854_));
 sg13g2_buf_2 _15893_ (.A(net714),
    .X(_06900_));
 sg13g2_a22oi_1 _15894_ (.Y(_06901_),
    .B1(_06899_),
    .B2(_06900_),
    .A2(_06896_),
    .A1(_06865_));
 sg13g2_inv_1 _15895_ (.Y(_00317_),
    .A(_06901_));
 sg13g2_buf_1 _15896_ (.A(\grid.cell_14_1.se ),
    .X(_06902_));
 sg13g2_buf_1 _15897_ (.A(net1164),
    .X(_06903_));
 sg13g2_buf_1 _15898_ (.A(_06903_),
    .X(_06904_));
 sg13g2_buf_1 _15899_ (.A(net613),
    .X(_06905_));
 sg13g2_nand4_1 _15900_ (.B(net626),
    .C(net311),
    .A(net157),
    .Y(_06906_),
    .D(_06850_));
 sg13g2_xnor2_1 _15901_ (.Y(_06907_),
    .A(_06539_),
    .B(net1164));
 sg13g2_nand2_1 _15902_ (.Y(_06908_),
    .A(net960),
    .B(net952));
 sg13g2_mux2_1 _15903_ (.A0(_06907_),
    .A1(_06908_),
    .S(_06128_),
    .X(_06909_));
 sg13g2_nor2_1 _15904_ (.A(net326),
    .B(_06909_),
    .Y(_06910_));
 sg13g2_nor2_1 _15905_ (.A(net967),
    .B(_06908_),
    .Y(_06911_));
 sg13g2_buf_1 _15906_ (.A(_06849_),
    .X(_06912_));
 sg13g2_o21ai_1 _15907_ (.B1(net612),
    .Y(_06913_),
    .A1(_06910_),
    .A2(_06911_));
 sg13g2_inv_1 _15908_ (.Y(_06914_),
    .A(net1164));
 sg13g2_xnor2_1 _15909_ (.Y(_06915_),
    .A(net951),
    .B(_06566_));
 sg13g2_xnor2_1 _15910_ (.Y(_06916_),
    .A(_06858_),
    .B(_06915_));
 sg13g2_xor2_1 _15911_ (.B(net1167),
    .A(_06095_),
    .X(_06917_));
 sg13g2_nor2_1 _15912_ (.A(_06894_),
    .B(_06917_),
    .Y(_06918_));
 sg13g2_nand3_1 _15913_ (.B(_06916_),
    .C(_06918_),
    .A(_06512_),
    .Y(_06919_));
 sg13g2_nand4_1 _15914_ (.B(_06906_),
    .C(_06913_),
    .A(net171),
    .Y(_06920_),
    .D(_06919_));
 sg13g2_inv_1 _15915_ (.Y(_06921_),
    .A(_06894_));
 sg13g2_nor2_1 _15916_ (.A(net971),
    .B(_06921_),
    .Y(_06922_));
 sg13g2_xnor2_1 _15917_ (.Y(_06923_),
    .A(net1167),
    .B(_06916_));
 sg13g2_a22oi_1 _15918_ (.Y(_06924_),
    .B1(_06512_),
    .B2(_06916_),
    .A2(_06921_),
    .A1(net971));
 sg13g2_o21ai_1 _15919_ (.B1(_06924_),
    .Y(_06925_),
    .A1(_06922_),
    .A2(_06923_));
 sg13g2_nand3_1 _15920_ (.B(_06542_),
    .C(net951),
    .A(net616),
    .Y(_06926_));
 sg13g2_nand4_1 _15921_ (.B(net636),
    .C(net960),
    .A(net1165),
    .Y(_06927_),
    .D(net952));
 sg13g2_a21oi_1 _15922_ (.A1(_06926_),
    .A2(_06927_),
    .Y(_06928_),
    .B1(net640));
 sg13g2_nor4_1 _15923_ (.A(net325),
    .B(_06548_),
    .C(_06904_),
    .D(_06224_),
    .Y(_06929_));
 sg13g2_nand2_1 _15924_ (.Y(_06930_),
    .A(net973),
    .B(net969));
 sg13g2_nand2b_1 _15925_ (.Y(_06931_),
    .B(net1164),
    .A_N(_06199_));
 sg13g2_o21ai_1 _15926_ (.B1(_06931_),
    .Y(_06932_),
    .A1(net952),
    .A2(_06930_));
 sg13g2_nor2_1 _15927_ (.A(net952),
    .B(_06199_),
    .Y(_06933_));
 sg13g2_nor3_1 _15928_ (.A(net960),
    .B(_06930_),
    .C(_06933_),
    .Y(_06934_));
 sg13g2_a21oi_1 _15929_ (.A1(_06548_),
    .A2(_06932_),
    .Y(_06935_),
    .B1(_06934_));
 sg13g2_nor2_1 _15930_ (.A(_06839_),
    .B(_06935_),
    .Y(_06936_));
 sg13g2_nor2b_1 _15931_ (.A(net1164),
    .B_N(_06199_),
    .Y(_06937_));
 sg13g2_a21oi_1 _15932_ (.A1(_06541_),
    .A2(_06931_),
    .Y(_06938_),
    .B1(_06937_));
 sg13g2_nand2_1 _15933_ (.Y(_06939_),
    .A(_06902_),
    .B(_06199_));
 sg13g2_o21ai_1 _15934_ (.B1(_06540_),
    .Y(_06940_),
    .A1(_06902_),
    .A2(_06199_));
 sg13g2_a21o_1 _15935_ (.A2(_06940_),
    .A1(_06939_),
    .B1(_06930_),
    .X(_06941_));
 sg13g2_o21ai_1 _15936_ (.B1(_06941_),
    .Y(_06942_),
    .A1(net636),
    .A2(_06938_));
 sg13g2_and2_1 _15937_ (.A(_06839_),
    .B(_06942_),
    .X(_06943_));
 sg13g2_nor4_1 _15938_ (.A(_06928_),
    .B(_06929_),
    .C(_06936_),
    .D(_06943_),
    .Y(_06944_));
 sg13g2_xnor2_1 _15939_ (.Y(_06945_),
    .A(_06925_),
    .B(_06944_));
 sg13g2_xor2_1 _15940_ (.B(_06917_),
    .A(_06857_),
    .X(_06946_));
 sg13g2_xnor2_1 _15941_ (.Y(_06947_),
    .A(_06916_),
    .B(_06946_));
 sg13g2_nor3_1 _15942_ (.A(_06920_),
    .B(_06945_),
    .C(_06947_),
    .Y(_06948_));
 sg13g2_o21ai_1 _15943_ (.B1(_02787_),
    .Y(_06949_),
    .A1(_06920_),
    .A2(_06945_));
 sg13g2_o21ai_1 _15944_ (.B1(_06949_),
    .Y(_06950_),
    .A1(_06556_),
    .A2(_06948_));
 sg13g2_o21ai_1 _15945_ (.B1(_05679_),
    .Y(_06951_),
    .A1(_03164_),
    .A2(_06854_));
 sg13g2_a21oi_1 _15946_ (.A1(_06854_),
    .A2(_06950_),
    .Y(_00318_),
    .B1(_06951_));
 sg13g2_nor3_1 _15947_ (.A(net375),
    .B(_05185_),
    .C(net159),
    .Y(_06952_));
 sg13g2_buf_1 _15948_ (.A(_06952_),
    .X(_06953_));
 sg13g2_nand2_1 _15949_ (.Y(_06954_),
    .A(net716),
    .B(_06953_));
 sg13g2_buf_2 _15950_ (.A(\grid.cell_14_2.se ),
    .X(_06955_));
 sg13g2_buf_1 _15951_ (.A(_06955_),
    .X(_06956_));
 sg13g2_inv_2 _15952_ (.Y(_06957_),
    .A(net950));
 sg13g2_inv_2 _15953_ (.Y(_06958_),
    .A(net959));
 sg13g2_nor2_1 _15954_ (.A(_06957_),
    .B(_06958_),
    .Y(_06959_));
 sg13g2_nor2b_1 _15955_ (.A(net959),
    .B_N(net950),
    .Y(_06960_));
 sg13g2_nor2b_1 _15956_ (.A(net950),
    .B_N(net959),
    .Y(_06961_));
 sg13g2_o21ai_1 _15957_ (.B1(net636),
    .Y(_06962_),
    .A1(_06960_),
    .A2(_06961_));
 sg13g2_o21ai_1 _15958_ (.B1(_06962_),
    .Y(_06963_),
    .A1(net635),
    .A2(_06959_));
 sg13g2_nand2_1 _15959_ (.Y(_06964_),
    .A(net325),
    .B(net635));
 sg13g2_buf_1 _15960_ (.A(net950),
    .X(_06965_));
 sg13g2_nor2_1 _15961_ (.A(_06965_),
    .B(net623),
    .Y(_06966_));
 sg13g2_a22oi_1 _15962_ (.Y(_06967_),
    .B1(_06964_),
    .B2(_06966_),
    .A2(_06963_),
    .A1(_06263_));
 sg13g2_o21ai_1 _15963_ (.B1(net324),
    .Y(_06968_),
    .A1(net326),
    .A2(_06914_));
 sg13g2_nand3_1 _15964_ (.B(_06968_),
    .C(_06966_),
    .A(_06263_),
    .Y(_06969_));
 sg13g2_o21ai_1 _15965_ (.B1(_06969_),
    .Y(_06970_),
    .A1(net311),
    .A2(_06967_));
 sg13g2_buf_1 _15966_ (.A(_00231_),
    .X(_06971_));
 sg13g2_buf_1 _15967_ (.A(_06971_),
    .X(_06972_));
 sg13g2_nand2_1 _15968_ (.Y(_06973_),
    .A(_06128_),
    .B(net949));
 sg13g2_xor2_1 _15969_ (.B(net1164),
    .A(net969),
    .X(_06974_));
 sg13g2_xnor2_1 _15970_ (.Y(_06975_),
    .A(_06955_),
    .B(_06593_));
 sg13g2_xnor2_1 _15971_ (.Y(_06976_),
    .A(_06974_),
    .B(_06975_));
 sg13g2_xnor2_1 _15972_ (.Y(_06977_),
    .A(net963),
    .B(_06976_));
 sg13g2_buf_1 _15973_ (.A(_06605_),
    .X(_06978_));
 sg13g2_inv_2 _15974_ (.Y(_06979_),
    .A(_06971_));
 sg13g2_nand2_1 _15975_ (.Y(_06980_),
    .A(net640),
    .B(_06979_));
 sg13g2_o21ai_1 _15976_ (.B1(_06980_),
    .Y(_06981_),
    .A1(net948),
    .A2(_06976_));
 sg13g2_a21oi_1 _15977_ (.A1(_06973_),
    .A2(_06977_),
    .Y(_06982_),
    .B1(_06981_));
 sg13g2_xor2_1 _15978_ (.B(_06982_),
    .A(_06970_),
    .X(_06983_));
 sg13g2_nand2_1 _15979_ (.Y(_06984_),
    .A(_06956_),
    .B(net623));
 sg13g2_o21ai_1 _15980_ (.B1(_06962_),
    .Y(_06985_),
    .A1(net325),
    .A2(_06984_));
 sg13g2_nand2_1 _15981_ (.Y(_06986_),
    .A(net324),
    .B(_06985_));
 sg13g2_o21ai_1 _15982_ (.B1(_06986_),
    .Y(_06987_),
    .A1(_06263_),
    .A2(_06984_));
 sg13g2_nor3_1 _15983_ (.A(net326),
    .B(net311),
    .C(_06598_),
    .Y(_06988_));
 sg13g2_buf_1 _15984_ (.A(net611),
    .X(_06989_));
 sg13g2_xor2_1 _15985_ (.B(net963),
    .A(net640),
    .X(_06990_));
 sg13g2_nor4_1 _15986_ (.A(net949),
    .B(net948),
    .C(_06990_),
    .D(_06976_),
    .Y(_06991_));
 sg13g2_a221oi_1 _15987_ (.B2(net310),
    .C1(_06991_),
    .B1(_06988_),
    .A1(_06905_),
    .Y(_06992_),
    .A2(_06987_));
 sg13g2_buf_1 _15988_ (.A(net168),
    .X(_06993_));
 sg13g2_a21oi_1 _15989_ (.A1(_06983_),
    .A2(_06992_),
    .Y(_06994_),
    .B1(net101));
 sg13g2_xor2_1 _15990_ (.B(_06977_),
    .A(_06858_),
    .X(_06995_));
 sg13g2_a21oi_1 _15991_ (.A1(net77),
    .A2(_06995_),
    .Y(_06996_),
    .B1(net626));
 sg13g2_or3_1 _15992_ (.A(_06855_),
    .B(_06994_),
    .C(_06996_),
    .X(_06997_));
 sg13g2_o21ai_1 _15993_ (.B1(_06997_),
    .Y(_00319_),
    .A1(net27),
    .A2(_06954_));
 sg13g2_buf_1 _15994_ (.A(\grid.cell_14_3.se ),
    .X(_06998_));
 sg13g2_inv_2 _15995_ (.Y(_06999_),
    .A(net1163));
 sg13g2_nor2_1 _15996_ (.A(_06957_),
    .B(_06700_),
    .Y(_07000_));
 sg13g2_nand2b_1 _15997_ (.Y(_07001_),
    .B(_07000_),
    .A_N(_06257_));
 sg13g2_nand3_1 _15998_ (.B(net622),
    .C(net324),
    .A(_06957_),
    .Y(_07002_));
 sg13g2_o21ai_1 _15999_ (.B1(_07002_),
    .Y(_07003_),
    .A1(_06957_),
    .A2(_06692_));
 sg13g2_a221oi_1 _16000_ (.B2(net633),
    .C1(_06999_),
    .B1(_07003_),
    .A1(_06310_),
    .Y(_07004_),
    .A2(_07000_));
 sg13g2_a21oi_1 _16001_ (.A1(_06999_),
    .A2(_07001_),
    .Y(_07005_),
    .B1(_07004_));
 sg13g2_xnor2_1 _16002_ (.Y(_07006_),
    .A(_06998_),
    .B(net1166));
 sg13g2_xnor2_1 _16003_ (.Y(_07007_),
    .A(_06539_),
    .B(net968));
 sg13g2_xnor2_1 _16004_ (.Y(_07008_),
    .A(_06955_),
    .B(net1169));
 sg13g2_xnor2_1 _16005_ (.Y(_07009_),
    .A(_07007_),
    .B(_07008_));
 sg13g2_xnor2_1 _16006_ (.Y(_07010_),
    .A(_07006_),
    .B(_07009_));
 sg13g2_buf_1 _16007_ (.A(_07010_),
    .X(_07011_));
 sg13g2_xnor2_1 _16008_ (.Y(_07012_),
    .A(_06974_),
    .B(_07011_));
 sg13g2_a21oi_1 _16009_ (.A1(net126),
    .A2(_07012_),
    .Y(_07013_),
    .B1(net318));
 sg13g2_buf_1 _16010_ (.A(net1163),
    .X(_07014_));
 sg13g2_xnor2_1 _16011_ (.Y(_07015_),
    .A(_06692_),
    .B(_07008_));
 sg13g2_xnor2_1 _16012_ (.Y(_07016_),
    .A(net947),
    .B(_07015_));
 sg13g2_nand2_1 _16013_ (.Y(_07017_),
    .A(_06653_),
    .B(_07016_));
 sg13g2_buf_1 _16014_ (.A(_00230_),
    .X(_07018_));
 sg13g2_nor2_1 _16015_ (.A(net1162),
    .B(_07011_),
    .Y(_07019_));
 sg13g2_and2_1 _16016_ (.A(_06653_),
    .B(_07016_),
    .X(_07020_));
 sg13g2_o21ai_1 _16017_ (.B1(_07011_),
    .Y(_07021_),
    .A1(net1162),
    .A2(_07020_));
 sg13g2_a21oi_1 _16018_ (.A1(net326),
    .A2(_07011_),
    .Y(_07022_),
    .B1(net1162));
 sg13g2_nor2_1 _16019_ (.A(_07017_),
    .B(_07022_),
    .Y(_07023_));
 sg13g2_a221oi_1 _16020_ (.B2(net157),
    .C1(_07023_),
    .B1(_07021_),
    .A1(_07017_),
    .Y(_07024_),
    .A2(_07019_));
 sg13g2_nand2_1 _16021_ (.Y(_07025_),
    .A(net1162),
    .B(_07011_));
 sg13g2_o21ai_1 _16022_ (.B1(_07025_),
    .Y(_07026_),
    .A1(net157),
    .A2(_07019_));
 sg13g2_nand2_1 _16023_ (.Y(_07027_),
    .A(_07017_),
    .B(_07026_));
 sg13g2_nor4_1 _16024_ (.A(net947),
    .B(net611),
    .C(net958),
    .D(net634),
    .Y(_07028_));
 sg13g2_nor2_1 _16025_ (.A(_06999_),
    .B(_06700_),
    .Y(_07029_));
 sg13g2_nand2_1 _16026_ (.Y(_07030_),
    .A(_07014_),
    .B(net950));
 sg13g2_o21ai_1 _16027_ (.B1(_07030_),
    .Y(_07031_),
    .A1(net634),
    .A2(net635));
 sg13g2_nor4_1 _16028_ (.A(_07000_),
    .B(_07028_),
    .C(_07029_),
    .D(_07031_),
    .Y(_07032_));
 sg13g2_buf_1 _16029_ (.A(net947),
    .X(_07033_));
 sg13g2_nor3_1 _16030_ (.A(net610),
    .B(net310),
    .C(net622),
    .Y(_07034_));
 sg13g2_a22oi_1 _16031_ (.Y(_07035_),
    .B1(_07034_),
    .B2(_06257_),
    .A2(_07032_),
    .A1(_06304_));
 sg13g2_mux2_1 _16032_ (.A0(_07024_),
    .A1(_07027_),
    .S(_07035_),
    .X(_07036_));
 sg13g2_or4_1 _16033_ (.A(_06953_),
    .B(_07005_),
    .C(_07013_),
    .D(_07036_),
    .X(_07037_));
 sg13g2_a21oi_1 _16034_ (.A1(_06633_),
    .A2(_06331_),
    .Y(_07038_),
    .B1(_06953_));
 sg13g2_a21o_1 _16035_ (.A2(_06953_),
    .A1(net48),
    .B1(_07038_),
    .X(_07039_));
 sg13g2_a21oi_1 _16036_ (.A1(_07037_),
    .A2(_07039_),
    .Y(_00320_),
    .B1(net350));
 sg13g2_buf_2 _16037_ (.A(\grid.cell_14_4.se ),
    .X(_07040_));
 sg13g2_buf_1 _16038_ (.A(net1161),
    .X(_07041_));
 sg13g2_nor4_1 _16039_ (.A(net946),
    .B(net947),
    .C(_06672_),
    .D(_06295_),
    .Y(_07042_));
 sg13g2_inv_1 _16040_ (.Y(_07043_),
    .A(net1161));
 sg13g2_buf_1 _16041_ (.A(_07043_),
    .X(_07044_));
 sg13g2_a21oi_1 _16042_ (.A1(_07044_),
    .A2(_06999_),
    .Y(_07045_),
    .B1(_06677_));
 sg13g2_nand2_1 _16043_ (.Y(_07046_),
    .A(_07041_),
    .B(net947));
 sg13g2_o21ai_1 _16044_ (.B1(_07046_),
    .Y(_07047_),
    .A1(_06295_),
    .A2(net966));
 sg13g2_nor3_1 _16045_ (.A(_07042_),
    .B(_07045_),
    .C(_07047_),
    .Y(_07048_));
 sg13g2_buf_1 _16046_ (.A(net946),
    .X(_07049_));
 sg13g2_nor3_1 _16047_ (.A(net608),
    .B(net610),
    .C(net316),
    .Y(_07050_));
 sg13g2_a22oi_1 _16048_ (.Y(_07051_),
    .B1(_07050_),
    .B2(_06298_),
    .A2(_07048_),
    .A1(net1168));
 sg13g2_buf_1 _16049_ (.A(_00046_),
    .X(_07052_));
 sg13g2_nand2_1 _16050_ (.Y(_07053_),
    .A(net1160),
    .B(_06187_));
 sg13g2_xnor2_1 _16051_ (.Y(_07054_),
    .A(net1161),
    .B(net1163));
 sg13g2_xnor2_1 _16052_ (.Y(_07055_),
    .A(_06686_),
    .B(_07054_));
 sg13g2_xnor2_1 _16053_ (.Y(_07056_),
    .A(_06253_),
    .B(_07055_));
 sg13g2_xnor2_1 _16054_ (.Y(_07057_),
    .A(net318),
    .B(_07056_));
 sg13g2_nand2b_1 _16055_ (.Y(_07058_),
    .B(net324),
    .A_N(net1160));
 sg13g2_o21ai_1 _16056_ (.B1(_07058_),
    .Y(_07059_),
    .A1(_06691_),
    .A2(_07056_));
 sg13g2_a21oi_1 _16057_ (.A1(_07053_),
    .A2(_07057_),
    .Y(_07060_),
    .B1(_07059_));
 sg13g2_xnor2_1 _16058_ (.Y(_07061_),
    .A(_07051_),
    .B(_07060_));
 sg13g2_nor2_1 _16059_ (.A(_06691_),
    .B(_07056_),
    .Y(_07062_));
 sg13g2_nor2b_1 _16060_ (.A(net1160),
    .B_N(_06593_),
    .Y(_07063_));
 sg13g2_nand2_1 _16061_ (.Y(_07064_),
    .A(net610),
    .B(net621));
 sg13g2_xnor2_1 _16062_ (.Y(_07065_),
    .A(net957),
    .B(net966));
 sg13g2_nor2_1 _16063_ (.A(_06999_),
    .B(_07065_),
    .Y(_07066_));
 sg13g2_nor3_1 _16064_ (.A(_07033_),
    .B(_06677_),
    .C(net634),
    .Y(_07067_));
 sg13g2_o21ai_1 _16065_ (.B1(net323),
    .Y(_07068_),
    .A1(_07066_),
    .A2(_07067_));
 sg13g2_o21ai_1 _16066_ (.B1(_07068_),
    .Y(_07069_),
    .A1(net1168),
    .A2(_07064_));
 sg13g2_nor3_1 _16067_ (.A(net608),
    .B(_06298_),
    .C(_07064_),
    .Y(_07070_));
 sg13g2_a221oi_1 _16068_ (.B2(_07049_),
    .C1(_07070_),
    .B1(_07069_),
    .A1(_07062_),
    .Y(_07071_),
    .A2(_07063_));
 sg13g2_a21oi_1 _16069_ (.A1(_07061_),
    .A2(_07071_),
    .Y(_07072_),
    .B1(net101));
 sg13g2_xnor2_1 _16070_ (.Y(_07073_),
    .A(_06975_),
    .B(_07056_));
 sg13g2_a21oi_1 _16071_ (.A1(net77),
    .A2(_07073_),
    .Y(_07074_),
    .B1(net622));
 sg13g2_or3_1 _16072_ (.A(_06855_),
    .B(_07072_),
    .C(_07074_),
    .X(_07075_));
 sg13g2_o21ai_1 _16073_ (.B1(_07075_),
    .Y(_00321_),
    .A1(_04942_),
    .A2(_06954_));
 sg13g2_buf_1 _16074_ (.A(\grid.cell_14_5.se ),
    .X(_07076_));
 sg13g2_xnor2_1 _16075_ (.Y(_07077_),
    .A(net1159),
    .B(_06713_));
 sg13g2_buf_2 _16076_ (.A(_07077_),
    .X(_07078_));
 sg13g2_xnor2_1 _16077_ (.Y(_07079_),
    .A(_06351_),
    .B(_07078_));
 sg13g2_xnor2_1 _16078_ (.Y(_07080_),
    .A(_07040_),
    .B(_07079_));
 sg13g2_and2_1 _16079_ (.A(_06743_),
    .B(_07080_),
    .X(_07081_));
 sg13g2_buf_2 _16080_ (.A(_00078_),
    .X(_07082_));
 sg13g2_xor2_1 _16081_ (.B(net633),
    .A(net622),
    .X(_07083_));
 sg13g2_nor2_1 _16082_ (.A(_07082_),
    .B(_07083_),
    .Y(_07084_));
 sg13g2_nand2_1 _16083_ (.Y(_07085_),
    .A(net946),
    .B(net956));
 sg13g2_xnor2_1 _16084_ (.Y(_07086_),
    .A(net956),
    .B(net632));
 sg13g2_nor2_1 _16085_ (.A(net609),
    .B(_07086_),
    .Y(_07087_));
 sg13g2_nor3_1 _16086_ (.A(net946),
    .B(_06732_),
    .C(_06295_),
    .Y(_07088_));
 sg13g2_o21ai_1 _16087_ (.B1(net322),
    .Y(_07089_),
    .A1(_07087_),
    .A2(_07088_));
 sg13g2_o21ai_1 _16088_ (.B1(_07089_),
    .Y(_07090_),
    .A1(_06392_),
    .A2(_07085_));
 sg13g2_buf_1 _16089_ (.A(net1159),
    .X(_07091_));
 sg13g2_buf_1 _16090_ (.A(net945),
    .X(_07092_));
 sg13g2_nand2_1 _16091_ (.Y(_07093_),
    .A(net322),
    .B(net323));
 sg13g2_nor3_1 _16092_ (.A(net607),
    .B(_07093_),
    .C(_07085_),
    .Y(_07094_));
 sg13g2_a221oi_1 _16093_ (.B2(net607),
    .C1(_07094_),
    .B1(_07090_),
    .A1(_07081_),
    .Y(_07095_),
    .A2(_07084_));
 sg13g2_nor2_1 _16094_ (.A(net631),
    .B(net632),
    .Y(_07096_));
 sg13g2_buf_1 _16095_ (.A(net1159),
    .X(_07097_));
 sg13g2_nor4_1 _16096_ (.A(net944),
    .B(_07041_),
    .C(_06728_),
    .D(net631),
    .Y(_07098_));
 sg13g2_nand2_1 _16097_ (.Y(_07099_),
    .A(net944),
    .B(net956));
 sg13g2_nand2_1 _16098_ (.Y(_07100_),
    .A(_07085_),
    .B(_07099_));
 sg13g2_inv_1 _16099_ (.Y(_07101_),
    .A(net1159));
 sg13g2_buf_1 _16100_ (.A(_07101_),
    .X(_07102_));
 sg13g2_nor2_1 _16101_ (.A(net606),
    .B(net609),
    .Y(_07103_));
 sg13g2_nor4_1 _16102_ (.A(_07096_),
    .B(_07098_),
    .C(_07100_),
    .D(_07103_),
    .Y(_07104_));
 sg13g2_nor3_1 _16103_ (.A(_07091_),
    .B(_07049_),
    .C(net315),
    .Y(_07105_));
 sg13g2_a22oi_1 _16104_ (.Y(_07106_),
    .B1(_07105_),
    .B2(_07093_),
    .A2(_07104_),
    .A1(_06392_));
 sg13g2_nand2_1 _16105_ (.Y(_07107_),
    .A(_07082_),
    .B(net634));
 sg13g2_xnor2_1 _16106_ (.Y(_07108_),
    .A(net620),
    .B(_07080_));
 sg13g2_nor2_1 _16107_ (.A(_07082_),
    .B(net634),
    .Y(_07109_));
 sg13g2_a221oi_1 _16108_ (.B2(_07108_),
    .C1(_07109_),
    .B1(_07107_),
    .A1(_06743_),
    .Y(_07110_),
    .A2(_07080_));
 sg13g2_xnor2_1 _16109_ (.Y(_07111_),
    .A(_07106_),
    .B(_07110_));
 sg13g2_a21oi_1 _16110_ (.A1(_07095_),
    .A2(_07111_),
    .Y(_07112_),
    .B1(net101));
 sg13g2_xnor2_1 _16111_ (.Y(_07113_),
    .A(net634),
    .B(_07006_));
 sg13g2_xnor2_1 _16112_ (.Y(_07114_),
    .A(_07080_),
    .B(_07113_));
 sg13g2_a21oi_1 _16113_ (.A1(net77),
    .A2(_07114_),
    .Y(_07115_),
    .B1(net316));
 sg13g2_or3_1 _16114_ (.A(_06855_),
    .B(_07112_),
    .C(_07115_),
    .X(_07116_));
 sg13g2_o21ai_1 _16115_ (.B1(_07116_),
    .Y(_00322_),
    .A1(net46),
    .A2(_06954_));
 sg13g2_buf_1 _16116_ (.A(net117),
    .X(_07117_));
 sg13g2_nand2_1 _16117_ (.Y(_07118_),
    .A(_06729_),
    .B(net73));
 sg13g2_buf_2 _16118_ (.A(_00140_),
    .X(_07119_));
 sg13g2_o21ai_1 _16119_ (.B1(_06417_),
    .Y(_07120_),
    .A1(_07119_),
    .A2(_06879_));
 sg13g2_inv_1 _16120_ (.Y(_07121_),
    .A(_07119_));
 sg13g2_nand2_1 _16121_ (.Y(_07122_),
    .A(_07121_),
    .B(net155));
 sg13g2_o21ai_1 _16122_ (.B1(_07122_),
    .Y(_07123_),
    .A1(net155),
    .A2(_07120_));
 sg13g2_o21ai_1 _16123_ (.B1(_06879_),
    .Y(_07124_),
    .A1(net945),
    .A2(net155));
 sg13g2_nor2_1 _16124_ (.A(net944),
    .B(_06879_),
    .Y(_07125_));
 sg13g2_a21oi_1 _16125_ (.A1(_07119_),
    .A2(_07124_),
    .Y(_07126_),
    .B1(_07125_));
 sg13g2_nor2_1 _16126_ (.A(_07121_),
    .B(net944),
    .Y(_07127_));
 sg13g2_nand2_1 _16127_ (.Y(_07128_),
    .A(net614),
    .B(net639));
 sg13g2_nand2_1 _16128_ (.Y(_07129_),
    .A(_06871_),
    .B(_07128_));
 sg13g2_nor2b_1 _16129_ (.A(_07119_),
    .B_N(net615),
    .Y(_07130_));
 sg13g2_a22oi_1 _16130_ (.Y(_07131_),
    .B1(_07130_),
    .B2(_06491_),
    .A2(_07129_),
    .A1(_07127_));
 sg13g2_and2_1 _16131_ (.A(_07097_),
    .B(_06859_),
    .X(_07132_));
 sg13g2_a21oi_1 _16132_ (.A1(_06491_),
    .A2(_07132_),
    .Y(_07133_),
    .B1(_07125_));
 sg13g2_mux2_1 _16133_ (.A0(_07131_),
    .A1(_07133_),
    .S(net631),
    .X(_07134_));
 sg13g2_o21ai_1 _16134_ (.B1(_07134_),
    .Y(_07135_),
    .A1(net321),
    .A2(_07126_));
 sg13g2_a21oi_1 _16135_ (.A1(net607),
    .A2(_07123_),
    .Y(_07136_),
    .B1(_07135_));
 sg13g2_buf_1 _16136_ (.A(_00110_),
    .X(_07137_));
 sg13g2_inv_1 _16137_ (.Y(_07138_),
    .A(_07137_));
 sg13g2_xnor2_1 _16138_ (.Y(_07139_),
    .A(_06394_),
    .B(_06845_));
 sg13g2_xnor2_1 _16139_ (.Y(_07140_),
    .A(_07097_),
    .B(_07139_));
 sg13g2_xnor2_1 _16140_ (.Y(_07141_),
    .A(_06677_),
    .B(_07140_));
 sg13g2_o21ai_1 _16141_ (.B1(_07141_),
    .Y(_07142_),
    .A1(_07138_),
    .A2(net323));
 sg13g2_nand2_1 _16142_ (.Y(_07143_),
    .A(_06785_),
    .B(_07140_));
 sg13g2_nand2_1 _16143_ (.Y(_07144_),
    .A(_07138_),
    .B(net323));
 sg13g2_nand3_1 _16144_ (.B(_07143_),
    .C(_07144_),
    .A(_07142_),
    .Y(_07145_));
 sg13g2_xor2_1 _16145_ (.B(_07145_),
    .A(_07136_),
    .X(_07146_));
 sg13g2_buf_1 _16146_ (.A(_06888_),
    .X(_07147_));
 sg13g2_xor2_1 _16147_ (.B(net630),
    .A(_06796_),
    .X(_07148_));
 sg13g2_nand2_1 _16148_ (.Y(_07149_),
    .A(net313),
    .B(_07148_));
 sg13g2_o21ai_1 _16149_ (.B1(_07149_),
    .Y(_07150_),
    .A1(_07147_),
    .A2(_06823_));
 sg13g2_a22oi_1 _16150_ (.Y(_07151_),
    .B1(_07150_),
    .B2(net321),
    .A2(_06844_),
    .A1(_07121_));
 sg13g2_a21oi_1 _16151_ (.A1(_06417_),
    .A2(_06844_),
    .Y(_07152_),
    .B1(net607));
 sg13g2_a21oi_1 _16152_ (.A1(_07092_),
    .A2(_07151_),
    .Y(_07153_),
    .B1(_07152_));
 sg13g2_inv_1 _16153_ (.Y(_07154_),
    .A(_06686_));
 sg13g2_nor3_1 _16154_ (.A(_07137_),
    .B(_07154_),
    .C(_07143_),
    .Y(_07155_));
 sg13g2_xnor2_1 _16155_ (.Y(_07156_),
    .A(_07040_),
    .B(_06670_));
 sg13g2_xnor2_1 _16156_ (.Y(_07157_),
    .A(_06295_),
    .B(_07156_));
 sg13g2_xnor2_1 _16157_ (.Y(_07158_),
    .A(_07140_),
    .B(_07157_));
 sg13g2_nor2_1 _16158_ (.A(net315),
    .B(_07158_),
    .Y(_07159_));
 sg13g2_nor4_1 _16159_ (.A(net125),
    .B(_07153_),
    .C(_07155_),
    .D(_07159_),
    .Y(_07160_));
 sg13g2_a22oi_1 _16160_ (.Y(_07161_),
    .B1(_07146_),
    .B2(_07160_),
    .A2(_06853_),
    .A1(_06810_));
 sg13g2_a221oi_1 _16161_ (.B2(_07161_),
    .C1(net617),
    .B1(_07118_),
    .A1(net24),
    .Y(_00323_),
    .A2(_06853_));
 sg13g2_nand2_1 _16162_ (.Y(_07162_),
    .A(_05678_),
    .B(_06953_));
 sg13g2_nand2_1 _16163_ (.Y(_07163_),
    .A(_06859_),
    .B(net619));
 sg13g2_nor2_1 _16164_ (.A(_06870_),
    .B(net956),
    .Y(_07164_));
 sg13g2_nand2_1 _16165_ (.Y(_07165_),
    .A(_07121_),
    .B(_07164_));
 sg13g2_nand3_1 _16166_ (.B(_07163_),
    .C(_07165_),
    .A(_06417_),
    .Y(_07166_));
 sg13g2_o21ai_1 _16167_ (.B1(_07166_),
    .Y(_07167_),
    .A1(_07119_),
    .A2(_07163_));
 sg13g2_o21ai_1 _16168_ (.B1(_07128_),
    .Y(_07168_),
    .A1(net313),
    .A2(net618));
 sg13g2_nand2_1 _16169_ (.Y(_07169_),
    .A(_07127_),
    .B(_07168_));
 sg13g2_nand3_1 _16170_ (.B(net321),
    .C(_07130_),
    .A(net619),
    .Y(_07170_));
 sg13g2_nand3_1 _16171_ (.B(_07169_),
    .C(_07170_),
    .A(net322),
    .Y(_07171_));
 sg13g2_nand2_1 _16172_ (.Y(_07172_),
    .A(net606),
    .B(_07164_));
 sg13g2_nand3_1 _16173_ (.B(net321),
    .C(_07132_),
    .A(net619),
    .Y(_07173_));
 sg13g2_nand3_1 _16174_ (.B(_07172_),
    .C(_07173_),
    .A(net631),
    .Y(_07174_));
 sg13g2_and2_1 _16175_ (.A(_06870_),
    .B(_06713_),
    .X(_07175_));
 sg13g2_buf_1 _16176_ (.A(_07175_),
    .X(_07176_));
 sg13g2_nor2_1 _16177_ (.A(net945),
    .B(_07176_),
    .Y(_07177_));
 sg13g2_o21ai_1 _16178_ (.B1(_07119_),
    .Y(_07178_),
    .A1(_07164_),
    .A2(_07177_));
 sg13g2_a21oi_1 _16179_ (.A1(_07172_),
    .A2(_07178_),
    .Y(_07179_),
    .B1(net321));
 sg13g2_a221oi_1 _16180_ (.B2(_07174_),
    .C1(_07179_),
    .B1(_07171_),
    .A1(_07092_),
    .Y(_07180_),
    .A2(_07167_));
 sg13g2_xnor2_1 _16181_ (.Y(_07181_),
    .A(_06394_),
    .B(_07078_));
 sg13g2_xnor2_1 _16182_ (.Y(_07182_),
    .A(net955),
    .B(_07181_));
 sg13g2_xnor2_1 _16183_ (.Y(_07183_),
    .A(_06917_),
    .B(_07182_));
 sg13g2_nor2_1 _16184_ (.A(_06894_),
    .B(_07183_),
    .Y(_07184_));
 sg13g2_xor2_1 _16185_ (.B(_07182_),
    .A(net1167),
    .X(_07185_));
 sg13g2_a22oi_1 _16186_ (.Y(_07186_),
    .B1(_07185_),
    .B2(net971),
    .A2(_07182_),
    .A1(_06512_));
 sg13g2_nor2b_1 _16187_ (.A(_07184_),
    .B_N(_07186_),
    .Y(_07187_));
 sg13g2_xnor2_1 _16188_ (.Y(_07188_),
    .A(_07186_),
    .B(_07184_));
 sg13g2_nand2_1 _16189_ (.Y(_07189_),
    .A(net1159),
    .B(net955));
 sg13g2_nor2b_1 _16190_ (.A(_07091_),
    .B_N(net629),
    .Y(_07190_));
 sg13g2_a221oi_1 _16191_ (.B2(_07190_),
    .C1(_07176_),
    .B1(_07164_),
    .A1(net631),
    .Y(_07191_),
    .A2(net629));
 sg13g2_nand4_1 _16192_ (.B(_07099_),
    .C(_07189_),
    .A(_07119_),
    .Y(_07192_),
    .D(_07191_));
 sg13g2_o21ai_1 _16193_ (.B1(_07192_),
    .Y(_07193_),
    .A1(_06417_),
    .A2(_07172_));
 sg13g2_buf_1 _16194_ (.A(net163),
    .X(_07194_));
 sg13g2_a221oi_1 _16195_ (.B2(_07193_),
    .C1(net100),
    .B1(_07188_),
    .A1(_07180_),
    .Y(_07195_),
    .A2(_07187_));
 sg13g2_xor2_1 _16196_ (.B(_07182_),
    .A(_06946_),
    .X(_07196_));
 sg13g2_a21oi_1 _16197_ (.A1(net109),
    .A2(_07196_),
    .Y(_07197_),
    .B1(_06797_));
 sg13g2_or3_1 _16198_ (.A(_06953_),
    .B(_07195_),
    .C(_07197_),
    .X(_07198_));
 sg13g2_a21oi_1 _16199_ (.A1(_07162_),
    .A2(_07198_),
    .Y(_00324_),
    .B1(net350));
 sg13g2_buf_1 _16200_ (.A(net120),
    .X(_07199_));
 sg13g2_nor3_1 _16201_ (.A(net375),
    .B(_05750_),
    .C(net159),
    .Y(_07200_));
 sg13g2_buf_1 _16202_ (.A(_07200_),
    .X(_07201_));
 sg13g2_a22oi_1 _16203_ (.Y(_07202_),
    .B1(net59),
    .B2(_01806_),
    .A2(net72),
    .A1(net953));
 sg13g2_buf_2 _16204_ (.A(\grid.cell_15_0.se ),
    .X(_07203_));
 sg13g2_buf_1 _16205_ (.A(_07203_),
    .X(_07204_));
 sg13g2_buf_1 _16206_ (.A(_07204_),
    .X(_07205_));
 sg13g2_nand2_1 _16207_ (.Y(_07206_),
    .A(net624),
    .B(net156));
 sg13g2_buf_2 _16208_ (.A(\grid.cell_15_0.sw ),
    .X(_07207_));
 sg13g2_buf_1 _16209_ (.A(_07207_),
    .X(_07208_));
 sg13g2_buf_1 _16210_ (.A(net942),
    .X(_07209_));
 sg13g2_buf_1 _16211_ (.A(net604),
    .X(_07210_));
 sg13g2_buf_1 _16212_ (.A(_07210_),
    .X(_07211_));
 sg13g2_nor2_1 _16213_ (.A(net153),
    .B(net154),
    .Y(_07212_));
 sg13g2_and2_1 _16214_ (.A(net942),
    .B(net614),
    .X(_07213_));
 sg13g2_buf_1 _16215_ (.A(_07213_),
    .X(_07214_));
 sg13g2_xnor2_1 _16216_ (.Y(_07215_),
    .A(_07207_),
    .B(_06840_));
 sg13g2_buf_2 _16217_ (.A(_07215_),
    .X(_07216_));
 sg13g2_nand2b_1 _16218_ (.Y(_07217_),
    .B(net963),
    .A_N(_07216_));
 sg13g2_o21ai_1 _16219_ (.B1(_07217_),
    .Y(_07218_),
    .A1(net156),
    .A2(_07214_));
 sg13g2_a22oi_1 _16220_ (.Y(_07219_),
    .B1(_07218_),
    .B2(net948),
    .A2(_07212_),
    .A1(_07206_));
 sg13g2_nand2_1 _16221_ (.Y(_07220_),
    .A(net963),
    .B(net943));
 sg13g2_nand2_1 _16222_ (.Y(_07221_),
    .A(net156),
    .B(_07220_));
 sg13g2_nand3_1 _16223_ (.B(_07221_),
    .C(_07212_),
    .A(net948),
    .Y(_07222_));
 sg13g2_o21ai_1 _16224_ (.B1(_07222_),
    .Y(_07223_),
    .A1(net605),
    .A2(_07219_));
 sg13g2_xnor2_1 _16225_ (.Y(_07224_),
    .A(_06478_),
    .B(_07203_));
 sg13g2_xor2_1 _16226_ (.B(_07224_),
    .A(_07216_),
    .X(_07225_));
 sg13g2_xnor2_1 _16227_ (.Y(_07226_),
    .A(net314),
    .B(_07225_));
 sg13g2_nor2_1 _16228_ (.A(_06972_),
    .B(_07226_),
    .Y(_07227_));
 sg13g2_xnor2_1 _16229_ (.Y(_07228_),
    .A(net1165),
    .B(_07224_));
 sg13g2_inv_1 _16230_ (.Y(_07229_),
    .A(_07207_));
 sg13g2_xnor2_1 _16231_ (.Y(_07230_),
    .A(_07229_),
    .B(_06845_));
 sg13g2_xnor2_1 _16232_ (.Y(_07231_),
    .A(_07228_),
    .B(_07230_));
 sg13g2_buf_2 _16233_ (.A(_07231_),
    .X(_07232_));
 sg13g2_buf_1 _16234_ (.A(_00229_),
    .X(_07233_));
 sg13g2_inv_1 _16235_ (.Y(_07234_),
    .A(net1158));
 sg13g2_o21ai_1 _16236_ (.B1(_07234_),
    .Y(_07235_),
    .A1(net961),
    .A2(_07232_));
 sg13g2_nor2_1 _16237_ (.A(net1158),
    .B(_07227_),
    .Y(_07236_));
 sg13g2_a22oi_1 _16238_ (.Y(_07237_),
    .B1(_07236_),
    .B2(_07232_),
    .A2(_07235_),
    .A1(_07227_));
 sg13g2_o21ai_1 _16239_ (.B1(net961),
    .Y(_07238_),
    .A1(_07232_),
    .A2(_07236_));
 sg13g2_nand2_1 _16240_ (.Y(_07239_),
    .A(_07237_),
    .B(_07238_));
 sg13g2_or2_1 _16241_ (.X(_07240_),
    .B(net955),
    .A(_07207_));
 sg13g2_buf_1 _16242_ (.A(_07240_),
    .X(_07241_));
 sg13g2_nor2_1 _16243_ (.A(net948),
    .B(_07241_),
    .Y(_07242_));
 sg13g2_nand2b_1 _16244_ (.Y(_07243_),
    .B(net604),
    .A_N(net615));
 sg13g2_buf_1 _16245_ (.A(_07229_),
    .X(_07244_));
 sg13g2_nand2_1 _16246_ (.Y(_07245_),
    .A(net603),
    .B(net314));
 sg13g2_a21oi_1 _16247_ (.A1(_07243_),
    .A2(_07245_),
    .Y(_07246_),
    .B1(net963));
 sg13g2_nand2b_1 _16248_ (.Y(_07247_),
    .B(net614),
    .A_N(_07208_));
 sg13g2_nand2_1 _16249_ (.Y(_07248_),
    .A(net615),
    .B(_06606_));
 sg13g2_nand2_1 _16250_ (.Y(_07249_),
    .A(net309),
    .B(_07248_));
 sg13g2_a21oi_1 _16251_ (.A1(_07247_),
    .A2(_07249_),
    .Y(_07250_),
    .B1(net156));
 sg13g2_or3_1 _16252_ (.A(_07242_),
    .B(_07246_),
    .C(_07250_),
    .X(_07251_));
 sg13g2_o21ai_1 _16253_ (.B1(_06875_),
    .Y(_07252_),
    .A1(_06888_),
    .A2(net948));
 sg13g2_nand3_1 _16254_ (.B(net314),
    .C(_07241_),
    .A(net628),
    .Y(_07253_));
 sg13g2_o21ai_1 _16255_ (.B1(_07253_),
    .Y(_07254_),
    .A1(net309),
    .A2(_07248_));
 sg13g2_a21oi_1 _16256_ (.A1(_07211_),
    .A2(_07252_),
    .Y(_07255_),
    .B1(_07254_));
 sg13g2_nor3_1 _16257_ (.A(net943),
    .B(net309),
    .C(_06871_),
    .Y(_07256_));
 sg13g2_inv_1 _16258_ (.Y(_07257_),
    .A(_07203_));
 sg13g2_nand2_1 _16259_ (.Y(_07258_),
    .A(net604),
    .B(net313));
 sg13g2_nor3_1 _16260_ (.A(_07257_),
    .B(_06606_),
    .C(_07258_),
    .Y(_07259_));
 sg13g2_o21ai_1 _16261_ (.B1(net624),
    .Y(_07260_),
    .A1(_07256_),
    .A2(_07259_));
 sg13g2_o21ai_1 _16262_ (.B1(_07260_),
    .Y(_07261_),
    .A1(net605),
    .A2(_07255_));
 sg13g2_a21oi_1 _16263_ (.A1(net605),
    .A2(_07251_),
    .Y(_07262_),
    .B1(_07261_));
 sg13g2_inv_1 _16264_ (.Y(_07263_),
    .A(_07232_));
 sg13g2_a21oi_1 _16265_ (.A1(_07234_),
    .A2(_07232_),
    .Y(_07264_),
    .B1(net961));
 sg13g2_a21oi_1 _16266_ (.A1(net1158),
    .A2(_07263_),
    .Y(_07265_),
    .B1(_07264_));
 sg13g2_nor3_1 _16267_ (.A(_07227_),
    .B(_07262_),
    .C(_07265_),
    .Y(_07266_));
 sg13g2_a21oi_1 _16268_ (.A1(_07223_),
    .A2(_07239_),
    .Y(_07267_),
    .B1(_07266_));
 sg13g2_buf_2 _16269_ (.A(\grid.cell_15_0.s ),
    .X(_07268_));
 sg13g2_buf_1 _16270_ (.A(_07268_),
    .X(_07269_));
 sg13g2_xnor2_1 _16271_ (.Y(_07270_),
    .A(net961),
    .B(_07269_));
 sg13g2_xnor2_1 _16272_ (.Y(_07271_),
    .A(_07232_),
    .B(_07270_));
 sg13g2_a21oi_1 _16273_ (.A1(net78),
    .A2(_07271_),
    .Y(_07272_),
    .B1(net953));
 sg13g2_nor2_2 _16274_ (.A(_05750_),
    .B(_06063_),
    .Y(_07273_));
 sg13g2_nand2_2 _16275_ (.Y(_07274_),
    .A(_06114_),
    .B(_07273_));
 sg13g2_o21ai_1 _16276_ (.B1(net668),
    .Y(_07275_),
    .A1(_01806_),
    .A2(_07274_));
 sg13g2_a221oi_1 _16277_ (.B2(_07274_),
    .C1(_07275_),
    .B1(_07272_),
    .A1(_07202_),
    .Y(_00325_),
    .A2(_07267_));
 sg13g2_buf_1 _16278_ (.A(_03153_),
    .X(_07276_));
 sg13g2_nand2_1 _16279_ (.Y(_07277_),
    .A(net42),
    .B(net59));
 sg13g2_nand2_1 _16280_ (.Y(_07278_),
    .A(_06856_),
    .B(_06921_));
 sg13g2_buf_1 _16281_ (.A(\grid.cell_15_1.se ),
    .X(_07279_));
 sg13g2_xnor2_1 _16282_ (.Y(_07280_),
    .A(net1157),
    .B(_06907_));
 sg13g2_xor2_1 _16283_ (.B(_07280_),
    .A(_07224_),
    .X(_07281_));
 sg13g2_buf_1 _16284_ (.A(_07281_),
    .X(_07282_));
 sg13g2_nor2_1 _16285_ (.A(net1167),
    .B(_06894_),
    .Y(_07283_));
 sg13g2_or2_1 _16286_ (.X(_07284_),
    .B(_07283_),
    .A(_07282_));
 sg13g2_nor3_1 _16287_ (.A(_06856_),
    .B(_06921_),
    .C(_07282_),
    .Y(_07285_));
 sg13g2_a221oi_1 _16288_ (.B2(_06857_),
    .C1(_07285_),
    .B1(_07284_),
    .A1(net961),
    .Y(_07286_),
    .A2(_07278_));
 sg13g2_xnor2_1 _16289_ (.Y(_07287_),
    .A(_06856_),
    .B(_07282_));
 sg13g2_nor2_1 _16290_ (.A(_06894_),
    .B(_07282_),
    .Y(_07288_));
 sg13g2_a22oi_1 _16291_ (.Y(_07289_),
    .B1(_07288_),
    .B2(net1158),
    .A2(_07287_),
    .A1(net961));
 sg13g2_o21ai_1 _16292_ (.B1(_07289_),
    .Y(_07290_),
    .A1(net1158),
    .A2(_07286_));
 sg13g2_buf_1 _16293_ (.A(net1157),
    .X(_07291_));
 sg13g2_nor3_1 _16294_ (.A(net319),
    .B(net613),
    .C(net940),
    .Y(_07292_));
 sg13g2_a22oi_1 _16295_ (.Y(_07293_),
    .B1(_06904_),
    .B2(net940),
    .A2(net625),
    .A1(net628));
 sg13g2_nor2b_1 _16296_ (.A(_07292_),
    .B_N(_07293_),
    .Y(_07294_));
 sg13g2_nand2_1 _16297_ (.Y(_07295_),
    .A(_06478_),
    .B(_06539_));
 sg13g2_nor2_2 _16298_ (.A(_06903_),
    .B(net940),
    .Y(_07296_));
 sg13g2_a22oi_1 _16299_ (.Y(_07297_),
    .B1(_07295_),
    .B2(_07296_),
    .A2(_07294_),
    .A1(net948));
 sg13g2_nand2_1 _16300_ (.Y(_07298_),
    .A(net626),
    .B(_07220_));
 sg13g2_nand3_1 _16301_ (.B(_07296_),
    .C(_07298_),
    .A(net948),
    .Y(_07299_));
 sg13g2_o21ai_1 _16302_ (.B1(_07299_),
    .Y(_07300_),
    .A1(net605),
    .A2(_07297_));
 sg13g2_buf_1 _16303_ (.A(_07257_),
    .X(_07301_));
 sg13g2_inv_1 _16304_ (.Y(_07302_),
    .A(net1157));
 sg13g2_nor2_1 _16305_ (.A(_07302_),
    .B(_06605_),
    .Y(_07303_));
 sg13g2_nand2_1 _16306_ (.Y(_07304_),
    .A(_07302_),
    .B(_06605_));
 sg13g2_o21ai_1 _16307_ (.B1(_07304_),
    .Y(_07305_),
    .A1(net952),
    .A2(_07303_));
 sg13g2_nand2_1 _16308_ (.Y(_07306_),
    .A(_07291_),
    .B(_06978_));
 sg13g2_or2_1 _16309_ (.X(_07307_),
    .B(_06605_),
    .A(net1157));
 sg13g2_nand2_1 _16310_ (.Y(_07308_),
    .A(net952),
    .B(_07307_));
 sg13g2_a21oi_1 _16311_ (.A1(_07306_),
    .A2(_07308_),
    .Y(_07309_),
    .B1(_07295_));
 sg13g2_a21oi_1 _16312_ (.A1(net319),
    .A2(_07305_),
    .Y(_07310_),
    .B1(_07309_));
 sg13g2_nor2_1 _16313_ (.A(net1157),
    .B(_07295_),
    .Y(_07311_));
 sg13g2_or2_1 _16314_ (.X(_07312_),
    .B(_07311_),
    .A(_07303_));
 sg13g2_nor2_1 _16315_ (.A(net613),
    .B(_07295_),
    .Y(_07313_));
 sg13g2_a221oi_1 _16316_ (.B2(_07307_),
    .C1(_07301_),
    .B1(_07313_),
    .A1(net613),
    .Y(_07314_),
    .A2(_07312_));
 sg13g2_a21oi_1 _16317_ (.A1(net602),
    .A2(_07310_),
    .Y(_07315_),
    .B1(_07314_));
 sg13g2_nor2b_1 _16318_ (.A(net1158),
    .B_N(net1167),
    .Y(_07316_));
 sg13g2_nand3_1 _16319_ (.B(_06978_),
    .C(_07296_),
    .A(net319),
    .Y(_07317_));
 sg13g2_nand2b_1 _16320_ (.Y(_07318_),
    .B(_07317_),
    .A_N(_07316_));
 sg13g2_nand2_1 _16321_ (.Y(_07319_),
    .A(_07301_),
    .B(_07296_));
 sg13g2_nand2_1 _16322_ (.Y(_07320_),
    .A(_07203_),
    .B(_07291_));
 sg13g2_or2_1 _16323_ (.X(_07321_),
    .B(_07320_),
    .A(_06908_));
 sg13g2_a21oi_1 _16324_ (.A1(_07319_),
    .A2(_07321_),
    .Y(_07322_),
    .B1(net624));
 sg13g2_nor4_1 _16325_ (.A(_07288_),
    .B(_07315_),
    .C(_07318_),
    .D(_07322_),
    .Y(_07323_));
 sg13g2_nand2b_1 _16326_ (.Y(_07324_),
    .B(_07233_),
    .A_N(net961));
 sg13g2_nand2_1 _16327_ (.Y(_07325_),
    .A(_07287_),
    .B(_07324_));
 sg13g2_a221oi_1 _16328_ (.B2(_07325_),
    .C1(net100),
    .B1(_07323_),
    .A1(_07290_),
    .Y(_07326_),
    .A2(_07300_));
 sg13g2_xor2_1 _16329_ (.B(_07268_),
    .A(_06856_),
    .X(_07327_));
 sg13g2_xor2_1 _16330_ (.B(_07327_),
    .A(net1167),
    .X(_07328_));
 sg13g2_xnor2_1 _16331_ (.Y(_07329_),
    .A(_07282_),
    .B(_07328_));
 sg13g2_a21oi_1 _16332_ (.A1(net109),
    .A2(_07329_),
    .Y(_07330_),
    .B1(net612));
 sg13g2_or3_1 _16333_ (.A(net59),
    .B(_07326_),
    .C(_07330_),
    .X(_07331_));
 sg13g2_a21oi_1 _16334_ (.A1(_07277_),
    .A2(_07331_),
    .Y(_00326_),
    .B1(net350));
 sg13g2_buf_1 _16335_ (.A(\grid.cell_15_2.se ),
    .X(_07332_));
 sg13g2_buf_1 _16336_ (.A(net1156),
    .X(_07333_));
 sg13g2_buf_1 _16337_ (.A(net939),
    .X(_07334_));
 sg13g2_buf_1 _16338_ (.A(net940),
    .X(_07335_));
 sg13g2_buf_1 _16339_ (.A(net600),
    .X(_07336_));
 sg13g2_a21oi_1 _16340_ (.A1(net626),
    .A2(net308),
    .Y(_07337_),
    .B1(_06958_));
 sg13g2_nor4_1 _16341_ (.A(net601),
    .B(net310),
    .C(_06653_),
    .D(_07337_),
    .Y(_07338_));
 sg13g2_xnor2_1 _16342_ (.Y(_07339_),
    .A(net1156),
    .B(_06955_));
 sg13g2_nor2_1 _16343_ (.A(net319),
    .B(_07339_),
    .Y(_07340_));
 sg13g2_a21oi_1 _16344_ (.A1(net601),
    .A2(net310),
    .Y(_07341_),
    .B1(net318));
 sg13g2_o21ai_1 _16345_ (.B1(_06636_),
    .Y(_07342_),
    .A1(_07340_),
    .A2(_07341_));
 sg13g2_nor2_1 _16346_ (.A(net939),
    .B(_06956_),
    .Y(_07343_));
 sg13g2_o21ai_1 _16347_ (.B1(_07343_),
    .Y(_07344_),
    .A1(net319),
    .A2(_06958_));
 sg13g2_a21oi_1 _16348_ (.A1(_07342_),
    .A2(_07344_),
    .Y(_07345_),
    .B1(net308));
 sg13g2_buf_1 _16349_ (.A(_00228_),
    .X(_07346_));
 sg13g2_buf_1 _16350_ (.A(_07346_),
    .X(_07347_));
 sg13g2_xnor2_1 _16351_ (.Y(_07348_),
    .A(net959),
    .B(_07339_));
 sg13g2_xnor2_1 _16352_ (.Y(_07349_),
    .A(net960),
    .B(_07279_));
 sg13g2_xnor2_1 _16353_ (.Y(_07350_),
    .A(_07348_),
    .B(_07349_));
 sg13g2_buf_1 _16354_ (.A(_07350_),
    .X(_07351_));
 sg13g2_o21ai_1 _16355_ (.B1(_07351_),
    .Y(_07352_),
    .A1(net624),
    .A2(_06972_));
 sg13g2_nor2_1 _16356_ (.A(_06912_),
    .B(_06979_),
    .Y(_07353_));
 sg13g2_a21oi_1 _16357_ (.A1(net612),
    .A2(_06979_),
    .Y(_07354_),
    .B1(net628));
 sg13g2_a221oi_1 _16358_ (.B2(_07351_),
    .C1(_07354_),
    .B1(_07353_),
    .A1(_06912_),
    .Y(_07355_),
    .A2(_07352_));
 sg13g2_xnor2_1 _16359_ (.Y(_07356_),
    .A(net616),
    .B(_07351_));
 sg13g2_and2_1 _16360_ (.A(_06979_),
    .B(_07351_),
    .X(_07357_));
 sg13g2_a22oi_1 _16361_ (.Y(_07358_),
    .B1(_07357_),
    .B2(_07347_),
    .A2(_07356_),
    .A1(net624));
 sg13g2_o21ai_1 _16362_ (.B1(_07358_),
    .Y(_07359_),
    .A1(_07347_),
    .A2(_07355_));
 sg13g2_o21ai_1 _16363_ (.B1(_07359_),
    .Y(_07360_),
    .A1(_07338_),
    .A2(_07345_));
 sg13g2_inv_1 _16364_ (.Y(_07361_),
    .A(_07346_));
 sg13g2_buf_1 _16365_ (.A(_07361_),
    .X(_07362_));
 sg13g2_nand2_1 _16366_ (.Y(_07363_),
    .A(_06965_),
    .B(_06653_));
 sg13g2_buf_1 _16367_ (.A(net939),
    .X(_07364_));
 sg13g2_nor2_1 _16368_ (.A(net598),
    .B(_06957_),
    .Y(_07365_));
 sg13g2_a21oi_1 _16369_ (.A1(_07334_),
    .A2(_07363_),
    .Y(_07366_),
    .B1(_07365_));
 sg13g2_nand2_1 _16370_ (.Y(_07367_),
    .A(net939),
    .B(_06957_));
 sg13g2_o21ai_1 _16371_ (.B1(_07367_),
    .Y(_07368_),
    .A1(net939),
    .A2(_06958_));
 sg13g2_a22oi_1 _16372_ (.Y(_07369_),
    .B1(_07368_),
    .B2(net319),
    .A2(_07343_),
    .A1(_06653_));
 sg13g2_o21ai_1 _16373_ (.B1(_07369_),
    .Y(_07370_),
    .A1(net318),
    .A2(_07366_));
 sg13g2_nand2_1 _16374_ (.Y(_07371_),
    .A(_07336_),
    .B(_07370_));
 sg13g2_nand2_1 _16375_ (.Y(_07372_),
    .A(net318),
    .B(_07343_));
 sg13g2_nand4_1 _16376_ (.B(net598),
    .C(_06989_),
    .A(net600),
    .Y(_07373_),
    .D(_06636_));
 sg13g2_o21ai_1 _16377_ (.B1(_07373_),
    .Y(_07374_),
    .A1(net600),
    .A2(_07372_));
 sg13g2_inv_2 _16378_ (.Y(_07375_),
    .A(net1156));
 sg13g2_a21oi_1 _16379_ (.A1(_06957_),
    .A2(_06653_),
    .Y(_07376_),
    .B1(_06960_));
 sg13g2_nor3_1 _16380_ (.A(net625),
    .B(_06958_),
    .C(_07343_),
    .Y(_07377_));
 sg13g2_nor2_1 _16381_ (.A(net598),
    .B(_07363_),
    .Y(_07378_));
 sg13g2_nor2_1 _16382_ (.A(_07377_),
    .B(_07378_),
    .Y(_07379_));
 sg13g2_o21ai_1 _16383_ (.B1(_07379_),
    .Y(_07380_),
    .A1(_07375_),
    .A2(_07376_));
 sg13g2_buf_1 _16384_ (.A(_07302_),
    .X(_07381_));
 sg13g2_a22oi_1 _16385_ (.Y(_07382_),
    .B1(_07380_),
    .B2(_07381_),
    .A2(_07374_),
    .A1(net626));
 sg13g2_a221oi_1 _16386_ (.B2(_07382_),
    .C1(_07357_),
    .B1(_07371_),
    .A1(net624),
    .Y(_07383_),
    .A2(net599));
 sg13g2_o21ai_1 _16387_ (.B1(_07356_),
    .Y(_07384_),
    .A1(net624),
    .A2(net599));
 sg13g2_a221oi_1 _16388_ (.B2(_07384_),
    .C1(_06466_),
    .B1(_07383_),
    .A1(_05811_),
    .Y(_07385_),
    .A2(net59));
 sg13g2_xor2_1 _16389_ (.B(_07351_),
    .A(_07228_),
    .X(_07386_));
 sg13g2_a21oi_1 _16390_ (.A1(_05815_),
    .A2(_07386_),
    .Y(_07387_),
    .B1(net311));
 sg13g2_o21ai_1 _16391_ (.B1(_05355_),
    .Y(_07388_),
    .A1(_05811_),
    .A2(_07274_));
 sg13g2_a221oi_1 _16392_ (.B2(_07274_),
    .C1(_07388_),
    .B1(_07387_),
    .A1(_07360_),
    .Y(_00327_),
    .A2(_07385_));
 sg13g2_buf_2 _16393_ (.A(\grid.cell_15_3.se ),
    .X(_07389_));
 sg13g2_buf_1 _16394_ (.A(_07389_),
    .X(_07390_));
 sg13g2_buf_1 _16395_ (.A(net937),
    .X(_07391_));
 sg13g2_nor4_1 _16396_ (.A(net596),
    .B(net939),
    .C(net947),
    .D(net620),
    .Y(_07392_));
 sg13g2_a221oi_1 _16397_ (.B2(_06958_),
    .C1(_07392_),
    .B1(net958),
    .A1(_07364_),
    .Y(_07393_),
    .A2(net610));
 sg13g2_o21ai_1 _16398_ (.B1(net596),
    .Y(_07394_),
    .A1(_07333_),
    .A2(net947));
 sg13g2_and2_1 _16399_ (.A(_06691_),
    .B(_07394_),
    .X(_07395_));
 sg13g2_buf_1 _16400_ (.A(net596),
    .X(_07396_));
 sg13g2_nor3_1 _16401_ (.A(net307),
    .B(_07334_),
    .C(_07033_),
    .Y(_07397_));
 sg13g2_nand2_1 _16402_ (.Y(_07398_),
    .A(net958),
    .B(net318));
 sg13g2_a22oi_1 _16403_ (.Y(_07399_),
    .B1(_07397_),
    .B2(_07398_),
    .A2(_07395_),
    .A1(_07393_));
 sg13g2_buf_1 _16404_ (.A(_00227_),
    .X(_07400_));
 sg13g2_nand2_1 _16405_ (.Y(_07401_),
    .A(net319),
    .B(net1155));
 sg13g2_xnor2_1 _16406_ (.Y(_07402_),
    .A(net937),
    .B(_07006_));
 sg13g2_xor2_1 _16407_ (.B(net959),
    .A(net1156),
    .X(_07403_));
 sg13g2_xnor2_1 _16408_ (.Y(_07404_),
    .A(_07402_),
    .B(_07403_));
 sg13g2_xnor2_1 _16409_ (.Y(_07405_),
    .A(net613),
    .B(_07404_));
 sg13g2_inv_1 _16410_ (.Y(_07406_),
    .A(net1155));
 sg13g2_nand2_1 _16411_ (.Y(_07407_),
    .A(net625),
    .B(_07406_));
 sg13g2_o21ai_1 _16412_ (.B1(_07407_),
    .Y(_07408_),
    .A1(net1162),
    .A2(_07404_));
 sg13g2_a21oi_1 _16413_ (.A1(_07401_),
    .A2(_07405_),
    .Y(_07409_),
    .B1(_07408_));
 sg13g2_xnor2_1 _16414_ (.Y(_07410_),
    .A(_07399_),
    .B(_07409_));
 sg13g2_nor2_1 _16415_ (.A(_07018_),
    .B(_07404_),
    .Y(_07411_));
 sg13g2_and2_1 _16416_ (.A(_07406_),
    .B(_06907_),
    .X(_07412_));
 sg13g2_nand2_1 _16417_ (.Y(_07413_),
    .A(_07364_),
    .B(net610));
 sg13g2_xnor2_1 _16418_ (.Y(_07414_),
    .A(_07014_),
    .B(net623));
 sg13g2_nor2_1 _16419_ (.A(_07375_),
    .B(_07414_),
    .Y(_07415_));
 sg13g2_nor3_1 _16420_ (.A(_07333_),
    .B(_06999_),
    .C(_06958_),
    .Y(_07416_));
 sg13g2_o21ai_1 _16421_ (.B1(net622),
    .Y(_07417_),
    .A1(_07415_),
    .A2(_07416_));
 sg13g2_o21ai_1 _16422_ (.B1(_07417_),
    .Y(_07418_),
    .A1(_06691_),
    .A2(_07413_));
 sg13g2_nor3_1 _16423_ (.A(net307),
    .B(_07398_),
    .C(_07413_),
    .Y(_07419_));
 sg13g2_a221oi_1 _16424_ (.B2(_07396_),
    .C1(_07419_),
    .B1(_07418_),
    .A1(_07411_),
    .Y(_07420_),
    .A2(_07412_));
 sg13g2_a21oi_1 _16425_ (.A1(_07410_),
    .A2(_07420_),
    .Y(_07421_),
    .B1(net106));
 sg13g2_xnor2_1 _16426_ (.Y(_07422_),
    .A(_07280_),
    .B(_07404_));
 sg13g2_a21oi_1 _16427_ (.A1(_05739_),
    .A2(_07422_),
    .Y(_07423_),
    .B1(net310));
 sg13g2_or4_1 _16428_ (.A(net1057),
    .B(net59),
    .C(_07421_),
    .D(_07423_),
    .X(_07424_));
 sg13g2_o21ai_1 _16429_ (.B1(_07424_),
    .Y(_00328_),
    .A1(net26),
    .A2(_07274_));
 sg13g2_a21o_1 _16430_ (.A2(_04938_),
    .A1(net376),
    .B1(_04939_),
    .X(_07425_));
 sg13g2_buf_2 _16431_ (.A(_07425_),
    .X(_07426_));
 sg13g2_nand2_1 _16432_ (.Y(_07427_),
    .A(_07426_),
    .B(net59));
 sg13g2_buf_2 _16433_ (.A(_00049_),
    .X(_07428_));
 sg13g2_buf_1 _16434_ (.A(\grid.cell_15_4.se ),
    .X(_07429_));
 sg13g2_buf_1 _16435_ (.A(_07429_),
    .X(_07430_));
 sg13g2_xor2_1 _16436_ (.B(net1166),
    .A(_07389_),
    .X(_07431_));
 sg13g2_xnor2_1 _16437_ (.Y(_07432_),
    .A(_07156_),
    .B(_07431_));
 sg13g2_xnor2_1 _16438_ (.Y(_07433_),
    .A(net936),
    .B(_07432_));
 sg13g2_buf_1 _16439_ (.A(_07433_),
    .X(_07434_));
 sg13g2_o21ai_1 _16440_ (.B1(_06958_),
    .Y(_07435_),
    .A1(net611),
    .A2(_07434_));
 sg13g2_nor2_1 _16441_ (.A(net1160),
    .B(net623),
    .Y(_07436_));
 sg13g2_or2_1 _16442_ (.X(_07437_),
    .B(_07436_),
    .A(_07434_));
 sg13g2_a221oi_1 _16443_ (.B2(_06989_),
    .C1(_06961_),
    .B1(_07437_),
    .A1(net1160),
    .Y(_07438_),
    .A2(_07435_));
 sg13g2_xnor2_1 _16444_ (.Y(_07439_),
    .A(net611),
    .B(_07434_));
 sg13g2_nor2_1 _16445_ (.A(_07052_),
    .B(_07434_),
    .Y(_07440_));
 sg13g2_a22oi_1 _16446_ (.Y(_07441_),
    .B1(_07440_),
    .B2(_07428_),
    .A2(_07439_),
    .A1(net318));
 sg13g2_o21ai_1 _16447_ (.B1(_07441_),
    .Y(_07442_),
    .A1(_07428_),
    .A2(_07438_));
 sg13g2_inv_1 _16448_ (.Y(_07443_),
    .A(net936));
 sg13g2_nor2_1 _16449_ (.A(net596),
    .B(net946),
    .Y(_07444_));
 sg13g2_nand2_1 _16450_ (.Y(_07445_),
    .A(_07443_),
    .B(_07444_));
 sg13g2_nand3_1 _16451_ (.B(net621),
    .C(_07444_),
    .A(_07443_),
    .Y(_07446_));
 sg13g2_buf_1 _16452_ (.A(net936),
    .X(_07447_));
 sg13g2_buf_1 _16453_ (.A(net595),
    .X(_07448_));
 sg13g2_o21ai_1 _16454_ (.B1(net608),
    .Y(_07449_),
    .A1(net306),
    .A2(net307));
 sg13g2_and2_1 _16455_ (.A(net936),
    .B(net937),
    .X(_07450_));
 sg13g2_buf_1 _16456_ (.A(_07450_),
    .X(_07451_));
 sg13g2_a21oi_1 _16457_ (.A1(net621),
    .A2(net620),
    .Y(_07452_),
    .B1(_07451_));
 sg13g2_nand4_1 _16458_ (.B(_07446_),
    .C(_07449_),
    .A(_06721_),
    .Y(_07453_),
    .D(_07452_));
 sg13g2_o21ai_1 _16459_ (.B1(_07453_),
    .Y(_07454_),
    .A1(_06681_),
    .A2(_07445_));
 sg13g2_buf_1 _16460_ (.A(net306),
    .X(_07455_));
 sg13g2_nand2_1 _16461_ (.Y(_07456_),
    .A(net596),
    .B(net621));
 sg13g2_o21ai_1 _16462_ (.B1(_07456_),
    .Y(_07457_),
    .A1(_07391_),
    .A2(net609));
 sg13g2_nor2_1 _16463_ (.A(_06743_),
    .B(net620),
    .Y(_07458_));
 sg13g2_a22oi_1 _16464_ (.Y(_07459_),
    .B1(_07457_),
    .B2(_07458_),
    .A2(_07444_),
    .A1(net620));
 sg13g2_inv_1 _16465_ (.Y(_07460_),
    .A(_07428_));
 sg13g2_inv_1 _16466_ (.Y(_07461_),
    .A(_07389_));
 sg13g2_buf_1 _16467_ (.A(_07461_),
    .X(_07462_));
 sg13g2_nor3_1 _16468_ (.A(_06743_),
    .B(_07462_),
    .C(net609),
    .Y(_07463_));
 sg13g2_nor3_1 _16469_ (.A(_06721_),
    .B(net937),
    .C(net1161),
    .Y(_07464_));
 sg13g2_a21oi_1 _16470_ (.A1(net937),
    .A2(net1161),
    .Y(_07465_),
    .B1(_06681_));
 sg13g2_nor3_1 _16471_ (.A(_07463_),
    .B(_07464_),
    .C(_07465_),
    .Y(_07466_));
 sg13g2_mux2_1 _16472_ (.A0(_06721_),
    .A1(_07443_),
    .S(net620),
    .X(_07467_));
 sg13g2_nor4_1 _16473_ (.A(net594),
    .B(net609),
    .C(_06677_),
    .D(_07467_),
    .Y(_07468_));
 sg13g2_a221oi_1 _16474_ (.B2(net306),
    .C1(_07468_),
    .B1(_07466_),
    .A1(_07460_),
    .Y(_07469_),
    .A2(net623));
 sg13g2_o21ai_1 _16475_ (.B1(_07469_),
    .Y(_07470_),
    .A1(net152),
    .A2(_07459_));
 sg13g2_a21oi_1 _16476_ (.A1(_07391_),
    .A2(net946),
    .Y(_07471_),
    .B1(net306));
 sg13g2_o21ai_1 _16477_ (.B1(_06721_),
    .Y(_07472_),
    .A1(_07444_),
    .A2(_07471_));
 sg13g2_a21oi_1 _16478_ (.A1(_07445_),
    .A2(_07472_),
    .Y(_07473_),
    .B1(net316));
 sg13g2_nor3_1 _16479_ (.A(_07440_),
    .B(_07470_),
    .C(_07473_),
    .Y(_07474_));
 sg13g2_o21ai_1 _16480_ (.B1(_07439_),
    .Y(_07475_),
    .A1(_07460_),
    .A2(net318));
 sg13g2_a221oi_1 _16481_ (.B2(_07475_),
    .C1(net100),
    .B1(_07474_),
    .A1(_07442_),
    .Y(_07476_),
    .A2(_07454_));
 sg13g2_xnor2_1 _16482_ (.Y(_07477_),
    .A(_07348_),
    .B(_07434_));
 sg13g2_a21oi_1 _16483_ (.A1(net109),
    .A2(_07477_),
    .Y(_07478_),
    .B1(net610));
 sg13g2_or3_1 _16484_ (.A(_07201_),
    .B(_07476_),
    .C(_07478_),
    .X(_07479_));
 sg13g2_buf_1 _16485_ (.A(_00669_),
    .X(_07480_));
 sg13g2_a21oi_1 _16486_ (.A1(_07427_),
    .A2(_07479_),
    .Y(_00329_),
    .B1(net305));
 sg13g2_nand2_1 _16487_ (.Y(_07481_),
    .A(_06330_),
    .B(net59));
 sg13g2_buf_1 _16488_ (.A(\grid.cell_15_5.se ),
    .X(_07482_));
 sg13g2_buf_1 _16489_ (.A(_07482_),
    .X(_07483_));
 sg13g2_buf_1 _16490_ (.A(net935),
    .X(_07484_));
 sg13g2_nor4_1 _16491_ (.A(_07484_),
    .B(net595),
    .C(net944),
    .D(net618),
    .Y(_07485_));
 sg13g2_inv_2 _16492_ (.Y(_07486_),
    .A(net935));
 sg13g2_a21oi_1 _16493_ (.A1(_07486_),
    .A2(_07443_),
    .Y(_07487_),
    .B1(net606));
 sg13g2_nand2_1 _16494_ (.Y(_07488_),
    .A(net593),
    .B(net595));
 sg13g2_o21ai_1 _16495_ (.B1(_07488_),
    .Y(_07489_),
    .A1(net618),
    .A2(net621));
 sg13g2_nor3_1 _16496_ (.A(_07485_),
    .B(_07487_),
    .C(_07489_),
    .Y(_07490_));
 sg13g2_buf_1 _16497_ (.A(net593),
    .X(_07491_));
 sg13g2_nor3_1 _16498_ (.A(net304),
    .B(net152),
    .C(net945),
    .Y(_07492_));
 sg13g2_nand2_1 _16499_ (.Y(_07493_),
    .A(net315),
    .B(net621));
 sg13g2_a22oi_1 _16500_ (.Y(_07494_),
    .B1(_07492_),
    .B2(_07493_),
    .A2(_07490_),
    .A1(_06784_));
 sg13g2_buf_1 _16501_ (.A(_00081_),
    .X(_07495_));
 sg13g2_nand2_1 _16502_ (.Y(_07496_),
    .A(net1154),
    .B(net620));
 sg13g2_xor2_1 _16503_ (.B(_06670_),
    .A(net936),
    .X(_07497_));
 sg13g2_xnor2_1 _16504_ (.Y(_07498_),
    .A(_07078_),
    .B(_07497_));
 sg13g2_xnor2_1 _16505_ (.Y(_07499_),
    .A(net935),
    .B(_07498_));
 sg13g2_xnor2_1 _16506_ (.Y(_07500_),
    .A(net610),
    .B(_07499_));
 sg13g2_nand2b_1 _16507_ (.Y(_07501_),
    .B(net958),
    .A_N(net1154));
 sg13g2_o21ai_1 _16508_ (.B1(_07501_),
    .Y(_07502_),
    .A1(_07082_),
    .A2(_07499_));
 sg13g2_a21oi_1 _16509_ (.A1(_07496_),
    .A2(_07500_),
    .Y(_07503_),
    .B1(_07502_));
 sg13g2_xnor2_1 _16510_ (.Y(_07504_),
    .A(_07494_),
    .B(_07503_));
 sg13g2_buf_1 _16511_ (.A(net304),
    .X(_07505_));
 sg13g2_xor2_1 _16512_ (.B(net621),
    .A(net944),
    .X(_07506_));
 sg13g2_nor3_1 _16513_ (.A(net306),
    .B(_07102_),
    .C(_06677_),
    .Y(_07507_));
 sg13g2_a21oi_1 _16514_ (.A1(_07448_),
    .A2(_07506_),
    .Y(_07508_),
    .B1(_07507_));
 sg13g2_nand3_1 _16515_ (.B(_07455_),
    .C(net945),
    .A(_06785_),
    .Y(_07509_));
 sg13g2_o21ai_1 _16516_ (.B1(_07509_),
    .Y(_07510_),
    .A1(net618),
    .A2(_07508_));
 sg13g2_nand2b_1 _16517_ (.Y(_07511_),
    .B(net1159),
    .A_N(_07483_));
 sg13g2_nor2_1 _16518_ (.A(_07493_),
    .B(_07511_),
    .Y(_07512_));
 sg13g2_nand2b_1 _16519_ (.Y(_07513_),
    .B(_07006_),
    .A_N(_07495_));
 sg13g2_nor3_1 _16520_ (.A(_07082_),
    .B(_07499_),
    .C(_07513_),
    .Y(_07514_));
 sg13g2_a221oi_1 _16521_ (.B2(_07455_),
    .C1(_07514_),
    .B1(_07512_),
    .A1(net151),
    .Y(_07515_),
    .A2(_07510_));
 sg13g2_a21oi_1 _16522_ (.A1(_07504_),
    .A2(_07515_),
    .Y(_07516_),
    .B1(net102));
 sg13g2_xnor2_1 _16523_ (.Y(_07517_),
    .A(_07402_),
    .B(_07499_));
 sg13g2_a21oi_1 _16524_ (.A1(net109),
    .A2(_07517_),
    .Y(_07518_),
    .B1(net608));
 sg13g2_or3_1 _16525_ (.A(net59),
    .B(_07516_),
    .C(_07518_),
    .X(_07519_));
 sg13g2_a21oi_1 _16526_ (.A1(_07481_),
    .A2(_07519_),
    .Y(_00330_),
    .B1(net305));
 sg13g2_buf_1 _16527_ (.A(_00143_),
    .X(_07520_));
 sg13g2_nand2_1 _16528_ (.Y(_07521_),
    .A(net619),
    .B(net314));
 sg13g2_nor2_1 _16529_ (.A(_07521_),
    .B(_07214_),
    .Y(_07522_));
 sg13g2_o21ai_1 _16530_ (.B1(_07522_),
    .Y(_07523_),
    .A1(net1153),
    .A2(_07241_));
 sg13g2_o21ai_1 _16531_ (.B1(_07523_),
    .Y(_07524_),
    .A1(net1153),
    .A2(_07258_));
 sg13g2_o21ai_1 _16532_ (.B1(_07241_),
    .Y(_07525_),
    .A1(net304),
    .A2(_07214_));
 sg13g2_nor2_1 _16533_ (.A(net593),
    .B(_07241_),
    .Y(_07526_));
 sg13g2_a21oi_1 _16534_ (.A1(net1153),
    .A2(_07525_),
    .Y(_07527_),
    .B1(_07526_));
 sg13g2_nor2b_1 _16535_ (.A(net593),
    .B_N(_07520_),
    .Y(_07528_));
 sg13g2_nand2_1 _16536_ (.Y(_07529_),
    .A(_07208_),
    .B(net627));
 sg13g2_nand2_1 _16537_ (.Y(_07530_),
    .A(_07247_),
    .B(_07529_));
 sg13g2_nor2_1 _16538_ (.A(net1153),
    .B(net603),
    .Y(_07531_));
 sg13g2_a22oi_1 _16539_ (.Y(_07532_),
    .B1(_07531_),
    .B2(net155),
    .A2(_07530_),
    .A1(_07528_));
 sg13g2_nor2_1 _16540_ (.A(_07486_),
    .B(net603),
    .Y(_07533_));
 sg13g2_a21oi_1 _16541_ (.A1(net155),
    .A2(_07533_),
    .Y(_07534_),
    .B1(_07526_));
 sg13g2_mux2_1 _16542_ (.A0(_07532_),
    .A1(_07534_),
    .S(net618),
    .X(_07535_));
 sg13g2_o21ai_1 _16543_ (.B1(_07535_),
    .Y(_07536_),
    .A1(net156),
    .A2(_07527_));
 sg13g2_a21oi_1 _16544_ (.A1(net151),
    .A2(_07524_),
    .Y(_07537_),
    .B1(_07536_));
 sg13g2_buf_1 _16545_ (.A(_00113_),
    .X(_07538_));
 sg13g2_inv_1 _16546_ (.Y(_07539_),
    .A(_07538_));
 sg13g2_xnor2_1 _16547_ (.Y(_07540_),
    .A(_06786_),
    .B(_07216_));
 sg13g2_xnor2_1 _16548_ (.Y(_07541_),
    .A(net593),
    .B(_07540_));
 sg13g2_xnor2_1 _16549_ (.Y(_07542_),
    .A(_07044_),
    .B(_07541_));
 sg13g2_o21ai_1 _16550_ (.B1(_07542_),
    .Y(_07543_),
    .A1(_07539_),
    .A2(net316));
 sg13g2_and2_1 _16551_ (.A(_07138_),
    .B(_07541_),
    .X(_07544_));
 sg13g2_a21oi_1 _16552_ (.A1(_07539_),
    .A2(net316),
    .Y(_07545_),
    .B1(_07544_));
 sg13g2_nand2_1 _16553_ (.Y(_07546_),
    .A(_07543_),
    .B(_07545_));
 sg13g2_xor2_1 _16554_ (.B(_07546_),
    .A(_07537_),
    .X(_07547_));
 sg13g2_xnor2_1 _16555_ (.Y(_07548_),
    .A(net313),
    .B(net619));
 sg13g2_o21ai_1 _16556_ (.B1(net156),
    .Y(_07549_),
    .A1(net309),
    .A2(_07176_));
 sg13g2_a21o_1 _16557_ (.A2(_07548_),
    .A1(_07211_),
    .B1(_07549_),
    .X(_07550_));
 sg13g2_o21ai_1 _16558_ (.B1(_07550_),
    .Y(_07551_),
    .A1(net1153),
    .A2(_07258_));
 sg13g2_nor2_1 _16559_ (.A(net151),
    .B(_07529_),
    .Y(_07552_));
 sg13g2_buf_1 _16560_ (.A(net163),
    .X(_07553_));
 sg13g2_a221oi_1 _16561_ (.B2(_07176_),
    .C1(net99),
    .B1(_07552_),
    .A1(net151),
    .Y(_07554_),
    .A2(_07551_));
 sg13g2_nand3_1 _16562_ (.B(_07156_),
    .C(_07544_),
    .A(_07539_),
    .Y(_07555_));
 sg13g2_xnor2_1 _16563_ (.Y(_07556_),
    .A(_07448_),
    .B(net608));
 sg13g2_xnor2_1 _16564_ (.Y(_07557_),
    .A(net316),
    .B(_07556_));
 sg13g2_xnor2_1 _16565_ (.Y(_07558_),
    .A(_07541_),
    .B(_07557_));
 sg13g2_nand2_1 _16566_ (.Y(_07559_),
    .A(net606),
    .B(_07558_));
 sg13g2_nand4_1 _16567_ (.B(_07554_),
    .C(_07555_),
    .A(_07547_),
    .Y(_07560_),
    .D(_07559_));
 sg13g2_buf_1 _16568_ (.A(net120),
    .X(_07561_));
 sg13g2_buf_1 _16569_ (.A(_06810_),
    .X(_07562_));
 sg13g2_a22oi_1 _16570_ (.Y(_07563_),
    .B1(net25),
    .B2(_07273_),
    .A2(net71),
    .A1(net607));
 sg13g2_a221oi_1 _16571_ (.B2(_07563_),
    .C1(net617),
    .B1(_07560_),
    .A1(net24),
    .Y(_00331_),
    .A2(_07273_));
 sg13g2_xnor2_1 _16572_ (.Y(_07564_),
    .A(net935),
    .B(_07207_));
 sg13g2_xnor2_1 _16573_ (.Y(_07565_),
    .A(_07078_),
    .B(_07564_));
 sg13g2_xnor2_1 _16574_ (.Y(_07566_),
    .A(net627),
    .B(_07565_));
 sg13g2_xor2_1 _16575_ (.B(_07566_),
    .A(net953),
    .X(_07567_));
 sg13g2_a221oi_1 _16576_ (.B2(_07324_),
    .C1(_07316_),
    .B1(_07567_),
    .A1(_06921_),
    .Y(_07568_),
    .A2(_07566_));
 sg13g2_nor2_1 _16577_ (.A(_07244_),
    .B(net606),
    .Y(_07569_));
 sg13g2_nand2_1 _16578_ (.Y(_07570_),
    .A(_07244_),
    .B(net606));
 sg13g2_o21ai_1 _16579_ (.B1(_07570_),
    .Y(_07571_),
    .A1(_07491_),
    .A2(_07569_));
 sg13g2_nor2_1 _16580_ (.A(_07491_),
    .B(_07570_),
    .Y(_07572_));
 sg13g2_a21oi_1 _16581_ (.A1(net1153),
    .A2(_07571_),
    .Y(_07573_),
    .B1(_07572_));
 sg13g2_or2_1 _16582_ (.X(_07574_),
    .B(_07573_),
    .A(net156));
 sg13g2_nand2_1 _16583_ (.Y(_07575_),
    .A(_07209_),
    .B(net944));
 sg13g2_nor2_1 _16584_ (.A(net1153),
    .B(_07575_),
    .Y(_07576_));
 sg13g2_nor2_1 _16585_ (.A(net1153),
    .B(_07570_),
    .Y(_07577_));
 sg13g2_nor3_1 _16586_ (.A(_07521_),
    .B(_07569_),
    .C(_07577_),
    .Y(_07578_));
 sg13g2_o21ai_1 _16587_ (.B1(_07505_),
    .Y(_07579_),
    .A1(_07576_),
    .A2(_07578_));
 sg13g2_o21ai_1 _16588_ (.B1(_07529_),
    .Y(_07580_),
    .A1(_07209_),
    .A2(net606));
 sg13g2_and2_1 _16589_ (.A(net944),
    .B(net314),
    .X(_07581_));
 sg13g2_a22oi_1 _16590_ (.Y(_07582_),
    .B1(_07581_),
    .B2(_07531_),
    .A2(_07580_),
    .A1(_07528_));
 sg13g2_a21oi_1 _16591_ (.A1(_07533_),
    .A2(_07581_),
    .Y(_07583_),
    .B1(_07572_));
 sg13g2_mux2_1 _16592_ (.A0(_07582_),
    .A1(_07583_),
    .S(net618),
    .X(_07584_));
 sg13g2_nand3_1 _16593_ (.B(_07579_),
    .C(_07584_),
    .A(_07574_),
    .Y(_07585_));
 sg13g2_xor2_1 _16594_ (.B(_07585_),
    .A(_07568_),
    .X(_07586_));
 sg13g2_xnor2_1 _16595_ (.Y(_07587_),
    .A(net1167),
    .B(net953));
 sg13g2_and4_1 _16596_ (.A(_07234_),
    .B(_06921_),
    .C(_07566_),
    .D(_07587_),
    .X(_07588_));
 sg13g2_nand2b_1 _16597_ (.Y(_07589_),
    .B(net309),
    .A_N(_07078_));
 sg13g2_o21ai_1 _16598_ (.B1(_07589_),
    .Y(_07590_),
    .A1(_07210_),
    .A2(_07099_));
 sg13g2_a21oi_1 _16599_ (.A1(net156),
    .A2(_07590_),
    .Y(_07591_),
    .B1(_07576_));
 sg13g2_nor2_1 _16600_ (.A(_07486_),
    .B(_07591_),
    .Y(_07592_));
 sg13g2_nor3_1 _16601_ (.A(_07505_),
    .B(_07521_),
    .C(_07575_),
    .Y(_07593_));
 sg13g2_nor4_1 _16602_ (.A(net125),
    .B(_07588_),
    .C(_07592_),
    .D(_07593_),
    .Y(_07594_));
 sg13g2_xnor2_1 _16603_ (.Y(_07595_),
    .A(_07328_),
    .B(_07566_));
 sg13g2_nand2b_1 _16604_ (.Y(_07596_),
    .B(_07595_),
    .A_N(net154));
 sg13g2_nand3_1 _16605_ (.B(_07594_),
    .C(_07596_),
    .A(_07586_),
    .Y(_07597_));
 sg13g2_a22oi_1 _16606_ (.Y(_07598_),
    .B1(net76),
    .B2(_07273_),
    .A2(net71),
    .A1(_07147_));
 sg13g2_a221oi_1 _16607_ (.B2(_07598_),
    .C1(net617),
    .B1(_07597_),
    .A1(_06471_),
    .Y(_00332_),
    .A2(_07273_));
 sg13g2_or2_1 _16608_ (.X(_07599_),
    .B(net320),
    .A(_01935_));
 sg13g2_buf_2 _16609_ (.A(_07599_),
    .X(_07600_));
 sg13g2_or2_1 _16610_ (.X(_07601_),
    .B(net177),
    .A(_01870_));
 sg13g2_buf_2 _16611_ (.A(_07601_),
    .X(_07602_));
 sg13g2_nor2_1 _16612_ (.A(_07600_),
    .B(_07602_),
    .Y(_07603_));
 sg13g2_nand2_1 _16613_ (.Y(_07604_),
    .A(net158),
    .B(_07603_));
 sg13g2_buf_1 _16614_ (.A(_07604_),
    .X(_07605_));
 sg13g2_nand3_1 _16615_ (.B(_06425_),
    .C(_07605_),
    .A(net941),
    .Y(_07606_));
 sg13g2_o21ai_1 _16616_ (.B1(_07606_),
    .Y(_07607_),
    .A1(net50),
    .A2(_07605_));
 sg13g2_buf_2 _16617_ (.A(\grid.cell_16_0.sw ),
    .X(_07608_));
 sg13g2_buf_1 _16618_ (.A(_07608_),
    .X(_07609_));
 sg13g2_buf_1 _16619_ (.A(\grid.cell_16_0.se ),
    .X(_07610_));
 sg13g2_xnor2_1 _16620_ (.Y(_07611_),
    .A(net1165),
    .B(net1152));
 sg13g2_xnor2_1 _16621_ (.Y(_07612_),
    .A(net934),
    .B(_07611_));
 sg13g2_xnor2_1 _16622_ (.Y(_07613_),
    .A(_07216_),
    .B(_07612_));
 sg13g2_buf_1 _16623_ (.A(\grid.cell_16_0.s ),
    .X(_07614_));
 sg13g2_buf_1 _16624_ (.A(_07614_),
    .X(_07615_));
 sg13g2_xor2_1 _16625_ (.B(_07204_),
    .A(_06856_),
    .X(_07616_));
 sg13g2_xnor2_1 _16626_ (.Y(_07617_),
    .A(net933),
    .B(_07616_));
 sg13g2_xnor2_1 _16627_ (.Y(_07618_),
    .A(_07613_),
    .B(_07617_));
 sg13g2_a21oi_1 _16628_ (.A1(_06057_),
    .A2(_07618_),
    .Y(_07619_),
    .B1(net941));
 sg13g2_buf_1 _16629_ (.A(net934),
    .X(_07620_));
 sg13g2_nand2_2 _16630_ (.Y(_07621_),
    .A(net592),
    .B(net604));
 sg13g2_nor2_1 _16631_ (.A(net592),
    .B(_07229_),
    .Y(_07622_));
 sg13g2_inv_1 _16632_ (.Y(_07623_),
    .A(net934));
 sg13g2_buf_1 _16633_ (.A(_07623_),
    .X(_07624_));
 sg13g2_nor2_1 _16634_ (.A(net303),
    .B(net604),
    .Y(_07625_));
 sg13g2_o21ai_1 _16635_ (.B1(net954),
    .Y(_07626_),
    .A1(_07622_),
    .A2(_07625_));
 sg13g2_o21ai_1 _16636_ (.B1(_07626_),
    .Y(_07627_),
    .A1(net954),
    .A2(_07621_));
 sg13g2_nand2_1 _16637_ (.Y(_07628_),
    .A(net604),
    .B(_06979_));
 sg13g2_nor2_1 _16638_ (.A(_07624_),
    .B(_07628_),
    .Y(_07629_));
 sg13g2_a21oi_1 _16639_ (.A1(net154),
    .A2(_07627_),
    .Y(_07630_),
    .B1(_07629_));
 sg13g2_buf_1 _16640_ (.A(_07610_),
    .X(_07631_));
 sg13g2_buf_1 _16641_ (.A(net932),
    .X(_07632_));
 sg13g2_nand2b_1 _16642_ (.Y(_07633_),
    .B(net591),
    .A_N(_07630_));
 sg13g2_nor2_1 _16643_ (.A(net1152),
    .B(_07624_),
    .Y(_07634_));
 sg13g2_nand3_1 _16644_ (.B(_07214_),
    .C(_07634_),
    .A(net612),
    .Y(_07635_));
 sg13g2_nand4_1 _16645_ (.B(_07605_),
    .C(_07633_),
    .A(net1060),
    .Y(_07636_),
    .D(_07635_));
 sg13g2_buf_2 _16646_ (.A(_00226_),
    .X(_07637_));
 sg13g2_nand2_1 _16647_ (.Y(_07638_),
    .A(net599),
    .B(_07613_));
 sg13g2_nor3_1 _16648_ (.A(_07637_),
    .B(_07616_),
    .C(_07638_),
    .Y(_07639_));
 sg13g2_buf_1 _16649_ (.A(_07620_),
    .X(_07640_));
 sg13g2_buf_1 _16650_ (.A(net302),
    .X(_07641_));
 sg13g2_a21oi_1 _16651_ (.A1(net150),
    .A2(_07628_),
    .Y(_07642_),
    .B1(_07622_));
 sg13g2_a21o_1 _16652_ (.A2(net313),
    .A1(net303),
    .B1(_07625_),
    .X(_07643_));
 sg13g2_or2_1 _16653_ (.X(_07644_),
    .B(net942),
    .A(_07608_));
 sg13g2_buf_1 _16654_ (.A(_07644_),
    .X(_07645_));
 sg13g2_nor2_1 _16655_ (.A(net949),
    .B(_07645_),
    .Y(_07646_));
 sg13g2_a21oi_1 _16656_ (.A1(net616),
    .A2(_07643_),
    .Y(_07647_),
    .B1(_07646_));
 sg13g2_o21ai_1 _16657_ (.B1(_07647_),
    .Y(_07648_),
    .A1(net154),
    .A2(_07642_));
 sg13g2_nor2b_1 _16658_ (.A(net954),
    .B_N(net313),
    .Y(_07649_));
 sg13g2_o21ai_1 _16659_ (.B1(_07243_),
    .Y(_07650_),
    .A1(net309),
    .A2(net949));
 sg13g2_nor2_1 _16660_ (.A(net302),
    .B(_07628_),
    .Y(_07651_));
 sg13g2_a221oi_1 _16661_ (.B2(net150),
    .C1(_07651_),
    .B1(_07650_),
    .A1(_07645_),
    .Y(_07652_),
    .A2(_07649_));
 sg13g2_buf_1 _16662_ (.A(net1152),
    .X(_07653_));
 sg13g2_nor3_1 _16663_ (.A(_07653_),
    .B(net302),
    .C(_07247_),
    .Y(_07654_));
 sg13g2_nand2_1 _16664_ (.Y(_07655_),
    .A(net1152),
    .B(net592));
 sg13g2_nor3_1 _16665_ (.A(net603),
    .B(_06979_),
    .C(_07655_),
    .Y(_07656_));
 sg13g2_o21ai_1 _16666_ (.B1(net954),
    .Y(_07657_),
    .A1(_07654_),
    .A2(_07656_));
 sg13g2_o21ai_1 _16667_ (.B1(_07657_),
    .Y(_07658_),
    .A1(net591),
    .A2(_07652_));
 sg13g2_a21oi_1 _16668_ (.A1(net591),
    .A2(_07648_),
    .Y(_07659_),
    .B1(_07658_));
 sg13g2_nand2b_1 _16669_ (.Y(_07660_),
    .B(net953),
    .A_N(_07637_));
 sg13g2_xnor2_1 _16670_ (.Y(_07661_),
    .A(net943),
    .B(_07613_));
 sg13g2_nand2b_1 _16671_ (.Y(_07662_),
    .B(_07637_),
    .A_N(_06856_));
 sg13g2_nand2b_1 _16672_ (.Y(_07663_),
    .B(_07662_),
    .A_N(_07661_));
 sg13g2_nand3_1 _16673_ (.B(_07660_),
    .C(_07663_),
    .A(_07638_),
    .Y(_07664_));
 sg13g2_xor2_1 _16674_ (.B(_07664_),
    .A(_07659_),
    .X(_07665_));
 sg13g2_nor4_1 _16675_ (.A(_07619_),
    .B(_07636_),
    .C(_07639_),
    .D(_07665_),
    .Y(_07666_));
 sg13g2_a21o_1 _16676_ (.A2(_07607_),
    .A1(_06667_),
    .B1(_07666_),
    .X(_00333_));
 sg13g2_buf_1 _16677_ (.A(\grid.cell_16_1.se ),
    .X(_07667_));
 sg13g2_buf_1 _16678_ (.A(net1151),
    .X(_07668_));
 sg13g2_buf_1 _16679_ (.A(net930),
    .X(_07669_));
 sg13g2_or3_1 _16680_ (.A(_07653_),
    .B(net600),
    .C(net590),
    .X(_07670_));
 sg13g2_nand4_1 _16681_ (.B(net613),
    .C(net600),
    .A(net932),
    .Y(_07671_),
    .D(net590));
 sg13g2_a21oi_1 _16682_ (.A1(_07670_),
    .A2(_07671_),
    .Y(_07672_),
    .B1(net612));
 sg13g2_buf_1 _16683_ (.A(_07669_),
    .X(_07673_));
 sg13g2_nor4_1 _16684_ (.A(net311),
    .B(net308),
    .C(_07673_),
    .D(_06979_),
    .Y(_07674_));
 sg13g2_nand2_1 _16685_ (.Y(_07675_),
    .A(net1165),
    .B(net952));
 sg13g2_nand2b_1 _16686_ (.Y(_07676_),
    .B(net1151),
    .A_N(_06971_));
 sg13g2_o21ai_1 _16687_ (.B1(_07676_),
    .Y(_07677_),
    .A1(net930),
    .A2(_07675_));
 sg13g2_nor2_1 _16688_ (.A(net930),
    .B(net949),
    .Y(_07678_));
 sg13g2_nor3_1 _16689_ (.A(net600),
    .B(_07675_),
    .C(_07678_),
    .Y(_07679_));
 sg13g2_a21oi_1 _16690_ (.A1(_07335_),
    .A2(_07677_),
    .Y(_07680_),
    .B1(_07679_));
 sg13g2_nor2b_1 _16691_ (.A(_07680_),
    .B_N(net591),
    .Y(_07681_));
 sg13g2_nand2_1 _16692_ (.Y(_07682_),
    .A(_07302_),
    .B(_07676_));
 sg13g2_o21ai_1 _16693_ (.B1(_07682_),
    .Y(_07683_),
    .A1(net590),
    .A2(_06979_));
 sg13g2_nand2_1 _16694_ (.Y(_07684_),
    .A(net930),
    .B(net949));
 sg13g2_o21ai_1 _16695_ (.B1(net940),
    .Y(_07685_),
    .A1(net930),
    .A2(net949));
 sg13g2_a21oi_1 _16696_ (.A1(_07684_),
    .A2(_07685_),
    .Y(_07686_),
    .B1(_07675_));
 sg13g2_a21oi_1 _16697_ (.A1(net951),
    .A2(_07683_),
    .Y(_07687_),
    .B1(_07686_));
 sg13g2_nor2_1 _16698_ (.A(net591),
    .B(_07687_),
    .Y(_07688_));
 sg13g2_nor4_1 _16699_ (.A(_07672_),
    .B(_07674_),
    .C(_07681_),
    .D(_07688_),
    .Y(_07689_));
 sg13g2_xor2_1 _16700_ (.B(net1151),
    .A(net1157),
    .X(_07690_));
 sg13g2_xnor2_1 _16701_ (.Y(_07691_),
    .A(net951),
    .B(_07690_));
 sg13g2_xor2_1 _16702_ (.B(_07691_),
    .A(_07611_),
    .X(_07692_));
 sg13g2_xnor2_1 _16703_ (.Y(_07693_),
    .A(net941),
    .B(_07692_));
 sg13g2_o21ai_1 _16704_ (.B1(_07660_),
    .Y(_07694_),
    .A1(net1158),
    .A2(_07692_));
 sg13g2_a21oi_1 _16705_ (.A1(_07662_),
    .A2(_07693_),
    .Y(_07695_),
    .B1(_07694_));
 sg13g2_xnor2_1 _16706_ (.Y(_07696_),
    .A(_07689_),
    .B(_07695_));
 sg13g2_nand2_2 _16707_ (.Y(_07697_),
    .A(net940),
    .B(net590));
 sg13g2_nand2_1 _16708_ (.Y(_07698_),
    .A(net954),
    .B(_07690_));
 sg13g2_o21ai_1 _16709_ (.B1(_07698_),
    .Y(_07699_),
    .A1(net954),
    .A2(_07697_));
 sg13g2_nand2_1 _16710_ (.Y(_07700_),
    .A(net311),
    .B(_07699_));
 sg13g2_o21ai_1 _16711_ (.B1(_07700_),
    .Y(_07701_),
    .A1(net949),
    .A2(_07697_));
 sg13g2_inv_1 _16712_ (.Y(_07702_),
    .A(_07614_));
 sg13g2_xnor2_1 _16713_ (.Y(_07703_),
    .A(_07702_),
    .B(_07327_));
 sg13g2_xor2_1 _16714_ (.B(_07703_),
    .A(_07692_),
    .X(_07704_));
 sg13g2_nor3_1 _16715_ (.A(_07637_),
    .B(net1158),
    .C(_07327_),
    .Y(_07705_));
 sg13g2_nor2b_1 _16716_ (.A(_07692_),
    .B_N(_07705_),
    .Y(_07706_));
 sg13g2_nor3_1 _16717_ (.A(_07632_),
    .B(_07697_),
    .C(_07675_),
    .Y(_07707_));
 sg13g2_or3_1 _16718_ (.A(_05130_),
    .B(_07706_),
    .C(_07707_),
    .X(_07708_));
 sg13g2_a221oi_1 _16719_ (.B2(net602),
    .C1(_07708_),
    .B1(_07704_),
    .A1(_07632_),
    .Y(_07709_),
    .A2(_07701_));
 sg13g2_a22oi_1 _16720_ (.Y(_07710_),
    .B1(_07696_),
    .B2(_07709_),
    .A2(_06538_),
    .A1(net605));
 sg13g2_o21ai_1 _16721_ (.B1(net334),
    .Y(_07711_),
    .A1(_03164_),
    .A2(_07605_));
 sg13g2_a21oi_1 _16722_ (.A1(_07605_),
    .A2(_07710_),
    .Y(_00334_),
    .B1(_07711_));
 sg13g2_nor3_1 _16723_ (.A(_07600_),
    .B(_02032_),
    .C(_07602_),
    .Y(_07712_));
 sg13g2_buf_1 _16724_ (.A(_07712_),
    .X(_07713_));
 sg13g2_nand2_1 _16725_ (.Y(_07714_),
    .A(net33),
    .B(_07713_));
 sg13g2_buf_2 _16726_ (.A(_00225_),
    .X(_07715_));
 sg13g2_inv_2 _16727_ (.Y(_07716_),
    .A(_07715_));
 sg13g2_buf_2 _16728_ (.A(\grid.cell_16_2.se ),
    .X(_07717_));
 sg13g2_buf_1 _16729_ (.A(net1150),
    .X(_07718_));
 sg13g2_nand2_1 _16730_ (.Y(_07719_),
    .A(net929),
    .B(net1156));
 sg13g2_xnor2_1 _16731_ (.Y(_07720_),
    .A(_07717_),
    .B(_07332_));
 sg13g2_nor2_1 _16732_ (.A(net951),
    .B(_07720_),
    .Y(_07721_));
 sg13g2_nor2_1 _16733_ (.A(net952),
    .B(_07719_),
    .Y(_07722_));
 sg13g2_o21ai_1 _16734_ (.B1(net611),
    .Y(_07723_),
    .A1(_07721_),
    .A2(_07722_));
 sg13g2_o21ai_1 _16735_ (.B1(_07723_),
    .Y(_07724_),
    .A1(net1162),
    .A2(_07719_));
 sg13g2_nand2_1 _16736_ (.Y(_07725_),
    .A(net613),
    .B(net611));
 sg13g2_nor3_1 _16737_ (.A(_07669_),
    .B(_07725_),
    .C(_07719_),
    .Y(_07726_));
 sg13g2_a221oi_1 _16738_ (.B2(net301),
    .C1(_07726_),
    .B1(_07724_),
    .A1(net954),
    .Y(_07727_),
    .A2(_07716_));
 sg13g2_xnor2_1 _16739_ (.Y(_07728_),
    .A(_07667_),
    .B(_07717_));
 sg13g2_xnor2_1 _16740_ (.Y(_07729_),
    .A(_07339_),
    .B(_07728_));
 sg13g2_xnor2_1 _16741_ (.Y(_07730_),
    .A(net1164),
    .B(_07729_));
 sg13g2_xnor2_1 _16742_ (.Y(_07731_),
    .A(_07257_),
    .B(_07730_));
 sg13g2_buf_1 _16743_ (.A(_07715_),
    .X(_07732_));
 sg13g2_nand2_1 _16744_ (.Y(_07733_),
    .A(net616),
    .B(net928));
 sg13g2_and2_1 _16745_ (.A(net599),
    .B(_07730_),
    .X(_07734_));
 sg13g2_a21oi_1 _16746_ (.A1(_07731_),
    .A2(_07733_),
    .Y(_07735_),
    .B1(_07734_));
 sg13g2_and2_1 _16747_ (.A(_07727_),
    .B(_07735_),
    .X(_07736_));
 sg13g2_nand2_1 _16748_ (.Y(_07737_),
    .A(_07205_),
    .B(net599));
 sg13g2_nor2_1 _16749_ (.A(_07205_),
    .B(_07362_),
    .Y(_07738_));
 sg13g2_nand2_1 _16750_ (.Y(_07739_),
    .A(net616),
    .B(_07362_));
 sg13g2_a21oi_1 _16751_ (.A1(_07730_),
    .A2(_07739_),
    .Y(_07740_),
    .B1(net602));
 sg13g2_a221oi_1 _16752_ (.B2(_07730_),
    .C1(_07740_),
    .B1(_07738_),
    .A1(net612),
    .Y(_07741_),
    .A2(_07737_));
 sg13g2_a22oi_1 _16753_ (.Y(_07742_),
    .B1(_07731_),
    .B2(net612),
    .A2(_07734_),
    .A1(_07732_));
 sg13g2_o21ai_1 _16754_ (.B1(_07742_),
    .Y(_07743_),
    .A1(_07732_),
    .A2(_07741_));
 sg13g2_buf_1 _16755_ (.A(_07718_),
    .X(_07744_));
 sg13g2_nor2_1 _16756_ (.A(_07744_),
    .B(net598),
    .Y(_07745_));
 sg13g2_a21oi_1 _16757_ (.A1(net929),
    .A2(net939),
    .Y(_07746_),
    .B1(net611));
 sg13g2_or2_1 _16758_ (.X(_07747_),
    .B(_07746_),
    .A(_07721_));
 sg13g2_a22oi_1 _16759_ (.Y(_07748_),
    .B1(_07747_),
    .B2(net1162),
    .A2(_07725_),
    .A1(_07745_));
 sg13g2_inv_1 _16760_ (.Y(_07749_),
    .A(_07667_));
 sg13g2_o21ai_1 _16761_ (.B1(net310),
    .Y(_07750_),
    .A1(net951),
    .A2(_07749_));
 sg13g2_nand3_1 _16762_ (.B(_07750_),
    .C(_07745_),
    .A(net1162),
    .Y(_07751_));
 sg13g2_o21ai_1 _16763_ (.B1(_07751_),
    .Y(_07752_),
    .A1(_07673_),
    .A2(_07748_));
 sg13g2_mux2_1 _16764_ (.A0(_07736_),
    .A1(_07743_),
    .S(_07752_),
    .X(_07753_));
 sg13g2_xnor2_1 _16765_ (.Y(_07754_),
    .A(_07611_),
    .B(_07731_));
 sg13g2_a21oi_1 _16766_ (.A1(net116),
    .A2(_07754_),
    .Y(_07755_),
    .B1(net308));
 sg13g2_nor2_1 _16767_ (.A(_07713_),
    .B(_07755_),
    .Y(_07756_));
 sg13g2_o21ai_1 _16768_ (.B1(_07756_),
    .Y(_07757_),
    .A1(net74),
    .A2(_07753_));
 sg13g2_a21oi_1 _16769_ (.A1(_07714_),
    .A2(_07757_),
    .Y(_00335_),
    .B1(net305));
 sg13g2_nand2_1 _16770_ (.Y(_07758_),
    .A(net1056),
    .B(_07713_));
 sg13g2_buf_1 _16771_ (.A(_00224_),
    .X(_07759_));
 sg13g2_nand2_1 _16772_ (.Y(_07760_),
    .A(net1149),
    .B(net1155));
 sg13g2_buf_1 _16773_ (.A(\grid.cell_16_3.se ),
    .X(_07761_));
 sg13g2_xnor2_1 _16774_ (.Y(_07762_),
    .A(net1148),
    .B(_07389_));
 sg13g2_buf_2 _16775_ (.A(_07762_),
    .X(_07763_));
 sg13g2_xor2_1 _16776_ (.B(_06955_),
    .A(net1163),
    .X(_07764_));
 sg13g2_xnor2_1 _16777_ (.Y(_07765_),
    .A(_07763_),
    .B(_07764_));
 sg13g2_xnor2_1 _16778_ (.Y(_07766_),
    .A(net929),
    .B(_07765_));
 sg13g2_buf_1 _16779_ (.A(_07766_),
    .X(_07767_));
 sg13g2_nor2_1 _16780_ (.A(_07302_),
    .B(net1149),
    .Y(_07768_));
 sg13g2_nand2_1 _16781_ (.Y(_07769_),
    .A(net597),
    .B(net1149));
 sg13g2_o21ai_1 _16782_ (.B1(_07769_),
    .Y(_07770_),
    .A1(net613),
    .A2(_07768_));
 sg13g2_nand2_1 _16783_ (.Y(_07771_),
    .A(_07767_),
    .B(_07770_));
 sg13g2_o21ai_1 _16784_ (.B1(_07771_),
    .Y(_07772_),
    .A1(net311),
    .A2(_07760_));
 sg13g2_inv_1 _16785_ (.Y(_07773_),
    .A(net1149));
 sg13g2_a21oi_1 _16786_ (.A1(net600),
    .A2(_07767_),
    .Y(_07774_),
    .B1(_07773_));
 sg13g2_nand2_1 _16787_ (.Y(_07775_),
    .A(_07767_),
    .B(_07768_));
 sg13g2_o21ai_1 _16788_ (.B1(_07775_),
    .Y(_07776_),
    .A1(net951),
    .A2(_07774_));
 sg13g2_nor2_1 _16789_ (.A(net1148),
    .B(net1150),
    .Y(_07777_));
 sg13g2_nor2b_1 _16790_ (.A(net937),
    .B_N(net1163),
    .Y(_07778_));
 sg13g2_nor2b_1 _16791_ (.A(net950),
    .B_N(net1163),
    .Y(_07779_));
 sg13g2_a221oi_1 _16792_ (.B2(_07778_),
    .C1(_07779_),
    .B1(_07777_),
    .A1(net1150),
    .Y(_07780_),
    .A2(net937));
 sg13g2_o21ai_1 _16793_ (.B1(net1148),
    .Y(_07781_),
    .A1(net1150),
    .A2(_07390_));
 sg13g2_and2_1 _16794_ (.A(net1160),
    .B(_07781_),
    .X(_07782_));
 sg13g2_nor3_1 _16795_ (.A(net1148),
    .B(net1150),
    .C(_07390_),
    .Y(_07783_));
 sg13g2_a22oi_1 _16796_ (.Y(_07784_),
    .B1(_07783_),
    .B2(_07030_),
    .A2(_07782_),
    .A1(_07780_));
 sg13g2_buf_1 _16797_ (.A(_07784_),
    .X(_07785_));
 sg13g2_mux2_1 _16798_ (.A0(_07772_),
    .A1(_07776_),
    .S(_07785_),
    .X(_07786_));
 sg13g2_buf_1 _16799_ (.A(net1148),
    .X(_07787_));
 sg13g2_inv_2 _16800_ (.Y(_07788_),
    .A(_07787_));
 sg13g2_buf_1 _16801_ (.A(_07718_),
    .X(_07789_));
 sg13g2_xnor2_1 _16802_ (.Y(_07790_),
    .A(net596),
    .B(net611));
 sg13g2_a21oi_1 _16803_ (.A1(net307),
    .A2(net310),
    .Y(_07791_),
    .B1(_07744_));
 sg13g2_a21oi_1 _16804_ (.A1(net588),
    .A2(_07790_),
    .Y(_07792_),
    .B1(_07791_));
 sg13g2_nand2_1 _16805_ (.Y(_07793_),
    .A(net589),
    .B(net307));
 sg13g2_nor2_1 _16806_ (.A(net1160),
    .B(_07793_),
    .Y(_07794_));
 sg13g2_a21oi_1 _16807_ (.A1(net610),
    .A2(_07792_),
    .Y(_07795_),
    .B1(_07794_));
 sg13g2_nor2_1 _16808_ (.A(_07788_),
    .B(_07795_),
    .Y(_07796_));
 sg13g2_buf_1 _16809_ (.A(net927),
    .X(_07797_));
 sg13g2_buf_1 _16810_ (.A(net587),
    .X(_07798_));
 sg13g2_nor3_1 _16811_ (.A(_07798_),
    .B(_07030_),
    .C(_07793_),
    .Y(_07799_));
 sg13g2_nor3_1 _16812_ (.A(_07336_),
    .B(net1149),
    .C(net1155),
    .Y(_07800_));
 sg13g2_nor3_1 _16813_ (.A(_07381_),
    .B(_07406_),
    .C(_07785_),
    .Y(_07801_));
 sg13g2_o21ai_1 _16814_ (.B1(net951),
    .Y(_07802_),
    .A1(_07800_),
    .A2(_07801_));
 sg13g2_o21ai_1 _16815_ (.B1(_07400_),
    .Y(_07803_),
    .A1(net600),
    .A2(_07759_));
 sg13g2_nor3_1 _16816_ (.A(net597),
    .B(_07759_),
    .C(net1155),
    .Y(_07804_));
 sg13g2_a21o_1 _16817_ (.A2(_07785_),
    .A1(net597),
    .B1(_07804_),
    .X(_07805_));
 sg13g2_nor3_1 _16818_ (.A(net597),
    .B(_07785_),
    .C(_07760_),
    .Y(_07806_));
 sg13g2_a221oi_1 _16819_ (.B2(net311),
    .C1(_07806_),
    .B1(_07805_),
    .A1(_07785_),
    .Y(_07807_),
    .A2(_07803_));
 sg13g2_a21oi_1 _16820_ (.A1(_07802_),
    .A2(_07807_),
    .Y(_07808_),
    .B1(_07767_));
 sg13g2_nor4_1 _16821_ (.A(_07786_),
    .B(_07796_),
    .C(_07799_),
    .D(_07808_),
    .Y(_07809_));
 sg13g2_nand2_1 _16822_ (.Y(_07810_),
    .A(_13074_),
    .B(_07605_));
 sg13g2_xnor2_1 _16823_ (.Y(_07811_),
    .A(_07691_),
    .B(_07767_));
 sg13g2_a21oi_1 _16824_ (.A1(net114),
    .A2(_07811_),
    .Y(_07812_),
    .B1(net601));
 sg13g2_nor2_1 _16825_ (.A(_07810_),
    .B(_07812_),
    .Y(_07813_));
 sg13g2_o21ai_1 _16826_ (.B1(_07813_),
    .Y(_07814_),
    .A1(net81),
    .A2(_07809_));
 sg13g2_o21ai_1 _16827_ (.B1(_07814_),
    .Y(_00336_),
    .A1(net32),
    .A2(_07758_));
 sg13g2_buf_1 _16828_ (.A(\grid.cell_16_4.se ),
    .X(_07815_));
 sg13g2_xnor2_1 _16829_ (.Y(_07816_),
    .A(net1147),
    .B(_07429_));
 sg13g2_xor2_1 _16830_ (.B(_07816_),
    .A(_07054_),
    .X(_07817_));
 sg13g2_xnor2_1 _16831_ (.Y(_07818_),
    .A(net927),
    .B(_07817_));
 sg13g2_xnor2_1 _16832_ (.Y(_07819_),
    .A(net598),
    .B(_07818_));
 sg13g2_nor2_1 _16833_ (.A(_07428_),
    .B(_07818_),
    .Y(_07820_));
 sg13g2_a21oi_1 _16834_ (.A1(net310),
    .A2(_07819_),
    .Y(_07821_),
    .B1(_07820_));
 sg13g2_nor4_1 _16835_ (.A(net1147),
    .B(net1148),
    .C(net936),
    .D(net609),
    .Y(_07822_));
 sg13g2_a221oi_1 _16836_ (.B2(_06999_),
    .C1(_07822_),
    .B1(net1161),
    .A1(net927),
    .Y(_07823_),
    .A2(net595));
 sg13g2_buf_1 _16837_ (.A(net1147),
    .X(_07824_));
 sg13g2_o21ai_1 _16838_ (.B1(_07824_),
    .Y(_07825_),
    .A1(net927),
    .A2(_07430_));
 sg13g2_and2_1 _16839_ (.A(_07082_),
    .B(_07825_),
    .X(_07826_));
 sg13g2_nor3_1 _16840_ (.A(_07824_),
    .B(net927),
    .C(_07447_),
    .Y(_07827_));
 sg13g2_a22oi_1 _16841_ (.Y(_07828_),
    .B1(_07827_),
    .B2(_07046_),
    .A2(_07826_),
    .A1(_07823_));
 sg13g2_buf_1 _16842_ (.A(_00048_),
    .X(_07829_));
 sg13g2_xnor2_1 _16843_ (.Y(_07830_),
    .A(_07761_),
    .B(net1156));
 sg13g2_xnor2_1 _16844_ (.Y(_07831_),
    .A(net950),
    .B(_07830_));
 sg13g2_xnor2_1 _16845_ (.Y(_07832_),
    .A(_07817_),
    .B(_07831_));
 sg13g2_nor2_1 _16846_ (.A(net1146),
    .B(_07832_),
    .Y(_07833_));
 sg13g2_or2_1 _16847_ (.X(_07834_),
    .B(_07833_),
    .A(_07828_));
 sg13g2_buf_1 _16848_ (.A(net926),
    .X(_07835_));
 sg13g2_buf_1 _16849_ (.A(_07835_),
    .X(_07836_));
 sg13g2_nand2_1 _16850_ (.Y(_07837_),
    .A(net587),
    .B(net595));
 sg13g2_xnor2_1 _16851_ (.Y(_07838_),
    .A(_07430_),
    .B(net1163));
 sg13g2_a21oi_1 _16852_ (.A1(_07447_),
    .A2(net947),
    .Y(_07839_),
    .B1(_07787_));
 sg13g2_a21oi_1 _16853_ (.A1(net927),
    .A2(_07838_),
    .Y(_07840_),
    .B1(_07839_));
 sg13g2_nand2_1 _16854_ (.Y(_07841_),
    .A(net608),
    .B(_07840_));
 sg13g2_o21ai_1 _16855_ (.B1(_07841_),
    .Y(_07842_),
    .A1(_07082_),
    .A2(_07837_));
 sg13g2_nor3_1 _16856_ (.A(net299),
    .B(_07046_),
    .C(_07837_),
    .Y(_07843_));
 sg13g2_a221oi_1 _16857_ (.B2(_07833_),
    .C1(_07843_),
    .B1(_07828_),
    .A1(net299),
    .Y(_07844_),
    .A2(_07842_));
 sg13g2_and3_1 _16858_ (.X(_07845_),
    .A(_07821_),
    .B(_07834_),
    .C(_07844_));
 sg13g2_nor3_1 _16859_ (.A(_07828_),
    .B(_07833_),
    .C(_07821_),
    .Y(_07846_));
 sg13g2_nor3_1 _16860_ (.A(net107),
    .B(_07845_),
    .C(_07846_),
    .Y(_07847_));
 sg13g2_xnor2_1 _16861_ (.Y(_07848_),
    .A(net588),
    .B(_07339_));
 sg13g2_xnor2_1 _16862_ (.Y(_07849_),
    .A(_07818_),
    .B(_07848_));
 sg13g2_a21oi_1 _16863_ (.A1(_04650_),
    .A2(_07849_),
    .Y(_07850_),
    .B1(_07396_));
 sg13g2_nor3_1 _16864_ (.A(_07810_),
    .B(_07847_),
    .C(_07850_),
    .Y(_07851_));
 sg13g2_nor2_1 _16865_ (.A(net47),
    .B(_07758_),
    .Y(_07852_));
 sg13g2_or2_1 _16866_ (.X(_00337_),
    .B(_07852_),
    .A(_07851_));
 sg13g2_buf_2 _16867_ (.A(_00080_),
    .X(_07853_));
 sg13g2_xor2_1 _16868_ (.B(net1159),
    .A(_07482_),
    .X(_07854_));
 sg13g2_buf_1 _16869_ (.A(\grid.cell_16_5.se ),
    .X(_07855_));
 sg13g2_buf_1 _16870_ (.A(_07855_),
    .X(_07856_));
 sg13g2_xnor2_1 _16871_ (.Y(_07857_),
    .A(net925),
    .B(net1147));
 sg13g2_xnor2_1 _16872_ (.Y(_07858_),
    .A(_07854_),
    .B(_07857_));
 sg13g2_xor2_1 _16873_ (.B(_07858_),
    .A(_07054_),
    .X(_07859_));
 sg13g2_xnor2_1 _16874_ (.Y(_07860_),
    .A(_07462_),
    .B(_07859_));
 sg13g2_nor2_1 _16875_ (.A(_07853_),
    .B(_07860_),
    .Y(_07861_));
 sg13g2_nor2_1 _16876_ (.A(net594),
    .B(_06999_),
    .Y(_07862_));
 sg13g2_nand2b_1 _16877_ (.Y(_07863_),
    .B(net1154),
    .A_N(_07778_));
 sg13g2_xnor2_1 _16878_ (.Y(_07864_),
    .A(net609),
    .B(_07858_));
 sg13g2_mux2_1 _16879_ (.A0(_07862_),
    .A1(_07863_),
    .S(_07864_),
    .X(_07865_));
 sg13g2_inv_1 _16880_ (.Y(_07866_),
    .A(net925));
 sg13g2_buf_1 _16881_ (.A(_07866_),
    .X(_07867_));
 sg13g2_nor3_1 _16882_ (.A(net926),
    .B(_07484_),
    .C(_07103_),
    .Y(_07868_));
 sg13g2_buf_1 _16883_ (.A(net925),
    .X(_07869_));
 sg13g2_nor3_1 _16884_ (.A(net585),
    .B(net926),
    .C(_07511_),
    .Y(_07870_));
 sg13g2_inv_2 _16885_ (.Y(_07871_),
    .A(net1147));
 sg13g2_nor2_1 _16886_ (.A(_07871_),
    .B(_07486_),
    .Y(_07872_));
 sg13g2_nor2_1 _16887_ (.A(_07102_),
    .B(net1161),
    .Y(_07873_));
 sg13g2_nand2_1 _16888_ (.Y(_07874_),
    .A(net925),
    .B(net935));
 sg13g2_nand2_1 _16889_ (.Y(_07875_),
    .A(_07856_),
    .B(_07815_));
 sg13g2_nand3_1 _16890_ (.B(_07874_),
    .C(_07875_),
    .A(_07137_),
    .Y(_07876_));
 sg13g2_nor4_1 _16891_ (.A(_07870_),
    .B(_07872_),
    .C(_07873_),
    .D(_07876_),
    .Y(_07877_));
 sg13g2_a21oi_1 _16892_ (.A1(net298),
    .A2(_07868_),
    .Y(_07878_),
    .B1(_07877_));
 sg13g2_xnor2_1 _16893_ (.Y(_07879_),
    .A(_07865_),
    .B(_07878_));
 sg13g2_or4_1 _16894_ (.A(_07853_),
    .B(_07865_),
    .C(_07878_),
    .D(_07860_),
    .X(_07880_));
 sg13g2_o21ai_1 _16895_ (.B1(_07880_),
    .Y(_07881_),
    .A1(_07861_),
    .A2(_07879_));
 sg13g2_xnor2_1 _16896_ (.Y(_07882_),
    .A(net593),
    .B(net946));
 sg13g2_a21oi_1 _16897_ (.A1(net304),
    .A2(net946),
    .Y(_07883_),
    .B1(net586));
 sg13g2_a21oi_1 _16898_ (.A1(_07836_),
    .A2(_07882_),
    .Y(_07884_),
    .B1(_07883_));
 sg13g2_a221oi_1 _16899_ (.B2(net607),
    .C1(_07867_),
    .B1(_07884_),
    .A1(_07138_),
    .Y(_07885_),
    .A2(_07872_));
 sg13g2_buf_1 _16900_ (.A(net585),
    .X(_07886_));
 sg13g2_buf_1 _16901_ (.A(net297),
    .X(_07887_));
 sg13g2_a21oi_1 _16902_ (.A1(_07103_),
    .A2(_07872_),
    .Y(_07888_),
    .B1(_07887_));
 sg13g2_or2_1 _16903_ (.X(_07889_),
    .B(_07888_),
    .A(_07885_));
 sg13g2_a21oi_1 _16904_ (.A1(_07881_),
    .A2(_07889_),
    .Y(_07890_),
    .B1(net101));
 sg13g2_xor2_1 _16905_ (.B(_07859_),
    .A(_07763_),
    .X(_07891_));
 sg13g2_a21oi_1 _16906_ (.A1(net77),
    .A2(_07891_),
    .Y(_07892_),
    .B1(net152));
 sg13g2_or3_1 _16907_ (.A(_07810_),
    .B(_07890_),
    .C(_07892_),
    .X(_07893_));
 sg13g2_o21ai_1 _16908_ (.B1(_07893_),
    .Y(_00338_),
    .A1(_05003_),
    .A2(_07758_));
 sg13g2_buf_1 _16909_ (.A(_00142_),
    .X(_07894_));
 sg13g2_and2_1 _16910_ (.A(net934),
    .B(net942),
    .X(_07895_));
 sg13g2_buf_1 _16911_ (.A(_07895_),
    .X(_07896_));
 sg13g2_o21ai_1 _16912_ (.B1(_07645_),
    .Y(_07897_),
    .A1(net297),
    .A2(_07896_));
 sg13g2_nor2_1 _16913_ (.A(net585),
    .B(_07645_),
    .Y(_07898_));
 sg13g2_a21oi_1 _16914_ (.A1(net1145),
    .A2(_07897_),
    .Y(_07899_),
    .B1(_07898_));
 sg13g2_nor2_1 _16915_ (.A(_07189_),
    .B(_07896_),
    .Y(_07900_));
 sg13g2_o21ai_1 _16916_ (.B1(_07900_),
    .Y(_07901_),
    .A1(net1145),
    .A2(_07645_));
 sg13g2_o21ai_1 _16917_ (.B1(_07901_),
    .Y(_07902_),
    .A1(net1145),
    .A2(_07621_));
 sg13g2_nand2_1 _16918_ (.Y(_07903_),
    .A(net302),
    .B(_07214_));
 sg13g2_and2_1 _16919_ (.A(_07609_),
    .B(net955),
    .X(_07904_));
 sg13g2_nor2b_1 _16920_ (.A(_07869_),
    .B_N(net1145),
    .Y(_07905_));
 sg13g2_o21ai_1 _16921_ (.B1(_07905_),
    .Y(_07906_),
    .A1(_07622_),
    .A2(_07904_));
 sg13g2_o21ai_1 _16922_ (.B1(_07906_),
    .Y(_07907_),
    .A1(net1145),
    .A2(_07903_));
 sg13g2_nor2_1 _16923_ (.A(_07866_),
    .B(_07623_),
    .Y(_07908_));
 sg13g2_a21oi_1 _16924_ (.A1(_07214_),
    .A2(_07908_),
    .Y(_07909_),
    .B1(_07898_));
 sg13g2_nor2_1 _16925_ (.A(net607),
    .B(_07909_),
    .Y(_07910_));
 sg13g2_a221oi_1 _16926_ (.B2(net607),
    .C1(_07910_),
    .B1(_07907_),
    .A1(net149),
    .Y(_07911_),
    .A2(_07902_));
 sg13g2_o21ai_1 _16927_ (.B1(_07911_),
    .Y(_07912_),
    .A1(net154),
    .A2(_07899_));
 sg13g2_buf_1 _16928_ (.A(_00112_),
    .X(_07913_));
 sg13g2_inv_1 _16929_ (.Y(_07914_),
    .A(net1144));
 sg13g2_xnor2_1 _16930_ (.Y(_07915_),
    .A(net925),
    .B(_07608_));
 sg13g2_xnor2_1 _16931_ (.Y(_07916_),
    .A(_07216_),
    .B(_07915_));
 sg13g2_xnor2_1 _16932_ (.Y(_07917_),
    .A(net1159),
    .B(_07916_));
 sg13g2_xnor2_1 _16933_ (.Y(_07918_),
    .A(net152),
    .B(_07917_));
 sg13g2_a21oi_1 _16934_ (.A1(net1144),
    .A2(net609),
    .Y(_07919_),
    .B1(_07918_));
 sg13g2_a221oi_1 _16935_ (.B2(_07539_),
    .C1(_07919_),
    .B1(_07917_),
    .A1(_07914_),
    .Y(_07920_),
    .A2(net608));
 sg13g2_xor2_1 _16936_ (.B(_07920_),
    .A(_07912_),
    .X(_07921_));
 sg13g2_xnor2_1 _16937_ (.Y(_07922_),
    .A(net309),
    .B(net945));
 sg13g2_o21ai_1 _16938_ (.B1(net154),
    .Y(_07923_),
    .A1(net150),
    .A2(_07569_));
 sg13g2_a21o_1 _16939_ (.A2(_07922_),
    .A1(_07641_),
    .B1(_07923_),
    .X(_07924_));
 sg13g2_o21ai_1 _16940_ (.B1(_07924_),
    .Y(_07925_),
    .A1(_07894_),
    .A2(_07621_));
 sg13g2_nor2_1 _16941_ (.A(net149),
    .B(_07189_),
    .Y(_07926_));
 sg13g2_a221oi_1 _16942_ (.B2(_07896_),
    .C1(net99),
    .B1(_07926_),
    .A1(net149),
    .Y(_07927_),
    .A2(_07925_));
 sg13g2_nand4_1 _16943_ (.B(_07914_),
    .C(_07556_),
    .A(_07539_),
    .Y(_07928_),
    .D(_07917_));
 sg13g2_xnor2_1 _16944_ (.Y(_07929_),
    .A(net608),
    .B(_07816_));
 sg13g2_xnor2_1 _16945_ (.Y(_07930_),
    .A(_07917_),
    .B(_07929_));
 sg13g2_nand2_1 _16946_ (.Y(_07931_),
    .A(_07486_),
    .B(_07930_));
 sg13g2_nand4_1 _16947_ (.B(_07927_),
    .C(_07928_),
    .A(_07921_),
    .Y(_07932_),
    .D(_07931_));
 sg13g2_a22oi_1 _16948_ (.Y(_07933_),
    .B1(net25),
    .B2(_07603_),
    .A2(net71),
    .A1(net151));
 sg13g2_a221oi_1 _16949_ (.B2(_07933_),
    .C1(_06815_),
    .B1(_07932_),
    .A1(net24),
    .Y(_00339_),
    .A2(_07603_));
 sg13g2_nand2_1 _16950_ (.Y(_07934_),
    .A(net304),
    .B(net945));
 sg13g2_nand2_1 _16951_ (.Y(_07935_),
    .A(_07640_),
    .B(_07854_));
 sg13g2_o21ai_1 _16952_ (.B1(_07935_),
    .Y(_07936_),
    .A1(_07641_),
    .A2(_07934_));
 sg13g2_and2_1 _16953_ (.A(_07608_),
    .B(_07482_),
    .X(_07937_));
 sg13g2_buf_1 _16954_ (.A(_07937_),
    .X(_07938_));
 sg13g2_nor2b_1 _16955_ (.A(net1145),
    .B_N(_07938_),
    .Y(_07939_));
 sg13g2_a21oi_1 _16956_ (.A1(net154),
    .A2(_07936_),
    .Y(_07940_),
    .B1(_07939_));
 sg13g2_xor2_1 _16957_ (.B(_07915_),
    .A(_07854_),
    .X(_07941_));
 sg13g2_xnor2_1 _16958_ (.Y(_07942_),
    .A(net614),
    .B(_07941_));
 sg13g2_a221oi_1 _16959_ (.B2(_07705_),
    .C1(_03810_),
    .B1(_07942_),
    .A1(_07926_),
    .Y(_07943_),
    .A2(_07938_));
 sg13g2_o21ai_1 _16960_ (.B1(_07943_),
    .Y(_07944_),
    .A1(net298),
    .A2(_07940_));
 sg13g2_nor2_1 _16961_ (.A(_07620_),
    .B(net935),
    .Y(_07945_));
 sg13g2_nand2_1 _16962_ (.Y(_07946_),
    .A(_07867_),
    .B(_07945_));
 sg13g2_nor2_1 _16963_ (.A(_07869_),
    .B(_07938_),
    .Y(_07947_));
 sg13g2_o21ai_1 _16964_ (.B1(net1145),
    .Y(_07948_),
    .A1(_07945_),
    .A2(_07947_));
 sg13g2_a21oi_1 _16965_ (.A1(_07946_),
    .A2(_07948_),
    .Y(_07949_),
    .B1(net154));
 sg13g2_nor3_1 _16966_ (.A(_00142_),
    .B(_07609_),
    .C(_07483_),
    .Y(_07950_));
 sg13g2_nor3_1 _16967_ (.A(_07189_),
    .B(_07938_),
    .C(_07950_),
    .Y(_07951_));
 sg13g2_o21ai_1 _16968_ (.B1(_07886_),
    .Y(_07952_),
    .A1(_07939_),
    .A2(_07951_));
 sg13g2_inv_1 _16969_ (.Y(_07953_),
    .A(_07952_));
 sg13g2_a21o_1 _16970_ (.A2(net593),
    .A1(_07623_),
    .B1(_07904_),
    .X(_07954_));
 sg13g2_nor2b_1 _16971_ (.A(net1145),
    .B_N(net615),
    .Y(_07955_));
 sg13g2_a22oi_1 _16972_ (.Y(_07956_),
    .B1(_07955_),
    .B2(_07938_),
    .A2(_07954_),
    .A1(_07905_));
 sg13g2_nor2_1 _16973_ (.A(net606),
    .B(_07956_),
    .Y(_07957_));
 sg13g2_nand3_1 _16974_ (.B(net313),
    .C(_07908_),
    .A(net593),
    .Y(_07958_));
 sg13g2_a21oi_1 _16975_ (.A1(_07946_),
    .A2(_07958_),
    .Y(_07959_),
    .B1(net945));
 sg13g2_nor4_1 _16976_ (.A(_07949_),
    .B(_07953_),
    .C(_07957_),
    .D(_07959_),
    .Y(_07960_));
 sg13g2_xor2_1 _16977_ (.B(_07942_),
    .A(_07268_),
    .X(_07961_));
 sg13g2_nor2b_1 _16978_ (.A(_07637_),
    .B_N(net953),
    .Y(_07962_));
 sg13g2_a221oi_1 _16979_ (.B2(_07662_),
    .C1(_07962_),
    .B1(_07961_),
    .A1(_07234_),
    .Y(_07963_),
    .A2(_07942_));
 sg13g2_xor2_1 _16980_ (.B(_07963_),
    .A(_07960_),
    .X(_07964_));
 sg13g2_nor2_1 _16981_ (.A(_07944_),
    .B(_07964_),
    .Y(_07965_));
 sg13g2_nor2_1 _16982_ (.A(net603),
    .B(_07713_),
    .Y(_07966_));
 sg13g2_o21ai_1 _16983_ (.B1(_07966_),
    .Y(_07967_),
    .A1(net73),
    .A2(_07965_));
 sg13g2_xnor2_1 _16984_ (.Y(_07968_),
    .A(_07703_),
    .B(_07942_));
 sg13g2_nor2_1 _16985_ (.A(_07713_),
    .B(_07968_),
    .Y(_07969_));
 sg13g2_a22oi_1 _16986_ (.Y(_07970_),
    .B1(_07965_),
    .B2(_07969_),
    .A2(_07713_),
    .A1(_05678_));
 sg13g2_a21oi_1 _16987_ (.A1(_07967_),
    .A2(_07970_),
    .Y(_00340_),
    .B1(_07480_));
 sg13g2_a21oi_1 _16988_ (.A1(net1188),
    .A2(_01492_),
    .Y(_07971_),
    .B1(_05745_));
 sg13g2_buf_2 _16989_ (.A(_07971_),
    .X(_07972_));
 sg13g2_nor3_1 _16990_ (.A(_07972_),
    .B(net320),
    .C(_07602_),
    .Y(_07973_));
 sg13g2_buf_2 _16991_ (.A(_07973_),
    .X(_07974_));
 sg13g2_and2_1 _16992_ (.A(net158),
    .B(_07974_),
    .X(_07975_));
 sg13g2_buf_1 _16993_ (.A(_07975_),
    .X(_07976_));
 sg13g2_nand2_2 _16994_ (.Y(_07977_),
    .A(_12977_),
    .B(_07976_));
 sg13g2_buf_2 _16995_ (.A(\grid.cell_17_0.sw ),
    .X(_07978_));
 sg13g2_xnor2_1 _16996_ (.Y(_07979_),
    .A(_07978_),
    .B(_07608_));
 sg13g2_buf_2 _16997_ (.A(_07979_),
    .X(_07980_));
 sg13g2_buf_1 _16998_ (.A(\grid.cell_17_0.se ),
    .X(_07981_));
 sg13g2_xnor2_1 _16999_ (.Y(_07982_),
    .A(_07203_),
    .B(net1143));
 sg13g2_xnor2_1 _17000_ (.Y(_07983_),
    .A(_07207_),
    .B(_07982_));
 sg13g2_xnor2_1 _17001_ (.Y(_07984_),
    .A(_07980_),
    .B(_07983_));
 sg13g2_xor2_1 _17002_ (.B(_07983_),
    .A(_07980_),
    .X(_07985_));
 sg13g2_xnor2_1 _17003_ (.Y(_07986_),
    .A(net931),
    .B(_07985_));
 sg13g2_buf_1 _17004_ (.A(net1143),
    .X(_07987_));
 sg13g2_buf_1 _17005_ (.A(_07987_),
    .X(_07988_));
 sg13g2_buf_1 _17006_ (.A(_07978_),
    .X(_07989_));
 sg13g2_buf_1 _17007_ (.A(net923),
    .X(_07990_));
 sg13g2_buf_1 _17008_ (.A(net583),
    .X(_07991_));
 sg13g2_nand2b_1 _17009_ (.Y(_07992_),
    .B(net592),
    .A_N(_07346_));
 sg13g2_buf_1 _17010_ (.A(net583),
    .X(_07993_));
 sg13g2_nor2_1 _17011_ (.A(net295),
    .B(_07623_),
    .Y(_07994_));
 sg13g2_a21oi_1 _17012_ (.A1(net296),
    .A2(_07992_),
    .Y(_07995_),
    .B1(_07994_));
 sg13g2_nor2_1 _17013_ (.A(net296),
    .B(net302),
    .Y(_07996_));
 sg13g2_nand2b_1 _17014_ (.Y(_07997_),
    .B(net295),
    .A_N(net592));
 sg13g2_o21ai_1 _17015_ (.B1(_07997_),
    .Y(_07998_),
    .A1(net296),
    .A2(net603));
 sg13g2_a22oi_1 _17016_ (.Y(_07999_),
    .B1(_07998_),
    .B2(net602),
    .A2(_07996_),
    .A1(net599));
 sg13g2_o21ai_1 _17017_ (.B1(_07999_),
    .Y(_08000_),
    .A1(net153),
    .A2(_07995_));
 sg13g2_or2_1 _17018_ (.X(_08001_),
    .B(net934),
    .A(net923));
 sg13g2_buf_1 _17019_ (.A(_08001_),
    .X(_08002_));
 sg13g2_nor2_1 _17020_ (.A(_07203_),
    .B(net603),
    .Y(_08003_));
 sg13g2_nand2b_1 _17021_ (.Y(_08004_),
    .B(net592),
    .A_N(net942));
 sg13g2_o21ai_1 _17022_ (.B1(_08004_),
    .Y(_08005_),
    .A1(net592),
    .A2(net938));
 sg13g2_nor2_1 _17023_ (.A(net296),
    .B(_07992_),
    .Y(_08006_));
 sg13g2_a221oi_1 _17024_ (.B2(_07991_),
    .C1(_08006_),
    .B1(_08005_),
    .A1(_08002_),
    .Y(_08007_),
    .A2(_08003_));
 sg13g2_nor4_1 _17025_ (.A(net1143),
    .B(net296),
    .C(net302),
    .D(net603),
    .Y(_08008_));
 sg13g2_inv_2 _17026_ (.Y(_08009_),
    .A(net1143));
 sg13g2_nand2_1 _17027_ (.Y(_08010_),
    .A(net583),
    .B(net934));
 sg13g2_nor3_1 _17028_ (.A(_08009_),
    .B(net599),
    .C(_08010_),
    .Y(_08011_));
 sg13g2_o21ai_1 _17029_ (.B1(net943),
    .Y(_08012_),
    .A1(_08008_),
    .A2(_08011_));
 sg13g2_o21ai_1 _17030_ (.B1(_08012_),
    .Y(_08013_),
    .A1(net584),
    .A2(_08007_));
 sg13g2_a21oi_1 _17031_ (.A1(net584),
    .A2(_08000_),
    .Y(_08014_),
    .B1(_08013_));
 sg13g2_a221oi_1 _17032_ (.B2(net941),
    .C1(_08014_),
    .B1(_07986_),
    .A1(_07716_),
    .Y(_08015_),
    .A2(_07984_));
 sg13g2_nand2_1 _17033_ (.Y(_08016_),
    .A(net605),
    .B(net153));
 sg13g2_and2_1 _17034_ (.A(_07989_),
    .B(_07608_),
    .X(_08017_));
 sg13g2_buf_1 _17035_ (.A(_08017_),
    .X(_08018_));
 sg13g2_nand2b_1 _17036_ (.Y(_08019_),
    .B(net943),
    .A_N(_07980_));
 sg13g2_o21ai_1 _17037_ (.B1(_08019_),
    .Y(_08020_),
    .A1(net153),
    .A2(_08018_));
 sg13g2_a22oi_1 _17038_ (.Y(_08021_),
    .B1(_08020_),
    .B2(net938),
    .A2(_07996_),
    .A1(_08016_));
 sg13g2_o21ai_1 _17039_ (.B1(net153),
    .Y(_08022_),
    .A1(net602),
    .A2(_08009_));
 sg13g2_nand3_1 _17040_ (.B(_08022_),
    .C(_07996_),
    .A(net938),
    .Y(_08023_));
 sg13g2_o21ai_1 _17041_ (.B1(_08023_),
    .Y(_08024_),
    .A1(net584),
    .A2(_08021_));
 sg13g2_buf_1 _17042_ (.A(_00223_),
    .X(_08025_));
 sg13g2_nand2_1 _17043_ (.Y(_08026_),
    .A(net932),
    .B(_07716_));
 sg13g2_o21ai_1 _17044_ (.B1(_07984_),
    .Y(_08027_),
    .A1(_07268_),
    .A2(net928));
 sg13g2_nor3_1 _17045_ (.A(_07631_),
    .B(_07716_),
    .C(_07985_),
    .Y(_08028_));
 sg13g2_a221oi_1 _17046_ (.B2(_07631_),
    .C1(_08028_),
    .B1(_08027_),
    .A1(net941),
    .Y(_08029_),
    .A2(_08026_));
 sg13g2_nor2_1 _17047_ (.A(net928),
    .B(_07985_),
    .Y(_08030_));
 sg13g2_a22oi_1 _17048_ (.Y(_08031_),
    .B1(_08030_),
    .B2(net1142),
    .A2(_07986_),
    .A1(net941));
 sg13g2_o21ai_1 _17049_ (.B1(_08031_),
    .Y(_08032_),
    .A1(net1142),
    .A2(_08029_));
 sg13g2_mux2_1 _17050_ (.A0(_08015_),
    .A1(_08024_),
    .S(_08032_),
    .X(_08033_));
 sg13g2_buf_1 _17051_ (.A(\grid.cell_17_0.s ),
    .X(_08034_));
 sg13g2_buf_1 _17052_ (.A(_08034_),
    .X(_08035_));
 sg13g2_buf_1 _17053_ (.A(net922),
    .X(_08036_));
 sg13g2_xnor2_1 _17054_ (.Y(_08037_),
    .A(net941),
    .B(_08036_));
 sg13g2_xnor2_1 _17055_ (.Y(_08038_),
    .A(_07986_),
    .B(_08037_));
 sg13g2_a21oi_1 _17056_ (.A1(_02820_),
    .A2(_08038_),
    .Y(_08039_),
    .B1(net933));
 sg13g2_nand2_1 _17057_ (.Y(_08040_),
    .A(net158),
    .B(_07974_));
 sg13g2_nand2_1 _17058_ (.Y(_08041_),
    .A(net1059),
    .B(_08040_));
 sg13g2_nor2_1 _17059_ (.A(_08039_),
    .B(_08041_),
    .Y(_08042_));
 sg13g2_o21ai_1 _17060_ (.B1(_08042_),
    .Y(_08043_),
    .A1(net81),
    .A2(_08033_));
 sg13g2_o21ai_1 _17061_ (.B1(_08043_),
    .Y(_00341_),
    .A1(_01817_),
    .A2(_07977_));
 sg13g2_buf_2 _17062_ (.A(\grid.cell_17_1.se ),
    .X(_08044_));
 sg13g2_buf_1 _17063_ (.A(_08044_),
    .X(_08045_));
 sg13g2_nand2_1 _17064_ (.Y(_08046_),
    .A(net924),
    .B(net921));
 sg13g2_buf_1 _17065_ (.A(net921),
    .X(_08047_));
 sg13g2_nor2_1 _17066_ (.A(net930),
    .B(net581),
    .Y(_08048_));
 sg13g2_nand2_1 _17067_ (.Y(_08049_),
    .A(_08009_),
    .B(_08048_));
 sg13g2_o21ai_1 _17068_ (.B1(_08049_),
    .Y(_08050_),
    .A1(_07697_),
    .A2(_08046_));
 sg13g2_inv_1 _17069_ (.Y(_08051_),
    .A(_08044_));
 sg13g2_buf_1 _17070_ (.A(_08051_),
    .X(_08052_));
 sg13g2_nor2_1 _17071_ (.A(net580),
    .B(net938),
    .Y(_08053_));
 sg13g2_nor2_1 _17072_ (.A(net581),
    .B(_07320_),
    .Y(_08054_));
 sg13g2_o21ai_1 _17073_ (.B1(net301),
    .Y(_08055_),
    .A1(_08053_),
    .A2(_08054_));
 sg13g2_nor2_1 _17074_ (.A(net590),
    .B(_07320_),
    .Y(_08056_));
 sg13g2_o21ai_1 _17075_ (.B1(_08056_),
    .Y(_08057_),
    .A1(net581),
    .A2(net938));
 sg13g2_nand3_1 _17076_ (.B(_08055_),
    .C(_08057_),
    .A(net584),
    .Y(_08058_));
 sg13g2_nand2_1 _17077_ (.Y(_08059_),
    .A(net580),
    .B(net938));
 sg13g2_o21ai_1 _17078_ (.B1(_08059_),
    .Y(_08060_),
    .A1(_07668_),
    .A2(_08053_));
 sg13g2_nand2_1 _17079_ (.Y(_08061_),
    .A(net581),
    .B(net938));
 sg13g2_o21ai_1 _17080_ (.B1(_07668_),
    .Y(_08062_),
    .A1(net921),
    .A2(net938));
 sg13g2_a21oi_1 _17081_ (.A1(_08061_),
    .A2(_08062_),
    .Y(_08063_),
    .B1(_07320_));
 sg13g2_a21oi_1 _17082_ (.A1(net597),
    .A2(_08060_),
    .Y(_08064_),
    .B1(_08063_));
 sg13g2_nand2_1 _17083_ (.Y(_08065_),
    .A(_08009_),
    .B(_08064_));
 sg13g2_buf_1 _17084_ (.A(_08047_),
    .X(_08066_));
 sg13g2_nor4_1 _17085_ (.A(net308),
    .B(net301),
    .C(net294),
    .D(net599),
    .Y(_08067_));
 sg13g2_a221oi_1 _17086_ (.B2(_08065_),
    .C1(_08067_),
    .B1(_08058_),
    .A1(net602),
    .Y(_08068_),
    .A2(_08050_));
 sg13g2_nand2b_1 _17087_ (.Y(_08069_),
    .B(net1142),
    .A_N(_07269_));
 sg13g2_xnor2_1 _17088_ (.Y(_08070_),
    .A(_07981_),
    .B(net921));
 sg13g2_xor2_1 _17089_ (.B(_08070_),
    .A(_07690_),
    .X(_08071_));
 sg13g2_xnor2_1 _17090_ (.Y(_08072_),
    .A(_07257_),
    .B(_08071_));
 sg13g2_xnor2_1 _17091_ (.Y(_08073_),
    .A(net933),
    .B(_08072_));
 sg13g2_nand2b_1 _17092_ (.Y(_08074_),
    .B(_07268_),
    .A_N(net1142));
 sg13g2_o21ai_1 _17093_ (.B1(_08074_),
    .Y(_08075_),
    .A1(_07637_),
    .A2(_08072_));
 sg13g2_a21oi_1 _17094_ (.A1(_08069_),
    .A2(_08073_),
    .Y(_08076_),
    .B1(_08075_));
 sg13g2_xnor2_1 _17095_ (.Y(_08077_),
    .A(_08068_),
    .B(_08076_));
 sg13g2_nand2_1 _17096_ (.Y(_08078_),
    .A(net590),
    .B(_08047_));
 sg13g2_xor2_1 _17097_ (.B(_08044_),
    .A(net1151),
    .X(_08079_));
 sg13g2_nand2_1 _17098_ (.Y(_08080_),
    .A(net943),
    .B(_08079_));
 sg13g2_o21ai_1 _17099_ (.B1(_08080_),
    .Y(_08081_),
    .A1(net605),
    .A2(_08078_));
 sg13g2_a22oi_1 _17100_ (.Y(_08082_),
    .B1(_08081_),
    .B2(net308),
    .A2(_08053_),
    .A1(net301));
 sg13g2_or4_1 _17101_ (.A(net602),
    .B(_07988_),
    .C(_08052_),
    .D(_07697_),
    .X(_08083_));
 sg13g2_o21ai_1 _17102_ (.B1(_08083_),
    .Y(_08084_),
    .A1(_08009_),
    .A2(_08082_));
 sg13g2_xor2_1 _17103_ (.B(_07615_),
    .A(_07268_),
    .X(_08085_));
 sg13g2_or3_1 _17104_ (.A(_08025_),
    .B(_07637_),
    .C(_08085_),
    .X(_08086_));
 sg13g2_o21ai_1 _17105_ (.B1(net119),
    .Y(_08087_),
    .A1(_08072_),
    .A2(_08086_));
 sg13g2_xnor2_1 _17106_ (.Y(_08088_),
    .A(_07614_),
    .B(net922));
 sg13g2_xnor2_1 _17107_ (.Y(_08089_),
    .A(_07268_),
    .B(_08088_));
 sg13g2_xnor2_1 _17108_ (.Y(_08090_),
    .A(_08072_),
    .B(_08089_));
 sg13g2_nor2_1 _17109_ (.A(net591),
    .B(_08090_),
    .Y(_08091_));
 sg13g2_nor3_1 _17110_ (.A(_08084_),
    .B(_08087_),
    .C(_08091_),
    .Y(_08092_));
 sg13g2_a22oi_1 _17111_ (.Y(_08093_),
    .B1(_08077_),
    .B2(_08092_),
    .A2(_06538_),
    .A1(net591));
 sg13g2_o21ai_1 _17112_ (.B1(net334),
    .Y(_08094_),
    .A1(net49),
    .A2(_08040_));
 sg13g2_a21oi_1 _17113_ (.A1(_08040_),
    .A2(_08093_),
    .Y(_00342_),
    .B1(_08094_));
 sg13g2_buf_1 _17114_ (.A(\grid.cell_17_2.se ),
    .X(_08095_));
 sg13g2_buf_1 _17115_ (.A(_08095_),
    .X(_08096_));
 sg13g2_nand2_1 _17116_ (.Y(_08097_),
    .A(_08096_),
    .B(net929));
 sg13g2_inv_1 _17117_ (.Y(_08098_),
    .A(_08097_));
 sg13g2_xor2_1 _17118_ (.B(net1150),
    .A(_08095_),
    .X(_08099_));
 sg13g2_nand2_1 _17119_ (.Y(_08100_),
    .A(net1157),
    .B(_08099_));
 sg13g2_o21ai_1 _17120_ (.B1(_08100_),
    .Y(_08101_),
    .A1(net939),
    .A2(_08098_));
 sg13g2_nand2_1 _17121_ (.Y(_08102_),
    .A(net940),
    .B(net598));
 sg13g2_nor2_1 _17122_ (.A(_08096_),
    .B(net929),
    .Y(_08103_));
 sg13g2_a22oi_1 _17123_ (.Y(_08104_),
    .B1(_08102_),
    .B2(_08103_),
    .A2(_08101_),
    .A1(net1155));
 sg13g2_o21ai_1 _17124_ (.B1(net598),
    .Y(_08105_),
    .A1(net597),
    .A2(_08052_));
 sg13g2_nand3_1 _17125_ (.B(_08105_),
    .C(_08103_),
    .A(net1155),
    .Y(_08106_));
 sg13g2_o21ai_1 _17126_ (.B1(_08106_),
    .Y(_08107_),
    .A1(net294),
    .A2(_08104_));
 sg13g2_buf_2 _17127_ (.A(_00222_),
    .X(_08108_));
 sg13g2_nand2_1 _17128_ (.Y(_08109_),
    .A(net602),
    .B(_08108_));
 sg13g2_xor2_1 _17129_ (.B(_08044_),
    .A(net1157),
    .X(_08110_));
 sg13g2_xnor2_1 _17130_ (.Y(_08111_),
    .A(_07375_),
    .B(_08099_));
 sg13g2_xnor2_1 _17131_ (.Y(_08112_),
    .A(_08110_),
    .B(_08111_));
 sg13g2_xnor2_1 _17132_ (.Y(_08113_),
    .A(net931),
    .B(_08112_));
 sg13g2_inv_2 _17133_ (.Y(_08114_),
    .A(_08108_));
 sg13g2_nand2_1 _17134_ (.Y(_08115_),
    .A(net943),
    .B(_08114_));
 sg13g2_o21ai_1 _17135_ (.B1(_08115_),
    .Y(_08116_),
    .A1(net928),
    .A2(_08112_));
 sg13g2_a21oi_1 _17136_ (.A1(_08109_),
    .A2(_08113_),
    .Y(_08117_),
    .B1(_08116_));
 sg13g2_xor2_1 _17137_ (.B(_08117_),
    .A(_08107_),
    .X(_08118_));
 sg13g2_o21ai_1 _17138_ (.B1(_08100_),
    .Y(_08119_),
    .A1(net940),
    .A2(_08097_));
 sg13g2_nand2_1 _17139_ (.Y(_08120_),
    .A(net601),
    .B(_08119_));
 sg13g2_o21ai_1 _17140_ (.B1(_08120_),
    .Y(_08121_),
    .A1(net1155),
    .A2(_08097_));
 sg13g2_nor3_1 _17141_ (.A(net597),
    .B(net294),
    .C(_07719_),
    .Y(_08122_));
 sg13g2_buf_1 _17142_ (.A(net920),
    .X(_08123_));
 sg13g2_buf_1 _17143_ (.A(_08123_),
    .X(_08124_));
 sg13g2_xor2_1 _17144_ (.B(net932),
    .A(net943),
    .X(_08125_));
 sg13g2_nor4_1 _17145_ (.A(_08108_),
    .B(net928),
    .C(_08125_),
    .D(_08112_),
    .Y(_08126_));
 sg13g2_a221oi_1 _17146_ (.B2(_08124_),
    .C1(_08126_),
    .B1(_08122_),
    .A1(_08066_),
    .Y(_08127_),
    .A2(_08121_));
 sg13g2_a21oi_1 _17147_ (.A1(_08118_),
    .A2(_08127_),
    .Y(_08128_),
    .B1(_06993_));
 sg13g2_xnor2_1 _17148_ (.Y(_08129_),
    .A(_07982_),
    .B(_08113_));
 sg13g2_a21oi_1 _17149_ (.A1(net77),
    .A2(_08129_),
    .Y(_08130_),
    .B1(net301));
 sg13g2_or3_1 _17150_ (.A(_08041_),
    .B(_08128_),
    .C(_08130_),
    .X(_08131_));
 sg13g2_o21ai_1 _17151_ (.B1(_08131_),
    .Y(_00343_),
    .A1(_04088_),
    .A2(_07977_));
 sg13g2_buf_1 _17152_ (.A(\grid.cell_17_3.se ),
    .X(_08132_));
 sg13g2_xnor2_1 _17153_ (.Y(_08133_),
    .A(net1141),
    .B(net920));
 sg13g2_xnor2_1 _17154_ (.Y(_08134_),
    .A(_07830_),
    .B(_08133_));
 sg13g2_xnor2_1 _17155_ (.Y(_08135_),
    .A(net937),
    .B(_08134_));
 sg13g2_nand2_1 _17156_ (.Y(_08136_),
    .A(_07773_),
    .B(_08135_));
 sg13g2_buf_2 _17157_ (.A(_00221_),
    .X(_08137_));
 sg13g2_xnor2_1 _17158_ (.Y(_08138_),
    .A(net1151),
    .B(net1156));
 sg13g2_xnor2_1 _17159_ (.Y(_08139_),
    .A(_08133_),
    .B(_08138_));
 sg13g2_xnor2_1 _17160_ (.Y(_08140_),
    .A(_07763_),
    .B(_08139_));
 sg13g2_buf_1 _17161_ (.A(_08140_),
    .X(_08141_));
 sg13g2_nor2_1 _17162_ (.A(_08137_),
    .B(_08141_),
    .Y(_08142_));
 sg13g2_and2_1 _17163_ (.A(_07773_),
    .B(_08135_),
    .X(_08143_));
 sg13g2_o21ai_1 _17164_ (.B1(_08141_),
    .Y(_08144_),
    .A1(_08137_),
    .A2(_08143_));
 sg13g2_a21oi_1 _17165_ (.A1(net597),
    .A2(_08141_),
    .Y(_08145_),
    .B1(_08137_));
 sg13g2_nor2_1 _17166_ (.A(_08136_),
    .B(_08145_),
    .Y(_08146_));
 sg13g2_a221oi_1 _17167_ (.B2(net308),
    .C1(_08146_),
    .B1(_08144_),
    .A1(_08136_),
    .Y(_08147_),
    .A2(_08142_));
 sg13g2_nand2_1 _17168_ (.Y(_08148_),
    .A(_08137_),
    .B(_08141_));
 sg13g2_o21ai_1 _17169_ (.B1(_08148_),
    .Y(_08149_),
    .A1(net308),
    .A2(_08142_));
 sg13g2_nand2_1 _17170_ (.Y(_08150_),
    .A(_08136_),
    .B(_08149_));
 sg13g2_buf_1 _17171_ (.A(net1141),
    .X(_08151_));
 sg13g2_nor4_1 _17172_ (.A(_08151_),
    .B(net920),
    .C(_07797_),
    .D(net594),
    .Y(_08152_));
 sg13g2_a221oi_1 _17173_ (.B2(_07375_),
    .C1(_08152_),
    .B1(net307),
    .A1(net579),
    .Y(_08153_),
    .A2(net587));
 sg13g2_o21ai_1 _17174_ (.B1(_08151_),
    .Y(_08154_),
    .A1(net579),
    .A2(_07797_));
 sg13g2_and2_1 _17175_ (.A(_07428_),
    .B(_08154_),
    .X(_08155_));
 sg13g2_buf_1 _17176_ (.A(net919),
    .X(_08156_));
 sg13g2_nor3_1 _17177_ (.A(net578),
    .B(_08123_),
    .C(net300),
    .Y(_08157_));
 sg13g2_nand2_1 _17178_ (.Y(_08158_),
    .A(net307),
    .B(net601));
 sg13g2_a22oi_1 _17179_ (.Y(_08159_),
    .B1(_08157_),
    .B2(_08158_),
    .A2(_08155_),
    .A1(_08153_));
 sg13g2_mux2_1 _17180_ (.A0(_08147_),
    .A1(_08150_),
    .S(_08159_),
    .X(_08160_));
 sg13g2_xnor2_1 _17181_ (.Y(_08161_),
    .A(_08110_),
    .B(_08141_));
 sg13g2_a21oi_1 _17182_ (.A1(net111),
    .A2(_08161_),
    .Y(_08162_),
    .B1(_07789_));
 sg13g2_inv_1 _17183_ (.Y(_08163_),
    .A(net1141));
 sg13g2_buf_1 _17184_ (.A(_08163_),
    .X(_08164_));
 sg13g2_inv_1 _17185_ (.Y(_08165_),
    .A(net920));
 sg13g2_nand3_1 _17186_ (.B(net300),
    .C(net601),
    .A(_08165_),
    .Y(_08166_));
 sg13g2_o21ai_1 _17187_ (.B1(_08166_),
    .Y(_08167_),
    .A1(_08165_),
    .A2(_07830_));
 sg13g2_nand2_1 _17188_ (.Y(_08168_),
    .A(_08124_),
    .B(net300));
 sg13g2_nor2_1 _17189_ (.A(_07428_),
    .B(_08168_),
    .Y(_08169_));
 sg13g2_a21oi_1 _17190_ (.A1(net307),
    .A2(_08167_),
    .Y(_08170_),
    .B1(_08169_));
 sg13g2_buf_1 _17191_ (.A(net578),
    .X(_08171_));
 sg13g2_or3_1 _17192_ (.A(_08171_),
    .B(_08158_),
    .C(_08168_),
    .X(_08172_));
 sg13g2_o21ai_1 _17193_ (.B1(_08172_),
    .Y(_08173_),
    .A1(net577),
    .A2(_08170_));
 sg13g2_nor4_1 _17194_ (.A(_08041_),
    .B(_08160_),
    .C(_08162_),
    .D(_08173_),
    .Y(_08174_));
 sg13g2_nand4_1 _17195_ (.B(_07789_),
    .C(net115),
    .A(net1056),
    .Y(_08175_),
    .D(_08040_));
 sg13g2_o21ai_1 _17196_ (.B1(_08175_),
    .Y(_08176_),
    .A1(_04914_),
    .A2(_07977_));
 sg13g2_or2_1 _17197_ (.X(_00344_),
    .B(_08176_),
    .A(_08174_));
 sg13g2_nand2_1 _17198_ (.Y(_08177_),
    .A(_07426_),
    .B(_07976_));
 sg13g2_buf_2 _17199_ (.A(_00051_),
    .X(_08178_));
 sg13g2_buf_1 _17200_ (.A(\grid.cell_17_4.se ),
    .X(_08179_));
 sg13g2_xnor2_1 _17201_ (.Y(_08180_),
    .A(_08179_),
    .B(net1141));
 sg13g2_xnor2_1 _17202_ (.Y(_08181_),
    .A(_07461_),
    .B(_08180_));
 sg13g2_xnor2_1 _17203_ (.Y(_08182_),
    .A(_07816_),
    .B(_08181_));
 sg13g2_buf_1 _17204_ (.A(_08182_),
    .X(_08183_));
 sg13g2_o21ai_1 _17205_ (.B1(_07375_),
    .Y(_08184_),
    .A1(net929),
    .A2(_08183_));
 sg13g2_inv_1 _17206_ (.Y(_08185_),
    .A(net1146));
 sg13g2_a21o_1 _17207_ (.A2(_07375_),
    .A1(_08185_),
    .B1(_08183_),
    .X(_08186_));
 sg13g2_nor2_1 _17208_ (.A(net589),
    .B(_07375_),
    .Y(_08187_));
 sg13g2_a221oi_1 _17209_ (.B2(net588),
    .C1(_08187_),
    .B1(_08186_),
    .A1(net1146),
    .Y(_08188_),
    .A2(_08184_));
 sg13g2_xnor2_1 _17210_ (.Y(_08189_),
    .A(net589),
    .B(_08183_));
 sg13g2_nor2_1 _17211_ (.A(_07829_),
    .B(_08183_),
    .Y(_08190_));
 sg13g2_a22oi_1 _17212_ (.Y(_08191_),
    .B1(_08190_),
    .B2(_08178_),
    .A2(_08189_),
    .A1(net601));
 sg13g2_o21ai_1 _17213_ (.B1(_08191_),
    .Y(_08192_),
    .A1(_08178_),
    .A2(_08188_));
 sg13g2_buf_1 _17214_ (.A(_08179_),
    .X(_08193_));
 sg13g2_inv_1 _17215_ (.Y(_08194_),
    .A(net918));
 sg13g2_buf_1 _17216_ (.A(_08194_),
    .X(_08195_));
 sg13g2_nor2_1 _17217_ (.A(net919),
    .B(net926),
    .Y(_08196_));
 sg13g2_nand2_1 _17218_ (.Y(_08197_),
    .A(net291),
    .B(_08196_));
 sg13g2_nand3_1 _17219_ (.B(net152),
    .C(_08196_),
    .A(net291),
    .Y(_08198_));
 sg13g2_buf_1 _17220_ (.A(net918),
    .X(_08199_));
 sg13g2_o21ai_1 _17221_ (.B1(net299),
    .Y(_08200_),
    .A1(net576),
    .A2(net578));
 sg13g2_nor2_1 _17222_ (.A(_08194_),
    .B(_08163_),
    .Y(_08201_));
 sg13g2_a21oi_1 _17223_ (.A1(net306),
    .A2(net594),
    .Y(_08202_),
    .B1(_08201_));
 sg13g2_nand4_1 _17224_ (.B(_08198_),
    .C(_08200_),
    .A(net1154),
    .Y(_08203_),
    .D(_08202_));
 sg13g2_o21ai_1 _17225_ (.B1(_08203_),
    .Y(_08204_),
    .A1(_07451_),
    .A2(_08197_));
 sg13g2_buf_1 _17226_ (.A(_08199_),
    .X(_08205_));
 sg13g2_nand2_1 _17227_ (.Y(_08206_),
    .A(net919),
    .B(net595));
 sg13g2_o21ai_1 _17228_ (.B1(_08206_),
    .Y(_08207_),
    .A1(net919),
    .A2(_07871_));
 sg13g2_and2_1 _17229_ (.A(net1154),
    .B(net596),
    .X(_08208_));
 sg13g2_a22oi_1 _17230_ (.Y(_08209_),
    .B1(_08207_),
    .B2(_08208_),
    .A2(_08196_),
    .A1(net594));
 sg13g2_inv_1 _17231_ (.Y(_08210_),
    .A(_08178_));
 sg13g2_nand2_1 _17232_ (.Y(_08211_),
    .A(net918),
    .B(net594));
 sg13g2_o21ai_1 _17233_ (.B1(_08211_),
    .Y(_08212_),
    .A1(net1154),
    .A2(net594));
 sg13g2_and3_1 _17234_ (.X(_08213_),
    .A(net919),
    .B(net926),
    .C(net595));
 sg13g2_and3_1 _17235_ (.X(_08214_),
    .A(_00081_),
    .B(_08132_),
    .C(net926));
 sg13g2_nor3_1 _17236_ (.A(net1154),
    .B(net1141),
    .C(net926),
    .Y(_08215_));
 sg13g2_a21oi_1 _17237_ (.A1(net919),
    .A2(net926),
    .Y(_08216_),
    .B1(_07451_));
 sg13g2_nor4_1 _17238_ (.A(_08194_),
    .B(_08214_),
    .C(_08215_),
    .D(_08216_),
    .Y(_08217_));
 sg13g2_a221oi_1 _17239_ (.B2(_08213_),
    .C1(_08217_),
    .B1(_08212_),
    .A1(_08210_),
    .Y(_08218_),
    .A2(net598));
 sg13g2_o21ai_1 _17240_ (.B1(_08218_),
    .Y(_08219_),
    .A1(_08205_),
    .A2(_08209_));
 sg13g2_a21oi_1 _17241_ (.A1(net919),
    .A2(_07835_),
    .Y(_08220_),
    .B1(net576));
 sg13g2_o21ai_1 _17242_ (.B1(net1154),
    .Y(_08221_),
    .A1(_08196_),
    .A2(_08220_));
 sg13g2_a21oi_1 _17243_ (.A1(_08197_),
    .A2(_08221_),
    .Y(_08222_),
    .B1(net152));
 sg13g2_nor3_1 _17244_ (.A(_08190_),
    .B(_08219_),
    .C(_08222_),
    .Y(_08223_));
 sg13g2_o21ai_1 _17245_ (.B1(_08189_),
    .Y(_08224_),
    .A1(_08210_),
    .A2(net601));
 sg13g2_a221oi_1 _17246_ (.B2(_08224_),
    .C1(_07194_),
    .B1(_08223_),
    .A1(_08192_),
    .Y(_08225_),
    .A2(_08204_));
 sg13g2_xnor2_1 _17247_ (.Y(_08226_),
    .A(_08111_),
    .B(_08183_));
 sg13g2_a21oi_1 _17248_ (.A1(_06057_),
    .A2(_08226_),
    .Y(_08227_),
    .B1(_07798_));
 sg13g2_or3_1 _17249_ (.A(_07976_),
    .B(_08225_),
    .C(_08227_),
    .X(_08228_));
 sg13g2_a21oi_1 _17250_ (.A1(_08177_),
    .A2(_08228_),
    .Y(_00345_),
    .B1(_07480_));
 sg13g2_buf_1 _17251_ (.A(\grid.cell_17_5.se ),
    .X(_08229_));
 sg13g2_buf_1 _17252_ (.A(_08229_),
    .X(_08230_));
 sg13g2_buf_1 _17253_ (.A(net917),
    .X(_08231_));
 sg13g2_nor4_1 _17254_ (.A(net575),
    .B(net918),
    .C(net297),
    .D(_07486_),
    .Y(_08232_));
 sg13g2_inv_1 _17255_ (.Y(_08233_),
    .A(_08230_));
 sg13g2_buf_1 _17256_ (.A(_08233_),
    .X(_08234_));
 sg13g2_a21oi_1 _17257_ (.A1(net289),
    .A2(_08194_),
    .Y(_08235_),
    .B1(net298));
 sg13g2_nor2_1 _17258_ (.A(_07486_),
    .B(net306),
    .Y(_08236_));
 sg13g2_nor2_1 _17259_ (.A(net289),
    .B(_08194_),
    .Y(_08237_));
 sg13g2_nor4_1 _17260_ (.A(_08232_),
    .B(_08235_),
    .C(_08236_),
    .D(_08237_),
    .Y(_08238_));
 sg13g2_buf_1 _17261_ (.A(net575),
    .X(_08239_));
 sg13g2_nor3_1 _17262_ (.A(_08239_),
    .B(_08205_),
    .C(net149),
    .Y(_08240_));
 sg13g2_a22oi_1 _17263_ (.Y(_08241_),
    .B1(_08240_),
    .B2(_07488_),
    .A2(_08238_),
    .A1(_07538_));
 sg13g2_buf_1 _17264_ (.A(_00083_),
    .X(_08242_));
 sg13g2_nand2_1 _17265_ (.Y(_08243_),
    .A(_08242_),
    .B(net594));
 sg13g2_xor2_1 _17266_ (.B(_07482_),
    .A(_07855_),
    .X(_08244_));
 sg13g2_xnor2_1 _17267_ (.Y(_08245_),
    .A(_08193_),
    .B(net936));
 sg13g2_xor2_1 _17268_ (.B(_08245_),
    .A(_08244_),
    .X(_08246_));
 sg13g2_xnor2_1 _17269_ (.Y(_08247_),
    .A(_08233_),
    .B(_08246_));
 sg13g2_xnor2_1 _17270_ (.Y(_08248_),
    .A(net587),
    .B(_08247_));
 sg13g2_inv_1 _17271_ (.Y(_08249_),
    .A(net1140));
 sg13g2_nand2_1 _17272_ (.Y(_08250_),
    .A(_08249_),
    .B(net596));
 sg13g2_o21ai_1 _17273_ (.B1(_08250_),
    .Y(_08251_),
    .A1(_07853_),
    .A2(_08247_));
 sg13g2_a21oi_1 _17274_ (.A1(_08243_),
    .A2(_08248_),
    .Y(_08252_),
    .B1(_08251_));
 sg13g2_xnor2_1 _17275_ (.Y(_08253_),
    .A(_08241_),
    .B(_08252_));
 sg13g2_nor2_1 _17276_ (.A(_07853_),
    .B(_08247_),
    .Y(_08254_));
 sg13g2_and2_1 _17277_ (.A(_08249_),
    .B(_07763_),
    .X(_08255_));
 sg13g2_nand2_1 _17278_ (.Y(_08256_),
    .A(_08199_),
    .B(_07887_));
 sg13g2_xnor2_1 _17279_ (.Y(_08257_),
    .A(net585),
    .B(net595));
 sg13g2_nor2_1 _17280_ (.A(_08195_),
    .B(_08257_),
    .Y(_08258_));
 sg13g2_and3_1 _17281_ (.X(_08259_),
    .A(_08195_),
    .B(net297),
    .C(net306));
 sg13g2_o21ai_1 _17282_ (.B1(net151),
    .Y(_08260_),
    .A1(_08258_),
    .A2(_08259_));
 sg13g2_o21ai_1 _17283_ (.B1(_08260_),
    .Y(_08261_),
    .A1(_07538_),
    .A2(_08256_));
 sg13g2_buf_1 _17284_ (.A(net288),
    .X(_08262_));
 sg13g2_nor3_1 _17285_ (.A(net148),
    .B(_07488_),
    .C(_08256_),
    .Y(_08263_));
 sg13g2_a221oi_1 _17286_ (.B2(net148),
    .C1(_08263_),
    .B1(_08261_),
    .A1(_08254_),
    .Y(_08264_),
    .A2(_08255_));
 sg13g2_a21oi_1 _17287_ (.A1(_08253_),
    .A2(_08264_),
    .Y(_08265_),
    .B1(_06993_));
 sg13g2_xnor2_1 _17288_ (.Y(_08266_),
    .A(_08156_),
    .B(_07763_));
 sg13g2_xnor2_1 _17289_ (.Y(_08267_),
    .A(_08247_),
    .B(_08266_));
 sg13g2_a21oi_1 _17290_ (.A1(net77),
    .A2(_08267_),
    .Y(_08268_),
    .B1(net299));
 sg13g2_or3_1 _17291_ (.A(_08041_),
    .B(_08265_),
    .C(_08268_),
    .X(_08269_));
 sg13g2_o21ai_1 _17292_ (.B1(_08269_),
    .Y(_00346_),
    .A1(_05003_),
    .A2(_07977_));
 sg13g2_buf_1 _17293_ (.A(_00145_),
    .X(_08270_));
 sg13g2_o21ai_1 _17294_ (.B1(_08002_),
    .Y(_08271_),
    .A1(net288),
    .A2(_08018_));
 sg13g2_nor2_1 _17295_ (.A(net575),
    .B(_08002_),
    .Y(_08272_));
 sg13g2_a21oi_1 _17296_ (.A1(net1139),
    .A2(_08271_),
    .Y(_08273_),
    .B1(_08272_));
 sg13g2_nand2_1 _17297_ (.Y(_08274_),
    .A(net935),
    .B(net942));
 sg13g2_nor2_1 _17298_ (.A(_08274_),
    .B(_08018_),
    .Y(_08275_));
 sg13g2_o21ai_1 _17299_ (.B1(_08275_),
    .Y(_08276_),
    .A1(net1139),
    .A2(_08002_));
 sg13g2_o21ai_1 _17300_ (.B1(_08276_),
    .Y(_08277_),
    .A1(net1139),
    .A2(_08010_));
 sg13g2_nand2b_1 _17301_ (.Y(_08278_),
    .B(_07991_),
    .A_N(net1139));
 sg13g2_and2_1 _17302_ (.A(net583),
    .B(net942),
    .X(_08279_));
 sg13g2_nor2b_1 _17303_ (.A(net917),
    .B_N(_00145_),
    .Y(_08280_));
 sg13g2_o21ai_1 _17304_ (.B1(_08280_),
    .Y(_08281_),
    .A1(_07994_),
    .A2(_08279_));
 sg13g2_o21ai_1 _17305_ (.B1(_08281_),
    .Y(_08282_),
    .A1(_07621_),
    .A2(_08278_));
 sg13g2_and2_1 _17306_ (.A(net917),
    .B(_07978_),
    .X(_08283_));
 sg13g2_buf_1 _17307_ (.A(_08283_),
    .X(_08284_));
 sg13g2_a21oi_1 _17308_ (.A1(_07896_),
    .A2(_08284_),
    .Y(_08285_),
    .B1(_08272_));
 sg13g2_nor2_1 _17309_ (.A(net151),
    .B(_08285_),
    .Y(_08286_));
 sg13g2_a221oi_1 _17310_ (.B2(net151),
    .C1(_08286_),
    .B1(_08282_),
    .A1(net288),
    .Y(_08287_),
    .A2(_08277_));
 sg13g2_o21ai_1 _17311_ (.B1(_08287_),
    .Y(_08288_),
    .A1(net153),
    .A2(_08273_));
 sg13g2_xnor2_1 _17312_ (.Y(_08289_),
    .A(_07564_),
    .B(_07980_));
 sg13g2_xnor2_1 _17313_ (.Y(_08290_),
    .A(_08231_),
    .B(_08289_));
 sg13g2_xnor2_1 _17314_ (.Y(_08291_),
    .A(_07836_),
    .B(_08290_));
 sg13g2_buf_2 _17315_ (.A(_00115_),
    .X(_08292_));
 sg13g2_inv_2 _17316_ (.Y(_08293_),
    .A(_08292_));
 sg13g2_nor2_1 _17317_ (.A(_08293_),
    .B(net152),
    .Y(_08294_));
 sg13g2_and2_1 _17318_ (.A(_07914_),
    .B(_08290_),
    .X(_08295_));
 sg13g2_a21oi_1 _17319_ (.A1(_08293_),
    .A2(net152),
    .Y(_08296_),
    .B1(_08295_));
 sg13g2_o21ai_1 _17320_ (.B1(_08296_),
    .Y(_08297_),
    .A1(_08291_),
    .A2(_08294_));
 sg13g2_xnor2_1 _17321_ (.Y(_08298_),
    .A(_08288_),
    .B(_08297_));
 sg13g2_buf_1 _17322_ (.A(net296),
    .X(_08299_));
 sg13g2_xnor2_1 _17323_ (.Y(_08300_),
    .A(_07640_),
    .B(net304));
 sg13g2_o21ai_1 _17324_ (.B1(net309),
    .Y(_08301_),
    .A1(net147),
    .A2(_07938_));
 sg13g2_a21o_1 _17325_ (.A2(_08300_),
    .A1(net147),
    .B1(_08301_),
    .X(_08302_));
 sg13g2_o21ai_1 _17326_ (.B1(_08302_),
    .Y(_08303_),
    .A1(net1139),
    .A2(_08010_));
 sg13g2_nor2_1 _17327_ (.A(net148),
    .B(_08274_),
    .Y(_08304_));
 sg13g2_a221oi_1 _17328_ (.B2(_08018_),
    .C1(net99),
    .B1(_08304_),
    .A1(net148),
    .Y(_08305_),
    .A2(_08303_));
 sg13g2_nand3_1 _17329_ (.B(_07816_),
    .C(_08295_),
    .A(_08293_),
    .Y(_08306_));
 sg13g2_xnor2_1 _17330_ (.Y(_08307_),
    .A(_08245_),
    .B(_08291_));
 sg13g2_nand2_1 _17331_ (.Y(_08308_),
    .A(net298),
    .B(_08307_));
 sg13g2_nand4_1 _17332_ (.B(_08305_),
    .C(_08306_),
    .A(_08298_),
    .Y(_08309_),
    .D(_08308_));
 sg13g2_a22oi_1 _17333_ (.Y(_08310_),
    .B1(net25),
    .B2(_07974_),
    .A2(net71),
    .A1(net149));
 sg13g2_a221oi_1 _17334_ (.B2(_08310_),
    .C1(net617),
    .B1(_08309_),
    .A1(_06814_),
    .Y(_00347_),
    .A2(_07974_));
 sg13g2_nor2_1 _17335_ (.A(net583),
    .B(net925),
    .Y(_08311_));
 sg13g2_nand2_1 _17336_ (.Y(_08312_),
    .A(_08234_),
    .B(_08311_));
 sg13g2_inv_1 _17337_ (.Y(_08313_),
    .A(_07978_));
 sg13g2_nor2_1 _17338_ (.A(_08313_),
    .B(_07866_),
    .Y(_08314_));
 sg13g2_nor2_1 _17339_ (.A(_08231_),
    .B(_08314_),
    .Y(_08315_));
 sg13g2_o21ai_1 _17340_ (.B1(_08270_),
    .Y(_08316_),
    .A1(_08311_),
    .A2(_08315_));
 sg13g2_a21oi_1 _17341_ (.A1(_08312_),
    .A2(_08316_),
    .Y(_08317_),
    .B1(net153));
 sg13g2_nand2_1 _17342_ (.Y(_08318_),
    .A(net295),
    .B(net585));
 sg13g2_nor2_1 _17343_ (.A(net1139),
    .B(_08318_),
    .Y(_08319_));
 sg13g2_nor3_1 _17344_ (.A(net1139),
    .B(net296),
    .C(net297),
    .Y(_08320_));
 sg13g2_nor3_1 _17345_ (.A(_08274_),
    .B(_08314_),
    .C(_08320_),
    .Y(_08321_));
 sg13g2_o21ai_1 _17346_ (.B1(net288),
    .Y(_08322_),
    .A1(_08319_),
    .A2(_08321_));
 sg13g2_nand2b_1 _17347_ (.Y(_08323_),
    .B(net604),
    .A_N(net1139));
 sg13g2_nor2b_1 _17348_ (.A(_07990_),
    .B_N(net925),
    .Y(_08324_));
 sg13g2_o21ai_1 _17349_ (.B1(_08280_),
    .Y(_08325_),
    .A1(_08279_),
    .A2(_08324_));
 sg13g2_o21ai_1 _17350_ (.B1(_08325_),
    .Y(_08326_),
    .A1(_08318_),
    .A2(_08323_));
 sg13g2_nand3_1 _17351_ (.B(net604),
    .C(_08284_),
    .A(_07886_),
    .Y(_08327_));
 sg13g2_a21oi_1 _17352_ (.A1(_08312_),
    .A2(_08327_),
    .Y(_08328_),
    .B1(net304));
 sg13g2_a21oi_1 _17353_ (.A1(net304),
    .A2(_08326_),
    .Y(_08329_),
    .B1(_08328_));
 sg13g2_nand3b_1 _17354_ (.B(_08322_),
    .C(_08329_),
    .Y(_08330_),
    .A_N(_08317_));
 sg13g2_xnor2_1 _17355_ (.Y(_08331_),
    .A(net917),
    .B(_07978_));
 sg13g2_xnor2_1 _17356_ (.Y(_08332_),
    .A(_08244_),
    .B(_08331_));
 sg13g2_xnor2_1 _17357_ (.Y(_08333_),
    .A(net942),
    .B(_08332_));
 sg13g2_xnor2_1 _17358_ (.Y(_08334_),
    .A(_07615_),
    .B(_08333_));
 sg13g2_o21ai_1 _17359_ (.B1(_08074_),
    .Y(_08335_),
    .A1(_07637_),
    .A2(_08333_));
 sg13g2_a21oi_1 _17360_ (.A1(_08069_),
    .A2(_08334_),
    .Y(_08336_),
    .B1(_08335_));
 sg13g2_xnor2_1 _17361_ (.Y(_08337_),
    .A(_08330_),
    .B(_08336_));
 sg13g2_nand2_1 _17362_ (.Y(_08338_),
    .A(_08299_),
    .B(_08244_));
 sg13g2_o21ai_1 _17363_ (.B1(_08338_),
    .Y(_08339_),
    .A1(_08299_),
    .A2(_07874_));
 sg13g2_a21oi_1 _17364_ (.A1(net153),
    .A2(_08339_),
    .Y(_08340_),
    .B1(_08319_));
 sg13g2_a21oi_1 _17365_ (.A1(_07533_),
    .A2(_08314_),
    .Y(_08341_),
    .B1(_08262_));
 sg13g2_a21oi_1 _17366_ (.A1(_08262_),
    .A2(_08340_),
    .Y(_08342_),
    .B1(_08341_));
 sg13g2_o21ai_1 _17367_ (.B1(_05136_),
    .Y(_08343_),
    .A1(_08086_),
    .A2(_08333_));
 sg13g2_xnor2_1 _17368_ (.Y(_08344_),
    .A(_08089_),
    .B(_08333_));
 sg13g2_nor2_1 _17369_ (.A(net150),
    .B(_08344_),
    .Y(_08345_));
 sg13g2_or4_1 _17370_ (.A(_08337_),
    .B(_08342_),
    .C(_08343_),
    .D(_08345_),
    .X(_08346_));
 sg13g2_a22oi_1 _17371_ (.Y(_08347_),
    .B1(net76),
    .B2(_07974_),
    .A2(net71),
    .A1(net150));
 sg13g2_a221oi_1 _17372_ (.B2(_08347_),
    .C1(net617),
    .B1(_08346_),
    .A1(_06471_),
    .Y(_00348_),
    .A2(_07974_));
 sg13g2_nand2_1 _17373_ (.Y(_08348_),
    .A(_07972_),
    .B(net320));
 sg13g2_buf_2 _17374_ (.A(_08348_),
    .X(_08349_));
 sg13g2_nor3_1 _17375_ (.A(_02021_),
    .B(_08349_),
    .C(_07602_),
    .Y(_08350_));
 sg13g2_buf_1 _17376_ (.A(_08350_),
    .X(_08351_));
 sg13g2_buf_1 _17377_ (.A(_08351_),
    .X(_08352_));
 sg13g2_nand2_1 _17378_ (.Y(_08353_),
    .A(net44),
    .B(net41));
 sg13g2_buf_1 _17379_ (.A(_00220_),
    .X(_08354_));
 sg13g2_buf_1 _17380_ (.A(net1138),
    .X(_08355_));
 sg13g2_buf_1 _17381_ (.A(\grid.cell_18_0.se ),
    .X(_08356_));
 sg13g2_xor2_1 _17382_ (.B(_08356_),
    .A(net1152),
    .X(_08357_));
 sg13g2_buf_1 _17383_ (.A(\grid.cell_18_0.sw ),
    .X(_08358_));
 sg13g2_buf_1 _17384_ (.A(_08358_),
    .X(_08359_));
 sg13g2_xnor2_1 _17385_ (.Y(_08360_),
    .A(net915),
    .B(_07980_));
 sg13g2_xnor2_1 _17386_ (.Y(_08361_),
    .A(_08357_),
    .B(_08360_));
 sg13g2_nor2_1 _17387_ (.A(_08108_),
    .B(_08361_),
    .Y(_08362_));
 sg13g2_xnor2_1 _17388_ (.Y(_08363_),
    .A(_08009_),
    .B(_08357_));
 sg13g2_xnor2_1 _17389_ (.Y(_08364_),
    .A(_08360_),
    .B(_08363_));
 sg13g2_buf_1 _17390_ (.A(_08364_),
    .X(_08365_));
 sg13g2_o21ai_1 _17391_ (.B1(_08365_),
    .Y(_08366_),
    .A1(net916),
    .A2(_08362_));
 sg13g2_nor2_1 _17392_ (.A(net1138),
    .B(_08365_),
    .Y(_08367_));
 sg13g2_a21o_1 _17393_ (.A2(_08365_),
    .A1(_07702_),
    .B1(net1138),
    .X(_08368_));
 sg13g2_mux2_1 _17394_ (.A0(_08367_),
    .A1(_08368_),
    .S(_08362_),
    .X(_08369_));
 sg13g2_a21o_1 _17395_ (.A2(_08366_),
    .A1(net933),
    .B1(_08369_),
    .X(_08370_));
 sg13g2_buf_1 _17396_ (.A(_08356_),
    .X(_08371_));
 sg13g2_buf_1 _17397_ (.A(net914),
    .X(_08372_));
 sg13g2_buf_1 _17398_ (.A(net574),
    .X(_08373_));
 sg13g2_nor2_1 _17399_ (.A(net915),
    .B(_07989_),
    .Y(_08374_));
 sg13g2_buf_2 _17400_ (.A(_08374_),
    .X(_08375_));
 sg13g2_and2_1 _17401_ (.A(net915),
    .B(net923),
    .X(_08376_));
 sg13g2_buf_2 _17402_ (.A(_08376_),
    .X(_08377_));
 sg13g2_buf_1 _17403_ (.A(net915),
    .X(_08378_));
 sg13g2_nand2b_1 _17404_ (.Y(_08379_),
    .B(net573),
    .A_N(net923));
 sg13g2_nand2b_1 _17405_ (.Y(_08380_),
    .B(net923),
    .A_N(_08359_));
 sg13g2_buf_1 _17406_ (.A(_08380_),
    .X(_08381_));
 sg13g2_nand2_1 _17407_ (.Y(_08382_),
    .A(_08379_),
    .B(_08381_));
 sg13g2_nand2_1 _17408_ (.Y(_08383_),
    .A(net931),
    .B(_08382_));
 sg13g2_o21ai_1 _17409_ (.B1(_08383_),
    .Y(_08384_),
    .A1(net150),
    .A2(_08377_));
 sg13g2_a22oi_1 _17410_ (.Y(_08385_),
    .B1(_08384_),
    .B2(net928),
    .A2(_08375_),
    .A1(_07655_));
 sg13g2_a21oi_1 _17411_ (.A1(net932),
    .A2(net574),
    .Y(_08386_),
    .B1(net303));
 sg13g2_nand3b_1 _17412_ (.B(_08375_),
    .C(net928),
    .Y(_08387_),
    .A_N(_08386_));
 sg13g2_o21ai_1 _17413_ (.B1(_08387_),
    .Y(_08388_),
    .A1(net287),
    .A2(_08385_));
 sg13g2_nand2_1 _17414_ (.Y(_08389_),
    .A(net916),
    .B(_08365_));
 sg13g2_o21ai_1 _17415_ (.B1(_08389_),
    .Y(_08390_),
    .A1(net933),
    .A2(_08367_));
 sg13g2_inv_1 _17416_ (.Y(_08391_),
    .A(net914));
 sg13g2_buf_1 _17417_ (.A(net573),
    .X(_08392_));
 sg13g2_nand2_1 _17418_ (.Y(_08393_),
    .A(net286),
    .B(net296));
 sg13g2_nor3_1 _17419_ (.A(_08391_),
    .B(_07716_),
    .C(_08393_),
    .Y(_08394_));
 sg13g2_buf_1 _17420_ (.A(net286),
    .X(_08395_));
 sg13g2_nor4_1 _17421_ (.A(_08372_),
    .B(net146),
    .C(net147),
    .D(net303),
    .Y(_08396_));
 sg13g2_o21ai_1 _17422_ (.B1(net591),
    .Y(_08397_),
    .A1(_08394_),
    .A2(_08396_));
 sg13g2_nand2b_1 _17423_ (.Y(_08398_),
    .B(_07990_),
    .A_N(_07715_));
 sg13g2_nand2_1 _17424_ (.Y(_08399_),
    .A(net573),
    .B(_08398_));
 sg13g2_nand2_1 _17425_ (.Y(_08400_),
    .A(_08381_),
    .B(_08399_));
 sg13g2_inv_1 _17426_ (.Y(_08401_),
    .A(_08359_));
 sg13g2_buf_1 _17427_ (.A(_08401_),
    .X(_08402_));
 sg13g2_nand2_1 _17428_ (.Y(_08403_),
    .A(net285),
    .B(net592));
 sg13g2_a21oi_1 _17429_ (.A1(_08379_),
    .A2(_08403_),
    .Y(_08404_),
    .B1(net931));
 sg13g2_a221oi_1 _17430_ (.B2(net303),
    .C1(_08404_),
    .B1(_08400_),
    .A1(_07716_),
    .Y(_08405_),
    .A2(_08375_));
 sg13g2_inv_1 _17431_ (.Y(_08406_),
    .A(_08375_));
 sg13g2_o21ai_1 _17432_ (.B1(_07997_),
    .Y(_08407_),
    .A1(_07993_),
    .A2(_07715_));
 sg13g2_nor2_1 _17433_ (.A(net286),
    .B(_08398_),
    .Y(_08408_));
 sg13g2_a221oi_1 _17434_ (.B2(net286),
    .C1(_08408_),
    .B1(_08407_),
    .A1(_07634_),
    .Y(_08409_),
    .A2(_08406_));
 sg13g2_mux2_1 _17435_ (.A0(_08405_),
    .A1(_08409_),
    .S(_08391_),
    .X(_08410_));
 sg13g2_a21oi_1 _17436_ (.A1(_08397_),
    .A2(_08410_),
    .Y(_08411_),
    .B1(_08362_));
 sg13g2_a221oi_1 _17437_ (.B2(_08411_),
    .C1(_07194_),
    .B1(_08390_),
    .A1(_08370_),
    .Y(_08412_),
    .A2(_08388_));
 sg13g2_buf_1 _17438_ (.A(\grid.cell_18_0.s ),
    .X(_08413_));
 sg13g2_buf_1 _17439_ (.A(_08413_),
    .X(_08414_));
 sg13g2_buf_1 _17440_ (.A(net913),
    .X(_08415_));
 sg13g2_xor2_1 _17441_ (.B(_08415_),
    .A(net933),
    .X(_08416_));
 sg13g2_xnor2_1 _17442_ (.Y(_08417_),
    .A(_08365_),
    .B(_08416_));
 sg13g2_a21oi_1 _17443_ (.A1(net109),
    .A2(_08417_),
    .Y(_08418_),
    .B1(net582));
 sg13g2_or3_1 _17444_ (.A(net41),
    .B(_08412_),
    .C(_08418_),
    .X(_08419_));
 sg13g2_a21oi_1 _17445_ (.A1(_08353_),
    .A2(_08419_),
    .Y(_00349_),
    .B1(net305));
 sg13g2_xor2_1 _17446_ (.B(_08035_),
    .A(_07614_),
    .X(_08420_));
 sg13g2_buf_1 _17447_ (.A(\grid.cell_18_1.se ),
    .X(_08421_));
 sg13g2_inv_2 _17448_ (.Y(_08422_),
    .A(net1137));
 sg13g2_xnor2_1 _17449_ (.Y(_08423_),
    .A(_08422_),
    .B(_08079_));
 sg13g2_xnor2_1 _17450_ (.Y(_08424_),
    .A(_08357_),
    .B(_08423_));
 sg13g2_nor4_1 _17451_ (.A(_08355_),
    .B(net1142),
    .C(_08420_),
    .D(_08424_),
    .Y(_08425_));
 sg13g2_buf_1 _17452_ (.A(net1137),
    .X(_08426_));
 sg13g2_nand2_1 _17453_ (.Y(_08427_),
    .A(net921),
    .B(net912));
 sg13g2_nand2_1 _17454_ (.Y(_08428_),
    .A(net1152),
    .B(net1151));
 sg13g2_nor3_1 _17455_ (.A(net287),
    .B(_08427_),
    .C(_08428_),
    .Y(_08429_));
 sg13g2_nor2b_1 _17456_ (.A(_07715_),
    .B_N(net1137),
    .Y(_08430_));
 sg13g2_xor2_1 _17457_ (.B(net1137),
    .A(_08044_),
    .X(_08431_));
 sg13g2_nand2_1 _17458_ (.Y(_08432_),
    .A(net931),
    .B(_08431_));
 sg13g2_o21ai_1 _17459_ (.B1(_08432_),
    .Y(_08433_),
    .A1(net931),
    .A2(_08427_));
 sg13g2_a22oi_1 _17460_ (.Y(_08434_),
    .B1(_08433_),
    .B2(net301),
    .A2(_08430_),
    .A1(_08066_));
 sg13g2_nor2_1 _17461_ (.A(_08391_),
    .B(_08434_),
    .Y(_08435_));
 sg13g2_or3_1 _17462_ (.A(_08425_),
    .B(_08429_),
    .C(_08435_),
    .X(_08436_));
 sg13g2_nand2_1 _17463_ (.Y(_08437_),
    .A(_07702_),
    .B(_08354_));
 sg13g2_xnor2_1 _17464_ (.Y(_08438_),
    .A(_08035_),
    .B(_08424_));
 sg13g2_nand2b_1 _17465_ (.Y(_08439_),
    .B(net933),
    .A_N(_08354_));
 sg13g2_o21ai_1 _17466_ (.B1(_08439_),
    .Y(_08440_),
    .A1(net1142),
    .A2(_08424_));
 sg13g2_a21oi_1 _17467_ (.A1(_08437_),
    .A2(_08438_),
    .Y(_08441_),
    .B1(_08440_));
 sg13g2_buf_1 _17468_ (.A(net912),
    .X(_08442_));
 sg13g2_and2_1 _17469_ (.A(net1152),
    .B(net930),
    .X(_08443_));
 sg13g2_o21ai_1 _17470_ (.B1(_08443_),
    .Y(_08444_),
    .A1(net571),
    .A2(net928));
 sg13g2_nor2_1 _17471_ (.A(net912),
    .B(_08428_),
    .Y(_08445_));
 sg13g2_o21ai_1 _17472_ (.B1(net581),
    .Y(_08446_),
    .A1(_08430_),
    .A2(_08445_));
 sg13g2_o21ai_1 _17473_ (.B1(_08446_),
    .Y(_08447_),
    .A1(net294),
    .A2(_08444_));
 sg13g2_nand2b_1 _17474_ (.Y(_08448_),
    .B(_07715_),
    .A_N(net1137));
 sg13g2_o21ai_1 _17475_ (.B1(_08448_),
    .Y(_08449_),
    .A1(_08045_),
    .A2(_08430_));
 sg13g2_o21ai_1 _17476_ (.B1(_08045_),
    .Y(_08450_),
    .A1(net1137),
    .A2(_07715_));
 sg13g2_o21ai_1 _17477_ (.B1(_08450_),
    .Y(_08451_),
    .A1(_08422_),
    .A2(_07716_));
 sg13g2_a22oi_1 _17478_ (.Y(_08452_),
    .B1(_08451_),
    .B2(_08443_),
    .A2(_08449_),
    .A1(_07749_));
 sg13g2_nor2_1 _17479_ (.A(_08426_),
    .B(_07716_),
    .Y(_08453_));
 sg13g2_or3_1 _17480_ (.A(_08371_),
    .B(net921),
    .C(_08421_),
    .X(_08454_));
 sg13g2_nand4_1 _17481_ (.B(net1151),
    .C(net921),
    .A(_08372_),
    .Y(_08455_),
    .D(_08426_));
 sg13g2_a21oi_1 _17482_ (.A1(_08454_),
    .A2(_08455_),
    .Y(_08456_),
    .B1(net931));
 sg13g2_a21oi_1 _17483_ (.A1(_08048_),
    .A2(_08453_),
    .Y(_08457_),
    .B1(_08456_));
 sg13g2_o21ai_1 _17484_ (.B1(_08457_),
    .Y(_08458_),
    .A1(_08373_),
    .A2(_08452_));
 sg13g2_a21oi_1 _17485_ (.A1(_08373_),
    .A2(_08447_),
    .Y(_08459_),
    .B1(_08458_));
 sg13g2_xor2_1 _17486_ (.B(_08459_),
    .A(_08441_),
    .X(_08460_));
 sg13g2_o21ai_1 _17487_ (.B1(_05416_),
    .Y(_08461_),
    .A1(_08436_),
    .A2(_08460_));
 sg13g2_xnor2_1 _17488_ (.Y(_08462_),
    .A(net913),
    .B(_08088_));
 sg13g2_xnor2_1 _17489_ (.Y(_08463_),
    .A(_08424_),
    .B(_08462_));
 sg13g2_a21oi_1 _17490_ (.A1(_05619_),
    .A2(_08463_),
    .Y(_08464_),
    .B1(_07988_));
 sg13g2_nor2_1 _17491_ (.A(net41),
    .B(_08464_),
    .Y(_08465_));
 sg13g2_a22oi_1 _17492_ (.Y(_08466_),
    .B1(_08461_),
    .B2(_08465_),
    .A2(net41),
    .A1(net42));
 sg13g2_nor2_1 _17493_ (.A(net370),
    .B(_08466_),
    .Y(_00350_));
 sg13g2_nand2_1 _17494_ (.Y(_08467_),
    .A(_05354_),
    .B(_08351_));
 sg13g2_buf_2 _17495_ (.A(\grid.cell_18_2.se ),
    .X(_08468_));
 sg13g2_buf_1 _17496_ (.A(_08468_),
    .X(_08469_));
 sg13g2_inv_2 _17497_ (.Y(_08470_),
    .A(net911));
 sg13g2_nor2_1 _17498_ (.A(_08470_),
    .B(_08165_),
    .Y(_08471_));
 sg13g2_xnor2_1 _17499_ (.Y(_08472_),
    .A(_08468_),
    .B(_08095_));
 sg13g2_nand2b_1 _17500_ (.Y(_08473_),
    .B(net1151),
    .A_N(_08472_));
 sg13g2_o21ai_1 _17501_ (.B1(_08473_),
    .Y(_08474_),
    .A1(net929),
    .A2(_08471_));
 sg13g2_nand2_1 _17502_ (.Y(_08475_),
    .A(net590),
    .B(net929));
 sg13g2_buf_1 _17503_ (.A(net911),
    .X(_08476_));
 sg13g2_nor2_1 _17504_ (.A(net570),
    .B(net920),
    .Y(_08477_));
 sg13g2_a22oi_1 _17505_ (.Y(_08478_),
    .B1(_08475_),
    .B2(_08477_),
    .A2(_08474_),
    .A1(net1149));
 sg13g2_o21ai_1 _17506_ (.B1(net589),
    .Y(_08479_),
    .A1(_07749_),
    .A2(_08422_));
 sg13g2_nand3_1 _17507_ (.B(_08479_),
    .C(_08477_),
    .A(net1149),
    .Y(_08480_));
 sg13g2_o21ai_1 _17508_ (.B1(_08480_),
    .Y(_08481_),
    .A1(net571),
    .A2(_08478_));
 sg13g2_buf_1 _17509_ (.A(_00211_),
    .X(_08482_));
 sg13g2_inv_1 _17510_ (.Y(_08483_),
    .A(_08482_));
 sg13g2_nor2_1 _17511_ (.A(net932),
    .B(_08483_),
    .Y(_08484_));
 sg13g2_xnor2_1 _17512_ (.Y(_08485_),
    .A(_07728_),
    .B(_08472_));
 sg13g2_xnor2_1 _17513_ (.Y(_08486_),
    .A(_08421_),
    .B(_08485_));
 sg13g2_xnor2_1 _17514_ (.Y(_08487_),
    .A(net924),
    .B(_08486_));
 sg13g2_a22oi_1 _17515_ (.Y(_08488_),
    .B1(_08114_),
    .B2(_08486_),
    .A2(_08483_),
    .A1(net932));
 sg13g2_o21ai_1 _17516_ (.B1(_08488_),
    .Y(_08489_),
    .A1(_08484_),
    .A2(_08487_));
 sg13g2_xnor2_1 _17517_ (.Y(_08490_),
    .A(_08481_),
    .B(_08489_));
 sg13g2_nand2_1 _17518_ (.Y(_08491_),
    .A(net911),
    .B(net920));
 sg13g2_o21ai_1 _17519_ (.B1(_08473_),
    .Y(_08492_),
    .A1(net930),
    .A2(_08491_));
 sg13g2_nand2_1 _17520_ (.Y(_08493_),
    .A(net589),
    .B(_08492_));
 sg13g2_o21ai_1 _17521_ (.B1(_08493_),
    .Y(_08494_),
    .A1(net1149),
    .A2(_08491_));
 sg13g2_nor3_1 _17522_ (.A(_07749_),
    .B(_08442_),
    .C(_08097_),
    .Y(_08495_));
 sg13g2_buf_1 _17523_ (.A(net570),
    .X(_08496_));
 sg13g2_xnor2_1 _17524_ (.Y(_08497_),
    .A(net931),
    .B(net924));
 sg13g2_and4_1 _17525_ (.A(_08483_),
    .B(_08114_),
    .C(_08497_),
    .D(_08486_),
    .X(_08498_));
 sg13g2_a221oi_1 _17526_ (.B2(_08496_),
    .C1(_08498_),
    .B1(_08495_),
    .A1(_08442_),
    .Y(_08499_),
    .A2(_08494_));
 sg13g2_a21oi_1 _17527_ (.A1(_08490_),
    .A2(_08499_),
    .Y(_08500_),
    .B1(net106));
 sg13g2_xor2_1 _17528_ (.B(_08486_),
    .A(_08363_),
    .X(_08501_));
 sg13g2_a21oi_1 _17529_ (.A1(net111),
    .A2(_08501_),
    .Y(_08502_),
    .B1(net294));
 sg13g2_or4_1 _17530_ (.A(_00659_),
    .B(net41),
    .C(_08500_),
    .D(_08502_),
    .X(_08503_));
 sg13g2_o21ai_1 _17531_ (.B1(_08503_),
    .Y(_00351_),
    .A1(_04088_),
    .A2(_08467_));
 sg13g2_buf_1 _17532_ (.A(\grid.cell_18_3.se ),
    .X(_08504_));
 sg13g2_buf_1 _17533_ (.A(_08504_),
    .X(_08505_));
 sg13g2_buf_1 _17534_ (.A(net910),
    .X(_08506_));
 sg13g2_buf_1 _17535_ (.A(net569),
    .X(_08507_));
 sg13g2_nor2_1 _17536_ (.A(_08507_),
    .B(net284),
    .Y(_08508_));
 sg13g2_nor2_1 _17537_ (.A(_08156_),
    .B(_07788_),
    .Y(_08509_));
 sg13g2_nand2_1 _17538_ (.Y(_08510_),
    .A(net911),
    .B(net1141));
 sg13g2_o21ai_1 _17539_ (.B1(_08510_),
    .Y(_08511_),
    .A1(_07788_),
    .A2(net588));
 sg13g2_a21oi_1 _17540_ (.A1(_08508_),
    .A2(_08509_),
    .Y(_08512_),
    .B1(_08511_));
 sg13g2_o21ai_1 _17541_ (.B1(_08507_),
    .Y(_08513_),
    .A1(_08496_),
    .A2(net578));
 sg13g2_and2_1 _17542_ (.A(net1146),
    .B(_08513_),
    .X(_08514_));
 sg13g2_nor3_1 _17543_ (.A(net910),
    .B(net570),
    .C(net919),
    .Y(_08515_));
 sg13g2_nand2_1 _17544_ (.Y(_08516_),
    .A(net300),
    .B(net588));
 sg13g2_a22oi_1 _17545_ (.Y(_08517_),
    .B1(_08515_),
    .B2(_08516_),
    .A2(_08514_),
    .A1(_08512_));
 sg13g2_xor2_1 _17546_ (.B(net1148),
    .A(net910),
    .X(_08518_));
 sg13g2_xnor2_1 _17547_ (.Y(_08519_),
    .A(_08132_),
    .B(net1150));
 sg13g2_xnor2_1 _17548_ (.Y(_08520_),
    .A(_08518_),
    .B(_08519_));
 sg13g2_xnor2_1 _17549_ (.Y(_08521_),
    .A(net911),
    .B(_08520_));
 sg13g2_xnor2_1 _17550_ (.Y(_08522_),
    .A(net581),
    .B(_08521_));
 sg13g2_nor2_1 _17551_ (.A(_08137_),
    .B(_08521_),
    .Y(_08523_));
 sg13g2_a21oi_1 _17552_ (.A1(net301),
    .A2(_08522_),
    .Y(_08524_),
    .B1(_08523_));
 sg13g2_inv_1 _17553_ (.Y(_08525_),
    .A(_00210_));
 sg13g2_xnor2_1 _17554_ (.Y(_08526_),
    .A(_08079_),
    .B(_08521_));
 sg13g2_nand2_1 _17555_ (.Y(_08527_),
    .A(_08525_),
    .B(_08526_));
 sg13g2_xnor2_1 _17556_ (.Y(_08528_),
    .A(_08524_),
    .B(_08527_));
 sg13g2_inv_1 _17557_ (.Y(_08529_),
    .A(net910));
 sg13g2_buf_1 _17558_ (.A(_08529_),
    .X(_08530_));
 sg13g2_nand2_1 _17559_ (.Y(_08531_),
    .A(net911),
    .B(net927));
 sg13g2_o21ai_1 _17560_ (.B1(_08531_),
    .Y(_08532_),
    .A1(_08476_),
    .A2(_08163_));
 sg13g2_nand3_1 _17561_ (.B(_08530_),
    .C(_08532_),
    .A(net1146),
    .Y(_08533_));
 sg13g2_nand4_1 _17562_ (.B(_08476_),
    .C(net578),
    .A(_08185_),
    .Y(_08534_),
    .D(net587));
 sg13g2_nand3_1 _17563_ (.B(_08533_),
    .C(_08534_),
    .A(net588),
    .Y(_08535_));
 sg13g2_nor4_1 _17564_ (.A(_08530_),
    .B(_08470_),
    .C(_08163_),
    .D(_07788_),
    .Y(_08536_));
 sg13g2_or3_1 _17565_ (.A(net588),
    .B(_08515_),
    .C(_08536_),
    .X(_08537_));
 sg13g2_nor2_1 _17566_ (.A(_08469_),
    .B(net1141),
    .Y(_08538_));
 sg13g2_nand2_1 _17567_ (.Y(_08539_),
    .A(_08185_),
    .B(_08538_));
 sg13g2_nand4_1 _17568_ (.B(net589),
    .C(_08510_),
    .A(net587),
    .Y(_08540_),
    .D(_08539_));
 sg13g2_o21ai_1 _17569_ (.B1(_08540_),
    .Y(_08541_),
    .A1(net1146),
    .A2(_08510_));
 sg13g2_a21o_1 _17570_ (.A2(_08510_),
    .A1(net282),
    .B1(_08538_),
    .X(_08542_));
 sg13g2_a21oi_1 _17571_ (.A1(net1146),
    .A2(_08542_),
    .Y(_08543_),
    .B1(_08515_));
 sg13g2_nor2_1 _17572_ (.A(net300),
    .B(_08543_),
    .Y(_08544_));
 sg13g2_a221oi_1 _17573_ (.B2(net283),
    .C1(_08544_),
    .B1(_08541_),
    .A1(_08535_),
    .Y(_08545_),
    .A2(_08537_));
 sg13g2_a221oi_1 _17574_ (.B2(_08525_),
    .C1(_08523_),
    .B1(_08526_),
    .A1(net301),
    .Y(_08546_),
    .A2(_08522_));
 sg13g2_a21oi_1 _17575_ (.A1(_08545_),
    .A2(_08546_),
    .Y(_08547_),
    .B1(net99));
 sg13g2_o21ai_1 _17576_ (.B1(_08547_),
    .Y(_08548_),
    .A1(_08517_),
    .A2(_08528_));
 sg13g2_buf_1 _17577_ (.A(net171),
    .X(_08549_));
 sg13g2_xnor2_1 _17578_ (.Y(_08550_),
    .A(_08423_),
    .B(_08521_));
 sg13g2_a21oi_1 _17579_ (.A1(net98),
    .A2(_08550_),
    .Y(_08551_),
    .B1(net293));
 sg13g2_nor2_1 _17580_ (.A(net41),
    .B(_08551_),
    .Y(_08552_));
 sg13g2_a22oi_1 _17581_ (.Y(_08553_),
    .B1(_08548_),
    .B2(_08552_),
    .A2(net41),
    .A1(_06621_));
 sg13g2_nor2_1 _17582_ (.A(_02970_),
    .B(_08553_),
    .Y(_00352_));
 sg13g2_buf_1 _17583_ (.A(\grid.cell_18_4.se ),
    .X(_08554_));
 sg13g2_buf_1 _17584_ (.A(net1136),
    .X(_08555_));
 sg13g2_nor4_1 _17585_ (.A(net909),
    .B(net910),
    .C(net918),
    .D(_07871_),
    .Y(_08556_));
 sg13g2_a221oi_1 _17586_ (.B2(_07788_),
    .C1(_08556_),
    .B1(net586),
    .A1(_08506_),
    .Y(_08557_),
    .A2(net576));
 sg13g2_o21ai_1 _17587_ (.B1(net909),
    .Y(_08558_),
    .A1(net910),
    .A2(net918));
 sg13g2_and2_1 _17588_ (.A(_07853_),
    .B(_08558_),
    .X(_08559_));
 sg13g2_nor3_1 _17589_ (.A(net909),
    .B(_08506_),
    .C(net290),
    .Y(_08560_));
 sg13g2_nand2_1 _17590_ (.Y(_08561_),
    .A(net586),
    .B(net587));
 sg13g2_a22oi_1 _17591_ (.Y(_08562_),
    .B1(_08560_),
    .B2(_08561_),
    .A2(_08559_),
    .A1(_08557_));
 sg13g2_buf_1 _17592_ (.A(_00050_),
    .X(_08563_));
 sg13g2_inv_1 _17593_ (.Y(_08564_),
    .A(net589));
 sg13g2_nand2_1 _17594_ (.Y(_08565_),
    .A(net1135),
    .B(_08564_));
 sg13g2_xnor2_1 _17595_ (.Y(_08566_),
    .A(net1136),
    .B(_08179_));
 sg13g2_xnor2_1 _17596_ (.Y(_08567_),
    .A(net1147),
    .B(_08566_));
 sg13g2_xnor2_1 _17597_ (.Y(_08568_),
    .A(_08518_),
    .B(_08567_));
 sg13g2_xnor2_1 _17598_ (.Y(_08569_),
    .A(net579),
    .B(_08568_));
 sg13g2_nand2b_1 _17599_ (.Y(_08570_),
    .B(net589),
    .A_N(net1135));
 sg13g2_o21ai_1 _17600_ (.B1(_08570_),
    .Y(_08571_),
    .A1(_08178_),
    .A2(_08568_));
 sg13g2_a21oi_1 _17601_ (.A1(_08565_),
    .A2(_08569_),
    .Y(_08572_),
    .B1(_08571_));
 sg13g2_xnor2_1 _17602_ (.Y(_08573_),
    .A(_08562_),
    .B(_08572_));
 sg13g2_nor4_1 _17603_ (.A(_08178_),
    .B(net1135),
    .C(_08099_),
    .D(_08568_),
    .Y(_08574_));
 sg13g2_buf_1 _17604_ (.A(net909),
    .X(_08575_));
 sg13g2_nand2_1 _17605_ (.Y(_08576_),
    .A(_08505_),
    .B(net576));
 sg13g2_xnor2_1 _17606_ (.Y(_08577_),
    .A(net918),
    .B(net927));
 sg13g2_nor2_1 _17607_ (.A(_08529_),
    .B(_08577_),
    .Y(_08578_));
 sg13g2_nor3_1 _17608_ (.A(net910),
    .B(_08194_),
    .C(_07788_),
    .Y(_08579_));
 sg13g2_o21ai_1 _17609_ (.B1(net586),
    .Y(_08580_),
    .A1(_08578_),
    .A2(_08579_));
 sg13g2_o21ai_1 _17610_ (.B1(_08580_),
    .Y(_08581_),
    .A1(_07853_),
    .A2(_08576_));
 sg13g2_nor3_1 _17611_ (.A(net568),
    .B(_08561_),
    .C(_08576_),
    .Y(_08582_));
 sg13g2_a21oi_1 _17612_ (.A1(net568),
    .A2(_08581_),
    .Y(_08583_),
    .B1(_08582_));
 sg13g2_nor2b_1 _17613_ (.A(_08574_),
    .B_N(_08583_),
    .Y(_08584_));
 sg13g2_a21oi_1 _17614_ (.A1(_08573_),
    .A2(_08584_),
    .Y(_08585_),
    .B1(net105));
 sg13g2_buf_1 _17615_ (.A(net123),
    .X(_08586_));
 sg13g2_xnor2_1 _17616_ (.Y(_08587_),
    .A(net588),
    .B(_08472_));
 sg13g2_xnor2_1 _17617_ (.Y(_08588_),
    .A(_08568_),
    .B(_08587_));
 sg13g2_a21oi_1 _17618_ (.A1(net70),
    .A2(_08588_),
    .Y(_08589_),
    .B1(net292));
 sg13g2_nor4_1 _17619_ (.A(_06110_),
    .B(_08352_),
    .C(_08585_),
    .D(_08589_),
    .Y(_08590_));
 sg13g2_nor2_1 _17620_ (.A(net47),
    .B(_08467_),
    .Y(_08591_));
 sg13g2_or2_1 _17621_ (.X(_00353_),
    .B(_08591_),
    .A(_08590_));
 sg13g2_buf_1 _17622_ (.A(\grid.cell_18_5.se ),
    .X(_08592_));
 sg13g2_buf_1 _17623_ (.A(net1134),
    .X(_08593_));
 sg13g2_xnor2_1 _17624_ (.Y(_08594_),
    .A(net1136),
    .B(net1147));
 sg13g2_xnor2_1 _17625_ (.Y(_08595_),
    .A(_08229_),
    .B(_07855_));
 sg13g2_xnor2_1 _17626_ (.Y(_08596_),
    .A(_08594_),
    .B(_08595_));
 sg13g2_xnor2_1 _17627_ (.Y(_08597_),
    .A(net908),
    .B(_08596_));
 sg13g2_xnor2_1 _17628_ (.Y(_08598_),
    .A(_08164_),
    .B(_08597_));
 sg13g2_and2_1 _17629_ (.A(_08249_),
    .B(_08597_),
    .X(_08599_));
 sg13g2_buf_1 _17630_ (.A(_00082_),
    .X(_08600_));
 sg13g2_a21o_1 _17631_ (.A2(_08597_),
    .A1(_08164_),
    .B1(net587),
    .X(_08601_));
 sg13g2_o21ai_1 _17632_ (.B1(_08597_),
    .Y(_08602_),
    .A1(_08242_),
    .A2(net300));
 sg13g2_a221oi_1 _17633_ (.B2(_08171_),
    .C1(_08509_),
    .B1(_08602_),
    .A1(net1140),
    .Y(_08603_),
    .A2(_08601_));
 sg13g2_nor2_1 _17634_ (.A(net1133),
    .B(_08603_),
    .Y(_08604_));
 sg13g2_a221oi_1 _17635_ (.B2(net1133),
    .C1(_08604_),
    .B1(_08599_),
    .A1(net300),
    .Y(_08605_),
    .A2(_08598_));
 sg13g2_buf_1 _17636_ (.A(net908),
    .X(_08606_));
 sg13g2_buf_1 _17637_ (.A(net567),
    .X(_08607_));
 sg13g2_or2_1 _17638_ (.X(_08608_),
    .B(net917),
    .A(_08554_));
 sg13g2_buf_1 _17639_ (.A(_08608_),
    .X(_08609_));
 sg13g2_nor3_1 _17640_ (.A(net281),
    .B(net298),
    .C(_08609_),
    .Y(_08610_));
 sg13g2_inv_2 _17641_ (.Y(_08611_),
    .A(net1136));
 sg13g2_nor2_2 _17642_ (.A(_08611_),
    .B(net289),
    .Y(_08612_));
 sg13g2_inv_1 _17643_ (.Y(_08613_),
    .A(net908));
 sg13g2_nor2_1 _17644_ (.A(net566),
    .B(_08234_),
    .Y(_08614_));
 sg13g2_buf_1 _17645_ (.A(net567),
    .X(_08615_));
 sg13g2_nand2_1 _17646_ (.Y(_08616_),
    .A(net280),
    .B(net568));
 sg13g2_o21ai_1 _17647_ (.B1(_08616_),
    .Y(_08617_),
    .A1(net298),
    .A2(net299));
 sg13g2_nor4_1 _17648_ (.A(_08610_),
    .B(_08612_),
    .C(_08614_),
    .D(_08617_),
    .Y(_08618_));
 sg13g2_nor2_1 _17649_ (.A(_08606_),
    .B(_08609_),
    .Y(_08619_));
 sg13g2_a22oi_1 _17650_ (.Y(_08620_),
    .B1(_08619_),
    .B2(_07875_),
    .A2(_08618_),
    .A1(_07913_));
 sg13g2_mux2_1 _17651_ (.A0(net575),
    .A1(net585),
    .S(_08554_),
    .X(_08621_));
 sg13g2_nand3_1 _17652_ (.B(net586),
    .C(_08621_),
    .A(net1144),
    .Y(_08622_));
 sg13g2_o21ai_1 _17653_ (.B1(_08622_),
    .Y(_08623_),
    .A1(net586),
    .A2(_08609_));
 sg13g2_nand2_1 _17654_ (.Y(_08624_),
    .A(net566),
    .B(_08623_));
 sg13g2_a21oi_1 _17655_ (.A1(net297),
    .A2(net586),
    .Y(_08625_),
    .B1(_08612_));
 sg13g2_nor2_1 _17656_ (.A(net1144),
    .B(_08609_),
    .Y(_08626_));
 sg13g2_a21oi_1 _17657_ (.A1(net1144),
    .A2(_08612_),
    .Y(_08627_),
    .B1(_08626_));
 sg13g2_nand3b_1 _17658_ (.B(_08627_),
    .C(_08615_),
    .Y(_08628_),
    .A_N(_08625_));
 sg13g2_nand2_1 _17659_ (.Y(_08629_),
    .A(net567),
    .B(_07871_));
 sg13g2_o21ai_1 _17660_ (.B1(_08629_),
    .Y(_08630_),
    .A1(net1144),
    .A2(_07871_));
 sg13g2_nand3_1 _17661_ (.B(_08612_),
    .C(_08630_),
    .A(net149),
    .Y(_08631_));
 sg13g2_nand2b_1 _17662_ (.Y(_08632_),
    .B(net300),
    .A_N(_08600_));
 sg13g2_nand4_1 _17663_ (.B(_08628_),
    .C(_08631_),
    .A(_08624_),
    .Y(_08633_),
    .D(_08632_));
 sg13g2_o21ai_1 _17664_ (.B1(_08609_),
    .Y(_08634_),
    .A1(_08606_),
    .A2(_08612_));
 sg13g2_a21oi_1 _17665_ (.A1(net1144),
    .A2(_08634_),
    .Y(_08635_),
    .B1(_08619_));
 sg13g2_nor2_1 _17666_ (.A(net149),
    .B(_08635_),
    .Y(_08636_));
 sg13g2_nand2_1 _17667_ (.Y(_08637_),
    .A(_08600_),
    .B(_07788_));
 sg13g2_and2_1 _17668_ (.A(_08598_),
    .B(_08637_),
    .X(_08638_));
 sg13g2_nor4_1 _17669_ (.A(_08599_),
    .B(_08633_),
    .C(_08636_),
    .D(_08638_),
    .Y(_08639_));
 sg13g2_nor3_1 _17670_ (.A(net115),
    .B(_08351_),
    .C(_08639_),
    .Y(_08640_));
 sg13g2_o21ai_1 _17671_ (.B1(_08640_),
    .Y(_08641_),
    .A1(_08605_),
    .A2(_08620_));
 sg13g2_nor2_1 _17672_ (.A(_08349_),
    .B(_07602_),
    .Y(_08642_));
 sg13g2_xor2_1 _17673_ (.B(_08598_),
    .A(_08518_),
    .X(_08643_));
 sg13g2_a221oi_1 _17674_ (.B2(net111),
    .C1(net290),
    .B1(_08643_),
    .A1(_06114_),
    .Y(_08644_),
    .A2(_08642_));
 sg13g2_a21oi_1 _17675_ (.A1(_06762_),
    .A2(_08352_),
    .Y(_08645_),
    .B1(_08644_));
 sg13g2_and3_1 _17676_ (.X(_00354_),
    .A(_06667_),
    .B(_08641_),
    .C(_08645_));
 sg13g2_nand2_1 _17677_ (.Y(_08646_),
    .A(net566),
    .B(_08375_));
 sg13g2_nor2_1 _17678_ (.A(net908),
    .B(_08377_),
    .Y(_08647_));
 sg13g2_buf_1 _17679_ (.A(_00144_),
    .X(_08648_));
 sg13g2_o21ai_1 _17680_ (.B1(net1132),
    .Y(_08649_),
    .A1(_08375_),
    .A2(_08647_));
 sg13g2_a21oi_1 _17681_ (.A1(_08646_),
    .A2(_08649_),
    .Y(_08650_),
    .B1(net302));
 sg13g2_nand2b_1 _17682_ (.Y(_08651_),
    .B(_08377_),
    .A_N(net1132));
 sg13g2_nand2_1 _17683_ (.Y(_08652_),
    .A(net925),
    .B(net934));
 sg13g2_nor2_1 _17684_ (.A(_08652_),
    .B(_08377_),
    .Y(_08653_));
 sg13g2_o21ai_1 _17685_ (.B1(_08653_),
    .Y(_08654_),
    .A1(net1132),
    .A2(_08406_));
 sg13g2_a21oi_1 _17686_ (.A1(_08651_),
    .A2(_08654_),
    .Y(_08655_),
    .B1(net566));
 sg13g2_nor2b_1 _17687_ (.A(_08593_),
    .B_N(net1132),
    .Y(_08656_));
 sg13g2_nand2_1 _17688_ (.Y(_08657_),
    .A(net573),
    .B(net934));
 sg13g2_nand2_1 _17689_ (.Y(_08658_),
    .A(_08381_),
    .B(_08657_));
 sg13g2_nor2_1 _17690_ (.A(net1132),
    .B(net285),
    .Y(_08659_));
 sg13g2_a22oi_1 _17691_ (.Y(_08660_),
    .B1(_08659_),
    .B2(_08018_),
    .A2(_08658_),
    .A1(_08656_));
 sg13g2_nor2_1 _17692_ (.A(net298),
    .B(_08660_),
    .Y(_08661_));
 sg13g2_nand2_1 _17693_ (.Y(_08662_),
    .A(_08593_),
    .B(_08378_));
 sg13g2_or2_1 _17694_ (.X(_08663_),
    .B(_08662_),
    .A(_08010_));
 sg13g2_a21oi_1 _17695_ (.A1(_08646_),
    .A2(_08663_),
    .Y(_08664_),
    .B1(net297));
 sg13g2_nor4_2 _17696_ (.A(_08650_),
    .B(_08655_),
    .C(_08661_),
    .Y(_08665_),
    .D(_08664_));
 sg13g2_xnor2_1 _17697_ (.Y(_08666_),
    .A(_08592_),
    .B(net915));
 sg13g2_xnor2_1 _17698_ (.Y(_08667_),
    .A(_07980_),
    .B(_08666_));
 sg13g2_xnor2_1 _17699_ (.Y(_08668_),
    .A(net585),
    .B(_08667_));
 sg13g2_buf_1 _17700_ (.A(_08668_),
    .X(_08669_));
 sg13g2_nor2_1 _17701_ (.A(net291),
    .B(_08669_),
    .Y(_08670_));
 sg13g2_buf_1 _17702_ (.A(_00114_),
    .X(_08671_));
 sg13g2_inv_1 _17703_ (.Y(_08672_),
    .A(net1131));
 sg13g2_o21ai_1 _17704_ (.B1(_08672_),
    .Y(_08673_),
    .A1(net299),
    .A2(_08670_));
 sg13g2_nand2_1 _17705_ (.Y(_08674_),
    .A(net299),
    .B(_08670_));
 sg13g2_nand2_1 _17706_ (.Y(_08675_),
    .A(_08673_),
    .B(_08674_));
 sg13g2_xnor2_1 _17707_ (.Y(_08676_),
    .A(_08567_),
    .B(_08669_));
 sg13g2_o21ai_1 _17708_ (.B1(net289),
    .Y(_08677_),
    .A1(net170),
    .A2(_08676_));
 sg13g2_nand2b_1 _17709_ (.Y(_08678_),
    .B(_07993_),
    .A_N(net585));
 sg13g2_nand3b_1 _17710_ (.B(_08678_),
    .C(net286),
    .Y(_08679_),
    .A_N(_08324_));
 sg13g2_o21ai_1 _17711_ (.B1(_08679_),
    .Y(_08680_),
    .A1(net146),
    .A2(_08314_));
 sg13g2_o21ai_1 _17712_ (.B1(_08651_),
    .Y(_08681_),
    .A1(net303),
    .A2(_08680_));
 sg13g2_nor2_1 _17713_ (.A(net281),
    .B(_08652_),
    .Y(_08682_));
 sg13g2_a221oi_1 _17714_ (.B2(_08377_),
    .C1(_08351_),
    .B1(_08682_),
    .A1(net281),
    .Y(_08683_),
    .A2(_08681_));
 sg13g2_nand2_1 _17715_ (.Y(_08684_),
    .A(_08677_),
    .B(_08683_));
 sg13g2_a21oi_1 _17716_ (.A1(_08665_),
    .A2(_08675_),
    .Y(_08685_),
    .B1(_08684_));
 sg13g2_o21ai_1 _17717_ (.B1(_08670_),
    .Y(_08686_),
    .A1(_08672_),
    .A2(net299));
 sg13g2_nand4_1 _17718_ (.B(net1131),
    .C(_07871_),
    .A(_08292_),
    .Y(_08687_),
    .D(_08665_));
 sg13g2_nor2_1 _17719_ (.A(net1131),
    .B(_07871_),
    .Y(_08688_));
 sg13g2_nand2_1 _17720_ (.Y(_08689_),
    .A(_08292_),
    .B(net576));
 sg13g2_nand2_1 _17721_ (.Y(_08690_),
    .A(_08669_),
    .B(_08689_));
 sg13g2_o21ai_1 _17722_ (.B1(_08690_),
    .Y(_08691_),
    .A1(_08665_),
    .A2(_08688_));
 sg13g2_nor3_1 _17723_ (.A(net1131),
    .B(net291),
    .C(net586),
    .Y(_08692_));
 sg13g2_a21oi_1 _17724_ (.A1(net1131),
    .A2(_08669_),
    .Y(_08693_),
    .B1(_08692_));
 sg13g2_o21ai_1 _17725_ (.B1(_07871_),
    .Y(_08694_),
    .A1(_08293_),
    .A2(_08671_));
 sg13g2_nand3_1 _17726_ (.B(_08669_),
    .C(_08694_),
    .A(net291),
    .Y(_08695_));
 sg13g2_o21ai_1 _17727_ (.B1(_08695_),
    .Y(_08696_),
    .A1(_08292_),
    .A2(_08693_));
 sg13g2_nand2b_1 _17728_ (.Y(_08697_),
    .B(_08696_),
    .A_N(_08665_));
 sg13g2_nand4_1 _17729_ (.B(_08687_),
    .C(_08691_),
    .A(_08686_),
    .Y(_08698_),
    .D(_08697_));
 sg13g2_nor3_1 _17730_ (.A(net289),
    .B(net83),
    .C(_08351_),
    .Y(_08699_));
 sg13g2_a221oi_1 _17731_ (.B2(_08698_),
    .C1(_08699_),
    .B1(_08685_),
    .A1(net45),
    .Y(_08700_),
    .A2(net41));
 sg13g2_nor2_1 _17732_ (.A(_02970_),
    .B(_08700_),
    .Y(_00355_));
 sg13g2_and2_1 _17733_ (.A(_08378_),
    .B(net917),
    .X(_08701_));
 sg13g2_buf_1 _17734_ (.A(_08701_),
    .X(_08702_));
 sg13g2_nor2b_1 _17735_ (.A(net1132),
    .B_N(_08702_),
    .Y(_08703_));
 sg13g2_nor3_1 _17736_ (.A(net1132),
    .B(_08395_),
    .C(net288),
    .Y(_08704_));
 sg13g2_nor3_1 _17737_ (.A(_08652_),
    .B(_08702_),
    .C(_08704_),
    .Y(_08705_));
 sg13g2_o21ai_1 _17738_ (.B1(net281),
    .Y(_08706_),
    .A1(_08703_),
    .A2(_08705_));
 sg13g2_nor2_1 _17739_ (.A(net286),
    .B(net575),
    .Y(_08707_));
 sg13g2_nand2_1 _17740_ (.Y(_08708_),
    .A(net566),
    .B(_08707_));
 sg13g2_nor2_1 _17741_ (.A(net567),
    .B(_08702_),
    .Y(_08709_));
 sg13g2_o21ai_1 _17742_ (.B1(_08648_),
    .Y(_08710_),
    .A1(_08707_),
    .A2(_08709_));
 sg13g2_a21oi_1 _17743_ (.A1(_08708_),
    .A2(_08710_),
    .Y(_08711_),
    .B1(net150));
 sg13g2_o21ai_1 _17744_ (.B1(_08657_),
    .Y(_08712_),
    .A1(_08392_),
    .A2(net289));
 sg13g2_nor2_1 _17745_ (.A(net1132),
    .B(net303),
    .Y(_08713_));
 sg13g2_a22oi_1 _17746_ (.Y(_08714_),
    .B1(_08713_),
    .B2(_08702_),
    .A2(_08712_),
    .A1(_08656_));
 sg13g2_nor2_1 _17747_ (.A(net298),
    .B(_08714_),
    .Y(_08715_));
 sg13g2_nand4_1 _17748_ (.B(_08395_),
    .C(net288),
    .A(net567),
    .Y(_08716_),
    .D(net302));
 sg13g2_a21oi_1 _17749_ (.A1(_08708_),
    .A2(_08716_),
    .Y(_08717_),
    .B1(net149));
 sg13g2_nor3_1 _17750_ (.A(_08711_),
    .B(_08715_),
    .C(_08717_),
    .Y(_08718_));
 sg13g2_nand2_1 _17751_ (.Y(_08719_),
    .A(_08706_),
    .B(_08718_));
 sg13g2_xnor2_1 _17752_ (.Y(_08720_),
    .A(_08595_),
    .B(_08666_));
 sg13g2_xnor2_1 _17753_ (.Y(_08721_),
    .A(net303),
    .B(_08720_));
 sg13g2_xnor2_1 _17754_ (.Y(_08722_),
    .A(_08036_),
    .B(_08721_));
 sg13g2_o21ai_1 _17755_ (.B1(_08439_),
    .Y(_08723_),
    .A1(net1142),
    .A2(_08721_));
 sg13g2_a21oi_1 _17756_ (.A1(_08437_),
    .A2(_08722_),
    .Y(_08724_),
    .B1(_08723_));
 sg13g2_xor2_1 _17757_ (.B(_08724_),
    .A(_08719_),
    .X(_08725_));
 sg13g2_nand3_1 _17758_ (.B(net288),
    .C(net297),
    .A(_08402_),
    .Y(_08726_));
 sg13g2_o21ai_1 _17759_ (.B1(_08726_),
    .Y(_08727_),
    .A1(_08402_),
    .A2(_08595_));
 sg13g2_a21oi_1 _17760_ (.A1(net150),
    .A2(_08727_),
    .Y(_08728_),
    .B1(_08703_));
 sg13g2_a21oi_1 _17761_ (.A1(_07908_),
    .A2(_08702_),
    .Y(_08729_),
    .B1(net281));
 sg13g2_a21oi_1 _17762_ (.A1(net281),
    .A2(_08728_),
    .Y(_08730_),
    .B1(_08729_));
 sg13g2_nor4_1 _17763_ (.A(_08355_),
    .B(net1142),
    .C(_08420_),
    .D(_08721_),
    .Y(_08731_));
 sg13g2_xnor2_1 _17764_ (.Y(_08732_),
    .A(_08462_),
    .B(_08721_));
 sg13g2_nor2_1 _17765_ (.A(net147),
    .B(_08732_),
    .Y(_08733_));
 sg13g2_nor4_1 _17766_ (.A(net99),
    .B(_08730_),
    .C(_08731_),
    .D(_08733_),
    .Y(_08734_));
 sg13g2_nand2_1 _17767_ (.Y(_08735_),
    .A(_08725_),
    .B(_08734_));
 sg13g2_a22oi_1 _17768_ (.Y(_08736_),
    .B1(net76),
    .B2(_08642_),
    .A2(net71),
    .A1(net147));
 sg13g2_a221oi_1 _17769_ (.B2(_08736_),
    .C1(net617),
    .B1(_08735_),
    .A1(_06471_),
    .Y(_00356_),
    .A2(_08642_));
 sg13g2_buf_2 _17770_ (.A(net110),
    .X(_08737_));
 sg13g2_nand2_1 _17771_ (.Y(_08738_),
    .A(net584),
    .B(net147));
 sg13g2_buf_2 _17772_ (.A(\grid.cell_19_0.se ),
    .X(_08739_));
 sg13g2_inv_1 _17773_ (.Y(_08740_),
    .A(_08739_));
 sg13g2_buf_1 _17774_ (.A(_08740_),
    .X(_08741_));
 sg13g2_buf_2 _17775_ (.A(\grid.cell_19_0.sw ),
    .X(_08742_));
 sg13g2_xnor2_1 _17776_ (.Y(_08743_),
    .A(_08742_),
    .B(_08358_));
 sg13g2_buf_2 _17777_ (.A(_08743_),
    .X(_08744_));
 sg13g2_xnor2_1 _17778_ (.Y(_08745_),
    .A(net565),
    .B(_08744_));
 sg13g2_nor2_1 _17779_ (.A(net1143),
    .B(_08313_),
    .Y(_08746_));
 sg13g2_nor3_1 _17780_ (.A(_08114_),
    .B(_08745_),
    .C(_08746_),
    .Y(_08747_));
 sg13g2_a21oi_1 _17781_ (.A1(_08738_),
    .A2(_08745_),
    .Y(_08748_),
    .B1(_08747_));
 sg13g2_buf_1 _17782_ (.A(_08742_),
    .X(_08749_));
 sg13g2_buf_1 _17783_ (.A(net907),
    .X(_08750_));
 sg13g2_nand2b_1 _17784_ (.Y(_08751_),
    .B(net915),
    .A_N(_08108_));
 sg13g2_nor2b_1 _17785_ (.A(_08742_),
    .B_N(_08358_),
    .Y(_08752_));
 sg13g2_a21oi_1 _17786_ (.A1(net564),
    .A2(_08751_),
    .Y(_08753_),
    .B1(_08752_));
 sg13g2_nor2_1 _17787_ (.A(net295),
    .B(_08753_),
    .Y(_08754_));
 sg13g2_nand2b_1 _17788_ (.Y(_08755_),
    .B(_08742_),
    .A_N(_08358_));
 sg13g2_nand2b_1 _17789_ (.Y(_08756_),
    .B(net583),
    .A_N(_08750_));
 sg13g2_a21oi_1 _17790_ (.A1(_08755_),
    .A2(_08756_),
    .Y(_08757_),
    .B1(net1143));
 sg13g2_or2_1 _17791_ (.X(_08758_),
    .B(net915),
    .A(net907));
 sg13g2_buf_1 _17792_ (.A(_08758_),
    .X(_08759_));
 sg13g2_nor2_1 _17793_ (.A(_08108_),
    .B(_08759_),
    .Y(_08760_));
 sg13g2_nor4_1 _17794_ (.A(net565),
    .B(_08754_),
    .C(_08757_),
    .D(_08760_),
    .Y(_08761_));
 sg13g2_o21ai_1 _17795_ (.B1(_08379_),
    .Y(_08762_),
    .A1(net573),
    .A2(_08108_));
 sg13g2_buf_1 _17796_ (.A(net907),
    .X(_08763_));
 sg13g2_nor2_1 _17797_ (.A(net563),
    .B(_08751_),
    .Y(_08764_));
 sg13g2_a221oi_1 _17798_ (.B2(net563),
    .C1(_08764_),
    .B1(_08762_),
    .A1(_08746_),
    .Y(_08765_),
    .A2(_08759_));
 sg13g2_and2_1 _17799_ (.A(net565),
    .B(_08765_),
    .X(_08766_));
 sg13g2_buf_1 _17800_ (.A(_08739_),
    .X(_08767_));
 sg13g2_buf_1 _17801_ (.A(_08750_),
    .X(_08768_));
 sg13g2_nor3_1 _17802_ (.A(net906),
    .B(net279),
    .C(_08381_),
    .Y(_08769_));
 sg13g2_nand2_1 _17803_ (.Y(_08770_),
    .A(net563),
    .B(net573));
 sg13g2_nor3_1 _17804_ (.A(_08740_),
    .B(_08114_),
    .C(_08770_),
    .Y(_08771_));
 sg13g2_o21ai_1 _17805_ (.B1(net924),
    .Y(_08772_),
    .A1(_08769_),
    .A2(_08771_));
 sg13g2_o21ai_1 _17806_ (.B1(_08772_),
    .Y(_08773_),
    .A1(_08761_),
    .A2(_08766_));
 sg13g2_buf_1 _17807_ (.A(_00209_),
    .X(_08774_));
 sg13g2_buf_1 _17808_ (.A(_08774_),
    .X(_08775_));
 sg13g2_nor4_1 _17809_ (.A(net922),
    .B(net574),
    .C(net905),
    .D(_08744_),
    .Y(_08776_));
 sg13g2_nand3b_1 _17810_ (.B(net914),
    .C(net922),
    .Y(_08777_),
    .A_N(_08774_));
 sg13g2_nor2_1 _17811_ (.A(_08744_),
    .B(_08777_),
    .Y(_08778_));
 sg13g2_xor2_1 _17812_ (.B(_08739_),
    .A(net1143),
    .X(_08779_));
 sg13g2_xnor2_1 _17813_ (.Y(_08780_),
    .A(net295),
    .B(_08779_));
 sg13g2_o21ai_1 _17814_ (.B1(_08780_),
    .Y(_08781_),
    .A1(_08776_),
    .A2(_08778_));
 sg13g2_nand2b_1 _17815_ (.Y(_08782_),
    .B(_08755_),
    .A_N(_08752_));
 sg13g2_buf_1 _17816_ (.A(_08782_),
    .X(_08783_));
 sg13g2_nand2_1 _17817_ (.Y(_08784_),
    .A(net922),
    .B(_08391_));
 sg13g2_nor3_1 _17818_ (.A(_08775_),
    .B(_08783_),
    .C(_08784_),
    .Y(_08785_));
 sg13g2_inv_1 _17819_ (.Y(_08786_),
    .A(_08034_));
 sg13g2_nand2_1 _17820_ (.Y(_08787_),
    .A(_08786_),
    .B(net914));
 sg13g2_nor3_1 _17821_ (.A(net905),
    .B(_08783_),
    .C(_08787_),
    .Y(_08788_));
 sg13g2_o21ai_1 _17822_ (.B1(_08780_),
    .Y(_08789_),
    .A1(_08785_),
    .A2(_08788_));
 sg13g2_nor3_1 _17823_ (.A(_08775_),
    .B(_08744_),
    .C(_08784_),
    .Y(_08790_));
 sg13g2_nor3_1 _17824_ (.A(net905),
    .B(_08744_),
    .C(_08787_),
    .Y(_08791_));
 sg13g2_xnor2_1 _17825_ (.Y(_08792_),
    .A(_08313_),
    .B(_08779_));
 sg13g2_o21ai_1 _17826_ (.B1(_08792_),
    .Y(_08793_),
    .A1(_08790_),
    .A2(_08791_));
 sg13g2_nor4_1 _17827_ (.A(net922),
    .B(net914),
    .C(_08774_),
    .D(_08783_),
    .Y(_08794_));
 sg13g2_nor2_1 _17828_ (.A(_08783_),
    .B(_08777_),
    .Y(_08795_));
 sg13g2_o21ai_1 _17829_ (.B1(_08792_),
    .Y(_08796_),
    .A1(_08794_),
    .A2(_08795_));
 sg13g2_nand4_1 _17830_ (.B(_08789_),
    .C(_08793_),
    .A(_08781_),
    .Y(_08797_),
    .D(_08796_));
 sg13g2_xor2_1 _17831_ (.B(_08797_),
    .A(_08773_),
    .X(_08798_));
 sg13g2_xnor2_1 _17832_ (.Y(_08799_),
    .A(_08783_),
    .B(_08792_));
 sg13g2_xnor2_1 _17833_ (.Y(_08800_),
    .A(net574),
    .B(_08799_));
 sg13g2_nor2_1 _17834_ (.A(_08482_),
    .B(_08799_),
    .Y(_08801_));
 sg13g2_a21oi_1 _17835_ (.A1(net582),
    .A2(_08800_),
    .Y(_08802_),
    .B1(_08801_));
 sg13g2_buf_1 _17836_ (.A(net906),
    .X(_08803_));
 sg13g2_and2_1 _17837_ (.A(net907),
    .B(net573),
    .X(_08804_));
 sg13g2_buf_1 _17838_ (.A(_08804_),
    .X(_08805_));
 sg13g2_a21o_1 _17839_ (.A2(_08759_),
    .A1(net562),
    .B1(_08805_),
    .X(_08806_));
 sg13g2_nor4_1 _17840_ (.A(_08748_),
    .B(_08798_),
    .C(_08802_),
    .D(_08806_),
    .Y(_08807_));
 sg13g2_nand2_1 _17841_ (.Y(_08808_),
    .A(_08748_),
    .B(_08806_));
 sg13g2_and3_1 _17842_ (.X(_08809_),
    .A(_08798_),
    .B(_08802_),
    .C(_08808_));
 sg13g2_nor3_1 _17843_ (.A(net69),
    .B(_08807_),
    .C(_08809_),
    .Y(_08810_));
 sg13g2_buf_1 _17844_ (.A(\grid.cell_19_0.s ),
    .X(_08811_));
 sg13g2_buf_1 _17845_ (.A(_08811_),
    .X(_08812_));
 sg13g2_xnor2_1 _17846_ (.Y(_08813_),
    .A(_08786_),
    .B(_08800_));
 sg13g2_xnor2_1 _17847_ (.Y(_08814_),
    .A(net904),
    .B(_08813_));
 sg13g2_nor2_1 _17848_ (.A(net103),
    .B(_08814_),
    .Y(_08815_));
 sg13g2_nand2_1 _17849_ (.Y(_08816_),
    .A(_05175_),
    .B(_05748_));
 sg13g2_buf_2 _17850_ (.A(_08816_),
    .X(_08817_));
 sg13g2_nor2_1 _17851_ (.A(_07602_),
    .B(_08817_),
    .Y(_08818_));
 sg13g2_nor2_2 _17852_ (.A(_00648_),
    .B(_08818_),
    .Y(_08819_));
 sg13g2_o21ai_1 _17853_ (.B1(_08819_),
    .Y(_08820_),
    .A1(net572),
    .A2(_08815_));
 sg13g2_buf_1 _17854_ (.A(_08818_),
    .X(_08821_));
 sg13g2_nand3_1 _17855_ (.B(net44),
    .C(net58),
    .A(net637),
    .Y(_08822_));
 sg13g2_o21ai_1 _17856_ (.B1(_08822_),
    .Y(_00357_),
    .A1(_08810_),
    .A2(_08820_));
 sg13g2_buf_2 _17857_ (.A(\grid.cell_19_1.se ),
    .X(_08823_));
 sg13g2_buf_1 _17858_ (.A(_08823_),
    .X(_08824_));
 sg13g2_nand2_1 _17859_ (.Y(_08825_),
    .A(net912),
    .B(net903));
 sg13g2_xor2_1 _17860_ (.B(_08823_),
    .A(net1137),
    .X(_08826_));
 sg13g2_buf_2 _17861_ (.A(_08826_),
    .X(_08827_));
 sg13g2_nand2_1 _17862_ (.Y(_08828_),
    .A(net924),
    .B(_08827_));
 sg13g2_o21ai_1 _17863_ (.B1(_08828_),
    .Y(_08829_),
    .A1(net924),
    .A2(_08825_));
 sg13g2_nand2_1 _17864_ (.Y(_08830_),
    .A(net294),
    .B(_08829_));
 sg13g2_o21ai_1 _17865_ (.B1(_08830_),
    .Y(_08831_),
    .A1(_08108_),
    .A2(_08825_));
 sg13g2_nor2_1 _17866_ (.A(net562),
    .B(_08046_),
    .Y(_08832_));
 sg13g2_nor2_1 _17867_ (.A(net912),
    .B(_08824_),
    .Y(_08833_));
 sg13g2_a21oi_1 _17868_ (.A1(_08832_),
    .A2(_08833_),
    .Y(_08834_),
    .B1(net916));
 sg13g2_xor2_1 _17869_ (.B(net581),
    .A(net906),
    .X(_08835_));
 sg13g2_nand3_1 _17870_ (.B(_08767_),
    .C(net580),
    .A(_07987_),
    .Y(_08836_));
 sg13g2_o21ai_1 _17871_ (.B1(_08836_),
    .Y(_08837_),
    .A1(net584),
    .A2(_08835_));
 sg13g2_xnor2_1 _17872_ (.Y(_08838_),
    .A(_08741_),
    .B(_08070_));
 sg13g2_nand2_1 _17873_ (.Y(_08839_),
    .A(_08827_),
    .B(_08838_));
 sg13g2_o21ai_1 _17874_ (.B1(_08839_),
    .Y(_08840_),
    .A1(_08827_),
    .A2(_08837_));
 sg13g2_nor3_1 _17875_ (.A(_08803_),
    .B(_08046_),
    .C(_08825_),
    .Y(_08841_));
 sg13g2_a221oi_1 _17876_ (.B2(_08840_),
    .C1(_08841_),
    .B1(_08834_),
    .A1(_08803_),
    .Y(_08842_),
    .A2(_08831_));
 sg13g2_buf_1 _17877_ (.A(net905),
    .X(_08843_));
 sg13g2_inv_2 _17878_ (.Y(_08844_),
    .A(_08823_));
 sg13g2_xnor2_1 _17879_ (.Y(_08845_),
    .A(_08844_),
    .B(_08431_));
 sg13g2_xor2_1 _17880_ (.B(_08845_),
    .A(_08779_),
    .X(_08846_));
 sg13g2_buf_2 _17881_ (.A(_08846_),
    .X(_08847_));
 sg13g2_xnor2_1 _17882_ (.Y(_08848_),
    .A(net913),
    .B(_08847_));
 sg13g2_o21ai_1 _17883_ (.B1(_08786_),
    .Y(_08849_),
    .A1(net561),
    .A2(_08848_));
 sg13g2_nand2_1 _17884_ (.Y(_08850_),
    .A(net561),
    .B(_08848_));
 sg13g2_nand2_1 _17885_ (.Y(_08851_),
    .A(_08849_),
    .B(_08850_));
 sg13g2_a22oi_1 _17886_ (.Y(_08852_),
    .B1(_08827_),
    .B2(net924),
    .A2(_08825_),
    .A1(net580));
 sg13g2_nand2_1 _17887_ (.Y(_08853_),
    .A(_08046_),
    .B(_08833_));
 sg13g2_o21ai_1 _17888_ (.B1(_08853_),
    .Y(_08854_),
    .A1(_08114_),
    .A2(_08852_));
 sg13g2_buf_1 _17889_ (.A(net903),
    .X(_08855_));
 sg13g2_a21oi_1 _17890_ (.A1(net924),
    .A2(_08767_),
    .Y(_08856_),
    .B1(net580));
 sg13g2_nor4_1 _17891_ (.A(net571),
    .B(_08855_),
    .C(_08114_),
    .D(_08856_),
    .Y(_08857_));
 sg13g2_a21oi_1 _17892_ (.A1(_08741_),
    .A2(_08854_),
    .Y(_08858_),
    .B1(_08857_));
 sg13g2_nand2_1 _17893_ (.Y(_08859_),
    .A(net127),
    .B(_08858_));
 sg13g2_a21oi_1 _17894_ (.A1(_08842_),
    .A2(_08851_),
    .Y(_08860_),
    .B1(_08859_));
 sg13g2_xnor2_1 _17895_ (.Y(_08861_),
    .A(_08413_),
    .B(_08811_));
 sg13g2_xnor2_1 _17896_ (.Y(_08862_),
    .A(net922),
    .B(_08861_));
 sg13g2_xor2_1 _17897_ (.B(_08862_),
    .A(_08847_),
    .X(_08863_));
 sg13g2_a21oi_1 _17898_ (.A1(net70),
    .A2(_08863_),
    .Y(_08864_),
    .B1(net287));
 sg13g2_o21ai_1 _17899_ (.B1(_08847_),
    .Y(_08865_),
    .A1(net582),
    .A2(net1138));
 sg13g2_nand2_1 _17900_ (.Y(_08866_),
    .A(net572),
    .B(_08865_));
 sg13g2_nand2b_1 _17901_ (.Y(_08867_),
    .B(net572),
    .A_N(net1138));
 sg13g2_nor2b_1 _17902_ (.A(net572),
    .B_N(net1138),
    .Y(_08868_));
 sg13g2_a22oi_1 _17903_ (.Y(_08869_),
    .B1(_08868_),
    .B2(_08847_),
    .A2(_08867_),
    .A1(net582));
 sg13g2_a21oi_1 _17904_ (.A1(_08866_),
    .A2(_08869_),
    .Y(_08870_),
    .B1(net561));
 sg13g2_nand3b_1 _17905_ (.B(_08847_),
    .C(net561),
    .Y(_08871_),
    .A_N(net916));
 sg13g2_o21ai_1 _17906_ (.B1(_08871_),
    .Y(_08872_),
    .A1(_08786_),
    .A2(_08848_));
 sg13g2_nor4_1 _17907_ (.A(net120),
    .B(_08858_),
    .C(_08870_),
    .D(_08872_),
    .Y(_08873_));
 sg13g2_nor3_1 _17908_ (.A(_08860_),
    .B(_08864_),
    .C(_08873_),
    .Y(_08874_));
 sg13g2_and3_1 _17909_ (.X(_08875_),
    .A(net716),
    .B(_03153_),
    .C(net58));
 sg13g2_a21o_1 _17910_ (.A2(_08874_),
    .A1(_08819_),
    .B1(_08875_),
    .X(_00358_));
 sg13g2_nor2_1 _17911_ (.A(_00648_),
    .B(_02765_),
    .Y(_08876_));
 sg13g2_buf_2 _17912_ (.A(_08876_),
    .X(_08877_));
 sg13g2_or2_1 _17913_ (.X(_08878_),
    .B(_08817_),
    .A(_07602_));
 sg13g2_buf_1 _17914_ (.A(_08878_),
    .X(_08879_));
 sg13g2_buf_1 _17915_ (.A(\grid.cell_19_2.se ),
    .X(_08880_));
 sg13g2_buf_1 _17916_ (.A(_08880_),
    .X(_08881_));
 sg13g2_xnor2_1 _17917_ (.Y(_08882_),
    .A(_08371_),
    .B(net902));
 sg13g2_xnor2_1 _17918_ (.Y(_08883_),
    .A(_08044_),
    .B(net903));
 sg13g2_xnor2_1 _17919_ (.Y(_08884_),
    .A(_08882_),
    .B(_08883_));
 sg13g2_xnor2_1 _17920_ (.Y(_08885_),
    .A(_08472_),
    .B(_08884_));
 sg13g2_buf_1 _17921_ (.A(_08885_),
    .X(_08886_));
 sg13g2_xor2_1 _17922_ (.B(_08886_),
    .A(_08779_),
    .X(_08887_));
 sg13g2_o21ai_1 _17923_ (.B1(_08422_),
    .Y(_08888_),
    .A1(net125),
    .A2(_08887_));
 sg13g2_nand3_1 _17924_ (.B(_08879_),
    .C(_08888_),
    .A(_08877_),
    .Y(_08889_));
 sg13g2_nand3_1 _17925_ (.B(net33),
    .C(net58),
    .A(net637),
    .Y(_08890_));
 sg13g2_buf_1 _17926_ (.A(_08855_),
    .X(_08891_));
 sg13g2_buf_1 _17927_ (.A(net902),
    .X(_08892_));
 sg13g2_nor2_1 _17928_ (.A(net559),
    .B(net570),
    .Y(_08893_));
 sg13g2_nand2_1 _17929_ (.Y(_08894_),
    .A(net581),
    .B(net920));
 sg13g2_nand2_1 _17930_ (.Y(_08895_),
    .A(net902),
    .B(net911));
 sg13g2_inv_1 _17931_ (.Y(_08896_),
    .A(_08895_));
 sg13g2_xor2_1 _17932_ (.B(_08468_),
    .A(_08880_),
    .X(_08897_));
 sg13g2_nand2_1 _17933_ (.Y(_08898_),
    .A(net921),
    .B(_08897_));
 sg13g2_o21ai_1 _17934_ (.B1(_08898_),
    .Y(_08899_),
    .A1(net579),
    .A2(_08896_));
 sg13g2_a22oi_1 _17935_ (.Y(_08900_),
    .B1(_08899_),
    .B2(_08137_),
    .A2(_08894_),
    .A1(_08893_));
 sg13g2_o21ai_1 _17936_ (.B1(net579),
    .Y(_08901_),
    .A1(net580),
    .A2(_08844_));
 sg13g2_nand3_1 _17937_ (.B(_08901_),
    .C(_08893_),
    .A(_08137_),
    .Y(_08902_));
 sg13g2_o21ai_1 _17938_ (.B1(_08902_),
    .Y(_08903_),
    .A1(_08891_),
    .A2(_08900_));
 sg13g2_xnor2_1 _17939_ (.Y(_08904_),
    .A(_08165_),
    .B(_08897_));
 sg13g2_xor2_1 _17940_ (.B(_08904_),
    .A(_08883_),
    .X(_08905_));
 sg13g2_nor2_1 _17941_ (.A(_08482_),
    .B(_08905_),
    .Y(_08906_));
 sg13g2_buf_1 _17942_ (.A(_00208_),
    .X(_08907_));
 sg13g2_buf_1 _17943_ (.A(_08907_),
    .X(_08908_));
 sg13g2_a21o_1 _17944_ (.A2(_08886_),
    .A1(_08009_),
    .B1(net901),
    .X(_08909_));
 sg13g2_o21ai_1 _17945_ (.B1(_08886_),
    .Y(_08910_),
    .A1(net901),
    .A2(_08906_));
 sg13g2_nor3_1 _17946_ (.A(net901),
    .B(_08886_),
    .C(_08906_),
    .Y(_08911_));
 sg13g2_a221oi_1 _17947_ (.B2(net584),
    .C1(_08911_),
    .B1(_08910_),
    .A1(_08906_),
    .Y(_08912_),
    .A2(_08909_));
 sg13g2_o21ai_1 _17948_ (.B1(_08009_),
    .Y(_08913_),
    .A1(net901),
    .A2(_08886_));
 sg13g2_nand2_1 _17949_ (.Y(_08914_),
    .A(net901),
    .B(_08886_));
 sg13g2_a21oi_1 _17950_ (.A1(_08913_),
    .A2(_08914_),
    .Y(_08915_),
    .B1(_08906_));
 sg13g2_nor2_1 _17951_ (.A(_08903_),
    .B(_08915_),
    .Y(_08916_));
 sg13g2_a21oi_1 _17952_ (.A1(_08903_),
    .A2(_08912_),
    .Y(_08917_),
    .B1(_08916_));
 sg13g2_o21ai_1 _17953_ (.B1(_08898_),
    .Y(_08918_),
    .A1(net294),
    .A2(_08895_));
 sg13g2_nand2_1 _17954_ (.Y(_08919_),
    .A(net293),
    .B(_08918_));
 sg13g2_o21ai_1 _17955_ (.B1(_08919_),
    .Y(_08920_),
    .A1(_08137_),
    .A2(_08895_));
 sg13g2_nor2_1 _17956_ (.A(net278),
    .B(_08894_),
    .Y(_08921_));
 sg13g2_a22oi_1 _17957_ (.Y(_08922_),
    .B1(_08921_),
    .B2(_08896_),
    .A2(_08920_),
    .A1(net278));
 sg13g2_nand4_1 _17958_ (.B(_08888_),
    .C(_08917_),
    .A(_08819_),
    .Y(_08923_),
    .D(_08922_));
 sg13g2_nand3_1 _17959_ (.B(_08890_),
    .C(_08923_),
    .A(_08889_),
    .Y(_00359_));
 sg13g2_buf_1 _17960_ (.A(\grid.cell_19_3.se ),
    .X(_08924_));
 sg13g2_buf_1 _17961_ (.A(_08924_),
    .X(_08925_));
 sg13g2_buf_1 _17962_ (.A(net900),
    .X(_08926_));
 sg13g2_buf_1 _17963_ (.A(net558),
    .X(_08927_));
 sg13g2_buf_1 _17964_ (.A(net559),
    .X(_08928_));
 sg13g2_nand4_1 _17965_ (.B(net283),
    .C(net292),
    .A(net276),
    .Y(_08929_),
    .D(net293));
 sg13g2_o21ai_1 _17966_ (.B1(_08819_),
    .Y(_08930_),
    .A1(net277),
    .A2(_08929_));
 sg13g2_buf_2 _17967_ (.A(_00207_),
    .X(_08931_));
 sg13g2_xnor2_1 _17968_ (.Y(_08932_),
    .A(_08924_),
    .B(_08504_));
 sg13g2_xnor2_1 _17969_ (.Y(_08933_),
    .A(_08133_),
    .B(_08932_));
 sg13g2_xnor2_1 _17970_ (.Y(_08934_),
    .A(_08881_),
    .B(_08933_));
 sg13g2_nand2_1 _17971_ (.Y(_08935_),
    .A(_08525_),
    .B(_08934_));
 sg13g2_nor3_1 _17972_ (.A(_08931_),
    .B(_08431_),
    .C(_08935_),
    .Y(_08936_));
 sg13g2_xnor2_1 _17973_ (.Y(_08937_),
    .A(net559),
    .B(net569));
 sg13g2_a21oi_1 _17974_ (.A1(net276),
    .A2(net569),
    .Y(_08938_),
    .B1(net579));
 sg13g2_a21oi_1 _17975_ (.A1(net293),
    .A2(_08937_),
    .Y(_08939_),
    .B1(_08938_));
 sg13g2_nand2_1 _17976_ (.Y(_08940_),
    .A(net292),
    .B(_08939_));
 sg13g2_nand3_1 _17977_ (.B(_08928_),
    .C(net283),
    .A(_08210_),
    .Y(_08941_));
 sg13g2_inv_1 _17978_ (.Y(_08942_),
    .A(_08925_));
 sg13g2_a21oi_1 _17979_ (.A1(_08940_),
    .A2(_08941_),
    .Y(_08943_),
    .B1(_08942_));
 sg13g2_xor2_1 _17980_ (.B(_08934_),
    .A(_08845_),
    .X(_08944_));
 sg13g2_a21oi_1 _17981_ (.A1(net119),
    .A2(_08944_),
    .Y(_08945_),
    .B1(net284));
 sg13g2_nor4_1 _17982_ (.A(_08930_),
    .B(_08936_),
    .C(_08943_),
    .D(_08945_),
    .Y(_08946_));
 sg13g2_nor2_1 _17983_ (.A(net577),
    .B(net579),
    .Y(_08947_));
 sg13g2_nor4_1 _17984_ (.A(net558),
    .B(net559),
    .C(net569),
    .D(net577),
    .Y(_08948_));
 sg13g2_o21ai_1 _17985_ (.B1(net569),
    .Y(_08949_),
    .A1(net558),
    .A2(_08892_));
 sg13g2_inv_1 _17986_ (.Y(_08950_),
    .A(_08949_));
 sg13g2_and2_1 _17987_ (.A(_08924_),
    .B(_08880_),
    .X(_08951_));
 sg13g2_buf_1 _17988_ (.A(_08951_),
    .X(_08952_));
 sg13g2_nor4_1 _17989_ (.A(_08947_),
    .B(_08948_),
    .C(_08950_),
    .D(_08952_),
    .Y(_08953_));
 sg13g2_nor3_1 _17990_ (.A(net277),
    .B(_08928_),
    .C(net283),
    .Y(_08954_));
 sg13g2_nand2_1 _17991_ (.Y(_08955_),
    .A(net292),
    .B(net293));
 sg13g2_a22oi_1 _17992_ (.Y(_08956_),
    .B1(_08954_),
    .B2(_08955_),
    .A2(_08953_),
    .A1(_08178_));
 sg13g2_xnor2_1 _17993_ (.Y(_08957_),
    .A(net571),
    .B(_08934_));
 sg13g2_a21oi_1 _17994_ (.A1(net580),
    .A2(_08931_),
    .Y(_08958_),
    .B1(_08957_));
 sg13g2_o21ai_1 _17995_ (.B1(_08935_),
    .Y(_08959_),
    .A1(net580),
    .A2(_08931_));
 sg13g2_nor2_1 _17996_ (.A(_08958_),
    .B(_08959_),
    .Y(_08960_));
 sg13g2_xnor2_1 _17997_ (.Y(_08961_),
    .A(_08956_),
    .B(_08960_));
 sg13g2_nand3_1 _17998_ (.B(net102),
    .C(_08879_),
    .A(net284),
    .Y(_08962_));
 sg13g2_o21ai_1 _17999_ (.B1(_08962_),
    .Y(_08963_),
    .A1(net48),
    .A2(_08879_));
 sg13g2_a22oi_1 _18000_ (.Y(_08964_),
    .B1(_08963_),
    .B2(_06900_),
    .A2(_08961_),
    .A1(_08946_));
 sg13g2_inv_1 _18001_ (.Y(_00360_),
    .A(_08964_));
 sg13g2_buf_1 _18002_ (.A(_06110_),
    .X(_08965_));
 sg13g2_buf_2 _18003_ (.A(\grid.cell_19_4.se ),
    .X(_08966_));
 sg13g2_xor2_1 _18004_ (.B(net1136),
    .A(net1129),
    .X(_08967_));
 sg13g2_xnor2_1 _18005_ (.Y(_08968_),
    .A(net900),
    .B(_08180_));
 sg13g2_xnor2_1 _18006_ (.Y(_08969_),
    .A(_08967_),
    .B(_08968_));
 sg13g2_buf_1 _18007_ (.A(_08969_),
    .X(_08970_));
 sg13g2_xnor2_1 _18008_ (.Y(_08971_),
    .A(_08904_),
    .B(_08970_));
 sg13g2_a21oi_1 _18009_ (.A1(net116),
    .A2(_08971_),
    .Y(_08972_),
    .B1(net283));
 sg13g2_nor2_1 _18010_ (.A(net58),
    .B(_08972_),
    .Y(_08973_));
 sg13g2_a21oi_1 _18011_ (.A1(_07426_),
    .A2(_08821_),
    .Y(_08974_),
    .B1(_08973_));
 sg13g2_buf_2 _18012_ (.A(_00053_),
    .X(_08975_));
 sg13g2_o21ai_1 _18013_ (.B1(_08165_),
    .Y(_08976_),
    .A1(net284),
    .A2(_08970_));
 sg13g2_nor2_1 _18014_ (.A(net1135),
    .B(net579),
    .Y(_08977_));
 sg13g2_nor3_1 _18015_ (.A(_08470_),
    .B(_08970_),
    .C(_08977_),
    .Y(_08978_));
 sg13g2_nor2_1 _18016_ (.A(_08477_),
    .B(_08978_),
    .Y(_08979_));
 sg13g2_a21oi_1 _18017_ (.A1(net1135),
    .A2(_08976_),
    .Y(_08980_),
    .B1(_08979_));
 sg13g2_xnor2_1 _18018_ (.Y(_08981_),
    .A(net284),
    .B(_08970_));
 sg13g2_nor2_1 _18019_ (.A(_08563_),
    .B(_08970_),
    .Y(_08982_));
 sg13g2_a22oi_1 _18020_ (.Y(_08983_),
    .B1(_08982_),
    .B2(_08975_),
    .A2(_08981_),
    .A1(net293));
 sg13g2_o21ai_1 _18021_ (.B1(_08983_),
    .Y(_08984_),
    .A1(_08975_),
    .A2(_08980_));
 sg13g2_inv_1 _18022_ (.Y(_08985_),
    .A(net1129));
 sg13g2_nor2_2 _18023_ (.A(net558),
    .B(_08555_),
    .Y(_08986_));
 sg13g2_nand2_1 _18024_ (.Y(_08987_),
    .A(_08985_),
    .B(_08986_));
 sg13g2_nand3_1 _18025_ (.B(net290),
    .C(_08986_),
    .A(_08985_),
    .Y(_08988_));
 sg13g2_buf_1 _18026_ (.A(net1129),
    .X(_08989_));
 sg13g2_buf_1 _18027_ (.A(_08989_),
    .X(_08990_));
 sg13g2_o21ai_1 _18028_ (.B1(net568),
    .Y(_08991_),
    .A1(net556),
    .A2(net277));
 sg13g2_a22oi_1 _18029_ (.Y(_08992_),
    .B1(net290),
    .B2(net577),
    .A2(net277),
    .A1(net556));
 sg13g2_nand4_1 _18030_ (.B(_08988_),
    .C(_08991_),
    .A(net1140),
    .Y(_08993_),
    .D(_08992_));
 sg13g2_o21ai_1 _18031_ (.B1(_08993_),
    .Y(_08994_),
    .A1(_08201_),
    .A2(_08987_));
 sg13g2_nand2_1 _18032_ (.Y(_08995_),
    .A(net577),
    .B(_08986_));
 sg13g2_nand2_1 _18033_ (.Y(_08996_),
    .A(_08926_),
    .B(net576));
 sg13g2_o21ai_1 _18034_ (.B1(_08996_),
    .Y(_08997_),
    .A1(net277),
    .A2(_08611_));
 sg13g2_nand3_1 _18035_ (.B(net292),
    .C(_08997_),
    .A(net1140),
    .Y(_08998_));
 sg13g2_a21oi_1 _18036_ (.A1(_08995_),
    .A2(_08998_),
    .Y(_08999_),
    .B1(net556));
 sg13g2_nand3_1 _18037_ (.B(net277),
    .C(net568),
    .A(net1140),
    .Y(_09000_));
 sg13g2_nand2_1 _18038_ (.Y(_09001_),
    .A(_08926_),
    .B(_08555_));
 sg13g2_nand2_1 _18039_ (.Y(_09002_),
    .A(net576),
    .B(net578));
 sg13g2_a22oi_1 _18040_ (.Y(_09003_),
    .B1(_09001_),
    .B2(_09002_),
    .A2(_08986_),
    .A1(_08249_));
 sg13g2_nand3_1 _18041_ (.B(_09000_),
    .C(_09003_),
    .A(net556),
    .Y(_09004_));
 sg13g2_buf_1 _18042_ (.A(net1129),
    .X(_09005_));
 sg13g2_nand2_1 _18043_ (.Y(_09006_),
    .A(net898),
    .B(_08163_));
 sg13g2_o21ai_1 _18044_ (.B1(_09006_),
    .Y(_09007_),
    .A1(net1140),
    .A2(net577));
 sg13g2_nand4_1 _18045_ (.B(_08575_),
    .C(net290),
    .A(_08927_),
    .Y(_09008_),
    .D(_09007_));
 sg13g2_inv_1 _18046_ (.Y(_09009_),
    .A(_08975_));
 sg13g2_nand2_1 _18047_ (.Y(_09010_),
    .A(_09009_),
    .B(net293));
 sg13g2_nand3_1 _18048_ (.B(_09008_),
    .C(_09010_),
    .A(_09004_),
    .Y(_09011_));
 sg13g2_a21oi_1 _18049_ (.A1(_08927_),
    .A2(_08575_),
    .Y(_09012_),
    .B1(net899));
 sg13g2_o21ai_1 _18050_ (.B1(net1140),
    .Y(_09013_),
    .A1(_08986_),
    .A2(_09012_));
 sg13g2_a21oi_1 _18051_ (.A1(_08987_),
    .A2(_09013_),
    .Y(_09014_),
    .B1(net290));
 sg13g2_nor4_1 _18052_ (.A(_08982_),
    .B(_08999_),
    .C(_09011_),
    .D(_09014_),
    .Y(_09015_));
 sg13g2_o21ai_1 _18053_ (.B1(_08981_),
    .Y(_09016_),
    .A1(_09009_),
    .A2(net293));
 sg13g2_nand2_1 _18054_ (.Y(_09017_),
    .A(net70),
    .B(_08879_));
 sg13g2_a221oi_1 _18055_ (.B2(_09016_),
    .C1(_09017_),
    .B1(_09015_),
    .A1(_08984_),
    .Y(_09018_),
    .A2(_08994_));
 sg13g2_nor3_1 _18056_ (.A(net557),
    .B(_08974_),
    .C(_09018_),
    .Y(_00361_));
 sg13g2_buf_2 _18057_ (.A(_00085_),
    .X(_09019_));
 sg13g2_buf_2 _18058_ (.A(\grid.cell_19_5.se ),
    .X(_09020_));
 sg13g2_xnor2_1 _18059_ (.Y(_09021_),
    .A(_08592_),
    .B(net917));
 sg13g2_xnor2_1 _18060_ (.Y(_09022_),
    .A(_09020_),
    .B(_09021_));
 sg13g2_xnor2_1 _18061_ (.Y(_09023_),
    .A(_08966_),
    .B(net918));
 sg13g2_xnor2_1 _18062_ (.Y(_09024_),
    .A(_09022_),
    .B(_09023_));
 sg13g2_buf_1 _18063_ (.A(_09024_),
    .X(_09025_));
 sg13g2_a21o_1 _18064_ (.A2(_09025_),
    .A1(net282),
    .B1(net578),
    .X(_09026_));
 sg13g2_o21ai_1 _18065_ (.B1(_09025_),
    .Y(_09027_),
    .A1(net1133),
    .A2(net578));
 sg13g2_nor2_1 _18066_ (.A(net283),
    .B(net577),
    .Y(_09028_));
 sg13g2_a221oi_1 _18067_ (.B2(net283),
    .C1(_09028_),
    .B1(_09027_),
    .A1(net1133),
    .Y(_09029_),
    .A2(_09026_));
 sg13g2_xnor2_1 _18068_ (.Y(_09030_),
    .A(net282),
    .B(_09025_));
 sg13g2_nor2b_1 _18069_ (.A(net1133),
    .B_N(_09025_),
    .Y(_09031_));
 sg13g2_a22oi_1 _18070_ (.Y(_09032_),
    .B1(_09031_),
    .B2(_09019_),
    .A2(_09030_),
    .A1(net292));
 sg13g2_o21ai_1 _18071_ (.B1(_09032_),
    .Y(_09033_),
    .A1(_09019_),
    .A2(_09029_));
 sg13g2_inv_1 _18072_ (.Y(_09034_),
    .A(_09020_));
 sg13g2_buf_1 _18073_ (.A(_09034_),
    .X(_09035_));
 sg13g2_nor2_1 _18074_ (.A(net898),
    .B(net567),
    .Y(_09036_));
 sg13g2_nand2_1 _18075_ (.Y(_09037_),
    .A(net555),
    .B(_09036_));
 sg13g2_buf_1 _18076_ (.A(_09020_),
    .X(_09038_));
 sg13g2_nand2_1 _18077_ (.Y(_09039_),
    .A(_09038_),
    .B(net908));
 sg13g2_buf_1 _18078_ (.A(net897),
    .X(_09040_));
 sg13g2_buf_1 _18079_ (.A(net554),
    .X(_09041_));
 sg13g2_nand2_1 _18080_ (.Y(_09042_),
    .A(net275),
    .B(net899));
 sg13g2_nor4_1 _18081_ (.A(net554),
    .B(net899),
    .C(net280),
    .D(net289),
    .Y(_09043_));
 sg13g2_a221oi_1 _18082_ (.B2(net291),
    .C1(_09043_),
    .B1(net148),
    .A1(net556),
    .Y(_09044_),
    .A2(_08615_));
 sg13g2_nand4_1 _18083_ (.B(_09039_),
    .C(_09042_),
    .A(_08292_),
    .Y(_09045_),
    .D(_09044_));
 sg13g2_o21ai_1 _18084_ (.B1(_09045_),
    .Y(_09046_),
    .A1(_08237_),
    .A2(_09037_));
 sg13g2_nand2_1 _18085_ (.Y(_09047_),
    .A(net291),
    .B(_09036_));
 sg13g2_nand2_1 _18086_ (.Y(_09048_),
    .A(_09005_),
    .B(_08239_));
 sg13g2_o21ai_1 _18087_ (.B1(_09048_),
    .Y(_09049_),
    .A1(net899),
    .A2(_08613_));
 sg13g2_nand2b_1 _18088_ (.Y(_09050_),
    .B(_09049_),
    .A_N(_08689_));
 sg13g2_a21oi_1 _18089_ (.A1(_09047_),
    .A2(_09050_),
    .Y(_09051_),
    .B1(net275));
 sg13g2_mux2_1 _18090_ (.A0(_08293_),
    .A1(net554),
    .S(net291),
    .X(_09052_));
 sg13g2_nand4_1 _18091_ (.B(net281),
    .C(net148),
    .A(_08990_),
    .Y(_09053_),
    .D(_09052_));
 sg13g2_inv_1 _18092_ (.Y(_09054_),
    .A(_09019_));
 sg13g2_nand2_1 _18093_ (.Y(_09055_),
    .A(_09054_),
    .B(net292));
 sg13g2_nand3_1 _18094_ (.B(net899),
    .C(net280),
    .A(_08292_),
    .Y(_09056_));
 sg13g2_a21oi_1 _18095_ (.A1(_09005_),
    .A2(net567),
    .Y(_09057_),
    .B1(_08237_));
 sg13g2_a21oi_1 _18096_ (.A1(_08293_),
    .A2(_09036_),
    .Y(_09058_),
    .B1(_09057_));
 sg13g2_nand3_1 _18097_ (.B(_09056_),
    .C(_09058_),
    .A(net275),
    .Y(_09059_));
 sg13g2_nand3_1 _18098_ (.B(_09055_),
    .C(_09059_),
    .A(_09053_),
    .Y(_09060_));
 sg13g2_a21oi_1 _18099_ (.A1(_08989_),
    .A2(net280),
    .Y(_09061_),
    .B1(net275));
 sg13g2_o21ai_1 _18100_ (.B1(_08292_),
    .Y(_09062_),
    .A1(_09036_),
    .A2(_09061_));
 sg13g2_a21oi_1 _18101_ (.A1(_09037_),
    .A2(_09062_),
    .Y(_09063_),
    .B1(net148));
 sg13g2_nor4_1 _18102_ (.A(_09031_),
    .B(_09051_),
    .C(_09060_),
    .D(_09063_),
    .Y(_09064_));
 sg13g2_o21ai_1 _18103_ (.B1(_09030_),
    .Y(_09065_),
    .A1(_09054_),
    .A2(net292));
 sg13g2_a221oi_1 _18104_ (.B2(_09065_),
    .C1(_09017_),
    .B1(_09064_),
    .A1(_09033_),
    .Y(_09066_),
    .A2(_09046_));
 sg13g2_xnor2_1 _18105_ (.Y(_09067_),
    .A(net577),
    .B(_08932_));
 sg13g2_xnor2_1 _18106_ (.Y(_09068_),
    .A(_09025_),
    .B(_09067_));
 sg13g2_a21oi_1 _18107_ (.A1(net126),
    .A2(_09068_),
    .Y(_09069_),
    .B1(net568));
 sg13g2_nor2_1 _18108_ (.A(_08821_),
    .B(_09069_),
    .Y(_09070_));
 sg13g2_a21oi_1 _18109_ (.A1(_06330_),
    .A2(net58),
    .Y(_09071_),
    .B1(_09070_));
 sg13g2_nor3_1 _18110_ (.A(net557),
    .B(_09066_),
    .C(_09071_),
    .Y(_00362_));
 sg13g2_xnor2_1 _18111_ (.Y(_09072_),
    .A(_08331_),
    .B(_08744_));
 sg13g2_xnor2_1 _18112_ (.Y(_09073_),
    .A(_09038_),
    .B(_09072_));
 sg13g2_xnor2_1 _18113_ (.Y(_09074_),
    .A(net576),
    .B(_08967_));
 sg13g2_xnor2_1 _18114_ (.Y(_09075_),
    .A(_09073_),
    .B(_09074_));
 sg13g2_nor2_1 _18115_ (.A(_08607_),
    .B(_09075_),
    .Y(_09076_));
 sg13g2_buf_1 _18116_ (.A(_00117_),
    .X(_09077_));
 sg13g2_inv_1 _18117_ (.Y(_09078_),
    .A(_09077_));
 sg13g2_and4_1 _18118_ (.A(_08672_),
    .B(_09078_),
    .C(_08566_),
    .D(_09073_),
    .X(_09079_));
 sg13g2_nand2_1 _18119_ (.Y(_09080_),
    .A(net555),
    .B(_08284_));
 sg13g2_buf_1 _18120_ (.A(_00147_),
    .X(_09081_));
 sg13g2_nor2_1 _18121_ (.A(net1128),
    .B(_08770_),
    .Y(_09082_));
 sg13g2_buf_1 _18122_ (.A(net279),
    .X(_09083_));
 sg13g2_xnor2_1 _18123_ (.Y(_09084_),
    .A(_08392_),
    .B(net575));
 sg13g2_o21ai_1 _18124_ (.B1(net147),
    .Y(_09085_),
    .A1(net145),
    .A2(_08702_));
 sg13g2_a21oi_1 _18125_ (.A1(_09083_),
    .A2(_09084_),
    .Y(_09086_),
    .B1(_09085_));
 sg13g2_o21ai_1 _18126_ (.B1(_09041_),
    .Y(_09087_),
    .A1(_09082_),
    .A2(_09086_));
 sg13g2_o21ai_1 _18127_ (.B1(_09087_),
    .Y(_09088_),
    .A1(_08770_),
    .A2(_09080_));
 sg13g2_nor4_1 _18128_ (.A(net110),
    .B(_09076_),
    .C(_09079_),
    .D(_09088_),
    .Y(_09089_));
 sg13g2_o21ai_1 _18129_ (.B1(_08759_),
    .Y(_09090_),
    .A1(_09040_),
    .A2(_08805_));
 sg13g2_nor2_1 _18130_ (.A(_09040_),
    .B(_08759_),
    .Y(_09091_));
 sg13g2_a21oi_1 _18131_ (.A1(net1128),
    .A2(_09090_),
    .Y(_09092_),
    .B1(_09091_));
 sg13g2_nand2_1 _18132_ (.Y(_09093_),
    .A(net917),
    .B(net583));
 sg13g2_nor2_1 _18133_ (.A(_09093_),
    .B(_08805_),
    .Y(_09094_));
 sg13g2_o21ai_1 _18134_ (.B1(_09094_),
    .Y(_09095_),
    .A1(net1128),
    .A2(_08759_));
 sg13g2_nand2b_1 _18135_ (.Y(_09096_),
    .B(_09095_),
    .A_N(_09082_));
 sg13g2_nand2b_1 _18136_ (.Y(_09097_),
    .B(net279),
    .A_N(_09081_));
 sg13g2_and2_1 _18137_ (.A(_08768_),
    .B(net295),
    .X(_09098_));
 sg13g2_nor2b_1 _18138_ (.A(_09020_),
    .B_N(net1128),
    .Y(_09099_));
 sg13g2_o21ai_1 _18139_ (.B1(_09099_),
    .Y(_09100_),
    .A1(_08752_),
    .A2(_09098_));
 sg13g2_o21ai_1 _18140_ (.B1(_09100_),
    .Y(_09101_),
    .A1(_08393_),
    .A2(_09097_));
 sg13g2_and2_1 _18141_ (.A(_09020_),
    .B(_08742_),
    .X(_09102_));
 sg13g2_buf_1 _18142_ (.A(_09102_),
    .X(_09103_));
 sg13g2_a21oi_1 _18143_ (.A1(_08377_),
    .A2(_09103_),
    .Y(_09104_),
    .B1(_09091_));
 sg13g2_nor2_1 _18144_ (.A(net288),
    .B(_09104_),
    .Y(_09105_));
 sg13g2_a221oi_1 _18145_ (.B2(net148),
    .C1(_09105_),
    .B1(_09101_),
    .A1(_09041_),
    .Y(_09106_),
    .A2(_09096_));
 sg13g2_o21ai_1 _18146_ (.B1(_09106_),
    .Y(_09107_),
    .A1(net147),
    .A2(_09092_));
 sg13g2_xnor2_1 _18147_ (.Y(_09108_),
    .A(_08611_),
    .B(_09073_));
 sg13g2_o21ai_1 _18148_ (.B1(_09108_),
    .Y(_09109_),
    .A1(_09078_),
    .A2(net290));
 sg13g2_a22oi_1 _18149_ (.Y(_09110_),
    .B1(_09073_),
    .B2(_08672_),
    .A2(net290),
    .A1(_09078_));
 sg13g2_nand2_1 _18150_ (.Y(_09111_),
    .A(_09109_),
    .B(_09110_));
 sg13g2_xnor2_1 _18151_ (.Y(_09112_),
    .A(_09107_),
    .B(_09111_));
 sg13g2_a221oi_1 _18152_ (.B2(_09112_),
    .C1(net58),
    .B1(_09089_),
    .A1(_08607_),
    .Y(_09113_),
    .A2(net69));
 sg13g2_o21ai_1 _18153_ (.B1(net356),
    .Y(_09114_),
    .A1(net31),
    .A2(_08879_));
 sg13g2_nor2_1 _18154_ (.A(_09113_),
    .B(_09114_),
    .Y(_00363_));
 sg13g2_xor2_1 _18155_ (.B(net295),
    .A(net563),
    .X(_09115_));
 sg13g2_xnor2_1 _18156_ (.Y(_09116_),
    .A(_09022_),
    .B(_09115_));
 sg13g2_buf_2 _18157_ (.A(_09116_),
    .X(_09117_));
 sg13g2_nor2_1 _18158_ (.A(net907),
    .B(net1134),
    .Y(_09118_));
 sg13g2_nand2_1 _18159_ (.Y(_09119_),
    .A(_09034_),
    .B(_09118_));
 sg13g2_a21oi_1 _18160_ (.A1(net907),
    .A2(net1134),
    .Y(_09120_),
    .B1(_09020_));
 sg13g2_o21ai_1 _18161_ (.B1(_09081_),
    .Y(_09121_),
    .A1(_09118_),
    .A2(_09120_));
 sg13g2_a21oi_1 _18162_ (.A1(_09119_),
    .A2(_09121_),
    .Y(_09122_),
    .B1(net295));
 sg13g2_and2_1 _18163_ (.A(_08742_),
    .B(net1134),
    .X(_09123_));
 sg13g2_buf_1 _18164_ (.A(_09123_),
    .X(_09124_));
 sg13g2_nand2b_1 _18165_ (.Y(_09125_),
    .B(_09124_),
    .A_N(net1128));
 sg13g2_nand2_1 _18166_ (.Y(_09126_),
    .A(_08749_),
    .B(net1134));
 sg13g2_or3_1 _18167_ (.A(net1128),
    .B(_08742_),
    .C(net1134),
    .X(_09127_));
 sg13g2_nand3_1 _18168_ (.B(_09126_),
    .C(_09127_),
    .A(_08284_),
    .Y(_09128_));
 sg13g2_a21oi_1 _18169_ (.A1(_09125_),
    .A2(_09128_),
    .Y(_09129_),
    .B1(_09034_));
 sg13g2_mux2_1 _18170_ (.A0(net1134),
    .A1(net923),
    .S(_08749_),
    .X(_09130_));
 sg13g2_nor2b_1 _18171_ (.A(net1128),
    .B_N(net923),
    .Y(_09131_));
 sg13g2_a22oi_1 _18172_ (.Y(_09132_),
    .B1(_09131_),
    .B2(_09124_),
    .A2(_09130_),
    .A1(_09099_));
 sg13g2_nor2_1 _18173_ (.A(net289),
    .B(_09132_),
    .Y(_09133_));
 sg13g2_nand3_1 _18174_ (.B(net583),
    .C(_09103_),
    .A(net908),
    .Y(_09134_));
 sg13g2_a21oi_1 _18175_ (.A1(_09119_),
    .A2(_09134_),
    .Y(_09135_),
    .B1(net575));
 sg13g2_nor4_2 _18176_ (.A(_09122_),
    .B(_09129_),
    .C(_09133_),
    .Y(_09136_),
    .D(_09135_));
 sg13g2_nand2_1 _18177_ (.Y(_09137_),
    .A(_08415_),
    .B(net1138));
 sg13g2_or3_1 _18178_ (.A(net913),
    .B(net905),
    .C(net1138),
    .X(_09138_));
 sg13g2_o21ai_1 _18179_ (.B1(_09138_),
    .Y(_09139_),
    .A1(_09136_),
    .A2(_09137_));
 sg13g2_nor2b_1 _18180_ (.A(net922),
    .B_N(net905),
    .Y(_09140_));
 sg13g2_o21ai_1 _18181_ (.B1(net916),
    .Y(_09141_),
    .A1(net572),
    .A2(_09140_));
 sg13g2_nand3_1 _18182_ (.B(net561),
    .C(net916),
    .A(net572),
    .Y(_09142_));
 sg13g2_nor2_1 _18183_ (.A(_09136_),
    .B(_09142_),
    .Y(_09143_));
 sg13g2_a221oi_1 _18184_ (.B2(_09136_),
    .C1(_09143_),
    .B1(_09141_),
    .A1(_08786_),
    .Y(_09144_),
    .A2(_09139_));
 sg13g2_or2_1 _18185_ (.X(_09145_),
    .B(_09144_),
    .A(_09117_));
 sg13g2_nand2_1 _18186_ (.Y(_09146_),
    .A(net567),
    .B(net575));
 sg13g2_mux2_1 _18187_ (.A0(_09146_),
    .A1(_09021_),
    .S(_09083_),
    .X(_09147_));
 sg13g2_o21ai_1 _18188_ (.B1(_09125_),
    .Y(_09148_),
    .A1(_08313_),
    .A2(_09147_));
 sg13g2_or2_1 _18189_ (.X(_09149_),
    .B(_09148_),
    .A(_09035_));
 sg13g2_o21ai_1 _18190_ (.B1(_09035_),
    .Y(_09150_),
    .A1(_09093_),
    .A2(_09126_));
 sg13g2_xor2_1 _18191_ (.B(_09117_),
    .A(_08862_),
    .X(_09151_));
 sg13g2_nor2b_1 _18192_ (.A(net905),
    .B_N(_08414_),
    .Y(_09152_));
 sg13g2_nand3b_1 _18193_ (.B(_09152_),
    .C(net582),
    .Y(_09153_),
    .A_N(net916));
 sg13g2_o21ai_1 _18194_ (.B1(net118),
    .Y(_09154_),
    .A1(_09117_),
    .A2(_09153_));
 sg13g2_a221oi_1 _18195_ (.B2(net285),
    .C1(_09154_),
    .B1(_09151_),
    .A1(_09149_),
    .Y(_09155_),
    .A2(_09150_));
 sg13g2_nand2_1 _18196_ (.Y(_09156_),
    .A(net572),
    .B(_09117_));
 sg13g2_a21oi_1 _18197_ (.A1(_09117_),
    .A2(_09152_),
    .Y(_09157_),
    .B1(net582));
 sg13g2_a21oi_1 _18198_ (.A1(_08843_),
    .A2(_09156_),
    .Y(_09158_),
    .B1(_09157_));
 sg13g2_nand2b_1 _18199_ (.Y(_09159_),
    .B(_08843_),
    .A_N(_08414_));
 sg13g2_o21ai_1 _18200_ (.B1(_09159_),
    .Y(_09160_),
    .A1(net582),
    .A2(_09152_));
 sg13g2_a22oi_1 _18201_ (.Y(_09161_),
    .B1(_09160_),
    .B2(_09117_),
    .A2(_09140_),
    .A1(net916));
 sg13g2_nor2_1 _18202_ (.A(_09136_),
    .B(_09161_),
    .Y(_09162_));
 sg13g2_a21oi_1 _18203_ (.A1(_09136_),
    .A2(_09158_),
    .Y(_09163_),
    .B1(_09162_));
 sg13g2_nand3_1 _18204_ (.B(_09155_),
    .C(_09163_),
    .A(_09145_),
    .Y(_09164_));
 sg13g2_a21oi_1 _18205_ (.A1(net146),
    .A2(net69),
    .Y(_09165_),
    .B1(net58));
 sg13g2_a221oi_1 _18206_ (.B2(_09165_),
    .C1(net617),
    .B1(_09164_),
    .A1(net121),
    .Y(_00364_),
    .A2(net58));
 sg13g2_nor2_1 _18207_ (.A(_01870_),
    .B(_06474_),
    .Y(_09166_));
 sg13g2_nand2_1 _18208_ (.Y(_09167_),
    .A(net327),
    .B(_09166_));
 sg13g2_buf_2 _18209_ (.A(_09167_),
    .X(_09168_));
 sg13g2_buf_1 _18210_ (.A(\grid.cell_1_0.sw ),
    .X(_09169_));
 sg13g2_buf_1 _18211_ (.A(_09169_),
    .X(_09170_));
 sg13g2_or2_1 _18212_ (.X(_09171_),
    .B(net1041),
    .A(net896));
 sg13g2_buf_1 _18213_ (.A(_09171_),
    .X(_09172_));
 sg13g2_buf_1 _18214_ (.A(\grid.cell_1_0.se ),
    .X(_09173_));
 sg13g2_buf_1 _18215_ (.A(_09173_),
    .X(_09174_));
 sg13g2_inv_1 _18216_ (.Y(_09175_),
    .A(net895));
 sg13g2_buf_1 _18217_ (.A(_09175_),
    .X(_09176_));
 sg13g2_nand2_1 _18218_ (.Y(_09177_),
    .A(net274),
    .B(net684));
 sg13g2_buf_1 _18219_ (.A(_00219_),
    .X(_09178_));
 sg13g2_buf_1 _18220_ (.A(_09178_),
    .X(_09179_));
 sg13g2_inv_2 _18221_ (.Y(_09180_),
    .A(_09170_));
 sg13g2_nor2_1 _18222_ (.A(net274),
    .B(_09180_),
    .Y(_09181_));
 sg13g2_nand3_1 _18223_ (.B(net894),
    .C(_09181_),
    .A(net174),
    .Y(_09182_));
 sg13g2_o21ai_1 _18224_ (.B1(_09182_),
    .Y(_09183_),
    .A1(_09172_),
    .A2(_09177_));
 sg13g2_buf_1 _18225_ (.A(_09170_),
    .X(_09184_));
 sg13g2_buf_1 _18226_ (.A(net553),
    .X(_09185_));
 sg13g2_inv_1 _18227_ (.Y(_09186_),
    .A(_09178_));
 sg13g2_nand2_1 _18228_ (.Y(_09187_),
    .A(net709),
    .B(net893));
 sg13g2_nor2_2 _18229_ (.A(net553),
    .B(_02561_),
    .Y(_09188_));
 sg13g2_a21oi_1 _18230_ (.A1(net273),
    .A2(_09187_),
    .Y(_09189_),
    .B1(_09188_));
 sg13g2_nor2_1 _18231_ (.A(net553),
    .B(net374),
    .Y(_09190_));
 sg13g2_buf_1 _18232_ (.A(_09180_),
    .X(_09191_));
 sg13g2_nor2_1 _18233_ (.A(_09180_),
    .B(net709),
    .Y(_09192_));
 sg13g2_a21o_1 _18234_ (.A2(_05060_),
    .A1(net272),
    .B1(_09192_),
    .X(_09193_));
 sg13g2_a22oi_1 _18235_ (.Y(_09194_),
    .B1(_09193_),
    .B2(_04352_),
    .A2(_09190_),
    .A1(net893));
 sg13g2_o21ai_1 _18236_ (.B1(_09194_),
    .Y(_09195_),
    .A1(net359),
    .A2(_09189_));
 sg13g2_buf_1 _18237_ (.A(net895),
    .X(_09196_));
 sg13g2_buf_1 _18238_ (.A(net552),
    .X(_09197_));
 sg13g2_inv_1 _18239_ (.Y(_09198_),
    .A(_02237_));
 sg13g2_nor2_1 _18240_ (.A(net1186),
    .B(_09198_),
    .Y(_09199_));
 sg13g2_mux2_1 _18241_ (.A0(_09198_),
    .A1(net893),
    .S(net373),
    .X(_09200_));
 sg13g2_buf_1 _18242_ (.A(net553),
    .X(_09201_));
 sg13g2_nor2_1 _18243_ (.A(net273),
    .B(_09187_),
    .Y(_09202_));
 sg13g2_a221oi_1 _18244_ (.B2(net270),
    .C1(_09202_),
    .B1(_09200_),
    .A1(_09172_),
    .Y(_09203_),
    .A2(_09199_));
 sg13g2_nor2_1 _18245_ (.A(net271),
    .B(_09203_),
    .Y(_09204_));
 sg13g2_a221oi_1 _18246_ (.B2(net271),
    .C1(_09204_),
    .B1(_09195_),
    .A1(net710),
    .Y(_09205_),
    .A2(_09183_));
 sg13g2_buf_1 _18247_ (.A(_00213_),
    .X(_09206_));
 sg13g2_nand2b_1 _18248_ (.Y(_09207_),
    .B(net1127),
    .A_N(_02874_));
 sg13g2_xnor2_1 _18249_ (.Y(_09208_),
    .A(net1186),
    .B(net895));
 sg13g2_xnor2_1 _18250_ (.Y(_09209_),
    .A(_02259_),
    .B(_09208_));
 sg13g2_xnor2_1 _18251_ (.Y(_09210_),
    .A(_09180_),
    .B(_09209_));
 sg13g2_xnor2_1 _18252_ (.Y(_09211_),
    .A(net711),
    .B(_09210_));
 sg13g2_nand2b_1 _18253_ (.Y(_09212_),
    .B(_02863_),
    .A_N(net1127));
 sg13g2_o21ai_1 _18254_ (.B1(_09212_),
    .Y(_09213_),
    .A1(net1047),
    .A2(_09210_));
 sg13g2_a21oi_1 _18255_ (.A1(_09207_),
    .A2(_09211_),
    .Y(_09214_),
    .B1(_09213_));
 sg13g2_xor2_1 _18256_ (.B(_09214_),
    .A(_09205_),
    .X(_09215_));
 sg13g2_buf_2 _18257_ (.A(\grid.cell_1_0.s ),
    .X(_09216_));
 sg13g2_inv_1 _18258_ (.Y(_09217_),
    .A(_09216_));
 sg13g2_xnor2_1 _18259_ (.Y(_09218_),
    .A(net892),
    .B(_03283_));
 sg13g2_xnor2_1 _18260_ (.Y(_09219_),
    .A(_09210_),
    .B(_09218_));
 sg13g2_nor2_1 _18261_ (.A(net708),
    .B(_09219_),
    .Y(_09220_));
 sg13g2_nor4_1 _18262_ (.A(net1127),
    .B(_02108_),
    .C(_03283_),
    .D(_09210_),
    .Y(_09221_));
 sg13g2_nand2_2 _18263_ (.Y(_09222_),
    .A(net553),
    .B(net709));
 sg13g2_o21ai_1 _18264_ (.B1(net1046),
    .Y(_09223_),
    .A1(_09188_),
    .A2(_09192_));
 sg13g2_o21ai_1 _18265_ (.B1(_09223_),
    .Y(_09224_),
    .A1(net1042),
    .A2(_09222_));
 sg13g2_nor2_1 _18266_ (.A(net272),
    .B(_09187_),
    .Y(_09225_));
 sg13g2_a21oi_1 _18267_ (.A1(net359),
    .A2(_09224_),
    .Y(_09226_),
    .B1(_09225_));
 sg13g2_and2_1 _18268_ (.A(net896),
    .B(_02237_),
    .X(_09227_));
 sg13g2_buf_1 _18269_ (.A(_09227_),
    .X(_09228_));
 sg13g2_and2_1 _18270_ (.A(net1041),
    .B(_09228_),
    .X(_09229_));
 sg13g2_buf_1 _18271_ (.A(_09229_),
    .X(_09230_));
 sg13g2_a21oi_1 _18272_ (.A1(net710),
    .A2(_09230_),
    .Y(_09231_),
    .B1(net271));
 sg13g2_a21oi_1 _18273_ (.A1(net271),
    .A2(_09226_),
    .Y(_09232_),
    .B1(_09231_));
 sg13g2_nor4_1 _18274_ (.A(net107),
    .B(_09220_),
    .C(_09221_),
    .D(_09232_),
    .Y(_09233_));
 sg13g2_a22oi_1 _18275_ (.Y(_09234_),
    .B1(_09215_),
    .B2(_09233_),
    .A2(net75),
    .A1(net708));
 sg13g2_buf_1 _18276_ (.A(_01806_),
    .X(_09235_));
 sg13g2_o21ai_1 _18277_ (.B1(net334),
    .Y(_09236_),
    .A1(net40),
    .A2(_09168_));
 sg13g2_a21oi_1 _18278_ (.A1(_09168_),
    .A2(_09234_),
    .Y(_00365_),
    .B1(_09236_));
 sg13g2_buf_2 _18279_ (.A(\grid.cell_1_1.se ),
    .X(_09237_));
 sg13g2_buf_1 _18280_ (.A(net1126),
    .X(_09238_));
 sg13g2_buf_1 _18281_ (.A(net891),
    .X(_09239_));
 sg13g2_nand2_1 _18282_ (.Y(_09240_),
    .A(net1186),
    .B(net705));
 sg13g2_nand2b_1 _18283_ (.Y(_09241_),
    .B(net891),
    .A_N(_09178_));
 sg13g2_o21ai_1 _18284_ (.B1(_09241_),
    .Y(_09242_),
    .A1(net551),
    .A2(_09240_));
 sg13g2_nor2_1 _18285_ (.A(net551),
    .B(net894),
    .Y(_09243_));
 sg13g2_nor3_1 _18286_ (.A(net369),
    .B(_09240_),
    .C(_09243_),
    .Y(_09244_));
 sg13g2_a21o_1 _18287_ (.A2(_09242_),
    .A1(net369),
    .B1(_09244_),
    .X(_09245_));
 sg13g2_nand2_1 _18288_ (.Y(_09246_),
    .A(net701),
    .B(_09241_));
 sg13g2_o21ai_1 _18289_ (.B1(_09246_),
    .Y(_09247_),
    .A1(net551),
    .A2(net893));
 sg13g2_nand2_1 _18290_ (.Y(_09248_),
    .A(net551),
    .B(net894));
 sg13g2_o21ai_1 _18291_ (.B1(net1033),
    .Y(_09249_),
    .A1(net551),
    .A2(_09179_));
 sg13g2_a21oi_1 _18292_ (.A1(_09248_),
    .A2(_09249_),
    .Y(_09250_),
    .B1(_09240_));
 sg13g2_a21oi_1 _18293_ (.A1(_03530_),
    .A2(_09247_),
    .Y(_09251_),
    .B1(_09250_));
 sg13g2_nor2_1 _18294_ (.A(net1033),
    .B(net891),
    .Y(_09252_));
 sg13g2_nor2_1 _18295_ (.A(net705),
    .B(_09186_),
    .Y(_09253_));
 sg13g2_nand2_1 _18296_ (.Y(_09254_),
    .A(net274),
    .B(_09252_));
 sg13g2_nand4_1 _18297_ (.B(net705),
    .C(net1033),
    .A(net895),
    .Y(_09255_),
    .D(net551));
 sg13g2_a21oi_1 _18298_ (.A1(_09254_),
    .A2(_09255_),
    .Y(_09256_),
    .B1(_02366_));
 sg13g2_a21oi_1 _18299_ (.A1(_09252_),
    .A2(_09253_),
    .Y(_09257_),
    .B1(_09256_));
 sg13g2_o21ai_1 _18300_ (.B1(_09257_),
    .Y(_09258_),
    .A1(net552),
    .A2(_09251_));
 sg13g2_a21oi_1 _18301_ (.A1(net271),
    .A2(_09245_),
    .Y(_09259_),
    .B1(_09258_));
 sg13g2_xnor2_1 _18302_ (.Y(_09260_),
    .A(net891),
    .B(_03207_));
 sg13g2_xor2_1 _18303_ (.B(_09260_),
    .A(_09208_),
    .X(_09261_));
 sg13g2_xnor2_1 _18304_ (.Y(_09262_),
    .A(net708),
    .B(_09261_));
 sg13g2_o21ai_1 _18305_ (.B1(_09212_),
    .Y(_09263_),
    .A1(_00212_),
    .A2(_09261_));
 sg13g2_a21oi_1 _18306_ (.A1(_09207_),
    .A2(_09262_),
    .Y(_09264_),
    .B1(_09263_));
 sg13g2_xnor2_1 _18307_ (.Y(_09265_),
    .A(_09259_),
    .B(_09264_));
 sg13g2_buf_1 _18308_ (.A(_09216_),
    .X(_09266_));
 sg13g2_xnor2_1 _18309_ (.Y(_09267_),
    .A(net890),
    .B(_05137_));
 sg13g2_xor2_1 _18310_ (.B(_09267_),
    .A(_09261_),
    .X(_09268_));
 sg13g2_inv_1 _18311_ (.Y(_09269_),
    .A(_05137_));
 sg13g2_nor3_1 _18312_ (.A(_00212_),
    .B(net1127),
    .C(_09269_),
    .Y(_09270_));
 sg13g2_nand2b_1 _18313_ (.Y(_09271_),
    .B(_09270_),
    .A_N(_09261_));
 sg13g2_xor2_1 _18314_ (.B(net551),
    .A(net1033),
    .X(_09272_));
 sg13g2_nand2_1 _18315_ (.Y(_09273_),
    .A(_03185_),
    .B(net1126));
 sg13g2_nor2_1 _18316_ (.A(_02130_),
    .B(_09273_),
    .Y(_09274_));
 sg13g2_a21oi_1 _18317_ (.A1(_02130_),
    .A2(_09272_),
    .Y(_09275_),
    .B1(_09274_));
 sg13g2_nor2_1 _18318_ (.A(_03530_),
    .B(_09275_),
    .Y(_09276_));
 sg13g2_nor2_1 _18319_ (.A(_09179_),
    .B(_09273_),
    .Y(_09277_));
 sg13g2_o21ai_1 _18320_ (.B1(net271),
    .Y(_09278_),
    .A1(_09276_),
    .A2(_09277_));
 sg13g2_inv_2 _18321_ (.Y(_09279_),
    .A(_09237_));
 sg13g2_buf_1 _18322_ (.A(_09279_),
    .X(_09280_));
 sg13g2_or4_1 _18323_ (.A(_04352_),
    .B(net552),
    .C(net550),
    .D(_03347_),
    .X(_09281_));
 sg13g2_nand4_1 _18324_ (.B(_09271_),
    .C(_09278_),
    .A(net119),
    .Y(_09282_),
    .D(_09281_));
 sg13g2_a21oi_1 _18325_ (.A1(_02087_),
    .A2(_09268_),
    .Y(_09283_),
    .B1(_09282_));
 sg13g2_a22oi_1 _18326_ (.Y(_09284_),
    .B1(_09265_),
    .B2(_09283_),
    .A2(net75),
    .A1(net711));
 sg13g2_o21ai_1 _18327_ (.B1(net334),
    .Y(_09285_),
    .A1(net49),
    .A2(_09168_));
 sg13g2_a21oi_1 _18328_ (.A1(_09168_),
    .A2(_09284_),
    .Y(_00366_),
    .B1(_09285_));
 sg13g2_nand3_1 _18329_ (.B(net108),
    .C(_09166_),
    .A(net1060),
    .Y(_09286_));
 sg13g2_buf_1 _18330_ (.A(_09286_),
    .X(_09287_));
 sg13g2_buf_1 _18331_ (.A(_00218_),
    .X(_09288_));
 sg13g2_inv_2 _18332_ (.Y(_09289_),
    .A(net1125));
 sg13g2_nor2_1 _18333_ (.A(_02119_),
    .B(net1047),
    .Y(_09290_));
 sg13g2_buf_2 _18334_ (.A(\grid.cell_1_2.se ),
    .X(_09291_));
 sg13g2_xnor2_1 _18335_ (.Y(_09292_),
    .A(_09291_),
    .B(_04965_));
 sg13g2_xor2_1 _18336_ (.B(net1126),
    .A(_03174_),
    .X(_09293_));
 sg13g2_xnor2_1 _18337_ (.Y(_09294_),
    .A(_09292_),
    .B(_09293_));
 sg13g2_buf_1 _18338_ (.A(_09294_),
    .X(_09295_));
 sg13g2_o21ai_1 _18339_ (.B1(net1045),
    .Y(_09296_),
    .A1(_09290_),
    .A2(_09295_));
 sg13g2_nand2b_1 _18340_ (.Y(_09297_),
    .B(_02312_),
    .A_N(_09295_));
 sg13g2_nand3_1 _18341_ (.B(_09296_),
    .C(_09297_),
    .A(_02140_),
    .Y(_09298_));
 sg13g2_xnor2_1 _18342_ (.Y(_09299_),
    .A(net1045),
    .B(_09295_));
 sg13g2_nor3_1 _18343_ (.A(net1047),
    .B(_09289_),
    .C(_09295_),
    .Y(_09300_));
 sg13g2_a221oi_1 _18344_ (.B2(_02377_),
    .C1(_09300_),
    .B1(_09299_),
    .A1(_09289_),
    .Y(_09301_),
    .A2(_09298_));
 sg13g2_inv_1 _18345_ (.Y(_09302_),
    .A(_03433_));
 sg13g2_buf_1 _18346_ (.A(_09291_),
    .X(_09303_));
 sg13g2_nand2_1 _18347_ (.Y(_09304_),
    .A(net1029),
    .B(net889));
 sg13g2_xor2_1 _18348_ (.B(_09291_),
    .A(net1029),
    .X(_09305_));
 sg13g2_and2_1 _18349_ (.A(_03326_),
    .B(_09305_),
    .X(_09306_));
 sg13g2_a21oi_1 _18350_ (.A1(net700),
    .A2(_09304_),
    .Y(_09307_),
    .B1(_09306_));
 sg13g2_inv_1 _18351_ (.Y(_09308_),
    .A(_09303_));
 sg13g2_buf_1 _18352_ (.A(_09308_),
    .X(_09309_));
 sg13g2_nand2_1 _18353_ (.Y(_09310_),
    .A(net1034),
    .B(net1031));
 sg13g2_nand3_1 _18354_ (.B(net269),
    .C(_09310_),
    .A(_04236_),
    .Y(_09311_));
 sg13g2_o21ai_1 _18355_ (.B1(_09311_),
    .Y(_09312_),
    .A1(_09302_),
    .A2(_09307_));
 sg13g2_buf_1 _18356_ (.A(net889),
    .X(_09313_));
 sg13g2_a21oi_1 _18357_ (.A1(net705),
    .A2(_09239_),
    .Y(_09314_),
    .B1(net700));
 sg13g2_nor4_1 _18358_ (.A(net366),
    .B(net549),
    .C(_09302_),
    .D(_09314_),
    .Y(_09315_));
 sg13g2_a21oi_1 _18359_ (.A1(net550),
    .A2(_09312_),
    .Y(_09316_),
    .B1(_09315_));
 sg13g2_nor2_1 _18360_ (.A(net163),
    .B(_09316_),
    .Y(_09317_));
 sg13g2_and2_1 _18361_ (.A(_09301_),
    .B(_09317_),
    .X(_09318_));
 sg13g2_buf_1 _18362_ (.A(net551),
    .X(_09319_));
 sg13g2_nor2_1 _18363_ (.A(_03369_),
    .B(_09304_),
    .Y(_09320_));
 sg13g2_o21ai_1 _18364_ (.B1(_04283_),
    .Y(_09321_),
    .A1(_09306_),
    .A2(_09320_));
 sg13g2_o21ai_1 _18365_ (.B1(_09321_),
    .Y(_09322_),
    .A1(_03433_),
    .A2(_09304_));
 sg13g2_nor2_1 _18366_ (.A(_09310_),
    .B(_09304_),
    .Y(_09323_));
 sg13g2_a22oi_1 _18367_ (.Y(_09324_),
    .B1(_09323_),
    .B2(net550),
    .A2(_09289_),
    .A1(_02366_));
 sg13g2_o21ai_1 _18368_ (.B1(_09324_),
    .Y(_09325_),
    .A1(_02108_),
    .A2(_09295_));
 sg13g2_a21oi_1 _18369_ (.A1(_09319_),
    .A2(_09322_),
    .Y(_09326_),
    .B1(_09325_));
 sg13g2_o21ai_1 _18370_ (.B1(_09299_),
    .Y(_09327_),
    .A1(_02377_),
    .A2(_09289_));
 sg13g2_nand2_1 _18371_ (.Y(_09328_),
    .A(net118),
    .B(_09316_));
 sg13g2_a21oi_1 _18372_ (.A1(_09326_),
    .A2(_09327_),
    .Y(_09329_),
    .B1(_09328_));
 sg13g2_xnor2_1 _18373_ (.Y(_09330_),
    .A(_09208_),
    .B(_09299_));
 sg13g2_a21oi_1 _18374_ (.A1(net113),
    .A2(_09330_),
    .Y(_09331_),
    .B1(net369));
 sg13g2_nand2_1 _18375_ (.Y(_09332_),
    .A(net1059),
    .B(_09168_));
 sg13g2_or4_1 _18376_ (.A(_09318_),
    .B(_09329_),
    .C(_09331_),
    .D(_09332_),
    .X(_09333_));
 sg13g2_o21ai_1 _18377_ (.B1(_09333_),
    .Y(_00367_),
    .A1(net27),
    .A2(_09287_));
 sg13g2_buf_2 _18378_ (.A(\grid.cell_1_3.se ),
    .X(_09334_));
 sg13g2_nand2_2 _18379_ (.Y(_09335_),
    .A(_09334_),
    .B(net889));
 sg13g2_inv_2 _18380_ (.Y(_09336_),
    .A(_09334_));
 sg13g2_xnor2_1 _18381_ (.Y(_09337_),
    .A(_04142_),
    .B(net889));
 sg13g2_nor2_1 _18382_ (.A(_09336_),
    .B(_09337_),
    .Y(_09338_));
 sg13g2_buf_1 _18383_ (.A(_09334_),
    .X(_09339_));
 sg13g2_nor3_1 _18384_ (.A(net888),
    .B(net700),
    .C(net269),
    .Y(_09340_));
 sg13g2_o21ai_1 _18385_ (.B1(_04768_),
    .Y(_09341_),
    .A1(_09338_),
    .A2(_09340_));
 sg13g2_o21ai_1 _18386_ (.B1(_09341_),
    .Y(_09342_),
    .A1(net1181),
    .A2(_09335_));
 sg13g2_inv_1 _18387_ (.Y(_09343_),
    .A(_04440_));
 sg13g2_xnor2_1 _18388_ (.Y(_09344_),
    .A(_09334_),
    .B(_09291_));
 sg13g2_xnor2_1 _18389_ (.Y(_09345_),
    .A(_04862_),
    .B(_09344_));
 sg13g2_xnor2_1 _18390_ (.Y(_09346_),
    .A(_04142_),
    .B(_09345_));
 sg13g2_and2_1 _18391_ (.A(_09343_),
    .B(_09346_),
    .X(_09347_));
 sg13g2_inv_1 _18392_ (.Y(_09348_),
    .A(_00215_));
 sg13g2_and2_1 _18393_ (.A(net1124),
    .B(_03207_),
    .X(_09349_));
 sg13g2_nand2_2 _18394_ (.Y(_09350_),
    .A(net1028),
    .B(net1031));
 sg13g2_nor3_1 _18395_ (.A(_04885_),
    .B(_09335_),
    .C(_09350_),
    .Y(_09351_));
 sg13g2_a221oi_1 _18396_ (.B2(_09349_),
    .C1(_09351_),
    .B1(_09347_),
    .A1(net693),
    .Y(_09352_),
    .A2(_09342_));
 sg13g2_inv_1 _18397_ (.Y(_09353_),
    .A(_09344_));
 sg13g2_a22oi_1 _18398_ (.Y(_09354_),
    .B1(_09353_),
    .B2(_04283_),
    .A2(_09335_),
    .A1(_04830_));
 sg13g2_nor2_1 _18399_ (.A(net888),
    .B(net889),
    .Y(_09355_));
 sg13g2_o21ai_1 _18400_ (.B1(_09355_),
    .Y(_09356_),
    .A1(_04830_),
    .A2(_04969_));
 sg13g2_o21ai_1 _18401_ (.B1(_09356_),
    .Y(_09357_),
    .A1(net1026),
    .A2(_09354_));
 sg13g2_buf_1 _18402_ (.A(net888),
    .X(_09358_));
 sg13g2_nor3_1 _18403_ (.A(net1026),
    .B(net548),
    .C(net549),
    .Y(_09359_));
 sg13g2_a22oi_1 _18404_ (.Y(_09360_),
    .B1(_09359_),
    .B2(_09350_),
    .A2(_09357_),
    .A1(_04120_));
 sg13g2_nor2_1 _18405_ (.A(_03369_),
    .B(net1124),
    .Y(_09361_));
 sg13g2_xnor2_1 _18406_ (.Y(_09362_),
    .A(_03380_),
    .B(_09346_));
 sg13g2_a22oi_1 _18407_ (.Y(_09363_),
    .B1(_09346_),
    .B2(_09343_),
    .A2(net1124),
    .A1(_04674_));
 sg13g2_o21ai_1 _18408_ (.B1(_09363_),
    .Y(_09364_),
    .A1(_09361_),
    .A2(_09362_));
 sg13g2_xor2_1 _18409_ (.B(_09364_),
    .A(_09360_),
    .X(_09365_));
 sg13g2_a21oi_1 _18410_ (.A1(_09352_),
    .A2(_09365_),
    .Y(_09366_),
    .B1(net101));
 sg13g2_xor2_1 _18411_ (.B(_09346_),
    .A(_09260_),
    .X(_09367_));
 sg13g2_a21oi_1 _18412_ (.A1(net77),
    .A2(_09367_),
    .Y(_09368_),
    .B1(net366));
 sg13g2_or3_1 _18413_ (.A(_09332_),
    .B(_09366_),
    .C(_09368_),
    .X(_09369_));
 sg13g2_o21ai_1 _18414_ (.B1(_09369_),
    .Y(_00368_),
    .A1(net32),
    .A2(_09287_));
 sg13g2_buf_2 _18415_ (.A(\grid.cell_1_4.se ),
    .X(_09370_));
 sg13g2_buf_1 _18416_ (.A(_09370_),
    .X(_09371_));
 sg13g2_nand2_1 _18417_ (.Y(_09372_),
    .A(net887),
    .B(_09339_));
 sg13g2_buf_1 _18418_ (.A(net887),
    .X(_09373_));
 sg13g2_nand2_1 _18419_ (.Y(_09374_),
    .A(net1028),
    .B(net888));
 sg13g2_xor2_1 _18420_ (.B(_09334_),
    .A(net1180),
    .X(_09375_));
 sg13g2_nand2_1 _18421_ (.Y(_09376_),
    .A(net887),
    .B(_09375_));
 sg13g2_o21ai_1 _18422_ (.B1(_09376_),
    .Y(_09377_),
    .A1(net547),
    .A2(_09374_));
 sg13g2_nand2_1 _18423_ (.Y(_09378_),
    .A(net685),
    .B(_09377_));
 sg13g2_o21ai_1 _18424_ (.B1(_09378_),
    .Y(_09379_),
    .A1(_04857_),
    .A2(_09372_));
 sg13g2_nor2_1 _18425_ (.A(_04959_),
    .B(_09374_),
    .Y(_09380_));
 sg13g2_buf_1 _18426_ (.A(net547),
    .X(_09381_));
 sg13g2_buf_2 _18427_ (.A(_00035_),
    .X(_09382_));
 sg13g2_xnor2_1 _18428_ (.Y(_09383_),
    .A(_09370_),
    .B(_04963_));
 sg13g2_xnor2_1 _18429_ (.Y(_09384_),
    .A(_09375_),
    .B(_09383_));
 sg13g2_nor4_1 _18430_ (.A(_04870_),
    .B(_09382_),
    .C(_04385_),
    .D(_09384_),
    .Y(_09385_));
 sg13g2_a221oi_1 _18431_ (.B2(net267),
    .C1(_09385_),
    .B1(_09380_),
    .A1(net692),
    .Y(_09386_),
    .A2(_09379_));
 sg13g2_xor2_1 _18432_ (.B(_09334_),
    .A(_09370_),
    .X(_09387_));
 sg13g2_a22oi_1 _18433_ (.Y(_09388_),
    .B1(_09387_),
    .B2(_04758_),
    .A2(_09372_),
    .A1(_05101_));
 sg13g2_a21oi_1 _18434_ (.A1(_04943_),
    .A2(_04729_),
    .Y(_09389_),
    .B1(_05101_));
 sg13g2_or3_1 _18435_ (.A(net887),
    .B(net888),
    .C(_09389_),
    .X(_09390_));
 sg13g2_o21ai_1 _18436_ (.B1(_09390_),
    .Y(_09391_),
    .A1(_04944_),
    .A2(_09388_));
 sg13g2_nand2_1 _18437_ (.Y(_09392_),
    .A(_04951_),
    .B(_04768_));
 sg13g2_nor3_1 _18438_ (.A(net692),
    .B(net547),
    .C(net548),
    .Y(_09393_));
 sg13g2_a22oi_1 _18439_ (.Y(_09394_),
    .B1(_09392_),
    .B2(_09393_),
    .A2(_09391_),
    .A1(_04857_));
 sg13g2_nand2_1 _18440_ (.Y(_09395_),
    .A(_09382_),
    .B(_04152_));
 sg13g2_xnor2_1 _18441_ (.Y(_09396_),
    .A(_04495_),
    .B(_09384_));
 sg13g2_nand2b_1 _18442_ (.Y(_09397_),
    .B(net697),
    .A_N(_09382_));
 sg13g2_o21ai_1 _18443_ (.B1(_09397_),
    .Y(_09398_),
    .A1(_04870_),
    .A2(_09384_));
 sg13g2_a21oi_1 _18444_ (.A1(_09395_),
    .A2(_09396_),
    .Y(_09399_),
    .B1(_09398_));
 sg13g2_xnor2_1 _18445_ (.Y(_09400_),
    .A(_09394_),
    .B(_09399_));
 sg13g2_a21oi_1 _18446_ (.A1(_09386_),
    .A2(_09400_),
    .Y(_09401_),
    .B1(net101));
 sg13g2_buf_1 _18447_ (.A(_04642_),
    .X(_09402_));
 sg13g2_xnor2_1 _18448_ (.Y(_09403_),
    .A(_09292_),
    .B(_09384_));
 sg13g2_a21oi_1 _18449_ (.A1(_09402_),
    .A2(_09403_),
    .Y(_09404_),
    .B1(net693));
 sg13g2_or3_1 _18450_ (.A(_09332_),
    .B(_09401_),
    .C(_09404_),
    .X(_09405_));
 sg13g2_o21ai_1 _18451_ (.B1(_09405_),
    .Y(_00369_),
    .A1(net34),
    .A2(_09287_));
 sg13g2_nand2_1 _18452_ (.Y(_09406_),
    .A(_05018_),
    .B(net1023));
 sg13g2_buf_1 _18453_ (.A(\grid.cell_1_5.se ),
    .X(_09407_));
 sg13g2_buf_1 _18454_ (.A(net1123),
    .X(_09408_));
 sg13g2_buf_1 _18455_ (.A(net886),
    .X(_09409_));
 sg13g2_nor3_1 _18456_ (.A(net546),
    .B(net362),
    .C(net547),
    .Y(_09410_));
 sg13g2_inv_1 _18457_ (.Y(_09411_),
    .A(net1123));
 sg13g2_buf_1 _18458_ (.A(_09411_),
    .X(_09412_));
 sg13g2_inv_2 _18459_ (.Y(_09413_),
    .A(net887));
 sg13g2_nand4_1 _18460_ (.B(_05104_),
    .C(net1019),
    .A(net545),
    .Y(_09414_),
    .D(_09413_));
 sg13g2_o21ai_1 _18461_ (.B1(net547),
    .Y(_09415_),
    .A1(net1123),
    .A2(net690));
 sg13g2_a22oi_1 _18462_ (.Y(_09416_),
    .B1(net1019),
    .B2(_05101_),
    .A2(net690),
    .A1(net886));
 sg13g2_and4_1 _18463_ (.A(_04946_),
    .B(_09414_),
    .C(_09415_),
    .D(_09416_),
    .X(_09417_));
 sg13g2_a21oi_1 _18464_ (.A1(_09406_),
    .A2(_09410_),
    .Y(_09418_),
    .B1(_09417_));
 sg13g2_buf_2 _18465_ (.A(_00067_),
    .X(_09419_));
 sg13g2_nand2_1 _18466_ (.Y(_09420_),
    .A(_09419_),
    .B(_04830_));
 sg13g2_xor2_1 _18467_ (.B(net1022),
    .A(net1123),
    .X(_09421_));
 sg13g2_xnor2_1 _18468_ (.Y(_09422_),
    .A(net1179),
    .B(_09370_));
 sg13g2_xor2_1 _18469_ (.B(_09422_),
    .A(_09421_),
    .X(_09423_));
 sg13g2_xnor2_1 _18470_ (.Y(_09424_),
    .A(_05120_),
    .B(_09423_));
 sg13g2_xnor2_1 _18471_ (.Y(_09425_),
    .A(net693),
    .B(_09424_));
 sg13g2_nand2b_1 _18472_ (.Y(_09426_),
    .B(_04758_),
    .A_N(_09419_));
 sg13g2_o21ai_1 _18473_ (.B1(_09426_),
    .Y(_09427_),
    .A1(_04970_),
    .A2(_09424_));
 sg13g2_a21oi_1 _18474_ (.A1(_09420_),
    .A2(_09425_),
    .Y(_09428_),
    .B1(_09427_));
 sg13g2_xor2_1 _18475_ (.B(_09428_),
    .A(_09418_),
    .X(_09429_));
 sg13g2_nand2b_1 _18476_ (.Y(_09430_),
    .B(_04862_),
    .A_N(_09419_));
 sg13g2_nor3_1 _18477_ (.A(_04970_),
    .B(_09424_),
    .C(_09430_),
    .Y(_09431_));
 sg13g2_nand3_1 _18478_ (.B(net1023),
    .C(net547),
    .A(net357),
    .Y(_09432_));
 sg13g2_o21ai_1 _18479_ (.B1(_09432_),
    .Y(_09433_),
    .A1(net357),
    .A2(_09422_));
 sg13g2_nor2_1 _18480_ (.A(_04946_),
    .B(net357),
    .Y(_09434_));
 sg13g2_a22oi_1 _18481_ (.Y(_09435_),
    .B1(_09434_),
    .B2(net267),
    .A2(_09433_),
    .A1(net360));
 sg13g2_nor2_1 _18482_ (.A(net886),
    .B(net357),
    .Y(_09436_));
 sg13g2_nand4_1 _18483_ (.B(net685),
    .C(net267),
    .A(net360),
    .Y(_09437_),
    .D(_09436_));
 sg13g2_o21ai_1 _18484_ (.B1(_09437_),
    .Y(_09438_),
    .A1(net545),
    .A2(_09435_));
 sg13g2_nor3_1 _18485_ (.A(_09429_),
    .B(_09431_),
    .C(_09438_),
    .Y(_09439_));
 sg13g2_xnor2_1 _18486_ (.Y(_09440_),
    .A(net548),
    .B(_04862_));
 sg13g2_xnor2_1 _18487_ (.Y(_09441_),
    .A(_09424_),
    .B(_09440_));
 sg13g2_a21oi_1 _18488_ (.A1(_05517_),
    .A2(_09441_),
    .Y(_09442_),
    .B1(_04945_));
 sg13g2_nor2_1 _18489_ (.A(_09332_),
    .B(_09442_),
    .Y(_09443_));
 sg13g2_o21ai_1 _18490_ (.B1(_09443_),
    .Y(_09444_),
    .A1(net81),
    .A2(_09439_));
 sg13g2_o21ai_1 _18491_ (.B1(_09444_),
    .Y(_00370_),
    .A1(net46),
    .A2(_09287_));
 sg13g2_and2_1 _18492_ (.A(net896),
    .B(_02421_),
    .X(_09445_));
 sg13g2_o21ai_1 _18493_ (.B1(_09172_),
    .Y(_09446_),
    .A1(net886),
    .A2(_09445_));
 sg13g2_nor2_1 _18494_ (.A(net1123),
    .B(_09172_),
    .Y(_09447_));
 sg13g2_a21oi_1 _18495_ (.A1(net689),
    .A2(_09446_),
    .Y(_09448_),
    .B1(_09447_));
 sg13g2_nand2_2 _18496_ (.Y(_09449_),
    .A(_05016_),
    .B(_05059_));
 sg13g2_nor2_1 _18497_ (.A(_09445_),
    .B(_09449_),
    .Y(_09450_));
 sg13g2_o21ai_1 _18498_ (.B1(_09450_),
    .Y(_09451_),
    .A1(net1178),
    .A2(_09172_));
 sg13g2_o21ai_1 _18499_ (.B1(_09451_),
    .Y(_09452_),
    .A1(net1021),
    .A2(_09222_));
 sg13g2_nand2b_1 _18500_ (.Y(_09453_),
    .B(_09230_),
    .A_N(net1178));
 sg13g2_nor2b_1 _18501_ (.A(net1123),
    .B_N(_05008_),
    .Y(_09454_));
 sg13g2_o21ai_1 _18502_ (.B1(_09454_),
    .Y(_09455_),
    .A1(_09188_),
    .A2(_09228_));
 sg13g2_nand2_1 _18503_ (.Y(_09456_),
    .A(_09453_),
    .B(_09455_));
 sg13g2_a21oi_1 _18504_ (.A1(net886),
    .A2(_09230_),
    .Y(_09457_),
    .B1(_09447_));
 sg13g2_nor2_1 _18505_ (.A(net360),
    .B(_09457_),
    .Y(_09458_));
 sg13g2_a221oi_1 _18506_ (.B2(net360),
    .C1(_09458_),
    .B1(_09456_),
    .A1(net546),
    .Y(_09459_),
    .A2(_09452_));
 sg13g2_o21ai_1 _18507_ (.B1(_09459_),
    .Y(_09460_),
    .A1(net359),
    .A2(_09448_));
 sg13g2_inv_1 _18508_ (.Y(_09461_),
    .A(_00099_));
 sg13g2_xnor2_1 _18509_ (.Y(_09462_),
    .A(net1123),
    .B(_09169_));
 sg13g2_xnor2_1 _18510_ (.Y(_09463_),
    .A(_05016_),
    .B(_02237_));
 sg13g2_xnor2_1 _18511_ (.Y(_09464_),
    .A(_09462_),
    .B(_09463_));
 sg13g2_xnor2_1 _18512_ (.Y(_09465_),
    .A(net709),
    .B(_09464_));
 sg13g2_xnor2_1 _18513_ (.Y(_09466_),
    .A(net691),
    .B(_09465_));
 sg13g2_o21ai_1 _18514_ (.B1(_09466_),
    .Y(_09467_),
    .A1(_09461_),
    .A2(_05051_));
 sg13g2_a22oi_1 _18515_ (.Y(_09468_),
    .B1(_09465_),
    .B2(_05025_),
    .A2(_05051_),
    .A1(_09461_));
 sg13g2_nand2_1 _18516_ (.Y(_09469_),
    .A(_09467_),
    .B(_09468_));
 sg13g2_xnor2_1 _18517_ (.Y(_09470_),
    .A(_09460_),
    .B(_09469_));
 sg13g2_buf_1 _18518_ (.A(net546),
    .X(_09471_));
 sg13g2_xor2_1 _18519_ (.B(net374),
    .A(net686),
    .X(_09472_));
 sg13g2_a21oi_1 _18520_ (.A1(net686),
    .A2(net374),
    .Y(_09473_),
    .B1(net273));
 sg13g2_nor2_1 _18521_ (.A(_09198_),
    .B(_09473_),
    .Y(_09474_));
 sg13g2_o21ai_1 _18522_ (.B1(_09474_),
    .Y(_09475_),
    .A1(net272),
    .A2(_09472_));
 sg13g2_o21ai_1 _18523_ (.B1(_09475_),
    .Y(_09476_),
    .A1(net689),
    .A2(_09222_));
 sg13g2_nor2_1 _18524_ (.A(net266),
    .B(net683),
    .Y(_09477_));
 sg13g2_a221oi_1 _18525_ (.B2(_09230_),
    .C1(net99),
    .B1(_09477_),
    .A1(net266),
    .Y(_09478_),
    .A2(_09476_));
 sg13g2_nand4_1 _18526_ (.B(_09461_),
    .C(_04963_),
    .A(_05025_),
    .Y(_09479_),
    .D(_09465_));
 sg13g2_xnor2_1 _18527_ (.Y(_09480_),
    .A(_09383_),
    .B(_09465_));
 sg13g2_nand2_1 _18528_ (.Y(_09481_),
    .A(net357),
    .B(_09480_));
 sg13g2_nand4_1 _18529_ (.B(_09478_),
    .C(_09479_),
    .A(_09470_),
    .Y(_09482_),
    .D(_09481_));
 sg13g2_a22oi_1 _18530_ (.Y(_09483_),
    .B1(_07562_),
    .B2(_09166_),
    .A2(net71),
    .A1(net362));
 sg13g2_a221oi_1 _18531_ (.B2(_09483_),
    .C1(net617),
    .B1(_09482_),
    .A1(_06814_),
    .Y(_00371_),
    .A2(_09166_));
 sg13g2_nand3_1 _18532_ (.B(net104),
    .C(_09168_),
    .A(_02626_),
    .Y(_09484_));
 sg13g2_o21ai_1 _18533_ (.B1(_09484_),
    .Y(_09485_),
    .A1(net121),
    .A2(_09168_));
 sg13g2_nand4_1 _18534_ (.B(net362),
    .C(_05071_),
    .A(net545),
    .Y(_09486_),
    .D(_09228_));
 sg13g2_nand2_1 _18535_ (.Y(_09487_),
    .A(net896),
    .B(net1022));
 sg13g2_nor2_1 _18536_ (.A(net272),
    .B(_05026_),
    .Y(_09488_));
 sg13g2_nor2_1 _18537_ (.A(net273),
    .B(_05041_),
    .Y(_09489_));
 sg13g2_o21ai_1 _18538_ (.B1(_05073_),
    .Y(_09490_),
    .A1(_09488_),
    .A2(_09489_));
 sg13g2_o21ai_1 _18539_ (.B1(_09490_),
    .Y(_09491_),
    .A1(net689),
    .A2(_09487_));
 sg13g2_xnor2_1 _18540_ (.Y(_09492_),
    .A(net690),
    .B(_09464_));
 sg13g2_a22oi_1 _18541_ (.Y(_09493_),
    .B1(_09492_),
    .B2(_09270_),
    .A2(_09491_),
    .A1(net266));
 sg13g2_nand4_1 _18542_ (.B(_09168_),
    .C(_09486_),
    .A(_05354_),
    .Y(_09494_),
    .D(_09493_));
 sg13g2_xor2_1 _18543_ (.B(_09492_),
    .A(_09267_),
    .X(_09495_));
 sg13g2_a21oi_1 _18544_ (.A1(net84),
    .A2(_09495_),
    .Y(_09496_),
    .B1(_02626_));
 sg13g2_nor2_1 _18545_ (.A(net553),
    .B(_05104_),
    .Y(_09497_));
 sg13g2_o21ai_1 _18546_ (.B1(_09454_),
    .Y(_09498_),
    .A1(_09228_),
    .A2(_09497_));
 sg13g2_nand3b_1 _18547_ (.B(net362),
    .C(_09228_),
    .Y(_09499_),
    .A_N(_05009_));
 sg13g2_nand3_1 _18548_ (.B(_09498_),
    .C(_09499_),
    .A(_05071_),
    .Y(_09500_));
 sg13g2_nor2_1 _18549_ (.A(net553),
    .B(net1022),
    .Y(_09501_));
 sg13g2_nand2_1 _18550_ (.Y(_09502_),
    .A(net545),
    .B(_09501_));
 sg13g2_nand3_1 _18551_ (.B(net690),
    .C(_09228_),
    .A(net886),
    .Y(_09503_));
 sg13g2_nand3_1 _18552_ (.B(_09502_),
    .C(_09503_),
    .A(_05121_),
    .Y(_09504_));
 sg13g2_nand2b_1 _18553_ (.Y(_09505_),
    .B(_09501_),
    .A_N(_05008_));
 sg13g2_nand4_1 _18554_ (.B(_05060_),
    .C(_09487_),
    .A(net686),
    .Y(_09506_),
    .D(_09505_));
 sg13g2_o21ai_1 _18555_ (.B1(_09506_),
    .Y(_09507_),
    .A1(net689),
    .A2(_09487_));
 sg13g2_a21oi_1 _18556_ (.A1(net553),
    .A2(net690),
    .Y(_09508_),
    .B1(net886));
 sg13g2_o21ai_1 _18557_ (.B1(_05009_),
    .Y(_09509_),
    .A1(_09501_),
    .A2(_09508_));
 sg13g2_a21oi_1 _18558_ (.A1(_09502_),
    .A2(_09509_),
    .Y(_09510_),
    .B1(_05073_));
 sg13g2_a221oi_1 _18559_ (.B2(net266),
    .C1(_09510_),
    .B1(_09507_),
    .A1(_09500_),
    .Y(_09511_),
    .A2(_09504_));
 sg13g2_xnor2_1 _18560_ (.Y(_09512_),
    .A(_02183_),
    .B(_09492_));
 sg13g2_inv_1 _18561_ (.Y(_09513_),
    .A(_09492_));
 sg13g2_o21ai_1 _18562_ (.B1(_09212_),
    .Y(_09514_),
    .A1(_00212_),
    .A2(_09513_));
 sg13g2_a21oi_1 _18563_ (.A1(_09207_),
    .A2(_09512_),
    .Y(_09515_),
    .B1(_09514_));
 sg13g2_xor2_1 _18564_ (.B(_09515_),
    .A(_09511_),
    .X(_09516_));
 sg13g2_nor3_1 _18565_ (.A(_09494_),
    .B(_09496_),
    .C(_09516_),
    .Y(_09517_));
 sg13g2_a21o_1 _18566_ (.A2(_09485_),
    .A1(net317),
    .B1(_09517_),
    .X(_00372_));
 sg13g2_nor2b_1 _18567_ (.A(net1190),
    .B_N(net1049),
    .Y(_09518_));
 sg13g2_a22oi_1 _18568_ (.Y(_09519_),
    .B1(_09518_),
    .B2(net1053),
    .A2(_06061_),
    .A1(_01849_));
 sg13g2_buf_2 _18569_ (.A(_09519_),
    .X(_09520_));
 sg13g2_or2_1 _18570_ (.X(_09521_),
    .B(_09520_),
    .A(net177));
 sg13g2_buf_2 _18571_ (.A(_09521_),
    .X(_09522_));
 sg13g2_nor3_1 _18572_ (.A(_07600_),
    .B(net176),
    .C(_09522_),
    .Y(_09523_));
 sg13g2_buf_2 _18573_ (.A(_09523_),
    .X(_09524_));
 sg13g2_buf_2 _18574_ (.A(\grid.cell_20_0.sw ),
    .X(_09525_));
 sg13g2_inv_1 _18575_ (.Y(_09526_),
    .A(_09525_));
 sg13g2_buf_1 _18576_ (.A(_09526_),
    .X(_09527_));
 sg13g2_buf_1 _18577_ (.A(\grid.cell_20_0.se ),
    .X(_09528_));
 sg13g2_xnor2_1 _18578_ (.Y(_09529_),
    .A(net914),
    .B(_09528_));
 sg13g2_xnor2_1 _18579_ (.Y(_09530_),
    .A(_08744_),
    .B(_09529_));
 sg13g2_xnor2_1 _18580_ (.Y(_09531_),
    .A(net544),
    .B(_09530_));
 sg13g2_xnor2_1 _18581_ (.Y(_09532_),
    .A(net906),
    .B(_09531_));
 sg13g2_buf_1 _18582_ (.A(_00206_),
    .X(_09533_));
 sg13g2_nand2b_1 _18583_ (.Y(_09534_),
    .B(_09533_),
    .A_N(net913));
 sg13g2_inv_1 _18584_ (.Y(_09535_),
    .A(_09533_));
 sg13g2_nand2_1 _18585_ (.Y(_09536_),
    .A(net913),
    .B(_09535_));
 sg13g2_o21ai_1 _18586_ (.B1(_09536_),
    .Y(_09537_),
    .A1(_08908_),
    .A2(_09531_));
 sg13g2_a21oi_1 _18587_ (.A1(_09532_),
    .A2(_09534_),
    .Y(_09538_),
    .B1(_09537_));
 sg13g2_buf_1 _18588_ (.A(_09528_),
    .X(_09539_));
 sg13g2_buf_1 _18589_ (.A(_09525_),
    .X(_09540_));
 sg13g2_and2_1 _18590_ (.A(net884),
    .B(net907),
    .X(_09541_));
 sg13g2_buf_1 _18591_ (.A(_09541_),
    .X(_09542_));
 sg13g2_and3_1 _18592_ (.X(_09543_),
    .A(net885),
    .B(_08482_),
    .C(net265));
 sg13g2_buf_1 _18593_ (.A(net884),
    .X(_09544_));
 sg13g2_buf_1 _18594_ (.A(net543),
    .X(_09545_));
 sg13g2_nor4_1 _18595_ (.A(_09539_),
    .B(net264),
    .C(net279),
    .D(net285),
    .Y(_09546_));
 sg13g2_o21ai_1 _18596_ (.B1(net287),
    .Y(_09547_),
    .A1(_09543_),
    .A2(_09546_));
 sg13g2_nor2_1 _18597_ (.A(net884),
    .B(net564),
    .Y(_09548_));
 sg13g2_nand2b_1 _18598_ (.Y(_09549_),
    .B(net564),
    .A_N(_08482_));
 sg13g2_nor2b_1 _18599_ (.A(net884),
    .B_N(net564),
    .Y(_09550_));
 sg13g2_a21o_1 _18600_ (.A2(_09549_),
    .A1(net543),
    .B1(_09550_),
    .X(_09551_));
 sg13g2_nand2b_1 _18601_ (.Y(_09552_),
    .B(_09540_),
    .A_N(net564));
 sg13g2_nand2b_1 _18602_ (.Y(_09553_),
    .B(net573),
    .A_N(net543));
 sg13g2_a21oi_1 _18603_ (.A1(_09552_),
    .A2(_09553_),
    .Y(_09554_),
    .B1(net574));
 sg13g2_a221oi_1 _18604_ (.B2(net285),
    .C1(_09554_),
    .B1(_09551_),
    .A1(_08483_),
    .Y(_09555_),
    .A2(_09548_));
 sg13g2_nor2_1 _18605_ (.A(net914),
    .B(net285),
    .Y(_09556_));
 sg13g2_inv_1 _18606_ (.Y(_09557_),
    .A(_09548_));
 sg13g2_o21ai_1 _18607_ (.B1(_08755_),
    .Y(_09558_),
    .A1(_08763_),
    .A2(_08482_));
 sg13g2_nor2_1 _18608_ (.A(net264),
    .B(_09549_),
    .Y(_09559_));
 sg13g2_a221oi_1 _18609_ (.B2(net264),
    .C1(_09559_),
    .B1(_09558_),
    .A1(_09556_),
    .Y(_09560_),
    .A2(_09557_));
 sg13g2_inv_2 _18610_ (.Y(_09561_),
    .A(net885));
 sg13g2_mux2_1 _18611_ (.A0(_09555_),
    .A1(_09560_),
    .S(_09561_),
    .X(_09562_));
 sg13g2_xor2_1 _18612_ (.B(net906),
    .A(net913),
    .X(_09563_));
 sg13g2_nor2_1 _18613_ (.A(_09533_),
    .B(_09563_),
    .Y(_09564_));
 sg13g2_nor2_1 _18614_ (.A(_08908_),
    .B(_09531_),
    .Y(_09565_));
 sg13g2_xor2_1 _18615_ (.B(net564),
    .A(net543),
    .X(_09566_));
 sg13g2_mux2_1 _18616_ (.A0(net265),
    .A1(_09566_),
    .S(net574),
    .X(_09567_));
 sg13g2_nor2_1 _18617_ (.A(net544),
    .B(_09549_),
    .Y(_09568_));
 sg13g2_a21oi_1 _18618_ (.A1(net146),
    .A2(_09567_),
    .Y(_09569_),
    .B1(_09568_));
 sg13g2_nor2_1 _18619_ (.A(net885),
    .B(_09527_),
    .Y(_09570_));
 sg13g2_nand3_1 _18620_ (.B(_08805_),
    .C(_09570_),
    .A(net574),
    .Y(_09571_));
 sg13g2_o21ai_1 _18621_ (.B1(_09571_),
    .Y(_09572_),
    .A1(_09561_),
    .A2(_09569_));
 sg13g2_a221oi_1 _18622_ (.B2(_09565_),
    .C1(_09572_),
    .B1(_09564_),
    .A1(_09547_),
    .Y(_09573_),
    .A2(_09562_));
 sg13g2_nand2_1 _18623_ (.Y(_09574_),
    .A(_09538_),
    .B(_09573_));
 sg13g2_nand2_1 _18624_ (.Y(_09575_),
    .A(_09547_),
    .B(_09562_));
 sg13g2_and2_1 _18625_ (.A(_09565_),
    .B(_09564_),
    .X(_09576_));
 sg13g2_or4_1 _18626_ (.A(_09575_),
    .B(_09572_),
    .C(_09538_),
    .D(_09576_),
    .X(_09577_));
 sg13g2_nand3_1 _18627_ (.B(_09574_),
    .C(_09577_),
    .A(net82),
    .Y(_09578_));
 sg13g2_buf_1 _18628_ (.A(\grid.cell_20_0.s ),
    .X(_09579_));
 sg13g2_buf_1 _18629_ (.A(_09579_),
    .X(_09580_));
 sg13g2_xnor2_1 _18630_ (.Y(_09581_),
    .A(_09580_),
    .B(_09563_));
 sg13g2_xor2_1 _18631_ (.B(_09581_),
    .A(_09531_),
    .X(_09582_));
 sg13g2_a21oi_1 _18632_ (.A1(net98),
    .A2(_09582_),
    .Y(_09583_),
    .B1(net904));
 sg13g2_nor2_1 _18633_ (.A(_09524_),
    .B(_09583_),
    .Y(_09584_));
 sg13g2_a22oi_1 _18634_ (.Y(_09585_),
    .B1(_09578_),
    .B2(_09584_),
    .A2(_09524_),
    .A1(net40));
 sg13g2_nor2_1 _18635_ (.A(net370),
    .B(_09585_),
    .Y(_00373_));
 sg13g2_buf_1 _18636_ (.A(\grid.cell_20_1.se ),
    .X(_09586_));
 sg13g2_inv_2 _18637_ (.Y(_09587_),
    .A(net1122));
 sg13g2_xnor2_1 _18638_ (.Y(_09588_),
    .A(_09587_),
    .B(_08827_));
 sg13g2_xor2_1 _18639_ (.B(_09588_),
    .A(_09529_),
    .X(_09589_));
 sg13g2_xnor2_1 _18640_ (.Y(_09590_),
    .A(_08812_),
    .B(_09589_));
 sg13g2_o21ai_1 _18641_ (.B1(_09536_),
    .Y(_09591_),
    .A1(net905),
    .A2(_09589_));
 sg13g2_a21oi_1 _18642_ (.A1(_09534_),
    .A2(_09590_),
    .Y(_09592_),
    .B1(_09591_));
 sg13g2_a21oi_1 _18643_ (.A1(_08391_),
    .A2(net912),
    .Y(_09593_),
    .B1(_08483_));
 sg13g2_nand2_1 _18644_ (.Y(_09594_),
    .A(net574),
    .B(net912));
 sg13g2_xnor2_1 _18645_ (.Y(_09595_),
    .A(_08824_),
    .B(net1122));
 sg13g2_xnor2_1 _18646_ (.Y(_09596_),
    .A(_09561_),
    .B(_09595_));
 sg13g2_mux2_1 _18647_ (.A0(_09593_),
    .A1(_09594_),
    .S(_09596_),
    .X(_09597_));
 sg13g2_xnor2_1 _18648_ (.Y(_09598_),
    .A(_09592_),
    .B(_09597_));
 sg13g2_buf_1 _18649_ (.A(net1122),
    .X(_09599_));
 sg13g2_buf_1 _18650_ (.A(_09599_),
    .X(_09600_));
 sg13g2_nand2_1 _18651_ (.Y(_09601_),
    .A(net278),
    .B(net542));
 sg13g2_buf_1 _18652_ (.A(net885),
    .X(_09602_));
 sg13g2_o21ai_1 _18653_ (.B1(_09602_),
    .Y(_09603_),
    .A1(net560),
    .A2(net542));
 sg13g2_xor2_1 _18654_ (.B(_08811_),
    .A(net913),
    .X(_09604_));
 sg13g2_or4_1 _18655_ (.A(_09533_),
    .B(net561),
    .C(_09604_),
    .D(_09589_),
    .X(_09605_));
 sg13g2_nand3_1 _18656_ (.B(_09603_),
    .C(_09605_),
    .A(_09601_),
    .Y(_09606_));
 sg13g2_inv_1 _18657_ (.Y(_09607_),
    .A(_09597_));
 sg13g2_a21oi_1 _18658_ (.A1(_09601_),
    .A2(_09603_),
    .Y(_09608_),
    .B1(_09607_));
 sg13g2_a21oi_1 _18659_ (.A1(_09592_),
    .A2(_09608_),
    .Y(_09609_),
    .B1(net99));
 sg13g2_o21ai_1 _18660_ (.B1(_09609_),
    .Y(_09610_),
    .A1(_09598_),
    .A2(_09606_));
 sg13g2_xnor2_1 _18661_ (.Y(_09611_),
    .A(_09580_),
    .B(_08861_));
 sg13g2_xnor2_1 _18662_ (.Y(_09612_),
    .A(_09589_),
    .B(_09611_));
 sg13g2_a21oi_1 _18663_ (.A1(net98),
    .A2(_09612_),
    .Y(_09613_),
    .B1(net562));
 sg13g2_nor2_1 _18664_ (.A(_09524_),
    .B(_09613_),
    .Y(_09614_));
 sg13g2_a22oi_1 _18665_ (.Y(_09615_),
    .B1(_09610_),
    .B2(_09614_),
    .A2(_09524_),
    .A1(net49));
 sg13g2_nor2_1 _18666_ (.A(net370),
    .B(_09615_),
    .Y(_00374_));
 sg13g2_nor2_2 _18667_ (.A(_07600_),
    .B(_09522_),
    .Y(_09616_));
 sg13g2_nand2_2 _18668_ (.Y(_09617_),
    .A(net158),
    .B(_09616_));
 sg13g2_nand3_1 _18669_ (.B(net104),
    .C(_09617_),
    .A(net278),
    .Y(_09618_));
 sg13g2_o21ai_1 _18670_ (.B1(_09618_),
    .Y(_09619_),
    .A1(net35),
    .A2(_09617_));
 sg13g2_buf_1 _18671_ (.A(_00205_),
    .X(_09620_));
 sg13g2_inv_2 _18672_ (.Y(_09621_),
    .A(net1121));
 sg13g2_buf_1 _18673_ (.A(\grid.cell_20_2.se ),
    .X(_09622_));
 sg13g2_xor2_1 _18674_ (.B(_08880_),
    .A(_09622_),
    .X(_09623_));
 sg13g2_xnor2_1 _18675_ (.Y(_09624_),
    .A(_08470_),
    .B(_09623_));
 sg13g2_xnor2_1 _18676_ (.Y(_09625_),
    .A(net1137),
    .B(net1122));
 sg13g2_xnor2_1 _18677_ (.Y(_09626_),
    .A(_09624_),
    .B(_09625_));
 sg13g2_xnor2_1 _18678_ (.Y(_09627_),
    .A(net565),
    .B(_09626_));
 sg13g2_o21ai_1 _18679_ (.B1(_09627_),
    .Y(_09628_),
    .A1(net287),
    .A2(_09621_));
 sg13g2_inv_1 _18680_ (.Y(_09629_),
    .A(net901));
 sg13g2_a22oi_1 _18681_ (.Y(_09630_),
    .B1(_09629_),
    .B2(_09626_),
    .A2(_09621_),
    .A1(net287));
 sg13g2_and2_1 _18682_ (.A(_09628_),
    .B(_09630_),
    .X(_09631_));
 sg13g2_buf_1 _18683_ (.A(_09622_),
    .X(_09632_));
 sg13g2_buf_1 _18684_ (.A(net881),
    .X(_09633_));
 sg13g2_buf_1 _18685_ (.A(_09633_),
    .X(_09634_));
 sg13g2_nor2_1 _18686_ (.A(_09634_),
    .B(net559),
    .Y(_09635_));
 sg13g2_nand2_1 _18687_ (.Y(_09636_),
    .A(net571),
    .B(net570));
 sg13g2_and2_1 _18688_ (.A(_09632_),
    .B(_08881_),
    .X(_09637_));
 sg13g2_buf_1 _18689_ (.A(_09637_),
    .X(_09638_));
 sg13g2_nand2_1 _18690_ (.Y(_09639_),
    .A(net912),
    .B(_09623_));
 sg13g2_o21ai_1 _18691_ (.B1(_09639_),
    .Y(_09640_),
    .A1(net284),
    .A2(_09638_));
 sg13g2_a22oi_1 _18692_ (.Y(_09641_),
    .B1(_09640_),
    .B2(_00210_),
    .A2(_09636_),
    .A1(_09635_));
 sg13g2_buf_1 _18693_ (.A(_09587_),
    .X(_09642_));
 sg13g2_o21ai_1 _18694_ (.B1(net284),
    .Y(_09643_),
    .A1(_08422_),
    .A2(_09642_));
 sg13g2_nand3_1 _18695_ (.B(_09643_),
    .C(_09635_),
    .A(_00210_),
    .Y(_09644_));
 sg13g2_o21ai_1 _18696_ (.B1(_09644_),
    .Y(_09645_),
    .A1(_09600_),
    .A2(_09641_));
 sg13g2_xnor2_1 _18697_ (.Y(_09646_),
    .A(_09631_),
    .B(_09645_));
 sg13g2_nand2b_1 _18698_ (.Y(_09647_),
    .B(_09638_),
    .A_N(_09636_));
 sg13g2_nand2_1 _18699_ (.Y(_09648_),
    .A(net540),
    .B(_08892_));
 sg13g2_o21ai_1 _18700_ (.B1(_09639_),
    .Y(_09649_),
    .A1(net571),
    .A2(_09648_));
 sg13g2_a221oi_1 _18701_ (.B2(net284),
    .C1(_09642_),
    .B1(_09649_),
    .A1(_08525_),
    .Y(_09650_),
    .A2(_09638_));
 sg13g2_a21o_1 _18702_ (.A2(_09647_),
    .A1(net539),
    .B1(_09650_),
    .X(_09651_));
 sg13g2_xnor2_1 _18703_ (.Y(_09652_),
    .A(net287),
    .B(net562));
 sg13g2_nand4_1 _18704_ (.B(_09629_),
    .C(_09626_),
    .A(_09621_),
    .Y(_09653_),
    .D(_09652_));
 sg13g2_nand4_1 _18705_ (.B(_09617_),
    .C(_09651_),
    .A(net1002),
    .Y(_09654_),
    .D(_09653_));
 sg13g2_xnor2_1 _18706_ (.Y(_09655_),
    .A(_09529_),
    .B(_09627_));
 sg13g2_a21oi_1 _18707_ (.A1(net83),
    .A2(_09655_),
    .Y(_09656_),
    .B1(_08891_));
 sg13g2_nor3_1 _18708_ (.A(_09646_),
    .B(_09654_),
    .C(_09656_),
    .Y(_09657_));
 sg13g2_a21o_1 _18709_ (.A2(_09619_),
    .A1(net317),
    .B1(_09657_),
    .X(_00375_));
 sg13g2_nand2_1 _18710_ (.Y(_09658_),
    .A(net716),
    .B(_09524_));
 sg13g2_buf_2 _18711_ (.A(\grid.cell_20_3.se ),
    .X(_09659_));
 sg13g2_buf_1 _18712_ (.A(_09659_),
    .X(_09660_));
 sg13g2_buf_1 _18713_ (.A(net880),
    .X(_09661_));
 sg13g2_buf_1 _18714_ (.A(_09661_),
    .X(_09662_));
 sg13g2_nand2_1 _18715_ (.Y(_09663_),
    .A(net540),
    .B(_08925_));
 sg13g2_nand2_1 _18716_ (.Y(_09664_),
    .A(net900),
    .B(net570));
 sg13g2_xor2_1 _18717_ (.B(net911),
    .A(net900),
    .X(_09665_));
 sg13g2_nand2_1 _18718_ (.Y(_09666_),
    .A(net540),
    .B(_09665_));
 sg13g2_o21ai_1 _18719_ (.B1(_09666_),
    .Y(_09667_),
    .A1(_09633_),
    .A2(_09664_));
 sg13g2_nand2_1 _18720_ (.Y(_09668_),
    .A(net569),
    .B(_09667_));
 sg13g2_o21ai_1 _18721_ (.B1(_09668_),
    .Y(_09669_),
    .A1(net1135),
    .A2(_09663_));
 sg13g2_nor2_1 _18722_ (.A(_09662_),
    .B(_09663_),
    .Y(_09670_));
 sg13g2_nor2_1 _18723_ (.A(net282),
    .B(_08470_),
    .Y(_09671_));
 sg13g2_buf_1 _18724_ (.A(_00204_),
    .X(_09672_));
 sg13g2_xor2_1 _18725_ (.B(_08468_),
    .A(_09632_),
    .X(_09673_));
 sg13g2_xnor2_1 _18726_ (.Y(_09674_),
    .A(_08932_),
    .B(_09673_));
 sg13g2_xnor2_1 _18727_ (.Y(_09675_),
    .A(net880),
    .B(_09674_));
 sg13g2_nor4_1 _18728_ (.A(net1120),
    .B(_08931_),
    .C(_08827_),
    .D(_09675_),
    .Y(_09676_));
 sg13g2_a221oi_1 _18729_ (.B2(_09671_),
    .C1(_09676_),
    .B1(_09670_),
    .A1(net262),
    .Y(_09677_),
    .A2(_09669_));
 sg13g2_nor4_1 _18730_ (.A(net880),
    .B(net540),
    .C(net900),
    .D(_08529_),
    .Y(_09678_));
 sg13g2_inv_2 _18731_ (.Y(_09679_),
    .A(net880));
 sg13g2_o21ai_1 _18732_ (.B1(_09663_),
    .Y(_09680_),
    .A1(_09679_),
    .A2(_08942_));
 sg13g2_nand2_1 _18733_ (.Y(_09681_),
    .A(_09660_),
    .B(net881));
 sg13g2_o21ai_1 _18734_ (.B1(_09681_),
    .Y(_09682_),
    .A1(net282),
    .A2(net570));
 sg13g2_nor3_1 _18735_ (.A(_09678_),
    .B(_09680_),
    .C(_09682_),
    .Y(_09683_));
 sg13g2_nor3_1 _18736_ (.A(_09634_),
    .B(net558),
    .C(_09671_),
    .Y(_09684_));
 sg13g2_a22oi_1 _18737_ (.Y(_09685_),
    .B1(_09684_),
    .B2(_09679_),
    .A2(_09683_),
    .A1(net1135));
 sg13g2_nand2_1 _18738_ (.Y(_09686_),
    .A(_08422_),
    .B(_09672_));
 sg13g2_xnor2_1 _18739_ (.Y(_09687_),
    .A(net560),
    .B(_09675_));
 sg13g2_nand2b_1 _18740_ (.Y(_09688_),
    .B(net571),
    .A_N(_09672_));
 sg13g2_o21ai_1 _18741_ (.B1(_09688_),
    .Y(_09689_),
    .A1(_08931_),
    .A2(_09675_));
 sg13g2_a21oi_1 _18742_ (.A1(_09686_),
    .A2(_09687_),
    .Y(_09690_),
    .B1(_09689_));
 sg13g2_xnor2_1 _18743_ (.Y(_09691_),
    .A(_09685_),
    .B(_09690_));
 sg13g2_a21oi_1 _18744_ (.A1(_09677_),
    .A2(_09691_),
    .Y(_09692_),
    .B1(net106));
 sg13g2_xnor2_1 _18745_ (.Y(_09693_),
    .A(_09588_),
    .B(_09675_));
 sg13g2_a21oi_1 _18746_ (.A1(net111),
    .A2(_09693_),
    .Y(_09694_),
    .B1(net276));
 sg13g2_or4_1 _18747_ (.A(net1057),
    .B(_09524_),
    .C(_09692_),
    .D(_09694_),
    .X(_09695_));
 sg13g2_o21ai_1 _18748_ (.B1(_09695_),
    .Y(_00376_),
    .A1(net32),
    .A2(_09658_));
 sg13g2_buf_1 _18749_ (.A(\grid.cell_20_4.se ),
    .X(_09696_));
 sg13g2_buf_1 _18750_ (.A(_09696_),
    .X(_09697_));
 sg13g2_buf_1 _18751_ (.A(net879),
    .X(_09698_));
 sg13g2_nor4_1 _18752_ (.A(net537),
    .B(net880),
    .C(net898),
    .D(_08611_),
    .Y(_09699_));
 sg13g2_a221oi_1 _18753_ (.B2(net282),
    .C1(_09699_),
    .B1(net909),
    .A1(net538),
    .Y(_09700_),
    .A2(net899));
 sg13g2_o21ai_1 _18754_ (.B1(net537),
    .Y(_09701_),
    .A1(net538),
    .A2(net898));
 sg13g2_and2_1 _18755_ (.A(net1133),
    .B(_09701_),
    .X(_09702_));
 sg13g2_nor3_1 _18756_ (.A(net537),
    .B(net262),
    .C(net899),
    .Y(_09703_));
 sg13g2_nand2_1 _18757_ (.Y(_09704_),
    .A(net909),
    .B(net569));
 sg13g2_a22oi_1 _18758_ (.Y(_09705_),
    .B1(_09703_),
    .B2(_09704_),
    .A2(_09702_),
    .A1(_09700_));
 sg13g2_buf_2 _18759_ (.A(_00052_),
    .X(_09706_));
 sg13g2_nand2_1 _18760_ (.Y(_09707_),
    .A(_09706_),
    .B(_08470_));
 sg13g2_xnor2_1 _18761_ (.Y(_09708_),
    .A(_09696_),
    .B(_09659_));
 sg13g2_xor2_1 _18762_ (.B(_09708_),
    .A(_08967_),
    .X(_09709_));
 sg13g2_xnor2_1 _18763_ (.Y(_09710_),
    .A(_08529_),
    .B(_09709_));
 sg13g2_xnor2_1 _18764_ (.Y(_09711_),
    .A(net559),
    .B(_09710_));
 sg13g2_nand2b_1 _18765_ (.Y(_09712_),
    .B(net570),
    .A_N(_09706_));
 sg13g2_o21ai_1 _18766_ (.B1(_09712_),
    .Y(_09713_),
    .A1(_08975_),
    .A2(_09710_));
 sg13g2_a21oi_1 _18767_ (.A1(_09707_),
    .A2(_09711_),
    .Y(_09714_),
    .B1(_09713_));
 sg13g2_xor2_1 _18768_ (.B(_09714_),
    .A(_09705_),
    .X(_09715_));
 sg13g2_nor4_1 _18769_ (.A(_08975_),
    .B(_09706_),
    .C(_08897_),
    .D(_09710_),
    .Y(_09716_));
 sg13g2_buf_1 _18770_ (.A(_09698_),
    .X(_09717_));
 sg13g2_nand2_1 _18771_ (.Y(_09718_),
    .A(net538),
    .B(net898));
 sg13g2_xnor2_1 _18772_ (.Y(_09719_),
    .A(_08966_),
    .B(net910));
 sg13g2_nor2_1 _18773_ (.A(_09679_),
    .B(_09719_),
    .Y(_09720_));
 sg13g2_nor3_1 _18774_ (.A(_09660_),
    .B(_08985_),
    .C(net282),
    .Y(_09721_));
 sg13g2_o21ai_1 _18775_ (.B1(net568),
    .Y(_09722_),
    .A1(_09720_),
    .A2(_09721_));
 sg13g2_o21ai_1 _18776_ (.B1(_09722_),
    .Y(_09723_),
    .A1(net1133),
    .A2(_09718_));
 sg13g2_nor3_1 _18777_ (.A(_09717_),
    .B(_09704_),
    .C(_09718_),
    .Y(_09724_));
 sg13g2_a21oi_1 _18778_ (.A1(_09717_),
    .A2(_09723_),
    .Y(_09725_),
    .B1(_09724_));
 sg13g2_nand2b_1 _18779_ (.Y(_09726_),
    .B(_09725_),
    .A_N(_09716_));
 sg13g2_o21ai_1 _18780_ (.B1(net83),
    .Y(_09727_),
    .A1(_09715_),
    .A2(_09726_));
 sg13g2_xor2_1 _18781_ (.B(_09710_),
    .A(_09624_),
    .X(_09728_));
 sg13g2_o21ai_1 _18782_ (.B1(_08942_),
    .Y(_09729_),
    .A1(net115),
    .A2(_09728_));
 sg13g2_nand4_1 _18783_ (.B(_09617_),
    .C(_09727_),
    .A(net637),
    .Y(_09730_),
    .D(_09729_));
 sg13g2_o21ai_1 _18784_ (.B1(_09730_),
    .Y(_00377_),
    .A1(net34),
    .A2(_09658_));
 sg13g2_buf_1 _18785_ (.A(\grid.cell_20_5.se ),
    .X(_09731_));
 sg13g2_buf_1 _18786_ (.A(_09731_),
    .X(_09732_));
 sg13g2_buf_1 _18787_ (.A(net878),
    .X(_09733_));
 sg13g2_nor4_1 _18788_ (.A(net536),
    .B(net879),
    .C(net897),
    .D(net566),
    .Y(_09734_));
 sg13g2_nand2_1 _18789_ (.Y(_09735_),
    .A(net879),
    .B(net897));
 sg13g2_nand2_1 _18790_ (.Y(_09736_),
    .A(net536),
    .B(net897));
 sg13g2_nand2_1 _18791_ (.Y(_09737_),
    .A(_09735_),
    .B(_09736_));
 sg13g2_nor2_1 _18792_ (.A(net566),
    .B(net909),
    .Y(_09738_));
 sg13g2_and2_1 _18793_ (.A(net536),
    .B(net879),
    .X(_09739_));
 sg13g2_buf_1 _18794_ (.A(_09739_),
    .X(_09740_));
 sg13g2_nor4_1 _18795_ (.A(_09734_),
    .B(_09737_),
    .C(_09738_),
    .D(_09740_),
    .Y(_09741_));
 sg13g2_buf_1 _18796_ (.A(net878),
    .X(_09742_));
 sg13g2_buf_1 _18797_ (.A(net535),
    .X(_09743_));
 sg13g2_nor3_1 _18798_ (.A(net260),
    .B(_09698_),
    .C(net275),
    .Y(_09744_));
 sg13g2_a22oi_1 _18799_ (.Y(_09745_),
    .B1(_09744_),
    .B2(_08616_),
    .A2(_09741_),
    .A1(net1131));
 sg13g2_buf_2 _18800_ (.A(_00084_),
    .X(_09746_));
 sg13g2_nand2_1 _18801_ (.Y(_09747_),
    .A(_09746_),
    .B(net282));
 sg13g2_xor2_1 _18802_ (.B(net1134),
    .A(_09020_),
    .X(_09748_));
 sg13g2_xnor2_1 _18803_ (.Y(_09749_),
    .A(net879),
    .B(net1136));
 sg13g2_xnor2_1 _18804_ (.Y(_09750_),
    .A(_09748_),
    .B(_09749_));
 sg13g2_xnor2_1 _18805_ (.Y(_09751_),
    .A(_09733_),
    .B(_09750_));
 sg13g2_xnor2_1 _18806_ (.Y(_09752_),
    .A(net558),
    .B(_09751_));
 sg13g2_nand2b_1 _18807_ (.Y(_09753_),
    .B(net569),
    .A_N(_09746_));
 sg13g2_o21ai_1 _18808_ (.B1(_09753_),
    .Y(_09754_),
    .A1(_09019_),
    .A2(_09751_));
 sg13g2_a21oi_1 _18809_ (.A1(_09747_),
    .A2(_09752_),
    .Y(_09755_),
    .B1(_09754_));
 sg13g2_xnor2_1 _18810_ (.Y(_09756_),
    .A(_09745_),
    .B(_09755_));
 sg13g2_nor2_1 _18811_ (.A(_09019_),
    .B(_09751_),
    .Y(_09757_));
 sg13g2_nor2b_1 _18812_ (.A(_09746_),
    .B_N(_08932_),
    .Y(_09758_));
 sg13g2_inv_1 _18813_ (.Y(_09759_),
    .A(net879));
 sg13g2_xnor2_1 _18814_ (.Y(_09760_),
    .A(net897),
    .B(net1136));
 sg13g2_nor2_1 _18815_ (.A(net534),
    .B(_09760_),
    .Y(_09761_));
 sg13g2_nor3_1 _18816_ (.A(net537),
    .B(net555),
    .C(_08611_),
    .Y(_09762_));
 sg13g2_o21ai_1 _18817_ (.B1(net280),
    .Y(_09763_),
    .A1(_09761_),
    .A2(_09762_));
 sg13g2_o21ai_1 _18818_ (.B1(_09763_),
    .Y(_09764_),
    .A1(net1131),
    .A2(_09735_));
 sg13g2_buf_1 _18819_ (.A(net260),
    .X(_09765_));
 sg13g2_nor3_1 _18820_ (.A(_09765_),
    .B(_08616_),
    .C(_09735_),
    .Y(_09766_));
 sg13g2_a221oi_1 _18821_ (.B2(_09765_),
    .C1(_09766_),
    .B1(_09764_),
    .A1(_09757_),
    .Y(_09767_),
    .A2(_09758_));
 sg13g2_a21oi_1 _18822_ (.A1(_09756_),
    .A2(_09767_),
    .Y(_09768_),
    .B1(net102));
 sg13g2_xnor2_1 _18823_ (.Y(_09769_),
    .A(_09659_),
    .B(_08924_));
 sg13g2_xnor2_1 _18824_ (.Y(_09770_),
    .A(net283),
    .B(_09769_));
 sg13g2_xnor2_1 _18825_ (.Y(_09771_),
    .A(_09751_),
    .B(_09770_));
 sg13g2_a21oi_1 _18826_ (.A1(_05814_),
    .A2(_09771_),
    .Y(_09772_),
    .B1(_08990_));
 sg13g2_or4_1 _18827_ (.A(net1057),
    .B(_09524_),
    .C(_09768_),
    .D(_09772_),
    .X(_09773_));
 sg13g2_o21ai_1 _18828_ (.B1(_09773_),
    .Y(_00378_),
    .A1(net46),
    .A2(_09658_));
 sg13g2_buf_2 _18829_ (.A(_00146_),
    .X(_09774_));
 sg13g2_inv_1 _18830_ (.Y(_09775_),
    .A(_09774_));
 sg13g2_xor2_1 _18831_ (.B(net908),
    .A(_08768_),
    .X(_09776_));
 sg13g2_nor2_1 _18832_ (.A(net544),
    .B(_09776_),
    .Y(_09777_));
 sg13g2_a21oi_1 _18833_ (.A1(net544),
    .A2(_09126_),
    .Y(_09778_),
    .B1(_09777_));
 sg13g2_a22oi_1 _18834_ (.Y(_09779_),
    .B1(_09778_),
    .B2(net146),
    .A2(net265),
    .A1(_09775_));
 sg13g2_nor2_1 _18835_ (.A(_09527_),
    .B(net285),
    .Y(_09780_));
 sg13g2_a21oi_1 _18836_ (.A1(_09124_),
    .A2(_09780_),
    .Y(_09781_),
    .B1(net144));
 sg13g2_a21oi_1 _18837_ (.A1(net144),
    .A2(_09779_),
    .Y(_09782_),
    .B1(_09781_));
 sg13g2_buf_1 _18838_ (.A(_00116_),
    .X(_09783_));
 sg13g2_xnor2_1 _18839_ (.Y(_09784_),
    .A(_09732_),
    .B(_09525_));
 sg13g2_xnor2_1 _18840_ (.Y(_09785_),
    .A(_08744_),
    .B(_09784_));
 sg13g2_xnor2_1 _18841_ (.Y(_09786_),
    .A(net566),
    .B(_09785_));
 sg13g2_nor4_1 _18842_ (.A(_09077_),
    .B(_09783_),
    .C(_08967_),
    .D(_09786_),
    .Y(_09787_));
 sg13g2_xnor2_1 _18843_ (.Y(_09788_),
    .A(_09697_),
    .B(net1129));
 sg13g2_xnor2_1 _18844_ (.Y(_09789_),
    .A(net909),
    .B(_09788_));
 sg13g2_xnor2_1 _18845_ (.Y(_09790_),
    .A(_09786_),
    .B(_09789_));
 sg13g2_nor2_1 _18846_ (.A(net275),
    .B(_09790_),
    .Y(_09791_));
 sg13g2_nor4_1 _18847_ (.A(net125),
    .B(_09782_),
    .C(_09787_),
    .D(_09791_),
    .Y(_09792_));
 sg13g2_o21ai_1 _18848_ (.B1(_09557_),
    .Y(_09793_),
    .A1(net260),
    .A2(net265));
 sg13g2_nor3_1 _18849_ (.A(net536),
    .B(net264),
    .C(net279),
    .Y(_09794_));
 sg13g2_a21oi_1 _18850_ (.A1(_09774_),
    .A2(_09793_),
    .Y(_09795_),
    .B1(_09794_));
 sg13g2_nor3_1 _18851_ (.A(_09774_),
    .B(net543),
    .C(_08763_),
    .Y(_09796_));
 sg13g2_nor3_1 _18852_ (.A(_08662_),
    .B(net265),
    .C(_09796_),
    .Y(_09797_));
 sg13g2_a21o_1 _18853_ (.A2(_09542_),
    .A1(_09775_),
    .B1(_09797_),
    .X(_09798_));
 sg13g2_buf_1 _18854_ (.A(net543),
    .X(_09799_));
 sg13g2_nand2_1 _18855_ (.Y(_09800_),
    .A(_09775_),
    .B(_09799_));
 sg13g2_nor2_1 _18856_ (.A(_09775_),
    .B(net536),
    .Y(_09801_));
 sg13g2_o21ai_1 _18857_ (.B1(_09801_),
    .Y(_09802_),
    .A1(_09550_),
    .A2(_09780_));
 sg13g2_o21ai_1 _18858_ (.B1(_09802_),
    .Y(_09803_),
    .A1(_08770_),
    .A2(_09800_));
 sg13g2_and2_1 _18859_ (.A(net878),
    .B(_09525_),
    .X(_09804_));
 sg13g2_buf_1 _18860_ (.A(_09804_),
    .X(_09805_));
 sg13g2_a21oi_1 _18861_ (.A1(_08805_),
    .A2(_09805_),
    .Y(_09806_),
    .B1(_09794_));
 sg13g2_nor2_1 _18862_ (.A(net280),
    .B(_09806_),
    .Y(_09807_));
 sg13g2_a221oi_1 _18863_ (.B2(net281),
    .C1(_09807_),
    .B1(_09803_),
    .A1(net260),
    .Y(_09808_),
    .A2(_09798_));
 sg13g2_o21ai_1 _18864_ (.B1(_09808_),
    .Y(_09809_),
    .A1(net146),
    .A2(_09795_));
 sg13g2_nand2_1 _18865_ (.Y(_09810_),
    .A(net1119),
    .B(_08611_));
 sg13g2_xnor2_1 _18866_ (.Y(_09811_),
    .A(net556),
    .B(_09786_));
 sg13g2_inv_1 _18867_ (.Y(_09812_),
    .A(_09783_));
 sg13g2_nand2_1 _18868_ (.Y(_09813_),
    .A(_09812_),
    .B(net568));
 sg13g2_o21ai_1 _18869_ (.B1(_09813_),
    .Y(_09814_),
    .A1(_09077_),
    .A2(_09786_));
 sg13g2_a21oi_1 _18870_ (.A1(_09810_),
    .A2(_09811_),
    .Y(_09815_),
    .B1(_09814_));
 sg13g2_xor2_1 _18871_ (.B(_09815_),
    .A(_09809_),
    .X(_09816_));
 sg13g2_a22oi_1 _18872_ (.Y(_09817_),
    .B1(_09792_),
    .B2(_09816_),
    .A2(net72),
    .A1(net275));
 sg13g2_buf_1 _18873_ (.A(_06110_),
    .X(_09818_));
 sg13g2_a221oi_1 _18874_ (.B2(_09817_),
    .C1(net533),
    .B1(_09617_),
    .A1(net24),
    .Y(_00379_),
    .A2(_09616_));
 sg13g2_nor2_1 _18875_ (.A(_09544_),
    .B(net897),
    .Y(_09819_));
 sg13g2_nand2b_1 _18876_ (.Y(_09820_),
    .B(_09819_),
    .A_N(net535));
 sg13g2_nor2_1 _18877_ (.A(net544),
    .B(_09034_),
    .Y(_09821_));
 sg13g2_nor2_1 _18878_ (.A(net535),
    .B(_09821_),
    .Y(_09822_));
 sg13g2_o21ai_1 _18879_ (.B1(_09774_),
    .Y(_09823_),
    .A1(_09819_),
    .A2(_09822_));
 sg13g2_a21oi_1 _18880_ (.A1(_09820_),
    .A2(_09823_),
    .Y(_09824_),
    .B1(net146));
 sg13g2_nand2_1 _18881_ (.Y(_09825_),
    .A(net264),
    .B(net897));
 sg13g2_nor2_1 _18882_ (.A(_09774_),
    .B(_09825_),
    .Y(_09826_));
 sg13g2_nor3_1 _18883_ (.A(_09774_),
    .B(net264),
    .C(net554),
    .Y(_09827_));
 sg13g2_nor3_1 _18884_ (.A(_08662_),
    .B(_09821_),
    .C(_09827_),
    .Y(_09828_));
 sg13g2_o21ai_1 _18885_ (.B1(_09743_),
    .Y(_09829_),
    .A1(_09826_),
    .A2(_09828_));
 sg13g2_nand2_1 _18886_ (.Y(_09830_),
    .A(_09775_),
    .B(net286));
 sg13g2_nor2_1 _18887_ (.A(_09544_),
    .B(net555),
    .Y(_09831_));
 sg13g2_o21ai_1 _18888_ (.B1(_09801_),
    .Y(_09832_),
    .A1(_09780_),
    .A2(_09831_));
 sg13g2_o21ai_1 _18889_ (.B1(_09832_),
    .Y(_09833_),
    .A1(_09825_),
    .A2(_09830_));
 sg13g2_nand3_1 _18890_ (.B(net286),
    .C(_09805_),
    .A(net554),
    .Y(_09834_));
 sg13g2_a21oi_1 _18891_ (.A1(_09820_),
    .A2(_09834_),
    .Y(_09835_),
    .B1(net280));
 sg13g2_a21oi_1 _18892_ (.A1(net280),
    .A2(_09833_),
    .Y(_09836_),
    .B1(_09835_));
 sg13g2_nand3b_1 _18893_ (.B(_09829_),
    .C(_09836_),
    .Y(_09837_),
    .A_N(_09824_));
 sg13g2_xor2_1 _18894_ (.B(_09784_),
    .A(_09748_),
    .X(_09838_));
 sg13g2_xnor2_1 _18895_ (.Y(_09839_),
    .A(net285),
    .B(_09838_));
 sg13g2_xnor2_1 _18896_ (.Y(_09840_),
    .A(_08812_),
    .B(_09839_));
 sg13g2_o21ai_1 _18897_ (.B1(_09536_),
    .Y(_09841_),
    .A1(net561),
    .A2(_09839_));
 sg13g2_a21oi_1 _18898_ (.A1(_09534_),
    .A2(_09840_),
    .Y(_09842_),
    .B1(_09841_));
 sg13g2_xnor2_1 _18899_ (.Y(_09843_),
    .A(_09837_),
    .B(_09842_));
 sg13g2_xnor2_1 _18900_ (.Y(_09844_),
    .A(_09611_),
    .B(_09839_));
 sg13g2_nor4_1 _18901_ (.A(_09533_),
    .B(net561),
    .C(_09604_),
    .D(_09839_),
    .Y(_09845_));
 sg13g2_nand2_1 _18902_ (.Y(_09846_),
    .A(_09545_),
    .B(_09748_));
 sg13g2_o21ai_1 _18903_ (.B1(_09846_),
    .Y(_09847_),
    .A1(net259),
    .A2(_09039_));
 sg13g2_a21oi_1 _18904_ (.A1(net146),
    .A2(_09847_),
    .Y(_09848_),
    .B1(_09826_));
 sg13g2_nor2b_1 _18905_ (.A(_09848_),
    .B_N(_09743_),
    .Y(_09849_));
 sg13g2_nor3_1 _18906_ (.A(net144),
    .B(_08662_),
    .C(_09825_),
    .Y(_09850_));
 sg13g2_nor4_1 _18907_ (.A(net170),
    .B(_09845_),
    .C(_09849_),
    .D(_09850_),
    .Y(_09851_));
 sg13g2_o21ai_1 _18908_ (.B1(_09851_),
    .Y(_09852_),
    .A1(net145),
    .A2(_09844_));
 sg13g2_or2_1 _18909_ (.X(_09853_),
    .B(_09852_),
    .A(_09843_));
 sg13g2_a22oi_1 _18910_ (.Y(_09854_),
    .B1(net76),
    .B2(_09616_),
    .A2(net72),
    .A1(net145));
 sg13g2_a221oi_1 _18911_ (.B2(_09854_),
    .C1(net533),
    .B1(_09853_),
    .A1(_06471_),
    .Y(_00380_),
    .A2(_09616_));
 sg13g2_or4_1 _18912_ (.A(_07972_),
    .B(_06472_),
    .C(_02021_),
    .D(_09522_),
    .X(_09855_));
 sg13g2_buf_1 _18913_ (.A(_09855_),
    .X(_09856_));
 sg13g2_buf_1 _18914_ (.A(\grid.cell_21_0.sw ),
    .X(_09857_));
 sg13g2_xor2_1 _18915_ (.B(_09525_),
    .A(net1118),
    .X(_09858_));
 sg13g2_buf_2 _18916_ (.A(_09858_),
    .X(_09859_));
 sg13g2_buf_2 _18917_ (.A(\grid.cell_21_0.se ),
    .X(_09860_));
 sg13g2_xnor2_1 _18918_ (.Y(_09861_),
    .A(_08739_),
    .B(_09860_));
 sg13g2_xor2_1 _18919_ (.B(_09861_),
    .A(_09859_),
    .X(_09862_));
 sg13g2_xnor2_1 _18920_ (.Y(_09863_),
    .A(net563),
    .B(_09862_));
 sg13g2_xnor2_1 _18921_ (.Y(_09864_),
    .A(_09561_),
    .B(_09863_));
 sg13g2_buf_2 _18922_ (.A(\grid.cell_21_0.s ),
    .X(_09865_));
 sg13g2_xor2_1 _18923_ (.B(_09865_),
    .A(net904),
    .X(_09866_));
 sg13g2_xor2_1 _18924_ (.B(_09866_),
    .A(_09864_),
    .X(_09867_));
 sg13g2_nor2_1 _18925_ (.A(net883),
    .B(_09867_),
    .Y(_09868_));
 sg13g2_buf_1 _18926_ (.A(_09860_),
    .X(_09869_));
 sg13g2_buf_1 _18927_ (.A(net877),
    .X(_09870_));
 sg13g2_buf_1 _18928_ (.A(net1118),
    .X(_09871_));
 sg13g2_buf_1 _18929_ (.A(net876),
    .X(_09872_));
 sg13g2_nand2b_1 _18930_ (.Y(_09873_),
    .B(_09550_),
    .A_N(net531));
 sg13g2_and2_1 _18931_ (.A(net1118),
    .B(_09525_),
    .X(_09874_));
 sg13g2_buf_2 _18932_ (.A(_09874_),
    .X(_09875_));
 sg13g2_nand3_1 _18933_ (.B(net1130),
    .C(_09875_),
    .A(_09869_),
    .Y(_09876_));
 sg13g2_o21ai_1 _18934_ (.B1(_09876_),
    .Y(_09877_),
    .A1(net532),
    .A2(_09873_));
 sg13g2_nand2b_1 _18935_ (.Y(_09878_),
    .B(net884),
    .A_N(net1118));
 sg13g2_buf_1 _18936_ (.A(_09878_),
    .X(_09879_));
 sg13g2_buf_1 _18937_ (.A(net876),
    .X(_09880_));
 sg13g2_nand2b_1 _18938_ (.Y(_09881_),
    .B(_09540_),
    .A_N(net1130));
 sg13g2_nand2_1 _18939_ (.Y(_09882_),
    .A(net530),
    .B(_09881_));
 sg13g2_a21oi_1 _18940_ (.A1(_09879_),
    .A2(_09882_),
    .Y(_09883_),
    .B1(net279));
 sg13g2_nand2b_1 _18941_ (.Y(_09884_),
    .B(net530),
    .A_N(net543));
 sg13g2_nand2b_1 _18942_ (.Y(_09885_),
    .B(net563),
    .A_N(net530));
 sg13g2_a21oi_1 _18943_ (.A1(_09884_),
    .A2(_09885_),
    .Y(_09886_),
    .B1(net906));
 sg13g2_nor3_1 _18944_ (.A(net531),
    .B(net264),
    .C(net1130),
    .Y(_09887_));
 sg13g2_or3_1 _18945_ (.A(_09883_),
    .B(_09886_),
    .C(_09887_),
    .X(_09888_));
 sg13g2_buf_1 _18946_ (.A(net877),
    .X(_09889_));
 sg13g2_o21ai_1 _18947_ (.B1(_09552_),
    .Y(_09890_),
    .A1(net543),
    .A2(_08907_));
 sg13g2_or2_1 _18948_ (.X(_09891_),
    .B(_09525_),
    .A(_09857_));
 sg13g2_buf_1 _18949_ (.A(_09891_),
    .X(_09892_));
 sg13g2_nor2b_1 _18950_ (.A(_08739_),
    .B_N(net563),
    .Y(_09893_));
 sg13g2_nor2_1 _18951_ (.A(net531),
    .B(_09881_),
    .Y(_09894_));
 sg13g2_a221oi_1 _18952_ (.B2(_09893_),
    .C1(_09894_),
    .B1(_09892_),
    .A1(net531),
    .Y(_09895_),
    .A2(_09890_));
 sg13g2_nor2_1 _18953_ (.A(net529),
    .B(_09895_),
    .Y(_09896_));
 sg13g2_a221oi_1 _18954_ (.B2(net529),
    .C1(_09896_),
    .B1(_09888_),
    .A1(net562),
    .Y(_09897_),
    .A2(_09877_));
 sg13g2_inv_1 _18955_ (.Y(_09898_),
    .A(_08811_));
 sg13g2_buf_1 _18956_ (.A(_00203_),
    .X(_09899_));
 sg13g2_nand2_1 _18957_ (.Y(_09900_),
    .A(_09898_),
    .B(net1117));
 sg13g2_nor2_1 _18958_ (.A(_09898_),
    .B(net1117),
    .Y(_09901_));
 sg13g2_a221oi_1 _18959_ (.B2(_09900_),
    .C1(_09901_),
    .B1(_09864_),
    .A1(_09621_),
    .Y(_09902_),
    .A2(_09863_));
 sg13g2_xnor2_1 _18960_ (.Y(_09903_),
    .A(_09897_),
    .B(_09902_));
 sg13g2_mux2_1 _18961_ (.A0(_09859_),
    .A1(_09875_),
    .S(net565),
    .X(_09904_));
 sg13g2_a22oi_1 _18962_ (.Y(_09905_),
    .B1(_09904_),
    .B2(net145),
    .A2(_09875_),
    .A1(_09629_));
 sg13g2_nand2b_1 _18963_ (.Y(_09906_),
    .B(net529),
    .A_N(_09905_));
 sg13g2_nor2b_1 _18964_ (.A(net877),
    .B_N(net1118),
    .Y(_09907_));
 sg13g2_nand3_1 _18965_ (.B(net265),
    .C(_09907_),
    .A(net562),
    .Y(_09908_));
 sg13g2_nand3_1 _18966_ (.B(_09906_),
    .C(_09908_),
    .A(net118),
    .Y(_09909_));
 sg13g2_inv_1 _18967_ (.Y(_09910_),
    .A(net1117));
 sg13g2_xnor2_1 _18968_ (.Y(_09911_),
    .A(net904),
    .B(net541));
 sg13g2_and4_1 _18969_ (.A(_09910_),
    .B(_09621_),
    .C(_09863_),
    .D(_09911_),
    .X(_09912_));
 sg13g2_nor4_1 _18970_ (.A(_09868_),
    .B(_09903_),
    .C(_09909_),
    .D(_09912_),
    .Y(_09913_));
 sg13g2_a21oi_1 _18971_ (.A1(net883),
    .A2(net73),
    .Y(_09914_),
    .B1(_09913_));
 sg13g2_o21ai_1 _18972_ (.B1(net334),
    .Y(_09915_),
    .A1(net40),
    .A2(net57));
 sg13g2_a21oi_1 _18973_ (.A1(net57),
    .A2(_09914_),
    .Y(_00381_),
    .B1(_09915_));
 sg13g2_buf_1 _18974_ (.A(net320),
    .X(_09916_));
 sg13g2_nor4_1 _18975_ (.A(_07972_),
    .B(net143),
    .C(net375),
    .D(_09522_),
    .Y(_09917_));
 sg13g2_buf_1 _18976_ (.A(_09917_),
    .X(_09918_));
 sg13g2_nand2_1 _18977_ (.Y(_09919_),
    .A(net42),
    .B(net56));
 sg13g2_buf_2 _18978_ (.A(\grid.cell_21_1.se ),
    .X(_09920_));
 sg13g2_xnor2_1 _18979_ (.Y(_09921_),
    .A(_08823_),
    .B(_09920_));
 sg13g2_xnor2_1 _18980_ (.Y(_09922_),
    .A(_09586_),
    .B(_09921_));
 sg13g2_xor2_1 _18981_ (.B(_09922_),
    .A(_09861_),
    .X(_09923_));
 sg13g2_nor2_1 _18982_ (.A(_09533_),
    .B(_09923_),
    .Y(_09924_));
 sg13g2_xor2_1 _18983_ (.B(_09920_),
    .A(net1122),
    .X(_09925_));
 sg13g2_xor2_1 _18984_ (.B(_08823_),
    .A(_08739_),
    .X(_09926_));
 sg13g2_xnor2_1 _18985_ (.Y(_09927_),
    .A(_09579_),
    .B(_09860_));
 sg13g2_xnor2_1 _18986_ (.Y(_09928_),
    .A(_09926_),
    .B(_09927_));
 sg13g2_xnor2_1 _18987_ (.Y(_09929_),
    .A(_09925_),
    .B(_09928_));
 sg13g2_buf_1 _18988_ (.A(_09929_),
    .X(_09930_));
 sg13g2_o21ai_1 _18989_ (.B1(_09930_),
    .Y(_09931_),
    .A1(net1117),
    .A2(_09924_));
 sg13g2_nor2_1 _18990_ (.A(net1117),
    .B(_09930_),
    .Y(_09932_));
 sg13g2_a21o_1 _18991_ (.A2(_09930_),
    .A1(_09898_),
    .B1(net1117),
    .X(_09933_));
 sg13g2_mux2_1 _18992_ (.A0(_09932_),
    .A1(_09933_),
    .S(_09924_),
    .X(_09934_));
 sg13g2_a21o_1 _18993_ (.A2(_09931_),
    .A1(net904),
    .B1(_09934_),
    .X(_09935_));
 sg13g2_buf_1 _18994_ (.A(_09920_),
    .X(_09936_));
 sg13g2_inv_1 _18995_ (.Y(_09937_),
    .A(net875));
 sg13g2_buf_1 _18996_ (.A(_09937_),
    .X(_09938_));
 sg13g2_nor2_1 _18997_ (.A(net539),
    .B(net258),
    .Y(_09939_));
 sg13g2_nand2_1 _18998_ (.Y(_09940_),
    .A(net906),
    .B(_09925_));
 sg13g2_o21ai_1 _18999_ (.B1(_09940_),
    .Y(_09941_),
    .A1(net560),
    .A2(_09939_));
 sg13g2_nand2_1 _19000_ (.Y(_09942_),
    .A(_08739_),
    .B(net903));
 sg13g2_buf_1 _19001_ (.A(net875),
    .X(_09943_));
 sg13g2_nor2_2 _19002_ (.A(net882),
    .B(net528),
    .Y(_09944_));
 sg13g2_a22oi_1 _19003_ (.Y(_09945_),
    .B1(_09942_),
    .B2(_09944_),
    .A2(_09941_),
    .A1(net901));
 sg13g2_nand2_1 _19004_ (.Y(_09946_),
    .A(net901),
    .B(_09944_));
 sg13g2_inv_1 _19005_ (.Y(_09947_),
    .A(_09869_));
 sg13g2_o21ai_1 _19006_ (.B1(net560),
    .Y(_09948_),
    .A1(net565),
    .A2(_09947_));
 sg13g2_nand2b_1 _19007_ (.Y(_09949_),
    .B(_09948_),
    .A_N(_09946_));
 sg13g2_o21ai_1 _19008_ (.B1(_09949_),
    .Y(_09950_),
    .A1(_09889_),
    .A2(_09945_));
 sg13g2_nand2b_1 _19009_ (.Y(_09951_),
    .B(net875),
    .A_N(net1130));
 sg13g2_o21ai_1 _19010_ (.B1(_09951_),
    .Y(_09952_),
    .A1(net875),
    .A2(_09942_));
 sg13g2_nor2_1 _19011_ (.A(net875),
    .B(net1130),
    .Y(_09953_));
 sg13g2_nor3_1 _19012_ (.A(net882),
    .B(_09942_),
    .C(_09953_),
    .Y(_09954_));
 sg13g2_a21oi_1 _19013_ (.A1(net882),
    .A2(_09952_),
    .Y(_09955_),
    .B1(_09954_));
 sg13g2_nor2b_1 _19014_ (.A(net875),
    .B_N(net1130),
    .Y(_09956_));
 sg13g2_a21oi_1 _19015_ (.A1(_09587_),
    .A2(_09951_),
    .Y(_09957_),
    .B1(_09956_));
 sg13g2_nor2_1 _19016_ (.A(net903),
    .B(_09957_),
    .Y(_09958_));
 sg13g2_nand2_1 _19017_ (.Y(_09959_),
    .A(net875),
    .B(net1130));
 sg13g2_o21ai_1 _19018_ (.B1(net1122),
    .Y(_09960_),
    .A1(_09936_),
    .A2(net1130));
 sg13g2_a21oi_1 _19019_ (.A1(_09959_),
    .A2(_09960_),
    .Y(_09961_),
    .B1(_09942_));
 sg13g2_nor3_1 _19020_ (.A(net532),
    .B(_09958_),
    .C(_09961_),
    .Y(_09962_));
 sg13g2_a21oi_1 _19021_ (.A1(_09889_),
    .A2(_09955_),
    .Y(_09963_),
    .B1(_09962_));
 sg13g2_nand2_1 _19022_ (.Y(_09964_),
    .A(_09947_),
    .B(_09944_));
 sg13g2_nand3_1 _19023_ (.B(net560),
    .C(_09939_),
    .A(net532),
    .Y(_09965_));
 sg13g2_a21oi_1 _19024_ (.A1(_09964_),
    .A2(_09965_),
    .Y(_09966_),
    .B1(net562));
 sg13g2_nor2_1 _19025_ (.A(net278),
    .B(_09946_),
    .Y(_09967_));
 sg13g2_nor4_1 _19026_ (.A(_09924_),
    .B(_09963_),
    .C(_09966_),
    .D(_09967_),
    .Y(_09968_));
 sg13g2_nand2_1 _19027_ (.Y(_09969_),
    .A(_09899_),
    .B(_09930_));
 sg13g2_o21ai_1 _19028_ (.B1(_09969_),
    .Y(_09970_),
    .A1(net904),
    .A2(_09932_));
 sg13g2_a221oi_1 _19029_ (.B2(_09970_),
    .C1(net100),
    .B1(_09968_),
    .A1(_09935_),
    .Y(_09971_),
    .A2(_09950_));
 sg13g2_xnor2_1 _19030_ (.Y(_09972_),
    .A(_09866_),
    .B(_09930_));
 sg13g2_a21oi_1 _19031_ (.A1(net109),
    .A2(_09972_),
    .Y(_09973_),
    .B1(_09602_));
 sg13g2_or3_1 _19032_ (.A(net56),
    .B(_09971_),
    .C(_09973_),
    .X(_09974_));
 sg13g2_a21oi_1 _19033_ (.A1(_09919_),
    .A2(_09974_),
    .Y(_00382_),
    .B1(net305));
 sg13g2_nand2_1 _19034_ (.Y(_09975_),
    .A(net33),
    .B(net56));
 sg13g2_buf_1 _19035_ (.A(net528),
    .X(_09976_));
 sg13g2_buf_2 _19036_ (.A(\grid.cell_21_2.se ),
    .X(_09977_));
 sg13g2_xor2_1 _19037_ (.B(net881),
    .A(_09977_),
    .X(_09978_));
 sg13g2_and2_1 _19038_ (.A(net903),
    .B(_09978_),
    .X(_09979_));
 sg13g2_buf_1 _19039_ (.A(_09977_),
    .X(_09980_));
 sg13g2_nand2_1 _19040_ (.Y(_09981_),
    .A(net874),
    .B(net881));
 sg13g2_nor2_1 _19041_ (.A(net903),
    .B(_09981_),
    .Y(_09982_));
 sg13g2_o21ai_1 _19042_ (.B1(net276),
    .Y(_09983_),
    .A1(_09979_),
    .A2(_09982_));
 sg13g2_or2_1 _19043_ (.X(_09984_),
    .B(_09981_),
    .A(_08931_));
 sg13g2_nand3_1 _19044_ (.B(_09983_),
    .C(_09984_),
    .A(net257),
    .Y(_09985_));
 sg13g2_buf_1 _19045_ (.A(net874),
    .X(_09986_));
 sg13g2_buf_1 _19046_ (.A(_09986_),
    .X(_09987_));
 sg13g2_nand2_1 _19047_ (.Y(_09988_),
    .A(net560),
    .B(net256));
 sg13g2_o21ai_1 _19048_ (.B1(_09938_),
    .Y(_09989_),
    .A1(_09648_),
    .A2(_09988_));
 sg13g2_buf_1 _19049_ (.A(_00202_),
    .X(_09990_));
 sg13g2_buf_1 _19050_ (.A(_09990_),
    .X(_09991_));
 sg13g2_xor2_1 _19051_ (.B(_09977_),
    .A(_09528_),
    .X(_09992_));
 sg13g2_xnor2_1 _19052_ (.Y(_09993_),
    .A(_09921_),
    .B(_09992_));
 sg13g2_xnor2_1 _19053_ (.Y(_09994_),
    .A(_09623_),
    .B(_09993_));
 sg13g2_buf_1 _19054_ (.A(_09994_),
    .X(_09995_));
 sg13g2_nand2_1 _19055_ (.Y(_09996_),
    .A(net873),
    .B(_09995_));
 sg13g2_o21ai_1 _19056_ (.B1(net565),
    .Y(_09997_),
    .A1(net873),
    .A2(_09995_));
 sg13g2_xor2_1 _19057_ (.B(_09978_),
    .A(net902),
    .X(_09998_));
 sg13g2_xor2_1 _19058_ (.B(_09998_),
    .A(_09921_),
    .X(_09999_));
 sg13g2_nor2_1 _19059_ (.A(_09620_),
    .B(_09999_),
    .Y(_10000_));
 sg13g2_a221oi_1 _19060_ (.B2(_09997_),
    .C1(_10000_),
    .B1(_09996_),
    .A1(_09985_),
    .Y(_10001_),
    .A2(_09989_));
 sg13g2_o21ai_1 _19061_ (.B1(_09995_),
    .Y(_10002_),
    .A1(net873),
    .A2(_10000_));
 sg13g2_nor2_1 _19062_ (.A(_09991_),
    .B(_09995_),
    .Y(_10003_));
 sg13g2_a21o_1 _19063_ (.A2(_09995_),
    .A1(net565),
    .B1(net873),
    .X(_10004_));
 sg13g2_mux2_1 _19064_ (.A0(_10003_),
    .A1(_10004_),
    .S(_10000_),
    .X(_10005_));
 sg13g2_a21o_1 _19065_ (.A2(_10002_),
    .A1(net562),
    .B1(_10005_),
    .X(_10006_));
 sg13g2_a21oi_1 _19066_ (.A1(net527),
    .A2(net540),
    .Y(_10007_),
    .B1(net902));
 sg13g2_or2_1 _19067_ (.X(_10008_),
    .B(_10007_),
    .A(_09979_));
 sg13g2_nand2_1 _19068_ (.Y(_10009_),
    .A(net560),
    .B(net276));
 sg13g2_nor2_1 _19069_ (.A(_09986_),
    .B(net263),
    .Y(_10010_));
 sg13g2_a22oi_1 _19070_ (.Y(_10011_),
    .B1(_10009_),
    .B2(_10010_),
    .A2(_10008_),
    .A1(_08931_));
 sg13g2_o21ai_1 _19071_ (.B1(net276),
    .Y(_10012_),
    .A1(_08844_),
    .A2(_09938_));
 sg13g2_nand3_1 _19072_ (.B(_10012_),
    .C(_10010_),
    .A(_08931_),
    .Y(_10013_));
 sg13g2_o21ai_1 _19073_ (.B1(_10013_),
    .Y(_10014_),
    .A1(net257),
    .A2(_10011_));
 sg13g2_mux2_1 _19074_ (.A0(_10001_),
    .A1(_10006_),
    .S(_10014_),
    .X(_10015_));
 sg13g2_xor2_1 _19075_ (.B(_09995_),
    .A(_09861_),
    .X(_10016_));
 sg13g2_a21oi_1 _19076_ (.A1(net116),
    .A2(_10016_),
    .Y(_10017_),
    .B1(_09600_));
 sg13g2_nor2_1 _19077_ (.A(net56),
    .B(_10017_),
    .Y(_10018_));
 sg13g2_o21ai_1 _19078_ (.B1(_10018_),
    .Y(_10019_),
    .A1(net74),
    .A2(_10015_));
 sg13g2_a21oi_1 _19079_ (.A1(_09975_),
    .A2(_10019_),
    .Y(_00383_),
    .B1(net305));
 sg13g2_nand2_1 _19080_ (.Y(_10020_),
    .A(_06621_),
    .B(net56));
 sg13g2_buf_1 _19081_ (.A(\grid.cell_21_3.se ),
    .X(_10021_));
 sg13g2_buf_1 _19082_ (.A(net1116),
    .X(_10022_));
 sg13g2_inv_2 _19083_ (.Y(_10023_),
    .A(_10022_));
 sg13g2_xnor2_1 _19084_ (.Y(_10024_),
    .A(net880),
    .B(net559));
 sg13g2_a21oi_1 _19085_ (.A1(net538),
    .A2(net559),
    .Y(_10025_),
    .B1(net527));
 sg13g2_a21oi_1 _19086_ (.A1(_09987_),
    .A2(_10024_),
    .Y(_10026_),
    .B1(_10025_));
 sg13g2_inv_1 _19087_ (.Y(_10027_),
    .A(net527));
 sg13g2_nor2_1 _19088_ (.A(_10027_),
    .B(_09679_),
    .Y(_10028_));
 sg13g2_a22oi_1 _19089_ (.Y(_10029_),
    .B1(_10028_),
    .B2(_09009_),
    .A2(_10026_),
    .A1(net277));
 sg13g2_nor2_1 _19090_ (.A(_10022_),
    .B(_09679_),
    .Y(_10030_));
 sg13g2_nand3_1 _19091_ (.B(_08952_),
    .C(_10030_),
    .A(_09987_),
    .Y(_10031_));
 sg13g2_o21ai_1 _19092_ (.B1(_10031_),
    .Y(_10032_),
    .A1(_10023_),
    .A2(_10029_));
 sg13g2_nor2b_1 _19093_ (.A(_09659_),
    .B_N(net900),
    .Y(_10033_));
 sg13g2_nor2_1 _19094_ (.A(net1116),
    .B(_09977_),
    .Y(_10034_));
 sg13g2_nor2b_1 _19095_ (.A(net902),
    .B_N(net900),
    .Y(_10035_));
 sg13g2_a221oi_1 _19096_ (.B2(_10034_),
    .C1(_10035_),
    .B1(_10033_),
    .A1(net874),
    .Y(_10036_),
    .A2(_09659_));
 sg13g2_o21ai_1 _19097_ (.B1(net1116),
    .Y(_10037_),
    .A1(_09977_),
    .A2(_09659_));
 sg13g2_and2_1 _19098_ (.A(_08975_),
    .B(_10037_),
    .X(_10038_));
 sg13g2_nor4_1 _19099_ (.A(net1116),
    .B(net874),
    .C(net880),
    .D(_08952_),
    .Y(_10039_));
 sg13g2_a21o_1 _19100_ (.A2(_10038_),
    .A1(_10036_),
    .B1(_10039_),
    .X(_10040_));
 sg13g2_buf_1 _19101_ (.A(_10040_),
    .X(_10041_));
 sg13g2_xor2_1 _19102_ (.B(net902),
    .A(_09980_),
    .X(_10042_));
 sg13g2_xnor2_1 _19103_ (.Y(_10043_),
    .A(_09769_),
    .B(_10042_));
 sg13g2_xnor2_1 _19104_ (.Y(_10044_),
    .A(net872),
    .B(_10043_));
 sg13g2_buf_1 _19105_ (.A(_10044_),
    .X(_10045_));
 sg13g2_buf_1 _19106_ (.A(_00201_),
    .X(_10046_));
 sg13g2_inv_1 _19107_ (.Y(_10047_),
    .A(net1115));
 sg13g2_a21oi_1 _19108_ (.A1(net542),
    .A2(_10045_),
    .Y(_10048_),
    .B1(_10047_));
 sg13g2_nor2_1 _19109_ (.A(_09587_),
    .B(net1115),
    .Y(_10049_));
 sg13g2_a21oi_1 _19110_ (.A1(_10045_),
    .A2(_10049_),
    .Y(_10050_),
    .B1(net278));
 sg13g2_nor3_1 _19111_ (.A(_10041_),
    .B(_10048_),
    .C(_10050_),
    .Y(_10051_));
 sg13g2_nand2_1 _19112_ (.Y(_10052_),
    .A(net1115),
    .B(_00204_));
 sg13g2_nand2_1 _19113_ (.Y(_10053_),
    .A(net539),
    .B(net1115));
 sg13g2_o21ai_1 _19114_ (.B1(_10053_),
    .Y(_10054_),
    .A1(net903),
    .A2(_10049_));
 sg13g2_nand2_1 _19115_ (.Y(_10055_),
    .A(_10045_),
    .B(_10054_));
 sg13g2_o21ai_1 _19116_ (.B1(_10055_),
    .Y(_10056_),
    .A1(net278),
    .A2(_10052_));
 sg13g2_and2_1 _19117_ (.A(_10041_),
    .B(_10056_),
    .X(_10057_));
 sg13g2_nor3_1 _19118_ (.A(net542),
    .B(_10046_),
    .C(net1120),
    .Y(_10058_));
 sg13g2_and3_1 _19119_ (.X(_10059_),
    .A(net542),
    .B(net1120),
    .C(_10041_));
 sg13g2_o21ai_1 _19120_ (.B1(_08844_),
    .Y(_10060_),
    .A1(_10058_),
    .A2(_10059_));
 sg13g2_nand3b_1 _19121_ (.B(net882),
    .C(_10047_),
    .Y(_10061_),
    .A_N(net1120));
 sg13g2_o21ai_1 _19122_ (.B1(_10061_),
    .Y(_10062_),
    .A1(net542),
    .A2(_10041_));
 sg13g2_o21ai_1 _19123_ (.B1(net1120),
    .Y(_10063_),
    .A1(_09599_),
    .A2(_10046_));
 sg13g2_nor2_1 _19124_ (.A(net539),
    .B(_10052_),
    .Y(_10064_));
 sg13g2_mux2_1 _19125_ (.A0(_10063_),
    .A1(_10064_),
    .S(_10041_),
    .X(_10065_));
 sg13g2_a21oi_1 _19126_ (.A1(net278),
    .A2(_10062_),
    .Y(_10066_),
    .B1(_10065_));
 sg13g2_a21oi_1 _19127_ (.A1(_10060_),
    .A2(_10066_),
    .Y(_10067_),
    .B1(_10045_));
 sg13g2_nor4_1 _19128_ (.A(_10032_),
    .B(_10051_),
    .C(_10057_),
    .D(_10067_),
    .Y(_10068_));
 sg13g2_xnor2_1 _19129_ (.Y(_10069_),
    .A(_09922_),
    .B(_10045_));
 sg13g2_a21oi_1 _19130_ (.A1(net116),
    .A2(_10069_),
    .Y(_10070_),
    .B1(net263));
 sg13g2_nor2_1 _19131_ (.A(net56),
    .B(_10070_),
    .Y(_10071_));
 sg13g2_o21ai_1 _19132_ (.B1(_10071_),
    .Y(_10072_),
    .A1(net74),
    .A2(_10068_));
 sg13g2_a21oi_1 _19133_ (.A1(_10020_),
    .A2(_10072_),
    .Y(_00384_),
    .B1(net305));
 sg13g2_nand3_1 _19134_ (.B(net104),
    .C(net57),
    .A(_09662_),
    .Y(_10073_));
 sg13g2_o21ai_1 _19135_ (.B1(_10073_),
    .Y(_10074_),
    .A1(net47),
    .A2(net57));
 sg13g2_buf_1 _19136_ (.A(_00055_),
    .X(_10075_));
 sg13g2_xor2_1 _19137_ (.B(net900),
    .A(net872),
    .X(_10076_));
 sg13g2_buf_1 _19138_ (.A(\grid.cell_21_4.se ),
    .X(_10077_));
 sg13g2_buf_1 _19139_ (.A(_10077_),
    .X(_10078_));
 sg13g2_xnor2_1 _19140_ (.Y(_10079_),
    .A(net871),
    .B(_09788_));
 sg13g2_xnor2_1 _19141_ (.Y(_10080_),
    .A(_10076_),
    .B(_10079_));
 sg13g2_nor4_1 _19142_ (.A(_09706_),
    .B(_10075_),
    .C(_09623_),
    .D(_10080_),
    .Y(_10081_));
 sg13g2_buf_1 _19143_ (.A(net871),
    .X(_10082_));
 sg13g2_buf_1 _19144_ (.A(net526),
    .X(_10083_));
 sg13g2_nand2_1 _19145_ (.Y(_10084_),
    .A(net872),
    .B(net879));
 sg13g2_nor2_1 _19146_ (.A(net558),
    .B(_10084_),
    .Y(_10085_));
 sg13g2_xnor2_1 _19147_ (.Y(_10086_),
    .A(net872),
    .B(net879));
 sg13g2_nor2_1 _19148_ (.A(_08942_),
    .B(_10086_),
    .Y(_10087_));
 sg13g2_o21ai_1 _19149_ (.B1(net556),
    .Y(_10088_),
    .A1(_10085_),
    .A2(_10087_));
 sg13g2_o21ai_1 _19150_ (.B1(_10088_),
    .Y(_10089_),
    .A1(_09019_),
    .A2(_10084_));
 sg13g2_nand2_1 _19151_ (.Y(_10090_),
    .A(net255),
    .B(_10089_));
 sg13g2_nand2_1 _19152_ (.Y(_10091_),
    .A(net899),
    .B(net277));
 sg13g2_or3_1 _19153_ (.A(net255),
    .B(_10091_),
    .C(_10084_),
    .X(_10092_));
 sg13g2_nand4_1 _19154_ (.B(_09856_),
    .C(_10090_),
    .A(net1060),
    .Y(_10093_),
    .D(_10092_));
 sg13g2_xnor2_1 _19155_ (.Y(_10094_),
    .A(_09998_),
    .B(_10080_));
 sg13g2_a21oi_1 _19156_ (.A1(net70),
    .A2(_10094_),
    .Y(_10095_),
    .B1(net262));
 sg13g2_buf_1 _19157_ (.A(net872),
    .X(_10096_));
 sg13g2_buf_1 _19158_ (.A(_10096_),
    .X(_10097_));
 sg13g2_nor4_1 _19159_ (.A(net526),
    .B(net525),
    .C(net537),
    .D(_08985_),
    .Y(_10098_));
 sg13g2_a221oi_1 _19160_ (.B2(_08942_),
    .C1(_10098_),
    .B1(net556),
    .A1(net254),
    .Y(_10099_),
    .A2(net261));
 sg13g2_o21ai_1 _19161_ (.B1(net255),
    .Y(_10100_),
    .A1(_10096_),
    .A2(net537));
 sg13g2_and2_1 _19162_ (.A(_09019_),
    .B(_10100_),
    .X(_10101_));
 sg13g2_nor3_1 _19163_ (.A(_10083_),
    .B(_10097_),
    .C(net261),
    .Y(_10102_));
 sg13g2_a22oi_1 _19164_ (.Y(_10103_),
    .B1(_10102_),
    .B2(_10091_),
    .A2(_10101_),
    .A1(_10099_));
 sg13g2_nand2b_1 _19165_ (.Y(_10104_),
    .B(_10075_),
    .A_N(net276));
 sg13g2_xnor2_1 _19166_ (.Y(_10105_),
    .A(net263),
    .B(_10080_));
 sg13g2_inv_1 _19167_ (.Y(_10106_),
    .A(_10075_));
 sg13g2_nand2_1 _19168_ (.Y(_10107_),
    .A(_10106_),
    .B(net276));
 sg13g2_o21ai_1 _19169_ (.B1(_10107_),
    .Y(_10108_),
    .A1(_09706_),
    .A2(_10080_));
 sg13g2_a21oi_1 _19170_ (.A1(_10104_),
    .A2(_10105_),
    .Y(_10109_),
    .B1(_10108_));
 sg13g2_xor2_1 _19171_ (.B(_10109_),
    .A(_10103_),
    .X(_10110_));
 sg13g2_nor4_1 _19172_ (.A(_10081_),
    .B(_10093_),
    .C(_10095_),
    .D(_10110_),
    .Y(_10111_));
 sg13g2_a21o_1 _19173_ (.A2(_10074_),
    .A1(net317),
    .B1(_10111_),
    .X(_00385_));
 sg13g2_nand2_1 _19174_ (.Y(_10112_),
    .A(_06330_),
    .B(_09918_));
 sg13g2_buf_2 _19175_ (.A(\grid.cell_21_5.se ),
    .X(_10113_));
 sg13g2_buf_1 _19176_ (.A(_10113_),
    .X(_10114_));
 sg13g2_buf_1 _19177_ (.A(_10114_),
    .X(_10115_));
 sg13g2_buf_1 _19178_ (.A(net524),
    .X(_10116_));
 sg13g2_nor4_1 _19179_ (.A(net253),
    .B(net526),
    .C(net535),
    .D(net555),
    .Y(_10117_));
 sg13g2_nand2_1 _19180_ (.Y(_10118_),
    .A(net526),
    .B(net536));
 sg13g2_nand2_1 _19181_ (.Y(_10119_),
    .A(net524),
    .B(net536));
 sg13g2_nand2_1 _19182_ (.Y(_10120_),
    .A(_10118_),
    .B(_10119_));
 sg13g2_nand2_1 _19183_ (.Y(_10121_),
    .A(net524),
    .B(net871));
 sg13g2_o21ai_1 _19184_ (.B1(_10121_),
    .Y(_10122_),
    .A1(net555),
    .A2(net898));
 sg13g2_nor3_1 _19185_ (.A(_10117_),
    .B(_10120_),
    .C(_10122_),
    .Y(_10123_));
 sg13g2_nor3_1 _19186_ (.A(net253),
    .B(net255),
    .C(net260),
    .Y(_10124_));
 sg13g2_a22oi_1 _19187_ (.Y(_10125_),
    .B1(_10124_),
    .B2(_09042_),
    .A2(_10123_),
    .A1(_09077_));
 sg13g2_xor2_1 _19188_ (.B(_09020_),
    .A(net878),
    .X(_10126_));
 sg13g2_xnor2_1 _19189_ (.Y(_10127_),
    .A(net871),
    .B(net1129));
 sg13g2_xnor2_1 _19190_ (.Y(_10128_),
    .A(_10126_),
    .B(_10127_));
 sg13g2_xnor2_1 _19191_ (.Y(_10129_),
    .A(net524),
    .B(_10128_));
 sg13g2_xnor2_1 _19192_ (.Y(_10130_),
    .A(_09661_),
    .B(_10129_));
 sg13g2_buf_1 _19193_ (.A(_00087_),
    .X(_10131_));
 sg13g2_nand2_1 _19194_ (.Y(_10132_),
    .A(net1114),
    .B(_08942_));
 sg13g2_inv_1 _19195_ (.Y(_10133_),
    .A(net1114));
 sg13g2_nand2_1 _19196_ (.Y(_10134_),
    .A(_10133_),
    .B(net558));
 sg13g2_o21ai_1 _19197_ (.B1(_10134_),
    .Y(_10135_),
    .A1(_09746_),
    .A2(_10129_));
 sg13g2_a21oi_1 _19198_ (.A1(_10130_),
    .A2(_10132_),
    .Y(_10136_),
    .B1(_10135_));
 sg13g2_xnor2_1 _19199_ (.Y(_10137_),
    .A(_10125_),
    .B(_10136_));
 sg13g2_nor2_1 _19200_ (.A(_09746_),
    .B(_10129_),
    .Y(_10138_));
 sg13g2_and2_1 _19201_ (.A(_10133_),
    .B(_09769_),
    .X(_10139_));
 sg13g2_inv_1 _19202_ (.Y(_10140_),
    .A(net871));
 sg13g2_xnor2_1 _19203_ (.Y(_10141_),
    .A(_09733_),
    .B(net1129));
 sg13g2_nor2_1 _19204_ (.A(_10140_),
    .B(_10141_),
    .Y(_10142_));
 sg13g2_and3_1 _19205_ (.X(_10143_),
    .A(_10140_),
    .B(_09742_),
    .C(net898));
 sg13g2_o21ai_1 _19206_ (.B1(net275),
    .Y(_10144_),
    .A1(_10142_),
    .A2(_10143_));
 sg13g2_o21ai_1 _19207_ (.B1(_10144_),
    .Y(_10145_),
    .A1(_09077_),
    .A2(_10118_));
 sg13g2_buf_1 _19208_ (.A(net253),
    .X(_10146_));
 sg13g2_nor3_1 _19209_ (.A(net142),
    .B(_09042_),
    .C(_10118_),
    .Y(_10147_));
 sg13g2_a221oi_1 _19210_ (.B2(net142),
    .C1(_10147_),
    .B1(_10145_),
    .A1(_10138_),
    .Y(_10148_),
    .A2(_10139_));
 sg13g2_a21o_1 _19211_ (.A2(_10148_),
    .A1(_10137_),
    .B1(net124),
    .X(_10149_));
 sg13g2_buf_1 _19212_ (.A(net168),
    .X(_10150_));
 sg13g2_xnor2_1 _19213_ (.Y(_10151_),
    .A(_10076_),
    .B(_10130_));
 sg13g2_o21ai_1 _19214_ (.B1(net534),
    .Y(_10152_),
    .A1(net97),
    .A2(_10151_));
 sg13g2_nand3_1 _19215_ (.B(_10149_),
    .C(_10152_),
    .A(net57),
    .Y(_10153_));
 sg13g2_a21oi_1 _19216_ (.A1(_10112_),
    .A2(_10153_),
    .Y(_00386_),
    .B1(net305));
 sg13g2_buf_1 _19217_ (.A(_00149_),
    .X(_10154_));
 sg13g2_nor2b_1 _19218_ (.A(net1113),
    .B_N(_09875_),
    .Y(_10155_));
 sg13g2_buf_1 _19219_ (.A(net531),
    .X(_10156_));
 sg13g2_xnor2_1 _19220_ (.Y(_10157_),
    .A(_09545_),
    .B(net554));
 sg13g2_o21ai_1 _19221_ (.B1(net145),
    .Y(_10158_),
    .A1(_09872_),
    .A2(_09821_));
 sg13g2_a21oi_1 _19222_ (.A1(net252),
    .A2(_10157_),
    .Y(_10159_),
    .B1(_10158_));
 sg13g2_o21ai_1 _19223_ (.B1(net142),
    .Y(_10160_),
    .A1(_10155_),
    .A2(_10159_));
 sg13g2_inv_2 _19224_ (.Y(_10161_),
    .A(net870));
 sg13g2_nand3_1 _19225_ (.B(_09103_),
    .C(_09875_),
    .A(_10161_),
    .Y(_10162_));
 sg13g2_nand3_1 _19226_ (.B(_10160_),
    .C(_10162_),
    .A(net171),
    .Y(_10163_));
 sg13g2_buf_1 _19227_ (.A(_00119_),
    .X(_10164_));
 sg13g2_buf_1 _19228_ (.A(_10164_),
    .X(_10165_));
 sg13g2_inv_1 _19229_ (.Y(_10166_),
    .A(_09788_));
 sg13g2_xnor2_1 _19230_ (.Y(_10167_),
    .A(_10113_),
    .B(_08742_));
 sg13g2_xor2_1 _19231_ (.B(_10167_),
    .A(_09859_),
    .X(_10168_));
 sg13g2_xnor2_1 _19232_ (.Y(_10169_),
    .A(_09034_),
    .B(_10168_));
 sg13g2_nor4_1 _19233_ (.A(net1119),
    .B(net869),
    .C(_10166_),
    .D(_10169_),
    .Y(_10170_));
 sg13g2_nand2_1 _19234_ (.Y(_10171_),
    .A(net869),
    .B(_08985_));
 sg13g2_xnor2_1 _19235_ (.Y(_10172_),
    .A(net537),
    .B(_10169_));
 sg13g2_nand2b_1 _19236_ (.Y(_10173_),
    .B(net898),
    .A_N(_10164_));
 sg13g2_o21ai_1 _19237_ (.B1(_10173_),
    .Y(_10174_),
    .A1(net1119),
    .A2(_10169_));
 sg13g2_a21oi_1 _19238_ (.A1(_10171_),
    .A2(_10172_),
    .Y(_10175_),
    .B1(_10174_));
 sg13g2_o21ai_1 _19239_ (.B1(_09892_),
    .Y(_10176_),
    .A1(net524),
    .A2(_09875_));
 sg13g2_nor2_1 _19240_ (.A(_10115_),
    .B(_09892_),
    .Y(_10177_));
 sg13g2_a21oi_1 _19241_ (.A1(net1113),
    .A2(_10176_),
    .Y(_10178_),
    .B1(_10177_));
 sg13g2_or2_1 _19242_ (.X(_10179_),
    .B(_10178_),
    .A(net145));
 sg13g2_o21ai_1 _19243_ (.B1(_09103_),
    .Y(_10180_),
    .A1(net1113),
    .A2(_09892_));
 sg13g2_nor2_1 _19244_ (.A(_09875_),
    .B(_10180_),
    .Y(_10181_));
 sg13g2_o21ai_1 _19245_ (.B1(_10116_),
    .Y(_10182_),
    .A1(_10155_),
    .A2(_10181_));
 sg13g2_nor2b_1 _19246_ (.A(_10114_),
    .B_N(net1113),
    .Y(_10183_));
 sg13g2_nand2_1 _19247_ (.Y(_10184_),
    .A(net530),
    .B(net564));
 sg13g2_nand2_1 _19248_ (.Y(_10185_),
    .A(_09879_),
    .B(_10184_));
 sg13g2_nor2b_1 _19249_ (.A(net1113),
    .B_N(net530),
    .Y(_10186_));
 sg13g2_a22oi_1 _19250_ (.Y(_10187_),
    .B1(_10186_),
    .B2(net265),
    .A2(_10185_),
    .A1(_10183_));
 sg13g2_and2_1 _19251_ (.A(net870),
    .B(net876),
    .X(_10188_));
 sg13g2_buf_1 _19252_ (.A(_10188_),
    .X(_10189_));
 sg13g2_a21oi_1 _19253_ (.A1(net265),
    .A2(_10189_),
    .Y(_10190_),
    .B1(_10177_));
 sg13g2_mux2_1 _19254_ (.A0(_10187_),
    .A1(_10190_),
    .S(net555),
    .X(_10191_));
 sg13g2_nand3_1 _19255_ (.B(_10182_),
    .C(_10191_),
    .A(_10179_),
    .Y(_10192_));
 sg13g2_xnor2_1 _19256_ (.Y(_10193_),
    .A(_10175_),
    .B(_10192_));
 sg13g2_nor3_1 _19257_ (.A(_10163_),
    .B(_10170_),
    .C(_10193_),
    .Y(_10194_));
 sg13g2_and2_1 _19258_ (.A(net144),
    .B(net57),
    .X(_10195_));
 sg13g2_o21ai_1 _19259_ (.B1(_10195_),
    .Y(_10196_),
    .A1(net75),
    .A2(_10194_));
 sg13g2_xor2_1 _19260_ (.B(_10169_),
    .A(_10079_),
    .X(_10197_));
 sg13g2_nor2_1 _19261_ (.A(net56),
    .B(_10197_),
    .Y(_10198_));
 sg13g2_a22oi_1 _19262_ (.Y(_10199_),
    .B1(_10194_),
    .B2(_10198_),
    .A2(net56),
    .A1(net45));
 sg13g2_buf_1 _19263_ (.A(_06110_),
    .X(_10200_));
 sg13g2_a21oi_1 _19264_ (.A1(_10196_),
    .A2(_10199_),
    .Y(_00387_),
    .B1(_10200_));
 sg13g2_xor2_1 _19265_ (.B(_10167_),
    .A(_10126_),
    .X(_10201_));
 sg13g2_xnor2_1 _19266_ (.Y(_10202_),
    .A(_09880_),
    .B(_10201_));
 sg13g2_xor2_1 _19267_ (.B(_10202_),
    .A(net883),
    .X(_10203_));
 sg13g2_xnor2_1 _19268_ (.Y(_10204_),
    .A(_09866_),
    .B(_10203_));
 sg13g2_nand2_1 _19269_ (.Y(_10205_),
    .A(net544),
    .B(_10204_));
 sg13g2_and2_1 _19270_ (.A(_09871_),
    .B(net878),
    .X(_10206_));
 sg13g2_buf_1 _19271_ (.A(_10206_),
    .X(_10207_));
 sg13g2_nor2b_1 _19272_ (.A(_10154_),
    .B_N(_10207_),
    .Y(_10208_));
 sg13g2_nand2_1 _19273_ (.Y(_10209_),
    .A(net554),
    .B(net279));
 sg13g2_nor3_1 _19274_ (.A(_10154_),
    .B(_09872_),
    .C(net535),
    .Y(_10210_));
 sg13g2_nor3_1 _19275_ (.A(_10209_),
    .B(_10207_),
    .C(_10210_),
    .Y(_10211_));
 sg13g2_o21ai_1 _19276_ (.B1(_10116_),
    .Y(_10212_),
    .A1(_10208_),
    .A2(_10211_));
 sg13g2_nor2_1 _19277_ (.A(_09871_),
    .B(net878),
    .Y(_10213_));
 sg13g2_nand2_1 _19278_ (.Y(_10214_),
    .A(_10161_),
    .B(_10213_));
 sg13g2_a21oi_1 _19279_ (.A1(_09880_),
    .A2(net878),
    .Y(_10215_),
    .B1(_10115_));
 sg13g2_o21ai_1 _19280_ (.B1(net1113),
    .Y(_10216_),
    .A1(_10213_),
    .A2(_10215_));
 sg13g2_a21oi_1 _19281_ (.A1(_10214_),
    .A2(_10216_),
    .Y(_10217_),
    .B1(net145));
 sg13g2_mux2_1 _19282_ (.A0(net878),
    .A1(net564),
    .S(net876),
    .X(_10218_));
 sg13g2_nor2b_1 _19283_ (.A(net1113),
    .B_N(net563),
    .Y(_10219_));
 sg13g2_a22oi_1 _19284_ (.Y(_10220_),
    .B1(_10219_),
    .B2(_10207_),
    .A2(_10218_),
    .A1(_10183_));
 sg13g2_nor2_1 _19285_ (.A(net555),
    .B(_10220_),
    .Y(_10221_));
 sg13g2_nand3_1 _19286_ (.B(net279),
    .C(_10189_),
    .A(net535),
    .Y(_10222_));
 sg13g2_a21oi_1 _19287_ (.A1(_10214_),
    .A2(_10222_),
    .Y(_10223_),
    .B1(net554));
 sg13g2_nor3_1 _19288_ (.A(_10217_),
    .B(_10221_),
    .C(_10223_),
    .Y(_10224_));
 sg13g2_nand2_1 _19289_ (.Y(_10225_),
    .A(_10212_),
    .B(_10224_));
 sg13g2_a221oi_1 _19290_ (.B2(_09900_),
    .C1(_09901_),
    .B1(_10203_),
    .A1(_09535_),
    .Y(_10226_),
    .A2(_10202_));
 sg13g2_xnor2_1 _19291_ (.Y(_10227_),
    .A(_10225_),
    .B(_10226_));
 sg13g2_nand2_1 _19292_ (.Y(_10228_),
    .A(net252),
    .B(_10126_));
 sg13g2_o21ai_1 _19293_ (.B1(_10228_),
    .Y(_10229_),
    .A1(_10156_),
    .A2(_09736_));
 sg13g2_a21oi_1 _19294_ (.A1(net145),
    .A2(_10229_),
    .Y(_10230_),
    .B1(_10208_));
 sg13g2_a21oi_1 _19295_ (.A1(_09103_),
    .A2(_10207_),
    .Y(_10231_),
    .B1(net142));
 sg13g2_a21oi_1 _19296_ (.A1(_10146_),
    .A2(_10230_),
    .Y(_10232_),
    .B1(_10231_));
 sg13g2_xnor2_1 _19297_ (.Y(_10233_),
    .A(net904),
    .B(net883));
 sg13g2_and4_1 _19298_ (.A(_09910_),
    .B(_09535_),
    .C(_10202_),
    .D(_10233_),
    .X(_10234_));
 sg13g2_nor4_1 _19299_ (.A(net107),
    .B(_10227_),
    .C(_10232_),
    .D(_10234_),
    .Y(_10235_));
 sg13g2_a22oi_1 _19300_ (.Y(_10236_),
    .B1(_10205_),
    .B2(_10235_),
    .A2(net75),
    .A1(_09799_));
 sg13g2_buf_2 _19301_ (.A(net1056),
    .X(_10237_));
 sg13g2_o21ai_1 _19302_ (.B1(_10237_),
    .Y(_10238_),
    .A1(net80),
    .A2(net57));
 sg13g2_a21oi_1 _19303_ (.A1(net57),
    .A2(_10236_),
    .Y(_00388_),
    .B1(_10238_));
 sg13g2_nand2_2 _19304_ (.Y(_10239_),
    .A(_05175_),
    .B(_05183_));
 sg13g2_or2_1 _19305_ (.X(_10240_),
    .B(_10239_),
    .A(_09522_));
 sg13g2_buf_2 _19306_ (.A(_10240_),
    .X(_10241_));
 sg13g2_inv_1 _19307_ (.Y(_10242_),
    .A(_10241_));
 sg13g2_buf_1 _19308_ (.A(_10242_),
    .X(_10243_));
 sg13g2_buf_1 _19309_ (.A(_09865_),
    .X(_10244_));
 sg13g2_buf_2 _19310_ (.A(\grid.cell_22_0.sw ),
    .X(_10245_));
 sg13g2_buf_1 _19311_ (.A(_10245_),
    .X(_10246_));
 sg13g2_buf_1 _19312_ (.A(\grid.cell_22_0.se ),
    .X(_10247_));
 sg13g2_buf_1 _19313_ (.A(_10247_),
    .X(_10248_));
 sg13g2_xnor2_1 _19314_ (.Y(_10249_),
    .A(_09528_),
    .B(net866));
 sg13g2_xor2_1 _19315_ (.B(_10249_),
    .A(_09859_),
    .X(_10250_));
 sg13g2_xnor2_1 _19316_ (.Y(_10251_),
    .A(net867),
    .B(_10250_));
 sg13g2_buf_1 _19317_ (.A(\grid.cell_22_0.s ),
    .X(_10252_));
 sg13g2_inv_1 _19318_ (.Y(_10253_),
    .A(net1112));
 sg13g2_xnor2_1 _19319_ (.Y(_10254_),
    .A(_10253_),
    .B(_09927_));
 sg13g2_xnor2_1 _19320_ (.Y(_10255_),
    .A(_10251_),
    .B(_10254_));
 sg13g2_buf_1 _19321_ (.A(net866),
    .X(_10256_));
 sg13g2_buf_1 _19322_ (.A(net521),
    .X(_10257_));
 sg13g2_nor2_1 _19323_ (.A(net867),
    .B(net530),
    .Y(_10258_));
 sg13g2_inv_1 _19324_ (.Y(_10259_),
    .A(_10258_));
 sg13g2_nor2_1 _19325_ (.A(net1121),
    .B(_10259_),
    .Y(_10260_));
 sg13g2_nand2b_1 _19326_ (.Y(_10261_),
    .B(_10245_),
    .A_N(net1118));
 sg13g2_inv_1 _19327_ (.Y(_10262_),
    .A(_10245_));
 sg13g2_buf_1 _19328_ (.A(_10262_),
    .X(_10263_));
 sg13g2_nand2_1 _19329_ (.Y(_10264_),
    .A(net520),
    .B(net264));
 sg13g2_a21oi_1 _19330_ (.A1(_10261_),
    .A2(_10264_),
    .Y(_10265_),
    .B1(net885));
 sg13g2_nand2_1 _19331_ (.Y(_10266_),
    .A(net520),
    .B(net876));
 sg13g2_buf_1 _19332_ (.A(_10246_),
    .X(_10267_));
 sg13g2_nand2b_1 _19333_ (.Y(_10268_),
    .B(net876),
    .A_N(net1121));
 sg13g2_nand2_1 _19334_ (.Y(_10269_),
    .A(net519),
    .B(_10268_));
 sg13g2_a21oi_1 _19335_ (.A1(_10266_),
    .A2(_10269_),
    .Y(_10270_),
    .B1(net259));
 sg13g2_or3_1 _19336_ (.A(_10260_),
    .B(_10265_),
    .C(_10270_),
    .X(_10271_));
 sg13g2_o21ai_1 _19337_ (.B1(_09884_),
    .Y(_10272_),
    .A1(net531),
    .A2(net1121));
 sg13g2_nor2_1 _19338_ (.A(net519),
    .B(_10268_),
    .Y(_10273_));
 sg13g2_a221oi_1 _19339_ (.B2(net519),
    .C1(_10273_),
    .B1(_10272_),
    .A1(_09570_),
    .Y(_10274_),
    .A2(_10259_));
 sg13g2_inv_1 _19340_ (.Y(_10275_),
    .A(_10248_));
 sg13g2_nand2_1 _19341_ (.Y(_10276_),
    .A(net867),
    .B(net876));
 sg13g2_nor3_1 _19342_ (.A(_10275_),
    .B(_09621_),
    .C(_10276_),
    .Y(_10277_));
 sg13g2_nor3_1 _19343_ (.A(net866),
    .B(_10267_),
    .C(_09879_),
    .Y(_10278_));
 sg13g2_o21ai_1 _19344_ (.B1(net541),
    .Y(_10279_),
    .A1(_10277_),
    .A2(_10278_));
 sg13g2_o21ai_1 _19345_ (.B1(_10279_),
    .Y(_10280_),
    .A1(net251),
    .A2(_10274_));
 sg13g2_a21oi_1 _19346_ (.A1(net251),
    .A2(_10271_),
    .Y(_10281_),
    .B1(_10280_));
 sg13g2_inv_1 _19347_ (.Y(_10282_),
    .A(net873));
 sg13g2_buf_2 _19348_ (.A(_00200_),
    .X(_10283_));
 sg13g2_nand2b_1 _19349_ (.Y(_10284_),
    .B(_10283_),
    .A_N(_09579_));
 sg13g2_xnor2_1 _19350_ (.Y(_10285_),
    .A(_09947_),
    .B(_10251_));
 sg13g2_nor2b_1 _19351_ (.A(_10283_),
    .B_N(_09579_),
    .Y(_10286_));
 sg13g2_a221oi_1 _19352_ (.B2(_10285_),
    .C1(_10286_),
    .B1(_10284_),
    .A1(_10282_),
    .Y(_10287_),
    .A2(_10251_));
 sg13g2_xnor2_1 _19353_ (.Y(_10288_),
    .A(_10281_),
    .B(_10287_));
 sg13g2_inv_2 _19354_ (.Y(_10289_),
    .A(_10283_));
 sg13g2_nand4_1 _19355_ (.B(_10282_),
    .C(_09927_),
    .A(_10289_),
    .Y(_10290_),
    .D(_10251_));
 sg13g2_and2_1 _19356_ (.A(_10246_),
    .B(net876),
    .X(_10291_));
 sg13g2_buf_2 _19357_ (.A(_10291_),
    .X(_10292_));
 sg13g2_o21ai_1 _19358_ (.B1(net259),
    .Y(_10293_),
    .A1(net541),
    .A2(_10292_));
 sg13g2_nand3_1 _19359_ (.B(_10261_),
    .C(_10266_),
    .A(net885),
    .Y(_10294_));
 sg13g2_nor2b_1 _19360_ (.A(_10293_),
    .B_N(_10294_),
    .Y(_10295_));
 sg13g2_nor2_1 _19361_ (.A(net1121),
    .B(_10276_),
    .Y(_10296_));
 sg13g2_o21ai_1 _19362_ (.B1(net251),
    .Y(_10297_),
    .A1(_10295_),
    .A2(_10296_));
 sg13g2_buf_1 _19363_ (.A(_10275_),
    .X(_10298_));
 sg13g2_nand4_1 _19364_ (.B(_10298_),
    .C(net259),
    .A(net541),
    .Y(_10299_),
    .D(_10292_));
 sg13g2_nand4_1 _19365_ (.B(_10290_),
    .C(_10297_),
    .A(net127),
    .Y(_10300_),
    .D(_10299_));
 sg13g2_nor2_1 _19366_ (.A(_10288_),
    .B(_10300_),
    .Y(_10301_));
 sg13g2_o21ai_1 _19367_ (.B1(_10301_),
    .Y(_10302_),
    .A1(net868),
    .A2(_10255_));
 sg13g2_a21oi_1 _19368_ (.A1(net868),
    .A2(net69),
    .Y(_10303_),
    .B1(net30));
 sg13g2_a221oi_1 _19369_ (.B2(_10303_),
    .C1(_09818_),
    .B1(_10302_),
    .A1(net50),
    .Y(_00389_),
    .A2(net30));
 sg13g2_buf_1 _19370_ (.A(\grid.cell_22_1.se ),
    .X(_10304_));
 sg13g2_buf_1 _19371_ (.A(_10304_),
    .X(_10305_));
 sg13g2_buf_1 _19372_ (.A(net865),
    .X(_10306_));
 sg13g2_buf_1 _19373_ (.A(net518),
    .X(_10307_));
 sg13g2_nor2_1 _19374_ (.A(_09561_),
    .B(_09587_),
    .Y(_10308_));
 sg13g2_o21ai_1 _19375_ (.B1(_10308_),
    .Y(_10309_),
    .A1(net249),
    .A2(net1121));
 sg13g2_nor2b_1 _19376_ (.A(net1121),
    .B_N(net865),
    .Y(_10310_));
 sg13g2_inv_1 _19377_ (.Y(_10311_),
    .A(net865));
 sg13g2_and2_1 _19378_ (.A(net517),
    .B(_10308_),
    .X(_10312_));
 sg13g2_o21ai_1 _19379_ (.B1(net257),
    .Y(_10313_),
    .A1(_10310_),
    .A2(_10312_));
 sg13g2_o21ai_1 _19380_ (.B1(_10313_),
    .Y(_10314_),
    .A1(net257),
    .A2(_10309_));
 sg13g2_nor2_1 _19381_ (.A(_10305_),
    .B(_09621_),
    .Y(_10315_));
 sg13g2_nor2_1 _19382_ (.A(net875),
    .B(_10310_),
    .Y(_10316_));
 sg13g2_or2_1 _19383_ (.X(_10317_),
    .B(_10316_),
    .A(_10315_));
 sg13g2_o21ai_1 _19384_ (.B1(net528),
    .Y(_10318_),
    .A1(net518),
    .A2(net1121));
 sg13g2_o21ai_1 _19385_ (.B1(_10318_),
    .Y(_10319_),
    .A1(net517),
    .A2(_09621_));
 sg13g2_a22oi_1 _19386_ (.Y(_10320_),
    .B1(_10319_),
    .B2(_10308_),
    .A2(_10317_),
    .A1(net539));
 sg13g2_nor3_1 _19387_ (.A(net866),
    .B(net528),
    .C(net518),
    .Y(_10321_));
 sg13g2_nand4_1 _19388_ (.B(net882),
    .C(net528),
    .A(_10256_),
    .Y(_10322_),
    .D(_10306_));
 sg13g2_nand2b_1 _19389_ (.Y(_10323_),
    .B(_10322_),
    .A_N(_10321_));
 sg13g2_a22oi_1 _19390_ (.Y(_10324_),
    .B1(_10323_),
    .B2(_09561_),
    .A2(_10315_),
    .A1(_09944_));
 sg13g2_o21ai_1 _19391_ (.B1(_10324_),
    .Y(_10325_),
    .A1(_10257_),
    .A2(_10320_));
 sg13g2_a21oi_1 _19392_ (.A1(_10257_),
    .A2(_10314_),
    .Y(_10326_),
    .B1(_10325_));
 sg13g2_xnor2_1 _19393_ (.Y(_10327_),
    .A(net517),
    .B(_09925_));
 sg13g2_xor2_1 _19394_ (.B(_10327_),
    .A(_10249_),
    .X(_10328_));
 sg13g2_xnor2_1 _19395_ (.Y(_10329_),
    .A(_10244_),
    .B(_10328_));
 sg13g2_nand2_1 _19396_ (.Y(_10330_),
    .A(net883),
    .B(_10289_));
 sg13g2_o21ai_1 _19397_ (.B1(_10330_),
    .Y(_10331_),
    .A1(net1117),
    .A2(_10328_));
 sg13g2_a21oi_1 _19398_ (.A1(_10284_),
    .A2(_10329_),
    .Y(_10332_),
    .B1(_10331_));
 sg13g2_xnor2_1 _19399_ (.Y(_10333_),
    .A(_10326_),
    .B(_10332_));
 sg13g2_nand2_1 _19400_ (.Y(_10334_),
    .A(_09943_),
    .B(_10306_));
 sg13g2_xor2_1 _19401_ (.B(net865),
    .A(_09920_),
    .X(_10335_));
 sg13g2_nand2_1 _19402_ (.Y(_10336_),
    .A(net885),
    .B(_10335_));
 sg13g2_o21ai_1 _19403_ (.B1(_10336_),
    .Y(_10337_),
    .A1(net541),
    .A2(_10334_));
 sg13g2_a22oi_1 _19404_ (.Y(_10338_),
    .B1(_10337_),
    .B2(net542),
    .A2(_10310_),
    .A1(net257));
 sg13g2_nand4_1 _19405_ (.B(net250),
    .C(net249),
    .A(net541),
    .Y(_10339_),
    .D(_09939_));
 sg13g2_o21ai_1 _19406_ (.B1(_10339_),
    .Y(_10340_),
    .A1(_10298_),
    .A2(_10338_));
 sg13g2_xor2_1 _19407_ (.B(_09865_),
    .A(net883),
    .X(_10341_));
 sg13g2_nor3_1 _19408_ (.A(_10283_),
    .B(net1117),
    .C(_10341_),
    .Y(_10342_));
 sg13g2_nor2b_1 _19409_ (.A(_10328_),
    .B_N(_10342_),
    .Y(_10343_));
 sg13g2_xnor2_1 _19410_ (.Y(_10344_),
    .A(_09865_),
    .B(net1112));
 sg13g2_xnor2_1 _19411_ (.Y(_10345_),
    .A(net883),
    .B(_10344_));
 sg13g2_xnor2_1 _19412_ (.Y(_10346_),
    .A(_10328_),
    .B(_10345_));
 sg13g2_nor2_1 _19413_ (.A(net529),
    .B(_10346_),
    .Y(_10347_));
 sg13g2_nor4_1 _19414_ (.A(net120),
    .B(_10340_),
    .C(_10343_),
    .D(_10347_),
    .Y(_10348_));
 sg13g2_a221oi_1 _19415_ (.B2(_10348_),
    .C1(net30),
    .B1(_10333_),
    .A1(net529),
    .Y(_10349_),
    .A2(net69));
 sg13g2_o21ai_1 _19416_ (.B1(net356),
    .Y(_10350_),
    .A1(net49),
    .A2(_10241_));
 sg13g2_nor2_1 _19417_ (.A(_10349_),
    .B(_10350_),
    .Y(_00390_));
 sg13g2_nand2_1 _19418_ (.Y(_10351_),
    .A(net714),
    .B(net30));
 sg13g2_buf_1 _19419_ (.A(\grid.cell_22_2.se ),
    .X(_10352_));
 sg13g2_buf_1 _19420_ (.A(_10352_),
    .X(_10353_));
 sg13g2_nand2_1 _19421_ (.Y(_10354_),
    .A(net864),
    .B(net874));
 sg13g2_nor2b_1 _19422_ (.A(net864),
    .B_N(net874),
    .Y(_10355_));
 sg13g2_nor2b_1 _19423_ (.A(net874),
    .B_N(net864),
    .Y(_10356_));
 sg13g2_o21ai_1 _19424_ (.B1(net1122),
    .Y(_10357_),
    .A1(_10355_),
    .A2(_10356_));
 sg13g2_o21ai_1 _19425_ (.B1(_10357_),
    .Y(_10358_),
    .A1(net882),
    .A2(_10354_));
 sg13g2_nand2_1 _19426_ (.Y(_10359_),
    .A(net263),
    .B(_10358_));
 sg13g2_o21ai_1 _19427_ (.B1(_10359_),
    .Y(_10360_),
    .A1(net1120),
    .A2(_10354_));
 sg13g2_nor3_1 _19428_ (.A(net539),
    .B(net249),
    .C(_09981_),
    .Y(_10361_));
 sg13g2_buf_1 _19429_ (.A(net864),
    .X(_10362_));
 sg13g2_buf_1 _19430_ (.A(net516),
    .X(_10363_));
 sg13g2_buf_2 _19431_ (.A(_00197_),
    .X(_10364_));
 sg13g2_buf_1 _19432_ (.A(_10364_),
    .X(_10365_));
 sg13g2_xor2_1 _19433_ (.B(net881),
    .A(_10353_),
    .X(_10366_));
 sg13g2_xnor2_1 _19434_ (.Y(_10367_),
    .A(_10305_),
    .B(_09977_));
 sg13g2_xnor2_1 _19435_ (.Y(_10368_),
    .A(_10366_),
    .B(_10367_));
 sg13g2_xnor2_1 _19436_ (.Y(_10369_),
    .A(net1122),
    .B(_10368_));
 sg13g2_xor2_1 _19437_ (.B(_09870_),
    .A(net541),
    .X(_10370_));
 sg13g2_nor4_1 _19438_ (.A(net863),
    .B(_09991_),
    .C(_10369_),
    .D(_10370_),
    .Y(_10371_));
 sg13g2_a221oi_1 _19439_ (.B2(net248),
    .C1(_10371_),
    .B1(_10361_),
    .A1(net249),
    .Y(_10372_),
    .A2(_10360_));
 sg13g2_inv_1 _19440_ (.Y(_10373_),
    .A(_10354_));
 sg13g2_o21ai_1 _19441_ (.B1(_10357_),
    .Y(_10374_),
    .A1(net540),
    .A2(_10373_));
 sg13g2_nand2_1 _19442_ (.Y(_10375_),
    .A(net882),
    .B(net540));
 sg13g2_nor2_1 _19443_ (.A(net516),
    .B(net527),
    .Y(_10376_));
 sg13g2_a22oi_1 _19444_ (.Y(_10377_),
    .B1(_10375_),
    .B2(_10376_),
    .A2(_10374_),
    .A1(net1120));
 sg13g2_o21ai_1 _19445_ (.B1(net263),
    .Y(_10378_),
    .A1(net539),
    .A2(net517));
 sg13g2_nand3_1 _19446_ (.B(_10378_),
    .C(_10376_),
    .A(net1120),
    .Y(_10379_));
 sg13g2_o21ai_1 _19447_ (.B1(_10379_),
    .Y(_10380_),
    .A1(_10307_),
    .A2(_10377_));
 sg13g2_xnor2_1 _19448_ (.Y(_10381_),
    .A(_09870_),
    .B(_10369_));
 sg13g2_nand2_1 _19449_ (.Y(_10382_),
    .A(_09561_),
    .B(_10365_));
 sg13g2_inv_2 _19450_ (.Y(_10383_),
    .A(_10364_));
 sg13g2_nand2_1 _19451_ (.Y(_10384_),
    .A(net885),
    .B(_10383_));
 sg13g2_o21ai_1 _19452_ (.B1(_10384_),
    .Y(_10385_),
    .A1(net873),
    .A2(_10369_));
 sg13g2_a21oi_1 _19453_ (.A1(_10381_),
    .A2(_10382_),
    .Y(_10386_),
    .B1(_10385_));
 sg13g2_xor2_1 _19454_ (.B(_10386_),
    .A(_10380_),
    .X(_10387_));
 sg13g2_a21oi_1 _19455_ (.A1(_10372_),
    .A2(_10387_),
    .Y(_10388_),
    .B1(net102));
 sg13g2_xnor2_1 _19456_ (.Y(_10389_),
    .A(_10249_),
    .B(_10381_));
 sg13g2_a21oi_1 _19457_ (.A1(net111),
    .A2(_10389_),
    .Y(_10390_),
    .B1(_09976_));
 sg13g2_or4_1 _19458_ (.A(net1057),
    .B(net30),
    .C(_10388_),
    .D(_10390_),
    .X(_10391_));
 sg13g2_o21ai_1 _19459_ (.B1(_10391_),
    .Y(_00391_),
    .A1(net27),
    .A2(_10351_));
 sg13g2_inv_1 _19460_ (.Y(_10392_),
    .A(net864));
 sg13g2_nor2_1 _19461_ (.A(_09706_),
    .B(net515),
    .Y(_10393_));
 sg13g2_xnor2_1 _19462_ (.Y(_10394_),
    .A(net1116),
    .B(net881));
 sg13g2_a21oi_1 _19463_ (.A1(net872),
    .A2(net881),
    .Y(_10395_),
    .B1(net864));
 sg13g2_a21oi_1 _19464_ (.A1(net864),
    .A2(_10394_),
    .Y(_10396_),
    .B1(_10395_));
 sg13g2_a22oi_1 _19465_ (.Y(_10397_),
    .B1(_10396_),
    .B2(net538),
    .A2(_10393_),
    .A1(net872));
 sg13g2_buf_2 _19466_ (.A(\grid.cell_22_3.se ),
    .X(_10398_));
 sg13g2_buf_1 _19467_ (.A(_10398_),
    .X(_10399_));
 sg13g2_buf_1 _19468_ (.A(net862),
    .X(_10400_));
 sg13g2_buf_1 _19469_ (.A(net514),
    .X(_10401_));
 sg13g2_nand2b_1 _19470_ (.Y(_10402_),
    .B(net247),
    .A_N(_10397_));
 sg13g2_nor2_1 _19471_ (.A(net862),
    .B(_10023_),
    .Y(_10403_));
 sg13g2_nand4_1 _19472_ (.B(net538),
    .C(net263),
    .A(net248),
    .Y(_10404_),
    .D(_10403_));
 sg13g2_buf_2 _19473_ (.A(_00194_),
    .X(_10405_));
 sg13g2_xnor2_1 _19474_ (.Y(_10406_),
    .A(net1116),
    .B(_09659_));
 sg13g2_xnor2_1 _19475_ (.Y(_10407_),
    .A(_10398_),
    .B(_10406_));
 sg13g2_xnor2_1 _19476_ (.Y(_10408_),
    .A(_10366_),
    .B(_10407_));
 sg13g2_or4_1 _19477_ (.A(_10405_),
    .B(net1115),
    .C(_09925_),
    .D(_10408_),
    .X(_10409_));
 sg13g2_nand4_1 _19478_ (.B(_10402_),
    .C(_10404_),
    .A(_12956_),
    .Y(_10410_),
    .D(_10409_));
 sg13g2_nor2_1 _19479_ (.A(net862),
    .B(net516),
    .Y(_10411_));
 sg13g2_nor2_1 _19480_ (.A(_09679_),
    .B(net540),
    .Y(_10412_));
 sg13g2_a221oi_1 _19481_ (.B2(_10411_),
    .C1(_10412_),
    .B1(_10030_),
    .A1(_10362_),
    .Y(_10413_),
    .A2(net525));
 sg13g2_o21ai_1 _19482_ (.B1(net514),
    .Y(_10414_),
    .A1(_10362_),
    .A2(net872));
 sg13g2_and2_1 _19483_ (.A(_09706_),
    .B(_10414_),
    .X(_10415_));
 sg13g2_nor3_1 _19484_ (.A(net514),
    .B(net248),
    .C(net525),
    .Y(_10416_));
 sg13g2_a22oi_1 _19485_ (.Y(_10417_),
    .B1(_10416_),
    .B2(_09681_),
    .A2(_10415_),
    .A1(_10413_));
 sg13g2_nand2_1 _19486_ (.Y(_10418_),
    .A(net539),
    .B(_10405_));
 sg13g2_xnor2_1 _19487_ (.Y(_10419_),
    .A(net528),
    .B(_10408_));
 sg13g2_nand2b_1 _19488_ (.Y(_10420_),
    .B(net882),
    .A_N(_10405_));
 sg13g2_o21ai_1 _19489_ (.B1(_10420_),
    .Y(_10421_),
    .A1(net1115),
    .A2(_10408_));
 sg13g2_a21oi_1 _19490_ (.A1(_10418_),
    .A2(_10419_),
    .Y(_10422_),
    .B1(_10421_));
 sg13g2_xnor2_1 _19491_ (.Y(_10423_),
    .A(_10417_),
    .B(_10422_));
 sg13g2_nor2b_1 _19492_ (.A(_10410_),
    .B_N(_10423_),
    .Y(_10424_));
 sg13g2_xor2_1 _19493_ (.B(_10408_),
    .A(_10327_),
    .X(_10425_));
 sg13g2_nor3_1 _19494_ (.A(_05407_),
    .B(_10425_),
    .C(_10410_),
    .Y(_10426_));
 sg13g2_a21o_1 _19495_ (.A2(_10426_),
    .A1(_10423_),
    .B1(net256),
    .X(_10427_));
 sg13g2_o21ai_1 _19496_ (.B1(_10427_),
    .Y(_10428_),
    .A1(_08877_),
    .A2(_10424_));
 sg13g2_nand2b_1 _19497_ (.Y(_10429_),
    .B(net30),
    .A_N(net26));
 sg13g2_o21ai_1 _19498_ (.B1(_10429_),
    .Y(_00392_),
    .A1(_10243_),
    .A2(_10428_));
 sg13g2_buf_1 _19499_ (.A(\grid.cell_22_4.se ),
    .X(_10430_));
 sg13g2_buf_1 _19500_ (.A(_10430_),
    .X(_10431_));
 sg13g2_nor2_1 _19501_ (.A(net861),
    .B(net514),
    .Y(_10432_));
 sg13g2_nor2_1 _19502_ (.A(net526),
    .B(net534),
    .Y(_10433_));
 sg13g2_nand2_1 _19503_ (.Y(_10434_),
    .A(net862),
    .B(_10078_));
 sg13g2_o21ai_1 _19504_ (.B1(_10434_),
    .Y(_10435_),
    .A1(net534),
    .A2(net538));
 sg13g2_a21oi_1 _19505_ (.A1(_10432_),
    .A2(_10433_),
    .Y(_10436_),
    .B1(_10435_));
 sg13g2_o21ai_1 _19506_ (.B1(_10431_),
    .Y(_10437_),
    .A1(net514),
    .A2(_10082_));
 sg13g2_and2_1 _19507_ (.A(_09746_),
    .B(_10437_),
    .X(_10438_));
 sg13g2_buf_1 _19508_ (.A(net861),
    .X(_10439_));
 sg13g2_nor3_1 _19509_ (.A(net513),
    .B(_10400_),
    .C(_10082_),
    .Y(_10440_));
 sg13g2_nand2_1 _19510_ (.Y(_10441_),
    .A(net537),
    .B(net538));
 sg13g2_a22oi_1 _19511_ (.Y(_10442_),
    .B1(_10440_),
    .B2(_10441_),
    .A2(_10438_),
    .A1(_10436_));
 sg13g2_xnor2_1 _19512_ (.Y(_10443_),
    .A(_10430_),
    .B(_10077_));
 sg13g2_xnor2_1 _19513_ (.Y(_10444_),
    .A(_09708_),
    .B(_10443_));
 sg13g2_xnor2_1 _19514_ (.Y(_10445_),
    .A(_10399_),
    .B(_10444_));
 sg13g2_xnor2_1 _19515_ (.Y(_10446_),
    .A(_10027_),
    .B(_10445_));
 sg13g2_buf_1 _19516_ (.A(_00054_),
    .X(_10447_));
 sg13g2_nand2b_1 _19517_ (.Y(_10448_),
    .B(net1111),
    .A_N(net263));
 sg13g2_nor2b_1 _19518_ (.A(net1111),
    .B_N(net263),
    .Y(_10449_));
 sg13g2_a221oi_1 _19519_ (.B2(_10448_),
    .C1(_10449_),
    .B1(_10446_),
    .A1(_10106_),
    .Y(_10450_),
    .A2(_10445_));
 sg13g2_xnor2_1 _19520_ (.Y(_10451_),
    .A(_10442_),
    .B(_10450_));
 sg13g2_and2_1 _19521_ (.A(_10106_),
    .B(_10445_),
    .X(_10452_));
 sg13g2_nor2_1 _19522_ (.A(net1111),
    .B(_09978_),
    .Y(_10453_));
 sg13g2_inv_1 _19523_ (.Y(_10454_),
    .A(_10399_));
 sg13g2_xnor2_1 _19524_ (.Y(_10455_),
    .A(_10078_),
    .B(net880));
 sg13g2_nor2_1 _19525_ (.A(_10454_),
    .B(_10455_),
    .Y(_10456_));
 sg13g2_nor3_1 _19526_ (.A(_10400_),
    .B(_10140_),
    .C(_09679_),
    .Y(_10457_));
 sg13g2_o21ai_1 _19527_ (.B1(net261),
    .Y(_10458_),
    .A1(_10456_),
    .A2(_10457_));
 sg13g2_o21ai_1 _19528_ (.B1(_10458_),
    .Y(_10459_),
    .A1(_09746_),
    .A2(_10434_));
 sg13g2_buf_1 _19529_ (.A(net513),
    .X(_10460_));
 sg13g2_nor3_1 _19530_ (.A(net246),
    .B(_10441_),
    .C(_10434_),
    .Y(_10461_));
 sg13g2_a221oi_1 _19531_ (.B2(net246),
    .C1(_10461_),
    .B1(_10459_),
    .A1(_10452_),
    .Y(_10462_),
    .A2(_10453_));
 sg13g2_a21oi_1 _19532_ (.A1(_10451_),
    .A2(_10462_),
    .Y(_10463_),
    .B1(net102));
 sg13g2_xor2_1 _19533_ (.B(_10446_),
    .A(_10366_),
    .X(_10464_));
 sg13g2_a21oi_1 _19534_ (.A1(net111),
    .A2(_10464_),
    .Y(_10465_),
    .B1(_10097_));
 sg13g2_or4_1 _19535_ (.A(net1057),
    .B(_10243_),
    .C(_10463_),
    .D(_10465_),
    .X(_10466_));
 sg13g2_o21ai_1 _19536_ (.B1(_10466_),
    .Y(_00393_),
    .A1(net34),
    .A2(_10351_));
 sg13g2_buf_2 _19537_ (.A(_00086_),
    .X(_10467_));
 sg13g2_xor2_1 _19538_ (.B(_09731_),
    .A(_10113_),
    .X(_10468_));
 sg13g2_buf_2 _19539_ (.A(\grid.cell_22_5.se ),
    .X(_10469_));
 sg13g2_xnor2_1 _19540_ (.Y(_10470_),
    .A(_10469_),
    .B(_10430_));
 sg13g2_xor2_1 _19541_ (.B(_10470_),
    .A(_10468_),
    .X(_10471_));
 sg13g2_xnor2_1 _19542_ (.Y(_10472_),
    .A(_09697_),
    .B(_10471_));
 sg13g2_buf_1 _19543_ (.A(_10472_),
    .X(_10473_));
 sg13g2_a21o_1 _19544_ (.A2(_10473_),
    .A1(_10023_),
    .B1(net262),
    .X(_10474_));
 sg13g2_o21ai_1 _19545_ (.B1(_10473_),
    .Y(_10475_),
    .A1(net1114),
    .A2(net262));
 sg13g2_a221oi_1 _19546_ (.B2(net254),
    .C1(_10030_),
    .B1(_10475_),
    .A1(net1114),
    .Y(_10476_),
    .A2(_10474_));
 sg13g2_xnor2_1 _19547_ (.Y(_10477_),
    .A(_10023_),
    .B(_10473_));
 sg13g2_and2_1 _19548_ (.A(_10133_),
    .B(_10473_),
    .X(_10478_));
 sg13g2_a22oi_1 _19549_ (.Y(_10479_),
    .B1(_10478_),
    .B2(_10467_),
    .A2(_10477_),
    .A1(net262));
 sg13g2_o21ai_1 _19550_ (.B1(_10479_),
    .Y(_10480_),
    .A1(_10467_),
    .A2(_10476_));
 sg13g2_inv_1 _19551_ (.Y(_10481_),
    .A(_10469_));
 sg13g2_buf_1 _19552_ (.A(_10481_),
    .X(_10482_));
 sg13g2_nor2_2 _19553_ (.A(net861),
    .B(net253),
    .Y(_10483_));
 sg13g2_nand2_1 _19554_ (.Y(_10484_),
    .A(net512),
    .B(_10483_));
 sg13g2_nand3_1 _19555_ (.B(net144),
    .C(_10483_),
    .A(net512),
    .Y(_10485_));
 sg13g2_buf_1 _19556_ (.A(_10469_),
    .X(_10486_));
 sg13g2_buf_1 _19557_ (.A(net860),
    .X(_10487_));
 sg13g2_o21ai_1 _19558_ (.B1(_10146_),
    .Y(_10488_),
    .A1(net511),
    .A2(net246));
 sg13g2_a22oi_1 _19559_ (.Y(_10489_),
    .B1(net144),
    .B2(net534),
    .A2(net246),
    .A1(net511));
 sg13g2_nand4_1 _19560_ (.B(_10485_),
    .C(_10488_),
    .A(net1119),
    .Y(_10490_),
    .D(_10489_));
 sg13g2_o21ai_1 _19561_ (.B1(_10490_),
    .Y(_10491_),
    .A1(_09740_),
    .A2(_10484_));
 sg13g2_nand2_1 _19562_ (.Y(_10492_),
    .A(net534),
    .B(_10483_));
 sg13g2_nand2_1 _19563_ (.Y(_10493_),
    .A(net513),
    .B(_09742_));
 sg13g2_o21ai_1 _19564_ (.B1(_10493_),
    .Y(_10494_),
    .A1(_10439_),
    .A2(_10161_));
 sg13g2_nand3_1 _19565_ (.B(net261),
    .C(_10494_),
    .A(net1119),
    .Y(_10495_));
 sg13g2_buf_1 _19566_ (.A(net511),
    .X(_10496_));
 sg13g2_a21oi_1 _19567_ (.A1(_10492_),
    .A2(_10495_),
    .Y(_10497_),
    .B1(net245));
 sg13g2_nand3_1 _19568_ (.B(net246),
    .C(net253),
    .A(net1119),
    .Y(_10498_));
 sg13g2_a21oi_1 _19569_ (.A1(_10439_),
    .A2(net253),
    .Y(_10499_),
    .B1(_09740_));
 sg13g2_a21oi_1 _19570_ (.A1(_09812_),
    .A2(_10483_),
    .Y(_10500_),
    .B1(_10499_));
 sg13g2_nand3_1 _19571_ (.B(_10498_),
    .C(_10500_),
    .A(_10487_),
    .Y(_10501_));
 sg13g2_buf_1 _19572_ (.A(net860),
    .X(_10502_));
 sg13g2_mux2_1 _19573_ (.A0(_09812_),
    .A1(net510),
    .S(net534),
    .X(_10503_));
 sg13g2_nand4_1 _19574_ (.B(net142),
    .C(net144),
    .A(_10460_),
    .Y(_10504_),
    .D(_10503_));
 sg13g2_inv_1 _19575_ (.Y(_10505_),
    .A(_10467_));
 sg13g2_nand2_1 _19576_ (.Y(_10506_),
    .A(_10505_),
    .B(net262));
 sg13g2_nand3_1 _19577_ (.B(_10504_),
    .C(_10506_),
    .A(_10501_),
    .Y(_10507_));
 sg13g2_a21oi_1 _19578_ (.A1(_10460_),
    .A2(net253),
    .Y(_10508_),
    .B1(net510));
 sg13g2_o21ai_1 _19579_ (.B1(net1119),
    .Y(_10509_),
    .A1(_10483_),
    .A2(_10508_));
 sg13g2_a21oi_1 _19580_ (.A1(_10484_),
    .A2(_10509_),
    .Y(_10510_),
    .B1(net144));
 sg13g2_nor4_1 _19581_ (.A(_10478_),
    .B(_10497_),
    .C(_10507_),
    .D(_10510_),
    .Y(_10511_));
 sg13g2_o21ai_1 _19582_ (.B1(_10477_),
    .Y(_10512_),
    .A1(_10505_),
    .A2(net262));
 sg13g2_a221oi_1 _19583_ (.B2(_10512_),
    .C1(net73),
    .B1(_10511_),
    .A1(_10480_),
    .Y(_10513_),
    .A2(_10491_));
 sg13g2_buf_1 _19584_ (.A(_10140_),
    .X(_10514_));
 sg13g2_xor2_1 _19585_ (.B(_10473_),
    .A(_10407_),
    .X(_10515_));
 sg13g2_nand2_1 _19586_ (.Y(_10516_),
    .A(net126),
    .B(_10515_));
 sg13g2_nand3_1 _19587_ (.B(_10241_),
    .C(_10516_),
    .A(net244),
    .Y(_10517_));
 sg13g2_nand2_1 _19588_ (.Y(_10518_),
    .A(_05002_),
    .B(_10242_));
 sg13g2_nand3_1 _19589_ (.B(_10517_),
    .C(_10518_),
    .A(net637),
    .Y(_10519_));
 sg13g2_a21oi_1 _19590_ (.A1(_10241_),
    .A2(_10513_),
    .Y(_00394_),
    .B1(_10519_));
 sg13g2_buf_1 _19591_ (.A(_00118_),
    .X(_10520_));
 sg13g2_xnor2_1 _19592_ (.Y(_10521_),
    .A(_10469_),
    .B(_10245_));
 sg13g2_xor2_1 _19593_ (.B(_10521_),
    .A(_09859_),
    .X(_10522_));
 sg13g2_xnor2_1 _19594_ (.Y(_10523_),
    .A(net536),
    .B(_10522_));
 sg13g2_buf_1 _19595_ (.A(_10523_),
    .X(_10524_));
 sg13g2_a21o_1 _19596_ (.A2(_10524_),
    .A1(_10514_),
    .B1(net261),
    .X(_10525_));
 sg13g2_o21ai_1 _19597_ (.B1(_10524_),
    .Y(_10526_),
    .A1(net869),
    .A2(net261));
 sg13g2_a221oi_1 _19598_ (.B2(_10083_),
    .C1(_10433_),
    .B1(_10526_),
    .A1(_10165_),
    .Y(_10527_),
    .A2(_10525_));
 sg13g2_xnor2_1 _19599_ (.Y(_10528_),
    .A(_10514_),
    .B(_10524_));
 sg13g2_nor2b_1 _19600_ (.A(_10165_),
    .B_N(_10524_),
    .Y(_10529_));
 sg13g2_a22oi_1 _19601_ (.Y(_10530_),
    .B1(_10529_),
    .B2(net1110),
    .A2(_10528_),
    .A1(net261));
 sg13g2_o21ai_1 _19602_ (.B1(_10530_),
    .Y(_10531_),
    .A1(net1110),
    .A2(_10527_));
 sg13g2_nand2_1 _19603_ (.Y(_10532_),
    .A(net512),
    .B(_10258_));
 sg13g2_buf_1 _19604_ (.A(_00148_),
    .X(_10533_));
 sg13g2_buf_1 _19605_ (.A(_10267_),
    .X(_10534_));
 sg13g2_nor3_1 _19606_ (.A(_10487_),
    .B(_10534_),
    .C(_09879_),
    .Y(_10535_));
 sg13g2_o21ai_1 _19607_ (.B1(_10276_),
    .Y(_10536_),
    .A1(net260),
    .A2(net544));
 sg13g2_nor2_1 _19608_ (.A(_10535_),
    .B(_10536_),
    .Y(_10537_));
 sg13g2_o21ai_1 _19609_ (.B1(net245),
    .Y(_10538_),
    .A1(_10534_),
    .A2(net252));
 sg13g2_nand3_1 _19610_ (.B(_10537_),
    .C(_10538_),
    .A(net1109),
    .Y(_10539_));
 sg13g2_o21ai_1 _19611_ (.B1(_10539_),
    .Y(_10540_),
    .A1(_09805_),
    .A2(_10532_));
 sg13g2_nand2_1 _19612_ (.Y(_10541_),
    .A(_10531_),
    .B(_10540_));
 sg13g2_nand2_1 _19613_ (.Y(_10542_),
    .A(_10263_),
    .B(_10213_));
 sg13g2_o21ai_1 _19614_ (.B1(_10266_),
    .Y(_10543_),
    .A1(_10263_),
    .A2(net544));
 sg13g2_nand3_1 _19615_ (.B(net260),
    .C(_10543_),
    .A(net1109),
    .Y(_10544_));
 sg13g2_a21oi_1 _19616_ (.A1(_10542_),
    .A2(_10544_),
    .Y(_10545_),
    .B1(net245));
 sg13g2_nor2_1 _19617_ (.A(net510),
    .B(_10292_),
    .Y(_10546_));
 sg13g2_o21ai_1 _19618_ (.B1(_10533_),
    .Y(_10547_),
    .A1(_10258_),
    .A2(_10546_));
 sg13g2_a21oi_1 _19619_ (.A1(_10532_),
    .A2(_10547_),
    .Y(_10548_),
    .B1(net259));
 sg13g2_inv_1 _19620_ (.Y(_10549_),
    .A(_00148_));
 sg13g2_mux2_1 _19621_ (.A0(_10502_),
    .A1(_10549_),
    .S(net260),
    .X(_10550_));
 sg13g2_nand3_1 _19622_ (.B(_10292_),
    .C(_10550_),
    .A(net259),
    .Y(_10551_));
 sg13g2_o21ai_1 _19623_ (.B1(_10551_),
    .Y(_10552_),
    .A1(net1110),
    .A2(net534));
 sg13g2_nand2_1 _19624_ (.Y(_10553_),
    .A(net1109),
    .B(_10292_));
 sg13g2_o21ai_1 _19625_ (.B1(_10553_),
    .Y(_10554_),
    .A1(net1109),
    .A2(_10259_));
 sg13g2_o21ai_1 _19626_ (.B1(net245),
    .Y(_10555_),
    .A1(_09805_),
    .A2(_10292_));
 sg13g2_nor2_1 _19627_ (.A(_10554_),
    .B(_10555_),
    .Y(_10556_));
 sg13g2_nor4_1 _19628_ (.A(_10545_),
    .B(_10548_),
    .C(_10552_),
    .D(_10556_),
    .Y(_10557_));
 sg13g2_nand2_1 _19629_ (.Y(_10558_),
    .A(net1110),
    .B(_09759_));
 sg13g2_a21oi_1 _19630_ (.A1(_10528_),
    .A2(_10558_),
    .Y(_10559_),
    .B1(_10529_));
 sg13g2_nand2_1 _19631_ (.Y(_10560_),
    .A(net84),
    .B(_10241_));
 sg13g2_a21oi_1 _19632_ (.A1(_10557_),
    .A2(_10559_),
    .Y(_10561_),
    .B1(_10560_));
 sg13g2_nand2_1 _19633_ (.Y(_10562_),
    .A(net45),
    .B(net30));
 sg13g2_xnor2_1 _19634_ (.Y(_10563_),
    .A(net261),
    .B(_10443_));
 sg13g2_xnor2_1 _19635_ (.Y(_10564_),
    .A(_10524_),
    .B(_10563_));
 sg13g2_nor2_1 _19636_ (.A(net107),
    .B(_10564_),
    .Y(_10565_));
 sg13g2_o21ai_1 _19637_ (.B1(_10241_),
    .Y(_10566_),
    .A1(net142),
    .A2(_10565_));
 sg13g2_a221oi_1 _19638_ (.B2(_10566_),
    .C1(net533),
    .B1(_10562_),
    .A1(_10541_),
    .Y(_00395_),
    .A2(_10561_));
 sg13g2_nand2_1 _19639_ (.Y(_10567_),
    .A(net519),
    .B(_10468_));
 sg13g2_o21ai_1 _19640_ (.B1(_10567_),
    .Y(_10568_),
    .A1(net243),
    .A2(_10119_));
 sg13g2_nand2_1 _19641_ (.Y(_10569_),
    .A(net867),
    .B(net870));
 sg13g2_nor2_1 _19642_ (.A(net1109),
    .B(_10569_),
    .Y(_10570_));
 sg13g2_a21oi_1 _19643_ (.A1(net259),
    .A2(_10568_),
    .Y(_10571_),
    .B1(_10570_));
 sg13g2_buf_1 _19644_ (.A(_10245_),
    .X(_10572_));
 sg13g2_and2_1 _19645_ (.A(net859),
    .B(net870),
    .X(_10573_));
 sg13g2_a21oi_1 _19646_ (.A1(_09805_),
    .A2(_10573_),
    .Y(_10574_),
    .B1(net511));
 sg13g2_a21oi_1 _19647_ (.A1(net245),
    .A2(_10571_),
    .Y(_10575_),
    .B1(_10574_));
 sg13g2_xor2_1 _19648_ (.B(_10521_),
    .A(_10468_),
    .X(_10576_));
 sg13g2_xnor2_1 _19649_ (.Y(_10577_),
    .A(net884),
    .B(_10576_));
 sg13g2_a21oi_1 _19650_ (.A1(_10342_),
    .A2(_10577_),
    .Y(_10578_),
    .B1(net163));
 sg13g2_nand3_1 _19651_ (.B(net870),
    .C(net884),
    .A(net859),
    .Y(_10579_));
 sg13g2_mux2_1 _19652_ (.A0(net870),
    .A1(net884),
    .S(net859),
    .X(_10580_));
 sg13g2_nand3_1 _19653_ (.B(net512),
    .C(_10580_),
    .A(net1109),
    .Y(_10581_));
 sg13g2_o21ai_1 _19654_ (.B1(_10581_),
    .Y(_10582_),
    .A1(net1109),
    .A2(_10579_));
 sg13g2_nor2_1 _19655_ (.A(_10572_),
    .B(net870),
    .Y(_10583_));
 sg13g2_nand2_1 _19656_ (.Y(_10584_),
    .A(net512),
    .B(_10583_));
 sg13g2_or2_1 _19657_ (.X(_10585_),
    .B(_10579_),
    .A(_10482_));
 sg13g2_a21oi_1 _19658_ (.A1(_10584_),
    .A2(_10585_),
    .Y(_10586_),
    .B1(net535));
 sg13g2_a21oi_1 _19659_ (.A1(net535),
    .A2(_10582_),
    .Y(_10587_),
    .B1(_10586_));
 sg13g2_nand2_1 _19660_ (.Y(_10588_),
    .A(_09805_),
    .B(_10569_));
 sg13g2_a21oi_1 _19661_ (.A1(_10549_),
    .A2(_10583_),
    .Y(_10589_),
    .B1(_10588_));
 sg13g2_o21ai_1 _19662_ (.B1(net510),
    .Y(_10590_),
    .A1(_10570_),
    .A2(_10589_));
 sg13g2_nor2_1 _19663_ (.A(net860),
    .B(_10573_),
    .Y(_10591_));
 sg13g2_o21ai_1 _19664_ (.B1(net1109),
    .Y(_10592_),
    .A1(_10583_),
    .A2(_10591_));
 sg13g2_a21o_1 _19665_ (.A2(_10592_),
    .A1(_10584_),
    .B1(net259),
    .X(_10593_));
 sg13g2_nand3_1 _19666_ (.B(_10590_),
    .C(_10593_),
    .A(_10587_),
    .Y(_10594_));
 sg13g2_inv_1 _19667_ (.Y(_10595_),
    .A(_09865_));
 sg13g2_xnor2_1 _19668_ (.Y(_10596_),
    .A(_10595_),
    .B(_10577_));
 sg13g2_a221oi_1 _19669_ (.B2(_10284_),
    .C1(_10286_),
    .B1(_10596_),
    .A1(_09910_),
    .Y(_10597_),
    .A2(_10577_));
 sg13g2_xor2_1 _19670_ (.B(_10597_),
    .A(_10594_),
    .X(_10598_));
 sg13g2_nand3b_1 _19671_ (.B(_10578_),
    .C(_10598_),
    .Y(_10599_),
    .A_N(_10575_));
 sg13g2_xnor2_1 _19672_ (.Y(_10600_),
    .A(_10345_),
    .B(_10577_));
 sg13g2_nor2_1 _19673_ (.A(_10156_),
    .B(_10242_),
    .Y(_10601_));
 sg13g2_o21ai_1 _19674_ (.B1(_10601_),
    .Y(_10602_),
    .A1(_10599_),
    .A2(_10600_));
 sg13g2_nand2_1 _19675_ (.Y(_10603_),
    .A(net121),
    .B(net30));
 sg13g2_nand3_1 _19676_ (.B(_10241_),
    .C(_10599_),
    .A(net82),
    .Y(_10604_));
 sg13g2_and4_1 _19677_ (.A(net312),
    .B(_10602_),
    .C(_10603_),
    .D(_10604_),
    .X(_00396_));
 sg13g2_nor2_1 _19678_ (.A(_08817_),
    .B(_09522_),
    .Y(_10605_));
 sg13g2_buf_2 _19679_ (.A(_10605_),
    .X(_10606_));
 sg13g2_buf_1 _19680_ (.A(\grid.cell_23_0.se ),
    .X(_10607_));
 sg13g2_xnor2_1 _19681_ (.Y(_10608_),
    .A(_09860_),
    .B(_10607_));
 sg13g2_buf_2 _19682_ (.A(\grid.cell_23_0.sw ),
    .X(_10609_));
 sg13g2_xnor2_1 _19683_ (.Y(_10610_),
    .A(_10609_),
    .B(_10245_));
 sg13g2_xnor2_1 _19684_ (.Y(_10611_),
    .A(_10608_),
    .B(_10610_));
 sg13g2_xor2_1 _19685_ (.B(_10611_),
    .A(net531),
    .X(_10612_));
 sg13g2_buf_2 _19686_ (.A(_10612_),
    .X(_10613_));
 sg13g2_inv_1 _19687_ (.Y(_10614_),
    .A(_10607_));
 sg13g2_buf_1 _19688_ (.A(_10614_),
    .X(_10615_));
 sg13g2_inv_2 _19689_ (.Y(_10616_),
    .A(_10609_));
 sg13g2_nand2_1 _19690_ (.Y(_10617_),
    .A(_10616_),
    .B(_10262_));
 sg13g2_nor2_1 _19691_ (.A(net873),
    .B(_10617_),
    .Y(_10618_));
 sg13g2_buf_1 _19692_ (.A(_10609_),
    .X(_10619_));
 sg13g2_nand2b_1 _19693_ (.Y(_10620_),
    .B(net858),
    .A_N(net859));
 sg13g2_nand2_1 _19694_ (.Y(_10621_),
    .A(_10616_),
    .B(net1118));
 sg13g2_a21oi_1 _19695_ (.A1(_10620_),
    .A2(_10621_),
    .Y(_10622_),
    .B1(net877));
 sg13g2_nand2_1 _19696_ (.Y(_10623_),
    .A(_10616_),
    .B(net859));
 sg13g2_nand2b_1 _19697_ (.Y(_10624_),
    .B(_10245_),
    .A_N(_09990_));
 sg13g2_nand2_1 _19698_ (.Y(_10625_),
    .A(net858),
    .B(_10624_));
 sg13g2_a21oi_1 _19699_ (.A1(_10623_),
    .A2(_10625_),
    .Y(_10626_),
    .B1(net530));
 sg13g2_nor4_1 _19700_ (.A(net509),
    .B(_10618_),
    .C(_10622_),
    .D(_10626_),
    .Y(_10627_));
 sg13g2_o21ai_1 _19701_ (.B1(_10261_),
    .Y(_10628_),
    .A1(net859),
    .A2(_09990_));
 sg13g2_nor2_1 _19702_ (.A(net858),
    .B(_10624_),
    .Y(_10629_));
 sg13g2_a221oi_1 _19703_ (.B2(_10619_),
    .C1(_10629_),
    .B1(_10628_),
    .A1(_09907_),
    .Y(_10630_),
    .A2(_10617_));
 sg13g2_and2_1 _19704_ (.A(net509),
    .B(_10630_),
    .X(_10631_));
 sg13g2_nand2_1 _19705_ (.Y(_10632_),
    .A(_10619_),
    .B(net859));
 sg13g2_nor3_1 _19706_ (.A(_10615_),
    .B(_10282_),
    .C(_10632_),
    .Y(_10633_));
 sg13g2_buf_1 _19707_ (.A(_10607_),
    .X(_10634_));
 sg13g2_buf_1 _19708_ (.A(net858),
    .X(_10635_));
 sg13g2_nor3_1 _19709_ (.A(net857),
    .B(net508),
    .C(_10266_),
    .Y(_10636_));
 sg13g2_o21ai_1 _19710_ (.B1(net877),
    .Y(_10637_),
    .A1(_10633_),
    .A2(_10636_));
 sg13g2_o21ai_1 _19711_ (.B1(_10637_),
    .Y(_10638_),
    .A1(_10627_),
    .A2(_10631_));
 sg13g2_buf_1 _19712_ (.A(_10638_),
    .X(_10639_));
 sg13g2_nand2_1 _19713_ (.Y(_10640_),
    .A(net251),
    .B(net863));
 sg13g2_buf_1 _19714_ (.A(_00198_),
    .X(_10641_));
 sg13g2_inv_1 _19715_ (.Y(_10642_),
    .A(net1108));
 sg13g2_nand3_1 _19716_ (.B(_10383_),
    .C(_10642_),
    .A(net250),
    .Y(_10643_));
 sg13g2_o21ai_1 _19717_ (.B1(_10643_),
    .Y(_10644_),
    .A1(_10639_),
    .A2(_10640_));
 sg13g2_nor2_1 _19718_ (.A(_09865_),
    .B(net856),
    .Y(_10645_));
 sg13g2_o21ai_1 _19719_ (.B1(_10365_),
    .Y(_10646_),
    .A1(net251),
    .A2(_10645_));
 sg13g2_nand2_1 _19720_ (.Y(_10647_),
    .A(net863),
    .B(net1108));
 sg13g2_nor3_1 _19721_ (.A(net250),
    .B(_10639_),
    .C(_10647_),
    .Y(_10648_));
 sg13g2_a221oi_1 _19722_ (.B2(_10639_),
    .C1(_10648_),
    .B1(_10646_),
    .A1(_10595_),
    .Y(_10649_),
    .A2(_10644_));
 sg13g2_buf_1 _19723_ (.A(net1112),
    .X(_10650_));
 sg13g2_buf_1 _19724_ (.A(\grid.cell_23_0.s ),
    .X(_10651_));
 sg13g2_xnor2_1 _19725_ (.Y(_10652_),
    .A(net1107),
    .B(net866));
 sg13g2_xnor2_1 _19726_ (.Y(_10653_),
    .A(net868),
    .B(_10652_));
 sg13g2_xnor2_1 _19727_ (.Y(_10654_),
    .A(_10613_),
    .B(_10653_));
 sg13g2_nor2_1 _19728_ (.A(net855),
    .B(_10654_),
    .Y(_10655_));
 sg13g2_buf_1 _19729_ (.A(net857),
    .X(_10656_));
 sg13g2_buf_1 _19730_ (.A(net507),
    .X(_10657_));
 sg13g2_buf_1 _19731_ (.A(net508),
    .X(_10658_));
 sg13g2_nand3_1 _19732_ (.B(net241),
    .C(_10292_),
    .A(net529),
    .Y(_10659_));
 sg13g2_o21ai_1 _19733_ (.B1(net167),
    .Y(_10660_),
    .A1(net242),
    .A2(_10659_));
 sg13g2_nor2_1 _19734_ (.A(_10275_),
    .B(net1108),
    .Y(_10661_));
 sg13g2_nand3_1 _19735_ (.B(_10383_),
    .C(_10661_),
    .A(net868),
    .Y(_10662_));
 sg13g2_nand2b_1 _19736_ (.Y(_10663_),
    .B(net877),
    .A_N(_10610_));
 sg13g2_o21ai_1 _19737_ (.B1(_10663_),
    .Y(_10664_),
    .A1(net532),
    .A2(_10632_));
 sg13g2_buf_1 _19738_ (.A(_10616_),
    .X(_10665_));
 sg13g2_nor2_1 _19739_ (.A(net506),
    .B(_10624_),
    .Y(_10666_));
 sg13g2_a21oi_1 _19740_ (.A1(net252),
    .A2(_10664_),
    .Y(_10667_),
    .B1(_10666_));
 sg13g2_nand2b_1 _19741_ (.Y(_10668_),
    .B(_10657_),
    .A_N(_10667_));
 sg13g2_o21ai_1 _19742_ (.B1(_10668_),
    .Y(_10669_),
    .A1(_10613_),
    .A2(_10662_));
 sg13g2_nand2_1 _19743_ (.Y(_10670_),
    .A(net250),
    .B(net1108));
 sg13g2_o21ai_1 _19744_ (.B1(_10670_),
    .Y(_10671_),
    .A1(_09865_),
    .A2(_10661_));
 sg13g2_nand2_1 _19745_ (.Y(_10672_),
    .A(_10613_),
    .B(_10671_));
 sg13g2_o21ai_1 _19746_ (.B1(_10672_),
    .Y(_10673_),
    .A1(net868),
    .A2(_10647_));
 sg13g2_a21oi_1 _19747_ (.A1(_10256_),
    .A2(_10613_),
    .Y(_10674_),
    .B1(net856));
 sg13g2_a21oi_1 _19748_ (.A1(_10613_),
    .A2(_10661_),
    .Y(_10675_),
    .B1(net868));
 sg13g2_nor2_1 _19749_ (.A(_10674_),
    .B(_10675_),
    .Y(_10676_));
 sg13g2_mux2_1 _19750_ (.A0(_10673_),
    .A1(_10676_),
    .S(_10639_),
    .X(_10677_));
 sg13g2_nor4_1 _19751_ (.A(_10655_),
    .B(_10660_),
    .C(_10669_),
    .D(_10677_),
    .Y(_10678_));
 sg13g2_o21ai_1 _19752_ (.B1(_10678_),
    .Y(_10679_),
    .A1(_10613_),
    .A2(_10649_));
 sg13g2_a21oi_1 _19753_ (.A1(_10650_),
    .A2(net69),
    .Y(_10680_),
    .B1(_10606_));
 sg13g2_a221oi_1 _19754_ (.B2(_10680_),
    .C1(net533),
    .B1(_10679_),
    .A1(net50),
    .Y(_00397_),
    .A2(_10606_));
 sg13g2_nand2_1 _19755_ (.Y(_10681_),
    .A(net42),
    .B(_10606_));
 sg13g2_or2_1 _19756_ (.X(_10682_),
    .B(_09522_),
    .A(_08817_));
 sg13g2_buf_1 _19757_ (.A(_10682_),
    .X(_10683_));
 sg13g2_buf_1 _19758_ (.A(_10683_),
    .X(_10684_));
 sg13g2_buf_2 _19759_ (.A(\grid.cell_23_1.se ),
    .X(_10685_));
 sg13g2_buf_1 _19760_ (.A(_10685_),
    .X(_10686_));
 sg13g2_nand2_1 _19761_ (.Y(_10687_),
    .A(net518),
    .B(net854));
 sg13g2_xor2_1 _19762_ (.B(_10685_),
    .A(_10304_),
    .X(_10688_));
 sg13g2_and2_1 _19763_ (.A(net877),
    .B(_10688_),
    .X(_10689_));
 sg13g2_nor2_1 _19764_ (.A(net532),
    .B(_10687_),
    .Y(_10690_));
 sg13g2_o21ai_1 _19765_ (.B1(net257),
    .Y(_10691_),
    .A1(_10689_),
    .A2(_10690_));
 sg13g2_o21ai_1 _19766_ (.B1(_10691_),
    .Y(_10692_),
    .A1(net873),
    .A2(_10687_));
 sg13g2_nand2_1 _19767_ (.Y(_10693_),
    .A(net877),
    .B(net528));
 sg13g2_nor2_1 _19768_ (.A(_10656_),
    .B(_10693_),
    .Y(_10694_));
 sg13g2_nor2_1 _19769_ (.A(net518),
    .B(net854),
    .Y(_10695_));
 sg13g2_a21oi_1 _19770_ (.A1(_10694_),
    .A2(_10695_),
    .Y(_10696_),
    .B1(_10283_));
 sg13g2_xor2_1 _19771_ (.B(net528),
    .A(net857),
    .X(_10697_));
 sg13g2_nand3_1 _19772_ (.B(_10634_),
    .C(net258),
    .A(net532),
    .Y(_10698_));
 sg13g2_o21ai_1 _19773_ (.B1(_10698_),
    .Y(_10699_),
    .A1(net532),
    .A2(_10697_));
 sg13g2_xnor2_1 _19774_ (.Y(_10700_),
    .A(net258),
    .B(_10608_));
 sg13g2_nand2_1 _19775_ (.Y(_10701_),
    .A(_10688_),
    .B(_10700_));
 sg13g2_o21ai_1 _19776_ (.B1(_10701_),
    .Y(_10702_),
    .A1(_10688_),
    .A2(_10699_));
 sg13g2_nor3_1 _19777_ (.A(net507),
    .B(_10687_),
    .C(_10693_),
    .Y(_10703_));
 sg13g2_a221oi_1 _19778_ (.B2(_10702_),
    .C1(_10703_),
    .B1(_10696_),
    .A1(_10657_),
    .Y(_10704_),
    .A2(_10692_));
 sg13g2_inv_2 _19779_ (.Y(_10705_),
    .A(_10685_));
 sg13g2_xnor2_1 _19780_ (.Y(_10706_),
    .A(_10705_),
    .B(_10335_));
 sg13g2_xnor2_1 _19781_ (.Y(_10707_),
    .A(_10608_),
    .B(_10706_));
 sg13g2_buf_2 _19782_ (.A(_10707_),
    .X(_10708_));
 sg13g2_xnor2_1 _19783_ (.Y(_10709_),
    .A(net1112),
    .B(_10708_));
 sg13g2_inv_1 _19784_ (.Y(_10710_),
    .A(_10709_));
 sg13g2_o21ai_1 _19785_ (.B1(_10595_),
    .Y(_10711_),
    .A1(net1108),
    .A2(_10709_));
 sg13g2_o21ai_1 _19786_ (.B1(_10711_),
    .Y(_10712_),
    .A1(net856),
    .A2(_10710_));
 sg13g2_a21oi_1 _19787_ (.A1(net258),
    .A2(_10687_),
    .Y(_10713_),
    .B1(_10689_));
 sg13g2_nand2_1 _19788_ (.Y(_10714_),
    .A(_10693_),
    .B(_10695_));
 sg13g2_o21ai_1 _19789_ (.B1(_10714_),
    .Y(_10715_),
    .A1(_10282_),
    .A2(_10713_));
 sg13g2_buf_1 _19790_ (.A(net854),
    .X(_10716_));
 sg13g2_a21oi_1 _19791_ (.A1(net532),
    .A2(_10634_),
    .Y(_10717_),
    .B1(net258));
 sg13g2_nor4_1 _19792_ (.A(net249),
    .B(_10716_),
    .C(_10282_),
    .D(_10717_),
    .Y(_10718_));
 sg13g2_a21oi_1 _19793_ (.A1(_10615_),
    .A2(_10715_),
    .Y(_10719_),
    .B1(_10718_));
 sg13g2_nand2_1 _19794_ (.Y(_10720_),
    .A(net119),
    .B(_10719_));
 sg13g2_a21o_1 _19795_ (.A2(_10712_),
    .A1(_10704_),
    .B1(_10720_),
    .X(_10721_));
 sg13g2_xnor2_1 _19796_ (.Y(_10722_),
    .A(net1107),
    .B(_10344_));
 sg13g2_xor2_1 _19797_ (.B(_10722_),
    .A(_10708_),
    .X(_10723_));
 sg13g2_nand2_1 _19798_ (.Y(_10724_),
    .A(net119),
    .B(_10723_));
 sg13g2_nor2_1 _19799_ (.A(net856),
    .B(_10283_),
    .Y(_10725_));
 sg13g2_nand2_1 _19800_ (.Y(_10726_),
    .A(_10595_),
    .B(_10289_));
 sg13g2_a21o_1 _19801_ (.A2(_10726_),
    .A1(_10708_),
    .B1(_10253_),
    .X(_10727_));
 sg13g2_nor2_1 _19802_ (.A(net855),
    .B(_10289_),
    .Y(_10728_));
 sg13g2_a21oi_1 _19803_ (.A1(_10650_),
    .A2(_10289_),
    .Y(_10729_),
    .B1(_10595_));
 sg13g2_a21oi_1 _19804_ (.A1(_10708_),
    .A2(_10728_),
    .Y(_10730_),
    .B1(_10729_));
 sg13g2_a21oi_1 _19805_ (.A1(_10727_),
    .A2(_10730_),
    .Y(_10731_),
    .B1(_10641_));
 sg13g2_a221oi_1 _19806_ (.B2(_10708_),
    .C1(_10731_),
    .B1(_10725_),
    .A1(net868),
    .Y(_10732_),
    .A2(_10710_));
 sg13g2_nor2_1 _19807_ (.A(net166),
    .B(_10719_),
    .Y(_10733_));
 sg13g2_a22oi_1 _19808_ (.Y(_10734_),
    .B1(_10732_),
    .B2(_10733_),
    .A2(_10724_),
    .A1(net250));
 sg13g2_nand3_1 _19809_ (.B(_10721_),
    .C(_10734_),
    .A(net39),
    .Y(_10735_));
 sg13g2_a21oi_1 _19810_ (.A1(_10681_),
    .A2(_10735_),
    .Y(_00398_),
    .B1(net523));
 sg13g2_o21ai_1 _19811_ (.B1(net256),
    .Y(_10736_),
    .A1(net258),
    .A2(_10705_));
 sg13g2_buf_1 _19812_ (.A(\grid.cell_23_2.se ),
    .X(_10737_));
 sg13g2_buf_1 _19813_ (.A(_10737_),
    .X(_10738_));
 sg13g2_inv_2 _19814_ (.Y(_10739_),
    .A(net853));
 sg13g2_nand2_1 _19815_ (.Y(_10740_),
    .A(_10739_),
    .B(net515));
 sg13g2_nor2_1 _19816_ (.A(_10047_),
    .B(_10740_),
    .Y(_10741_));
 sg13g2_nor2_1 _19817_ (.A(net258),
    .B(_10027_),
    .Y(_10742_));
 sg13g2_xnor2_1 _19818_ (.Y(_10743_),
    .A(_10737_),
    .B(_10352_));
 sg13g2_buf_2 _19819_ (.A(_10743_),
    .X(_10744_));
 sg13g2_nor2_1 _19820_ (.A(_09937_),
    .B(_10744_),
    .Y(_10745_));
 sg13g2_buf_1 _19821_ (.A(_10738_),
    .X(_10746_));
 sg13g2_a21oi_1 _19822_ (.A1(net504),
    .A2(net516),
    .Y(_10747_),
    .B1(net527));
 sg13g2_o21ai_1 _19823_ (.B1(net1115),
    .Y(_10748_),
    .A1(_10745_),
    .A2(_10747_));
 sg13g2_o21ai_1 _19824_ (.B1(_10748_),
    .Y(_10749_),
    .A1(_10740_),
    .A2(_10742_));
 sg13g2_a22oi_1 _19825_ (.Y(_10750_),
    .B1(_10749_),
    .B2(_10705_),
    .A2(_10741_),
    .A1(_10736_));
 sg13g2_xnor2_1 _19826_ (.Y(_10751_),
    .A(_09977_),
    .B(_10744_));
 sg13g2_xnor2_1 _19827_ (.Y(_10752_),
    .A(_09920_),
    .B(_10685_));
 sg13g2_xnor2_1 _19828_ (.Y(_10753_),
    .A(_10751_),
    .B(_10752_));
 sg13g2_and2_1 _19829_ (.A(_10383_),
    .B(_10753_),
    .X(_10754_));
 sg13g2_buf_1 _19830_ (.A(_10754_),
    .X(_10755_));
 sg13g2_xnor2_1 _19831_ (.Y(_10756_),
    .A(net866),
    .B(_10753_));
 sg13g2_buf_1 _19832_ (.A(_10756_),
    .X(_10757_));
 sg13g2_buf_1 _19833_ (.A(_00195_),
    .X(_10758_));
 sg13g2_buf_1 _19834_ (.A(_10758_),
    .X(_10759_));
 sg13g2_a21o_1 _19835_ (.A2(_10757_),
    .A1(_09947_),
    .B1(net852),
    .X(_10760_));
 sg13g2_o21ai_1 _19836_ (.B1(_10757_),
    .Y(_10761_),
    .A1(net852),
    .A2(_10755_));
 sg13g2_nor3_1 _19837_ (.A(net852),
    .B(_10757_),
    .C(_10755_),
    .Y(_10762_));
 sg13g2_a221oi_1 _19838_ (.B2(net529),
    .C1(_10762_),
    .B1(_10761_),
    .A1(_10755_),
    .Y(_10763_),
    .A2(_10760_));
 sg13g2_or2_1 _19839_ (.X(_10764_),
    .B(_10763_),
    .A(_10750_));
 sg13g2_nand2_1 _19840_ (.Y(_10765_),
    .A(_10759_),
    .B(_10757_));
 sg13g2_o21ai_1 _19841_ (.B1(_09947_),
    .Y(_10766_),
    .A1(_10759_),
    .A2(_10757_));
 sg13g2_buf_1 _19842_ (.A(net505),
    .X(_10767_));
 sg13g2_nor3_1 _19843_ (.A(net258),
    .B(net240),
    .C(_10354_),
    .Y(_10768_));
 sg13g2_nand2_1 _19844_ (.Y(_10769_),
    .A(net853),
    .B(net864));
 sg13g2_nor2_1 _19845_ (.A(_09943_),
    .B(_10769_),
    .Y(_10770_));
 sg13g2_o21ai_1 _19846_ (.B1(net527),
    .Y(_10771_),
    .A1(_10745_),
    .A2(_10770_));
 sg13g2_o21ai_1 _19847_ (.B1(_10771_),
    .Y(_10772_),
    .A1(net1115),
    .A2(_10769_));
 sg13g2_a21o_1 _19848_ (.A2(_10772_),
    .A1(net240),
    .B1(_10755_),
    .X(_10773_));
 sg13g2_a221oi_1 _19849_ (.B2(net504),
    .C1(_10773_),
    .B1(_10768_),
    .A1(_10765_),
    .Y(_10774_),
    .A2(_10766_));
 sg13g2_a21oi_1 _19850_ (.A1(_10750_),
    .A2(_10774_),
    .Y(_10775_),
    .B1(net103));
 sg13g2_xnor2_1 _19851_ (.Y(_10776_),
    .A(_10608_),
    .B(_10757_));
 sg13g2_o21ai_1 _19852_ (.B1(_10311_),
    .Y(_10777_),
    .A1(net166),
    .A2(_10776_));
 sg13g2_nand3_1 _19853_ (.B(net39),
    .C(_10777_),
    .A(net714),
    .Y(_10778_));
 sg13g2_a21oi_1 _19854_ (.A1(_10764_),
    .A2(_10775_),
    .Y(_10779_),
    .B1(_10778_));
 sg13g2_nand3_1 _19855_ (.B(net33),
    .C(_10606_),
    .A(net334),
    .Y(_10780_));
 sg13g2_nand2b_1 _19856_ (.Y(_00399_),
    .B(_10780_),
    .A_N(_10779_));
 sg13g2_nand3_1 _19857_ (.B(net104),
    .C(net39),
    .A(_10363_),
    .Y(_10781_));
 sg13g2_o21ai_1 _19858_ (.B1(_10781_),
    .Y(_10782_),
    .A1(net48),
    .A2(net39));
 sg13g2_buf_1 _19859_ (.A(\grid.cell_23_3.se ),
    .X(_10783_));
 sg13g2_buf_1 _19860_ (.A(_10783_),
    .X(_10784_));
 sg13g2_buf_1 _19861_ (.A(net851),
    .X(_10785_));
 sg13g2_nand2_1 _19862_ (.Y(_10786_),
    .A(net862),
    .B(_10738_));
 sg13g2_nor2_1 _19863_ (.A(net527),
    .B(_10786_),
    .Y(_10787_));
 sg13g2_xnor2_1 _19864_ (.Y(_10788_),
    .A(net862),
    .B(net504));
 sg13g2_nor2_1 _19865_ (.A(_10027_),
    .B(_10788_),
    .Y(_10789_));
 sg13g2_o21ai_1 _19866_ (.B1(net525),
    .Y(_10790_),
    .A1(_10787_),
    .A2(_10789_));
 sg13g2_o21ai_1 _19867_ (.B1(_10790_),
    .Y(_10791_),
    .A1(_10075_),
    .A2(_10786_));
 sg13g2_nand2_1 _19868_ (.Y(_10792_),
    .A(net503),
    .B(_10791_));
 sg13g2_nand2_1 _19869_ (.Y(_10793_),
    .A(net525),
    .B(net256));
 sg13g2_or3_1 _19870_ (.A(net503),
    .B(_10793_),
    .C(_10786_),
    .X(_10794_));
 sg13g2_nand4_1 _19871_ (.B(_10683_),
    .C(_10792_),
    .A(net1060),
    .Y(_10795_),
    .D(_10794_));
 sg13g2_buf_1 _19872_ (.A(_00192_),
    .X(_10796_));
 sg13g2_xnor2_1 _19873_ (.Y(_10797_),
    .A(_10783_),
    .B(_10398_));
 sg13g2_xnor2_1 _19874_ (.Y(_10798_),
    .A(net1116),
    .B(_10797_));
 sg13g2_xnor2_1 _19875_ (.Y(_10799_),
    .A(net853),
    .B(net874));
 sg13g2_xnor2_1 _19876_ (.Y(_10800_),
    .A(_10798_),
    .B(_10799_));
 sg13g2_nand2b_1 _19877_ (.Y(_10801_),
    .B(_10800_),
    .A_N(_10405_));
 sg13g2_nor3_1 _19878_ (.A(_10796_),
    .B(_10335_),
    .C(_10801_),
    .Y(_10802_));
 sg13g2_xor2_1 _19879_ (.B(_10800_),
    .A(_10706_),
    .X(_10803_));
 sg13g2_a21oi_1 _19880_ (.A1(net70),
    .A2(_10803_),
    .Y(_10804_),
    .B1(net248));
 sg13g2_inv_1 _19881_ (.Y(_10805_),
    .A(_10783_));
 sg13g2_buf_1 _19882_ (.A(_10805_),
    .X(_10806_));
 sg13g2_nand4_1 _19883_ (.B(_10454_),
    .C(_10739_),
    .A(net502),
    .Y(_10807_),
    .D(net525));
 sg13g2_nand2_1 _19884_ (.Y(_10808_),
    .A(_10784_),
    .B(_10746_));
 sg13g2_nand3_1 _19885_ (.B(_10807_),
    .C(_10808_),
    .A(_10786_),
    .Y(_10809_));
 sg13g2_a221oi_1 _19886_ (.B2(_10027_),
    .C1(_10809_),
    .B1(net254),
    .A1(net503),
    .Y(_10810_),
    .A2(net247));
 sg13g2_nor3_1 _19887_ (.A(_10785_),
    .B(_10401_),
    .C(_10746_),
    .Y(_10811_));
 sg13g2_a22oi_1 _19888_ (.Y(_10812_),
    .B1(_10811_),
    .B2(_10793_),
    .A2(_10810_),
    .A1(_10075_));
 sg13g2_inv_1 _19889_ (.Y(_10813_),
    .A(_10796_));
 sg13g2_xnor2_1 _19890_ (.Y(_10814_),
    .A(net517),
    .B(_10800_));
 sg13g2_o21ai_1 _19891_ (.B1(_10814_),
    .Y(_10815_),
    .A1(net257),
    .A2(_10813_));
 sg13g2_nand2_1 _19892_ (.Y(_10816_),
    .A(net257),
    .B(_10813_));
 sg13g2_nand3_1 _19893_ (.B(_10815_),
    .C(_10816_),
    .A(_10801_),
    .Y(_10817_));
 sg13g2_xnor2_1 _19894_ (.Y(_10818_),
    .A(_10812_),
    .B(_10817_));
 sg13g2_nor4_1 _19895_ (.A(_10795_),
    .B(_10802_),
    .C(_10804_),
    .D(_10818_),
    .Y(_10819_));
 sg13g2_a21o_1 _19896_ (.A2(_10782_),
    .A1(net317),
    .B1(_10819_),
    .X(_00400_));
 sg13g2_buf_2 _19897_ (.A(\grid.cell_23_4.se ),
    .X(_10820_));
 sg13g2_xnor2_1 _19898_ (.Y(_10821_),
    .A(_10820_),
    .B(_10430_));
 sg13g2_xnor2_1 _19899_ (.Y(_10822_),
    .A(net871),
    .B(_10821_));
 sg13g2_xnor2_1 _19900_ (.Y(_10823_),
    .A(net851),
    .B(net1116));
 sg13g2_xnor2_1 _19901_ (.Y(_10824_),
    .A(_10822_),
    .B(_10823_));
 sg13g2_buf_1 _19902_ (.A(_10824_),
    .X(_10825_));
 sg13g2_xnor2_1 _19903_ (.Y(_10826_),
    .A(_10751_),
    .B(_10825_));
 sg13g2_o21ai_1 _19904_ (.B1(_10454_),
    .Y(_10827_),
    .A1(net166),
    .A2(_10826_));
 sg13g2_nand2_1 _19905_ (.Y(_10828_),
    .A(net39),
    .B(_10827_));
 sg13g2_o21ai_1 _19906_ (.B1(_10828_),
    .Y(_10829_),
    .A1(net47),
    .A2(net39));
 sg13g2_buf_1 _19907_ (.A(_10820_),
    .X(_10830_));
 sg13g2_buf_1 _19908_ (.A(_10830_),
    .X(_10831_));
 sg13g2_nor4_1 _19909_ (.A(_10831_),
    .B(net246),
    .C(net503),
    .D(net244),
    .Y(_10832_));
 sg13g2_inv_2 _19910_ (.Y(_10833_),
    .A(net861));
 sg13g2_nor2_2 _19911_ (.A(_10833_),
    .B(_10806_),
    .Y(_10834_));
 sg13g2_nor2_1 _19912_ (.A(net244),
    .B(net254),
    .Y(_10835_));
 sg13g2_o21ai_1 _19913_ (.B1(net850),
    .Y(_10836_),
    .A1(net861),
    .A2(net851));
 sg13g2_nand2_1 _19914_ (.Y(_10837_),
    .A(net1114),
    .B(_10836_));
 sg13g2_nor4_1 _19915_ (.A(_10832_),
    .B(_10834_),
    .C(_10835_),
    .D(_10837_),
    .Y(_10838_));
 sg13g2_inv_1 _19916_ (.Y(_10839_),
    .A(_10820_));
 sg13g2_buf_1 _19917_ (.A(_10839_),
    .X(_10840_));
 sg13g2_nand3_1 _19918_ (.B(_10833_),
    .C(net502),
    .A(net500),
    .Y(_10841_));
 sg13g2_buf_1 _19919_ (.A(_10841_),
    .X(_10842_));
 sg13g2_a21oi_1 _19920_ (.A1(net255),
    .A2(net254),
    .Y(_10843_),
    .B1(_10842_));
 sg13g2_buf_1 _19921_ (.A(_00056_),
    .X(_10844_));
 sg13g2_a21o_1 _19922_ (.A2(_10825_),
    .A1(net515),
    .B1(net527),
    .X(_10845_));
 sg13g2_o21ai_1 _19923_ (.B1(_10825_),
    .Y(_10846_),
    .A1(net1111),
    .A2(net256));
 sg13g2_a221oi_1 _19924_ (.B2(_10363_),
    .C1(_10355_),
    .B1(_10846_),
    .A1(_10447_),
    .Y(_10847_),
    .A2(_10845_));
 sg13g2_xnor2_1 _19925_ (.Y(_10848_),
    .A(_10392_),
    .B(_10825_));
 sg13g2_nor2b_1 _19926_ (.A(net1111),
    .B_N(_10825_),
    .Y(_10849_));
 sg13g2_a22oi_1 _19927_ (.Y(_10850_),
    .B1(_10849_),
    .B2(_10844_),
    .A2(_10848_),
    .A1(net256));
 sg13g2_o21ai_1 _19928_ (.B1(_10850_),
    .Y(_10851_),
    .A1(_10844_),
    .A2(_10847_));
 sg13g2_o21ai_1 _19929_ (.B1(_10851_),
    .Y(_10852_),
    .A1(_10838_),
    .A2(_10843_));
 sg13g2_inv_1 _19930_ (.Y(_10853_),
    .A(_10844_));
 sg13g2_o21ai_1 _19931_ (.B1(_10848_),
    .Y(_10854_),
    .A1(_10853_),
    .A2(net256));
 sg13g2_nand3_1 _19932_ (.B(net526),
    .C(_10834_),
    .A(net850),
    .Y(_10855_));
 sg13g2_a21oi_1 _19933_ (.A1(_10842_),
    .A2(_10855_),
    .Y(_10856_),
    .B1(net525));
 sg13g2_nor2_1 _19934_ (.A(net1114),
    .B(net500),
    .Y(_10857_));
 sg13g2_a22oi_1 _19935_ (.Y(_10858_),
    .B1(_10834_),
    .B2(_10857_),
    .A2(net256),
    .A1(_10853_));
 sg13g2_nand2b_1 _19936_ (.Y(_10859_),
    .B(_10858_),
    .A_N(_10856_));
 sg13g2_nor2b_1 _19937_ (.A(_10834_),
    .B_N(_10836_),
    .Y(_10860_));
 sg13g2_a21o_1 _19938_ (.A2(_10834_),
    .A1(net1114),
    .B1(net244),
    .X(_10861_));
 sg13g2_nand2_1 _19939_ (.Y(_10862_),
    .A(net513),
    .B(net244));
 sg13g2_nand3_1 _19940_ (.B(_10862_),
    .C(_10842_),
    .A(net525),
    .Y(_10863_));
 sg13g2_a221oi_1 _19941_ (.B2(net501),
    .C1(_10863_),
    .B1(_10861_),
    .A1(_10133_),
    .Y(_10864_),
    .A2(_10860_));
 sg13g2_nand2_1 _19942_ (.Y(_10865_),
    .A(net1114),
    .B(_10860_));
 sg13g2_a21oi_1 _19943_ (.A1(_10842_),
    .A2(_10865_),
    .Y(_10866_),
    .B1(net255));
 sg13g2_nor4_1 _19944_ (.A(_10849_),
    .B(_10859_),
    .C(_10864_),
    .D(_10866_),
    .Y(_10867_));
 sg13g2_nand2_1 _19945_ (.Y(_10868_),
    .A(_10854_),
    .B(_10867_));
 sg13g2_nand4_1 _19946_ (.B(_10684_),
    .C(_10852_),
    .A(net78),
    .Y(_10869_),
    .D(_10868_));
 sg13g2_and3_1 _19947_ (.X(_00401_),
    .A(net317),
    .B(_10829_),
    .C(_10869_));
 sg13g2_buf_2 _19948_ (.A(\grid.cell_23_5.se ),
    .X(_10870_));
 sg13g2_inv_1 _19949_ (.Y(_10871_),
    .A(_10870_));
 sg13g2_buf_1 _19950_ (.A(_10871_),
    .X(_10872_));
 sg13g2_nand2_1 _19951_ (.Y(_10873_),
    .A(net500),
    .B(net499));
 sg13g2_nor3_1 _19952_ (.A(net245),
    .B(_10161_),
    .C(_10873_),
    .Y(_10874_));
 sg13g2_buf_2 _19953_ (.A(_10870_),
    .X(_10875_));
 sg13g2_nand2_1 _19954_ (.Y(_10876_),
    .A(net850),
    .B(net849));
 sg13g2_o21ai_1 _19955_ (.B1(_10876_),
    .Y(_10877_),
    .A1(_10161_),
    .A2(net255));
 sg13g2_buf_1 _19956_ (.A(net849),
    .X(_10878_));
 sg13g2_o21ai_1 _19957_ (.B1(_10496_),
    .Y(_10879_),
    .A1(_10831_),
    .A2(net498));
 sg13g2_nand2_1 _19958_ (.Y(_10880_),
    .A(net869),
    .B(_10879_));
 sg13g2_nor3_1 _19959_ (.A(_10874_),
    .B(_10877_),
    .C(_10880_),
    .Y(_10881_));
 sg13g2_nor2_1 _19960_ (.A(_10502_),
    .B(net498),
    .Y(_10882_));
 sg13g2_and3_1 _19961_ (.X(_10883_),
    .A(net500),
    .B(_10121_),
    .C(_10882_));
 sg13g2_buf_2 _19962_ (.A(_00088_),
    .X(_10884_));
 sg13g2_xor2_1 _19963_ (.B(_10113_),
    .A(_10870_),
    .X(_10885_));
 sg13g2_xnor2_1 _19964_ (.Y(_10886_),
    .A(_10820_),
    .B(net871));
 sg13g2_xnor2_1 _19965_ (.Y(_10887_),
    .A(_10885_),
    .B(_10886_));
 sg13g2_xnor2_1 _19966_ (.Y(_10888_),
    .A(net860),
    .B(_10887_));
 sg13g2_buf_1 _19967_ (.A(_10888_),
    .X(_10889_));
 sg13g2_o21ai_1 _19968_ (.B1(_10023_),
    .Y(_10890_),
    .A1(net247),
    .A2(_10889_));
 sg13g2_a21o_1 _19969_ (.A2(_10023_),
    .A1(_10505_),
    .B1(_10889_),
    .X(_10891_));
 sg13g2_a221oi_1 _19970_ (.B2(net247),
    .C1(_10403_),
    .B1(_10891_),
    .A1(_10467_),
    .Y(_10892_),
    .A2(_10890_));
 sg13g2_xnor2_1 _19971_ (.Y(_10893_),
    .A(_10401_),
    .B(_10889_));
 sg13g2_nor2_1 _19972_ (.A(_10467_),
    .B(_10889_),
    .Y(_10894_));
 sg13g2_a22oi_1 _19973_ (.Y(_10895_),
    .B1(_10894_),
    .B2(_10884_),
    .A2(_10893_),
    .A1(net254));
 sg13g2_o21ai_1 _19974_ (.B1(_10895_),
    .Y(_10896_),
    .A1(_10884_),
    .A2(_10892_));
 sg13g2_o21ai_1 _19975_ (.B1(_10896_),
    .Y(_10897_),
    .A1(_10881_),
    .A2(_10883_));
 sg13g2_inv_1 _19976_ (.Y(_10898_),
    .A(_10884_));
 sg13g2_o21ai_1 _19977_ (.B1(_10893_),
    .Y(_10899_),
    .A1(_10898_),
    .A2(net254));
 sg13g2_nand2_1 _19978_ (.Y(_10900_),
    .A(net850),
    .B(net524));
 sg13g2_o21ai_1 _19979_ (.B1(_10900_),
    .Y(_10901_),
    .A1(_10830_),
    .A2(net499));
 sg13g2_nand3_1 _19980_ (.B(net526),
    .C(_10901_),
    .A(_10164_),
    .Y(_10902_));
 sg13g2_o21ai_1 _19981_ (.B1(_10902_),
    .Y(_10903_),
    .A1(net255),
    .A2(_10873_));
 sg13g2_nand2_1 _19982_ (.Y(_10904_),
    .A(_10482_),
    .B(_10903_));
 sg13g2_nor2_2 _19983_ (.A(net500),
    .B(_10872_),
    .Y(_10905_));
 sg13g2_nand2_1 _19984_ (.Y(_10906_),
    .A(_10121_),
    .B(_10876_));
 sg13g2_o21ai_1 _19985_ (.B1(_10906_),
    .Y(_10907_),
    .A1(_10164_),
    .A2(_10873_));
 sg13g2_a21oi_1 _19986_ (.A1(net869),
    .A2(_10905_),
    .Y(_10908_),
    .B1(_10907_));
 sg13g2_nand2_1 _19987_ (.Y(_10909_),
    .A(_10496_),
    .B(_10908_));
 sg13g2_nand2_1 _19988_ (.Y(_10910_),
    .A(_10486_),
    .B(net244));
 sg13g2_o21ai_1 _19989_ (.B1(_10910_),
    .Y(_10911_),
    .A1(net869),
    .A2(net244));
 sg13g2_nand3_1 _19990_ (.B(_10905_),
    .C(_10911_),
    .A(net142),
    .Y(_10912_));
 sg13g2_nand2_1 _19991_ (.Y(_10913_),
    .A(_10898_),
    .B(net254));
 sg13g2_nand4_1 _19992_ (.B(_10909_),
    .C(_10912_),
    .A(_10904_),
    .Y(_10914_),
    .D(_10913_));
 sg13g2_o21ai_1 _19993_ (.B1(_10873_),
    .Y(_10915_),
    .A1(net511),
    .A2(_10905_));
 sg13g2_a22oi_1 _19994_ (.Y(_10916_),
    .B1(_10915_),
    .B2(net869),
    .A2(_10882_),
    .A1(_10840_));
 sg13g2_nor2_1 _19995_ (.A(net142),
    .B(_10916_),
    .Y(_10917_));
 sg13g2_nor3_1 _19996_ (.A(_10894_),
    .B(_10914_),
    .C(_10917_),
    .Y(_10918_));
 sg13g2_nand2_1 _19997_ (.Y(_10919_),
    .A(net83),
    .B(_10684_));
 sg13g2_a21oi_1 _19998_ (.A1(_10899_),
    .A2(_10918_),
    .Y(_10920_),
    .B1(_10919_));
 sg13g2_xor2_1 _19999_ (.B(_10889_),
    .A(_10798_),
    .X(_10921_));
 sg13g2_o21ai_1 _20000_ (.B1(_10833_),
    .Y(_10922_),
    .A1(net105),
    .A2(_10921_));
 sg13g2_o21ai_1 _20001_ (.B1(net668),
    .Y(_10923_),
    .A1(_10606_),
    .A2(_10922_));
 sg13g2_a221oi_1 _20002_ (.B2(_10920_),
    .C1(_10923_),
    .B1(_10897_),
    .A1(net43),
    .Y(_00402_),
    .A2(_10606_));
 sg13g2_buf_2 _20003_ (.A(_00151_),
    .X(_10924_));
 sg13g2_and2_1 _20004_ (.A(net859),
    .B(_10870_),
    .X(_10925_));
 sg13g2_buf_1 _20005_ (.A(_10925_),
    .X(_10926_));
 sg13g2_nor2b_1 _20006_ (.A(_10924_),
    .B_N(_10926_),
    .Y(_10927_));
 sg13g2_nand2_1 _20007_ (.Y(_10928_),
    .A(net524),
    .B(net530));
 sg13g2_nor3_1 _20008_ (.A(_10924_),
    .B(net867),
    .C(net849),
    .Y(_10929_));
 sg13g2_nor3_1 _20009_ (.A(_10928_),
    .B(_10926_),
    .C(_10929_),
    .Y(_10930_));
 sg13g2_or2_1 _20010_ (.X(_10931_),
    .B(_10930_),
    .A(_10927_));
 sg13g2_nor2_1 _20011_ (.A(net867),
    .B(net849),
    .Y(_10932_));
 sg13g2_nand2_1 _20012_ (.Y(_10933_),
    .A(net506),
    .B(_10932_));
 sg13g2_nand4_1 _20013_ (.B(net519),
    .C(net498),
    .A(net508),
    .Y(_10934_),
    .D(net531));
 sg13g2_nand3_1 _20014_ (.B(_10933_),
    .C(_10934_),
    .A(_10161_),
    .Y(_10935_));
 sg13g2_o21ai_1 _20015_ (.B1(_10276_),
    .Y(_10936_),
    .A1(net519),
    .A2(_10871_));
 sg13g2_nand3_1 _20016_ (.B(net506),
    .C(_10936_),
    .A(_10924_),
    .Y(_10937_));
 sg13g2_nand3b_1 _20017_ (.B(net498),
    .C(_10292_),
    .Y(_10938_),
    .A_N(_10924_));
 sg13g2_nand3_1 _20018_ (.B(_10937_),
    .C(_10938_),
    .A(net253),
    .Y(_10939_));
 sg13g2_nor2_1 _20019_ (.A(_10635_),
    .B(_10926_),
    .Y(_10940_));
 sg13g2_o21ai_1 _20020_ (.B1(_10924_),
    .Y(_10941_),
    .A1(_10932_),
    .A2(_10940_));
 sg13g2_a21oi_1 _20021_ (.A1(_10933_),
    .A2(_10941_),
    .Y(_10942_),
    .B1(net252));
 sg13g2_a221oi_1 _20022_ (.B2(_10939_),
    .C1(_10942_),
    .B1(_10935_),
    .A1(net241),
    .Y(_10943_),
    .A2(_10931_));
 sg13g2_buf_2 _20023_ (.A(_00120_),
    .X(_10944_));
 sg13g2_nand2_1 _20024_ (.Y(_10945_),
    .A(_10944_),
    .B(net244));
 sg13g2_xor2_1 _20025_ (.B(_10885_),
    .A(net1118),
    .X(_10946_));
 sg13g2_xor2_1 _20026_ (.B(_10946_),
    .A(_10610_),
    .X(_10947_));
 sg13g2_xnor2_1 _20027_ (.Y(_10948_),
    .A(net513),
    .B(_10947_));
 sg13g2_nand2b_1 _20028_ (.Y(_10949_),
    .B(net526),
    .A_N(_10944_));
 sg13g2_o21ai_1 _20029_ (.B1(_10949_),
    .Y(_10950_),
    .A1(net1110),
    .A2(_10947_));
 sg13g2_a21oi_1 _20030_ (.A1(_10945_),
    .A2(_10948_),
    .Y(_10951_),
    .B1(_10950_));
 sg13g2_xor2_1 _20031_ (.B(_10951_),
    .A(_10943_),
    .X(_10952_));
 sg13g2_xnor2_1 _20032_ (.Y(_10953_),
    .A(_10822_),
    .B(_10947_));
 sg13g2_nand2_1 _20033_ (.Y(_10954_),
    .A(net849),
    .B(net524));
 sg13g2_nand2_1 _20034_ (.Y(_10955_),
    .A(net519),
    .B(_10885_));
 sg13g2_o21ai_1 _20035_ (.B1(_10955_),
    .Y(_10956_),
    .A1(net519),
    .A2(_10954_));
 sg13g2_a21o_1 _20036_ (.A2(_10956_),
    .A1(net252),
    .B1(_10927_),
    .X(_10957_));
 sg13g2_nor2_1 _20037_ (.A(_10928_),
    .B(_10623_),
    .Y(_10958_));
 sg13g2_nand2b_1 _20038_ (.Y(_10959_),
    .B(_10443_),
    .A_N(_10944_));
 sg13g2_nor3_1 _20039_ (.A(net1110),
    .B(_10947_),
    .C(_10959_),
    .Y(_10960_));
 sg13g2_a221oi_1 _20040_ (.B2(_10878_),
    .C1(_10960_),
    .B1(_10958_),
    .A1(net241),
    .Y(_10961_),
    .A2(_10957_));
 sg13g2_o21ai_1 _20041_ (.B1(_10961_),
    .Y(_10962_),
    .A1(net245),
    .A2(_10953_));
 sg13g2_nor3_1 _20042_ (.A(net103),
    .B(_10952_),
    .C(_10962_),
    .Y(_10963_));
 sg13g2_a21oi_1 _20043_ (.A1(net245),
    .A2(net73),
    .Y(_10964_),
    .B1(_10963_));
 sg13g2_o21ai_1 _20044_ (.B1(net522),
    .Y(_10965_),
    .A1(net31),
    .A2(net39));
 sg13g2_a21oi_1 _20045_ (.A1(net39),
    .A2(_10964_),
    .Y(_00403_),
    .B1(_10965_));
 sg13g2_nor2b_1 _20046_ (.A(_09522_),
    .B_N(_05748_),
    .Y(_10966_));
 sg13g2_a22oi_1 _20047_ (.Y(_10967_),
    .B1(net76),
    .B2(_10966_),
    .A2(net69),
    .A1(net243));
 sg13g2_nand2_1 _20048_ (.Y(_10968_),
    .A(net511),
    .B(_10878_));
 sg13g2_nand2_1 _20049_ (.Y(_10969_),
    .A(net510),
    .B(_10885_));
 sg13g2_o21ai_1 _20050_ (.B1(_10969_),
    .Y(_10970_),
    .A1(net511),
    .A2(_10954_));
 sg13g2_nand2_1 _20051_ (.Y(_10971_),
    .A(net252),
    .B(_10970_));
 sg13g2_o21ai_1 _20052_ (.B1(_10971_),
    .Y(_10972_),
    .A1(_10924_),
    .A2(_10968_));
 sg13g2_o21ai_1 _20053_ (.B1(net506),
    .Y(_10973_),
    .A1(_10928_),
    .A2(_10968_));
 sg13g2_o21ai_1 _20054_ (.B1(_10973_),
    .Y(_10974_),
    .A1(_10665_),
    .A2(_10972_));
 sg13g2_xor2_1 _20055_ (.B(_10469_),
    .A(_10609_),
    .X(_10975_));
 sg13g2_xor2_1 _20056_ (.B(_10975_),
    .A(_10946_),
    .X(_10976_));
 sg13g2_nand4_1 _20057_ (.B(_10289_),
    .C(_10344_),
    .A(net856),
    .Y(_10977_),
    .D(_10976_));
 sg13g2_xnor2_1 _20058_ (.Y(_10978_),
    .A(_10722_),
    .B(_10976_));
 sg13g2_xnor2_1 _20059_ (.Y(_10979_),
    .A(net1112),
    .B(_10976_));
 sg13g2_a22oi_1 _20060_ (.Y(_10980_),
    .B1(_10289_),
    .B2(_10976_),
    .A2(net856),
    .A1(net868));
 sg13g2_o21ai_1 _20061_ (.B1(_10980_),
    .Y(_10981_),
    .A1(_10645_),
    .A2(_10979_));
 sg13g2_nand2_1 _20062_ (.Y(_10982_),
    .A(net512),
    .B(_10871_));
 sg13g2_o21ai_1 _20063_ (.B1(net849),
    .Y(_10983_),
    .A1(_10635_),
    .A2(_10486_));
 sg13g2_o21ai_1 _20064_ (.B1(_10983_),
    .Y(_10984_),
    .A1(_10621_),
    .A2(_10982_));
 sg13g2_a221oi_1 _20065_ (.B2(net252),
    .C1(_10984_),
    .B1(_10161_),
    .A1(net241),
    .Y(_10985_),
    .A2(net510));
 sg13g2_nor2_1 _20066_ (.A(_10189_),
    .B(_10982_),
    .Y(_10986_));
 sg13g2_a22oi_1 _20067_ (.Y(_10987_),
    .B1(_10986_),
    .B2(_10665_),
    .A2(_10985_),
    .A1(_10924_));
 sg13g2_xnor2_1 _20068_ (.Y(_10988_),
    .A(_10981_),
    .B(_10987_));
 sg13g2_a21oi_1 _20069_ (.A1(net520),
    .A2(_10978_),
    .Y(_10989_),
    .B1(_10988_));
 sg13g2_nand4_1 _20070_ (.B(_10974_),
    .C(_10977_),
    .A(net82),
    .Y(_10990_),
    .D(_10989_));
 sg13g2_a221oi_1 _20071_ (.B2(_10990_),
    .C1(net533),
    .B1(_10967_),
    .A1(_06471_),
    .Y(_00404_),
    .A2(_10966_));
 sg13g2_nand2b_1 _20072_ (.Y(_10991_),
    .B(_05180_),
    .A_N(_01903_));
 sg13g2_buf_2 _20073_ (.A(_10991_),
    .X(_10992_));
 sg13g2_or2_1 _20074_ (.X(_10993_),
    .B(_10992_),
    .A(_07600_));
 sg13g2_buf_1 _20075_ (.A(_10993_),
    .X(_10994_));
 sg13g2_nor2_1 _20076_ (.A(net176),
    .B(_10994_),
    .Y(_10995_));
 sg13g2_buf_2 _20077_ (.A(_10995_),
    .X(_10996_));
 sg13g2_nand2_1 _20078_ (.Y(_10997_),
    .A(net44),
    .B(_10996_));
 sg13g2_buf_1 _20079_ (.A(\grid.cell_24_0.se ),
    .X(_10998_));
 sg13g2_buf_1 _20080_ (.A(net1106),
    .X(_10999_));
 sg13g2_buf_1 _20081_ (.A(net848),
    .X(_11000_));
 sg13g2_buf_2 _20082_ (.A(\grid.cell_24_0.sw ),
    .X(_11001_));
 sg13g2_buf_1 _20083_ (.A(_11001_),
    .X(_11002_));
 sg13g2_and2_1 _20084_ (.A(net847),
    .B(_10609_),
    .X(_11003_));
 sg13g2_buf_1 _20085_ (.A(_11003_),
    .X(_11004_));
 sg13g2_xor2_1 _20086_ (.B(_10609_),
    .A(_11001_),
    .X(_11005_));
 sg13g2_nand2_1 _20087_ (.Y(_11006_),
    .A(net521),
    .B(_11005_));
 sg13g2_o21ai_1 _20088_ (.B1(_11006_),
    .Y(_11007_),
    .A1(net243),
    .A2(_11004_));
 sg13g2_nand2_1 _20089_ (.Y(_11008_),
    .A(net521),
    .B(net243));
 sg13g2_nor2_1 _20090_ (.A(net847),
    .B(net858),
    .Y(_11009_));
 sg13g2_buf_1 _20091_ (.A(_11009_),
    .X(_11010_));
 sg13g2_a22oi_1 _20092_ (.Y(_11011_),
    .B1(_11008_),
    .B2(_11010_),
    .A2(_11007_),
    .A1(net863));
 sg13g2_inv_1 _20093_ (.Y(_11012_),
    .A(net1106));
 sg13g2_buf_1 _20094_ (.A(_11012_),
    .X(_11013_));
 sg13g2_o21ai_1 _20095_ (.B1(net243),
    .Y(_11014_),
    .A1(net250),
    .A2(net496));
 sg13g2_nand3_1 _20096_ (.B(_11014_),
    .C(_11010_),
    .A(net863),
    .Y(_11015_));
 sg13g2_o21ai_1 _20097_ (.B1(_11015_),
    .Y(_11016_),
    .A1(net497),
    .A2(_11011_));
 sg13g2_buf_2 _20098_ (.A(_00199_),
    .X(_11017_));
 sg13g2_inv_1 _20099_ (.Y(_11018_),
    .A(_10758_));
 sg13g2_buf_1 _20100_ (.A(_11018_),
    .X(_11019_));
 sg13g2_nand2_1 _20101_ (.Y(_11020_),
    .A(net857),
    .B(net495));
 sg13g2_xnor2_1 _20102_ (.Y(_11021_),
    .A(_10247_),
    .B(net1106));
 sg13g2_xor2_1 _20103_ (.B(_11021_),
    .A(_11005_),
    .X(_11022_));
 sg13g2_xnor2_1 _20104_ (.Y(_11023_),
    .A(net520),
    .B(_11022_));
 sg13g2_a21o_1 _20105_ (.A2(net495),
    .A1(_10253_),
    .B1(_11023_),
    .X(_11024_));
 sg13g2_nor3_1 _20106_ (.A(net857),
    .B(net495),
    .C(_11023_),
    .Y(_11025_));
 sg13g2_a221oi_1 _20107_ (.B2(net507),
    .C1(_11025_),
    .B1(_11024_),
    .A1(net855),
    .Y(_11026_),
    .A2(_11020_));
 sg13g2_xnor2_1 _20108_ (.Y(_11027_),
    .A(net857),
    .B(_11023_));
 sg13g2_nor2_1 _20109_ (.A(net852),
    .B(_11023_),
    .Y(_11028_));
 sg13g2_a22oi_1 _20110_ (.Y(_11029_),
    .B1(_11028_),
    .B2(_11017_),
    .A2(_11027_),
    .A1(net855));
 sg13g2_o21ai_1 _20111_ (.B1(_11029_),
    .Y(_11030_),
    .A1(_11017_),
    .A2(_11026_));
 sg13g2_inv_1 _20112_ (.Y(_11031_),
    .A(_11017_));
 sg13g2_o21ai_1 _20113_ (.B1(_11027_),
    .Y(_11032_),
    .A1(net855),
    .A2(_11031_));
 sg13g2_nand2b_1 _20114_ (.Y(_11033_),
    .B(_10609_),
    .A_N(_11001_));
 sg13g2_buf_1 _20115_ (.A(_11033_),
    .X(_11034_));
 sg13g2_buf_1 _20116_ (.A(net847),
    .X(_11035_));
 sg13g2_o21ai_1 _20117_ (.B1(net494),
    .Y(_11036_),
    .A1(_10616_),
    .A2(net863));
 sg13g2_a21oi_1 _20118_ (.A1(_11034_),
    .A2(_11036_),
    .Y(_11037_),
    .B1(net243));
 sg13g2_inv_2 _20119_ (.Y(_11038_),
    .A(net847));
 sg13g2_mux2_1 _20120_ (.A0(net508),
    .A1(net520),
    .S(_11038_),
    .X(_11039_));
 sg13g2_nand2_1 _20121_ (.Y(_11040_),
    .A(_10383_),
    .B(_11010_));
 sg13g2_o21ai_1 _20122_ (.B1(_11040_),
    .Y(_11041_),
    .A1(net521),
    .A2(_11039_));
 sg13g2_o21ai_1 _20123_ (.B1(net848),
    .Y(_11042_),
    .A1(_11037_),
    .A2(_11041_));
 sg13g2_nand2_1 _20124_ (.Y(_11043_),
    .A(_11012_),
    .B(_11038_));
 sg13g2_nor2_1 _20125_ (.A(_11012_),
    .B(_11038_),
    .Y(_11044_));
 sg13g2_nand3_1 _20126_ (.B(net863),
    .C(_11044_),
    .A(net508),
    .Y(_11045_));
 sg13g2_o21ai_1 _20127_ (.B1(_11045_),
    .Y(_11046_),
    .A1(_10623_),
    .A2(_11043_));
 sg13g2_nor3_1 _20128_ (.A(net866),
    .B(net520),
    .C(_11010_),
    .Y(_11047_));
 sg13g2_buf_1 _20129_ (.A(net494),
    .X(_11048_));
 sg13g2_o21ai_1 _20130_ (.B1(_10620_),
    .Y(_11049_),
    .A1(net508),
    .A2(_10364_));
 sg13g2_nor3_1 _20131_ (.A(_11035_),
    .B(_10616_),
    .C(_10364_),
    .Y(_11050_));
 sg13g2_a21oi_1 _20132_ (.A1(_11048_),
    .A2(_11049_),
    .Y(_11051_),
    .B1(_11050_));
 sg13g2_nand2b_1 _20133_ (.Y(_11052_),
    .B(_11051_),
    .A_N(_11047_));
 sg13g2_a22oi_1 _20134_ (.Y(_11053_),
    .B1(_11052_),
    .B2(net496),
    .A2(_11046_),
    .A1(net251));
 sg13g2_a221oi_1 _20135_ (.B2(_11053_),
    .C1(_11028_),
    .B1(_11042_),
    .A1(net855),
    .Y(_11054_),
    .A2(_11031_));
 sg13g2_a221oi_1 _20136_ (.B2(_11054_),
    .C1(net100),
    .B1(_11032_),
    .A1(_11016_),
    .Y(_11055_),
    .A2(_11030_));
 sg13g2_buf_1 _20137_ (.A(\grid.cell_24_0.s ),
    .X(_11056_));
 sg13g2_buf_1 _20138_ (.A(_11056_),
    .X(_11057_));
 sg13g2_xor2_1 _20139_ (.B(_11057_),
    .A(net1112),
    .X(_11058_));
 sg13g2_xor2_1 _20140_ (.B(_11058_),
    .A(_11027_),
    .X(_11059_));
 sg13g2_buf_1 _20141_ (.A(net1107),
    .X(_11060_));
 sg13g2_a21oi_1 _20142_ (.A1(net109),
    .A2(_11059_),
    .Y(_11061_),
    .B1(_11060_));
 sg13g2_or3_1 _20143_ (.A(_10996_),
    .B(_11055_),
    .C(_11061_),
    .X(_11062_));
 sg13g2_a21oi_1 _20144_ (.A1(_10997_),
    .A2(_11062_),
    .Y(_00405_),
    .B1(net523));
 sg13g2_nand2b_1 _20145_ (.Y(_11063_),
    .B(net327),
    .A_N(_10994_));
 sg13g2_buf_1 _20146_ (.A(_11063_),
    .X(_11064_));
 sg13g2_buf_1 _20147_ (.A(\grid.cell_24_1.se ),
    .X(_11065_));
 sg13g2_buf_1 _20148_ (.A(_11065_),
    .X(_11066_));
 sg13g2_buf_1 _20149_ (.A(net844),
    .X(_11067_));
 sg13g2_buf_1 _20150_ (.A(net493),
    .X(_11068_));
 sg13g2_nor2_1 _20151_ (.A(net238),
    .B(_10383_),
    .Y(_11069_));
 sg13g2_nor2b_1 _20152_ (.A(_10364_),
    .B_N(net844),
    .Y(_11070_));
 sg13g2_nand2_1 _20153_ (.Y(_11071_),
    .A(net866),
    .B(net865));
 sg13g2_nor2_1 _20154_ (.A(net493),
    .B(_11071_),
    .Y(_11072_));
 sg13g2_o21ai_1 _20155_ (.B1(net505),
    .Y(_11073_),
    .A1(_11070_),
    .A2(_11072_));
 sg13g2_nor2_1 _20156_ (.A(net854),
    .B(_11071_),
    .Y(_11074_));
 sg13g2_o21ai_1 _20157_ (.B1(_11074_),
    .Y(_11075_),
    .A1(net493),
    .A2(net863));
 sg13g2_nand3_1 _20158_ (.B(_11073_),
    .C(_11075_),
    .A(net848),
    .Y(_11076_));
 sg13g2_nand2b_1 _20159_ (.Y(_11077_),
    .B(_10364_),
    .A_N(net844));
 sg13g2_o21ai_1 _20160_ (.B1(_11077_),
    .Y(_11078_),
    .A1(_10686_),
    .A2(_11070_));
 sg13g2_nand2_1 _20161_ (.Y(_11079_),
    .A(_11066_),
    .B(_10364_));
 sg13g2_o21ai_1 _20162_ (.B1(_10686_),
    .Y(_11080_),
    .A1(_11066_),
    .A2(_10364_));
 sg13g2_a21oi_1 _20163_ (.A1(_11079_),
    .A2(_11080_),
    .Y(_11081_),
    .B1(_11071_));
 sg13g2_a21oi_1 _20164_ (.A1(net517),
    .A2(_11078_),
    .Y(_11082_),
    .B1(_11081_));
 sg13g2_nand2_1 _20165_ (.Y(_11083_),
    .A(_11013_),
    .B(_11082_));
 sg13g2_inv_1 _20166_ (.Y(_11084_),
    .A(net844));
 sg13g2_buf_1 _20167_ (.A(_11084_),
    .X(_11085_));
 sg13g2_nand3_1 _20168_ (.B(_10705_),
    .C(net237),
    .A(_11012_),
    .Y(_11086_));
 sg13g2_nand4_1 _20169_ (.B(net518),
    .C(net854),
    .A(_10998_),
    .Y(_11087_),
    .D(_11067_));
 sg13g2_a21oi_1 _20170_ (.A1(_11086_),
    .A2(_11087_),
    .Y(_11088_),
    .B1(net251));
 sg13g2_a221oi_1 _20171_ (.B2(_11083_),
    .C1(_11088_),
    .B1(_11076_),
    .A1(_10695_),
    .Y(_11089_),
    .A2(_11069_));
 sg13g2_nor2_1 _20172_ (.A(net1112),
    .B(_11031_),
    .Y(_11090_));
 sg13g2_xnor2_1 _20173_ (.Y(_11091_),
    .A(_11084_),
    .B(_10688_));
 sg13g2_xnor2_1 _20174_ (.Y(_11092_),
    .A(_11021_),
    .B(_11091_));
 sg13g2_xnor2_1 _20175_ (.Y(_11093_),
    .A(net1107),
    .B(_11092_));
 sg13g2_nor2_1 _20176_ (.A(_10253_),
    .B(_11017_),
    .Y(_11094_));
 sg13g2_a21oi_1 _20177_ (.A1(net856),
    .A2(_11092_),
    .Y(_11095_),
    .B1(_11094_));
 sg13g2_o21ai_1 _20178_ (.B1(_11095_),
    .Y(_11096_),
    .A1(_11090_),
    .A2(_11093_));
 sg13g2_xnor2_1 _20179_ (.Y(_11097_),
    .A(_11089_),
    .B(_11096_));
 sg13g2_xnor2_1 _20180_ (.Y(_11098_),
    .A(_11058_),
    .B(_11093_));
 sg13g2_nor2_1 _20181_ (.A(net242),
    .B(_11098_),
    .Y(_11099_));
 sg13g2_buf_1 _20182_ (.A(net493),
    .X(_11100_));
 sg13g2_xnor2_1 _20183_ (.Y(_11101_),
    .A(net505),
    .B(net236));
 sg13g2_a21oi_1 _20184_ (.A1(net505),
    .A2(net236),
    .Y(_11102_),
    .B1(net521));
 sg13g2_a21oi_1 _20185_ (.A1(net251),
    .A2(_11101_),
    .Y(_11103_),
    .B1(_11102_));
 sg13g2_a22oi_1 _20186_ (.Y(_11104_),
    .B1(_11103_),
    .B2(net249),
    .A2(_11070_),
    .A1(_10767_));
 sg13g2_xor2_1 _20187_ (.B(net1107),
    .A(net1112),
    .X(_11105_));
 sg13g2_nor3_1 _20188_ (.A(net1108),
    .B(_11017_),
    .C(_11105_),
    .Y(_11106_));
 sg13g2_nand4_1 _20189_ (.B(net249),
    .C(net505),
    .A(net521),
    .Y(_11107_),
    .D(net236));
 sg13g2_o21ai_1 _20190_ (.B1(net172),
    .Y(_11108_),
    .A1(_10999_),
    .A2(_11107_));
 sg13g2_a21oi_1 _20191_ (.A1(_11092_),
    .A2(_11106_),
    .Y(_11109_),
    .B1(_11108_));
 sg13g2_o21ai_1 _20192_ (.B1(_11109_),
    .Y(_11110_),
    .A1(_11013_),
    .A2(_11104_));
 sg13g2_nor3_1 _20193_ (.A(_11097_),
    .B(_11099_),
    .C(_11110_),
    .Y(_11111_));
 sg13g2_a21oi_1 _20194_ (.A1(net242),
    .A2(net73),
    .Y(_11112_),
    .B1(_11111_));
 sg13g2_buf_2 _20195_ (.A(_03153_),
    .X(_11113_));
 sg13g2_o21ai_1 _20196_ (.B1(net522),
    .Y(_11114_),
    .A1(net38),
    .A2(_11064_));
 sg13g2_a21oi_1 _20197_ (.A1(_11064_),
    .A2(_11112_),
    .Y(_00406_),
    .B1(_11114_));
 sg13g2_nand2_1 _20198_ (.Y(_11115_),
    .A(net716),
    .B(_10996_));
 sg13g2_buf_1 _20199_ (.A(_11068_),
    .X(_11116_));
 sg13g2_buf_1 _20200_ (.A(\grid.cell_24_2.se ),
    .X(_11117_));
 sg13g2_nand2_1 _20201_ (.Y(_11118_),
    .A(net853),
    .B(net1105));
 sg13g2_xor2_1 _20202_ (.B(net1105),
    .A(_10737_),
    .X(_11119_));
 sg13g2_nand2_1 _20203_ (.Y(_11120_),
    .A(net865),
    .B(_11119_));
 sg13g2_o21ai_1 _20204_ (.B1(_11120_),
    .Y(_11121_),
    .A1(net518),
    .A2(_11118_));
 sg13g2_nand2_1 _20205_ (.Y(_11122_),
    .A(net248),
    .B(_11121_));
 sg13g2_o21ai_1 _20206_ (.B1(_11122_),
    .Y(_11123_),
    .A1(_10405_),
    .A2(_11118_));
 sg13g2_xnor2_1 _20207_ (.Y(_11124_),
    .A(_11065_),
    .B(net1105));
 sg13g2_xnor2_1 _20208_ (.Y(_11125_),
    .A(_10744_),
    .B(_11124_));
 sg13g2_xnor2_1 _20209_ (.Y(_11126_),
    .A(net865),
    .B(_11125_));
 sg13g2_and2_1 _20210_ (.A(_11019_),
    .B(_11126_),
    .X(_11127_));
 sg13g2_buf_1 _20211_ (.A(_00196_),
    .X(_11128_));
 sg13g2_buf_1 _20212_ (.A(_11128_),
    .X(_11129_));
 sg13g2_xor2_1 _20213_ (.B(net507),
    .A(net521),
    .X(_11130_));
 sg13g2_nor2_1 _20214_ (.A(_11129_),
    .B(_11130_),
    .Y(_11131_));
 sg13g2_nand2_1 _20215_ (.Y(_11132_),
    .A(net518),
    .B(net516));
 sg13g2_nor3_1 _20216_ (.A(net141),
    .B(_11118_),
    .C(_11132_),
    .Y(_11133_));
 sg13g2_a221oi_1 _20217_ (.B2(_11131_),
    .C1(_11133_),
    .B1(_11127_),
    .A1(net141),
    .Y(_11134_),
    .A2(_11123_));
 sg13g2_xnor2_1 _20218_ (.Y(_11135_),
    .A(net509),
    .B(_11126_));
 sg13g2_nand2_1 _20219_ (.Y(_11136_),
    .A(net250),
    .B(_11129_));
 sg13g2_nor2_1 _20220_ (.A(net250),
    .B(net843),
    .Y(_11137_));
 sg13g2_a221oi_1 _20221_ (.B2(_11136_),
    .C1(_11137_),
    .B1(_11135_),
    .A1(_11019_),
    .Y(_11138_),
    .A2(_11126_));
 sg13g2_buf_1 _20222_ (.A(net1105),
    .X(_11139_));
 sg13g2_nor2_1 _20223_ (.A(net504),
    .B(net842),
    .Y(_11140_));
 sg13g2_inv_1 _20224_ (.Y(_11141_),
    .A(_11118_));
 sg13g2_o21ai_1 _20225_ (.B1(_11120_),
    .Y(_11142_),
    .A1(net516),
    .A2(_11141_));
 sg13g2_a22oi_1 _20226_ (.Y(_11143_),
    .B1(_11142_),
    .B2(_10405_),
    .A2(_11140_),
    .A1(_11132_));
 sg13g2_o21ai_1 _20227_ (.B1(net248),
    .Y(_11144_),
    .A1(net517),
    .A2(net237));
 sg13g2_nand3_1 _20228_ (.B(_11144_),
    .C(_11140_),
    .A(_10405_),
    .Y(_11145_));
 sg13g2_o21ai_1 _20229_ (.B1(_11145_),
    .Y(_11146_),
    .A1(_11068_),
    .A2(_11143_));
 sg13g2_xor2_1 _20230_ (.B(_11146_),
    .A(_11138_),
    .X(_11147_));
 sg13g2_a21oi_1 _20231_ (.A1(_11134_),
    .A2(_11147_),
    .Y(_11148_),
    .B1(net117));
 sg13g2_xnor2_1 _20232_ (.Y(_11149_),
    .A(_11021_),
    .B(_11135_));
 sg13g2_a21oi_1 _20233_ (.A1(net122),
    .A2(_11149_),
    .Y(_11150_),
    .B1(_10767_));
 sg13g2_nand2_1 _20234_ (.Y(_11151_),
    .A(net1059),
    .B(_11064_));
 sg13g2_or3_1 _20235_ (.A(_11148_),
    .B(_11150_),
    .C(_11151_),
    .X(_11152_));
 sg13g2_o21ai_1 _20236_ (.B1(_11152_),
    .Y(_00407_),
    .A1(net27),
    .A2(_11115_));
 sg13g2_buf_1 _20237_ (.A(_00193_),
    .X(_11153_));
 sg13g2_buf_2 _20238_ (.A(\grid.cell_24_3.se ),
    .X(_11154_));
 sg13g2_xnor2_1 _20239_ (.Y(_11155_),
    .A(_11154_),
    .B(_11117_));
 sg13g2_xnor2_1 _20240_ (.Y(_11156_),
    .A(_10797_),
    .B(_11155_));
 sg13g2_xnor2_1 _20241_ (.Y(_11157_),
    .A(net515),
    .B(_11156_));
 sg13g2_nor4_1 _20242_ (.A(_10796_),
    .B(net1104),
    .C(_10688_),
    .D(_11157_),
    .Y(_11158_));
 sg13g2_buf_1 _20243_ (.A(_11154_),
    .X(_11159_));
 sg13g2_inv_1 _20244_ (.Y(_11160_),
    .A(net841));
 sg13g2_buf_1 _20245_ (.A(_11160_),
    .X(_11161_));
 sg13g2_inv_2 _20246_ (.Y(_11162_),
    .A(net1105));
 sg13g2_nand2_1 _20247_ (.Y(_11163_),
    .A(net235),
    .B(_11162_));
 sg13g2_a21oi_1 _20248_ (.A1(net851),
    .A2(net516),
    .Y(_11164_),
    .B1(_10454_));
 sg13g2_nor2_1 _20249_ (.A(net515),
    .B(_11155_),
    .Y(_11165_));
 sg13g2_a21oi_1 _20250_ (.A1(net841),
    .A2(_11117_),
    .Y(_11166_),
    .B1(net862));
 sg13g2_o21ai_1 _20251_ (.B1(_10806_),
    .Y(_11167_),
    .A1(_11165_),
    .A2(_11166_));
 sg13g2_o21ai_1 _20252_ (.B1(_11167_),
    .Y(_11168_),
    .A1(_11163_),
    .A2(_11164_));
 sg13g2_nor2_1 _20253_ (.A(net503),
    .B(_11163_),
    .Y(_11169_));
 sg13g2_nand2_1 _20254_ (.Y(_11170_),
    .A(net247),
    .B(net248));
 sg13g2_a22oi_1 _20255_ (.Y(_11171_),
    .B1(_11169_),
    .B2(_11170_),
    .A2(_11168_),
    .A1(net1111));
 sg13g2_nand2_1 _20256_ (.Y(_11172_),
    .A(net517),
    .B(_11153_));
 sg13g2_xnor2_1 _20257_ (.Y(_11173_),
    .A(net505),
    .B(_11157_));
 sg13g2_inv_1 _20258_ (.Y(_11174_),
    .A(net1104));
 sg13g2_nand2_1 _20259_ (.Y(_11175_),
    .A(net249),
    .B(_11174_));
 sg13g2_o21ai_1 _20260_ (.B1(_11175_),
    .Y(_11176_),
    .A1(_10796_),
    .A2(_11157_));
 sg13g2_a21oi_1 _20261_ (.A1(_11172_),
    .A2(_11173_),
    .Y(_11177_),
    .B1(_11176_));
 sg13g2_xor2_1 _20262_ (.B(_11177_),
    .A(_11171_),
    .X(_11178_));
 sg13g2_buf_1 _20263_ (.A(net841),
    .X(_11179_));
 sg13g2_buf_1 _20264_ (.A(net842),
    .X(_11180_));
 sg13g2_nand2_1 _20265_ (.Y(_11181_),
    .A(net492),
    .B(net491));
 sg13g2_or2_1 _20266_ (.X(_11182_),
    .B(_11181_),
    .A(net1111));
 sg13g2_xor2_1 _20267_ (.B(net516),
    .A(net841),
    .X(_11183_));
 sg13g2_nor2_1 _20268_ (.A(net515),
    .B(_11139_),
    .Y(_11184_));
 sg13g2_a22oi_1 _20269_ (.Y(_11185_),
    .B1(_11184_),
    .B2(net492),
    .A2(_11183_),
    .A1(net491));
 sg13g2_nand2b_1 _20270_ (.Y(_11186_),
    .B(net247),
    .A_N(_11185_));
 sg13g2_a21oi_1 _20271_ (.A1(_11182_),
    .A2(_11186_),
    .Y(_11187_),
    .B1(net502));
 sg13g2_nand4_1 _20272_ (.B(net492),
    .C(net248),
    .A(net247),
    .Y(_11188_),
    .D(_11180_));
 sg13g2_o21ai_1 _20273_ (.B1(net1054),
    .Y(_11189_),
    .A1(net503),
    .A2(_11188_));
 sg13g2_nor4_1 _20274_ (.A(_11158_),
    .B(_11178_),
    .C(_11187_),
    .D(_11189_),
    .Y(_11190_));
 sg13g2_xnor2_1 _20275_ (.Y(_11191_),
    .A(_11091_),
    .B(_11157_));
 sg13g2_a21oi_1 _20276_ (.A1(net114),
    .A2(_11191_),
    .Y(_11192_),
    .B1(net504));
 sg13g2_nor2_1 _20277_ (.A(_10996_),
    .B(_11192_),
    .Y(_11193_));
 sg13g2_o21ai_1 _20278_ (.B1(_11193_),
    .Y(_11194_),
    .A1(_08877_),
    .A2(_11190_));
 sg13g2_o21ai_1 _20279_ (.B1(_11194_),
    .Y(_00408_),
    .A1(net26),
    .A2(_11064_));
 sg13g2_buf_1 _20280_ (.A(\grid.cell_24_4.se ),
    .X(_11195_));
 sg13g2_buf_1 _20281_ (.A(net1103),
    .X(_11196_));
 sg13g2_nand2_1 _20282_ (.Y(_11197_),
    .A(net840),
    .B(_11159_));
 sg13g2_nand2_1 _20283_ (.Y(_11198_),
    .A(net862),
    .B(_11159_));
 sg13g2_xor2_1 _20284_ (.B(_11154_),
    .A(_10398_),
    .X(_11199_));
 sg13g2_nand2_1 _20285_ (.Y(_11200_),
    .A(net840),
    .B(_11199_));
 sg13g2_o21ai_1 _20286_ (.B1(_11200_),
    .Y(_11201_),
    .A1(_11196_),
    .A2(_11198_));
 sg13g2_nand2_1 _20287_ (.Y(_11202_),
    .A(net246),
    .B(_11201_));
 sg13g2_o21ai_1 _20288_ (.B1(_11202_),
    .Y(_11203_),
    .A1(_10467_),
    .A2(_11197_));
 sg13g2_xnor2_1 _20289_ (.Y(_11204_),
    .A(net1103),
    .B(_10821_));
 sg13g2_xor2_1 _20290_ (.B(_11204_),
    .A(_11199_),
    .X(_11205_));
 sg13g2_and2_1 _20291_ (.A(_10853_),
    .B(_11205_),
    .X(_11206_));
 sg13g2_buf_2 _20292_ (.A(_00057_),
    .X(_11207_));
 sg13g2_nor2b_1 _20293_ (.A(_11207_),
    .B_N(_10744_),
    .Y(_11208_));
 sg13g2_inv_1 _20294_ (.Y(_11209_),
    .A(net1103));
 sg13g2_buf_1 _20295_ (.A(_11209_),
    .X(_11210_));
 sg13g2_nor4_1 _20296_ (.A(net501),
    .B(_10833_),
    .C(net490),
    .D(_11198_),
    .Y(_11211_));
 sg13g2_a221oi_1 _20297_ (.B2(_11208_),
    .C1(_11211_),
    .B1(_11206_),
    .A1(net501),
    .Y(_11212_),
    .A2(_11203_));
 sg13g2_xor2_1 _20298_ (.B(_11154_),
    .A(net1103),
    .X(_11213_));
 sg13g2_a22oi_1 _20299_ (.Y(_11214_),
    .B1(_11213_),
    .B2(net514),
    .A2(_11197_),
    .A1(_10833_));
 sg13g2_o21ai_1 _20300_ (.B1(net861),
    .Y(_11215_),
    .A1(_10840_),
    .A2(_10454_));
 sg13g2_nand3_1 _20301_ (.B(net235),
    .C(_11215_),
    .A(net490),
    .Y(_11216_));
 sg13g2_o21ai_1 _20302_ (.B1(_11216_),
    .Y(_11217_),
    .A1(net850),
    .A2(_11214_));
 sg13g2_buf_1 _20303_ (.A(net840),
    .X(_11218_));
 sg13g2_nor3_1 _20304_ (.A(net501),
    .B(_11218_),
    .C(_11179_),
    .Y(_11219_));
 sg13g2_nand2_1 _20305_ (.Y(_11220_),
    .A(net246),
    .B(net247));
 sg13g2_a22oi_1 _20306_ (.Y(_11221_),
    .B1(_11219_),
    .B2(_11220_),
    .A2(_11217_),
    .A1(_10467_));
 sg13g2_nand2_1 _20307_ (.Y(_11222_),
    .A(_11207_),
    .B(net515));
 sg13g2_xnor2_1 _20308_ (.Y(_11223_),
    .A(_10739_),
    .B(_11205_));
 sg13g2_nor2_1 _20309_ (.A(_11207_),
    .B(net515),
    .Y(_11224_));
 sg13g2_a221oi_1 _20310_ (.B2(_11223_),
    .C1(_11224_),
    .B1(_11222_),
    .A1(_10853_),
    .Y(_11225_),
    .A2(_11205_));
 sg13g2_xnor2_1 _20311_ (.Y(_11226_),
    .A(_11221_),
    .B(_11225_));
 sg13g2_a21oi_1 _20312_ (.A1(_11212_),
    .A2(_11226_),
    .Y(_11227_),
    .B1(net101));
 sg13g2_xnor2_1 _20313_ (.Y(_11228_),
    .A(_11162_),
    .B(_10744_));
 sg13g2_xnor2_1 _20314_ (.Y(_11229_),
    .A(_11205_),
    .B(_11228_));
 sg13g2_a21oi_1 _20315_ (.A1(_09402_),
    .A2(_11229_),
    .Y(_11230_),
    .B1(_10785_));
 sg13g2_or3_1 _20316_ (.A(_11151_),
    .B(_11227_),
    .C(_11230_),
    .X(_11231_));
 sg13g2_o21ai_1 _20317_ (.B1(_11231_),
    .Y(_00409_),
    .A1(net34),
    .A2(_11115_));
 sg13g2_buf_1 _20318_ (.A(_00089_),
    .X(_11232_));
 sg13g2_inv_1 _20319_ (.Y(_11233_),
    .A(_11232_));
 sg13g2_nor2_1 _20320_ (.A(_11233_),
    .B(net514),
    .Y(_11234_));
 sg13g2_buf_8 _20321_ (.A(\grid.cell_24_5.se ),
    .X(_11235_));
 sg13g2_xnor2_1 _20322_ (.Y(_11236_),
    .A(_11235_),
    .B(_10870_));
 sg13g2_xnor2_1 _20323_ (.Y(_11237_),
    .A(_10470_),
    .B(_11236_));
 sg13g2_xnor2_1 _20324_ (.Y(_11238_),
    .A(net1103),
    .B(_11237_));
 sg13g2_xnor2_1 _20325_ (.Y(_11239_),
    .A(net851),
    .B(_11238_));
 sg13g2_a22oi_1 _20326_ (.Y(_11240_),
    .B1(_11238_),
    .B2(_10898_),
    .A2(net514),
    .A1(_11233_));
 sg13g2_o21ai_1 _20327_ (.B1(_11240_),
    .Y(_11241_),
    .A1(_11234_),
    .A2(_11239_));
 sg13g2_buf_1 _20328_ (.A(_11235_),
    .X(_11242_));
 sg13g2_buf_1 _20329_ (.A(net839),
    .X(_11243_));
 sg13g2_xor2_1 _20330_ (.B(_10875_),
    .A(net1103),
    .X(_11244_));
 sg13g2_nand2_1 _20331_ (.Y(_11245_),
    .A(_11196_),
    .B(_10875_));
 sg13g2_a22oi_1 _20332_ (.Y(_11246_),
    .B1(_11245_),
    .B2(net512),
    .A2(_11244_),
    .A1(net861));
 sg13g2_inv_2 _20333_ (.Y(_11247_),
    .A(_11235_));
 sg13g2_o21ai_1 _20334_ (.B1(net860),
    .Y(_11248_),
    .A1(_11247_),
    .A2(_10833_));
 sg13g2_nand3_1 _20335_ (.B(_10872_),
    .C(_11248_),
    .A(net490),
    .Y(_11249_));
 sg13g2_o21ai_1 _20336_ (.B1(_11249_),
    .Y(_11250_),
    .A1(net488),
    .A2(_11246_));
 sg13g2_nor3_1 _20337_ (.A(net488),
    .B(_11218_),
    .C(net498),
    .Y(_11251_));
 sg13g2_nand2_1 _20338_ (.Y(_11252_),
    .A(net510),
    .B(net513));
 sg13g2_a22oi_1 _20339_ (.Y(_11253_),
    .B1(_11251_),
    .B2(_11252_),
    .A2(_11250_),
    .A1(net1110));
 sg13g2_xor2_1 _20340_ (.B(_11253_),
    .A(_11241_),
    .X(_11254_));
 sg13g2_buf_1 _20341_ (.A(net488),
    .X(_11255_));
 sg13g2_nand2_1 _20342_ (.Y(_11256_),
    .A(net861),
    .B(_11244_));
 sg13g2_o21ai_1 _20343_ (.B1(_11256_),
    .Y(_11257_),
    .A1(net513),
    .A2(_11245_));
 sg13g2_nand2_1 _20344_ (.Y(_11258_),
    .A(net511),
    .B(_11257_));
 sg13g2_o21ai_1 _20345_ (.B1(_11258_),
    .Y(_11259_),
    .A1(net1110),
    .A2(_11245_));
 sg13g2_and2_1 _20346_ (.A(_11233_),
    .B(_10797_),
    .X(_11260_));
 sg13g2_and2_1 _20347_ (.A(_10898_),
    .B(_11238_),
    .X(_11261_));
 sg13g2_nor3_1 _20348_ (.A(net234),
    .B(_11252_),
    .C(_11245_),
    .Y(_11262_));
 sg13g2_a221oi_1 _20349_ (.B2(_11261_),
    .C1(_11262_),
    .B1(_11260_),
    .A1(net234),
    .Y(_11263_),
    .A2(_11259_));
 sg13g2_a21oi_1 _20350_ (.A1(_11254_),
    .A2(_11263_),
    .Y(_11264_),
    .B1(net101));
 sg13g2_xnor2_1 _20351_ (.Y(_11265_),
    .A(net235),
    .B(_10797_));
 sg13g2_xnor2_1 _20352_ (.Y(_11266_),
    .A(_11238_),
    .B(_11265_));
 sg13g2_a21oi_1 _20353_ (.A1(net68),
    .A2(_11266_),
    .Y(_11267_),
    .B1(net501));
 sg13g2_or3_1 _20354_ (.A(_11151_),
    .B(_11264_),
    .C(_11267_),
    .X(_11268_));
 sg13g2_o21ai_1 _20355_ (.B1(_11268_),
    .Y(_00410_),
    .A1(net46),
    .A2(_11115_));
 sg13g2_nand2_1 _20356_ (.Y(_11269_),
    .A(_10658_),
    .B(net860));
 sg13g2_nand2_1 _20357_ (.Y(_11270_),
    .A(net239),
    .B(_10975_));
 sg13g2_o21ai_1 _20358_ (.B1(_11270_),
    .Y(_11271_),
    .A1(_11048_),
    .A2(_11269_));
 sg13g2_buf_2 _20359_ (.A(_00150_),
    .X(_11272_));
 sg13g2_nand2_1 _20360_ (.Y(_11273_),
    .A(net847),
    .B(net858));
 sg13g2_nor2_1 _20361_ (.A(_11272_),
    .B(_11273_),
    .Y(_11274_));
 sg13g2_a21oi_1 _20362_ (.A1(net243),
    .A2(_11271_),
    .Y(_11275_),
    .B1(_11274_));
 sg13g2_nand2_1 _20363_ (.Y(_11276_),
    .A(net860),
    .B(net867));
 sg13g2_nor3_1 _20364_ (.A(_11243_),
    .B(_11276_),
    .C(_11273_),
    .Y(_11277_));
 sg13g2_nor2_1 _20365_ (.A(net368),
    .B(_11277_),
    .Y(_11278_));
 sg13g2_o21ai_1 _20366_ (.B1(_11278_),
    .Y(_11279_),
    .A1(_11247_),
    .A2(_11275_));
 sg13g2_buf_2 _20367_ (.A(_00121_),
    .X(_11280_));
 sg13g2_inv_1 _20368_ (.Y(_11281_),
    .A(_10821_));
 sg13g2_xnor2_1 _20369_ (.Y(_11282_),
    .A(_11235_),
    .B(_11001_));
 sg13g2_xor2_1 _20370_ (.B(_11282_),
    .A(_10975_),
    .X(_11283_));
 sg13g2_xnor2_1 _20371_ (.Y(_11284_),
    .A(net520),
    .B(_11283_));
 sg13g2_nor4_1 _20372_ (.A(_10944_),
    .B(_11280_),
    .C(_11281_),
    .D(_11284_),
    .Y(_11285_));
 sg13g2_nand2_1 _20373_ (.Y(_11286_),
    .A(_11280_),
    .B(_10833_));
 sg13g2_xnor2_1 _20374_ (.Y(_11287_),
    .A(net850),
    .B(_11284_));
 sg13g2_nand2b_1 _20375_ (.Y(_11288_),
    .B(net513),
    .A_N(_11280_));
 sg13g2_o21ai_1 _20376_ (.B1(_11288_),
    .Y(_11289_),
    .A1(_10944_),
    .A2(_11284_));
 sg13g2_a21oi_1 _20377_ (.A1(_11286_),
    .A2(_11287_),
    .Y(_11290_),
    .B1(_11289_));
 sg13g2_nand2_1 _20378_ (.Y(_11291_),
    .A(net847),
    .B(net867));
 sg13g2_a21oi_1 _20379_ (.A1(_11034_),
    .A2(_11291_),
    .Y(_11292_),
    .B1(net839));
 sg13g2_nor3_1 _20380_ (.A(_11272_),
    .B(_11038_),
    .C(_10632_),
    .Y(_11293_));
 sg13g2_a21oi_1 _20381_ (.A1(_11272_),
    .A2(_11292_),
    .Y(_11294_),
    .B1(_11293_));
 sg13g2_nor2_1 _20382_ (.A(net512),
    .B(_11294_),
    .Y(_11295_));
 sg13g2_nand2_1 _20383_ (.Y(_11296_),
    .A(_11247_),
    .B(_11010_));
 sg13g2_nand2_1 _20384_ (.Y(_11297_),
    .A(_11235_),
    .B(net847));
 sg13g2_or2_1 _20385_ (.X(_11298_),
    .B(_11297_),
    .A(_10632_));
 sg13g2_a21oi_1 _20386_ (.A1(_11296_),
    .A2(_11298_),
    .Y(_11299_),
    .B1(net510));
 sg13g2_nor3_1 _20387_ (.A(_11272_),
    .B(net847),
    .C(net858),
    .Y(_11300_));
 sg13g2_nor3_1 _20388_ (.A(_11276_),
    .B(_11004_),
    .C(_11300_),
    .Y(_11301_));
 sg13g2_nor2_1 _20389_ (.A(_11274_),
    .B(_11301_),
    .Y(_11302_));
 sg13g2_nor2_1 _20390_ (.A(_11247_),
    .B(_11302_),
    .Y(_11303_));
 sg13g2_nor2_1 _20391_ (.A(net839),
    .B(_11004_),
    .Y(_11304_));
 sg13g2_o21ai_1 _20392_ (.B1(_11272_),
    .Y(_11305_),
    .A1(_11010_),
    .A2(_11304_));
 sg13g2_a21oi_1 _20393_ (.A1(_11296_),
    .A2(_11305_),
    .Y(_11306_),
    .B1(net243));
 sg13g2_nor4_1 _20394_ (.A(_11295_),
    .B(_11299_),
    .C(_11303_),
    .D(_11306_),
    .Y(_11307_));
 sg13g2_xor2_1 _20395_ (.B(_11307_),
    .A(_11290_),
    .X(_11308_));
 sg13g2_nor3_1 _20396_ (.A(_11279_),
    .B(_11285_),
    .C(_11308_),
    .Y(_11309_));
 sg13g2_nor2_1 _20397_ (.A(net499),
    .B(_10996_),
    .Y(_11310_));
 sg13g2_o21ai_1 _20398_ (.B1(_11310_),
    .Y(_11311_),
    .A1(net75),
    .A2(_11309_));
 sg13g2_xor2_1 _20399_ (.B(_11284_),
    .A(_11204_),
    .X(_11312_));
 sg13g2_nor2_1 _20400_ (.A(_10996_),
    .B(_11312_),
    .Y(_11313_));
 sg13g2_a22oi_1 _20401_ (.Y(_11314_),
    .B1(_11309_),
    .B2(_11313_),
    .A2(_10996_),
    .A1(net45));
 sg13g2_a21oi_1 _20402_ (.A1(_11311_),
    .A2(_11314_),
    .Y(_00411_),
    .B1(net523));
 sg13g2_xnor2_1 _20403_ (.Y(_11315_),
    .A(_10870_),
    .B(_11282_));
 sg13g2_o21ai_1 _20404_ (.B1(_11272_),
    .Y(_11316_),
    .A1(net860),
    .A2(net520));
 sg13g2_nand2_1 _20405_ (.Y(_11317_),
    .A(_11315_),
    .B(_11316_));
 sg13g2_o21ai_1 _20406_ (.B1(_11317_),
    .Y(_11318_),
    .A1(_11276_),
    .A2(_11315_));
 sg13g2_xnor2_1 _20407_ (.Y(_11319_),
    .A(_10521_),
    .B(_11315_));
 sg13g2_buf_2 _20408_ (.A(_11319_),
    .X(_11320_));
 sg13g2_a21oi_1 _20409_ (.A1(_11035_),
    .A2(net498),
    .Y(_11321_),
    .B1(net839));
 sg13g2_a21oi_2 _20410_ (.B1(_11321_),
    .Y(_11322_),
    .A2(net499),
    .A1(_11038_));
 sg13g2_nor4_1 _20411_ (.A(net855),
    .B(net845),
    .C(_11017_),
    .D(_11322_),
    .Y(_11323_));
 sg13g2_a21oi_1 _20412_ (.A1(_11320_),
    .A2(_11322_),
    .Y(_11324_),
    .B1(_11323_));
 sg13g2_nand3_1 _20413_ (.B(_11094_),
    .C(_11320_),
    .A(net845),
    .Y(_11325_));
 sg13g2_a21oi_1 _20414_ (.A1(_11324_),
    .A2(_11325_),
    .Y(_11326_),
    .B1(net1108));
 sg13g2_nand2_1 _20415_ (.Y(_11327_),
    .A(net856),
    .B(_11320_));
 sg13g2_nand3_1 _20416_ (.B(net1108),
    .C(_11320_),
    .A(net845),
    .Y(_11328_));
 sg13g2_or2_1 _20417_ (.X(_11329_),
    .B(_11320_),
    .A(net1107));
 sg13g2_a21oi_1 _20418_ (.A1(_11328_),
    .A2(_11329_),
    .Y(_11330_),
    .B1(_11094_));
 sg13g2_a21oi_1 _20419_ (.A1(_11090_),
    .A2(_11327_),
    .Y(_11331_),
    .B1(_11330_));
 sg13g2_xnor2_1 _20420_ (.Y(_11332_),
    .A(_10651_),
    .B(_11320_));
 sg13g2_inv_1 _20421_ (.Y(_11333_),
    .A(_11094_));
 sg13g2_o21ai_1 _20422_ (.B1(_11333_),
    .Y(_11334_),
    .A1(_11090_),
    .A2(_11332_));
 sg13g2_nand2_1 _20423_ (.Y(_11335_),
    .A(_11322_),
    .B(_11334_));
 sg13g2_o21ai_1 _20424_ (.B1(_11335_),
    .Y(_11336_),
    .A1(_11322_),
    .A2(_11331_));
 sg13g2_or3_1 _20425_ (.A(_11318_),
    .B(_11326_),
    .C(_11336_),
    .X(_11337_));
 sg13g2_nand2_1 _20426_ (.Y(_11338_),
    .A(_11318_),
    .B(_11327_));
 sg13g2_nor3_1 _20427_ (.A(_11322_),
    .B(_11334_),
    .C(_11338_),
    .Y(_11339_));
 sg13g2_nand2_1 _20428_ (.Y(_11340_),
    .A(net158),
    .B(_05677_));
 sg13g2_nor2_1 _20429_ (.A(_11340_),
    .B(_10994_),
    .Y(_11341_));
 sg13g2_nor3_1 _20430_ (.A(net103),
    .B(_11339_),
    .C(_11341_),
    .Y(_11342_));
 sg13g2_xnor2_1 _20431_ (.Y(_11343_),
    .A(_11058_),
    .B(_11332_));
 sg13g2_nand2_1 _20432_ (.Y(_11344_),
    .A(net78),
    .B(_11343_));
 sg13g2_nor2_1 _20433_ (.A(_10658_),
    .B(_11341_),
    .Y(_11345_));
 sg13g2_nand2_1 _20434_ (.Y(_11346_),
    .A(net327),
    .B(_05128_));
 sg13g2_buf_2 _20435_ (.A(_11346_),
    .X(_11347_));
 sg13g2_o21ai_1 _20436_ (.B1(net668),
    .Y(_11348_),
    .A1(_11347_),
    .A2(_10994_));
 sg13g2_a221oi_1 _20437_ (.B2(_11345_),
    .C1(_11348_),
    .B1(_11344_),
    .A1(_11337_),
    .Y(_00412_),
    .A2(_11342_));
 sg13g2_inv_1 _20438_ (.Y(_11349_),
    .A(_11128_));
 sg13g2_buf_1 _20439_ (.A(\grid.cell_25_0.sw ),
    .X(_11350_));
 sg13g2_buf_1 _20440_ (.A(net1102),
    .X(_11351_));
 sg13g2_buf_2 _20441_ (.A(\grid.cell_25_0.se ),
    .X(_11352_));
 sg13g2_xnor2_1 _20442_ (.Y(_11353_),
    .A(_10607_),
    .B(_11352_));
 sg13g2_xor2_1 _20443_ (.B(_11353_),
    .A(_11005_),
    .X(_11354_));
 sg13g2_xnor2_1 _20444_ (.Y(_11355_),
    .A(net837),
    .B(_11354_));
 sg13g2_xnor2_1 _20445_ (.Y(_11356_),
    .A(_11012_),
    .B(_11355_));
 sg13g2_a22oi_1 _20446_ (.Y(_11357_),
    .B1(_11356_),
    .B2(net845),
    .A2(_11355_),
    .A1(net838));
 sg13g2_or2_1 _20447_ (.X(_11358_),
    .B(net837),
    .A(_11002_));
 sg13g2_buf_1 _20448_ (.A(_11358_),
    .X(_11359_));
 sg13g2_buf_1 _20449_ (.A(_11352_),
    .X(_11360_));
 sg13g2_nand2b_1 _20450_ (.Y(_11361_),
    .B(net241),
    .A_N(net836));
 sg13g2_buf_1 _20451_ (.A(_11352_),
    .X(_11362_));
 sg13g2_buf_1 _20452_ (.A(net837),
    .X(_11363_));
 sg13g2_buf_1 _20453_ (.A(net487),
    .X(_11364_));
 sg13g2_nand4_1 _20454_ (.B(net239),
    .C(net852),
    .A(net835),
    .Y(_11365_),
    .D(net233));
 sg13g2_o21ai_1 _20455_ (.B1(_11365_),
    .Y(_11366_),
    .A1(_11359_),
    .A2(_11361_));
 sg13g2_buf_1 _20456_ (.A(net239),
    .X(_11367_));
 sg13g2_nand2_1 _20457_ (.Y(_11368_),
    .A(_11018_),
    .B(net487));
 sg13g2_nor2b_1 _20458_ (.A(net239),
    .B_N(net487),
    .Y(_11369_));
 sg13g2_a21oi_1 _20459_ (.A1(net140),
    .A2(_11368_),
    .Y(_11370_),
    .B1(_11369_));
 sg13g2_nor2_1 _20460_ (.A(net494),
    .B(net837),
    .Y(_11371_));
 sg13g2_o21ai_1 _20461_ (.B1(_11034_),
    .Y(_11372_),
    .A1(_11038_),
    .A2(net487));
 sg13g2_a22oi_1 _20462_ (.Y(_11373_),
    .B1(_11372_),
    .B2(net509),
    .A2(_11371_),
    .A1(net495));
 sg13g2_o21ai_1 _20463_ (.B1(_11373_),
    .Y(_11374_),
    .A1(net241),
    .A2(_11370_));
 sg13g2_buf_1 _20464_ (.A(net836),
    .X(_11375_));
 sg13g2_nor2b_1 _20465_ (.A(net857),
    .B_N(net508),
    .Y(_11376_));
 sg13g2_mux2_1 _20466_ (.A0(net495),
    .A1(_10616_),
    .S(net487),
    .X(_11377_));
 sg13g2_nor2_1 _20467_ (.A(net239),
    .B(_11368_),
    .Y(_11378_));
 sg13g2_a221oi_1 _20468_ (.B2(net140),
    .C1(_11378_),
    .B1(_11377_),
    .A1(_11359_),
    .Y(_11379_),
    .A2(_11376_));
 sg13g2_nor2_1 _20469_ (.A(net486),
    .B(_11379_),
    .Y(_11380_));
 sg13g2_a221oi_1 _20470_ (.B2(net486),
    .C1(_11380_),
    .B1(_11374_),
    .A1(net242),
    .Y(_11381_),
    .A2(_11366_));
 sg13g2_xor2_1 _20471_ (.B(_11356_),
    .A(net845),
    .X(_11382_));
 sg13g2_buf_2 _20472_ (.A(_00016_),
    .X(_11383_));
 sg13g2_inv_1 _20473_ (.Y(_11384_),
    .A(_11383_));
 sg13g2_a21o_1 _20474_ (.A2(net835),
    .A1(net507),
    .B1(net506),
    .X(_11385_));
 sg13g2_nor2_1 _20475_ (.A(net495),
    .B(_11359_),
    .Y(_11386_));
 sg13g2_or2_1 _20476_ (.X(_11387_),
    .B(_11034_),
    .A(net837));
 sg13g2_a21oi_1 _20477_ (.A1(net494),
    .A2(net487),
    .Y(_11388_),
    .B1(_11376_));
 sg13g2_nand3_1 _20478_ (.B(_11387_),
    .C(_11388_),
    .A(net852),
    .Y(_11389_));
 sg13g2_o21ai_1 _20479_ (.B1(_11371_),
    .Y(_11390_),
    .A1(net509),
    .A2(net506));
 sg13g2_a21oi_1 _20480_ (.A1(_11389_),
    .A2(_11390_),
    .Y(_11391_),
    .B1(net835));
 sg13g2_a21oi_1 _20481_ (.A1(_11385_),
    .A2(_11386_),
    .Y(_11392_),
    .B1(_11391_));
 sg13g2_nor2b_1 _20482_ (.A(_11357_),
    .B_N(_11392_),
    .Y(_11393_));
 sg13g2_a221oi_1 _20483_ (.B2(_11384_),
    .C1(_11393_),
    .B1(_11382_),
    .A1(_11357_),
    .Y(_11394_),
    .A2(_11381_));
 sg13g2_nand2_1 _20484_ (.Y(_11395_),
    .A(_11384_),
    .B(_11382_));
 sg13g2_nand2b_1 _20485_ (.Y(_11396_),
    .B(_11357_),
    .A_N(_11392_));
 sg13g2_o21ai_1 _20486_ (.B1(net85),
    .Y(_11397_),
    .A1(_11395_),
    .A2(_11396_));
 sg13g2_nor2_1 _20487_ (.A(_11394_),
    .B(_11397_),
    .Y(_11398_));
 sg13g2_buf_2 _20488_ (.A(\grid.cell_25_0.s ),
    .X(_11399_));
 sg13g2_inv_2 _20489_ (.Y(_11400_),
    .A(_11399_));
 sg13g2_xnor2_1 _20490_ (.Y(_11401_),
    .A(_11400_),
    .B(_11382_));
 sg13g2_a21oi_1 _20491_ (.A1(net112),
    .A2(_11401_),
    .Y(_11402_),
    .B1(net846));
 sg13g2_or4_1 _20492_ (.A(_07972_),
    .B(net320),
    .C(_02021_),
    .D(_10992_),
    .X(_11403_));
 sg13g2_buf_2 _20493_ (.A(_11403_),
    .X(_11404_));
 sg13g2_nand2_1 _20494_ (.Y(_11405_),
    .A(net1059),
    .B(_11404_));
 sg13g2_or2_1 _20495_ (.X(_11406_),
    .B(_11405_),
    .A(_11402_));
 sg13g2_buf_2 _20496_ (.A(_06472_),
    .X(_11407_));
 sg13g2_nor4_2 _20497_ (.A(_07972_),
    .B(net139),
    .C(net375),
    .Y(_11408_),
    .D(_10992_));
 sg13g2_nand2_2 _20498_ (.Y(_11409_),
    .A(net1059),
    .B(_11408_));
 sg13g2_nand2b_1 _20499_ (.Y(_11410_),
    .B(net44),
    .A_N(_11409_));
 sg13g2_o21ai_1 _20500_ (.B1(_11410_),
    .Y(_00413_),
    .A1(_11398_),
    .A2(_11406_));
 sg13g2_buf_1 _20501_ (.A(_06331_),
    .X(_11411_));
 sg13g2_buf_1 _20502_ (.A(\grid.cell_25_1.se ),
    .X(_11412_));
 sg13g2_buf_1 _20503_ (.A(_11412_),
    .X(_11413_));
 sg13g2_buf_1 _20504_ (.A(net834),
    .X(_11414_));
 sg13g2_buf_2 _20505_ (.A(_11414_),
    .X(_11415_));
 sg13g2_buf_1 _20506_ (.A(net232),
    .X(_11416_));
 sg13g2_nor4_1 _20507_ (.A(net240),
    .B(net238),
    .C(net138),
    .D(net495),
    .Y(_11417_));
 sg13g2_or3_1 _20508_ (.A(net836),
    .B(net236),
    .C(net232),
    .X(_11418_));
 sg13g2_nand4_1 _20509_ (.B(net505),
    .C(net238),
    .A(net835),
    .Y(_11419_),
    .D(net232));
 sg13g2_a21oi_1 _20510_ (.A1(_11418_),
    .A2(_11419_),
    .Y(_11420_),
    .B1(net242));
 sg13g2_nand2b_1 _20511_ (.Y(_11421_),
    .B(net834),
    .A_N(_10758_));
 sg13g2_nand2_1 _20512_ (.Y(_11422_),
    .A(_11084_),
    .B(_11421_));
 sg13g2_o21ai_1 _20513_ (.B1(_11422_),
    .Y(_11423_),
    .A1(net485),
    .A2(net495));
 sg13g2_nand2_1 _20514_ (.Y(_11424_),
    .A(net485),
    .B(net852));
 sg13g2_o21ai_1 _20515_ (.B1(_11067_),
    .Y(_11425_),
    .A1(net485),
    .A2(_10758_));
 sg13g2_nand2_1 _20516_ (.Y(_11426_),
    .A(net857),
    .B(_10685_));
 sg13g2_a21oi_1 _20517_ (.A1(_11424_),
    .A2(_11425_),
    .Y(_11427_),
    .B1(_11426_));
 sg13g2_a21oi_1 _20518_ (.A1(_10705_),
    .A2(_11423_),
    .Y(_11428_),
    .B1(_11427_));
 sg13g2_o21ai_1 _20519_ (.B1(_11421_),
    .Y(_11429_),
    .A1(net485),
    .A2(_11426_));
 sg13g2_nor2_1 _20520_ (.A(net834),
    .B(_10758_),
    .Y(_11430_));
 sg13g2_nor3_1 _20521_ (.A(net493),
    .B(_11426_),
    .C(_11430_),
    .Y(_11431_));
 sg13g2_a21oi_1 _20522_ (.A1(net236),
    .A2(_11429_),
    .Y(_11432_),
    .B1(_11431_));
 sg13g2_nand2b_1 _20523_ (.Y(_11433_),
    .B(net835),
    .A_N(_11432_));
 sg13g2_o21ai_1 _20524_ (.B1(_11433_),
    .Y(_11434_),
    .A1(net486),
    .A2(_11428_));
 sg13g2_nor3_1 _20525_ (.A(_11417_),
    .B(_11420_),
    .C(_11434_),
    .Y(_11435_));
 sg13g2_nand2b_1 _20526_ (.Y(_11436_),
    .B(_11383_),
    .A_N(net845));
 sg13g2_xnor2_1 _20527_ (.Y(_11437_),
    .A(_10685_),
    .B(net834));
 sg13g2_xnor2_1 _20528_ (.Y(_11438_),
    .A(net844),
    .B(_11437_));
 sg13g2_xor2_1 _20529_ (.B(_11438_),
    .A(_11353_),
    .X(_11439_));
 sg13g2_xnor2_1 _20530_ (.Y(_11440_),
    .A(net846),
    .B(_11439_));
 sg13g2_nor2b_1 _20531_ (.A(_11383_),
    .B_N(net845),
    .Y(_11441_));
 sg13g2_nor2_1 _20532_ (.A(_11017_),
    .B(_11439_),
    .Y(_11442_));
 sg13g2_or2_1 _20533_ (.X(_11443_),
    .B(_11442_),
    .A(_11441_));
 sg13g2_a21oi_1 _20534_ (.A1(_11436_),
    .A2(_11440_),
    .Y(_11444_),
    .B1(_11443_));
 sg13g2_xnor2_1 _20535_ (.Y(_11445_),
    .A(_11435_),
    .B(_11444_));
 sg13g2_inv_2 _20536_ (.Y(_11446_),
    .A(net834));
 sg13g2_nor2_1 _20537_ (.A(_11446_),
    .B(net852),
    .Y(_11447_));
 sg13g2_nand2_1 _20538_ (.Y(_11448_),
    .A(net236),
    .B(net232));
 sg13g2_xor2_1 _20539_ (.B(_11412_),
    .A(net844),
    .X(_11449_));
 sg13g2_nand2_1 _20540_ (.Y(_11450_),
    .A(net507),
    .B(_11449_));
 sg13g2_o21ai_1 _20541_ (.B1(_11450_),
    .Y(_11451_),
    .A1(net507),
    .A2(_11448_));
 sg13g2_a22oi_1 _20542_ (.Y(_11452_),
    .B1(_11451_),
    .B2(net240),
    .A2(_11447_),
    .A1(net141));
 sg13g2_nor2b_1 _20543_ (.A(_11452_),
    .B_N(net486),
    .Y(_11453_));
 sg13g2_xor2_1 _20544_ (.B(net846),
    .A(net1107),
    .X(_11454_));
 sg13g2_nor3_1 _20545_ (.A(_11017_),
    .B(_11383_),
    .C(_11454_),
    .Y(_11455_));
 sg13g2_nor2b_1 _20546_ (.A(_11439_),
    .B_N(_11455_),
    .Y(_11456_));
 sg13g2_nand4_1 _20547_ (.B(net240),
    .C(net141),
    .A(net242),
    .Y(_11457_),
    .D(net138));
 sg13g2_o21ai_1 _20548_ (.B1(net118),
    .Y(_11458_),
    .A1(net486),
    .A2(_11457_));
 sg13g2_xnor2_1 _20549_ (.Y(_11459_),
    .A(_11056_),
    .B(_11399_));
 sg13g2_xnor2_1 _20550_ (.Y(_11460_),
    .A(net845),
    .B(_11459_));
 sg13g2_xnor2_1 _20551_ (.Y(_11461_),
    .A(_11439_),
    .B(_11460_));
 sg13g2_nor2_1 _20552_ (.A(net497),
    .B(_11461_),
    .Y(_11462_));
 sg13g2_nor4_1 _20553_ (.A(_11453_),
    .B(_11456_),
    .C(_11458_),
    .D(_11462_),
    .Y(_11463_));
 sg13g2_a22oi_1 _20554_ (.Y(_11464_),
    .B1(_11445_),
    .B2(_11463_),
    .A2(net67),
    .A1(net497));
 sg13g2_o21ai_1 _20555_ (.B1(net522),
    .Y(_11465_),
    .A1(net38),
    .A2(_11404_));
 sg13g2_a21oi_1 _20556_ (.A1(_11404_),
    .A2(_11464_),
    .Y(_00414_),
    .B1(_11465_));
 sg13g2_buf_2 _20557_ (.A(\grid.cell_25_2.se ),
    .X(_11466_));
 sg13g2_inv_1 _20558_ (.Y(_11467_),
    .A(_11466_));
 sg13g2_xnor2_1 _20559_ (.Y(_11468_),
    .A(_11467_),
    .B(_11119_));
 sg13g2_xor2_1 _20560_ (.B(_11468_),
    .A(_11437_),
    .X(_11469_));
 sg13g2_buf_2 _20561_ (.A(_11469_),
    .X(_11470_));
 sg13g2_buf_2 _20562_ (.A(_00015_),
    .X(_11471_));
 sg13g2_buf_1 _20563_ (.A(_11471_),
    .X(_11472_));
 sg13g2_nor2_1 _20564_ (.A(net496),
    .B(net833),
    .Y(_11473_));
 sg13g2_nand2_1 _20565_ (.Y(_11474_),
    .A(net496),
    .B(net833));
 sg13g2_o21ai_1 _20566_ (.B1(_11474_),
    .Y(_11475_),
    .A1(net507),
    .A2(_11473_));
 sg13g2_inv_1 _20567_ (.Y(_11476_),
    .A(net833));
 sg13g2_nor2_1 _20568_ (.A(net838),
    .B(net484),
    .Y(_11477_));
 sg13g2_a22oi_1 _20569_ (.Y(_11478_),
    .B1(_11477_),
    .B2(net509),
    .A2(_11475_),
    .A1(_11470_));
 sg13g2_a21o_1 _20570_ (.A2(_11470_),
    .A1(net497),
    .B1(net484),
    .X(_11479_));
 sg13g2_a22oi_1 _20571_ (.Y(_11480_),
    .B1(_11479_),
    .B2(net242),
    .A2(_11473_),
    .A1(_11470_));
 sg13g2_buf_1 _20572_ (.A(_11466_),
    .X(_11481_));
 sg13g2_xor2_1 _20573_ (.B(net832),
    .A(net1105),
    .X(_11482_));
 sg13g2_nand2_1 _20574_ (.Y(_11483_),
    .A(net1105),
    .B(net832));
 sg13g2_buf_2 _20575_ (.A(_11483_),
    .X(_11484_));
 sg13g2_a22oi_1 _20576_ (.Y(_11485_),
    .B1(_11484_),
    .B2(_10739_),
    .A2(_11482_),
    .A1(net854));
 sg13g2_nand2_1 _20577_ (.Y(_11486_),
    .A(net854),
    .B(net853));
 sg13g2_nand3_1 _20578_ (.B(_11467_),
    .C(_11486_),
    .A(_11162_),
    .Y(_11487_));
 sg13g2_o21ai_1 _20579_ (.B1(_11487_),
    .Y(_11488_),
    .A1(_10813_),
    .A2(_11485_));
 sg13g2_buf_1 _20580_ (.A(net832),
    .X(_11489_));
 sg13g2_buf_1 _20581_ (.A(net483),
    .X(_11490_));
 sg13g2_a21oi_1 _20582_ (.A1(net854),
    .A2(net485),
    .Y(_11491_),
    .B1(_10739_));
 sg13g2_nor4_1 _20583_ (.A(net842),
    .B(_10813_),
    .C(net231),
    .D(_11491_),
    .Y(_11492_));
 sg13g2_a21oi_2 _20584_ (.B1(_11492_),
    .Y(_11493_),
    .A2(_11488_),
    .A1(_11446_));
 sg13g2_mux2_1 _20585_ (.A0(_11478_),
    .A1(_11480_),
    .S(_11493_),
    .X(_11494_));
 sg13g2_nand3_1 _20586_ (.B(net838),
    .C(_11473_),
    .A(net242),
    .Y(_11495_));
 sg13g2_or2_1 _20587_ (.X(_11496_),
    .B(_11495_),
    .A(_11470_));
 sg13g2_nand2_1 _20588_ (.Y(_11497_),
    .A(net505),
    .B(_11482_));
 sg13g2_o21ai_1 _20589_ (.B1(_11497_),
    .Y(_11498_),
    .A1(net240),
    .A2(_11484_));
 sg13g2_nand2_1 _20590_ (.Y(_11499_),
    .A(net504),
    .B(_11498_));
 sg13g2_o21ai_1 _20591_ (.B1(_11499_),
    .Y(_11500_),
    .A1(_10796_),
    .A2(_11484_));
 sg13g2_nor3_1 _20592_ (.A(net138),
    .B(_11484_),
    .C(_11486_),
    .Y(_11501_));
 sg13g2_nand2b_1 _20593_ (.Y(_11502_),
    .B(net1054),
    .A_N(_11501_));
 sg13g2_a21oi_1 _20594_ (.A1(net138),
    .A2(_11500_),
    .Y(_11503_),
    .B1(_11502_));
 sg13g2_xnor2_1 _20595_ (.Y(_11504_),
    .A(net848),
    .B(_11353_));
 sg13g2_xnor2_1 _20596_ (.Y(_11505_),
    .A(_11470_),
    .B(_11504_));
 sg13g2_nand2_1 _20597_ (.Y(_11506_),
    .A(net127),
    .B(_11505_));
 sg13g2_a22oi_1 _20598_ (.Y(_11507_),
    .B1(_11506_),
    .B2(_11085_),
    .A2(_11408_),
    .A1(_04067_));
 sg13g2_nand4_1 _20599_ (.B(_11496_),
    .C(_11503_),
    .A(_11494_),
    .Y(_11508_),
    .D(_11507_));
 sg13g2_nand2_1 _20600_ (.Y(_11509_),
    .A(net497),
    .B(_11477_));
 sg13g2_a21oi_1 _20601_ (.A1(net509),
    .A2(net833),
    .Y(_11510_),
    .B1(net497));
 sg13g2_nor2_1 _20602_ (.A(net838),
    .B(_11510_),
    .Y(_11511_));
 sg13g2_mux2_1 _20603_ (.A0(_11509_),
    .A1(_11511_),
    .S(_11493_),
    .X(_11512_));
 sg13g2_nand2_1 _20604_ (.Y(_11513_),
    .A(_11000_),
    .B(net843));
 sg13g2_nand3_1 _20605_ (.B(net838),
    .C(net484),
    .A(net496),
    .Y(_11514_));
 sg13g2_o21ai_1 _20606_ (.B1(_11514_),
    .Y(_11515_),
    .A1(_11493_),
    .A2(_11513_));
 sg13g2_nand2_1 _20607_ (.Y(_11516_),
    .A(net509),
    .B(_11515_));
 sg13g2_a21oi_1 _20608_ (.A1(_11512_),
    .A2(_11516_),
    .Y(_11517_),
    .B1(_11470_));
 sg13g2_nand3_1 _20609_ (.B(net110),
    .C(_11404_),
    .A(net141),
    .Y(_11518_));
 sg13g2_o21ai_1 _20610_ (.B1(_11518_),
    .Y(_11519_),
    .A1(net35),
    .A2(_11404_));
 sg13g2_nand2_1 _20611_ (.Y(_11520_),
    .A(net312),
    .B(_11519_));
 sg13g2_o21ai_1 _20612_ (.B1(_11520_),
    .Y(_00415_),
    .A1(_11508_),
    .A2(_11517_));
 sg13g2_buf_2 _20613_ (.A(\grid.cell_25_3.se ),
    .X(_11521_));
 sg13g2_buf_1 _20614_ (.A(_11521_),
    .X(_11522_));
 sg13g2_a21oi_1 _20615_ (.A1(net841),
    .A2(net853),
    .Y(_11523_),
    .B1(_10805_));
 sg13g2_nor3_1 _20616_ (.A(net832),
    .B(net831),
    .C(_11523_),
    .Y(_11524_));
 sg13g2_xor2_1 _20617_ (.B(_11521_),
    .A(_11466_),
    .X(_11525_));
 sg13g2_nand2_1 _20618_ (.Y(_11526_),
    .A(net853),
    .B(_11525_));
 sg13g2_nand2_2 _20619_ (.Y(_11527_),
    .A(_11466_),
    .B(_11521_));
 sg13g2_nand2_1 _20620_ (.Y(_11528_),
    .A(_10805_),
    .B(_11527_));
 sg13g2_a21oi_1 _20621_ (.A1(_11526_),
    .A2(_11528_),
    .Y(_11529_),
    .B1(net841));
 sg13g2_or2_1 _20622_ (.X(_11530_),
    .B(_11529_),
    .A(_11524_));
 sg13g2_buf_1 _20623_ (.A(net831),
    .X(_11531_));
 sg13g2_nor3_1 _20624_ (.A(net841),
    .B(net483),
    .C(net482),
    .Y(_11532_));
 sg13g2_a22oi_1 _20625_ (.Y(_11533_),
    .B1(_11532_),
    .B2(_10808_),
    .A2(_11530_),
    .A1(_10844_));
 sg13g2_buf_1 _20626_ (.A(_11533_),
    .X(_11534_));
 sg13g2_buf_1 _20627_ (.A(_00014_),
    .X(_11535_));
 sg13g2_buf_1 _20628_ (.A(_11535_),
    .X(_11536_));
 sg13g2_nor2_1 _20629_ (.A(net1104),
    .B(net830),
    .Y(_11537_));
 sg13g2_and2_1 _20630_ (.A(net141),
    .B(_11537_),
    .X(_11538_));
 sg13g2_a21oi_1 _20631_ (.A1(_11085_),
    .A2(_11534_),
    .Y(_11539_),
    .B1(_11538_));
 sg13g2_nand3_1 _20632_ (.B(net1104),
    .C(net830),
    .A(_11116_),
    .Y(_11540_));
 sg13g2_inv_1 _20633_ (.Y(_11541_),
    .A(net830));
 sg13g2_a21oi_1 _20634_ (.A1(net237),
    .A2(_11541_),
    .Y(_11542_),
    .B1(_11174_));
 sg13g2_mux2_1 _20635_ (.A0(_11540_),
    .A1(_11542_),
    .S(_11534_),
    .X(_11543_));
 sg13g2_o21ai_1 _20636_ (.B1(_11543_),
    .Y(_11544_),
    .A1(_10705_),
    .A2(_11539_));
 sg13g2_nand2_1 _20637_ (.Y(_11545_),
    .A(net237),
    .B(_11537_));
 sg13g2_nand3b_1 _20638_ (.B(net1104),
    .C(_11116_),
    .Y(_11546_),
    .A_N(_11534_));
 sg13g2_a21oi_1 _20639_ (.A1(_11545_),
    .A2(_11546_),
    .Y(_11547_),
    .B1(net240));
 sg13g2_xnor2_1 _20640_ (.Y(_11548_),
    .A(_10783_),
    .B(_11154_));
 sg13g2_xnor2_1 _20641_ (.Y(_11549_),
    .A(net831),
    .B(_11548_));
 sg13g2_xnor2_1 _20642_ (.Y(_11550_),
    .A(net853),
    .B(net832));
 sg13g2_xnor2_1 _20643_ (.Y(_11551_),
    .A(_11549_),
    .B(_11550_));
 sg13g2_buf_1 _20644_ (.A(_11551_),
    .X(_11552_));
 sg13g2_o21ai_1 _20645_ (.B1(_11552_),
    .Y(_11553_),
    .A1(_11544_),
    .A2(_11547_));
 sg13g2_nand2b_1 _20646_ (.Y(_11554_),
    .B(net236),
    .A_N(_11535_));
 sg13g2_nor2b_1 _20647_ (.A(net238),
    .B_N(_11535_),
    .Y(_11555_));
 sg13g2_a21oi_1 _20648_ (.A1(_10705_),
    .A2(_11554_),
    .Y(_11556_),
    .B1(_11555_));
 sg13g2_nand3_1 _20649_ (.B(net1104),
    .C(net830),
    .A(_10705_),
    .Y(_11557_));
 sg13g2_o21ai_1 _20650_ (.B1(_11557_),
    .Y(_11558_),
    .A1(_11552_),
    .A2(_11556_));
 sg13g2_o21ai_1 _20651_ (.B1(net830),
    .Y(_11559_),
    .A1(net237),
    .A2(_11552_));
 sg13g2_nand2_1 _20652_ (.Y(_11560_),
    .A(net240),
    .B(_11559_));
 sg13g2_o21ai_1 _20653_ (.B1(_11560_),
    .Y(_11561_),
    .A1(_11552_),
    .A2(_11554_));
 sg13g2_mux2_1 _20654_ (.A0(_11558_),
    .A1(_11561_),
    .S(_11534_),
    .X(_11562_));
 sg13g2_xor2_1 _20655_ (.B(_11552_),
    .A(_11438_),
    .X(_11563_));
 sg13g2_a21oi_1 _20656_ (.A1(net126),
    .A2(_11563_),
    .Y(_11564_),
    .B1(net491));
 sg13g2_o21ai_1 _20657_ (.B1(_11526_),
    .Y(_11565_),
    .A1(net504),
    .A2(_11527_));
 sg13g2_nor3_1 _20658_ (.A(net492),
    .B(_10739_),
    .C(_11527_),
    .Y(_11566_));
 sg13g2_a21oi_1 _20659_ (.A1(net492),
    .A2(_11565_),
    .Y(_11567_),
    .B1(_11566_));
 sg13g2_nor2_1 _20660_ (.A(net502),
    .B(_11567_),
    .Y(_11568_));
 sg13g2_nand4_1 _20661_ (.B(net492),
    .C(net231),
    .A(_10853_),
    .Y(_11569_),
    .D(net482));
 sg13g2_nand3_1 _20662_ (.B(_11404_),
    .C(_11569_),
    .A(net1002),
    .Y(_11570_));
 sg13g2_nor4_1 _20663_ (.A(_11562_),
    .B(_11564_),
    .C(_11568_),
    .D(_11570_),
    .Y(_11571_));
 sg13g2_nand4_1 _20664_ (.B(net491),
    .C(net104),
    .A(net1056),
    .Y(_11572_),
    .D(_11404_));
 sg13g2_o21ai_1 _20665_ (.B1(_11572_),
    .Y(_11573_),
    .A1(net32),
    .A2(_11409_));
 sg13g2_a21o_1 _20666_ (.A2(_11571_),
    .A1(_11553_),
    .B1(_11573_),
    .X(_00416_));
 sg13g2_buf_2 _20667_ (.A(\grid.cell_25_4.se ),
    .X(_11574_));
 sg13g2_xor2_1 _20668_ (.B(_11574_),
    .A(_11521_),
    .X(_11575_));
 sg13g2_buf_1 _20669_ (.A(_11574_),
    .X(_11576_));
 sg13g2_nand2_1 _20670_ (.Y(_11577_),
    .A(net831),
    .B(net829));
 sg13g2_nor2_1 _20671_ (.A(net851),
    .B(_11577_),
    .Y(_11578_));
 sg13g2_a21oi_1 _20672_ (.A1(net851),
    .A2(_11575_),
    .Y(_11579_),
    .B1(_11578_));
 sg13g2_inv_1 _20673_ (.Y(_11580_),
    .A(_11577_));
 sg13g2_nand3_1 _20674_ (.B(net503),
    .C(_11580_),
    .A(net490),
    .Y(_11581_));
 sg13g2_o21ai_1 _20675_ (.B1(_11581_),
    .Y(_11582_),
    .A1(_11210_),
    .A2(_11579_));
 sg13g2_nor2_1 _20676_ (.A(_10884_),
    .B(_11210_),
    .Y(_11583_));
 sg13g2_buf_1 _20677_ (.A(_00059_),
    .X(_11584_));
 sg13g2_xnor2_1 _20678_ (.Y(_11585_),
    .A(_10820_),
    .B(net1103));
 sg13g2_xor2_1 _20679_ (.B(_11585_),
    .A(_11575_),
    .X(_11586_));
 sg13g2_xnor2_1 _20680_ (.Y(_11587_),
    .A(net502),
    .B(_11586_));
 sg13g2_nor4_1 _20681_ (.A(_11207_),
    .B(net1101),
    .C(_11119_),
    .D(_11587_),
    .Y(_11588_));
 sg13g2_a221oi_1 _20682_ (.B2(_11580_),
    .C1(_11588_),
    .B1(_11583_),
    .A1(net501),
    .Y(_11589_),
    .A2(_11582_));
 sg13g2_a22oi_1 _20683_ (.Y(_11590_),
    .B1(_11577_),
    .B2(net500),
    .A2(_11575_),
    .A1(net851));
 sg13g2_inv_2 _20684_ (.Y(_11591_),
    .A(net831));
 sg13g2_inv_1 _20685_ (.Y(_11592_),
    .A(_11574_));
 sg13g2_buf_1 _20686_ (.A(_11592_),
    .X(_11593_));
 sg13g2_o21ai_1 _20687_ (.B1(net850),
    .Y(_11594_),
    .A1(_11209_),
    .A2(net502));
 sg13g2_nand3_1 _20688_ (.B(net481),
    .C(_11594_),
    .A(_11591_),
    .Y(_11595_));
 sg13g2_o21ai_1 _20689_ (.B1(_11595_),
    .Y(_11596_),
    .A1(net840),
    .A2(_11590_));
 sg13g2_buf_1 _20690_ (.A(net829),
    .X(_11597_));
 sg13g2_nor3_1 _20691_ (.A(net840),
    .B(net482),
    .C(net480),
    .Y(_11598_));
 sg13g2_nand2_1 _20692_ (.Y(_11599_),
    .A(net501),
    .B(net503));
 sg13g2_a22oi_1 _20693_ (.Y(_11600_),
    .B1(_11598_),
    .B2(_11599_),
    .A2(_11596_),
    .A1(_10884_));
 sg13g2_nand2_1 _20694_ (.Y(_11601_),
    .A(net1101),
    .B(_10739_));
 sg13g2_xnor2_1 _20695_ (.Y(_11602_),
    .A(_11139_),
    .B(_11587_));
 sg13g2_inv_1 _20696_ (.Y(_11603_),
    .A(net1101));
 sg13g2_nand2_1 _20697_ (.Y(_11604_),
    .A(_11603_),
    .B(net504));
 sg13g2_o21ai_1 _20698_ (.B1(_11604_),
    .Y(_11605_),
    .A1(_11207_),
    .A2(_11587_));
 sg13g2_a21oi_1 _20699_ (.A1(_11601_),
    .A2(_11602_),
    .Y(_11606_),
    .B1(_11605_));
 sg13g2_xnor2_1 _20700_ (.Y(_11607_),
    .A(_11600_),
    .B(_11606_));
 sg13g2_buf_1 _20701_ (.A(net168),
    .X(_11608_));
 sg13g2_a21oi_1 _20702_ (.A1(_11589_),
    .A2(_11607_),
    .Y(_11609_),
    .B1(net96));
 sg13g2_xnor2_1 _20703_ (.Y(_11610_),
    .A(_11468_),
    .B(_11587_));
 sg13g2_a21oi_1 _20704_ (.A1(net68),
    .A2(_11610_),
    .Y(_11611_),
    .B1(_11179_));
 sg13g2_or3_1 _20705_ (.A(_11405_),
    .B(_11609_),
    .C(_11611_),
    .X(_11612_));
 sg13g2_o21ai_1 _20706_ (.B1(_11612_),
    .Y(_00417_),
    .A1(net34),
    .A2(_11409_));
 sg13g2_buf_1 _20707_ (.A(\grid.cell_25_5.se ),
    .X(_11613_));
 sg13g2_buf_1 _20708_ (.A(net1100),
    .X(_11614_));
 sg13g2_nand2_2 _20709_ (.Y(_11615_),
    .A(net829),
    .B(net828));
 sg13g2_xnor2_1 _20710_ (.Y(_11616_),
    .A(_11574_),
    .B(net1100));
 sg13g2_nor2_1 _20711_ (.A(net500),
    .B(_11616_),
    .Y(_11617_));
 sg13g2_nor2_1 _20712_ (.A(net850),
    .B(_11615_),
    .Y(_11618_));
 sg13g2_o21ai_1 _20713_ (.B1(net498),
    .Y(_11619_),
    .A1(_11617_),
    .A2(_11618_));
 sg13g2_o21ai_1 _20714_ (.B1(_11619_),
    .Y(_11620_),
    .A1(_10944_),
    .A2(_11615_));
 sg13g2_xnor2_1 _20715_ (.Y(_11621_),
    .A(_11236_),
    .B(_11616_));
 sg13g2_xnor2_1 _20716_ (.Y(_11622_),
    .A(_10820_),
    .B(_11621_));
 sg13g2_and2_1 _20717_ (.A(_11233_),
    .B(_11622_),
    .X(_11623_));
 sg13g2_buf_2 _20718_ (.A(_00091_),
    .X(_11624_));
 sg13g2_nor2b_1 _20719_ (.A(_11624_),
    .B_N(_11548_),
    .Y(_11625_));
 sg13g2_nor3_1 _20720_ (.A(net234),
    .B(_10876_),
    .C(_11615_),
    .Y(_11626_));
 sg13g2_a221oi_1 _20721_ (.B2(_11625_),
    .C1(_11626_),
    .B1(_11623_),
    .A1(_11255_),
    .Y(_11627_),
    .A2(_11620_));
 sg13g2_a21oi_1 _20722_ (.A1(net499),
    .A2(_11615_),
    .Y(_11628_),
    .B1(_11617_));
 sg13g2_buf_1 _20723_ (.A(net828),
    .X(_11629_));
 sg13g2_a21oi_1 _20724_ (.A1(net839),
    .A2(_10820_),
    .Y(_11630_),
    .B1(_10871_));
 sg13g2_or3_1 _20725_ (.A(net829),
    .B(net479),
    .C(_11630_),
    .X(_11631_));
 sg13g2_o21ai_1 _20726_ (.B1(_11631_),
    .Y(_11632_),
    .A1(_11243_),
    .A2(_11628_));
 sg13g2_nor3_1 _20727_ (.A(net480),
    .B(net479),
    .C(_10905_),
    .Y(_11633_));
 sg13g2_a22oi_1 _20728_ (.Y(_11634_),
    .B1(_11633_),
    .B2(_11247_),
    .A2(_11632_),
    .A1(_10944_));
 sg13g2_nand2_1 _20729_ (.Y(_11635_),
    .A(_11624_),
    .B(net502));
 sg13g2_xnor2_1 _20730_ (.Y(_11636_),
    .A(net235),
    .B(_11622_));
 sg13g2_nor2_1 _20731_ (.A(_11624_),
    .B(net502),
    .Y(_11637_));
 sg13g2_a221oi_1 _20732_ (.B2(_11636_),
    .C1(_11637_),
    .B1(_11635_),
    .A1(_11233_),
    .Y(_11638_),
    .A2(_11622_));
 sg13g2_xnor2_1 _20733_ (.Y(_11639_),
    .A(_11634_),
    .B(_11638_));
 sg13g2_a21oi_1 _20734_ (.A1(_11627_),
    .A2(_11639_),
    .Y(_11640_),
    .B1(net96));
 sg13g2_xor2_1 _20735_ (.B(_11622_),
    .A(_11549_),
    .X(_11641_));
 sg13g2_a21oi_1 _20736_ (.A1(net68),
    .A2(_11641_),
    .Y(_11642_),
    .B1(net489));
 sg13g2_or3_1 _20737_ (.A(_11405_),
    .B(_11640_),
    .C(_11642_),
    .X(_11643_));
 sg13g2_o21ai_1 _20738_ (.B1(_11643_),
    .Y(_00418_),
    .A1(net46),
    .A2(_11409_));
 sg13g2_buf_2 _20739_ (.A(_00152_),
    .X(_11644_));
 sg13g2_nand2_1 _20740_ (.Y(_11645_),
    .A(net1100),
    .B(net1102));
 sg13g2_buf_1 _20741_ (.A(_11645_),
    .X(_11646_));
 sg13g2_nor2_2 _20742_ (.A(_11644_),
    .B(net478),
    .Y(_11647_));
 sg13g2_nor2_1 _20743_ (.A(net1100),
    .B(net1102),
    .Y(_11648_));
 sg13g2_buf_1 _20744_ (.A(_11648_),
    .X(_11649_));
 sg13g2_xnor2_1 _20745_ (.Y(_11650_),
    .A(_11644_),
    .B(net239));
 sg13g2_nand3_1 _20746_ (.B(net239),
    .C(net478),
    .A(_11644_),
    .Y(_11651_));
 sg13g2_o21ai_1 _20747_ (.B1(_11651_),
    .Y(_11652_),
    .A1(_11649_),
    .A2(_11650_));
 sg13g2_nor2_1 _20748_ (.A(net506),
    .B(net499),
    .Y(_11653_));
 sg13g2_o21ai_1 _20749_ (.B1(_11653_),
    .Y(_11654_),
    .A1(_11647_),
    .A2(_11652_));
 sg13g2_nand2_1 _20750_ (.Y(_11655_),
    .A(_11038_),
    .B(_11649_));
 sg13g2_o21ai_1 _20751_ (.B1(_11655_),
    .Y(_11656_),
    .A1(_11273_),
    .A2(net478));
 sg13g2_a21oi_1 _20752_ (.A1(net479),
    .A2(net837),
    .Y(_11657_),
    .B1(net494));
 sg13g2_o21ai_1 _20753_ (.B1(_11644_),
    .Y(_11658_),
    .A1(_11649_),
    .A2(_11657_));
 sg13g2_a21oi_1 _20754_ (.A1(_11655_),
    .A2(_11658_),
    .Y(_11659_),
    .B1(net241));
 sg13g2_a221oi_1 _20755_ (.B2(net499),
    .C1(_11659_),
    .B1(_11656_),
    .A1(net140),
    .Y(_11660_),
    .A2(_11647_));
 sg13g2_nand2_1 _20756_ (.Y(_11661_),
    .A(_11654_),
    .B(_11660_));
 sg13g2_buf_2 _20757_ (.A(_00123_),
    .X(_11662_));
 sg13g2_nand2_1 _20758_ (.Y(_11663_),
    .A(_11662_),
    .B(net500));
 sg13g2_xnor2_1 _20759_ (.Y(_11664_),
    .A(net1100),
    .B(net1102));
 sg13g2_xnor2_1 _20760_ (.Y(_11665_),
    .A(_10870_),
    .B(_11664_));
 sg13g2_xnor2_1 _20761_ (.Y(_11666_),
    .A(_11005_),
    .B(_11665_));
 sg13g2_xnor2_1 _20762_ (.Y(_11667_),
    .A(net489),
    .B(_11666_));
 sg13g2_inv_1 _20763_ (.Y(_11668_),
    .A(_11662_));
 sg13g2_nand2_1 _20764_ (.Y(_11669_),
    .A(_11668_),
    .B(net501));
 sg13g2_o21ai_1 _20765_ (.B1(_11669_),
    .Y(_11670_),
    .A1(_11280_),
    .A2(_11666_));
 sg13g2_a21oi_1 _20766_ (.A1(_11663_),
    .A2(_11667_),
    .Y(_11671_),
    .B1(_11670_));
 sg13g2_xor2_1 _20767_ (.B(_11671_),
    .A(_11661_),
    .X(_11672_));
 sg13g2_mux2_1 _20768_ (.A0(net478),
    .A1(_11664_),
    .S(net849),
    .X(_11673_));
 sg13g2_nor2_1 _20769_ (.A(net506),
    .B(_11673_),
    .Y(_11674_));
 sg13g2_or2_1 _20770_ (.X(_11675_),
    .B(_11674_),
    .A(_11647_));
 sg13g2_nor2_1 _20771_ (.A(_11034_),
    .B(net478),
    .Y(_11676_));
 sg13g2_nand2_1 _20772_ (.Y(_11677_),
    .A(_11668_),
    .B(_11585_));
 sg13g2_nor3_1 _20773_ (.A(_11280_),
    .B(_11666_),
    .C(_11677_),
    .Y(_11678_));
 sg13g2_a221oi_1 _20774_ (.B2(net498),
    .C1(_11678_),
    .B1(_11676_),
    .A1(net140),
    .Y(_11679_),
    .A2(_11675_));
 sg13g2_a21oi_1 _20775_ (.A1(_11672_),
    .A2(_11679_),
    .Y(_11680_),
    .B1(net79));
 sg13g2_xnor2_1 _20776_ (.Y(_11681_),
    .A(net480),
    .B(_11585_));
 sg13g2_xnor2_1 _20777_ (.Y(_11682_),
    .A(_11666_),
    .B(_11681_));
 sg13g2_a21oi_1 _20778_ (.A1(net122),
    .A2(_11682_),
    .Y(_11683_),
    .B1(net234));
 sg13g2_or2_1 _20779_ (.X(_11684_),
    .B(_11683_),
    .A(_11405_));
 sg13g2_nand2b_1 _20780_ (.Y(_11685_),
    .B(net31),
    .A_N(_11409_));
 sg13g2_o21ai_1 _20781_ (.B1(_11685_),
    .Y(_00419_),
    .A1(_11680_),
    .A2(_11684_));
 sg13g2_buf_1 _20782_ (.A(net479),
    .X(_11686_));
 sg13g2_nand3_1 _20783_ (.B(net233),
    .C(_11653_),
    .A(_11686_),
    .Y(_11687_));
 sg13g2_xnor2_1 _20784_ (.Y(_11688_),
    .A(_11235_),
    .B(net858));
 sg13g2_xnor2_1 _20785_ (.Y(_11689_),
    .A(_11665_),
    .B(_11688_));
 sg13g2_a22oi_1 _20786_ (.Y(_11690_),
    .B1(_11689_),
    .B2(_11455_),
    .A2(_11675_),
    .A1(net234));
 sg13g2_o21ai_1 _20787_ (.B1(_11690_),
    .Y(_11691_),
    .A1(net234),
    .A2(_11687_));
 sg13g2_xnor2_1 _20788_ (.Y(_11692_),
    .A(_11644_),
    .B(net839));
 sg13g2_nand3_1 _20789_ (.B(net488),
    .C(net478),
    .A(_11644_),
    .Y(_11693_));
 sg13g2_o21ai_1 _20790_ (.B1(_11693_),
    .Y(_11694_),
    .A1(_11649_),
    .A2(_11692_));
 sg13g2_o21ai_1 _20791_ (.B1(_11653_),
    .Y(_11695_),
    .A1(_11647_),
    .A2(_11694_));
 sg13g2_nand2_1 _20792_ (.Y(_11696_),
    .A(net839),
    .B(net508));
 sg13g2_nand2_1 _20793_ (.Y(_11697_),
    .A(_11247_),
    .B(_11649_));
 sg13g2_o21ai_1 _20794_ (.B1(_11697_),
    .Y(_11698_),
    .A1(net478),
    .A2(_11696_));
 sg13g2_a21oi_1 _20795_ (.A1(net828),
    .A2(net837),
    .Y(_11699_),
    .B1(net839));
 sg13g2_o21ai_1 _20796_ (.B1(_11644_),
    .Y(_11700_),
    .A1(_11649_),
    .A2(_11699_));
 sg13g2_a21oi_1 _20797_ (.A1(_11697_),
    .A2(_11700_),
    .Y(_11701_),
    .B1(net241));
 sg13g2_a221oi_1 _20798_ (.B2(net499),
    .C1(_11701_),
    .B1(_11698_),
    .A1(net488),
    .Y(_11702_),
    .A2(_11647_));
 sg13g2_nand2_1 _20799_ (.Y(_11703_),
    .A(_11695_),
    .B(_11702_));
 sg13g2_inv_1 _20800_ (.Y(_11704_),
    .A(net846));
 sg13g2_xnor2_1 _20801_ (.Y(_11705_),
    .A(_11704_),
    .B(_11689_));
 sg13g2_a221oi_1 _20802_ (.B2(_11436_),
    .C1(_11441_),
    .B1(_11705_),
    .A1(_11031_),
    .Y(_11706_),
    .A2(_11689_));
 sg13g2_xnor2_1 _20803_ (.Y(_11707_),
    .A(_11703_),
    .B(_11706_));
 sg13g2_o21ai_1 _20804_ (.B1(net82),
    .Y(_11708_),
    .A1(_11691_),
    .A2(_11707_));
 sg13g2_xor2_1 _20805_ (.B(_11689_),
    .A(_11460_),
    .X(_11709_));
 sg13g2_a21oi_1 _20806_ (.A1(net98),
    .A2(_11709_),
    .Y(_11710_),
    .B1(net140));
 sg13g2_nor2_1 _20807_ (.A(_11408_),
    .B(_11710_),
    .Y(_11711_));
 sg13g2_a22oi_1 _20808_ (.Y(_11712_),
    .B1(_11708_),
    .B2(_11711_),
    .A2(_11408_),
    .A1(net80));
 sg13g2_nor2_1 _20809_ (.A(net370),
    .B(_11712_),
    .Y(_00420_));
 sg13g2_or2_1 _20810_ (.X(_11713_),
    .B(_10992_),
    .A(_10239_));
 sg13g2_buf_1 _20811_ (.A(_11713_),
    .X(_11714_));
 sg13g2_buf_1 _20812_ (.A(_11399_),
    .X(_11715_));
 sg13g2_buf_2 _20813_ (.A(\grid.cell_26_0.se ),
    .X(_11716_));
 sg13g2_xnor2_1 _20814_ (.Y(_11717_),
    .A(net1106),
    .B(_11716_));
 sg13g2_buf_2 _20815_ (.A(\grid.cell_26_0.sw ),
    .X(_11718_));
 sg13g2_xnor2_1 _20816_ (.Y(_11719_),
    .A(net1102),
    .B(_11718_));
 sg13g2_buf_2 _20817_ (.A(_11719_),
    .X(_11720_));
 sg13g2_xnor2_1 _20818_ (.Y(_11721_),
    .A(_11717_),
    .B(_11720_));
 sg13g2_xnor2_1 _20819_ (.Y(_11722_),
    .A(net494),
    .B(_11721_));
 sg13g2_nand2_1 _20820_ (.Y(_11723_),
    .A(_11704_),
    .B(_00013_));
 sg13g2_xor2_1 _20821_ (.B(_11722_),
    .A(net486),
    .X(_11724_));
 sg13g2_buf_1 _20822_ (.A(_00013_),
    .X(_11725_));
 sg13g2_nor2_1 _20823_ (.A(_11704_),
    .B(net1099),
    .Y(_11726_));
 sg13g2_a221oi_1 _20824_ (.B2(_11724_),
    .C1(_11726_),
    .B1(_11723_),
    .A1(net484),
    .Y(_11727_),
    .A2(_11722_));
 sg13g2_buf_1 _20825_ (.A(_11716_),
    .X(_11728_));
 sg13g2_buf_1 _20826_ (.A(net826),
    .X(_11729_));
 sg13g2_nor2_1 _20827_ (.A(net1102),
    .B(_11718_),
    .Y(_11730_));
 sg13g2_buf_1 _20828_ (.A(_11730_),
    .X(_11731_));
 sg13g2_inv_1 _20829_ (.Y(_11732_),
    .A(_11731_));
 sg13g2_and2_1 _20830_ (.A(net1102),
    .B(_11718_),
    .X(_11733_));
 sg13g2_buf_2 _20831_ (.A(_11733_),
    .X(_11734_));
 sg13g2_nand3_1 _20832_ (.B(net140),
    .C(_11734_),
    .A(net477),
    .Y(_11735_));
 sg13g2_o21ai_1 _20833_ (.B1(_11735_),
    .Y(_11736_),
    .A1(net477),
    .A2(_11732_));
 sg13g2_buf_1 _20834_ (.A(_11718_),
    .X(_11737_));
 sg13g2_nand2_1 _20835_ (.Y(_11738_),
    .A(_11350_),
    .B(net825));
 sg13g2_buf_1 _20836_ (.A(_11738_),
    .X(_11739_));
 sg13g2_nor2_1 _20837_ (.A(net843),
    .B(_11739_),
    .Y(_11740_));
 sg13g2_buf_1 _20838_ (.A(net477),
    .X(_11741_));
 sg13g2_o21ai_1 _20839_ (.B1(_11732_),
    .Y(_11742_),
    .A1(net838),
    .A2(_11734_));
 sg13g2_inv_1 _20840_ (.Y(_11743_),
    .A(net826));
 sg13g2_buf_1 _20841_ (.A(_11743_),
    .X(_11744_));
 sg13g2_a22oi_1 _20842_ (.Y(_11745_),
    .B1(_11742_),
    .B2(net228),
    .A2(_11731_),
    .A1(net843));
 sg13g2_nor2_1 _20843_ (.A(net826),
    .B(_11739_),
    .Y(_11746_));
 sg13g2_xnor2_1 _20844_ (.Y(_11747_),
    .A(net826),
    .B(_11128_));
 sg13g2_nand3_1 _20845_ (.B(_11128_),
    .C(_11739_),
    .A(net826),
    .Y(_11748_));
 sg13g2_o21ai_1 _20846_ (.B1(_11748_),
    .Y(_11749_),
    .A1(_11731_),
    .A2(_11747_));
 sg13g2_o21ai_1 _20847_ (.B1(_11044_),
    .Y(_11750_),
    .A1(_11746_),
    .A2(_11749_));
 sg13g2_o21ai_1 _20848_ (.B1(_11750_),
    .Y(_11751_),
    .A1(net140),
    .A2(_11745_));
 sg13g2_a221oi_1 _20849_ (.B2(net229),
    .C1(_11751_),
    .B1(_11740_),
    .A1(net496),
    .Y(_11752_),
    .A2(_11736_));
 sg13g2_xnor2_1 _20850_ (.Y(_11753_),
    .A(_11727_),
    .B(_11752_));
 sg13g2_buf_1 _20851_ (.A(\grid.cell_26_0.s ),
    .X(_11754_));
 sg13g2_buf_1 _20852_ (.A(_11754_),
    .X(_11755_));
 sg13g2_xor2_1 _20853_ (.B(_11352_),
    .A(net846),
    .X(_11756_));
 sg13g2_xnor2_1 _20854_ (.Y(_11757_),
    .A(net824),
    .B(_11756_));
 sg13g2_xnor2_1 _20855_ (.Y(_11758_),
    .A(_11722_),
    .B(_11757_));
 sg13g2_nor2_1 _20856_ (.A(net827),
    .B(_11758_),
    .Y(_11759_));
 sg13g2_nand2_1 _20857_ (.Y(_11760_),
    .A(net484),
    .B(_11722_));
 sg13g2_nor3_1 _20858_ (.A(net1099),
    .B(_11756_),
    .C(_11760_),
    .Y(_11761_));
 sg13g2_nand2b_1 _20859_ (.Y(_11762_),
    .B(net1106),
    .A_N(_11720_));
 sg13g2_o21ai_1 _20860_ (.B1(_11762_),
    .Y(_11763_),
    .A1(net848),
    .A2(_11739_));
 sg13g2_a21oi_1 _20861_ (.A1(net140),
    .A2(_11763_),
    .Y(_11764_),
    .B1(_11740_));
 sg13g2_a21oi_1 _20862_ (.A1(_11044_),
    .A2(_11734_),
    .Y(_11765_),
    .B1(net229));
 sg13g2_a21oi_1 _20863_ (.A1(net229),
    .A2(_11764_),
    .Y(_11766_),
    .B1(_11765_));
 sg13g2_nor4_1 _20864_ (.A(net107),
    .B(_11759_),
    .C(_11761_),
    .D(_11766_),
    .Y(_11767_));
 sg13g2_a22oi_1 _20865_ (.Y(_11768_),
    .B1(_11753_),
    .B2(_11767_),
    .A2(net67),
    .A1(net827));
 sg13g2_o21ai_1 _20866_ (.B1(net522),
    .Y(_11769_),
    .A1(net40),
    .A2(net65));
 sg13g2_a21oi_1 _20867_ (.A1(net65),
    .A2(_11768_),
    .Y(_00421_),
    .B1(_11769_));
 sg13g2_buf_1 _20868_ (.A(\grid.cell_26_1.se ),
    .X(_11770_));
 sg13g2_xor2_1 _20869_ (.B(_11449_),
    .A(net1098),
    .X(_11771_));
 sg13g2_xor2_1 _20870_ (.B(_11771_),
    .A(_11717_),
    .X(_11772_));
 sg13g2_buf_2 _20871_ (.A(_11772_),
    .X(_11773_));
 sg13g2_xnor2_1 _20872_ (.Y(_11774_),
    .A(_11400_),
    .B(_11773_));
 sg13g2_o21ai_1 _20873_ (.B1(net846),
    .Y(_11775_),
    .A1(_11400_),
    .A2(_11383_));
 sg13g2_nor2_1 _20874_ (.A(net846),
    .B(_11383_),
    .Y(_11776_));
 sg13g2_o21ai_1 _20875_ (.B1(net827),
    .Y(_11777_),
    .A1(_11773_),
    .A2(_11776_));
 sg13g2_nand3b_1 _20876_ (.B(_11400_),
    .C(_11383_),
    .Y(_11778_),
    .A_N(_11773_));
 sg13g2_nand3_1 _20877_ (.B(_11777_),
    .C(_11778_),
    .A(_11775_),
    .Y(_11779_));
 sg13g2_o21ai_1 _20878_ (.B1(net1099),
    .Y(_11780_),
    .A1(_11383_),
    .A2(_11773_));
 sg13g2_o21ai_1 _20879_ (.B1(_11780_),
    .Y(_11781_),
    .A1(net1099),
    .A2(_11779_));
 sg13g2_o21ai_1 _20880_ (.B1(_11781_),
    .Y(_11782_),
    .A1(_11704_),
    .A2(_11774_));
 sg13g2_xor2_1 _20881_ (.B(net1098),
    .A(net834),
    .X(_11783_));
 sg13g2_buf_1 _20882_ (.A(net1098),
    .X(_11784_));
 sg13g2_buf_1 _20883_ (.A(net823),
    .X(_11785_));
 sg13g2_a21oi_1 _20884_ (.A1(net232),
    .A2(net476),
    .Y(_11786_),
    .B1(net236));
 sg13g2_a21o_1 _20885_ (.A2(_11783_),
    .A1(net848),
    .B1(_11786_),
    .X(_11787_));
 sg13g2_nand2_2 _20886_ (.Y(_11788_),
    .A(net1106),
    .B(net493));
 sg13g2_nor2_1 _20887_ (.A(net485),
    .B(net823),
    .Y(_11789_));
 sg13g2_a22oi_1 _20888_ (.Y(_11790_),
    .B1(_11788_),
    .B2(_11789_),
    .A2(_11787_),
    .A1(net843));
 sg13g2_o21ai_1 _20889_ (.B1(net141),
    .Y(_11791_),
    .A1(net496),
    .A2(net228));
 sg13g2_nand3_1 _20890_ (.B(_11789_),
    .C(_11791_),
    .A(net843),
    .Y(_11792_));
 sg13g2_o21ai_1 _20891_ (.B1(_11792_),
    .Y(_11793_),
    .A1(net229),
    .A2(_11790_));
 sg13g2_nand2_1 _20892_ (.Y(_11794_),
    .A(_11743_),
    .B(_11789_));
 sg13g2_buf_1 _20893_ (.A(net476),
    .X(_11795_));
 sg13g2_nand4_1 _20894_ (.B(net238),
    .C(net138),
    .A(net477),
    .Y(_11796_),
    .D(net227));
 sg13g2_a21oi_1 _20895_ (.A1(_11794_),
    .A2(_11796_),
    .Y(_11797_),
    .B1(net497));
 sg13g2_nor4_1 _20896_ (.A(net141),
    .B(net138),
    .C(net227),
    .D(net838),
    .Y(_11798_));
 sg13g2_nand2_1 _20897_ (.Y(_11799_),
    .A(net823),
    .B(net838));
 sg13g2_o21ai_1 _20898_ (.B1(_11799_),
    .Y(_11800_),
    .A1(net476),
    .A2(_11788_));
 sg13g2_nor2_1 _20899_ (.A(net476),
    .B(net843),
    .Y(_11801_));
 sg13g2_nor3_1 _20900_ (.A(net232),
    .B(_11788_),
    .C(_11801_),
    .Y(_11802_));
 sg13g2_a21oi_1 _20901_ (.A1(net138),
    .A2(_11800_),
    .Y(_11803_),
    .B1(_11802_));
 sg13g2_nor2_1 _20902_ (.A(net823),
    .B(_11349_),
    .Y(_11804_));
 sg13g2_a21oi_1 _20903_ (.A1(_11446_),
    .A2(_11799_),
    .Y(_11805_),
    .B1(_11804_));
 sg13g2_nor2_1 _20904_ (.A(net238),
    .B(_11805_),
    .Y(_11806_));
 sg13g2_nand2_1 _20905_ (.Y(_11807_),
    .A(net476),
    .B(net843));
 sg13g2_o21ai_1 _20906_ (.B1(net485),
    .Y(_11808_),
    .A1(net823),
    .A2(_11128_));
 sg13g2_a21oi_1 _20907_ (.A1(_11807_),
    .A2(_11808_),
    .Y(_11809_),
    .B1(_11788_));
 sg13g2_o21ai_1 _20908_ (.B1(net228),
    .Y(_11810_),
    .A1(_11806_),
    .A2(_11809_));
 sg13g2_o21ai_1 _20909_ (.B1(_11810_),
    .Y(_11811_),
    .A1(net228),
    .A2(_11803_));
 sg13g2_o21ai_1 _20910_ (.B1(_11384_),
    .Y(_11812_),
    .A1(_11788_),
    .A2(_11794_));
 sg13g2_xnor2_1 _20911_ (.Y(_11813_),
    .A(net237),
    .B(_11717_));
 sg13g2_xor2_1 _20912_ (.B(net493),
    .A(net826),
    .X(_11814_));
 sg13g2_nand3_1 _20913_ (.B(net826),
    .C(_11084_),
    .A(net1106),
    .Y(_11815_));
 sg13g2_o21ai_1 _20914_ (.B1(_11815_),
    .Y(_11816_),
    .A1(net1106),
    .A2(_11814_));
 sg13g2_nor2_1 _20915_ (.A(_11783_),
    .B(_11816_),
    .Y(_11817_));
 sg13g2_a21oi_1 _20916_ (.A1(_11783_),
    .A2(_11813_),
    .Y(_11818_),
    .B1(_11817_));
 sg13g2_nor2_1 _20917_ (.A(_11812_),
    .B(_11818_),
    .Y(_11819_));
 sg13g2_nor4_1 _20918_ (.A(_11797_),
    .B(_11798_),
    .C(_11811_),
    .D(_11819_),
    .Y(_11820_));
 sg13g2_nor2_1 _20919_ (.A(net1099),
    .B(_11774_),
    .Y(_11821_));
 sg13g2_nand2_1 _20920_ (.Y(_11822_),
    .A(net1099),
    .B(_11774_));
 sg13g2_o21ai_1 _20921_ (.B1(_11822_),
    .Y(_11823_),
    .A1(net846),
    .A2(_11821_));
 sg13g2_a221oi_1 _20922_ (.B2(_11823_),
    .C1(net69),
    .B1(_11820_),
    .A1(_11782_),
    .Y(_11824_),
    .A2(_11793_));
 sg13g2_xnor2_1 _20923_ (.Y(_11825_),
    .A(net824),
    .B(_11459_));
 sg13g2_xnor2_1 _20924_ (.Y(_11826_),
    .A(_11773_),
    .B(_11825_));
 sg13g2_a21oi_1 _20925_ (.A1(net112),
    .A2(_11826_),
    .Y(_11827_),
    .B1(net486));
 sg13g2_nand2_1 _20926_ (.Y(_11828_),
    .A(_12956_),
    .B(net65));
 sg13g2_or2_1 _20927_ (.X(_11829_),
    .B(_11828_),
    .A(_11827_));
 sg13g2_nor2_1 _20928_ (.A(_10239_),
    .B(_10992_),
    .Y(_11830_));
 sg13g2_nand2_1 _20929_ (.Y(_11831_),
    .A(net1056),
    .B(_11830_));
 sg13g2_nand2b_1 _20930_ (.Y(_11832_),
    .B(net42),
    .A_N(_11831_));
 sg13g2_o21ai_1 _20931_ (.B1(_11832_),
    .Y(_00422_),
    .A1(_11824_),
    .A2(_11829_));
 sg13g2_buf_1 _20932_ (.A(_00012_),
    .X(_11833_));
 sg13g2_inv_2 _20933_ (.Y(_11834_),
    .A(net1097));
 sg13g2_buf_2 _20934_ (.A(\grid.cell_26_2.se ),
    .X(_11835_));
 sg13g2_xnor2_1 _20935_ (.Y(_11836_),
    .A(_11466_),
    .B(_11835_));
 sg13g2_buf_2 _20936_ (.A(_11836_),
    .X(_11837_));
 sg13g2_xnor2_1 _20937_ (.Y(_11838_),
    .A(_11124_),
    .B(_11837_));
 sg13g2_xnor2_1 _20938_ (.Y(_11839_),
    .A(net1098),
    .B(_11838_));
 sg13g2_buf_1 _20939_ (.A(_11839_),
    .X(_11840_));
 sg13g2_xor2_1 _20940_ (.B(_11840_),
    .A(net836),
    .X(_11841_));
 sg13g2_o21ai_1 _20941_ (.B1(_11841_),
    .Y(_11842_),
    .A1(net497),
    .A2(_11834_));
 sg13g2_buf_1 _20942_ (.A(_11835_),
    .X(_11843_));
 sg13g2_and2_1 _20943_ (.A(net832),
    .B(net822),
    .X(_11844_));
 sg13g2_nand2_1 _20944_ (.Y(_11845_),
    .A(net832),
    .B(net822));
 sg13g2_nand2b_1 _20945_ (.Y(_11846_),
    .B(net844),
    .A_N(_11837_));
 sg13g2_o21ai_1 _20946_ (.B1(_11846_),
    .Y(_11847_),
    .A1(net493),
    .A2(_11845_));
 sg13g2_a22oi_1 _20947_ (.Y(_11848_),
    .B1(_11847_),
    .B2(net491),
    .A2(_11844_),
    .A1(_11174_));
 sg13g2_nand2b_1 _20948_ (.Y(_11849_),
    .B(net227),
    .A_N(_11848_));
 sg13g2_nand2_1 _20949_ (.Y(_11850_),
    .A(net484),
    .B(_11840_));
 sg13g2_buf_1 _20950_ (.A(net823),
    .X(_11851_));
 sg13g2_nor3_1 _20951_ (.A(net237),
    .B(net475),
    .C(_11484_),
    .Y(_11852_));
 sg13g2_buf_1 _20952_ (.A(net822),
    .X(_11853_));
 sg13g2_buf_1 _20953_ (.A(net474),
    .X(_11854_));
 sg13g2_a22oi_1 _20954_ (.Y(_11855_),
    .B1(_11852_),
    .B2(net226),
    .A2(_11834_),
    .A1(net848));
 sg13g2_and4_1 _20955_ (.A(_11842_),
    .B(_11849_),
    .C(_11850_),
    .D(_11855_),
    .X(_11856_));
 sg13g2_buf_1 _20956_ (.A(net1097),
    .X(_11857_));
 sg13g2_o21ai_1 _20957_ (.B1(_11840_),
    .Y(_11858_),
    .A1(net848),
    .A2(net833));
 sg13g2_nor2_1 _20958_ (.A(_11362_),
    .B(net484),
    .Y(_11859_));
 sg13g2_a21oi_1 _20959_ (.A1(net835),
    .A2(net484),
    .Y(_11860_),
    .B1(net496));
 sg13g2_a221oi_1 _20960_ (.B2(_11840_),
    .C1(_11860_),
    .B1(_11859_),
    .A1(_11375_),
    .Y(_11861_),
    .A2(_11858_));
 sg13g2_and2_1 _20961_ (.A(_11476_),
    .B(_11840_),
    .X(_11862_));
 sg13g2_a22oi_1 _20962_ (.Y(_11863_),
    .B1(_11862_),
    .B2(net821),
    .A2(_11841_),
    .A1(_11000_));
 sg13g2_o21ai_1 _20963_ (.B1(_11863_),
    .Y(_11864_),
    .A1(net821),
    .A2(_11861_));
 sg13g2_o21ai_1 _20964_ (.B1(_11846_),
    .Y(_11865_),
    .A1(net842),
    .A2(_11844_));
 sg13g2_nand2_1 _20965_ (.Y(_11866_),
    .A(net238),
    .B(net491));
 sg13g2_nor2_1 _20966_ (.A(net483),
    .B(net474),
    .Y(_11867_));
 sg13g2_a22oi_1 _20967_ (.Y(_11868_),
    .B1(_11866_),
    .B2(_11867_),
    .A2(_11865_),
    .A1(net1104));
 sg13g2_a21oi_1 _20968_ (.A1(net238),
    .A2(net475),
    .Y(_11869_),
    .B1(_11162_));
 sg13g2_nand3b_1 _20969_ (.B(_11867_),
    .C(net1104),
    .Y(_11870_),
    .A_N(_11869_));
 sg13g2_o21ai_1 _20970_ (.B1(_11870_),
    .Y(_11871_),
    .A1(net227),
    .A2(_11868_));
 sg13g2_mux2_1 _20971_ (.A0(_11856_),
    .A1(_11864_),
    .S(_11871_),
    .X(_11872_));
 sg13g2_xnor2_1 _20972_ (.Y(_11873_),
    .A(_11717_),
    .B(_11841_));
 sg13g2_a21oi_1 _20973_ (.A1(net114),
    .A2(_11873_),
    .Y(_11874_),
    .B1(_11416_));
 sg13g2_nor2_1 _20974_ (.A(_11828_),
    .B(_11874_),
    .Y(_11875_));
 sg13g2_o21ai_1 _20975_ (.B1(_11875_),
    .Y(_11876_),
    .A1(net81),
    .A2(_11872_));
 sg13g2_o21ai_1 _20976_ (.B1(_11876_),
    .Y(_00423_),
    .A1(net27),
    .A2(_11831_));
 sg13g2_buf_1 _20977_ (.A(\grid.cell_26_3.se ),
    .X(_11877_));
 sg13g2_buf_1 _20978_ (.A(_11877_),
    .X(_11878_));
 sg13g2_inv_2 _20979_ (.Y(_11879_),
    .A(net820));
 sg13g2_xnor2_1 _20980_ (.Y(_11880_),
    .A(_11835_),
    .B(_11521_));
 sg13g2_xnor2_1 _20981_ (.Y(_11881_),
    .A(_11155_),
    .B(_11880_));
 sg13g2_xnor2_1 _20982_ (.Y(_11882_),
    .A(_11879_),
    .B(_11881_));
 sg13g2_xnor2_1 _20983_ (.Y(_11883_),
    .A(_11771_),
    .B(_11882_));
 sg13g2_a21oi_1 _20984_ (.A1(net84),
    .A2(_11883_),
    .Y(_11884_),
    .B1(net231));
 sg13g2_buf_1 _20985_ (.A(net820),
    .X(_11885_));
 sg13g2_buf_1 _20986_ (.A(net473),
    .X(_11886_));
 sg13g2_nand2_1 _20987_ (.Y(_11887_),
    .A(net822),
    .B(net831));
 sg13g2_nand2b_1 _20988_ (.Y(_11888_),
    .B(net842),
    .A_N(_11880_));
 sg13g2_o21ai_1 _20989_ (.B1(_11888_),
    .Y(_11889_),
    .A1(net842),
    .A2(_11887_));
 sg13g2_nor3_1 _20990_ (.A(_11162_),
    .B(net473),
    .C(_11887_),
    .Y(_11890_));
 sg13g2_a21oi_1 _20991_ (.A1(net225),
    .A2(_11889_),
    .Y(_11891_),
    .B1(_11890_));
 sg13g2_nor2_1 _20992_ (.A(net235),
    .B(_11891_),
    .Y(_11892_));
 sg13g2_buf_1 _20993_ (.A(_00011_),
    .X(_11893_));
 sg13g2_nor4_1 _20994_ (.A(_11893_),
    .B(net830),
    .C(_11449_),
    .D(_11882_),
    .Y(_11894_));
 sg13g2_nor3_1 _20995_ (.A(_11207_),
    .B(_11879_),
    .C(_11887_),
    .Y(_11895_));
 sg13g2_nor4_1 _20996_ (.A(_11828_),
    .B(_11892_),
    .C(_11894_),
    .D(_11895_),
    .Y(_11896_));
 sg13g2_nand2_1 _20997_ (.Y(_11897_),
    .A(net237),
    .B(_11893_));
 sg13g2_xnor2_1 _20998_ (.Y(_11898_),
    .A(_11415_),
    .B(_11882_));
 sg13g2_inv_1 _20999_ (.Y(_11899_),
    .A(_11893_));
 sg13g2_nand2_1 _21000_ (.Y(_11900_),
    .A(_11100_),
    .B(_11899_));
 sg13g2_o21ai_1 _21001_ (.B1(_11900_),
    .Y(_11901_),
    .A1(net830),
    .A2(_11882_));
 sg13g2_a21oi_1 _21002_ (.A1(_11897_),
    .A2(_11898_),
    .Y(_11902_),
    .B1(_11901_));
 sg13g2_xor2_1 _21003_ (.B(_11877_),
    .A(_11521_),
    .X(_11903_));
 sg13g2_nand2_1 _21004_ (.Y(_11904_),
    .A(net831),
    .B(net820));
 sg13g2_a22oi_1 _21005_ (.Y(_11905_),
    .B1(_11904_),
    .B2(net235),
    .A2(_11903_),
    .A1(net842));
 sg13g2_a21oi_1 _21006_ (.A1(net1105),
    .A2(net822),
    .Y(_11906_),
    .B1(net235));
 sg13g2_or3_1 _21007_ (.A(net482),
    .B(net473),
    .C(_11906_),
    .X(_11907_));
 sg13g2_o21ai_1 _21008_ (.B1(_11907_),
    .Y(_11908_),
    .A1(net474),
    .A2(_11905_));
 sg13g2_nor3_1 _21009_ (.A(_11854_),
    .B(net482),
    .C(net473),
    .Y(_11909_));
 sg13g2_a22oi_1 _21010_ (.Y(_11910_),
    .B1(_11909_),
    .B2(_11181_),
    .A2(_11908_),
    .A1(_11207_));
 sg13g2_xnor2_1 _21011_ (.Y(_11911_),
    .A(_11902_),
    .B(_11910_));
 sg13g2_a22oi_1 _21012_ (.Y(_11912_),
    .B1(_11896_),
    .B2(_11911_),
    .A2(net65),
    .A1(_08877_));
 sg13g2_or2_1 _21013_ (.X(_11913_),
    .B(_11912_),
    .A(_11884_));
 sg13g2_o21ai_1 _21014_ (.B1(_11913_),
    .Y(_00424_),
    .A1(net26),
    .A2(net65));
 sg13g2_nand3_1 _21015_ (.B(net104),
    .C(net65),
    .A(net482),
    .Y(_11914_));
 sg13g2_o21ai_1 _21016_ (.B1(_11914_),
    .Y(_11915_),
    .A1(net47),
    .A2(net65));
 sg13g2_buf_1 _21017_ (.A(\grid.cell_26_4.se ),
    .X(_11916_));
 sg13g2_xor2_1 _21018_ (.B(net1096),
    .A(_11574_),
    .X(_11917_));
 sg13g2_buf_1 _21019_ (.A(net1096),
    .X(_11918_));
 sg13g2_nand2_1 _21020_ (.Y(_11919_),
    .A(net829),
    .B(net819));
 sg13g2_a22oi_1 _21021_ (.Y(_11920_),
    .B1(_11919_),
    .B2(_11209_),
    .A2(_11917_),
    .A1(net841));
 sg13g2_inv_2 _21022_ (.Y(_11921_),
    .A(_11916_));
 sg13g2_o21ai_1 _21023_ (.B1(net840),
    .Y(_11922_),
    .A1(_11160_),
    .A2(_11879_));
 sg13g2_nand3_1 _21024_ (.B(_11921_),
    .C(_11922_),
    .A(net481),
    .Y(_11923_));
 sg13g2_o21ai_1 _21025_ (.B1(_11923_),
    .Y(_11924_),
    .A1(net473),
    .A2(_11920_));
 sg13g2_nor3_1 _21026_ (.A(net473),
    .B(net829),
    .C(net819),
    .Y(_11925_));
 sg13g2_a22oi_1 _21027_ (.Y(_11926_),
    .B1(_11925_),
    .B2(_11197_),
    .A2(_11924_),
    .A1(_11232_));
 sg13g2_buf_1 _21028_ (.A(_11926_),
    .X(_11927_));
 sg13g2_buf_2 _21029_ (.A(_00058_),
    .X(_11928_));
 sg13g2_nor2_1 _21030_ (.A(_11928_),
    .B(_11484_),
    .Y(_11929_));
 sg13g2_o21ai_1 _21031_ (.B1(_11603_),
    .Y(_11930_),
    .A1(_11927_),
    .A2(_11929_));
 sg13g2_a21oi_1 _21032_ (.A1(_11928_),
    .A2(_11162_),
    .Y(_11931_),
    .B1(net231));
 sg13g2_nand2_1 _21033_ (.Y(_11932_),
    .A(_11927_),
    .B(_11931_));
 sg13g2_xnor2_1 _21034_ (.Y(_11933_),
    .A(net820),
    .B(_11574_));
 sg13g2_xor2_1 _21035_ (.B(_11933_),
    .A(_11213_),
    .X(_11934_));
 sg13g2_xnor2_1 _21036_ (.Y(_11935_),
    .A(_11921_),
    .B(_11934_));
 sg13g2_buf_2 _21037_ (.A(_11935_),
    .X(_11936_));
 sg13g2_a21oi_1 _21038_ (.A1(_11930_),
    .A2(_11932_),
    .Y(_11937_),
    .B1(_11936_));
 sg13g2_inv_1 _21039_ (.Y(_11938_),
    .A(_11928_));
 sg13g2_a21o_1 _21040_ (.A2(_11936_),
    .A1(net231),
    .B1(net491),
    .X(_11939_));
 sg13g2_nor2b_1 _21041_ (.A(_11484_),
    .B_N(_11936_),
    .Y(_11940_));
 sg13g2_a21oi_1 _21042_ (.A1(_11938_),
    .A2(_11939_),
    .Y(_11941_),
    .B1(_11940_));
 sg13g2_o21ai_1 _21043_ (.B1(_11928_),
    .Y(_11942_),
    .A1(net1101),
    .A2(_11936_));
 sg13g2_or3_1 _21044_ (.A(net1101),
    .B(_11928_),
    .C(net231),
    .X(_11943_));
 sg13g2_a21oi_1 _21045_ (.A1(_11942_),
    .A2(_11943_),
    .Y(_11944_),
    .B1(net491));
 sg13g2_nand3b_1 _21046_ (.B(_11490_),
    .C(net1101),
    .Y(_11945_),
    .A_N(_11936_));
 sg13g2_nand2b_1 _21047_ (.Y(_11946_),
    .B(_11936_),
    .A_N(_11490_));
 sg13g2_a22oi_1 _21048_ (.Y(_11947_),
    .B1(_11945_),
    .B2(_11946_),
    .A2(_11180_),
    .A1(_11938_));
 sg13g2_nor3_1 _21049_ (.A(_11927_),
    .B(_11944_),
    .C(_11947_),
    .Y(_11948_));
 sg13g2_a21oi_1 _21050_ (.A1(_11927_),
    .A2(_11941_),
    .Y(_11949_),
    .B1(_11948_));
 sg13g2_buf_1 _21051_ (.A(_11918_),
    .X(_11950_));
 sg13g2_nand4_1 _21052_ (.B(net225),
    .C(net480),
    .A(_11233_),
    .Y(_11951_),
    .D(net472));
 sg13g2_xnor2_1 _21053_ (.Y(_11952_),
    .A(net842),
    .B(_11837_));
 sg13g2_xnor2_1 _21054_ (.Y(_11953_),
    .A(_11936_),
    .B(_11952_));
 sg13g2_nand2_1 _21055_ (.Y(_11954_),
    .A(net172),
    .B(_11953_));
 sg13g2_nand3_1 _21056_ (.B(net225),
    .C(_11597_),
    .A(net492),
    .Y(_11955_));
 sg13g2_nor2_1 _21057_ (.A(net235),
    .B(_11933_),
    .Y(_11956_));
 sg13g2_nor3_1 _21058_ (.A(net492),
    .B(_11879_),
    .C(_11593_),
    .Y(_11957_));
 sg13g2_o21ai_1 _21059_ (.B1(net472),
    .Y(_11958_),
    .A1(_11956_),
    .A2(_11957_));
 sg13g2_o21ai_1 _21060_ (.B1(_11958_),
    .Y(_11959_),
    .A1(_11950_),
    .A2(_11955_));
 sg13g2_a22oi_1 _21061_ (.Y(_11960_),
    .B1(_11959_),
    .B2(net489),
    .A2(_11954_),
    .A1(_11591_));
 sg13g2_nand4_1 _21062_ (.B(_11714_),
    .C(_11951_),
    .A(net1056),
    .Y(_11961_),
    .D(_11960_));
 sg13g2_nor3_1 _21063_ (.A(_11937_),
    .B(_11949_),
    .C(_11961_),
    .Y(_11962_));
 sg13g2_a21o_1 _21064_ (.A2(_11915_),
    .A1(net312),
    .B1(_11962_),
    .X(_00425_));
 sg13g2_nand2_1 _21065_ (.Y(_11963_),
    .A(_06330_),
    .B(_11830_));
 sg13g2_nor2_1 _21066_ (.A(_11161_),
    .B(_11591_),
    .Y(_11964_));
 sg13g2_o21ai_1 _21067_ (.B1(_11624_),
    .Y(_11965_),
    .A1(_11161_),
    .A2(net831));
 sg13g2_buf_1 _21068_ (.A(\grid.cell_26_5.se ),
    .X(_11966_));
 sg13g2_xor2_1 _21069_ (.B(_11966_),
    .A(net1100),
    .X(_11967_));
 sg13g2_buf_2 _21070_ (.A(_11967_),
    .X(_11968_));
 sg13g2_xnor2_1 _21071_ (.Y(_11969_),
    .A(_11235_),
    .B(net1096));
 sg13g2_xnor2_1 _21072_ (.Y(_11970_),
    .A(_11968_),
    .B(_11969_));
 sg13g2_xnor2_1 _21073_ (.Y(_11971_),
    .A(_11209_),
    .B(_11970_));
 sg13g2_mux2_1 _21074_ (.A0(_11964_),
    .A1(_11965_),
    .S(_11971_),
    .X(_11972_));
 sg13g2_buf_1 _21075_ (.A(_11966_),
    .X(_11973_));
 sg13g2_nand2_1 _21076_ (.Y(_11974_),
    .A(net1100),
    .B(net818));
 sg13g2_a22oi_1 _21077_ (.Y(_11975_),
    .B1(_11968_),
    .B2(net840),
    .A2(_11974_),
    .A1(_11247_));
 sg13g2_nand2_1 _21078_ (.Y(_11976_),
    .A(net1103),
    .B(net1096));
 sg13g2_or2_1 _21079_ (.X(_11977_),
    .B(_11973_),
    .A(net1100));
 sg13g2_a21o_1 _21080_ (.A2(_11976_),
    .A1(_11242_),
    .B1(_11977_),
    .X(_11978_));
 sg13g2_o21ai_1 _21081_ (.B1(_11978_),
    .Y(_11979_),
    .A1(net819),
    .A2(_11975_));
 sg13g2_a21oi_1 _21082_ (.A1(_11242_),
    .A2(net840),
    .Y(_11980_),
    .B1(_11977_));
 sg13g2_a22oi_1 _21083_ (.Y(_11981_),
    .B1(_11980_),
    .B2(_11921_),
    .A2(_11979_),
    .A1(_11280_));
 sg13g2_or2_1 _21084_ (.X(_11982_),
    .B(_11981_),
    .A(_11972_));
 sg13g2_nand2_1 _21085_ (.Y(_11983_),
    .A(_11972_),
    .B(_11981_));
 sg13g2_buf_1 _21086_ (.A(_00090_),
    .X(_11984_));
 sg13g2_xnor2_1 _21087_ (.Y(_11985_),
    .A(_11213_),
    .B(_11970_));
 sg13g2_xnor2_1 _21088_ (.Y(_11986_),
    .A(_11591_),
    .B(_11985_));
 sg13g2_nor2_1 _21089_ (.A(_11984_),
    .B(_11986_),
    .Y(_11987_));
 sg13g2_a21o_1 _21090_ (.A2(_11983_),
    .A1(_11982_),
    .B1(_11987_),
    .X(_11988_));
 sg13g2_buf_1 _21091_ (.A(net818),
    .X(_11989_));
 sg13g2_buf_1 _21092_ (.A(net471),
    .X(_11990_));
 sg13g2_nand3_1 _21093_ (.B(net479),
    .C(net224),
    .A(net819),
    .Y(_11991_));
 sg13g2_nand2_1 _21094_ (.Y(_11992_),
    .A(net819),
    .B(_11968_));
 sg13g2_o21ai_1 _21095_ (.B1(_11992_),
    .Y(_11993_),
    .A1(net819),
    .A2(_11974_));
 sg13g2_nand2_1 _21096_ (.Y(_11994_),
    .A(net489),
    .B(_11993_));
 sg13g2_o21ai_1 _21097_ (.B1(_11994_),
    .Y(_11995_),
    .A1(net489),
    .A2(_11991_));
 sg13g2_nor2_1 _21098_ (.A(_11280_),
    .B(_11991_),
    .Y(_11996_));
 sg13g2_a221oi_1 _21099_ (.B2(_11982_),
    .C1(_11996_),
    .B1(_11987_),
    .A1(_11255_),
    .Y(_11997_),
    .A2(_11995_));
 sg13g2_a21o_1 _21100_ (.A2(_11997_),
    .A1(_11988_),
    .B1(net124),
    .X(_11998_));
 sg13g2_xor2_1 _21101_ (.B(_11985_),
    .A(_11903_),
    .X(_11999_));
 sg13g2_o21ai_1 _21102_ (.B1(net481),
    .Y(_12000_),
    .A1(net97),
    .A2(_11999_));
 sg13g2_nand3_1 _21103_ (.B(_11998_),
    .C(_12000_),
    .A(_11714_),
    .Y(_12001_));
 sg13g2_a21oi_1 _21104_ (.A1(_11963_),
    .A2(_12001_),
    .Y(_00426_),
    .B1(_10200_));
 sg13g2_buf_1 _21105_ (.A(_00153_),
    .X(_12002_));
 sg13g2_buf_1 _21106_ (.A(_12002_),
    .X(_12003_));
 sg13g2_inv_1 _21107_ (.Y(_12004_),
    .A(net818));
 sg13g2_nor2_1 _21108_ (.A(_12004_),
    .B(_11734_),
    .Y(_12005_));
 sg13g2_nor2_1 _21109_ (.A(net817),
    .B(_11739_),
    .Y(_12006_));
 sg13g2_a21oi_1 _21110_ (.A1(net817),
    .A2(_12005_),
    .Y(_12007_),
    .B1(_12006_));
 sg13g2_xor2_1 _21111_ (.B(net471),
    .A(_12002_),
    .X(_12008_));
 sg13g2_nand2_1 _21112_ (.Y(_12009_),
    .A(_11732_),
    .B(_12008_));
 sg13g2_a21oi_1 _21113_ (.A1(_12007_),
    .A2(_12009_),
    .Y(_12010_),
    .B1(_11297_));
 sg13g2_nand2_1 _21114_ (.Y(_12011_),
    .A(net471),
    .B(_11734_));
 sg13g2_nor2_1 _21115_ (.A(net817),
    .B(_12011_),
    .Y(_12012_));
 sg13g2_buf_1 _21116_ (.A(_12004_),
    .X(_12013_));
 sg13g2_nand2_1 _21117_ (.Y(_12014_),
    .A(net223),
    .B(_11731_));
 sg13g2_nand3_1 _21118_ (.B(net471),
    .C(_11734_),
    .A(net494),
    .Y(_12015_));
 sg13g2_a21oi_1 _21119_ (.A1(_12014_),
    .A2(_12015_),
    .Y(_12016_),
    .B1(net488));
 sg13g2_nor2_1 _21120_ (.A(net471),
    .B(_11734_),
    .Y(_12017_));
 sg13g2_o21ai_1 _21121_ (.B1(net817),
    .Y(_12018_),
    .A1(_11731_),
    .A2(_12017_));
 sg13g2_a21oi_1 _21122_ (.A1(_12014_),
    .A2(_12018_),
    .Y(_12019_),
    .B1(net239));
 sg13g2_nor4_2 _21123_ (.A(_12010_),
    .B(_12012_),
    .C(_12016_),
    .Y(_12020_),
    .D(_12019_));
 sg13g2_buf_1 _21124_ (.A(_00122_),
    .X(_12021_));
 sg13g2_a21oi_1 _21125_ (.A1(net1095),
    .A2(net490),
    .Y(_12022_),
    .B1(net480));
 sg13g2_nand2_1 _21126_ (.Y(_12023_),
    .A(_12020_),
    .B(_12022_));
 sg13g2_nor3_1 _21127_ (.A(net1095),
    .B(net490),
    .C(net481),
    .Y(_12024_));
 sg13g2_o21ai_1 _21128_ (.B1(_11668_),
    .Y(_12025_),
    .A1(_12020_),
    .A2(_12024_));
 sg13g2_xnor2_1 _21129_ (.Y(_12026_),
    .A(_11282_),
    .B(_11720_));
 sg13g2_xnor2_1 _21130_ (.Y(_12027_),
    .A(_12004_),
    .B(_12026_));
 sg13g2_buf_2 _21131_ (.A(_12027_),
    .X(_12028_));
 sg13g2_a21oi_1 _21132_ (.A1(_12023_),
    .A2(_12025_),
    .Y(_12029_),
    .B1(_12028_));
 sg13g2_xnor2_1 _21133_ (.Y(_12030_),
    .A(net490),
    .B(_11917_));
 sg13g2_xnor2_1 _21134_ (.Y(_12031_),
    .A(_12028_),
    .B(_12030_));
 sg13g2_nor2_1 _21135_ (.A(net230),
    .B(_12031_),
    .Y(_12032_));
 sg13g2_buf_1 _21136_ (.A(_11737_),
    .X(_12033_));
 sg13g2_buf_1 _21137_ (.A(net470),
    .X(_12034_));
 sg13g2_nor2b_1 _21138_ (.A(net222),
    .B_N(net487),
    .Y(_12035_));
 sg13g2_xor2_1 _21139_ (.B(net487),
    .A(net224),
    .X(_12036_));
 sg13g2_a22oi_1 _21140_ (.Y(_12037_),
    .B1(_12036_),
    .B2(net222),
    .A2(_12035_),
    .A1(net224));
 sg13g2_mux2_1 _21141_ (.A0(_12011_),
    .A1(_12037_),
    .S(net234),
    .X(_12038_));
 sg13g2_nor2_1 _21142_ (.A(_05407_),
    .B(_12012_),
    .Y(_12039_));
 sg13g2_o21ai_1 _21143_ (.B1(_12039_),
    .Y(_12040_),
    .A1(_11038_),
    .A2(_12038_));
 sg13g2_nor3_1 _21144_ (.A(_11668_),
    .B(net481),
    .C(_12028_),
    .Y(_12041_));
 sg13g2_a21oi_1 _21145_ (.A1(net481),
    .A2(_12028_),
    .Y(_12042_),
    .B1(_12041_));
 sg13g2_nor2_1 _21146_ (.A(net1095),
    .B(net490),
    .Y(_12043_));
 sg13g2_o21ai_1 _21147_ (.B1(net1095),
    .Y(_12044_),
    .A1(_11662_),
    .A2(_12028_));
 sg13g2_or3_1 _21148_ (.A(_11662_),
    .B(net1095),
    .C(net829),
    .X(_12045_));
 sg13g2_a21o_1 _21149_ (.A2(_12045_),
    .A1(_12044_),
    .B1(net489),
    .X(_12046_));
 sg13g2_o21ai_1 _21150_ (.B1(_12046_),
    .Y(_12047_),
    .A1(_12042_),
    .A2(_12043_));
 sg13g2_a21oi_1 _21151_ (.A1(net480),
    .A2(_12028_),
    .Y(_12048_),
    .B1(net489));
 sg13g2_nand3_1 _21152_ (.B(net480),
    .C(_12028_),
    .A(net489),
    .Y(_12049_));
 sg13g2_o21ai_1 _21153_ (.B1(_12049_),
    .Y(_12050_),
    .A1(net1095),
    .A2(_12048_));
 sg13g2_mux2_1 _21154_ (.A0(_12047_),
    .A1(_12050_),
    .S(_12020_),
    .X(_12051_));
 sg13g2_or4_1 _21155_ (.A(_12029_),
    .B(_12032_),
    .C(_12040_),
    .D(_12051_),
    .X(_12052_));
 sg13g2_a21oi_1 _21156_ (.A1(net230),
    .A2(net73),
    .Y(_12053_),
    .B1(_11830_));
 sg13g2_o21ai_1 _21157_ (.B1(net522),
    .Y(_12054_),
    .A1(net31),
    .A2(net65));
 sg13g2_a21oi_1 _21158_ (.A1(_12052_),
    .A2(_12053_),
    .Y(_00427_),
    .B1(_12054_));
 sg13g2_xor2_1 _21159_ (.B(_11968_),
    .A(_11282_),
    .X(_12055_));
 sg13g2_xnor2_1 _21160_ (.Y(_12056_),
    .A(net825),
    .B(_12055_));
 sg13g2_xnor2_1 _21161_ (.Y(_12057_),
    .A(_11400_),
    .B(_12056_));
 sg13g2_a221oi_1 _21162_ (.B2(_11723_),
    .C1(_11726_),
    .B1(_12057_),
    .A1(_11384_),
    .Y(_12058_),
    .A2(_12056_));
 sg13g2_nor2_1 _21163_ (.A(net471),
    .B(net470),
    .Y(_12059_));
 sg13g2_xor2_1 _21164_ (.B(_11614_),
    .A(net817),
    .X(_12060_));
 sg13g2_nand2b_1 _21165_ (.Y(_12061_),
    .B(_12060_),
    .A_N(_12059_));
 sg13g2_nand2_1 _21166_ (.Y(_12062_),
    .A(net817),
    .B(net828));
 sg13g2_nand2_1 _21167_ (.Y(_12063_),
    .A(net818),
    .B(net825));
 sg13g2_mux2_1 _21168_ (.A0(net817),
    .A1(_12062_),
    .S(_12063_),
    .X(_12064_));
 sg13g2_a21oi_1 _21169_ (.A1(_12061_),
    .A2(_12064_),
    .Y(_12065_),
    .B1(_11297_));
 sg13g2_and2_1 _21170_ (.A(_11966_),
    .B(net825),
    .X(_12066_));
 sg13g2_buf_1 _21171_ (.A(_12066_),
    .X(_12067_));
 sg13g2_nand2_1 _21172_ (.Y(_12068_),
    .A(net828),
    .B(_12067_));
 sg13g2_nor2_1 _21173_ (.A(_12003_),
    .B(_12068_),
    .Y(_12069_));
 sg13g2_nand2b_1 _21174_ (.Y(_12070_),
    .B(_12059_),
    .A_N(_11629_));
 sg13g2_nand3_1 _21175_ (.B(_11629_),
    .C(_12067_),
    .A(net494),
    .Y(_12071_));
 sg13g2_a21oi_1 _21176_ (.A1(_12070_),
    .A2(_12071_),
    .Y(_12072_),
    .B1(net488));
 sg13g2_nor2_1 _21177_ (.A(_11614_),
    .B(_12067_),
    .Y(_12073_));
 sg13g2_o21ai_1 _21178_ (.B1(net817),
    .Y(_12074_),
    .A1(_12059_),
    .A2(_12073_));
 sg13g2_a21oi_1 _21179_ (.A1(_12070_),
    .A2(_12074_),
    .Y(_12075_),
    .B1(_11367_));
 sg13g2_nor4_1 _21180_ (.A(_12065_),
    .B(_12069_),
    .C(_12072_),
    .D(_12075_),
    .Y(_12076_));
 sg13g2_xnor2_1 _21181_ (.Y(_12077_),
    .A(_12058_),
    .B(_12076_));
 sg13g2_and2_1 _21182_ (.A(net470),
    .B(_11968_),
    .X(_12078_));
 sg13g2_nor2_1 _21183_ (.A(net222),
    .B(_11974_),
    .Y(_12079_));
 sg13g2_o21ai_1 _21184_ (.B1(net488),
    .Y(_12080_),
    .A1(_12078_),
    .A2(_12079_));
 sg13g2_o21ai_1 _21185_ (.B1(_12080_),
    .Y(_12081_),
    .A1(net234),
    .A2(_12068_));
 sg13g2_nand2_1 _21186_ (.Y(_12082_),
    .A(_11367_),
    .B(_12081_));
 sg13g2_inv_1 _21187_ (.Y(_12083_),
    .A(net1099));
 sg13g2_nand4_1 _21188_ (.B(_11384_),
    .C(_11459_),
    .A(_12083_),
    .Y(_12084_),
    .D(_12056_));
 sg13g2_nor2_1 _21189_ (.A(net163),
    .B(_12069_),
    .Y(_12085_));
 sg13g2_and4_1 _21190_ (.A(_12077_),
    .B(_12082_),
    .C(_12084_),
    .D(_12085_),
    .X(_12086_));
 sg13g2_nor2_1 _21191_ (.A(net79),
    .B(_12086_),
    .Y(_12087_));
 sg13g2_nor3_1 _21192_ (.A(_08349_),
    .B(_11347_),
    .C(_10992_),
    .Y(_12088_));
 sg13g2_nor2_1 _21193_ (.A(net1057),
    .B(_12088_),
    .Y(_12089_));
 sg13g2_nand2_1 _21194_ (.Y(_12090_),
    .A(_11364_),
    .B(_12089_));
 sg13g2_nor3_1 _21195_ (.A(_08349_),
    .B(_11340_),
    .C(_10992_),
    .Y(_12091_));
 sg13g2_xnor2_1 _21196_ (.Y(_12092_),
    .A(_11825_),
    .B(_12056_));
 sg13g2_nor3_1 _21197_ (.A(net1057),
    .B(_12088_),
    .C(_12092_),
    .Y(_12093_));
 sg13g2_a22oi_1 _21198_ (.Y(_12094_),
    .B1(_12086_),
    .B2(_12093_),
    .A2(_12091_),
    .A1(_12089_));
 sg13g2_o21ai_1 _21199_ (.B1(_12094_),
    .Y(_00428_),
    .A1(_12087_),
    .A2(_12090_));
 sg13g2_buf_2 _21200_ (.A(\grid.cell_27_0.sw ),
    .X(_12095_));
 sg13g2_nor2b_1 _21201_ (.A(_12095_),
    .B_N(_11471_),
    .Y(_12096_));
 sg13g2_buf_1 _21202_ (.A(\grid.cell_27_0.se ),
    .X(_12097_));
 sg13g2_buf_2 _21203_ (.A(_12097_),
    .X(_12098_));
 sg13g2_buf_1 _21204_ (.A(net816),
    .X(_12099_));
 sg13g2_buf_1 _21205_ (.A(_12095_),
    .X(_12100_));
 sg13g2_buf_1 _21206_ (.A(net815),
    .X(_12101_));
 sg13g2_nand2_1 _21207_ (.Y(_12102_),
    .A(_11352_),
    .B(_11350_));
 sg13g2_nand2b_1 _21208_ (.Y(_12103_),
    .B(_12095_),
    .A_N(_11471_));
 sg13g2_o21ai_1 _21209_ (.B1(_12103_),
    .Y(_12104_),
    .A1(net468),
    .A2(_12102_));
 sg13g2_nor2_1 _21210_ (.A(net815),
    .B(_11471_),
    .Y(_12105_));
 sg13g2_nor3_1 _21211_ (.A(net470),
    .B(_12102_),
    .C(_12105_),
    .Y(_12106_));
 sg13g2_a21oi_1 _21212_ (.A1(net470),
    .A2(_12104_),
    .Y(_12107_),
    .B1(_12106_));
 sg13g2_nand2_1 _21213_ (.Y(_12108_),
    .A(net469),
    .B(_12107_));
 sg13g2_inv_2 _21214_ (.Y(_12109_),
    .A(net825));
 sg13g2_a21oi_1 _21215_ (.A1(_12109_),
    .A2(_12103_),
    .Y(_12110_),
    .B1(_12096_));
 sg13g2_nor2_1 _21216_ (.A(net837),
    .B(_12110_),
    .Y(_12111_));
 sg13g2_nand2_1 _21217_ (.Y(_12112_),
    .A(net815),
    .B(_11471_));
 sg13g2_o21ai_1 _21218_ (.B1(net825),
    .Y(_12113_),
    .A1(net815),
    .A2(_11471_));
 sg13g2_a21oi_1 _21219_ (.A1(_12112_),
    .A2(_12113_),
    .Y(_12114_),
    .B1(_12102_));
 sg13g2_or3_1 _21220_ (.A(net469),
    .B(_12111_),
    .C(_12114_),
    .X(_12115_));
 sg13g2_nor2_2 _21221_ (.A(_11737_),
    .B(net468),
    .Y(_12116_));
 sg13g2_nand2b_1 _21222_ (.Y(_12117_),
    .B(_12116_),
    .A_N(net816));
 sg13g2_inv_2 _21223_ (.Y(_12118_),
    .A(net815));
 sg13g2_nor2_1 _21224_ (.A(_12109_),
    .B(_12118_),
    .Y(_12119_));
 sg13g2_nand3_1 _21225_ (.B(_11351_),
    .C(_12119_),
    .A(net816),
    .Y(_12120_));
 sg13g2_a21oi_1 _21226_ (.A1(_12117_),
    .A2(_12120_),
    .Y(_12121_),
    .B1(net836));
 sg13g2_a221oi_1 _21227_ (.B2(_12115_),
    .C1(_12121_),
    .B1(_12108_),
    .A1(_11731_),
    .Y(_12122_),
    .A2(_12096_));
 sg13g2_buf_1 _21228_ (.A(_12122_),
    .X(_12123_));
 sg13g2_buf_1 _21229_ (.A(_00010_),
    .X(_12124_));
 sg13g2_buf_1 _21230_ (.A(_12124_),
    .X(_12125_));
 sg13g2_nor2b_1 _21231_ (.A(net827),
    .B_N(net814),
    .Y(_12126_));
 sg13g2_o21ai_1 _21232_ (.B1(net821),
    .Y(_12127_),
    .A1(net229),
    .A2(_12126_));
 sg13g2_nand3_1 _21233_ (.B(net814),
    .C(net821),
    .A(net229),
    .Y(_12128_));
 sg13g2_nor2_1 _21234_ (.A(_12123_),
    .B(_12128_),
    .Y(_12129_));
 sg13g2_a21oi_1 _21235_ (.A1(_12123_),
    .A2(_12127_),
    .Y(_12130_),
    .B1(_12129_));
 sg13g2_nor3_1 _21236_ (.A(net228),
    .B(_11834_),
    .C(_12123_),
    .Y(_12131_));
 sg13g2_nor3_1 _21237_ (.A(net229),
    .B(net814),
    .C(net821),
    .Y(_12132_));
 sg13g2_o21ai_1 _21238_ (.B1(_11400_),
    .Y(_12133_),
    .A1(_12131_),
    .A2(_12132_));
 sg13g2_xnor2_1 _21239_ (.Y(_12134_),
    .A(_11352_),
    .B(net816));
 sg13g2_xnor2_1 _21240_ (.Y(_12135_),
    .A(_11720_),
    .B(_12134_));
 sg13g2_xnor2_1 _21241_ (.Y(_12136_),
    .A(net467),
    .B(_12135_));
 sg13g2_buf_2 _21242_ (.A(_12136_),
    .X(_12137_));
 sg13g2_a21oi_1 _21243_ (.A1(_12130_),
    .A2(_12133_),
    .Y(_12138_),
    .B1(_12137_));
 sg13g2_nor2_1 _21244_ (.A(net228),
    .B(net814),
    .Y(_12139_));
 sg13g2_nand2_1 _21245_ (.Y(_12140_),
    .A(net477),
    .B(_12137_));
 sg13g2_nand2_1 _21246_ (.Y(_12141_),
    .A(net814),
    .B(_12140_));
 sg13g2_a22oi_1 _21247_ (.Y(_12142_),
    .B1(_12141_),
    .B2(net827),
    .A2(_12139_),
    .A1(_12137_));
 sg13g2_nand2_1 _21248_ (.Y(_12143_),
    .A(net228),
    .B(net814));
 sg13g2_o21ai_1 _21249_ (.B1(_12143_),
    .Y(_12144_),
    .A1(net827),
    .A2(_12139_));
 sg13g2_a221oi_1 _21250_ (.B2(_12137_),
    .C1(_12123_),
    .B1(_12144_),
    .A1(net821),
    .Y(_12145_),
    .A2(_12126_));
 sg13g2_a21oi_1 _21251_ (.A1(_12123_),
    .A2(_12142_),
    .Y(_12146_),
    .B1(_12145_));
 sg13g2_nor2_1 _21252_ (.A(net467),
    .B(net833),
    .Y(_12147_));
 sg13g2_nand2_1 _21253_ (.Y(_12148_),
    .A(net825),
    .B(net815));
 sg13g2_buf_1 _21254_ (.A(_12148_),
    .X(_12149_));
 sg13g2_xor2_1 _21255_ (.B(_12095_),
    .A(_11718_),
    .X(_12150_));
 sg13g2_nand2_1 _21256_ (.Y(_12151_),
    .A(net835),
    .B(_12150_));
 sg13g2_o21ai_1 _21257_ (.B1(_12151_),
    .Y(_12152_),
    .A1(net835),
    .A2(_12149_));
 sg13g2_a22oi_1 _21258_ (.Y(_12153_),
    .B1(_12152_),
    .B2(net233),
    .A2(_12147_),
    .A1(net222));
 sg13g2_buf_1 _21259_ (.A(net469),
    .X(_12154_));
 sg13g2_nor2b_1 _21260_ (.A(_12153_),
    .B_N(net221),
    .Y(_12155_));
 sg13g2_nor3_1 _21261_ (.A(net221),
    .B(_12102_),
    .C(_12149_),
    .Y(_12156_));
 sg13g2_nor2b_1 _21262_ (.A(_10992_),
    .B_N(_05748_),
    .Y(_12157_));
 sg13g2_buf_2 _21263_ (.A(_12157_),
    .X(_12158_));
 sg13g2_nand2_1 _21264_ (.Y(_12159_),
    .A(net327),
    .B(_12158_));
 sg13g2_buf_2 _21265_ (.A(_12159_),
    .X(_12160_));
 sg13g2_nand2_1 _21266_ (.Y(_12161_),
    .A(net1194),
    .B(_12160_));
 sg13g2_nand3_1 _21267_ (.B(_11834_),
    .C(_12139_),
    .A(net827),
    .Y(_12162_));
 sg13g2_buf_2 _21268_ (.A(\grid.cell_27_0.s ),
    .X(_12163_));
 sg13g2_xnor2_1 _21269_ (.Y(_12164_),
    .A(_12163_),
    .B(_11716_));
 sg13g2_xnor2_1 _21270_ (.Y(_12165_),
    .A(_11400_),
    .B(_12164_));
 sg13g2_xnor2_1 _21271_ (.Y(_12166_),
    .A(_12137_),
    .B(_12165_));
 sg13g2_inv_1 _21272_ (.Y(_12167_),
    .A(_11754_));
 sg13g2_o21ai_1 _21273_ (.B1(_12167_),
    .Y(_12168_),
    .A1(net170),
    .A2(_12166_));
 sg13g2_o21ai_1 _21274_ (.B1(_12168_),
    .Y(_12169_),
    .A1(_12137_),
    .A2(_12162_));
 sg13g2_nor4_1 _21275_ (.A(_12155_),
    .B(_12156_),
    .C(_12161_),
    .D(_12169_),
    .Y(_12170_));
 sg13g2_nand2b_1 _21276_ (.Y(_12171_),
    .B(_12170_),
    .A_N(_12146_));
 sg13g2_nand3_1 _21277_ (.B(net110),
    .C(_12160_),
    .A(net824),
    .Y(_12172_));
 sg13g2_o21ai_1 _21278_ (.B1(_12172_),
    .Y(_12173_),
    .A1(net50),
    .A2(_12160_));
 sg13g2_nand2_1 _21279_ (.Y(_12174_),
    .A(net312),
    .B(_12173_));
 sg13g2_o21ai_1 _21280_ (.B1(_12174_),
    .Y(_00429_),
    .A1(_12138_),
    .A2(_12171_));
 sg13g2_buf_8 _21281_ (.A(\grid.cell_27_1.se ),
    .X(_12175_));
 sg13g2_inv_2 _21282_ (.Y(_12176_),
    .A(_12175_));
 sg13g2_nand2_1 _21283_ (.Y(_12177_),
    .A(_12176_),
    .B(net833));
 sg13g2_nor3_1 _21284_ (.A(net138),
    .B(net227),
    .C(_12177_),
    .Y(_12178_));
 sg13g2_buf_1 _21285_ (.A(_12175_),
    .X(_12179_));
 sg13g2_buf_1 _21286_ (.A(net813),
    .X(_12180_));
 sg13g2_or3_1 _21287_ (.A(net221),
    .B(net475),
    .C(net466),
    .X(_12181_));
 sg13g2_nand2_1 _21288_ (.Y(_12182_),
    .A(net816),
    .B(net813));
 sg13g2_inv_1 _21289_ (.Y(_12183_),
    .A(_12182_));
 sg13g2_nand3_1 _21290_ (.B(net475),
    .C(_12183_),
    .A(net232),
    .Y(_12184_));
 sg13g2_a21oi_1 _21291_ (.A1(_12181_),
    .A2(_12184_),
    .Y(_12185_),
    .B1(_11375_));
 sg13g2_nor2_1 _21292_ (.A(_12176_),
    .B(net833),
    .Y(_12186_));
 sg13g2_o21ai_1 _21293_ (.B1(_12177_),
    .Y(_12187_),
    .A1(net476),
    .A2(_12186_));
 sg13g2_nand2_1 _21294_ (.Y(_12188_),
    .A(net466),
    .B(_11472_));
 sg13g2_o21ai_1 _21295_ (.B1(net823),
    .Y(_12189_),
    .A1(net813),
    .A2(_11472_));
 sg13g2_nand2_1 _21296_ (.Y(_12190_),
    .A(_11352_),
    .B(net834));
 sg13g2_a21oi_1 _21297_ (.A1(_12188_),
    .A2(_12189_),
    .Y(_12191_),
    .B1(_12190_));
 sg13g2_a21oi_1 _21298_ (.A1(_11446_),
    .A2(_12187_),
    .Y(_12192_),
    .B1(_12191_));
 sg13g2_nand2b_1 _21299_ (.Y(_12193_),
    .B(net813),
    .A_N(_11471_));
 sg13g2_o21ai_1 _21300_ (.B1(_12193_),
    .Y(_12194_),
    .A1(net466),
    .A2(_12190_));
 sg13g2_nor2_1 _21301_ (.A(net813),
    .B(_11471_),
    .Y(_12195_));
 sg13g2_nor3_1 _21302_ (.A(net823),
    .B(_12190_),
    .C(_12195_),
    .Y(_12196_));
 sg13g2_a21oi_1 _21303_ (.A1(net476),
    .A2(_12194_),
    .Y(_12197_),
    .B1(_12196_));
 sg13g2_nand2b_1 _21304_ (.Y(_12198_),
    .B(net221),
    .A_N(_12197_));
 sg13g2_o21ai_1 _21305_ (.B1(_12198_),
    .Y(_12199_),
    .A1(net221),
    .A2(_12192_));
 sg13g2_nor3_1 _21306_ (.A(_12178_),
    .B(_12185_),
    .C(_12199_),
    .Y(_12200_));
 sg13g2_nand2_1 _21307_ (.Y(_12201_),
    .A(_11400_),
    .B(net814));
 sg13g2_xnor2_1 _21308_ (.Y(_12202_),
    .A(_12176_),
    .B(_11783_));
 sg13g2_xor2_1 _21309_ (.B(_12202_),
    .A(_12134_),
    .X(_12203_));
 sg13g2_xnor2_1 _21310_ (.Y(_12204_),
    .A(net824),
    .B(_12203_));
 sg13g2_nand2b_1 _21311_ (.Y(_12205_),
    .B(net827),
    .A_N(_12125_));
 sg13g2_o21ai_1 _21312_ (.B1(_12205_),
    .Y(_12206_),
    .A1(net1099),
    .A2(_12203_));
 sg13g2_a21oi_1 _21313_ (.A1(_12201_),
    .A2(_12204_),
    .Y(_12207_),
    .B1(_12206_));
 sg13g2_xnor2_1 _21314_ (.Y(_12208_),
    .A(_12200_),
    .B(_12207_));
 sg13g2_xnor2_1 _21315_ (.Y(_12209_),
    .A(_11754_),
    .B(_12163_));
 sg13g2_xnor2_1 _21316_ (.Y(_12210_),
    .A(_11715_),
    .B(_12209_));
 sg13g2_xor2_1 _21317_ (.B(_12210_),
    .A(_12203_),
    .X(_12211_));
 sg13g2_buf_1 _21318_ (.A(net466),
    .X(_12212_));
 sg13g2_nand4_1 _21319_ (.B(net232),
    .C(net475),
    .A(net486),
    .Y(_12213_),
    .D(net220));
 sg13g2_nand2_1 _21320_ (.Y(_12214_),
    .A(_11784_),
    .B(net813));
 sg13g2_xor2_1 _21321_ (.B(_12175_),
    .A(net1098),
    .X(_12215_));
 sg13g2_nand2_1 _21322_ (.Y(_12216_),
    .A(net836),
    .B(_12215_));
 sg13g2_o21ai_1 _21323_ (.B1(_12216_),
    .Y(_12217_),
    .A1(net836),
    .A2(_12214_));
 sg13g2_a22oi_1 _21324_ (.Y(_12218_),
    .B1(_12217_),
    .B2(_11416_),
    .A2(_12186_),
    .A1(net475));
 sg13g2_mux2_1 _21325_ (.A0(_12213_),
    .A1(_12218_),
    .S(net221),
    .X(_12219_));
 sg13g2_xor2_1 _21326_ (.B(net824),
    .A(_11399_),
    .X(_12220_));
 sg13g2_nor3_1 _21327_ (.A(net814),
    .B(_11725_),
    .C(_12220_),
    .Y(_12221_));
 sg13g2_nand2b_1 _21328_ (.Y(_12222_),
    .B(_12221_),
    .A_N(_12203_));
 sg13g2_nand3_1 _21329_ (.B(_12219_),
    .C(_12222_),
    .A(net116),
    .Y(_12223_));
 sg13g2_a21oi_1 _21330_ (.A1(net228),
    .A2(_12211_),
    .Y(_12224_),
    .B1(_12223_));
 sg13g2_a22oi_1 _21331_ (.Y(_12225_),
    .B1(_12208_),
    .B2(_12224_),
    .A2(net67),
    .A1(net229));
 sg13g2_o21ai_1 _21332_ (.B1(net522),
    .Y(_12226_),
    .A1(net38),
    .A2(_12160_));
 sg13g2_a21oi_1 _21333_ (.A1(_12160_),
    .A2(_12225_),
    .Y(_00430_),
    .B1(_12226_));
 sg13g2_nand3_1 _21334_ (.B(net108),
    .C(_12158_),
    .A(net1002),
    .Y(_12227_));
 sg13g2_buf_1 _21335_ (.A(_12227_),
    .X(_12228_));
 sg13g2_buf_1 _21336_ (.A(\grid.cell_27_2.se ),
    .X(_12229_));
 sg13g2_nand2_1 _21337_ (.Y(_12230_),
    .A(net822),
    .B(net1094));
 sg13g2_xor2_1 _21338_ (.B(net1094),
    .A(net822),
    .X(_12231_));
 sg13g2_nand2_1 _21339_ (.Y(_12232_),
    .A(_11413_),
    .B(_12231_));
 sg13g2_o21ai_1 _21340_ (.B1(_12232_),
    .Y(_12233_),
    .A1(net485),
    .A2(_12230_));
 sg13g2_nand2_1 _21341_ (.Y(_12234_),
    .A(net231),
    .B(_12233_));
 sg13g2_o21ai_1 _21342_ (.B1(_12234_),
    .Y(_12235_),
    .A1(_11536_),
    .A2(_12230_));
 sg13g2_nand2_1 _21343_ (.Y(_12236_),
    .A(_11414_),
    .B(net483));
 sg13g2_nor2_1 _21344_ (.A(net220),
    .B(_12236_),
    .Y(_12237_));
 sg13g2_inv_1 _21345_ (.Y(_12238_),
    .A(_12230_));
 sg13g2_buf_1 _21346_ (.A(_00009_),
    .X(_12239_));
 sg13g2_buf_1 _21347_ (.A(_12239_),
    .X(_12240_));
 sg13g2_inv_1 _21348_ (.Y(_12241_),
    .A(net812));
 sg13g2_xnor2_1 _21349_ (.Y(_12242_),
    .A(net1094),
    .B(_11837_));
 sg13g2_xnor2_1 _21350_ (.Y(_12243_),
    .A(_11413_),
    .B(_12175_));
 sg13g2_xnor2_1 _21351_ (.Y(_12244_),
    .A(_12242_),
    .B(_12243_));
 sg13g2_xnor2_1 _21352_ (.Y(_12245_),
    .A(net836),
    .B(_11728_));
 sg13g2_and4_1 _21353_ (.A(_12241_),
    .B(_11834_),
    .C(_12244_),
    .D(_12245_),
    .X(_12246_));
 sg13g2_a221oi_1 _21354_ (.B2(_12238_),
    .C1(_12246_),
    .B1(_12237_),
    .A1(net220),
    .Y(_12247_),
    .A2(_12235_));
 sg13g2_xnor2_1 _21355_ (.Y(_12248_),
    .A(_11743_),
    .B(_12244_));
 sg13g2_nand2b_1 _21356_ (.Y(_12249_),
    .B(net812),
    .A_N(_11360_));
 sg13g2_nor2b_1 _21357_ (.A(net812),
    .B_N(_11360_),
    .Y(_12250_));
 sg13g2_a221oi_1 _21358_ (.B2(_12249_),
    .C1(_12250_),
    .B1(_12248_),
    .A1(_11834_),
    .Y(_12251_),
    .A2(_12244_));
 sg13g2_buf_1 _21359_ (.A(net1094),
    .X(_12252_));
 sg13g2_nor2_1 _21360_ (.A(net822),
    .B(net811),
    .Y(_12253_));
 sg13g2_o21ai_1 _21361_ (.B1(_12232_),
    .Y(_12254_),
    .A1(net483),
    .A2(_12238_));
 sg13g2_a22oi_1 _21362_ (.Y(_12255_),
    .B1(_12254_),
    .B2(_11536_),
    .A2(_12253_),
    .A1(_12236_));
 sg13g2_o21ai_1 _21363_ (.B1(net483),
    .Y(_12256_),
    .A1(_11446_),
    .A2(_12176_));
 sg13g2_nand3_1 _21364_ (.B(_12256_),
    .C(_12253_),
    .A(net830),
    .Y(_12257_));
 sg13g2_o21ai_1 _21365_ (.B1(_12257_),
    .Y(_12258_),
    .A1(net220),
    .A2(_12255_));
 sg13g2_xor2_1 _21366_ (.B(_12258_),
    .A(_12251_),
    .X(_12259_));
 sg13g2_a21oi_1 _21367_ (.A1(_12247_),
    .A2(_12259_),
    .Y(_12260_),
    .B1(net96));
 sg13g2_xnor2_1 _21368_ (.Y(_12261_),
    .A(_12134_),
    .B(_12248_));
 sg13g2_a21oi_1 _21369_ (.A1(net68),
    .A2(_12261_),
    .Y(_12262_),
    .B1(net227));
 sg13g2_or3_1 _21370_ (.A(_12161_),
    .B(_12260_),
    .C(_12262_),
    .X(_12263_));
 sg13g2_o21ai_1 _21371_ (.B1(_12263_),
    .Y(_00431_),
    .A1(net27),
    .A2(_12228_));
 sg13g2_buf_1 _21372_ (.A(net811),
    .X(_12264_));
 sg13g2_buf_1 _21373_ (.A(\grid.cell_27_3.se ),
    .X(_12265_));
 sg13g2_buf_1 _21374_ (.A(_12265_),
    .X(_12266_));
 sg13g2_nand2_2 _21375_ (.Y(_12267_),
    .A(net820),
    .B(net810));
 sg13g2_xor2_1 _21376_ (.B(net810),
    .A(net820),
    .X(_12268_));
 sg13g2_nand2_1 _21377_ (.Y(_12269_),
    .A(net483),
    .B(_12268_));
 sg13g2_o21ai_1 _21378_ (.B1(_12269_),
    .Y(_12270_),
    .A1(_11489_),
    .A2(_12267_));
 sg13g2_nand2_1 _21379_ (.Y(_12271_),
    .A(net482),
    .B(_12270_));
 sg13g2_o21ai_1 _21380_ (.B1(_12271_),
    .Y(_12272_),
    .A1(net1101),
    .A2(_12267_));
 sg13g2_xnor2_1 _21381_ (.Y(_12273_),
    .A(net1094),
    .B(_12265_));
 sg13g2_xor2_1 _21382_ (.B(_12273_),
    .A(_11903_),
    .X(_12274_));
 sg13g2_xnor2_1 _21383_ (.Y(_12275_),
    .A(net832),
    .B(_12274_));
 sg13g2_and2_1 _21384_ (.A(_11899_),
    .B(_12275_),
    .X(_12276_));
 sg13g2_buf_2 _21385_ (.A(_00008_),
    .X(_12277_));
 sg13g2_nor2_1 _21386_ (.A(_12277_),
    .B(_11783_),
    .Y(_12278_));
 sg13g2_nor3_1 _21387_ (.A(net465),
    .B(_11527_),
    .C(_12267_),
    .Y(_12279_));
 sg13g2_a221oi_1 _21388_ (.B2(_12278_),
    .C1(_12279_),
    .B1(_12276_),
    .A1(net465),
    .Y(_12280_),
    .A2(_12272_));
 sg13g2_a22oi_1 _21389_ (.Y(_12281_),
    .B1(_12267_),
    .B2(_11591_),
    .A2(_12268_),
    .A1(_11489_));
 sg13g2_buf_1 _21390_ (.A(net810),
    .X(_12282_));
 sg13g2_a21oi_1 _21391_ (.A1(_11481_),
    .A2(net1094),
    .Y(_12283_),
    .B1(_11591_));
 sg13g2_or3_1 _21392_ (.A(net473),
    .B(net464),
    .C(_12283_),
    .X(_12284_));
 sg13g2_o21ai_1 _21393_ (.B1(_12284_),
    .Y(_12285_),
    .A1(net811),
    .A2(_12281_));
 sg13g2_buf_1 _21394_ (.A(net464),
    .X(_12286_));
 sg13g2_nor3_1 _21395_ (.A(net811),
    .B(net473),
    .C(net219),
    .Y(_12287_));
 sg13g2_a22oi_1 _21396_ (.Y(_12288_),
    .B1(_12287_),
    .B2(_11527_),
    .A2(_12285_),
    .A1(net1101));
 sg13g2_nand2_1 _21397_ (.Y(_12289_),
    .A(_11446_),
    .B(_12277_));
 sg13g2_xor2_1 _21398_ (.B(_12275_),
    .A(_11785_),
    .X(_12290_));
 sg13g2_nor2_1 _21399_ (.A(_11446_),
    .B(_12277_),
    .Y(_12291_));
 sg13g2_a221oi_1 _21400_ (.B2(_12290_),
    .C1(_12291_),
    .B1(_12289_),
    .A1(_11899_),
    .Y(_12292_),
    .A2(_12275_));
 sg13g2_xnor2_1 _21401_ (.Y(_12293_),
    .A(_12288_),
    .B(_12292_));
 sg13g2_a21oi_1 _21402_ (.A1(_12280_),
    .A2(_12293_),
    .Y(_12294_),
    .B1(net96));
 sg13g2_xor2_1 _21403_ (.B(_12275_),
    .A(_12202_),
    .X(_12295_));
 sg13g2_a21oi_1 _21404_ (.A1(net68),
    .A2(_12295_),
    .Y(_12296_),
    .B1(net226));
 sg13g2_or3_1 _21405_ (.A(_12161_),
    .B(_12294_),
    .C(_12296_),
    .X(_12297_));
 sg13g2_o21ai_1 _21406_ (.B1(_12297_),
    .Y(_00432_),
    .A1(net32),
    .A2(_12228_));
 sg13g2_buf_1 _21407_ (.A(net47),
    .X(_12298_));
 sg13g2_xnor2_1 _21408_ (.Y(_12299_),
    .A(_11522_),
    .B(net810));
 sg13g2_buf_2 _21409_ (.A(\grid.cell_27_4.se ),
    .X(_12300_));
 sg13g2_inv_2 _21410_ (.Y(_12301_),
    .A(_12300_));
 sg13g2_xnor2_1 _21411_ (.Y(_12302_),
    .A(_12301_),
    .B(_11917_));
 sg13g2_xnor2_1 _21412_ (.Y(_12303_),
    .A(_12299_),
    .B(_12302_));
 sg13g2_xor2_1 _21413_ (.B(_12303_),
    .A(_11853_),
    .X(_12304_));
 sg13g2_buf_1 _21414_ (.A(_00061_),
    .X(_12305_));
 sg13g2_nand2b_1 _21415_ (.Y(_12306_),
    .B(net1093),
    .A_N(net483));
 sg13g2_nor2b_1 _21416_ (.A(net1093),
    .B_N(net231),
    .Y(_12307_));
 sg13g2_a221oi_1 _21417_ (.B2(_12306_),
    .C1(_12307_),
    .B1(_12304_),
    .A1(_11938_),
    .Y(_12308_),
    .A2(_12303_));
 sg13g2_buf_1 _21418_ (.A(_12300_),
    .X(_12309_));
 sg13g2_nand2_1 _21419_ (.Y(_12310_),
    .A(net819),
    .B(net809));
 sg13g2_xor2_1 _21420_ (.B(_12300_),
    .A(net1096),
    .X(_12311_));
 sg13g2_and2_1 _21421_ (.A(_11522_),
    .B(_12311_),
    .X(_12312_));
 sg13g2_a21oi_1 _21422_ (.A1(_11593_),
    .A2(_12310_),
    .Y(_12313_),
    .B1(_12312_));
 sg13g2_inv_2 _21423_ (.Y(_12314_),
    .A(net810));
 sg13g2_o21ai_1 _21424_ (.B1(net829),
    .Y(_12315_),
    .A1(_11591_),
    .A2(_12314_));
 sg13g2_nand3_1 _21425_ (.B(_12301_),
    .C(_12315_),
    .A(_11921_),
    .Y(_12316_));
 sg13g2_o21ai_1 _21426_ (.B1(_12316_),
    .Y(_12317_),
    .A1(net464),
    .A2(_12313_));
 sg13g2_buf_1 _21427_ (.A(_12309_),
    .X(_12318_));
 sg13g2_nor3_1 _21428_ (.A(_11950_),
    .B(_12318_),
    .C(_11580_),
    .Y(_12319_));
 sg13g2_a22oi_1 _21429_ (.Y(_12320_),
    .B1(_12319_),
    .B2(_12314_),
    .A2(_12317_),
    .A1(_11624_));
 sg13g2_xnor2_1 _21430_ (.Y(_12321_),
    .A(_12308_),
    .B(_12320_));
 sg13g2_nor2_1 _21431_ (.A(net482),
    .B(_12310_),
    .Y(_12322_));
 sg13g2_o21ai_1 _21432_ (.B1(_11597_),
    .Y(_12323_),
    .A1(_12312_),
    .A2(_12322_));
 sg13g2_o21ai_1 _21433_ (.B1(_12323_),
    .Y(_12324_),
    .A1(_11624_),
    .A2(_12310_));
 sg13g2_nor2b_1 _21434_ (.A(net1093),
    .B_N(_11837_),
    .Y(_12325_));
 sg13g2_and2_1 _21435_ (.A(_11938_),
    .B(_12303_),
    .X(_12326_));
 sg13g2_nor3_1 _21436_ (.A(net219),
    .B(_11577_),
    .C(_12310_),
    .Y(_12327_));
 sg13g2_a221oi_1 _21437_ (.B2(_12326_),
    .C1(_12327_),
    .B1(_12325_),
    .A1(net219),
    .Y(_12328_),
    .A2(_12324_));
 sg13g2_a21oi_1 _21438_ (.A1(_12321_),
    .A2(_12328_),
    .Y(_12329_),
    .B1(net96));
 sg13g2_xor2_1 _21439_ (.B(_12303_),
    .A(_12242_),
    .X(_12330_));
 sg13g2_a21oi_1 _21440_ (.A1(net68),
    .A2(_12330_),
    .Y(_12331_),
    .B1(_11886_));
 sg13g2_or3_1 _21441_ (.A(_12161_),
    .B(_12329_),
    .C(_12331_),
    .X(_12332_));
 sg13g2_o21ai_1 _21442_ (.B1(_12332_),
    .Y(_00433_),
    .A1(net29),
    .A2(_12228_));
 sg13g2_or2_1 _21443_ (.X(_12333_),
    .B(_12160_),
    .A(_05002_));
 sg13g2_buf_1 _21444_ (.A(\grid.cell_27_5.se ),
    .X(_12334_));
 sg13g2_xnor2_1 _21445_ (.Y(_12335_),
    .A(_12300_),
    .B(net1092));
 sg13g2_xnor2_1 _21446_ (.Y(_12336_),
    .A(_11616_),
    .B(_12335_));
 sg13g2_xnor2_1 _21447_ (.Y(_12337_),
    .A(net223),
    .B(_12336_));
 sg13g2_nor2_1 _21448_ (.A(_11984_),
    .B(_12337_),
    .Y(_12338_));
 sg13g2_xor2_1 _21449_ (.B(net1092),
    .A(_11966_),
    .X(_12339_));
 sg13g2_buf_2 _21450_ (.A(_12339_),
    .X(_12340_));
 sg13g2_buf_1 _21451_ (.A(net1092),
    .X(_12341_));
 sg13g2_a21oi_1 _21452_ (.A1(net818),
    .A2(net808),
    .Y(_12342_),
    .B1(_11613_));
 sg13g2_a21oi_1 _21453_ (.A1(_11576_),
    .A2(_12340_),
    .Y(_12343_),
    .B1(_12342_));
 sg13g2_nand2_1 _21454_ (.Y(_12344_),
    .A(_11576_),
    .B(net809));
 sg13g2_or2_1 _21455_ (.X(_12345_),
    .B(net1092),
    .A(net818));
 sg13g2_a21o_1 _21456_ (.A2(_12344_),
    .A1(net828),
    .B1(_12345_),
    .X(_12346_));
 sg13g2_o21ai_1 _21457_ (.B1(_12346_),
    .Y(_12347_),
    .A1(net809),
    .A2(_12343_));
 sg13g2_nor2_1 _21458_ (.A(net809),
    .B(_12345_),
    .Y(_12348_));
 sg13g2_a22oi_1 _21459_ (.Y(_12349_),
    .B1(_12348_),
    .B2(_11615_),
    .A2(_12347_),
    .A1(_11662_));
 sg13g2_and2_1 _21460_ (.A(net818),
    .B(net1092),
    .X(_12350_));
 sg13g2_buf_1 _21461_ (.A(_12350_),
    .X(_12351_));
 sg13g2_mux2_1 _21462_ (.A0(_12340_),
    .A1(_12351_),
    .S(_11592_),
    .X(_12352_));
 sg13g2_a22oi_1 _21463_ (.Y(_12353_),
    .B1(_12352_),
    .B2(net479),
    .A2(_12351_),
    .A1(_11668_));
 sg13g2_nand2b_1 _21464_ (.Y(_12354_),
    .B(net463),
    .A_N(_12353_));
 sg13g2_nand4_1 _21465_ (.B(_12301_),
    .C(net479),
    .A(net480),
    .Y(_12355_),
    .D(_12351_));
 sg13g2_nand3_1 _21466_ (.B(_12354_),
    .C(_12355_),
    .A(_12349_),
    .Y(_12356_));
 sg13g2_buf_2 _21467_ (.A(_00093_),
    .X(_12357_));
 sg13g2_xnor2_1 _21468_ (.Y(_12358_),
    .A(_12300_),
    .B(_11613_));
 sg13g2_xnor2_1 _21469_ (.Y(_12359_),
    .A(_12340_),
    .B(_12358_));
 sg13g2_xnor2_1 _21470_ (.Y(_12360_),
    .A(_11933_),
    .B(_12359_));
 sg13g2_nand2_1 _21471_ (.Y(_12361_),
    .A(_11531_),
    .B(_12360_));
 sg13g2_nor2_1 _21472_ (.A(_11531_),
    .B(_12360_),
    .Y(_12362_));
 sg13g2_a21oi_1 _21473_ (.A1(_12357_),
    .A2(_12361_),
    .Y(_12363_),
    .B1(_12362_));
 sg13g2_or3_1 _21474_ (.A(_12357_),
    .B(_12349_),
    .C(_12362_),
    .X(_12364_));
 sg13g2_o21ai_1 _21475_ (.B1(_12364_),
    .Y(_12365_),
    .A1(_12356_),
    .A2(_12363_));
 sg13g2_nor2b_1 _21476_ (.A(_12338_),
    .B_N(_12365_),
    .Y(_12366_));
 sg13g2_o21ai_1 _21477_ (.B1(_12338_),
    .Y(_12367_),
    .A1(_12357_),
    .A2(_12362_));
 sg13g2_a21oi_1 _21478_ (.A1(_12361_),
    .A2(_12367_),
    .Y(_12368_),
    .B1(_12349_));
 sg13g2_nand2b_1 _21479_ (.Y(_12369_),
    .B(net83),
    .A_N(_12368_));
 sg13g2_xnor2_1 _21480_ (.Y(_12370_),
    .A(_12299_),
    .B(_12360_));
 sg13g2_nand2_1 _21481_ (.Y(_12371_),
    .A(net126),
    .B(_12370_));
 sg13g2_a22oi_1 _21482_ (.Y(_12372_),
    .B1(_12371_),
    .B2(_11921_),
    .A2(_12158_),
    .A1(net108));
 sg13g2_o21ai_1 _21483_ (.B1(_12372_),
    .Y(_12373_),
    .A1(_12366_),
    .A2(_12369_));
 sg13g2_a21oi_1 _21484_ (.A1(_12333_),
    .A2(_12373_),
    .Y(_00434_),
    .B1(net523));
 sg13g2_buf_1 _21485_ (.A(_00155_),
    .X(_12374_));
 sg13g2_nor2_1 _21486_ (.A(net1091),
    .B(_12149_),
    .Y(_12375_));
 sg13g2_buf_1 _21487_ (.A(net808),
    .X(_12376_));
 sg13g2_nand3_1 _21488_ (.B(net462),
    .C(_12149_),
    .A(net1091),
    .Y(_12377_));
 sg13g2_nor2b_1 _21489_ (.A(_12375_),
    .B_N(_12377_),
    .Y(_12378_));
 sg13g2_xor2_1 _21490_ (.B(net462),
    .A(net1091),
    .X(_12379_));
 sg13g2_nand2b_1 _21491_ (.Y(_12380_),
    .B(_12379_),
    .A_N(_12116_));
 sg13g2_a21oi_1 _21492_ (.A1(_12378_),
    .A2(_12380_),
    .Y(_12381_),
    .B1(net478));
 sg13g2_inv_2 _21493_ (.Y(_12382_),
    .A(net1092));
 sg13g2_nand2_1 _21494_ (.Y(_12383_),
    .A(_12382_),
    .B(_12116_));
 sg13g2_nor2_1 _21495_ (.A(net462),
    .B(_12119_),
    .Y(_12384_));
 sg13g2_o21ai_1 _21496_ (.B1(net1091),
    .Y(_12385_),
    .A1(_12116_),
    .A2(_12384_));
 sg13g2_a21oi_1 _21497_ (.A1(_12383_),
    .A2(_12385_),
    .Y(_12386_),
    .B1(net233));
 sg13g2_buf_1 _21498_ (.A(net462),
    .X(_12387_));
 sg13g2_nand3_1 _21499_ (.B(_11363_),
    .C(_12119_),
    .A(net218),
    .Y(_12388_));
 sg13g2_a21oi_1 _21500_ (.A1(_12383_),
    .A2(_12388_),
    .Y(_12389_),
    .B1(net230));
 sg13g2_nor3_1 _21501_ (.A(_12374_),
    .B(_12382_),
    .C(_12149_),
    .Y(_12390_));
 sg13g2_nor4_1 _21502_ (.A(_12381_),
    .B(_12386_),
    .C(_12389_),
    .D(_12390_),
    .Y(_12391_));
 sg13g2_buf_2 _21503_ (.A(_00125_),
    .X(_12392_));
 sg13g2_xnor2_1 _21504_ (.Y(_12393_),
    .A(net1092),
    .B(_12095_));
 sg13g2_xnor2_1 _21505_ (.Y(_12394_),
    .A(_11720_),
    .B(_12393_));
 sg13g2_xnor2_1 _21506_ (.Y(_12395_),
    .A(net828),
    .B(_12394_));
 sg13g2_xnor2_1 _21507_ (.Y(_12396_),
    .A(net472),
    .B(_12395_));
 sg13g2_a21oi_1 _21508_ (.A1(_12392_),
    .A2(net481),
    .Y(_12397_),
    .B1(_12396_));
 sg13g2_nand2b_1 _21509_ (.Y(_12398_),
    .B(_12395_),
    .A_N(net1095));
 sg13g2_o21ai_1 _21510_ (.B1(_12398_),
    .Y(_12399_),
    .A1(_12392_),
    .A2(net481));
 sg13g2_nor2_1 _21511_ (.A(_12397_),
    .B(_12399_),
    .Y(_12400_));
 sg13g2_xnor2_1 _21512_ (.Y(_12401_),
    .A(_12391_),
    .B(_12400_));
 sg13g2_nand2_1 _21513_ (.Y(_12402_),
    .A(net479),
    .B(_12150_));
 sg13g2_o21ai_1 _21514_ (.B1(_12402_),
    .Y(_12403_),
    .A1(net230),
    .A2(_12149_));
 sg13g2_a21o_1 _21515_ (.A2(_12403_),
    .A1(net233),
    .B1(_12375_),
    .X(_12404_));
 sg13g2_nor3_1 _21516_ (.A(net218),
    .B(net467),
    .C(_11739_),
    .Y(_12405_));
 sg13g2_nor3_1 _21517_ (.A(_12392_),
    .B(_11917_),
    .C(_12398_),
    .Y(_12406_));
 sg13g2_a221oi_1 _21518_ (.B2(net230),
    .C1(_12406_),
    .B1(_12405_),
    .A1(net218),
    .Y(_12407_),
    .A2(_12404_));
 sg13g2_xnor2_1 _21519_ (.Y(_12408_),
    .A(_12302_),
    .B(_12395_));
 sg13g2_nand2_1 _21520_ (.Y(_12409_),
    .A(net223),
    .B(_12408_));
 sg13g2_nand4_1 _21521_ (.B(_12401_),
    .C(_12407_),
    .A(net82),
    .Y(_12410_),
    .D(_12409_));
 sg13g2_a22oi_1 _21522_ (.Y(_12411_),
    .B1(net25),
    .B2(_12158_),
    .A2(net72),
    .A1(net224));
 sg13g2_a221oi_1 _21523_ (.B2(_12411_),
    .C1(net533),
    .B1(_12410_),
    .A1(net24),
    .Y(_00435_),
    .A2(_12158_));
 sg13g2_nand2_1 _21524_ (.Y(_12412_),
    .A(net1092),
    .B(_12095_));
 sg13g2_buf_2 _21525_ (.A(_12412_),
    .X(_12413_));
 sg13g2_o21ai_1 _21526_ (.B1(net471),
    .Y(_12414_),
    .A1(net808),
    .A2(net468));
 sg13g2_nand2_1 _21527_ (.Y(_12415_),
    .A(_12413_),
    .B(_12414_));
 sg13g2_nand3b_1 _21528_ (.B(net233),
    .C(_12415_),
    .Y(_12416_),
    .A_N(net1091));
 sg13g2_nor2_1 _21529_ (.A(net471),
    .B(net462),
    .Y(_12417_));
 sg13g2_mux2_1 _21530_ (.A0(net808),
    .A1(_12413_),
    .S(_11989_),
    .X(_12418_));
 sg13g2_a22oi_1 _21531_ (.Y(_12419_),
    .B1(_12418_),
    .B2(_11363_),
    .A2(_12417_),
    .A1(net468));
 sg13g2_nand2b_1 _21532_ (.Y(_12420_),
    .B(net1091),
    .A_N(_12419_));
 sg13g2_nand3_1 _21533_ (.B(_12416_),
    .C(_12420_),
    .A(net230),
    .Y(_12421_));
 sg13g2_nand3_1 _21534_ (.B(_12382_),
    .C(net467),
    .A(net223),
    .Y(_12422_));
 sg13g2_buf_1 _21535_ (.A(net468),
    .X(_12423_));
 sg13g2_nand3_1 _21536_ (.B(net217),
    .C(_12351_),
    .A(net233),
    .Y(_12424_));
 sg13g2_nand3b_1 _21537_ (.B(_12422_),
    .C(_12424_),
    .Y(_12425_),
    .A_N(_11686_));
 sg13g2_nor2_1 _21538_ (.A(net1091),
    .B(_12413_),
    .Y(_12426_));
 sg13g2_nand3_1 _21539_ (.B(_12413_),
    .C(_12414_),
    .A(net1091),
    .Y(_12427_));
 sg13g2_a21oi_1 _21540_ (.A1(_12422_),
    .A2(_12427_),
    .Y(_12428_),
    .B1(_11364_));
 sg13g2_a221oi_1 _21541_ (.B2(net224),
    .C1(_12428_),
    .B1(_12426_),
    .A1(_12421_),
    .Y(_12429_),
    .A2(_12425_));
 sg13g2_xor2_1 _21542_ (.B(_12393_),
    .A(_11968_),
    .X(_12430_));
 sg13g2_xnor2_1 _21543_ (.Y(_12431_),
    .A(_11351_),
    .B(_12430_));
 sg13g2_xnor2_1 _21544_ (.Y(_12432_),
    .A(_12167_),
    .B(_12431_));
 sg13g2_inv_1 _21545_ (.Y(_12433_),
    .A(_12431_));
 sg13g2_o21ai_1 _21546_ (.B1(_12205_),
    .Y(_12434_),
    .A1(_11725_),
    .A2(_12433_));
 sg13g2_a21oi_1 _21547_ (.A1(_12201_),
    .A2(_12432_),
    .Y(_12435_),
    .B1(_12434_));
 sg13g2_xnor2_1 _21548_ (.Y(_12436_),
    .A(_12429_),
    .B(_12435_));
 sg13g2_nand2b_1 _21549_ (.Y(_12437_),
    .B(net230),
    .A_N(_12393_));
 sg13g2_o21ai_1 _21550_ (.B1(_12437_),
    .Y(_12438_),
    .A1(net230),
    .A2(_12413_));
 sg13g2_a21oi_1 _21551_ (.A1(net233),
    .A2(_12438_),
    .Y(_12439_),
    .B1(_12426_));
 sg13g2_nand2b_1 _21552_ (.Y(_12440_),
    .B(net224),
    .A_N(_12439_));
 sg13g2_xnor2_1 _21553_ (.Y(_12441_),
    .A(_12210_),
    .B(_12431_));
 sg13g2_nand2_1 _21554_ (.Y(_12442_),
    .A(_12109_),
    .B(_12441_));
 sg13g2_nor2_1 _21555_ (.A(_11646_),
    .B(_12413_),
    .Y(_12443_));
 sg13g2_a221oi_1 _21556_ (.B2(net223),
    .C1(net110),
    .B1(_12443_),
    .A1(_12221_),
    .Y(_12444_),
    .A2(_12431_));
 sg13g2_nand4_1 _21557_ (.B(_12440_),
    .C(_12442_),
    .A(_12436_),
    .Y(_12445_),
    .D(_12444_));
 sg13g2_a22oi_1 _21558_ (.Y(_12446_),
    .B1(net76),
    .B2(_12158_),
    .A2(net72),
    .A1(net222));
 sg13g2_a221oi_1 _21559_ (.B2(_12446_),
    .C1(net533),
    .B1(_12445_),
    .A1(_06471_),
    .Y(_00436_),
    .A2(_12158_));
 sg13g2_or2_1 _21560_ (.X(_12447_),
    .B(net159),
    .A(net177));
 sg13g2_buf_2 _21561_ (.A(_12447_),
    .X(_12448_));
 sg13g2_or3_1 _21562_ (.A(_07600_),
    .B(_02021_),
    .C(_12448_),
    .X(_12449_));
 sg13g2_buf_1 _21563_ (.A(_12449_),
    .X(_12450_));
 sg13g2_buf_1 _21564_ (.A(_12163_),
    .X(_12451_));
 sg13g2_buf_2 _21565_ (.A(\grid.cell_28_0.se ),
    .X(_12452_));
 sg13g2_buf_1 _21566_ (.A(_12452_),
    .X(_12453_));
 sg13g2_buf_1 _21567_ (.A(net806),
    .X(_12454_));
 sg13g2_buf_1 _21568_ (.A(\grid.cell_28_0.sw ),
    .X(_12455_));
 sg13g2_buf_1 _21569_ (.A(net1090),
    .X(_12456_));
 sg13g2_buf_1 _21570_ (.A(net805),
    .X(_12457_));
 sg13g2_buf_1 _21571_ (.A(net460),
    .X(_12458_));
 sg13g2_buf_1 _21572_ (.A(net216),
    .X(_12459_));
 sg13g2_nand2_1 _21573_ (.Y(_12460_),
    .A(_11728_),
    .B(net470));
 sg13g2_nand2_1 _21574_ (.Y(_12461_),
    .A(net460),
    .B(_11834_));
 sg13g2_o21ai_1 _21575_ (.B1(_12461_),
    .Y(_12462_),
    .A1(net137),
    .A2(_12460_));
 sg13g2_nor2_1 _21576_ (.A(net216),
    .B(net821),
    .Y(_12463_));
 sg13g2_nor3_1 _21577_ (.A(net217),
    .B(_12460_),
    .C(_12463_),
    .Y(_12464_));
 sg13g2_a21o_1 _21578_ (.A2(_12462_),
    .A1(net217),
    .B1(_12464_),
    .X(_12465_));
 sg13g2_nor2_1 _21579_ (.A(net460),
    .B(_11834_),
    .Y(_12466_));
 sg13g2_a21o_1 _21580_ (.A2(_12461_),
    .A1(net467),
    .B1(_12466_),
    .X(_12467_));
 sg13g2_nand2_1 _21581_ (.Y(_12468_),
    .A(net216),
    .B(net1097));
 sg13g2_buf_1 _21582_ (.A(net805),
    .X(_12469_));
 sg13g2_o21ai_1 _21583_ (.B1(net468),
    .Y(_12470_),
    .A1(net459),
    .A2(net1097));
 sg13g2_a21oi_1 _21584_ (.A1(_12468_),
    .A2(_12470_),
    .Y(_12471_),
    .B1(_12460_));
 sg13g2_a21oi_1 _21585_ (.A1(_12109_),
    .A2(_12467_),
    .Y(_12472_),
    .B1(_12471_));
 sg13g2_buf_1 _21586_ (.A(_12452_),
    .X(_12473_));
 sg13g2_or2_1 _21587_ (.X(_12474_),
    .B(net805),
    .A(net468));
 sg13g2_buf_1 _21588_ (.A(_12474_),
    .X(_12475_));
 sg13g2_nand4_1 _21589_ (.B(net470),
    .C(net217),
    .A(net804),
    .Y(_12476_),
    .D(net216));
 sg13g2_o21ai_1 _21590_ (.B1(_12476_),
    .Y(_12477_),
    .A1(net804),
    .A2(_12475_));
 sg13g2_a22oi_1 _21591_ (.Y(_12478_),
    .B1(_12477_),
    .B2(_11744_),
    .A2(_12466_),
    .A1(_12116_));
 sg13g2_o21ai_1 _21592_ (.B1(_12478_),
    .Y(_12479_),
    .A1(net461),
    .A2(_12472_));
 sg13g2_a21oi_1 _21593_ (.A1(net461),
    .A2(_12465_),
    .Y(_12480_),
    .B1(_12479_));
 sg13g2_xnor2_1 _21594_ (.Y(_12481_),
    .A(_11716_),
    .B(_12452_));
 sg13g2_xor2_1 _21595_ (.B(_12481_),
    .A(_12150_),
    .X(_12482_));
 sg13g2_xnor2_1 _21596_ (.Y(_12483_),
    .A(net460),
    .B(_12482_));
 sg13g2_xor2_1 _21597_ (.B(_12483_),
    .A(_12099_),
    .X(_12484_));
 sg13g2_buf_1 _21598_ (.A(_00007_),
    .X(_12485_));
 sg13g2_buf_1 _21599_ (.A(_12485_),
    .X(_12486_));
 sg13g2_nand2_1 _21600_ (.Y(_12487_),
    .A(_12167_),
    .B(net803));
 sg13g2_nor2_1 _21601_ (.A(_12167_),
    .B(net803),
    .Y(_12488_));
 sg13g2_a221oi_1 _21602_ (.B2(_12487_),
    .C1(_12488_),
    .B1(_12484_),
    .A1(_12241_),
    .Y(_12489_),
    .A2(_12483_));
 sg13g2_xnor2_1 _21603_ (.Y(_12490_),
    .A(_12480_),
    .B(_12489_));
 sg13g2_buf_1 _21604_ (.A(\grid.cell_28_0.s ),
    .X(_12491_));
 sg13g2_buf_1 _21605_ (.A(_12491_),
    .X(_12492_));
 sg13g2_xor2_1 _21606_ (.B(net802),
    .A(net824),
    .X(_12493_));
 sg13g2_xor2_1 _21607_ (.B(_12493_),
    .A(_12484_),
    .X(_12494_));
 sg13g2_nor2_1 _21608_ (.A(net807),
    .B(_12494_),
    .Y(_12495_));
 sg13g2_nand2_1 _21609_ (.Y(_12496_),
    .A(_12241_),
    .B(_12483_));
 sg13g2_xor2_1 _21610_ (.B(net221),
    .A(net824),
    .X(_12497_));
 sg13g2_nor3_1 _21611_ (.A(net803),
    .B(_12496_),
    .C(_12497_),
    .Y(_12498_));
 sg13g2_inv_1 _21612_ (.Y(_12499_),
    .A(net461));
 sg13g2_nand2_1 _21613_ (.Y(_12500_),
    .A(net815),
    .B(net1090));
 sg13g2_buf_1 _21614_ (.A(_12500_),
    .X(_12501_));
 sg13g2_xor2_1 _21615_ (.B(net1090),
    .A(_12095_),
    .X(_12502_));
 sg13g2_nand2_1 _21616_ (.Y(_12503_),
    .A(net477),
    .B(_12502_));
 sg13g2_o21ai_1 _21617_ (.B1(_12503_),
    .Y(_12504_),
    .A1(net477),
    .A2(_12501_));
 sg13g2_nor2_1 _21618_ (.A(net821),
    .B(_12501_),
    .Y(_12505_));
 sg13g2_a21oi_1 _21619_ (.A1(net222),
    .A2(_12504_),
    .Y(_12506_),
    .B1(_12505_));
 sg13g2_nor2b_1 _21620_ (.A(net804),
    .B_N(net459),
    .Y(_12507_));
 sg13g2_nand3_1 _21621_ (.B(_12119_),
    .C(_12507_),
    .A(_11741_),
    .Y(_12508_));
 sg13g2_o21ai_1 _21622_ (.B1(_12508_),
    .Y(_12509_),
    .A1(_12499_),
    .A2(_12506_));
 sg13g2_nor4_1 _21623_ (.A(net107),
    .B(_12495_),
    .C(_12498_),
    .D(_12509_),
    .Y(_12510_));
 sg13g2_a22oi_1 _21624_ (.Y(_12511_),
    .B1(_12490_),
    .B2(_12510_),
    .A2(net67),
    .A1(net807));
 sg13g2_o21ai_1 _21625_ (.B1(net522),
    .Y(_12512_),
    .A1(net40),
    .A2(net55));
 sg13g2_a21oi_1 _21626_ (.A1(net55),
    .A2(_12511_),
    .Y(_00437_),
    .B1(_12512_));
 sg13g2_nor3_1 _21627_ (.A(_07600_),
    .B(net375),
    .C(_12448_),
    .Y(_12513_));
 sg13g2_buf_1 _21628_ (.A(_12513_),
    .X(_12514_));
 sg13g2_nand2_1 _21629_ (.Y(_12515_),
    .A(net42),
    .B(net54));
 sg13g2_buf_8 _21630_ (.A(\grid.cell_28_1.se ),
    .X(_12516_));
 sg13g2_buf_1 _21631_ (.A(_12516_),
    .X(_12517_));
 sg13g2_buf_1 _21632_ (.A(net801),
    .X(_12518_));
 sg13g2_nand2_1 _21633_ (.Y(_12519_),
    .A(net826),
    .B(net1098));
 sg13g2_nand2b_1 _21634_ (.Y(_12520_),
    .B(_12516_),
    .A_N(net1097));
 sg13g2_o21ai_1 _21635_ (.B1(_12520_),
    .Y(_12521_),
    .A1(net458),
    .A2(_12519_));
 sg13g2_nor2_1 _21636_ (.A(net801),
    .B(net1097),
    .Y(_12522_));
 sg13g2_nor3_1 _21637_ (.A(net466),
    .B(_12519_),
    .C(_12522_),
    .Y(_12523_));
 sg13g2_a21oi_1 _21638_ (.A1(net466),
    .A2(_12521_),
    .Y(_12524_),
    .B1(_12523_));
 sg13g2_nor2b_1 _21639_ (.A(net801),
    .B_N(net1097),
    .Y(_12525_));
 sg13g2_a21oi_1 _21640_ (.A1(_12176_),
    .A2(_12520_),
    .Y(_12526_),
    .B1(_12525_));
 sg13g2_nor2_1 _21641_ (.A(_11785_),
    .B(_12526_),
    .Y(_12527_));
 sg13g2_nand2_1 _21642_ (.Y(_12528_),
    .A(net458),
    .B(_11833_));
 sg13g2_o21ai_1 _21643_ (.B1(net813),
    .Y(_12529_),
    .A1(net801),
    .A2(net1097));
 sg13g2_a21oi_1 _21644_ (.A1(_12528_),
    .A2(_12529_),
    .Y(_12530_),
    .B1(_12519_));
 sg13g2_nor3_1 _21645_ (.A(net806),
    .B(_12527_),
    .C(_12530_),
    .Y(_12531_));
 sg13g2_a21oi_1 _21646_ (.A1(net461),
    .A2(_12524_),
    .Y(_12532_),
    .B1(_12531_));
 sg13g2_inv_2 _21647_ (.Y(_12533_),
    .A(_12516_));
 sg13g2_xnor2_1 _21648_ (.Y(_12534_),
    .A(_12533_),
    .B(_12215_));
 sg13g2_xor2_1 _21649_ (.B(_12534_),
    .A(_12481_),
    .X(_12535_));
 sg13g2_nor2_1 _21650_ (.A(_12124_),
    .B(_12535_),
    .Y(_12536_));
 sg13g2_nor2_1 _21651_ (.A(net813),
    .B(net801),
    .Y(_12537_));
 sg13g2_nand2_1 _21652_ (.Y(_12538_),
    .A(_11857_),
    .B(_12537_));
 sg13g2_nor3_1 _21653_ (.A(net804),
    .B(net466),
    .C(net458),
    .Y(_12539_));
 sg13g2_nand2_1 _21654_ (.Y(_12540_),
    .A(_12452_),
    .B(net801));
 sg13g2_nor2_1 _21655_ (.A(_12214_),
    .B(_12540_),
    .Y(_12541_));
 sg13g2_o21ai_1 _21656_ (.B1(_11743_),
    .Y(_12542_),
    .A1(_12539_),
    .A2(_12541_));
 sg13g2_o21ai_1 _21657_ (.B1(_12542_),
    .Y(_12543_),
    .A1(net227),
    .A2(_12538_));
 sg13g2_nor3_1 _21658_ (.A(_12532_),
    .B(_12536_),
    .C(_12543_),
    .Y(_12544_));
 sg13g2_xnor2_1 _21659_ (.Y(_12545_),
    .A(_12175_),
    .B(_12516_));
 sg13g2_xnor2_1 _21660_ (.Y(_12546_),
    .A(_12452_),
    .B(net1098));
 sg13g2_xnor2_1 _21661_ (.Y(_12547_),
    .A(_12164_),
    .B(_12546_));
 sg13g2_xnor2_1 _21662_ (.Y(_12548_),
    .A(_12545_),
    .B(_12547_));
 sg13g2_buf_1 _21663_ (.A(_12548_),
    .X(_12549_));
 sg13g2_nor2_1 _21664_ (.A(_12485_),
    .B(_12549_),
    .Y(_12550_));
 sg13g2_nand2_1 _21665_ (.Y(_12551_),
    .A(net803),
    .B(_12549_));
 sg13g2_o21ai_1 _21666_ (.B1(_12551_),
    .Y(_12552_),
    .A1(net824),
    .A2(_12550_));
 sg13g2_o21ai_1 _21667_ (.B1(_12549_),
    .Y(_12553_),
    .A1(net803),
    .A2(_12536_));
 sg13g2_a21o_1 _21668_ (.A2(_12549_),
    .A1(_12167_),
    .B1(_12485_),
    .X(_12554_));
 sg13g2_mux2_1 _21669_ (.A0(_12550_),
    .A1(_12554_),
    .S(_12536_),
    .X(_12555_));
 sg13g2_a21o_1 _21670_ (.A2(_12553_),
    .A1(_11755_),
    .B1(_12555_),
    .X(_12556_));
 sg13g2_a21o_1 _21671_ (.A2(net458),
    .A1(net466),
    .B1(_11784_),
    .X(_12557_));
 sg13g2_o21ai_1 _21672_ (.B1(_12557_),
    .Y(_12558_),
    .A1(_11743_),
    .A2(_12545_));
 sg13g2_a22oi_1 _21673_ (.Y(_12559_),
    .B1(_12558_),
    .B2(_11857_),
    .A2(_12537_),
    .A1(_12519_));
 sg13g2_nand2_1 _21674_ (.Y(_12560_),
    .A(net477),
    .B(net806));
 sg13g2_a21o_1 _21675_ (.A2(_12560_),
    .A1(net227),
    .B1(_12538_),
    .X(_12561_));
 sg13g2_o21ai_1 _21676_ (.B1(_12561_),
    .Y(_12562_),
    .A1(net461),
    .A2(_12559_));
 sg13g2_a221oi_1 _21677_ (.B2(_12562_),
    .C1(net100),
    .B1(_12556_),
    .A1(_12544_),
    .Y(_12563_),
    .A2(_12552_));
 sg13g2_xnor2_1 _21678_ (.Y(_12564_),
    .A(_12493_),
    .B(_12549_));
 sg13g2_a21oi_1 _21679_ (.A1(net113),
    .A2(_12564_),
    .Y(_12565_),
    .B1(net221));
 sg13g2_or3_1 _21680_ (.A(net54),
    .B(_12563_),
    .C(_12565_),
    .X(_12566_));
 sg13g2_a21oi_1 _21681_ (.A1(_12515_),
    .A2(_12566_),
    .Y(_00438_),
    .B1(net523));
 sg13g2_buf_1 _21682_ (.A(net458),
    .X(_12567_));
 sg13g2_nand2_1 _21683_ (.Y(_12568_),
    .A(_11795_),
    .B(net215));
 sg13g2_buf_1 _21684_ (.A(\grid.cell_28_2.se ),
    .X(_12569_));
 sg13g2_buf_1 _21685_ (.A(net1089),
    .X(_12570_));
 sg13g2_nor2_1 _21686_ (.A(net465),
    .B(net800),
    .Y(_12571_));
 sg13g2_nand2_1 _21687_ (.Y(_12572_),
    .A(_11893_),
    .B(_12571_));
 sg13g2_a21oi_1 _21688_ (.A1(net226),
    .A2(_12568_),
    .Y(_12573_),
    .B1(_12572_));
 sg13g2_nand2_1 _21689_ (.Y(_12574_),
    .A(net475),
    .B(net474));
 sg13g2_nand2_1 _21690_ (.Y(_12575_),
    .A(_12252_),
    .B(net800));
 sg13g2_inv_1 _21691_ (.Y(_12576_),
    .A(_12575_));
 sg13g2_xor2_1 _21692_ (.B(net1089),
    .A(net1094),
    .X(_12577_));
 sg13g2_nand2_1 _21693_ (.Y(_12578_),
    .A(net476),
    .B(_12577_));
 sg13g2_o21ai_1 _21694_ (.B1(_12578_),
    .Y(_12579_),
    .A1(net474),
    .A2(_12576_));
 sg13g2_a22oi_1 _21695_ (.Y(_12580_),
    .B1(_12579_),
    .B2(_11893_),
    .A2(_12574_),
    .A1(_12571_));
 sg13g2_nor2_1 _21696_ (.A(net215),
    .B(_12580_),
    .Y(_12581_));
 sg13g2_nor2_1 _21697_ (.A(_12573_),
    .B(_12581_),
    .Y(_12582_));
 sg13g2_inv_2 _21698_ (.Y(_12583_),
    .A(net1094));
 sg13g2_xnor2_1 _21699_ (.Y(_12584_),
    .A(_11770_),
    .B(_12516_));
 sg13g2_xnor2_1 _21700_ (.Y(_12585_),
    .A(_11835_),
    .B(net1089));
 sg13g2_xnor2_1 _21701_ (.Y(_12586_),
    .A(_12584_),
    .B(_12585_));
 sg13g2_xnor2_1 _21702_ (.Y(_12587_),
    .A(_12583_),
    .B(_12586_));
 sg13g2_nor2_1 _21703_ (.A(net812),
    .B(_12587_),
    .Y(_12588_));
 sg13g2_xor2_1 _21704_ (.B(_11835_),
    .A(_12098_),
    .X(_12589_));
 sg13g2_xnor2_1 _21705_ (.Y(_12590_),
    .A(_12589_),
    .B(_12584_));
 sg13g2_xnor2_1 _21706_ (.Y(_12591_),
    .A(_12577_),
    .B(_12590_));
 sg13g2_buf_1 _21707_ (.A(_12591_),
    .X(_12592_));
 sg13g2_buf_2 _21708_ (.A(_00006_),
    .X(_12593_));
 sg13g2_buf_1 _21709_ (.A(_12593_),
    .X(_12594_));
 sg13g2_a21o_1 _21710_ (.A2(_12592_),
    .A1(_11744_),
    .B1(net799),
    .X(_12595_));
 sg13g2_o21ai_1 _21711_ (.B1(_12592_),
    .Y(_12596_),
    .A1(net799),
    .A2(_12588_));
 sg13g2_nor2_1 _21712_ (.A(net799),
    .B(_12592_),
    .Y(_12597_));
 sg13g2_nor2b_1 _21713_ (.A(_12588_),
    .B_N(_12597_),
    .Y(_12598_));
 sg13g2_a221oi_1 _21714_ (.B2(_11741_),
    .C1(_12598_),
    .B1(_12596_),
    .A1(_12588_),
    .Y(_12599_),
    .A2(_12595_));
 sg13g2_or2_1 _21715_ (.X(_12600_),
    .B(_12599_),
    .A(_12582_));
 sg13g2_nor3_1 _21716_ (.A(net215),
    .B(_12574_),
    .C(_12575_),
    .Y(_12601_));
 sg13g2_o21ai_1 _21717_ (.B1(_12578_),
    .Y(_12602_),
    .A1(net475),
    .A2(_12575_));
 sg13g2_a22oi_1 _21718_ (.Y(_12603_),
    .B1(_12602_),
    .B2(net226),
    .A2(_12576_),
    .A1(_11899_));
 sg13g2_nor2_1 _21719_ (.A(_12533_),
    .B(_12603_),
    .Y(_12604_));
 sg13g2_nor2_1 _21720_ (.A(_11729_),
    .B(_12597_),
    .Y(_12605_));
 sg13g2_a21oi_1 _21721_ (.A1(net799),
    .A2(_12592_),
    .Y(_12606_),
    .B1(_12605_));
 sg13g2_nor4_1 _21722_ (.A(_12588_),
    .B(_12601_),
    .C(_12604_),
    .D(_12606_),
    .Y(_12607_));
 sg13g2_a221oi_1 _21723_ (.B2(_12607_),
    .C1(net73),
    .B1(_12582_),
    .A1(_05811_),
    .Y(_12608_),
    .A2(net54));
 sg13g2_xor2_1 _21724_ (.B(_12592_),
    .A(_12481_),
    .X(_12609_));
 sg13g2_nand2_1 _21725_ (.Y(_12610_),
    .A(net111),
    .B(_12609_));
 sg13g2_nor2_1 _21726_ (.A(net220),
    .B(net54),
    .Y(_12611_));
 sg13g2_a22oi_1 _21727_ (.Y(_12612_),
    .B1(_12610_),
    .B2(_12611_),
    .A2(net54),
    .A1(net35));
 sg13g2_nand2_1 _21728_ (.Y(_12613_),
    .A(net312),
    .B(_12612_));
 sg13g2_a21oi_1 _21729_ (.A1(_12600_),
    .A2(_12608_),
    .Y(_00439_),
    .B1(_12613_));
 sg13g2_nand3_1 _21730_ (.B(net104),
    .C(net55),
    .A(_12264_),
    .Y(_12614_));
 sg13g2_o21ai_1 _21731_ (.B1(_12614_),
    .Y(_12615_),
    .A1(net48),
    .A2(_12450_));
 sg13g2_buf_1 _21732_ (.A(net800),
    .X(_12616_));
 sg13g2_buf_1 _21733_ (.A(\grid.cell_28_3.se ),
    .X(_12617_));
 sg13g2_buf_1 _21734_ (.A(net1088),
    .X(_12618_));
 sg13g2_nand2_1 _21735_ (.Y(_12619_),
    .A(net810),
    .B(net798));
 sg13g2_nand2_1 _21736_ (.Y(_12620_),
    .A(net226),
    .B(net225));
 sg13g2_or2_1 _21737_ (.X(_12621_),
    .B(_12620_),
    .A(_12619_));
 sg13g2_xor2_1 _21738_ (.B(net1088),
    .A(_12265_),
    .X(_12622_));
 sg13g2_nand2_1 _21739_ (.Y(_12623_),
    .A(net474),
    .B(_12622_));
 sg13g2_o21ai_1 _21740_ (.B1(_12623_),
    .Y(_12624_),
    .A1(net474),
    .A2(_12619_));
 sg13g2_nand2_1 _21741_ (.Y(_12625_),
    .A(net225),
    .B(_12624_));
 sg13g2_o21ai_1 _21742_ (.B1(_12625_),
    .Y(_12626_),
    .A1(_11928_),
    .A2(_12619_));
 sg13g2_nand2_1 _21743_ (.Y(_12627_),
    .A(net1197),
    .B(net55));
 sg13g2_a21oi_1 _21744_ (.A1(net457),
    .A2(_12626_),
    .Y(_12628_),
    .B1(_12627_));
 sg13g2_o21ai_1 _21745_ (.B1(_12628_),
    .Y(_12629_),
    .A1(net457),
    .A2(_12621_));
 sg13g2_buf_1 _21746_ (.A(_00005_),
    .X(_12630_));
 sg13g2_xnor2_1 _21747_ (.Y(_12631_),
    .A(_11879_),
    .B(_12622_));
 sg13g2_xor2_1 _21748_ (.B(_12631_),
    .A(_12585_),
    .X(_12632_));
 sg13g2_nor4_1 _21749_ (.A(_12630_),
    .B(_12277_),
    .C(_12215_),
    .D(_12632_),
    .Y(_12633_));
 sg13g2_xnor2_1 _21750_ (.Y(_12634_),
    .A(_12534_),
    .B(_12632_));
 sg13g2_a21oi_1 _21751_ (.A1(net70),
    .A2(_12634_),
    .Y(_12635_),
    .B1(net465));
 sg13g2_nand2b_1 _21752_ (.Y(_12636_),
    .B(_12630_),
    .A_N(_11795_));
 sg13g2_xnor2_1 _21753_ (.Y(_12637_),
    .A(net220),
    .B(_12632_));
 sg13g2_inv_1 _21754_ (.Y(_12638_),
    .A(_12630_));
 sg13g2_nand2_1 _21755_ (.Y(_12639_),
    .A(_11851_),
    .B(_12638_));
 sg13g2_o21ai_1 _21756_ (.B1(_12639_),
    .Y(_12640_),
    .A1(_12277_),
    .A2(_12632_));
 sg13g2_a21oi_1 _21757_ (.A1(_12636_),
    .A2(_12637_),
    .Y(_12641_),
    .B1(_12640_));
 sg13g2_a22oi_1 _21758_ (.Y(_12642_),
    .B1(_12619_),
    .B2(_11879_),
    .A2(_12622_),
    .A1(_11853_));
 sg13g2_a21oi_1 _21759_ (.A1(_11843_),
    .A2(net800),
    .Y(_12643_),
    .B1(_11879_));
 sg13g2_or3_1 _21760_ (.A(net464),
    .B(net798),
    .C(_12643_),
    .X(_12644_));
 sg13g2_o21ai_1 _21761_ (.B1(_12644_),
    .Y(_12645_),
    .A1(net457),
    .A2(_12642_));
 sg13g2_buf_1 _21762_ (.A(net798),
    .X(_12646_));
 sg13g2_nor3_1 _21763_ (.A(net457),
    .B(net219),
    .C(net456),
    .Y(_12647_));
 sg13g2_a22oi_1 _21764_ (.Y(_12648_),
    .B1(_12647_),
    .B2(_12620_),
    .A2(_12645_),
    .A1(_11928_));
 sg13g2_xor2_1 _21765_ (.B(_12648_),
    .A(_12641_),
    .X(_12649_));
 sg13g2_nor4_1 _21766_ (.A(_12629_),
    .B(_12633_),
    .C(_12635_),
    .D(_12649_),
    .Y(_12650_));
 sg13g2_a21o_1 _21767_ (.A2(_12615_),
    .A1(net312),
    .B1(_12650_),
    .X(_00440_));
 sg13g2_buf_2 _21768_ (.A(net715),
    .X(_12651_));
 sg13g2_buf_1 _21769_ (.A(\grid.cell_28_4.se ),
    .X(_12652_));
 sg13g2_buf_1 _21770_ (.A(_12652_),
    .X(_12653_));
 sg13g2_xor2_1 _21771_ (.B(_12311_),
    .A(net797),
    .X(_12654_));
 sg13g2_xnor2_1 _21772_ (.Y(_12655_),
    .A(net820),
    .B(net1088));
 sg13g2_xnor2_1 _21773_ (.Y(_12656_),
    .A(_12654_),
    .B(_12655_));
 sg13g2_nand2b_1 _21774_ (.Y(_12657_),
    .B(_12656_),
    .A_N(net1093));
 sg13g2_buf_2 _21775_ (.A(_00060_),
    .X(_12658_));
 sg13g2_inv_1 _21776_ (.Y(_12659_),
    .A(_12658_));
 sg13g2_nand2_1 _21777_ (.Y(_12660_),
    .A(_12659_),
    .B(net226));
 sg13g2_buf_1 _21778_ (.A(net797),
    .X(_12661_));
 sg13g2_nand2_1 _21779_ (.Y(_12662_),
    .A(net809),
    .B(_12661_));
 sg13g2_xor2_1 _21780_ (.B(_12652_),
    .A(_12300_),
    .X(_12663_));
 sg13g2_and2_1 _21781_ (.A(_11878_),
    .B(_12663_),
    .X(_12664_));
 sg13g2_nor2_1 _21782_ (.A(_11885_),
    .B(_12662_),
    .Y(_12665_));
 sg13g2_o21ai_1 _21783_ (.B1(net472),
    .Y(_12666_),
    .A1(_12664_),
    .A2(_12665_));
 sg13g2_o21ai_1 _21784_ (.B1(_12666_),
    .Y(_12667_),
    .A1(_11984_),
    .A2(_12662_));
 sg13g2_nand2_1 _21785_ (.Y(_12668_),
    .A(_11885_),
    .B(net472));
 sg13g2_nor3_1 _21786_ (.A(net456),
    .B(_12662_),
    .C(_12668_),
    .Y(_12669_));
 sg13g2_a21oi_1 _21787_ (.A1(net456),
    .A2(_12667_),
    .Y(_12670_),
    .B1(_12669_));
 sg13g2_xnor2_1 _21788_ (.Y(_12671_),
    .A(_12583_),
    .B(_12656_));
 sg13g2_o21ai_1 _21789_ (.B1(_12671_),
    .Y(_12672_),
    .A1(_12659_),
    .A2(net226));
 sg13g2_nand4_1 _21790_ (.B(_12660_),
    .C(_12670_),
    .A(_12657_),
    .Y(_12673_),
    .D(_12672_));
 sg13g2_a21oi_1 _21791_ (.A1(_11921_),
    .A2(_12662_),
    .Y(_12674_),
    .B1(_12664_));
 sg13g2_a21oi_1 _21792_ (.A1(net820),
    .A2(net798),
    .Y(_12675_),
    .B1(_11921_));
 sg13g2_or3_1 _21793_ (.A(net463),
    .B(net455),
    .C(_12675_),
    .X(_12676_));
 sg13g2_o21ai_1 _21794_ (.B1(_12676_),
    .Y(_12677_),
    .A1(net456),
    .A2(_12674_));
 sg13g2_buf_1 _21795_ (.A(net455),
    .X(_12678_));
 sg13g2_nor3_1 _21796_ (.A(net456),
    .B(net463),
    .C(net213),
    .Y(_12679_));
 sg13g2_a22oi_1 _21797_ (.Y(_12680_),
    .B1(_12679_),
    .B2(_12668_),
    .A2(_12677_),
    .A1(_11984_));
 sg13g2_and2_1 _21798_ (.A(net127),
    .B(_12680_),
    .X(_12681_));
 sg13g2_and2_1 _21799_ (.A(_11854_),
    .B(_12671_),
    .X(_12682_));
 sg13g2_nor2_1 _21800_ (.A(_12659_),
    .B(_12657_),
    .Y(_12683_));
 sg13g2_nor4_1 _21801_ (.A(net166),
    .B(_12680_),
    .C(_12682_),
    .D(_12683_),
    .Y(_12684_));
 sg13g2_a21oi_1 _21802_ (.A1(_12583_),
    .A2(_12656_),
    .Y(_12685_),
    .B1(net226));
 sg13g2_nand2b_1 _21803_ (.Y(_12686_),
    .B(net1093),
    .A_N(_12685_));
 sg13g2_or2_1 _21804_ (.X(_12687_),
    .B(net474),
    .A(net1093));
 sg13g2_nand3_1 _21805_ (.B(_12656_),
    .C(_12687_),
    .A(net465),
    .Y(_12688_));
 sg13g2_nand2b_1 _21806_ (.Y(_12689_),
    .B(_12688_),
    .A_N(_12253_));
 sg13g2_a21o_1 _21807_ (.A2(_12689_),
    .A1(_12686_),
    .B1(_12658_),
    .X(_12690_));
 sg13g2_a22oi_1 _21808_ (.Y(_12691_),
    .B1(_12684_),
    .B2(_12690_),
    .A2(_12681_),
    .A1(_12673_));
 sg13g2_xnor2_1 _21809_ (.Y(_12692_),
    .A(_12585_),
    .B(_12671_));
 sg13g2_a21oi_1 _21810_ (.A1(net98),
    .A2(_12692_),
    .Y(_12693_),
    .B1(_12286_));
 sg13g2_nor2_1 _21811_ (.A(net54),
    .B(_12693_),
    .Y(_12694_));
 sg13g2_a22oi_1 _21812_ (.Y(_12695_),
    .B1(_12691_),
    .B2(_12694_),
    .A2(_12514_),
    .A1(_07426_));
 sg13g2_nor2_1 _21813_ (.A(net214),
    .B(_12695_),
    .Y(_00441_));
 sg13g2_inv_1 _21814_ (.Y(_12696_),
    .A(_12357_));
 sg13g2_buf_1 _21815_ (.A(_00092_),
    .X(_12697_));
 sg13g2_inv_1 _21816_ (.Y(_12698_),
    .A(net1087));
 sg13g2_buf_1 _21817_ (.A(\grid.cell_28_5.se ),
    .X(_12699_));
 sg13g2_buf_1 _21818_ (.A(_12699_),
    .X(_12700_));
 sg13g2_xnor2_1 _21819_ (.Y(_12701_),
    .A(net797),
    .B(net796));
 sg13g2_xnor2_1 _21820_ (.Y(_12702_),
    .A(_12340_),
    .B(_12701_));
 sg13g2_xnor2_1 _21821_ (.Y(_12703_),
    .A(net1096),
    .B(_12702_));
 sg13g2_buf_1 _21822_ (.A(_12703_),
    .X(_12704_));
 sg13g2_nand2_1 _21823_ (.Y(_12705_),
    .A(_12698_),
    .B(net219));
 sg13g2_o21ai_1 _21824_ (.B1(_12705_),
    .Y(_12706_),
    .A1(_12698_),
    .A2(_12704_));
 sg13g2_nor2_1 _21825_ (.A(_12286_),
    .B(_12704_),
    .Y(_12707_));
 sg13g2_a21oi_1 _21826_ (.A1(_12357_),
    .A2(_12707_),
    .Y(_12708_),
    .B1(net225));
 sg13g2_and2_1 _21827_ (.A(net464),
    .B(_12704_),
    .X(_12709_));
 sg13g2_buf_1 _21828_ (.A(_12709_),
    .X(_12710_));
 sg13g2_nand2_1 _21829_ (.Y(_12711_),
    .A(net1087),
    .B(_11879_));
 sg13g2_xor2_1 _21830_ (.B(net796),
    .A(_12334_),
    .X(_12712_));
 sg13g2_nand2_2 _21831_ (.Y(_12713_),
    .A(net808),
    .B(net796));
 sg13g2_a22oi_1 _21832_ (.Y(_12714_),
    .B1(_12713_),
    .B2(_12013_),
    .A2(_12712_),
    .A1(_11918_));
 sg13g2_and2_1 _21833_ (.A(net1096),
    .B(net797),
    .X(_12715_));
 sg13g2_buf_1 _21834_ (.A(net796),
    .X(_12716_));
 sg13g2_nor2_1 _21835_ (.A(net808),
    .B(net454),
    .Y(_12717_));
 sg13g2_o21ai_1 _21836_ (.B1(_12717_),
    .Y(_12718_),
    .A1(_12013_),
    .A2(_12715_));
 sg13g2_o21ai_1 _21837_ (.B1(_12718_),
    .Y(_12719_),
    .A1(net455),
    .A2(_12714_));
 sg13g2_nand2_1 _21838_ (.Y(_12720_),
    .A(net819),
    .B(_11989_));
 sg13g2_buf_1 _21839_ (.A(net454),
    .X(_12721_));
 sg13g2_nor3_1 _21840_ (.A(net213),
    .B(_12387_),
    .C(net212),
    .Y(_12722_));
 sg13g2_a22oi_1 _21841_ (.Y(_12723_),
    .B1(_12720_),
    .B2(_12722_),
    .A2(_12719_),
    .A1(_12021_));
 sg13g2_buf_1 _21842_ (.A(_12723_),
    .X(_12724_));
 sg13g2_a221oi_1 _21843_ (.B2(_12711_),
    .C1(_12724_),
    .B1(_12710_),
    .A1(net225),
    .Y(_12725_),
    .A2(_12707_));
 sg13g2_o21ai_1 _21844_ (.B1(_12725_),
    .Y(_12726_),
    .A1(net1087),
    .A2(_12708_));
 sg13g2_a21oi_1 _21845_ (.A1(_12696_),
    .A2(_12706_),
    .Y(_12727_),
    .B1(_12726_));
 sg13g2_nor2_1 _21846_ (.A(net1087),
    .B(_12267_),
    .Y(_12728_));
 sg13g2_o21ai_1 _21847_ (.B1(_12696_),
    .Y(_12729_),
    .A1(_12724_),
    .A2(_12728_));
 sg13g2_nand3_1 _21848_ (.B(_12724_),
    .C(_12711_),
    .A(_12314_),
    .Y(_12730_));
 sg13g2_a21o_1 _21849_ (.A2(_12730_),
    .A1(_12729_),
    .B1(_12704_),
    .X(_12731_));
 sg13g2_nand2_1 _21850_ (.Y(_12732_),
    .A(net472),
    .B(_12712_));
 sg13g2_o21ai_1 _21851_ (.B1(_12732_),
    .Y(_12733_),
    .A1(net472),
    .A2(_12713_));
 sg13g2_nor2_1 _21852_ (.A(net1095),
    .B(_12713_),
    .Y(_12734_));
 sg13g2_a21oi_1 _21853_ (.A1(_11990_),
    .A2(_12733_),
    .Y(_12735_),
    .B1(_12734_));
 sg13g2_nor2b_1 _21854_ (.A(_12735_),
    .B_N(net213),
    .Y(_12736_));
 sg13g2_nor3_1 _21855_ (.A(net213),
    .B(_12713_),
    .C(_12720_),
    .Y(_12737_));
 sg13g2_xnor2_1 _21856_ (.Y(_12738_),
    .A(_12631_),
    .B(_12704_));
 sg13g2_a21oi_1 _21857_ (.A1(net123),
    .A2(_12738_),
    .Y(_12739_),
    .B1(net463));
 sg13g2_nor4_1 _21858_ (.A(_12627_),
    .B(_12736_),
    .C(_12737_),
    .D(_12739_),
    .Y(_12740_));
 sg13g2_nor2_1 _21859_ (.A(net225),
    .B(_12710_),
    .Y(_12741_));
 sg13g2_nand2_1 _21860_ (.Y(_12742_),
    .A(_11886_),
    .B(_12710_));
 sg13g2_o21ai_1 _21861_ (.B1(_12742_),
    .Y(_12743_),
    .A1(net1087),
    .A2(_12741_));
 sg13g2_nand2_1 _21862_ (.Y(_12744_),
    .A(_12724_),
    .B(_12743_));
 sg13g2_nand3_1 _21863_ (.B(_12740_),
    .C(_12744_),
    .A(_12731_),
    .Y(_12745_));
 sg13g2_nand3_1 _21864_ (.B(net110),
    .C(net55),
    .A(net463),
    .Y(_12746_));
 sg13g2_o21ai_1 _21865_ (.B1(_12746_),
    .Y(_12747_),
    .A1(_05002_),
    .A2(net55));
 sg13g2_nand2_1 _21866_ (.Y(_12748_),
    .A(net312),
    .B(_12747_));
 sg13g2_o21ai_1 _21867_ (.B1(_12748_),
    .Y(_00442_),
    .A1(_12727_),
    .A2(_12745_));
 sg13g2_nand2_1 _21868_ (.Y(_12749_),
    .A(net31),
    .B(net54));
 sg13g2_inv_1 _21869_ (.Y(_12750_),
    .A(_12392_));
 sg13g2_xnor2_1 _21870_ (.Y(_12751_),
    .A(_12699_),
    .B(net1090));
 sg13g2_xor2_1 _21871_ (.B(_12751_),
    .A(_12150_),
    .X(_12752_));
 sg13g2_xnor2_1 _21872_ (.Y(_12753_),
    .A(net818),
    .B(_12752_));
 sg13g2_xnor2_1 _21873_ (.Y(_12754_),
    .A(_12301_),
    .B(_12753_));
 sg13g2_a22oi_1 _21874_ (.Y(_12755_),
    .B1(_12754_),
    .B2(net472),
    .A2(_12753_),
    .A1(_12750_));
 sg13g2_buf_1 _21875_ (.A(_00124_),
    .X(_12756_));
 sg13g2_xnor2_1 _21876_ (.Y(_12757_),
    .A(_12311_),
    .B(_12753_));
 sg13g2_nor2_1 _21877_ (.A(_12756_),
    .B(_12757_),
    .Y(_12758_));
 sg13g2_buf_1 _21878_ (.A(_00154_),
    .X(_12759_));
 sg13g2_xor2_1 _21879_ (.B(net212),
    .A(net1086),
    .X(_12760_));
 sg13g2_nand3_1 _21880_ (.B(net212),
    .C(_12501_),
    .A(net1086),
    .Y(_12761_));
 sg13g2_o21ai_1 _21881_ (.B1(_12761_),
    .Y(_12762_),
    .A1(net1086),
    .A2(_12501_));
 sg13g2_a21oi_1 _21882_ (.A1(_12475_),
    .A2(_12760_),
    .Y(_12763_),
    .B1(_12762_));
 sg13g2_inv_1 _21883_ (.Y(_12764_),
    .A(net796));
 sg13g2_nor2_1 _21884_ (.A(net815),
    .B(net805),
    .Y(_12765_));
 sg13g2_nand2_1 _21885_ (.Y(_12766_),
    .A(_12764_),
    .B(_12765_));
 sg13g2_a21oi_1 _21886_ (.A1(net468),
    .A2(net805),
    .Y(_12767_),
    .B1(net454));
 sg13g2_o21ai_1 _21887_ (.B1(net1086),
    .Y(_12768_),
    .A1(_12765_),
    .A2(_12767_));
 sg13g2_a21oi_1 _21888_ (.A1(_12766_),
    .A2(_12768_),
    .Y(_12769_),
    .B1(net470));
 sg13g2_nand4_1 _21889_ (.B(_12033_),
    .C(_12101_),
    .A(net454),
    .Y(_12770_),
    .D(net460));
 sg13g2_a21oi_1 _21890_ (.A1(_12766_),
    .A2(_12770_),
    .Y(_12771_),
    .B1(net224));
 sg13g2_nor3_1 _21891_ (.A(net1086),
    .B(_12764_),
    .C(_12501_),
    .Y(_12772_));
 sg13g2_nor3_1 _21892_ (.A(_12769_),
    .B(_12771_),
    .C(_12772_),
    .Y(_12773_));
 sg13g2_o21ai_1 _21893_ (.B1(_12773_),
    .Y(_12774_),
    .A1(_12063_),
    .A2(_12763_));
 sg13g2_nor2_1 _21894_ (.A(_12758_),
    .B(_12774_),
    .Y(_12775_));
 sg13g2_buf_1 _21895_ (.A(net212),
    .X(_12776_));
 sg13g2_a22oi_1 _21896_ (.Y(_12777_),
    .B1(_12502_),
    .B2(_11990_),
    .A2(_12501_),
    .A1(_12109_));
 sg13g2_nor2_1 _21897_ (.A(net136),
    .B(_12777_),
    .Y(_12778_));
 sg13g2_nand2_1 _21898_ (.Y(_12779_),
    .A(net224),
    .B(net212));
 sg13g2_a21oi_1 _21899_ (.A1(net222),
    .A2(_12779_),
    .Y(_12780_),
    .B1(_12475_));
 sg13g2_o21ai_1 _21900_ (.B1(net1086),
    .Y(_12781_),
    .A1(_12778_),
    .A2(_12780_));
 sg13g2_o21ai_1 _21901_ (.B1(_12781_),
    .Y(_12782_),
    .A1(_12067_),
    .A2(_12766_));
 sg13g2_xnor2_1 _21902_ (.Y(_12783_),
    .A(_12755_),
    .B(_12758_));
 sg13g2_a221oi_1 _21903_ (.B2(_12783_),
    .C1(net100),
    .B1(_12782_),
    .A1(_12755_),
    .Y(_12784_),
    .A2(_12775_));
 sg13g2_xor2_1 _21904_ (.B(_12753_),
    .A(_12654_),
    .X(_12785_));
 sg13g2_a21oi_1 _21905_ (.A1(net113),
    .A2(_12785_),
    .Y(_12786_),
    .B1(net218));
 sg13g2_or3_1 _21906_ (.A(net54),
    .B(_12784_),
    .C(_12786_),
    .X(_12787_));
 sg13g2_a21oi_1 _21907_ (.A1(_12749_),
    .A2(_12787_),
    .Y(_00443_),
    .B1(net523));
 sg13g2_nand3_1 _21908_ (.B(net120),
    .C(net55),
    .A(net217),
    .Y(_12788_));
 sg13g2_o21ai_1 _21909_ (.B1(_12788_),
    .Y(_12789_),
    .A1(net121),
    .A2(net55));
 sg13g2_nand2_1 _21910_ (.Y(_12790_),
    .A(net796),
    .B(net1090));
 sg13g2_buf_2 _21911_ (.A(_12790_),
    .X(_12791_));
 sg13g2_o21ai_1 _21912_ (.B1(net462),
    .Y(_12792_),
    .A1(net212),
    .A2(net459));
 sg13g2_a21o_1 _21913_ (.A2(_12792_),
    .A1(_12791_),
    .B1(_12109_),
    .X(_12793_));
 sg13g2_mux2_1 _21914_ (.A0(net136),
    .A1(_12791_),
    .S(net462),
    .X(_12794_));
 sg13g2_a22oi_1 _21915_ (.Y(_12795_),
    .B1(_12794_),
    .B2(net222),
    .A2(_12717_),
    .A1(net137));
 sg13g2_mux2_1 _21916_ (.A0(_12793_),
    .A1(_12795_),
    .S(net1086),
    .X(_12796_));
 sg13g2_nand2_1 _21917_ (.Y(_12797_),
    .A(_12034_),
    .B(net216));
 sg13g2_or3_1 _21918_ (.A(net462),
    .B(net212),
    .C(net216),
    .X(_12798_));
 sg13g2_o21ai_1 _21919_ (.B1(_12798_),
    .Y(_12799_),
    .A1(_12713_),
    .A2(_12797_));
 sg13g2_nor2_1 _21920_ (.A(_12759_),
    .B(_12791_),
    .Y(_12800_));
 sg13g2_nand3_1 _21921_ (.B(_12791_),
    .C(_12792_),
    .A(net1086),
    .Y(_12801_));
 sg13g2_a21oi_1 _21922_ (.A1(_12798_),
    .A2(_12801_),
    .Y(_12802_),
    .B1(_12034_));
 sg13g2_a221oi_1 _21923_ (.B2(net218),
    .C1(_12802_),
    .B1(_12800_),
    .A1(net223),
    .Y(_12803_),
    .A2(_12799_));
 sg13g2_o21ai_1 _21924_ (.B1(_12803_),
    .Y(_12804_),
    .A1(net223),
    .A2(_12796_));
 sg13g2_xor2_1 _21925_ (.B(_12751_),
    .A(_12340_),
    .X(_12805_));
 sg13g2_xnor2_1 _21926_ (.Y(_12806_),
    .A(_12033_),
    .B(_12805_));
 sg13g2_xor2_1 _21927_ (.B(_12806_),
    .A(net807),
    .X(_12807_));
 sg13g2_nand2b_1 _21928_ (.Y(_12808_),
    .B(_12806_),
    .A_N(_12125_));
 sg13g2_nand2b_1 _21929_ (.Y(_12809_),
    .B(_12808_),
    .A_N(_12488_));
 sg13g2_a21oi_1 _21930_ (.A1(_12487_),
    .A2(_12807_),
    .Y(_12810_),
    .B1(_12809_));
 sg13g2_xor2_1 _21931_ (.B(_12810_),
    .A(_12804_),
    .X(_12811_));
 sg13g2_mux2_1 _21932_ (.A0(_12751_),
    .A1(_12791_),
    .S(net223),
    .X(_12812_));
 sg13g2_nor2_1 _21933_ (.A(_12109_),
    .B(_12812_),
    .Y(_12813_));
 sg13g2_o21ai_1 _21934_ (.B1(net218),
    .Y(_12814_),
    .A1(_12800_),
    .A2(_12813_));
 sg13g2_nand4_1 _21935_ (.B(net136),
    .C(net137),
    .A(_12382_),
    .Y(_12815_),
    .D(_12067_));
 sg13g2_nand4_1 _21936_ (.B(net127),
    .C(_12814_),
    .A(net1054),
    .Y(_12816_),
    .D(_12815_));
 sg13g2_nor3_1 _21937_ (.A(_07600_),
    .B(_11347_),
    .C(_12448_),
    .Y(_12817_));
 sg13g2_inv_1 _21938_ (.Y(_12818_),
    .A(_12209_));
 sg13g2_nor3_1 _21939_ (.A(net803),
    .B(_12818_),
    .C(_12808_),
    .Y(_12819_));
 sg13g2_inv_1 _21940_ (.Y(_12820_),
    .A(_12491_));
 sg13g2_xnor2_1 _21941_ (.Y(_12821_),
    .A(_12820_),
    .B(_12209_));
 sg13g2_xnor2_1 _21942_ (.Y(_12822_),
    .A(_12806_),
    .B(_12821_));
 sg13g2_nor2_1 _21943_ (.A(net217),
    .B(_12822_),
    .Y(_12823_));
 sg13g2_nor4_1 _21944_ (.A(_12816_),
    .B(_12817_),
    .C(_12819_),
    .D(_12823_),
    .Y(_12824_));
 sg13g2_a22oi_1 _21945_ (.Y(_12825_),
    .B1(_12811_),
    .B2(_12824_),
    .A2(_12789_),
    .A1(net356));
 sg13g2_inv_1 _21946_ (.Y(_00444_),
    .A(_12825_));
 sg13g2_nor3_2 _21947_ (.A(_07972_),
    .B(net320),
    .C(_12448_),
    .Y(_12826_));
 sg13g2_and2_1 _21948_ (.A(net327),
    .B(_12826_),
    .X(_12827_));
 sg13g2_buf_1 _21949_ (.A(_12827_),
    .X(_12828_));
 sg13g2_buf_1 _21950_ (.A(\grid.cell_29_0.se ),
    .X(_12829_));
 sg13g2_buf_2 _21951_ (.A(_12829_),
    .X(_12830_));
 sg13g2_inv_2 _21952_ (.Y(_12831_),
    .A(net795));
 sg13g2_buf_1 _21953_ (.A(\grid.cell_29_0.sw ),
    .X(_12832_));
 sg13g2_buf_1 _21954_ (.A(_12832_),
    .X(_12833_));
 sg13g2_buf_1 _21955_ (.A(net794),
    .X(_12834_));
 sg13g2_nor2_1 _21956_ (.A(net805),
    .B(net453),
    .Y(_12835_));
 sg13g2_nand2_1 _21957_ (.Y(_12836_),
    .A(_12831_),
    .B(_12835_));
 sg13g2_buf_1 _21958_ (.A(net794),
    .X(_12837_));
 sg13g2_nand4_1 _21959_ (.B(_12101_),
    .C(net459),
    .A(net795),
    .Y(_12838_),
    .D(net452));
 sg13g2_a21oi_1 _21960_ (.A1(_12836_),
    .A2(_12838_),
    .Y(_12839_),
    .B1(net469));
 sg13g2_nand2b_1 _21961_ (.Y(_12840_),
    .B(_12239_),
    .A_N(net794));
 sg13g2_nor2_1 _21962_ (.A(_12475_),
    .B(_12840_),
    .Y(_12841_));
 sg13g2_nand2_1 _21963_ (.Y(_12842_),
    .A(net816),
    .B(_12100_));
 sg13g2_nand2b_1 _21964_ (.Y(_12843_),
    .B(net453),
    .A_N(_12239_));
 sg13g2_o21ai_1 _21965_ (.B1(_12843_),
    .Y(_12844_),
    .A1(net452),
    .A2(_12842_));
 sg13g2_nor2_1 _21966_ (.A(net453),
    .B(net812),
    .Y(_12845_));
 sg13g2_nor3_1 _21967_ (.A(net460),
    .B(_12842_),
    .C(_12845_),
    .Y(_12846_));
 sg13g2_a21oi_1 _21968_ (.A1(net459),
    .A2(_12844_),
    .Y(_12847_),
    .B1(_12846_));
 sg13g2_nor2_1 _21969_ (.A(_12831_),
    .B(_12847_),
    .Y(_12848_));
 sg13g2_buf_2 _21970_ (.A(net795),
    .X(_12849_));
 sg13g2_nor2b_1 _21971_ (.A(_12239_),
    .B_N(net794),
    .Y(_12850_));
 sg13g2_o21ai_1 _21972_ (.B1(_12840_),
    .Y(_12851_),
    .A1(net805),
    .A2(_12850_));
 sg13g2_nand2_1 _21973_ (.Y(_12852_),
    .A(net453),
    .B(net812));
 sg13g2_o21ai_1 _21974_ (.B1(net805),
    .Y(_12853_),
    .A1(net453),
    .A2(net812));
 sg13g2_a21oi_1 _21975_ (.A1(_12852_),
    .A2(_12853_),
    .Y(_12854_),
    .B1(_12842_));
 sg13g2_a21oi_1 _21976_ (.A1(net467),
    .A2(_12851_),
    .Y(_12855_),
    .B1(_12854_));
 sg13g2_nor2_1 _21977_ (.A(net451),
    .B(_12855_),
    .Y(_12856_));
 sg13g2_nor4_1 _21978_ (.A(_12839_),
    .B(_12841_),
    .C(_12848_),
    .D(_12856_),
    .Y(_12857_));
 sg13g2_xnor2_1 _21979_ (.Y(_12858_),
    .A(_12097_),
    .B(_12829_));
 sg13g2_inv_1 _21980_ (.Y(_12859_),
    .A(_12832_));
 sg13g2_xnor2_1 _21981_ (.Y(_12860_),
    .A(_12859_),
    .B(_12502_));
 sg13g2_xor2_1 _21982_ (.B(_12860_),
    .A(_12858_),
    .X(_12861_));
 sg13g2_xnor2_1 _21983_ (.Y(_12862_),
    .A(net806),
    .B(_12861_));
 sg13g2_buf_1 _21984_ (.A(_00272_),
    .X(_12863_));
 sg13g2_buf_1 _21985_ (.A(_12863_),
    .X(_12864_));
 sg13g2_nand2b_1 _21986_ (.Y(_12865_),
    .B(net793),
    .A_N(_12163_));
 sg13g2_inv_2 _21987_ (.Y(_12866_),
    .A(_12863_));
 sg13g2_nand2_1 _21988_ (.Y(_12867_),
    .A(_12163_),
    .B(_12866_));
 sg13g2_o21ai_1 _21989_ (.B1(_12867_),
    .Y(_12868_),
    .A1(net799),
    .A2(_12861_));
 sg13g2_a21oi_1 _21990_ (.A1(_12862_),
    .A2(_12865_),
    .Y(_12869_),
    .B1(_12868_));
 sg13g2_xnor2_1 _21991_ (.Y(_12870_),
    .A(net1090),
    .B(_12832_));
 sg13g2_a21oi_1 _21992_ (.A1(net460),
    .A2(net452),
    .Y(_12871_),
    .B1(net816));
 sg13g2_a21oi_1 _21993_ (.A1(net469),
    .A2(_12870_),
    .Y(_12872_),
    .B1(_12871_));
 sg13g2_a22oi_1 _21994_ (.Y(_12873_),
    .B1(_12872_),
    .B2(net217),
    .A2(_12850_),
    .A1(net216));
 sg13g2_nand2_1 _21995_ (.Y(_12874_),
    .A(net1090),
    .B(net794));
 sg13g2_or3_1 _21996_ (.A(net451),
    .B(_12874_),
    .C(_12842_),
    .X(_12875_));
 sg13g2_o21ai_1 _21997_ (.B1(_12875_),
    .Y(_12876_),
    .A1(_12831_),
    .A2(_12873_));
 sg13g2_xor2_1 _21998_ (.B(net804),
    .A(_12163_),
    .X(_12877_));
 sg13g2_nor4_1 _21999_ (.A(net793),
    .B(net799),
    .C(_12877_),
    .D(_12861_),
    .Y(_12878_));
 sg13g2_nor2_1 _22000_ (.A(_12876_),
    .B(_12878_),
    .Y(_12879_));
 sg13g2_nand3_1 _22001_ (.B(_12869_),
    .C(_12879_),
    .A(_12857_),
    .Y(_12880_));
 sg13g2_or4_1 _22002_ (.A(_12857_),
    .B(_12876_),
    .C(_12869_),
    .D(_12878_),
    .X(_12881_));
 sg13g2_nand3_1 _22003_ (.B(_12880_),
    .C(_12881_),
    .A(net85),
    .Y(_12882_));
 sg13g2_buf_1 _22004_ (.A(\grid.cell_29_0.s ),
    .X(_12883_));
 sg13g2_buf_1 _22005_ (.A(net1085),
    .X(_12884_));
 sg13g2_xnor2_1 _22006_ (.Y(_12885_),
    .A(_12884_),
    .B(_12877_));
 sg13g2_xor2_1 _22007_ (.B(_12885_),
    .A(_12861_),
    .X(_12886_));
 sg13g2_a21oi_1 _22008_ (.A1(net98),
    .A2(_12886_),
    .Y(_12887_),
    .B1(net802));
 sg13g2_nor2_1 _22009_ (.A(net37),
    .B(_12887_),
    .Y(_12888_));
 sg13g2_a22oi_1 _22010_ (.Y(_12889_),
    .B1(_12882_),
    .B2(_12888_),
    .A2(net37),
    .A1(net40));
 sg13g2_nor2_1 _22011_ (.A(net214),
    .B(_12889_),
    .Y(_00445_));
 sg13g2_buf_1 _22012_ (.A(net451),
    .X(_12890_));
 sg13g2_buf_2 _22013_ (.A(\grid.cell_29_1.se ),
    .X(_12891_));
 sg13g2_buf_2 _22014_ (.A(_12891_),
    .X(_12892_));
 sg13g2_inv_2 _22015_ (.Y(_12893_),
    .A(_12892_));
 sg13g2_nor2_1 _22016_ (.A(_12533_),
    .B(_12893_),
    .Y(_12894_));
 sg13g2_xnor2_1 _22017_ (.Y(_12895_),
    .A(_12516_),
    .B(_12891_));
 sg13g2_nor2_1 _22018_ (.A(net469),
    .B(_12894_),
    .Y(_12896_));
 sg13g2_a21oi_1 _22019_ (.A1(net469),
    .A2(_12895_),
    .Y(_12897_),
    .B1(_12896_));
 sg13g2_a22oi_1 _22020_ (.Y(_12898_),
    .B1(_12897_),
    .B2(net220),
    .A2(_12894_),
    .A1(_12241_));
 sg13g2_a21oi_1 _22021_ (.A1(_12183_),
    .A2(_12894_),
    .Y(_12899_),
    .B1(net211));
 sg13g2_a21oi_1 _22022_ (.A1(net211),
    .A2(_12898_),
    .Y(_12900_),
    .B1(_12899_));
 sg13g2_xnor2_1 _22023_ (.Y(_12901_),
    .A(_12891_),
    .B(_12545_));
 sg13g2_xor2_1 _22024_ (.B(_12901_),
    .A(_12858_),
    .X(_12902_));
 sg13g2_xor2_1 _22025_ (.B(net802),
    .A(net807),
    .X(_12903_));
 sg13g2_nor4_1 _22026_ (.A(net793),
    .B(net803),
    .C(_12902_),
    .D(_12903_),
    .Y(_12904_));
 sg13g2_xnor2_1 _22027_ (.Y(_12905_),
    .A(_12491_),
    .B(_12902_));
 sg13g2_o21ai_1 _22028_ (.B1(_12867_),
    .Y(_12906_),
    .A1(_12485_),
    .A2(_12902_));
 sg13g2_a21oi_1 _22029_ (.A1(_12865_),
    .A2(_12905_),
    .Y(_12907_),
    .B1(_12906_));
 sg13g2_buf_2 _22030_ (.A(net791),
    .X(_12908_));
 sg13g2_o21ai_1 _22031_ (.B1(_12183_),
    .Y(_12909_),
    .A1(net450),
    .A2(net812));
 sg13g2_nor2b_1 _22032_ (.A(_12239_),
    .B_N(_12891_),
    .Y(_12910_));
 sg13g2_nor2_1 _22033_ (.A(net791),
    .B(_12182_),
    .Y(_12911_));
 sg13g2_o21ai_1 _22034_ (.B1(net458),
    .Y(_12912_),
    .A1(_12910_),
    .A2(_12911_));
 sg13g2_o21ai_1 _22035_ (.B1(_12912_),
    .Y(_12913_),
    .A1(net458),
    .A2(_12909_));
 sg13g2_nand2b_1 _22036_ (.Y(_12914_),
    .B(_12240_),
    .A_N(net791));
 sg13g2_o21ai_1 _22037_ (.B1(_12914_),
    .Y(_12915_),
    .A1(net801),
    .A2(_12910_));
 sg13g2_o21ai_1 _22038_ (.B1(net801),
    .Y(_12916_),
    .A1(net791),
    .A2(_12240_));
 sg13g2_o21ai_1 _22039_ (.B1(_12916_),
    .Y(_12917_),
    .A1(_12893_),
    .A2(_12241_));
 sg13g2_a22oi_1 _22040_ (.Y(_12918_),
    .B1(_12917_),
    .B2(_12183_),
    .A2(_12915_),
    .A1(_12176_));
 sg13g2_nor2_1 _22041_ (.A(net791),
    .B(_12241_),
    .Y(_12919_));
 sg13g2_or3_1 _22042_ (.A(net795),
    .B(_12516_),
    .C(_12891_),
    .X(_12920_));
 sg13g2_nand4_1 _22043_ (.B(_12179_),
    .C(_12516_),
    .A(net795),
    .Y(_12921_),
    .D(net791));
 sg13g2_a21oi_1 _22044_ (.A1(_12920_),
    .A2(_12921_),
    .Y(_12922_),
    .B1(net816));
 sg13g2_a21oi_1 _22045_ (.A1(_12537_),
    .A2(_12919_),
    .Y(_12923_),
    .B1(_12922_));
 sg13g2_o21ai_1 _22046_ (.B1(_12923_),
    .Y(_12924_),
    .A1(net451),
    .A2(_12918_));
 sg13g2_a21oi_1 _22047_ (.A1(net211),
    .A2(_12913_),
    .Y(_12925_),
    .B1(_12924_));
 sg13g2_xor2_1 _22048_ (.B(_12925_),
    .A(_12907_),
    .X(_12926_));
 sg13g2_nor4_1 _22049_ (.A(net166),
    .B(_12900_),
    .C(_12904_),
    .D(_12926_),
    .Y(_12927_));
 sg13g2_nor2b_1 _22050_ (.A(net37),
    .B_N(_12454_),
    .Y(_12928_));
 sg13g2_o21ai_1 _22051_ (.B1(_12928_),
    .Y(_12929_),
    .A1(net75),
    .A2(_12927_));
 sg13g2_xnor2_1 _22052_ (.Y(_12930_),
    .A(_12491_),
    .B(net1085));
 sg13g2_xnor2_1 _22053_ (.Y(_12931_),
    .A(_12451_),
    .B(_12930_));
 sg13g2_xor2_1 _22054_ (.B(_12931_),
    .A(_12902_),
    .X(_12932_));
 sg13g2_nor2_1 _22055_ (.A(net37),
    .B(_12932_),
    .Y(_12933_));
 sg13g2_a22oi_1 _22056_ (.Y(_12934_),
    .B1(_12927_),
    .B2(_12933_),
    .A2(net37),
    .A1(net38));
 sg13g2_a21oi_1 _22057_ (.A1(_12929_),
    .A2(_12934_),
    .Y(_00446_),
    .B1(net523));
 sg13g2_nand2_2 _22058_ (.Y(_12935_),
    .A(net714),
    .B(_12828_));
 sg13g2_buf_1 _22059_ (.A(net450),
    .X(_12936_));
 sg13g2_buf_2 _22060_ (.A(\grid.cell_29_2.se ),
    .X(_12937_));
 sg13g2_buf_1 _22061_ (.A(_12937_),
    .X(_12938_));
 sg13g2_nand2_1 _22062_ (.Y(_12939_),
    .A(net1089),
    .B(net790));
 sg13g2_xor2_1 _22063_ (.B(net790),
    .A(net1089),
    .X(_12940_));
 sg13g2_nand2_1 _22064_ (.Y(_12941_),
    .A(_12179_),
    .B(_12940_));
 sg13g2_o21ai_1 _22065_ (.B1(_12941_),
    .Y(_12942_),
    .A1(_12180_),
    .A2(_12939_));
 sg13g2_nand2_1 _22066_ (.Y(_12943_),
    .A(net465),
    .B(_12942_));
 sg13g2_o21ai_1 _22067_ (.B1(_12943_),
    .Y(_12944_),
    .A1(_12277_),
    .A2(_12939_));
 sg13g2_nand2_1 _22068_ (.Y(_12945_),
    .A(_12180_),
    .B(net811));
 sg13g2_nor2_1 _22069_ (.A(net210),
    .B(_12945_),
    .Y(_12946_));
 sg13g2_inv_1 _22070_ (.Y(_12947_),
    .A(_12939_));
 sg13g2_buf_1 _22071_ (.A(_00274_),
    .X(_12948_));
 sg13g2_inv_1 _22072_ (.Y(_12949_),
    .A(_12948_));
 sg13g2_inv_1 _22073_ (.Y(_12950_),
    .A(net799));
 sg13g2_xor2_1 _22074_ (.B(_12577_),
    .A(_12937_),
    .X(_12951_));
 sg13g2_xnor2_1 _22075_ (.Y(_12952_),
    .A(_12175_),
    .B(_12891_));
 sg13g2_xnor2_1 _22076_ (.Y(_12953_),
    .A(_12951_),
    .B(_12952_));
 sg13g2_xnor2_1 _22077_ (.Y(_12954_),
    .A(net469),
    .B(net806));
 sg13g2_and4_1 _22078_ (.A(_12949_),
    .B(_12950_),
    .C(_12953_),
    .D(_12954_),
    .X(_12955_));
 sg13g2_a221oi_1 _22079_ (.B2(_12947_),
    .C1(_12955_),
    .B1(_12946_),
    .A1(net210),
    .Y(_12957_),
    .A2(_12944_));
 sg13g2_xor2_1 _22080_ (.B(_12953_),
    .A(net804),
    .X(_12958_));
 sg13g2_nand2b_1 _22081_ (.Y(_12959_),
    .B(_12948_),
    .A_N(_12099_));
 sg13g2_nor2b_1 _22082_ (.A(_12948_),
    .B_N(_12154_),
    .Y(_12960_));
 sg13g2_a221oi_1 _22083_ (.B2(_12959_),
    .C1(_12960_),
    .B1(_12958_),
    .A1(_12950_),
    .Y(_12961_),
    .A2(_12953_));
 sg13g2_buf_1 _22084_ (.A(net790),
    .X(_12962_));
 sg13g2_nor2_1 _22085_ (.A(net800),
    .B(net449),
    .Y(_12963_));
 sg13g2_o21ai_1 _22086_ (.B1(_12941_),
    .Y(_12964_),
    .A1(net811),
    .A2(_12947_));
 sg13g2_a22oi_1 _22087_ (.Y(_12965_),
    .B1(_12964_),
    .B2(_12277_),
    .A2(_12963_),
    .A1(_12945_));
 sg13g2_o21ai_1 _22088_ (.B1(net811),
    .Y(_12966_),
    .A1(_12176_),
    .A2(_12893_));
 sg13g2_nand3_1 _22089_ (.B(_12966_),
    .C(_12963_),
    .A(_12277_),
    .Y(_12968_));
 sg13g2_o21ai_1 _22090_ (.B1(_12968_),
    .Y(_12969_),
    .A1(net210),
    .A2(_12965_));
 sg13g2_xor2_1 _22091_ (.B(_12969_),
    .A(_12961_),
    .X(_12970_));
 sg13g2_a21oi_1 _22092_ (.A1(_12957_),
    .A2(_12970_),
    .Y(_12971_),
    .B1(net117));
 sg13g2_xnor2_1 _22093_ (.Y(_12972_),
    .A(_12858_),
    .B(_12958_));
 sg13g2_a21oi_1 _22094_ (.A1(net122),
    .A2(_12972_),
    .Y(_12973_),
    .B1(net215));
 sg13g2_nand2b_1 _22095_ (.Y(_12974_),
    .B(net1194),
    .A_N(_12828_));
 sg13g2_buf_1 _22096_ (.A(_12974_),
    .X(_12975_));
 sg13g2_or3_1 _22097_ (.A(_12971_),
    .B(_12973_),
    .C(_12975_),
    .X(_12976_));
 sg13g2_o21ai_1 _22098_ (.B1(_12976_),
    .Y(_00447_),
    .A1(net35),
    .A2(_12935_));
 sg13g2_buf_1 _22099_ (.A(_00273_),
    .X(_12978_));
 sg13g2_inv_2 _22100_ (.Y(_12979_),
    .A(_12978_));
 sg13g2_nor2_1 _22101_ (.A(_12212_),
    .B(_12979_),
    .Y(_12980_));
 sg13g2_buf_2 _22102_ (.A(\grid.cell_29_3.se ),
    .X(_12981_));
 sg13g2_xnor2_1 _22103_ (.Y(_12982_),
    .A(net1088),
    .B(net1084));
 sg13g2_buf_2 _22104_ (.A(_12982_),
    .X(_12983_));
 sg13g2_xnor2_1 _22105_ (.Y(_12984_),
    .A(_12273_),
    .B(_12983_));
 sg13g2_xnor2_1 _22106_ (.Y(_12985_),
    .A(net790),
    .B(_12984_));
 sg13g2_xnor2_1 _22107_ (.Y(_12986_),
    .A(net215),
    .B(_12985_));
 sg13g2_a22oi_1 _22108_ (.Y(_12987_),
    .B1(_12638_),
    .B2(_12985_),
    .A2(_12979_),
    .A1(net220));
 sg13g2_o21ai_1 _22109_ (.B1(_12987_),
    .Y(_12989_),
    .A1(_12980_),
    .A2(_12986_));
 sg13g2_nand2_2 _22110_ (.Y(_12990_),
    .A(net1088),
    .B(net1084));
 sg13g2_nor2_1 _22111_ (.A(_12583_),
    .B(_12983_),
    .Y(_12991_));
 sg13g2_a21oi_1 _22112_ (.A1(_12314_),
    .A2(_12990_),
    .Y(_12992_),
    .B1(_12991_));
 sg13g2_buf_1 _22113_ (.A(net1084),
    .X(_12993_));
 sg13g2_a21oi_1 _22114_ (.A1(_12229_),
    .A2(net790),
    .Y(_12994_),
    .B1(_12314_));
 sg13g2_or3_1 _22115_ (.A(net798),
    .B(net789),
    .C(_12994_),
    .X(_12995_));
 sg13g2_o21ai_1 _22116_ (.B1(_12995_),
    .Y(_12996_),
    .A1(net449),
    .A2(_12992_));
 sg13g2_nand2_1 _22117_ (.Y(_12997_),
    .A(net811),
    .B(net464));
 sg13g2_nor3_1 _22118_ (.A(net449),
    .B(net456),
    .C(net789),
    .Y(_12998_));
 sg13g2_a22oi_1 _22119_ (.Y(_13000_),
    .B1(_12997_),
    .B2(_12998_),
    .A2(_12996_),
    .A1(net1093));
 sg13g2_xor2_1 _22120_ (.B(_13000_),
    .A(_12989_),
    .X(_13001_));
 sg13g2_nor2_1 _22121_ (.A(_12252_),
    .B(_12990_),
    .Y(_13002_));
 sg13g2_o21ai_1 _22122_ (.B1(net219),
    .Y(_13003_),
    .A1(_12991_),
    .A2(_13002_));
 sg13g2_o21ai_1 _22123_ (.B1(_13003_),
    .Y(_13004_),
    .A1(net1093),
    .A2(_12990_));
 sg13g2_and2_1 _22124_ (.A(_12979_),
    .B(_12545_),
    .X(_13005_));
 sg13g2_and2_1 _22125_ (.A(_12638_),
    .B(_12985_),
    .X(_13006_));
 sg13g2_nor3_1 _22126_ (.A(net449),
    .B(_12990_),
    .C(_12997_),
    .Y(_13007_));
 sg13g2_a221oi_1 _22127_ (.B2(_13006_),
    .C1(_13007_),
    .B1(_13005_),
    .A1(net449),
    .Y(_13008_),
    .A2(_13004_));
 sg13g2_a21oi_1 _22128_ (.A1(_13001_),
    .A2(_13008_),
    .Y(_13009_),
    .B1(net96));
 sg13g2_xor2_1 _22129_ (.B(_12985_),
    .A(_12901_),
    .X(_13011_));
 sg13g2_a21oi_1 _22130_ (.A1(net68),
    .A2(_13011_),
    .Y(_13012_),
    .B1(net457));
 sg13g2_or3_1 _22131_ (.A(_12975_),
    .B(_13009_),
    .C(_13012_),
    .X(_13013_));
 sg13g2_o21ai_1 _22132_ (.B1(_13013_),
    .Y(_00448_),
    .A1(net32),
    .A2(_12935_));
 sg13g2_buf_2 _22133_ (.A(\grid.cell_29_4.se ),
    .X(_13014_));
 sg13g2_xor2_1 _22134_ (.B(_13014_),
    .A(_12652_),
    .X(_13015_));
 sg13g2_buf_1 _22135_ (.A(_13014_),
    .X(_13016_));
 sg13g2_nand2_1 _22136_ (.Y(_13017_),
    .A(net797),
    .B(net788));
 sg13g2_a22oi_1 _22137_ (.Y(_13018_),
    .B1(_13017_),
    .B2(_12301_),
    .A2(_13015_),
    .A1(net810));
 sg13g2_inv_2 _22138_ (.Y(_13019_),
    .A(_13014_));
 sg13g2_inv_1 _22139_ (.Y(_13021_),
    .A(net1084));
 sg13g2_o21ai_1 _22140_ (.B1(net809),
    .Y(_13022_),
    .A1(_12314_),
    .A2(_13021_));
 sg13g2_nand3b_1 _22141_ (.B(_13019_),
    .C(_13022_),
    .Y(_13023_),
    .A_N(net455));
 sg13g2_o21ai_1 _22142_ (.B1(_13023_),
    .Y(_13024_),
    .A1(net789),
    .A2(_13018_));
 sg13g2_buf_1 _22143_ (.A(net788),
    .X(_13025_));
 sg13g2_nor2_1 _22144_ (.A(_12314_),
    .B(_12301_),
    .Y(_13026_));
 sg13g2_nor4_1 _22145_ (.A(net789),
    .B(_12678_),
    .C(net448),
    .D(_13026_),
    .Y(_13027_));
 sg13g2_a21o_1 _22146_ (.A2(_13024_),
    .A1(_12357_),
    .B1(_13027_),
    .X(_13028_));
 sg13g2_buf_2 _22147_ (.A(_00063_),
    .X(_13029_));
 sg13g2_xnor2_1 _22148_ (.Y(_13030_),
    .A(_12266_),
    .B(net1084));
 sg13g2_xnor2_1 _22149_ (.Y(_13032_),
    .A(_13019_),
    .B(_12663_));
 sg13g2_xor2_1 _22150_ (.B(_13032_),
    .A(_13030_),
    .X(_13033_));
 sg13g2_buf_1 _22151_ (.A(_13033_),
    .X(_13034_));
 sg13g2_o21ai_1 _22152_ (.B1(_12583_),
    .Y(_13035_),
    .A1(net800),
    .A2(_13034_));
 sg13g2_a21o_1 _22153_ (.A2(_12583_),
    .A1(_12659_),
    .B1(_13034_),
    .X(_13036_));
 sg13g2_nor2_1 _22154_ (.A(_12583_),
    .B(net800),
    .Y(_13037_));
 sg13g2_a221oi_1 _22155_ (.B2(net457),
    .C1(_13037_),
    .B1(_13036_),
    .A1(_12658_),
    .Y(_13038_),
    .A2(_13035_));
 sg13g2_xnor2_1 _22156_ (.Y(_13039_),
    .A(net800),
    .B(_13034_));
 sg13g2_nor2_1 _22157_ (.A(_12658_),
    .B(_13034_),
    .Y(_13040_));
 sg13g2_a22oi_1 _22158_ (.Y(_13041_),
    .B1(_13040_),
    .B2(_13029_),
    .A2(_13039_),
    .A1(net465));
 sg13g2_o21ai_1 _22159_ (.B1(_13041_),
    .Y(_13043_),
    .A1(_13029_),
    .A2(_13038_));
 sg13g2_and2_1 _22160_ (.A(net455),
    .B(net788),
    .X(_13044_));
 sg13g2_buf_1 _22161_ (.A(_13044_),
    .X(_13045_));
 sg13g2_nand2_1 _22162_ (.Y(_13046_),
    .A(net810),
    .B(_13015_));
 sg13g2_o21ai_1 _22163_ (.B1(_13046_),
    .Y(_13047_),
    .A1(net464),
    .A2(_13017_));
 sg13g2_a22oi_1 _22164_ (.Y(_13048_),
    .B1(_13047_),
    .B2(net463),
    .A2(_13045_),
    .A1(_12696_));
 sg13g2_nand3_1 _22165_ (.B(_13045_),
    .C(_13026_),
    .A(_13021_),
    .Y(_13049_));
 sg13g2_o21ai_1 _22166_ (.B1(_13049_),
    .Y(_13050_),
    .A1(_13021_),
    .A2(_13048_));
 sg13g2_nor3_1 _22167_ (.A(_13028_),
    .B(_13040_),
    .C(_13050_),
    .Y(_13051_));
 sg13g2_inv_1 _22168_ (.Y(_13052_),
    .A(_13029_));
 sg13g2_a21o_1 _22169_ (.A2(_13039_),
    .A1(_12264_),
    .B1(_13052_),
    .X(_13054_));
 sg13g2_o21ai_1 _22170_ (.B1(_13054_),
    .Y(_13055_),
    .A1(net465),
    .A2(_13039_));
 sg13g2_a221oi_1 _22171_ (.B2(_13055_),
    .C1(net106),
    .B1(_13051_),
    .A1(_13028_),
    .Y(_13056_),
    .A2(_13043_));
 sg13g2_xnor2_1 _22172_ (.Y(_13057_),
    .A(_12951_),
    .B(_13034_));
 sg13g2_a21oi_1 _22173_ (.A1(net68),
    .A2(_13057_),
    .Y(_13058_),
    .B1(net456));
 sg13g2_or3_1 _22174_ (.A(_12975_),
    .B(_13056_),
    .C(_13058_),
    .X(_13059_));
 sg13g2_o21ai_1 _22175_ (.B1(_13059_),
    .Y(_00449_),
    .A1(net29),
    .A2(_12935_));
 sg13g2_buf_2 _22176_ (.A(\grid.cell_29_5.se ),
    .X(_13060_));
 sg13g2_xor2_1 _22177_ (.B(_13060_),
    .A(net796),
    .X(_13061_));
 sg13g2_buf_1 _22178_ (.A(_13060_),
    .X(_13062_));
 sg13g2_nand2_1 _22179_ (.Y(_13064_),
    .A(net796),
    .B(net787));
 sg13g2_buf_1 _22180_ (.A(_13064_),
    .X(_13065_));
 sg13g2_a22oi_1 _22181_ (.Y(_13066_),
    .B1(_13065_),
    .B2(_12382_),
    .A2(_13061_),
    .A1(net809));
 sg13g2_nand2_1 _22182_ (.Y(_13067_),
    .A(net809),
    .B(net788));
 sg13g2_or2_1 _22183_ (.X(_13068_),
    .B(net787),
    .A(_12700_));
 sg13g2_a21o_1 _22184_ (.A2(_13067_),
    .A1(_12341_),
    .B1(_13068_),
    .X(_13069_));
 sg13g2_o21ai_1 _22185_ (.B1(_13069_),
    .Y(_13070_),
    .A1(net448),
    .A2(_13066_));
 sg13g2_nand2_1 _22186_ (.Y(_13071_),
    .A(_12309_),
    .B(_12376_));
 sg13g2_nor2_1 _22187_ (.A(net448),
    .B(_13068_),
    .Y(_13072_));
 sg13g2_and2_1 _22188_ (.A(_13071_),
    .B(_13072_),
    .X(_13073_));
 sg13g2_a21oi_1 _22189_ (.A1(_12392_),
    .A2(_13070_),
    .Y(_13075_),
    .B1(_13073_));
 sg13g2_xor2_1 _22190_ (.B(_13014_),
    .A(_12617_),
    .X(_13076_));
 sg13g2_xnor2_1 _22191_ (.Y(_13077_),
    .A(_12699_),
    .B(_13060_));
 sg13g2_xnor2_1 _22192_ (.Y(_13078_),
    .A(_12335_),
    .B(_13077_));
 sg13g2_xnor2_1 _22193_ (.Y(_13079_),
    .A(_13076_),
    .B(_13078_));
 sg13g2_buf_2 _22194_ (.A(_13079_),
    .X(_13080_));
 sg13g2_nand2_1 _22195_ (.Y(_13081_),
    .A(net448),
    .B(_13078_));
 sg13g2_or2_1 _22196_ (.X(_13082_),
    .B(_13078_),
    .A(net788));
 sg13g2_a221oi_1 _22197_ (.B2(_13082_),
    .C1(net1087),
    .B1(_13081_),
    .A1(net464),
    .Y(_13083_),
    .A2(_13080_));
 sg13g2_xnor2_1 _22198_ (.Y(_13084_),
    .A(net448),
    .B(_13078_));
 sg13g2_a22oi_1 _22199_ (.Y(_13086_),
    .B1(_13084_),
    .B2(_12698_),
    .A2(_13080_),
    .A1(_12282_));
 sg13g2_buf_1 _22200_ (.A(_00095_),
    .X(_13087_));
 sg13g2_inv_1 _22201_ (.Y(_13088_),
    .A(_13087_));
 sg13g2_o21ai_1 _22202_ (.B1(_13088_),
    .Y(_13089_),
    .A1(_12282_),
    .A2(_13080_));
 sg13g2_mux2_1 _22203_ (.A0(_13083_),
    .A1(_13086_),
    .S(_13089_),
    .X(_13090_));
 sg13g2_nor2_1 _22204_ (.A(net219),
    .B(_13080_),
    .Y(_13091_));
 sg13g2_a21oi_1 _22205_ (.A1(net219),
    .A2(_13080_),
    .Y(_13092_),
    .B1(_13088_));
 sg13g2_a221oi_1 _22206_ (.B2(_12698_),
    .C1(_13073_),
    .B1(_13084_),
    .A1(_12392_),
    .Y(_13093_),
    .A2(_13070_));
 sg13g2_o21ai_1 _22207_ (.B1(_13093_),
    .Y(_13094_),
    .A1(_13091_),
    .A2(_13092_));
 sg13g2_o21ai_1 _22208_ (.B1(_13094_),
    .Y(_13095_),
    .A1(_13075_),
    .A2(_13090_));
 sg13g2_nor2_1 _22209_ (.A(_12301_),
    .B(_13077_),
    .Y(_13097_));
 sg13g2_nor2_1 _22210_ (.A(_12318_),
    .B(_13065_),
    .Y(_13098_));
 sg13g2_o21ai_1 _22211_ (.B1(_12387_),
    .Y(_13099_),
    .A1(_13097_),
    .A2(_13098_));
 sg13g2_o21ai_1 _22212_ (.B1(_13099_),
    .Y(_13100_),
    .A1(_12392_),
    .A2(_13065_));
 sg13g2_o21ai_1 _22213_ (.B1(_13019_),
    .Y(_13101_),
    .A1(_13065_),
    .A2(_13071_));
 sg13g2_o21ai_1 _22214_ (.B1(_13101_),
    .Y(_13102_),
    .A1(_13019_),
    .A2(_13100_));
 sg13g2_a21oi_1 _22215_ (.A1(_13095_),
    .A2(_13102_),
    .Y(_13103_),
    .B1(_11608_));
 sg13g2_buf_1 _22216_ (.A(net123),
    .X(_13104_));
 sg13g2_xnor2_1 _22217_ (.Y(_13105_),
    .A(_13030_),
    .B(_13080_));
 sg13g2_a21oi_1 _22218_ (.A1(net66),
    .A2(_13105_),
    .Y(_13106_),
    .B1(_12678_));
 sg13g2_or3_1 _22219_ (.A(_12975_),
    .B(_13103_),
    .C(_13106_),
    .X(_13107_));
 sg13g2_o21ai_1 _22220_ (.B1(_13107_),
    .Y(_00450_),
    .A1(net43),
    .A2(_12935_));
 sg13g2_buf_1 _22221_ (.A(net787),
    .X(_13108_));
 sg13g2_inv_1 _22222_ (.Y(_13109_),
    .A(net447));
 sg13g2_nand2_1 _22223_ (.Y(_13110_),
    .A(_13109_),
    .B(_12835_));
 sg13g2_buf_2 _22224_ (.A(net452),
    .X(_13111_));
 sg13g2_buf_2 _22225_ (.A(net447),
    .X(_13112_));
 sg13g2_a21oi_1 _22226_ (.A1(net459),
    .A2(net209),
    .Y(_13113_),
    .B1(net208));
 sg13g2_buf_2 _22227_ (.A(_00157_),
    .X(_13114_));
 sg13g2_o21ai_1 _22228_ (.B1(_13114_),
    .Y(_13115_),
    .A1(_12835_),
    .A2(_13113_));
 sg13g2_a21oi_1 _22229_ (.A1(_13110_),
    .A2(_13115_),
    .Y(_13117_),
    .B1(net217));
 sg13g2_nor2_1 _22230_ (.A(_13114_),
    .B(_12874_),
    .Y(_13118_));
 sg13g2_xnor2_1 _22231_ (.Y(_13119_),
    .A(_13114_),
    .B(net208));
 sg13g2_nand3_1 _22232_ (.B(net447),
    .C(_12874_),
    .A(_13114_),
    .Y(_13120_));
 sg13g2_nor2b_1 _22233_ (.A(_13118_),
    .B_N(_13120_),
    .Y(_13121_));
 sg13g2_o21ai_1 _22234_ (.B1(_13121_),
    .Y(_13122_),
    .A1(_12835_),
    .A2(_13119_));
 sg13g2_nor2_1 _22235_ (.A(_12382_),
    .B(net467),
    .Y(_13123_));
 sg13g2_nand4_1 _22236_ (.B(_12423_),
    .C(net216),
    .A(net208),
    .Y(_13124_),
    .D(net209));
 sg13g2_a21oi_1 _22237_ (.A1(_13110_),
    .A2(_13124_),
    .Y(_13125_),
    .B1(net218));
 sg13g2_a221oi_1 _22238_ (.B2(_13123_),
    .C1(_13125_),
    .B1(_13122_),
    .A1(net208),
    .Y(_13126_),
    .A2(_13118_));
 sg13g2_nand2b_1 _22239_ (.Y(_13128_),
    .B(_13126_),
    .A_N(_13117_));
 sg13g2_buf_1 _22240_ (.A(_00127_),
    .X(_13129_));
 sg13g2_inv_2 _22241_ (.Y(_13130_),
    .A(_13129_));
 sg13g2_xnor2_1 _22242_ (.Y(_13131_),
    .A(net808),
    .B(net787));
 sg13g2_xnor2_1 _22243_ (.Y(_13132_),
    .A(_12860_),
    .B(_13131_));
 sg13g2_xor2_1 _22244_ (.B(_13132_),
    .A(net213),
    .X(_13133_));
 sg13g2_o21ai_1 _22245_ (.B1(_13133_),
    .Y(_13134_),
    .A1(_13130_),
    .A2(net463));
 sg13g2_nand2b_1 _22246_ (.Y(_13135_),
    .B(_13132_),
    .A_N(_12756_));
 sg13g2_nand2_1 _22247_ (.Y(_13136_),
    .A(_13130_),
    .B(net463));
 sg13g2_nand3_1 _22248_ (.B(_13135_),
    .C(_13136_),
    .A(_13134_),
    .Y(_13137_));
 sg13g2_xor2_1 _22249_ (.B(_13137_),
    .A(_13128_),
    .X(_13139_));
 sg13g2_xor2_1 _22250_ (.B(_13132_),
    .A(_13032_),
    .X(_13140_));
 sg13g2_nor3_1 _22251_ (.A(_13129_),
    .B(_12663_),
    .C(_13135_),
    .Y(_13141_));
 sg13g2_a21oi_1 _22252_ (.A1(net459),
    .A2(net452),
    .Y(_13142_),
    .B1(_12376_));
 sg13g2_a21oi_1 _22253_ (.A1(net218),
    .A2(_12870_),
    .Y(_13143_),
    .B1(_13142_));
 sg13g2_a21oi_1 _22254_ (.A1(_12423_),
    .A2(_13143_),
    .Y(_13144_),
    .B1(_13118_));
 sg13g2_nor2_1 _22255_ (.A(_13109_),
    .B(_13144_),
    .Y(_13145_));
 sg13g2_nor3_1 _22256_ (.A(net208),
    .B(_12413_),
    .C(_12874_),
    .Y(_13146_));
 sg13g2_nor4_1 _22257_ (.A(net170),
    .B(_13141_),
    .C(_13145_),
    .D(_13146_),
    .Y(_13147_));
 sg13g2_o21ai_1 _22258_ (.B1(_13147_),
    .Y(_13148_),
    .A1(net136),
    .A2(_13140_));
 sg13g2_or2_1 _22259_ (.X(_13150_),
    .B(_13148_),
    .A(_13139_));
 sg13g2_a22oi_1 _22260_ (.Y(_13151_),
    .B1(net25),
    .B2(_12826_),
    .A2(net72),
    .A1(net136));
 sg13g2_a221oi_1 _22261_ (.B2(_13151_),
    .C1(net533),
    .B1(_13150_),
    .A1(net24),
    .Y(_00451_),
    .A2(_12826_));
 sg13g2_xnor2_1 _22262_ (.Y(_13152_),
    .A(net794),
    .B(_13077_));
 sg13g2_xnor2_1 _22263_ (.Y(_13153_),
    .A(_12393_),
    .B(_13152_));
 sg13g2_buf_1 _22264_ (.A(_13153_),
    .X(_13154_));
 sg13g2_nand2b_1 _22265_ (.Y(_13155_),
    .B(_13154_),
    .A_N(net803));
 sg13g2_o21ai_1 _22266_ (.B1(_13114_),
    .Y(_13156_),
    .A1(net808),
    .A2(net467));
 sg13g2_mux2_1 _22267_ (.A0(_13123_),
    .A1(_13156_),
    .S(_13152_),
    .X(_13157_));
 sg13g2_a21oi_1 _22268_ (.A1(net447),
    .A2(net453),
    .Y(_13158_),
    .B1(net454));
 sg13g2_a21oi_1 _22269_ (.A1(_13109_),
    .A2(_12859_),
    .Y(_13160_),
    .B1(_13158_));
 sg13g2_and2_1 _22270_ (.A(_13157_),
    .B(_13160_),
    .X(_13161_));
 sg13g2_nor2_1 _22271_ (.A(_13157_),
    .B(_13160_),
    .Y(_13162_));
 sg13g2_or2_1 _22272_ (.X(_13163_),
    .B(_13162_),
    .A(_13161_));
 sg13g2_and2_1 _22273_ (.A(_13155_),
    .B(_13163_),
    .X(_13164_));
 sg13g2_xnor2_1 _22274_ (.Y(_13165_),
    .A(net802),
    .B(_13154_));
 sg13g2_nand2b_1 _22275_ (.Y(_13166_),
    .B(net807),
    .A_N(_13165_));
 sg13g2_o21ai_1 _22276_ (.B1(_13166_),
    .Y(_13167_),
    .A1(_12866_),
    .A2(_13164_));
 sg13g2_nor2b_1 _22277_ (.A(net807),
    .B_N(_13165_),
    .Y(_13168_));
 sg13g2_nand2b_1 _22278_ (.Y(_13169_),
    .B(net802),
    .A_N(_12485_));
 sg13g2_o21ai_1 _22279_ (.B1(_13154_),
    .Y(_13171_),
    .A1(net807),
    .A2(_12486_));
 sg13g2_and3_1 _22280_ (.X(_13172_),
    .A(_12820_),
    .B(_12486_),
    .C(_13154_));
 sg13g2_a221oi_1 _22281_ (.B2(net802),
    .C1(_13172_),
    .B1(_13171_),
    .A1(net807),
    .Y(_13173_),
    .A2(_13169_));
 sg13g2_nor2_1 _22282_ (.A(net793),
    .B(_13173_),
    .Y(_13174_));
 sg13g2_mux2_1 _22283_ (.A0(_13168_),
    .A1(_13174_),
    .S(_13163_),
    .X(_13175_));
 sg13g2_xor2_1 _22284_ (.B(_13154_),
    .A(_12931_),
    .X(_13176_));
 sg13g2_a21oi_1 _22285_ (.A1(net123),
    .A2(_13176_),
    .Y(_13177_),
    .B1(net137));
 sg13g2_a21oi_1 _22286_ (.A1(_13166_),
    .A2(_13155_),
    .Y(_13178_),
    .B1(_13162_));
 sg13g2_nor4_1 _22287_ (.A(net37),
    .B(_13177_),
    .C(_13161_),
    .D(_13178_),
    .Y(_13179_));
 sg13g2_o21ai_1 _22288_ (.B1(_13179_),
    .Y(_13180_),
    .A1(_13167_),
    .A2(_13175_));
 sg13g2_a21oi_1 _22289_ (.A1(net137),
    .A2(net105),
    .Y(_13182_),
    .B1(net37));
 sg13g2_a21o_1 _22290_ (.A2(net37),
    .A1(net121),
    .B1(_13182_),
    .X(_13183_));
 sg13g2_a21oi_1 _22291_ (.A1(_13180_),
    .A2(_13183_),
    .Y(_00452_),
    .B1(net523));
 sg13g2_nand2b_1 _22292_ (.Y(_13184_),
    .B(_01913_),
    .A_N(_01870_));
 sg13g2_buf_1 _22293_ (.A(_13184_),
    .X(_13185_));
 sg13g2_or2_1 _22294_ (.X(_13186_),
    .B(_13185_),
    .A(_10239_));
 sg13g2_buf_1 _22295_ (.A(_13186_),
    .X(_13187_));
 sg13g2_buf_1 _22296_ (.A(\grid.cell_2_0.se ),
    .X(_13188_));
 sg13g2_buf_1 _22297_ (.A(net1083),
    .X(_13189_));
 sg13g2_buf_1 _22298_ (.A(_13189_),
    .X(_13190_));
 sg13g2_buf_2 _22299_ (.A(\grid.cell_2_0.sw ),
    .X(_13192_));
 sg13g2_buf_1 _22300_ (.A(_13192_),
    .X(_13193_));
 sg13g2_inv_2 _22301_ (.Y(_13194_),
    .A(_13193_));
 sg13g2_buf_1 _22302_ (.A(net785),
    .X(_13195_));
 sg13g2_nand2_1 _22303_ (.Y(_13196_),
    .A(net1044),
    .B(net445));
 sg13g2_nand2_1 _22304_ (.Y(_13197_),
    .A(_09184_),
    .B(_13196_));
 sg13g2_o21ai_1 _22305_ (.B1(_13197_),
    .Y(_13198_),
    .A1(net273),
    .A2(_13194_));
 sg13g2_nand2_1 _22306_ (.Y(_13199_),
    .A(_09180_),
    .B(_13194_));
 sg13g2_nor2_1 _22307_ (.A(_09180_),
    .B(net445),
    .Y(_13200_));
 sg13g2_o21ai_1 _22308_ (.B1(_02087_),
    .Y(_13201_),
    .A1(_09188_),
    .A2(_13200_));
 sg13g2_o21ai_1 _22309_ (.B1(_13201_),
    .Y(_13203_),
    .A1(net1047),
    .A2(_13199_));
 sg13g2_a21o_1 _22310_ (.A2(_13198_),
    .A1(net373),
    .B1(_13203_),
    .X(_13204_));
 sg13g2_nor2_1 _22311_ (.A(net1045),
    .B(net373),
    .Y(_13205_));
 sg13g2_mux2_1 _22312_ (.A0(net373),
    .A1(net1044),
    .S(_13194_),
    .X(_13206_));
 sg13g2_nor2_1 _22313_ (.A(net273),
    .B(_13196_),
    .Y(_13207_));
 sg13g2_a221oi_1 _22314_ (.B2(net270),
    .C1(_13207_),
    .B1(_13206_),
    .A1(_13199_),
    .Y(_13208_),
    .A2(_13205_));
 sg13g2_nand2_2 _22315_ (.Y(_13209_),
    .A(net1083),
    .B(net445));
 sg13g2_nor3_1 _22316_ (.A(_09191_),
    .B(net1044),
    .C(_13209_),
    .Y(_13210_));
 sg13g2_nor3_1 _22317_ (.A(net1083),
    .B(net373),
    .C(_13199_),
    .Y(_13211_));
 sg13g2_o21ai_1 _22318_ (.B1(net711),
    .Y(_13212_),
    .A1(_13210_),
    .A2(_13211_));
 sg13g2_o21ai_1 _22319_ (.B1(_13212_),
    .Y(_13214_),
    .A1(net446),
    .A2(_13208_));
 sg13g2_a21oi_1 _22320_ (.A1(net446),
    .A2(_13204_),
    .Y(_13215_),
    .B1(_13214_));
 sg13g2_buf_1 _22321_ (.A(_00271_),
    .X(_13216_));
 sg13g2_buf_1 _22322_ (.A(_13216_),
    .X(_13217_));
 sg13g2_nand2_1 _22323_ (.Y(_13218_),
    .A(_02183_),
    .B(net784));
 sg13g2_xor2_1 _22324_ (.B(net1083),
    .A(_02076_),
    .X(_13219_));
 sg13g2_xnor2_1 _22325_ (.Y(_13220_),
    .A(net896),
    .B(_13192_));
 sg13g2_xor2_1 _22326_ (.B(_13220_),
    .A(_13219_),
    .X(_13221_));
 sg13g2_xnor2_1 _22327_ (.Y(_13222_),
    .A(net373),
    .B(_13221_));
 sg13g2_xnor2_1 _22328_ (.Y(_13223_),
    .A(net552),
    .B(_13222_));
 sg13g2_nand2b_1 _22329_ (.Y(_13225_),
    .B(net708),
    .A_N(net784));
 sg13g2_o21ai_1 _22330_ (.B1(_13225_),
    .Y(_13226_),
    .A1(net1125),
    .A2(_13222_));
 sg13g2_a21oi_1 _22331_ (.A1(_13218_),
    .A2(_13223_),
    .Y(_13227_),
    .B1(_13226_));
 sg13g2_xor2_1 _22332_ (.B(_13227_),
    .A(_13215_),
    .X(_13228_));
 sg13g2_buf_2 _22333_ (.A(\grid.cell_2_0.s ),
    .X(_13229_));
 sg13g2_inv_2 _22334_ (.Y(_13230_),
    .A(_13229_));
 sg13g2_xnor2_1 _22335_ (.Y(_13231_),
    .A(_02464_),
    .B(net552));
 sg13g2_xnor2_1 _22336_ (.Y(_13232_),
    .A(_13230_),
    .B(_13231_));
 sg13g2_xnor2_1 _22337_ (.Y(_13233_),
    .A(_13222_),
    .B(_13232_));
 sg13g2_nor2b_1 _22338_ (.A(net784),
    .B_N(_13231_),
    .Y(_13234_));
 sg13g2_nor2_1 _22339_ (.A(net1125),
    .B(_13222_),
    .Y(_13236_));
 sg13g2_inv_1 _22340_ (.Y(_13237_),
    .A(_13188_));
 sg13g2_buf_1 _22341_ (.A(_13237_),
    .X(_13238_));
 sg13g2_nand2_1 _22342_ (.Y(_13239_),
    .A(_09185_),
    .B(net445));
 sg13g2_nand2b_1 _22343_ (.Y(_13240_),
    .B(_02151_),
    .A_N(_13220_));
 sg13g2_o21ai_1 _22344_ (.B1(_13240_),
    .Y(_13241_),
    .A1(net711),
    .A2(_13239_));
 sg13g2_nor2_1 _22345_ (.A(net1047),
    .B(_13239_),
    .Y(_13242_));
 sg13g2_a21oi_1 _22346_ (.A1(net174),
    .A2(_13241_),
    .Y(_13243_),
    .B1(_13242_));
 sg13g2_buf_1 _22347_ (.A(net445),
    .X(_13244_));
 sg13g2_nor3_1 _22348_ (.A(_02087_),
    .B(net786),
    .C(_09222_),
    .Y(_13245_));
 sg13g2_a21oi_1 _22349_ (.A1(net207),
    .A2(_13245_),
    .Y(_13247_),
    .B1(_05130_));
 sg13g2_o21ai_1 _22350_ (.B1(_13247_),
    .Y(_13248_),
    .A1(net444),
    .A2(_13243_));
 sg13g2_a221oi_1 _22351_ (.B2(_13236_),
    .C1(_13248_),
    .B1(_13234_),
    .A1(net892),
    .Y(_13249_),
    .A2(_13233_));
 sg13g2_a22oi_1 _22352_ (.Y(_13250_),
    .B1(_13228_),
    .B2(_13249_),
    .A2(net67),
    .A1(_09266_));
 sg13g2_o21ai_1 _22353_ (.B1(net522),
    .Y(_13251_),
    .A1(net40),
    .A2(net53));
 sg13g2_a21oi_1 _22354_ (.A1(net53),
    .A2(_13250_),
    .Y(_00453_),
    .B1(_13251_));
 sg13g2_buf_8 _22355_ (.A(\grid.cell_2_1.se ),
    .X(_13252_));
 sg13g2_xnor2_1 _22356_ (.Y(_13253_),
    .A(_03185_),
    .B(_13252_));
 sg13g2_xor2_1 _22357_ (.B(_13253_),
    .A(_13219_),
    .X(_13254_));
 sg13g2_xnor2_1 _22358_ (.Y(_13255_),
    .A(net891),
    .B(_13254_));
 sg13g2_buf_2 _22359_ (.A(_13255_),
    .X(_13257_));
 sg13g2_xnor2_1 _22360_ (.Y(_13258_),
    .A(net892),
    .B(_13257_));
 sg13g2_nand2_1 _22361_ (.Y(_13259_),
    .A(net708),
    .B(_13258_));
 sg13g2_buf_1 _22362_ (.A(_13252_),
    .X(_13260_));
 sg13g2_nand2_1 _22363_ (.Y(_13261_),
    .A(_02076_),
    .B(_03185_));
 sg13g2_nand2b_1 _22364_ (.Y(_13262_),
    .B(_13252_),
    .A_N(_02097_));
 sg13g2_o21ai_1 _22365_ (.B1(_13262_),
    .Y(_13263_),
    .A1(net783),
    .A2(_13261_));
 sg13g2_inv_2 _22366_ (.Y(_13264_),
    .A(_13260_));
 sg13g2_nand2_1 _22367_ (.Y(_13265_),
    .A(_13264_),
    .B(net1044));
 sg13g2_nor2_1 _22368_ (.A(net1126),
    .B(_13261_),
    .Y(_13266_));
 sg13g2_a221oi_1 _22369_ (.B2(_13266_),
    .C1(_13237_),
    .B1(_13265_),
    .A1(_09238_),
    .Y(_13268_),
    .A2(_13263_));
 sg13g2_nor2b_1 _22370_ (.A(net783),
    .B_N(_02097_),
    .Y(_13269_));
 sg13g2_a21o_1 _22371_ (.A2(_13262_),
    .A1(_09279_),
    .B1(_13269_),
    .X(_13270_));
 sg13g2_o21ai_1 _22372_ (.B1(net1126),
    .Y(_13271_),
    .A1(net783),
    .A2(_02097_));
 sg13g2_o21ai_1 _22373_ (.B1(_13271_),
    .Y(_13272_),
    .A1(_13264_),
    .A2(net1044));
 sg13g2_inv_1 _22374_ (.Y(_13273_),
    .A(_13261_));
 sg13g2_a221oi_1 _22375_ (.B2(_13273_),
    .C1(net1083),
    .B1(_13272_),
    .A1(net701),
    .Y(_13274_),
    .A2(_13270_));
 sg13g2_nand2_1 _22376_ (.Y(_13275_),
    .A(net1083),
    .B(_13252_));
 sg13g2_buf_2 _22377_ (.A(_13275_),
    .X(_13276_));
 sg13g2_or3_1 _22378_ (.A(net1083),
    .B(net1126),
    .C(net783),
    .X(_13277_));
 sg13g2_o21ai_1 _22379_ (.B1(_13277_),
    .Y(_13279_),
    .A1(_09273_),
    .A2(_13276_));
 sg13g2_a22oi_1 _22380_ (.Y(_13280_),
    .B1(_13269_),
    .B2(_09252_),
    .A2(_13279_),
    .A1(_02087_));
 sg13g2_o21ai_1 _22381_ (.B1(_13280_),
    .Y(_13281_),
    .A1(_13268_),
    .A2(_13274_));
 sg13g2_buf_1 _22382_ (.A(_13281_),
    .X(_13282_));
 sg13g2_o21ai_1 _22383_ (.B1(net1040),
    .Y(_13283_),
    .A1(net892),
    .A2(net1127));
 sg13g2_o21ai_1 _22384_ (.B1(_13283_),
    .Y(_13284_),
    .A1(net892),
    .A2(_13257_));
 sg13g2_nand3_1 _22385_ (.B(net1127),
    .C(_13257_),
    .A(net892),
    .Y(_13285_));
 sg13g2_nand2b_1 _22386_ (.Y(_13286_),
    .B(_13285_),
    .A_N(_13284_));
 sg13g2_nand3b_1 _22387_ (.B(_13282_),
    .C(_13286_),
    .Y(_13287_),
    .A_N(net784));
 sg13g2_nand2b_1 _22388_ (.Y(_13288_),
    .B(_13257_),
    .A_N(net1127));
 sg13g2_nand2_1 _22389_ (.Y(_13290_),
    .A(_13282_),
    .B(_13288_));
 sg13g2_nand2_1 _22390_ (.Y(_13291_),
    .A(net784),
    .B(_13290_));
 sg13g2_nand2_1 _22391_ (.Y(_13292_),
    .A(net890),
    .B(_13257_));
 sg13g2_a21oi_1 _22392_ (.A1(net1127),
    .A2(_13282_),
    .Y(_13293_),
    .B1(_13292_));
 sg13g2_nor3_1 _22393_ (.A(net890),
    .B(_13257_),
    .C(_13282_),
    .Y(_13294_));
 sg13g2_o21ai_1 _22394_ (.B1(_02183_),
    .Y(_13295_),
    .A1(_13293_),
    .A2(_13294_));
 sg13g2_nand4_1 _22395_ (.B(_13287_),
    .C(_13291_),
    .A(_13259_),
    .Y(_13296_),
    .D(_13295_));
 sg13g2_a21oi_1 _22396_ (.A1(_13259_),
    .A2(_13288_),
    .Y(_13297_),
    .B1(_13282_));
 sg13g2_buf_1 _22397_ (.A(_13260_),
    .X(_13298_));
 sg13g2_buf_1 _22398_ (.A(net443),
    .X(_13299_));
 sg13g2_nand3_1 _22399_ (.B(net444),
    .C(net206),
    .A(net711),
    .Y(_13301_));
 sg13g2_o21ai_1 _22400_ (.B1(_05267_),
    .Y(_13302_),
    .A1(_09273_),
    .A2(_13301_));
 sg13g2_nor2_1 _22401_ (.A(_09280_),
    .B(_13264_),
    .Y(_13303_));
 sg13g2_xor2_1 _22402_ (.B(_13252_),
    .A(_09237_),
    .X(_13304_));
 sg13g2_mux2_1 _22403_ (.A0(_13303_),
    .A1(_13304_),
    .S(_02151_),
    .X(_13305_));
 sg13g2_a22oi_1 _22404_ (.Y(_13306_),
    .B1(_13305_),
    .B2(net369),
    .A2(_13303_),
    .A1(_02302_));
 sg13g2_nor2_1 _22405_ (.A(net444),
    .B(_13306_),
    .Y(_13307_));
 sg13g2_xnor2_1 _22406_ (.Y(_13308_),
    .A(_09216_),
    .B(_13229_));
 sg13g2_xnor2_1 _22407_ (.Y(_13309_),
    .A(_02464_),
    .B(_13308_));
 sg13g2_xor2_1 _22408_ (.B(_13309_),
    .A(_13257_),
    .X(_13310_));
 sg13g2_nor2_1 _22409_ (.A(net271),
    .B(_13310_),
    .Y(_00607_));
 sg13g2_nor4_1 _22410_ (.A(_13297_),
    .B(_13302_),
    .C(_13307_),
    .D(_00607_),
    .Y(_00608_));
 sg13g2_a22oi_1 _22411_ (.Y(_00609_),
    .B1(_13296_),
    .B2(_00608_),
    .A2(net67),
    .A1(_09197_));
 sg13g2_o21ai_1 _22412_ (.B1(_10237_),
    .Y(_00610_),
    .A1(_11113_),
    .A2(net53));
 sg13g2_a21oi_1 _22413_ (.A1(net53),
    .A2(_00609_),
    .Y(_00454_),
    .B1(_00610_));
 sg13g2_nor2_1 _22414_ (.A(_10239_),
    .B(_13185_),
    .Y(_00611_));
 sg13g2_nand2_1 _22415_ (.Y(_00612_),
    .A(net33),
    .B(_00611_));
 sg13g2_buf_2 _22416_ (.A(\grid.cell_2_2.se ),
    .X(_00613_));
 sg13g2_buf_1 _22417_ (.A(_00613_),
    .X(_00614_));
 sg13g2_xor2_1 _22418_ (.B(_09305_),
    .A(net782),
    .X(_00615_));
 sg13g2_xnor2_1 _22419_ (.Y(_00617_),
    .A(_13253_),
    .B(_00615_));
 sg13g2_nand2_1 _22420_ (.Y(_00618_),
    .A(_09289_),
    .B(_00617_));
 sg13g2_buf_1 _22421_ (.A(_00270_),
    .X(_00619_));
 sg13g2_xnor2_1 _22422_ (.Y(_00620_),
    .A(_09291_),
    .B(_00613_));
 sg13g2_xnor2_1 _22423_ (.Y(_00621_),
    .A(net895),
    .B(net1029));
 sg13g2_xnor2_1 _22424_ (.Y(_00622_),
    .A(_00620_),
    .B(_00621_));
 sg13g2_xnor2_1 _22425_ (.Y(_00623_),
    .A(_13253_),
    .B(_00622_));
 sg13g2_buf_1 _22426_ (.A(_00623_),
    .X(_00624_));
 sg13g2_nor2_1 _22427_ (.A(net1082),
    .B(_00624_),
    .Y(_00625_));
 sg13g2_buf_1 _22428_ (.A(net1082),
    .X(_00626_));
 sg13g2_a21oi_1 _22429_ (.A1(_09289_),
    .A2(_00617_),
    .Y(_00628_),
    .B1(net781));
 sg13g2_nand2b_1 _22430_ (.Y(_00629_),
    .B(_00624_),
    .A_N(_00628_));
 sg13g2_a21oi_1 _22431_ (.A1(_02087_),
    .A2(_00624_),
    .Y(_00630_),
    .B1(net781));
 sg13g2_nor2_1 _22432_ (.A(_00618_),
    .B(_00630_),
    .Y(_00631_));
 sg13g2_a221oi_1 _22433_ (.B2(_02162_),
    .C1(_00631_),
    .B1(_00629_),
    .A1(_00618_),
    .Y(_00632_),
    .A2(_00625_));
 sg13g2_nand2_1 _22434_ (.Y(_00633_),
    .A(net889),
    .B(net782));
 sg13g2_nor2_1 _22435_ (.A(_03682_),
    .B(_00620_),
    .Y(_00634_));
 sg13g2_nor2_1 _22436_ (.A(_03337_),
    .B(_00633_),
    .Y(_00635_));
 sg13g2_o21ai_1 _22437_ (.B1(net366),
    .Y(_00636_),
    .A1(_00634_),
    .A2(_00635_));
 sg13g2_o21ai_1 _22438_ (.B1(_00636_),
    .Y(_00637_),
    .A1(_04440_),
    .A2(_00633_));
 sg13g2_nand2_1 _22439_ (.Y(_00638_),
    .A(_03337_),
    .B(net699));
 sg13g2_nor3_1 _22440_ (.A(net206),
    .B(_00638_),
    .C(_00633_),
    .Y(_00639_));
 sg13g2_a21oi_1 _22441_ (.A1(net206),
    .A2(_00637_),
    .Y(_00640_),
    .B1(_00639_));
 sg13g2_nand2_1 _22442_ (.Y(_00641_),
    .A(net781),
    .B(_00624_));
 sg13g2_o21ai_1 _22443_ (.B1(_00641_),
    .Y(_00642_),
    .A1(_02162_),
    .A2(_00625_));
 sg13g2_nand3_1 _22444_ (.B(_00640_),
    .C(_00642_),
    .A(_00618_),
    .Y(_00643_));
 sg13g2_buf_1 _22445_ (.A(net782),
    .X(_00644_));
 sg13g2_a21oi_1 _22446_ (.A1(_03380_),
    .A2(net443),
    .Y(_00645_),
    .B1(_04236_));
 sg13g2_nor4_1 _22447_ (.A(_09313_),
    .B(_09343_),
    .C(net442),
    .D(_00645_),
    .Y(_00646_));
 sg13g2_buf_1 _22448_ (.A(net782),
    .X(_00647_));
 sg13g2_inv_1 _22449_ (.Y(_00649_),
    .A(net441));
 sg13g2_nand3_1 _22450_ (.B(_00649_),
    .C(_00638_),
    .A(net269),
    .Y(_00650_));
 sg13g2_a21oi_1 _22451_ (.A1(net889),
    .A2(net441),
    .Y(_00651_),
    .B1(net699));
 sg13g2_o21ai_1 _22452_ (.B1(_04440_),
    .Y(_00652_),
    .A1(_00634_),
    .A2(_00651_));
 sg13g2_a21oi_1 _22453_ (.A1(_00650_),
    .A2(_00652_),
    .Y(_00653_),
    .B1(net206));
 sg13g2_nor2_1 _22454_ (.A(_00646_),
    .B(_00653_),
    .Y(_00654_));
 sg13g2_mux2_1 _22455_ (.A0(_00632_),
    .A1(_00643_),
    .S(_00654_),
    .X(_00655_));
 sg13g2_xor2_1 _22456_ (.B(_00624_),
    .A(_13219_),
    .X(_00656_));
 sg13g2_o21ai_1 _22457_ (.B1(net550),
    .Y(_00657_),
    .A1(net166),
    .A2(_00656_));
 sg13g2_nand2_1 _22458_ (.Y(_00658_),
    .A(_13187_),
    .B(_00657_));
 sg13g2_a21o_1 _22459_ (.A2(_00655_),
    .A1(net78),
    .B1(_00658_),
    .X(_00660_));
 sg13g2_buf_1 _22460_ (.A(_06110_),
    .X(_00661_));
 sg13g2_a21oi_1 _22461_ (.A1(_00612_),
    .A2(_00660_),
    .Y(_00455_),
    .B1(net440));
 sg13g2_nand2_1 _22462_ (.Y(_00662_),
    .A(net716),
    .B(_00611_));
 sg13g2_nor2_1 _22463_ (.A(net696),
    .B(_04236_),
    .Y(_00663_));
 sg13g2_buf_2 _22464_ (.A(\grid.cell_2_3.se ),
    .X(_00664_));
 sg13g2_buf_1 _22465_ (.A(_00664_),
    .X(_00665_));
 sg13g2_or3_1 _22466_ (.A(net888),
    .B(net441),
    .C(net780),
    .X(_00666_));
 sg13g2_a21oi_1 _22467_ (.A1(net888),
    .A2(_04217_),
    .Y(_00667_),
    .B1(_04712_));
 sg13g2_nor3_1 _22468_ (.A(net441),
    .B(net780),
    .C(_00667_),
    .Y(_00668_));
 sg13g2_xor2_1 _22469_ (.B(_00664_),
    .A(_00613_),
    .X(_00670_));
 sg13g2_nand2_1 _22470_ (.Y(_00671_),
    .A(net699),
    .B(_00670_));
 sg13g2_nand2_1 _22471_ (.Y(_00672_),
    .A(net782),
    .B(_00665_));
 sg13g2_buf_2 _22472_ (.A(_00672_),
    .X(_00673_));
 sg13g2_nand2_1 _22473_ (.Y(_00674_),
    .A(_04712_),
    .B(_00673_));
 sg13g2_a21oi_1 _22474_ (.A1(_00671_),
    .A2(_00674_),
    .Y(_00675_),
    .B1(net888));
 sg13g2_o21ai_1 _22475_ (.B1(_04870_),
    .Y(_00676_),
    .A1(_00668_),
    .A2(_00675_));
 sg13g2_o21ai_1 _22476_ (.B1(_00676_),
    .Y(_00677_),
    .A1(_00663_),
    .A2(_00666_));
 sg13g2_buf_2 _22477_ (.A(_00269_),
    .X(_00678_));
 sg13g2_nand2_1 _22478_ (.Y(_00679_),
    .A(net268),
    .B(net1124));
 sg13g2_nor2_1 _22479_ (.A(net268),
    .B(net1124),
    .Y(_00681_));
 sg13g2_xnor2_1 _22480_ (.Y(_00682_),
    .A(_04705_),
    .B(_09334_));
 sg13g2_xor2_1 _22481_ (.B(_00682_),
    .A(_00670_),
    .X(_00683_));
 sg13g2_xnor2_1 _22482_ (.Y(_00684_),
    .A(_04206_),
    .B(_00683_));
 sg13g2_nand2_1 _22483_ (.Y(_00685_),
    .A(_03682_),
    .B(_09348_));
 sg13g2_a21oi_1 _22484_ (.A1(_00684_),
    .A2(_00685_),
    .Y(_00686_),
    .B1(net550));
 sg13g2_a221oi_1 _22485_ (.B2(_00684_),
    .C1(_00686_),
    .B1(_00681_),
    .A1(net369),
    .Y(_00687_),
    .A2(_00679_));
 sg13g2_xnor2_1 _22486_ (.Y(_00688_),
    .A(_09279_),
    .B(_00684_));
 sg13g2_and2_1 _22487_ (.A(net1124),
    .B(_00684_),
    .X(_00689_));
 sg13g2_a22oi_1 _22488_ (.Y(_00690_),
    .B1(_00689_),
    .B2(_00678_),
    .A2(_00688_),
    .A1(net369));
 sg13g2_o21ai_1 _22489_ (.B1(_00690_),
    .Y(_00692_),
    .A1(_00678_),
    .A2(_00687_));
 sg13g2_o21ai_1 _22490_ (.B1(_00671_),
    .Y(_00693_),
    .A1(_04495_),
    .A2(_00673_));
 sg13g2_nor3_1 _22491_ (.A(net548),
    .B(_04236_),
    .C(_00673_),
    .Y(_00694_));
 sg13g2_a21oi_1 _22492_ (.A1(net548),
    .A2(_00693_),
    .Y(_00695_),
    .B1(_00694_));
 sg13g2_nor2_1 _22493_ (.A(net696),
    .B(_00695_),
    .Y(_00696_));
 sg13g2_nor3_1 _22494_ (.A(_04870_),
    .B(_09336_),
    .C(_00673_),
    .Y(_00697_));
 sg13g2_nor4_1 _22495_ (.A(_00677_),
    .B(_00696_),
    .C(_00689_),
    .D(_00697_),
    .Y(_00698_));
 sg13g2_inv_1 _22496_ (.Y(_00699_),
    .A(_00678_));
 sg13g2_a21o_1 _22497_ (.A2(_00688_),
    .A1(_00699_),
    .B1(_03756_),
    .X(_00700_));
 sg13g2_o21ai_1 _22498_ (.B1(_00700_),
    .Y(_00701_),
    .A1(_00699_),
    .A2(_00688_));
 sg13g2_a22oi_1 _22499_ (.Y(_00703_),
    .B1(_00698_),
    .B2(_00701_),
    .A2(_00692_),
    .A1(_00677_));
 sg13g2_xnor2_1 _22500_ (.Y(_00704_),
    .A(_13253_),
    .B(_00688_));
 sg13g2_a21oi_1 _22501_ (.A1(net123),
    .A2(_00704_),
    .Y(_00705_),
    .B1(_09313_));
 sg13g2_nand2_1 _22502_ (.Y(_00706_),
    .A(_12967_),
    .B(net53));
 sg13g2_or2_1 _22503_ (.X(_00707_),
    .B(_00706_),
    .A(_00705_));
 sg13g2_a21o_1 _22504_ (.A2(_00703_),
    .A1(net78),
    .B1(_00707_),
    .X(_00708_));
 sg13g2_o21ai_1 _22505_ (.B1(_00708_),
    .Y(_00456_),
    .A1(net32),
    .A2(_00662_));
 sg13g2_buf_2 _22506_ (.A(\grid.cell_2_4.se ),
    .X(_00709_));
 sg13g2_buf_1 _22507_ (.A(_00709_),
    .X(_00710_));
 sg13g2_nand2_2 _22508_ (.Y(_00711_),
    .A(net780),
    .B(net779));
 sg13g2_xor2_1 _22509_ (.B(_00709_),
    .A(_00664_),
    .X(_00713_));
 sg13g2_nand2_1 _22510_ (.Y(_00714_),
    .A(net1026),
    .B(_00713_));
 sg13g2_o21ai_1 _22511_ (.B1(_00714_),
    .Y(_00715_),
    .A1(_04885_),
    .A2(_00711_));
 sg13g2_nor2_1 _22512_ (.A(_09381_),
    .B(net696),
    .Y(_00716_));
 sg13g2_inv_1 _22513_ (.Y(_00717_),
    .A(net780));
 sg13g2_inv_2 _22514_ (.Y(_00718_),
    .A(net779));
 sg13g2_nor2_1 _22515_ (.A(net439),
    .B(_00718_),
    .Y(_00719_));
 sg13g2_a22oi_1 _22516_ (.Y(_00720_),
    .B1(_00716_),
    .B2(_00719_),
    .A2(_00715_),
    .A1(net267));
 sg13g2_nor2_1 _22517_ (.A(net691),
    .B(_00720_),
    .Y(_00721_));
 sg13g2_nor3_1 _22518_ (.A(_04970_),
    .B(_09413_),
    .C(_00711_),
    .Y(_00722_));
 sg13g2_buf_1 _22519_ (.A(_00034_),
    .X(_00724_));
 sg13g2_xnor2_1 _22520_ (.Y(_00725_),
    .A(_04943_),
    .B(_09370_));
 sg13g2_xor2_1 _22521_ (.B(_00725_),
    .A(_00713_),
    .X(_00726_));
 sg13g2_xnor2_1 _22522_ (.Y(_00727_),
    .A(_04712_),
    .B(_00726_));
 sg13g2_nor4_1 _22523_ (.A(_09382_),
    .B(_00724_),
    .C(_09305_),
    .D(_00727_),
    .Y(_00728_));
 sg13g2_a22oi_1 _22524_ (.Y(_00729_),
    .B1(_00711_),
    .B2(net691),
    .A2(_00713_),
    .A1(_04884_));
 sg13g2_o21ai_1 _22525_ (.B1(net1025),
    .Y(_00730_),
    .A1(_09413_),
    .A2(_04721_));
 sg13g2_nand3_1 _22526_ (.B(_00718_),
    .C(_00730_),
    .A(net439),
    .Y(_00731_));
 sg13g2_o21ai_1 _22527_ (.B1(_00731_),
    .Y(_00732_),
    .A1(_09373_),
    .A2(_00729_));
 sg13g2_nand2_1 _22528_ (.Y(_00733_),
    .A(net692),
    .B(net693));
 sg13g2_buf_1 _22529_ (.A(net780),
    .X(_00735_));
 sg13g2_buf_1 _22530_ (.A(net779),
    .X(_00736_));
 sg13g2_nor3_1 _22531_ (.A(_09373_),
    .B(net438),
    .C(net437),
    .Y(_00737_));
 sg13g2_a22oi_1 _22532_ (.Y(_00738_),
    .B1(_00733_),
    .B2(_00737_),
    .A2(_00732_),
    .A1(_04970_));
 sg13g2_nand2_1 _22533_ (.Y(_00739_),
    .A(_00724_),
    .B(_04236_));
 sg13g2_xnor2_1 _22534_ (.Y(_00740_),
    .A(net549),
    .B(_00727_));
 sg13g2_inv_1 _22535_ (.Y(_00741_),
    .A(_00724_));
 sg13g2_nand2_1 _22536_ (.Y(_00742_),
    .A(_00741_),
    .B(net366));
 sg13g2_o21ai_1 _22537_ (.B1(_00742_),
    .Y(_00743_),
    .A1(_09382_),
    .A2(_00727_));
 sg13g2_a21oi_1 _22538_ (.A1(_00739_),
    .A2(_00740_),
    .Y(_00744_),
    .B1(_00743_));
 sg13g2_xor2_1 _22539_ (.B(_00744_),
    .A(_00738_),
    .X(_00746_));
 sg13g2_nor4_1 _22540_ (.A(_00721_),
    .B(_00722_),
    .C(_00728_),
    .D(_00746_),
    .Y(_00747_));
 sg13g2_xnor2_1 _22541_ (.Y(_00748_),
    .A(_00615_),
    .B(_00727_));
 sg13g2_a21oi_1 _22542_ (.A1(net114),
    .A2(_00748_),
    .Y(_00749_),
    .B1(_09358_));
 sg13g2_nor2_1 _22543_ (.A(_00706_),
    .B(_00749_),
    .Y(_00750_));
 sg13g2_o21ai_1 _22544_ (.B1(_00750_),
    .Y(_00751_),
    .A1(net81),
    .A2(_00747_));
 sg13g2_o21ai_1 _22545_ (.B1(_00751_),
    .Y(_00457_),
    .A1(net29),
    .A2(_00662_));
 sg13g2_buf_1 _22546_ (.A(\grid.cell_2_5.se ),
    .X(_00752_));
 sg13g2_buf_1 _22547_ (.A(_00752_),
    .X(_00753_));
 sg13g2_nand2_1 _22548_ (.Y(_00754_),
    .A(_00710_),
    .B(net778));
 sg13g2_buf_1 _22549_ (.A(_00754_),
    .X(_00756_));
 sg13g2_xor2_1 _22550_ (.B(_00752_),
    .A(_00709_),
    .X(_00757_));
 sg13g2_nand2_1 _22551_ (.Y(_00758_),
    .A(net1025),
    .B(_00757_));
 sg13g2_o21ai_1 _22552_ (.B1(_00758_),
    .Y(_00759_),
    .A1(_04944_),
    .A2(_00756_));
 sg13g2_nand2_1 _22553_ (.Y(_00760_),
    .A(_05007_),
    .B(_00759_));
 sg13g2_o21ai_1 _22554_ (.B1(_00760_),
    .Y(_00761_),
    .A1(_05024_),
    .A2(_00756_));
 sg13g2_nor3_1 _22555_ (.A(net266),
    .B(net357),
    .C(_00756_),
    .Y(_00762_));
 sg13g2_buf_2 _22556_ (.A(_00066_),
    .X(_00763_));
 sg13g2_inv_1 _22557_ (.Y(_00764_),
    .A(_00682_));
 sg13g2_xnor2_1 _22558_ (.Y(_00765_),
    .A(_09421_),
    .B(_00757_));
 sg13g2_xnor2_1 _22559_ (.Y(_00767_),
    .A(net691),
    .B(_00765_));
 sg13g2_nor4_1 _22560_ (.A(_09419_),
    .B(_00763_),
    .C(_00764_),
    .D(_00767_),
    .Y(_00768_));
 sg13g2_a221oi_1 _22561_ (.B2(net692),
    .C1(_00768_),
    .B1(_00762_),
    .A1(net266),
    .Y(_00769_),
    .A2(_00761_));
 sg13g2_a22oi_1 _22562_ (.Y(_00770_),
    .B1(_00756_),
    .B2(_05104_),
    .A2(_00757_),
    .A1(net1025));
 sg13g2_inv_2 _22563_ (.Y(_00771_),
    .A(net778));
 sg13g2_o21ai_1 _22564_ (.B1(net690),
    .Y(_00772_),
    .A1(_09411_),
    .A2(_04958_));
 sg13g2_nand3_1 _22565_ (.B(_00771_),
    .C(_00772_),
    .A(_00718_),
    .Y(_00773_));
 sg13g2_o21ai_1 _22566_ (.B1(_00773_),
    .Y(_00774_),
    .A1(_09408_),
    .A2(_00770_));
 sg13g2_nand2_1 _22567_ (.Y(_00775_),
    .A(_05007_),
    .B(_04945_));
 sg13g2_buf_1 _22568_ (.A(net778),
    .X(_00776_));
 sg13g2_buf_1 _22569_ (.A(_00776_),
    .X(_00778_));
 sg13g2_nor3_1 _22570_ (.A(net546),
    .B(net779),
    .C(net205),
    .Y(_00779_));
 sg13g2_a22oi_1 _22571_ (.Y(_00780_),
    .B1(_00775_),
    .B2(_00779_),
    .A2(_00774_),
    .A1(_05024_));
 sg13g2_nand2_1 _22572_ (.Y(_00781_),
    .A(_00763_),
    .B(_04721_));
 sg13g2_xnor2_1 _22573_ (.Y(_00782_),
    .A(net548),
    .B(_00767_));
 sg13g2_nand2b_1 _22574_ (.Y(_00783_),
    .B(_04884_),
    .A_N(_00763_));
 sg13g2_o21ai_1 _22575_ (.B1(_00783_),
    .Y(_00784_),
    .A1(_09419_),
    .A2(_00767_));
 sg13g2_a21oi_1 _22576_ (.A1(_00781_),
    .A2(_00782_),
    .Y(_00785_),
    .B1(_00784_));
 sg13g2_xnor2_1 _22577_ (.Y(_00786_),
    .A(_00780_),
    .B(_00785_));
 sg13g2_a21oi_1 _22578_ (.A1(_00769_),
    .A2(_00786_),
    .Y(_00787_),
    .B1(_11608_));
 sg13g2_xnor2_1 _22579_ (.Y(_00789_),
    .A(net438),
    .B(_00682_));
 sg13g2_xnor2_1 _22580_ (.Y(_00790_),
    .A(_00767_),
    .B(_00789_));
 sg13g2_a21oi_1 _22581_ (.A1(net66),
    .A2(_00790_),
    .Y(_00791_),
    .B1(net267));
 sg13g2_or3_1 _22582_ (.A(_00706_),
    .B(_00787_),
    .C(_00791_),
    .X(_00792_));
 sg13g2_o21ai_1 _22583_ (.B1(_00792_),
    .Y(_00458_),
    .A1(_06762_),
    .A2(_00662_));
 sg13g2_nand2_1 _22584_ (.Y(_00793_),
    .A(net31),
    .B(_00611_));
 sg13g2_nand2_1 _22585_ (.Y(_00794_),
    .A(_05006_),
    .B(net374));
 sg13g2_nand2_1 _22586_ (.Y(_00795_),
    .A(_00771_),
    .B(_13194_));
 sg13g2_xor2_1 _22587_ (.B(_09184_),
    .A(_05102_),
    .X(_00796_));
 sg13g2_nand2_1 _22588_ (.Y(_00797_),
    .A(net778),
    .B(_13193_));
 sg13g2_buf_2 _22589_ (.A(_00797_),
    .X(_00799_));
 sg13g2_and2_1 _22590_ (.A(net1177),
    .B(_00799_),
    .X(_00800_));
 sg13g2_nor2_2 _22591_ (.A(net1177),
    .B(_00799_),
    .Y(_00801_));
 sg13g2_a221oi_1 _22592_ (.B2(net273),
    .C1(_00801_),
    .B1(_00800_),
    .A1(_00795_),
    .Y(_00802_),
    .A2(_00796_));
 sg13g2_nor2_1 _22593_ (.A(net778),
    .B(net785),
    .Y(_00803_));
 sg13g2_nand2_1 _22594_ (.Y(_00804_),
    .A(_09180_),
    .B(_00803_));
 sg13g2_o21ai_1 _22595_ (.B1(_00804_),
    .Y(_00805_),
    .A1(_09222_),
    .A2(_00799_));
 sg13g2_a21oi_1 _22596_ (.A1(net778),
    .A2(net785),
    .Y(_00806_),
    .B1(net896));
 sg13g2_o21ai_1 _22597_ (.B1(net1177),
    .Y(_00807_),
    .A1(_00803_),
    .A2(_00806_));
 sg13g2_a21oi_1 _22598_ (.A1(_00804_),
    .A2(_00807_),
    .Y(_00808_),
    .B1(_02442_));
 sg13g2_a221oi_1 _22599_ (.B2(_05105_),
    .C1(_00808_),
    .B1(_00805_),
    .A1(net270),
    .Y(_00810_),
    .A2(_00801_));
 sg13g2_o21ai_1 _22600_ (.B1(_00810_),
    .Y(_00811_),
    .A1(_00794_),
    .A2(_00802_));
 sg13g2_nor2_1 _22601_ (.A(net205),
    .B(_13199_),
    .Y(_00812_));
 sg13g2_xnor2_1 _22602_ (.Y(_00813_),
    .A(_00752_),
    .B(_13192_));
 sg13g2_nor2_1 _22603_ (.A(_05104_),
    .B(_00813_),
    .Y(_00814_));
 sg13g2_a21oi_1 _22604_ (.A1(_02572_),
    .A2(_00799_),
    .Y(_00815_),
    .B1(_00814_));
 sg13g2_a21o_1 _22605_ (.A2(_09487_),
    .A1(_02432_),
    .B1(_00795_),
    .X(_00816_));
 sg13g2_o21ai_1 _22606_ (.B1(_00816_),
    .Y(_00817_),
    .A1(net273),
    .A2(_00815_));
 sg13g2_a22oi_1 _22607_ (.Y(_00818_),
    .B1(_00817_),
    .B2(net1177),
    .A2(_00794_),
    .A1(_00812_));
 sg13g2_xnor2_1 _22608_ (.Y(_00819_),
    .A(net1041),
    .B(_00813_));
 sg13g2_xnor2_1 _22609_ (.Y(_00821_),
    .A(net896),
    .B(_05005_));
 sg13g2_xnor2_1 _22610_ (.Y(_00822_),
    .A(_00819_),
    .B(_00821_));
 sg13g2_xnor2_1 _22611_ (.Y(_00823_),
    .A(net547),
    .B(_00822_));
 sg13g2_nand2_1 _22612_ (.Y(_00824_),
    .A(_09461_),
    .B(_00822_));
 sg13g2_o21ai_1 _22613_ (.B1(_00824_),
    .Y(_00825_),
    .A1(_04958_),
    .A2(_00823_));
 sg13g2_mux2_1 _22614_ (.A0(_00811_),
    .A1(_00818_),
    .S(_00825_),
    .X(_00826_));
 sg13g2_buf_1 _22615_ (.A(_00098_),
    .X(_00827_));
 sg13g2_xnor2_1 _22616_ (.Y(_00828_),
    .A(_00725_),
    .B(_00822_));
 sg13g2_nand2b_1 _22617_ (.Y(_00829_),
    .B(_00828_),
    .A_N(_00827_));
 sg13g2_nand2b_1 _22618_ (.Y(_00830_),
    .B(_00829_),
    .A_N(_00826_));
 sg13g2_nor3_1 _22619_ (.A(_00825_),
    .B(_00818_),
    .C(_00829_),
    .Y(_00831_));
 sg13g2_nor2_1 _22620_ (.A(net117),
    .B(_00831_),
    .Y(_00832_));
 sg13g2_xnor2_1 _22621_ (.Y(_00833_),
    .A(net437),
    .B(_00828_));
 sg13g2_o21ai_1 _22622_ (.B1(net545),
    .Y(_00834_),
    .A1(_04915_),
    .A2(_00833_));
 sg13g2_nand2_1 _22623_ (.Y(_00835_),
    .A(net53),
    .B(_00834_));
 sg13g2_a21o_1 _22624_ (.A2(_00832_),
    .A1(_00830_),
    .B1(_00835_),
    .X(_00836_));
 sg13g2_a21oi_1 _22625_ (.A1(_00793_),
    .A2(_00836_),
    .Y(_00459_),
    .B1(net440));
 sg13g2_nand3_1 _22626_ (.B(net120),
    .C(net53),
    .A(_09201_),
    .Y(_00837_));
 sg13g2_o21ai_1 _22627_ (.B1(_00837_),
    .Y(_00838_),
    .A1(net121),
    .A2(net53));
 sg13g2_nor2_1 _22628_ (.A(_11347_),
    .B(_13185_),
    .Y(_00839_));
 sg13g2_xnor2_1 _22629_ (.Y(_00841_),
    .A(_09421_),
    .B(_00819_));
 sg13g2_xor2_1 _22630_ (.B(_00841_),
    .A(_13309_),
    .X(_00842_));
 sg13g2_xor2_1 _22631_ (.B(net890),
    .A(_02475_),
    .X(_00843_));
 sg13g2_nor4_1 _22632_ (.A(_09206_),
    .B(net784),
    .C(_00841_),
    .D(_00843_),
    .Y(_00844_));
 sg13g2_xor2_1 _22633_ (.B(net436),
    .A(_05005_),
    .X(_00845_));
 sg13g2_nand2_1 _22634_ (.Y(_00846_),
    .A(net445),
    .B(_00845_));
 sg13g2_nand3_1 _22635_ (.B(net436),
    .C(_13194_),
    .A(_05006_),
    .Y(_00847_));
 sg13g2_a21oi_1 _22636_ (.A1(_00846_),
    .A2(_00847_),
    .Y(_00848_),
    .B1(_02572_));
 sg13g2_o21ai_1 _22637_ (.B1(net546),
    .Y(_00849_),
    .A1(_00801_),
    .A2(_00848_));
 sg13g2_nand4_1 _22638_ (.B(net205),
    .C(net207),
    .A(net174),
    .Y(_00850_),
    .D(_09436_));
 sg13g2_nand4_1 _22639_ (.B(net171),
    .C(_00849_),
    .A(net1197),
    .Y(_00852_),
    .D(_00850_));
 sg13g2_or2_1 _22640_ (.X(_00853_),
    .B(_00852_),
    .A(_00844_));
 sg13g2_a221oi_1 _22641_ (.B2(net272),
    .C1(_00853_),
    .B1(_00842_),
    .A1(_05183_),
    .Y(_00854_),
    .A2(_00839_));
 sg13g2_xor2_1 _22642_ (.B(net546),
    .A(net1177),
    .X(_00855_));
 sg13g2_a221oi_1 _22643_ (.B2(_00795_),
    .C1(_00801_),
    .B1(_00855_),
    .A1(net266),
    .Y(_00856_),
    .A2(_00800_));
 sg13g2_nand4_1 _22644_ (.B(_02442_),
    .C(net205),
    .A(net886),
    .Y(_00857_),
    .D(net207));
 sg13g2_o21ai_1 _22645_ (.B1(_00857_),
    .Y(_00858_),
    .A1(net546),
    .A2(_00795_));
 sg13g2_a21o_1 _22646_ (.A2(_00799_),
    .A1(net545),
    .B1(_00803_),
    .X(_00859_));
 sg13g2_a22oi_1 _22647_ (.Y(_00860_),
    .B1(_00859_),
    .B2(net1177),
    .A2(_00803_),
    .A1(net545));
 sg13g2_nor2_1 _22648_ (.A(net174),
    .B(_00860_),
    .Y(_00861_));
 sg13g2_a221oi_1 _22649_ (.B2(_05105_),
    .C1(_00861_),
    .B1(_00858_),
    .A1(net266),
    .Y(_00863_),
    .A2(_00801_));
 sg13g2_o21ai_1 _22650_ (.B1(_00863_),
    .Y(_00864_),
    .A1(_00794_),
    .A2(_00856_));
 sg13g2_xnor2_1 _22651_ (.Y(_00865_),
    .A(net890),
    .B(_00841_));
 sg13g2_o21ai_1 _22652_ (.B1(_13225_),
    .Y(_00866_),
    .A1(_09206_),
    .A2(_00841_));
 sg13g2_a21oi_1 _22653_ (.A1(_13218_),
    .A2(_00865_),
    .Y(_00867_),
    .B1(_00866_));
 sg13g2_xor2_1 _22654_ (.B(_00867_),
    .A(_00864_),
    .X(_00868_));
 sg13g2_a22oi_1 _22655_ (.Y(_00869_),
    .B1(_00854_),
    .B2(_00868_),
    .A2(_00838_),
    .A1(net356));
 sg13g2_inv_1 _22656_ (.Y(_00460_),
    .A(_00869_));
 sg13g2_nor2_1 _22657_ (.A(_08349_),
    .B(_12448_),
    .Y(_00870_));
 sg13g2_nand2_1 _22658_ (.Y(_00871_),
    .A(net327),
    .B(_00870_));
 sg13g2_buf_1 _22659_ (.A(_00871_),
    .X(_00873_));
 sg13g2_nor2_1 _22660_ (.A(net40),
    .B(_00873_),
    .Y(_00874_));
 sg13g2_buf_1 _22661_ (.A(net371),
    .X(_00875_));
 sg13g2_and2_1 _22662_ (.A(net1039),
    .B(_12832_),
    .X(_00876_));
 sg13g2_buf_1 _22663_ (.A(_00876_),
    .X(_00877_));
 sg13g2_xnor2_1 _22664_ (.Y(_00878_),
    .A(net372),
    .B(net209));
 sg13g2_o21ai_1 _22665_ (.B1(_12458_),
    .Y(_00879_),
    .A1(net804),
    .A2(_00877_));
 sg13g2_a21oi_1 _22666_ (.A1(net806),
    .A2(_00878_),
    .Y(_00880_),
    .B1(_00879_));
 sg13g2_a21oi_1 _22667_ (.A1(_12950_),
    .A2(_00877_),
    .Y(_00881_),
    .B1(_00880_));
 sg13g2_and3_1 _22668_ (.X(_00882_),
    .A(net1039),
    .B(_12455_),
    .C(_12832_));
 sg13g2_buf_1 _22669_ (.A(_00882_),
    .X(_00884_));
 sg13g2_a21oi_1 _22670_ (.A1(net461),
    .A2(_00884_),
    .Y(_00885_),
    .B1(net135));
 sg13g2_a21oi_1 _22671_ (.A1(net135),
    .A2(_00881_),
    .Y(_00886_),
    .B1(_00885_));
 sg13g2_xnor2_1 _22672_ (.Y(_00887_),
    .A(_12452_),
    .B(_12829_));
 sg13g2_xor2_1 _22673_ (.B(_12870_),
    .A(_02226_),
    .X(_00888_));
 sg13g2_xnor2_1 _22674_ (.Y(_00889_),
    .A(_00887_),
    .B(_00888_));
 sg13g2_buf_2 _22675_ (.A(_00889_),
    .X(_00890_));
 sg13g2_xor2_1 _22676_ (.B(net1184),
    .A(net802),
    .X(_00891_));
 sg13g2_xnor2_1 _22677_ (.Y(_00892_),
    .A(_00890_),
    .B(_00891_));
 sg13g2_nor2_1 _22678_ (.A(net792),
    .B(_00892_),
    .Y(_00893_));
 sg13g2_nor3_1 _22679_ (.A(net102),
    .B(_00886_),
    .C(_00893_),
    .Y(_00894_));
 sg13g2_nand2_1 _22680_ (.Y(_00895_),
    .A(net1043),
    .B(_00890_));
 sg13g2_o21ai_1 _22681_ (.B1(_12820_),
    .Y(_00896_),
    .A1(net1043),
    .A2(_00890_));
 sg13g2_xor2_1 _22682_ (.B(_00888_),
    .A(_12452_),
    .X(_00897_));
 sg13g2_nor2_1 _22683_ (.A(_12948_),
    .B(_00897_),
    .Y(_00898_));
 sg13g2_a21oi_1 _22684_ (.A1(_00895_),
    .A2(_00896_),
    .Y(_00899_),
    .B1(_00898_));
 sg13g2_o21ai_1 _22685_ (.B1(_00890_),
    .Y(_00900_),
    .A1(net1043),
    .A2(_00898_));
 sg13g2_nor2_1 _22686_ (.A(net1043),
    .B(_00890_),
    .Y(_00901_));
 sg13g2_a21o_1 _22687_ (.A2(_00890_),
    .A1(_12820_),
    .B1(net1043),
    .X(_00902_));
 sg13g2_mux2_1 _22688_ (.A0(_00901_),
    .A1(_00902_),
    .S(_00898_),
    .X(_00903_));
 sg13g2_a21o_1 _22689_ (.A2(_00900_),
    .A1(net802),
    .B1(_00903_),
    .X(_00905_));
 sg13g2_nor2b_1 _22690_ (.A(_12593_),
    .B_N(net453),
    .Y(_00906_));
 sg13g2_nor2_1 _22691_ (.A(net175),
    .B(_00906_),
    .Y(_00907_));
 sg13g2_a21oi_1 _22692_ (.A1(net175),
    .A2(net209),
    .Y(_00908_),
    .B1(_00907_));
 sg13g2_nor2b_1 _22693_ (.A(net453),
    .B_N(net707),
    .Y(_00909_));
 sg13g2_a21oi_1 _22694_ (.A1(_02604_),
    .A2(_12457_),
    .Y(_00910_),
    .B1(_00909_));
 sg13g2_nor2_1 _22695_ (.A(_12473_),
    .B(_00910_),
    .Y(_00911_));
 sg13g2_nor3_1 _22696_ (.A(net372),
    .B(net452),
    .C(_12593_),
    .Y(_00912_));
 sg13g2_nor2_1 _22697_ (.A(_00911_),
    .B(_00912_),
    .Y(_00913_));
 sg13g2_o21ai_1 _22698_ (.B1(_00913_),
    .Y(_00914_),
    .A1(net137),
    .A2(_00908_));
 sg13g2_nor2_1 _22699_ (.A(net1038),
    .B(_02583_),
    .Y(_00916_));
 sg13g2_buf_2 _22700_ (.A(_00916_),
    .X(_00917_));
 sg13g2_nand2_1 _22701_ (.Y(_00918_),
    .A(_12458_),
    .B(_00917_));
 sg13g2_nand4_1 _22702_ (.B(net173),
    .C(net209),
    .A(net706),
    .Y(_00919_),
    .D(net799));
 sg13g2_o21ai_1 _22703_ (.B1(_00919_),
    .Y(_00920_),
    .A1(net209),
    .A2(_00918_));
 sg13g2_mux2_1 _22704_ (.A0(_12593_),
    .A1(_12457_),
    .S(net452),
    .X(_00921_));
 sg13g2_nand2_1 _22705_ (.Y(_00922_),
    .A(net372),
    .B(_00921_));
 sg13g2_o21ai_1 _22706_ (.B1(_00922_),
    .Y(_00923_),
    .A1(net173),
    .A2(_00906_));
 sg13g2_nor2_1 _22707_ (.A(net1039),
    .B(_12833_),
    .Y(_00924_));
 sg13g2_nand2b_1 _22708_ (.Y(_00925_),
    .B(_12507_),
    .A_N(_00924_));
 sg13g2_a21oi_1 _22709_ (.A1(_00923_),
    .A2(_00925_),
    .Y(_00927_),
    .B1(net371));
 sg13g2_a221oi_1 _22710_ (.B2(net461),
    .C1(_00927_),
    .B1(_00920_),
    .A1(net135),
    .Y(_00928_),
    .A2(_00914_));
 sg13g2_mux2_1 _22711_ (.A0(_00899_),
    .A1(_00905_),
    .S(_00928_),
    .X(_00929_));
 sg13g2_nor3_1 _22712_ (.A(net176),
    .B(_08349_),
    .C(_12448_),
    .Y(_00930_));
 sg13g2_a221oi_1 _22713_ (.B2(_00929_),
    .C1(_00930_),
    .B1(_00894_),
    .A1(net792),
    .Y(_00931_),
    .A2(net71));
 sg13g2_nor3_1 _22714_ (.A(net557),
    .B(_00874_),
    .C(_00931_),
    .Y(_00461_));
 sg13g2_or3_1 _22715_ (.A(net706),
    .B(net450),
    .C(net367),
    .X(_00932_));
 sg13g2_nand4_1 _22716_ (.B(net215),
    .C(net450),
    .A(net371),
    .Y(_00933_),
    .D(net367));
 sg13g2_a21oi_1 _22717_ (.A1(_00932_),
    .A2(_00933_),
    .Y(_00934_),
    .B1(net461));
 sg13g2_nand2b_1 _22718_ (.Y(_00935_),
    .B(_12593_),
    .A_N(net702));
 sg13g2_nor3_1 _22719_ (.A(_12567_),
    .B(net210),
    .C(_00935_),
    .Y(_00937_));
 sg13g2_nor2b_1 _22720_ (.A(_12593_),
    .B_N(net702),
    .Y(_00938_));
 sg13g2_nor2_1 _22721_ (.A(net702),
    .B(_12540_),
    .Y(_00939_));
 sg13g2_or2_1 _22722_ (.X(_00940_),
    .B(_00939_),
    .A(_00938_));
 sg13g2_nor2_1 _22723_ (.A(net703),
    .B(_12594_),
    .Y(_00941_));
 sg13g2_nor3_1 _22724_ (.A(net450),
    .B(_12540_),
    .C(_00941_),
    .Y(_00942_));
 sg13g2_a21oi_1 _22725_ (.A1(net210),
    .A2(_00940_),
    .Y(_00943_),
    .B1(_00942_));
 sg13g2_nor2b_1 _22726_ (.A(_00943_),
    .B_N(net371),
    .Y(_00944_));
 sg13g2_o21ai_1 _22727_ (.B1(_00935_),
    .Y(_00945_),
    .A1(net450),
    .A2(_00938_));
 sg13g2_nand2_1 _22728_ (.Y(_00946_),
    .A(net703),
    .B(_12594_));
 sg13g2_o21ai_1 _22729_ (.B1(net450),
    .Y(_00948_),
    .A1(net702),
    .A2(_12593_));
 sg13g2_a21oi_1 _22730_ (.A1(_00946_),
    .A2(_00948_),
    .Y(_00949_),
    .B1(_12540_));
 sg13g2_a21oi_1 _22731_ (.A1(_12533_),
    .A2(_00945_),
    .Y(_00950_),
    .B1(_00949_));
 sg13g2_nor2_1 _22732_ (.A(net135),
    .B(_00950_),
    .Y(_00951_));
 sg13g2_nor4_1 _22733_ (.A(_00934_),
    .B(_00937_),
    .C(_00944_),
    .D(_00951_),
    .Y(_00952_));
 sg13g2_nand2_1 _22734_ (.Y(_00953_),
    .A(_12820_),
    .B(net1043));
 sg13g2_xor2_1 _22735_ (.B(_12895_),
    .A(_03240_),
    .X(_00954_));
 sg13g2_xnor2_1 _22736_ (.Y(_00955_),
    .A(net804),
    .B(_00954_));
 sg13g2_xnor2_1 _22737_ (.Y(_00956_),
    .A(net792),
    .B(_00955_));
 sg13g2_nand2_1 _22738_ (.Y(_00957_),
    .A(_12492_),
    .B(_02518_));
 sg13g2_o21ai_1 _22739_ (.B1(_00957_),
    .Y(_00959_),
    .A1(_12864_),
    .A2(_00955_));
 sg13g2_a21oi_1 _22740_ (.A1(_00953_),
    .A2(_00956_),
    .Y(_00960_),
    .B1(_00959_));
 sg13g2_xnor2_1 _22741_ (.Y(_00961_),
    .A(_00952_),
    .B(_00960_));
 sg13g2_xnor2_1 _22742_ (.Y(_00962_),
    .A(net450),
    .B(net367));
 sg13g2_a21oi_1 _22743_ (.A1(_12936_),
    .A2(net367),
    .Y(_00963_),
    .B1(_12453_));
 sg13g2_a21oi_1 _22744_ (.A1(_12453_),
    .A2(_00962_),
    .Y(_00964_),
    .B1(_00963_));
 sg13g2_a22oi_1 _22745_ (.Y(_00965_),
    .B1(_00964_),
    .B2(_12567_),
    .A2(_00938_),
    .A1(net210));
 sg13g2_nor2b_1 _22746_ (.A(_00965_),
    .B_N(net135),
    .Y(_00966_));
 sg13g2_and3_1 _22747_ (.X(_00967_),
    .A(_02518_),
    .B(_12866_),
    .C(_12930_));
 sg13g2_nor2b_1 _22748_ (.A(_00955_),
    .B_N(_00967_),
    .Y(_00968_));
 sg13g2_nand3_1 _22749_ (.B(net169),
    .C(_12894_),
    .A(_12454_),
    .Y(_00970_));
 sg13g2_o21ai_1 _22750_ (.B1(net118),
    .Y(_00971_),
    .A1(net135),
    .A2(_00970_));
 sg13g2_xnor2_1 _22751_ (.Y(_00972_),
    .A(net1184),
    .B(_12930_));
 sg13g2_xnor2_1 _22752_ (.Y(_00973_),
    .A(_00955_),
    .B(_00972_));
 sg13g2_nor2_1 _22753_ (.A(net211),
    .B(_00973_),
    .Y(_00974_));
 sg13g2_nor4_1 _22754_ (.A(_00966_),
    .B(_00968_),
    .C(_00971_),
    .D(_00974_),
    .Y(_00975_));
 sg13g2_a22oi_1 _22755_ (.Y(_00976_),
    .B1(_00961_),
    .B2(_00975_),
    .A2(net67),
    .A1(net211));
 sg13g2_buf_1 _22756_ (.A(_00788_),
    .X(_00977_));
 sg13g2_o21ai_1 _22757_ (.B1(net435),
    .Y(_00978_),
    .A1(net38),
    .A2(_00873_));
 sg13g2_a21oi_1 _22758_ (.A1(_00873_),
    .A2(_00976_),
    .Y(_00462_),
    .B1(_00978_));
 sg13g2_nand2_2 _22759_ (.Y(_00980_),
    .A(net714),
    .B(_00930_));
 sg13g2_and2_1 _22760_ (.A(net1030),
    .B(net790),
    .X(_00981_));
 sg13g2_xor2_1 _22761_ (.B(_12937_),
    .A(net1030),
    .X(_00982_));
 sg13g2_nand2_1 _22762_ (.Y(_00983_),
    .A(_12517_),
    .B(_00982_));
 sg13g2_o21ai_1 _22763_ (.B1(_00983_),
    .Y(_00984_),
    .A1(_12570_),
    .A2(_00981_));
 sg13g2_nand2_1 _22764_ (.Y(_00985_),
    .A(_12518_),
    .B(_12570_));
 sg13g2_nor2_1 _22765_ (.A(net698),
    .B(net449),
    .Y(_00986_));
 sg13g2_a22oi_1 _22766_ (.Y(_00987_),
    .B1(_00985_),
    .B2(_00986_),
    .A2(_00984_),
    .A1(_12630_));
 sg13g2_inv_2 _22767_ (.Y(_00988_),
    .A(net1089));
 sg13g2_a21oi_1 _22768_ (.A1(_12518_),
    .A2(net703),
    .Y(_00989_),
    .B1(_00988_));
 sg13g2_nand3b_1 _22769_ (.B(_00986_),
    .C(_12630_),
    .Y(_00991_),
    .A_N(_00989_));
 sg13g2_o21ai_1 _22770_ (.B1(_00991_),
    .Y(_00992_),
    .A1(net367),
    .A2(_00987_));
 sg13g2_nand2b_1 _22771_ (.Y(_00993_),
    .B(_04363_),
    .A_N(net806));
 sg13g2_xor2_1 _22772_ (.B(net1089),
    .A(_04163_),
    .X(_00994_));
 sg13g2_xnor2_1 _22773_ (.Y(_00995_),
    .A(_03218_),
    .B(_12937_));
 sg13g2_xnor2_1 _22774_ (.Y(_00996_),
    .A(_00994_),
    .B(_00995_));
 sg13g2_xnor2_1 _22775_ (.Y(_00997_),
    .A(_12517_),
    .B(_00996_));
 sg13g2_xnor2_1 _22776_ (.Y(_00998_),
    .A(net451),
    .B(_00997_));
 sg13g2_nand2b_1 _22777_ (.Y(_00999_),
    .B(_12473_),
    .A_N(_04363_));
 sg13g2_o21ai_1 _22778_ (.B1(_00999_),
    .Y(_01000_),
    .A1(_12948_),
    .A2(_00997_));
 sg13g2_a21oi_1 _22779_ (.A1(_00993_),
    .A2(_00998_),
    .Y(_01002_),
    .B1(_01000_));
 sg13g2_xor2_1 _22780_ (.B(_01002_),
    .A(_00992_),
    .X(_01003_));
 sg13g2_nand2_1 _22781_ (.Y(_01004_),
    .A(net1030),
    .B(net790));
 sg13g2_o21ai_1 _22782_ (.B1(_00983_),
    .Y(_01005_),
    .A1(net458),
    .A2(_01004_));
 sg13g2_nand2_1 _22783_ (.Y(_01006_),
    .A(net457),
    .B(_01005_));
 sg13g2_o21ai_1 _22784_ (.B1(_01006_),
    .Y(_01007_),
    .A1(_12630_),
    .A2(_01004_));
 sg13g2_nor3_1 _22785_ (.A(_12533_),
    .B(net169),
    .C(_12939_),
    .Y(_01008_));
 sg13g2_nand2b_1 _22786_ (.Y(_01009_),
    .B(_00887_),
    .A_N(_04363_));
 sg13g2_nor3_1 _22787_ (.A(_12948_),
    .B(_00997_),
    .C(_01009_),
    .Y(_01010_));
 sg13g2_a221oi_1 _22788_ (.B2(net365),
    .C1(_01010_),
    .B1(_01008_),
    .A1(net169),
    .Y(_01011_),
    .A2(_01007_));
 sg13g2_a21oi_1 _22789_ (.A1(_01003_),
    .A2(_01011_),
    .Y(_01013_),
    .B1(net117));
 sg13g2_xnor2_1 _22790_ (.Y(_01014_),
    .A(net371),
    .B(_00887_));
 sg13g2_xnor2_1 _22791_ (.Y(_01015_),
    .A(_00997_),
    .B(_01014_));
 sg13g2_a21oi_1 _22792_ (.A1(net122),
    .A2(_01015_),
    .Y(_01016_),
    .B1(net210));
 sg13g2_nand2_1 _22793_ (.Y(_01017_),
    .A(net1059),
    .B(_00873_));
 sg13g2_or3_1 _22794_ (.A(_01013_),
    .B(_01016_),
    .C(_01017_),
    .X(_01018_));
 sg13g2_o21ai_1 _22795_ (.B1(_01018_),
    .Y(_00463_),
    .A1(net35),
    .A2(_00980_));
 sg13g2_or2_1 _22796_ (.X(_01019_),
    .B(net1084),
    .A(_04163_));
 sg13g2_buf_1 _22797_ (.A(_01019_),
    .X(_01020_));
 sg13g2_nand2_1 _22798_ (.Y(_01021_),
    .A(_04841_),
    .B(net798));
 sg13g2_o21ai_1 _22799_ (.B1(net789),
    .Y(_01023_),
    .A1(net694),
    .A2(net698));
 sg13g2_o21ai_1 _22800_ (.B1(_01023_),
    .Y(_01024_),
    .A1(_01020_),
    .A2(_01021_));
 sg13g2_a221oi_1 _22801_ (.B2(net798),
    .C1(_01024_),
    .B1(_00988_),
    .A1(net694),
    .Y(_01025_),
    .A2(_04264_));
 sg13g2_a21oi_1 _22802_ (.A1(_12616_),
    .A2(_12646_),
    .Y(_01026_),
    .B1(_01020_));
 sg13g2_a22oi_1 _22803_ (.Y(_01027_),
    .B1(_01026_),
    .B2(_04841_),
    .A2(_01025_),
    .A1(_12658_));
 sg13g2_nand2_1 _22804_ (.Y(_01028_),
    .A(_12533_),
    .B(_00251_));
 sg13g2_xor2_1 _22805_ (.B(_12983_),
    .A(_04861_),
    .X(_01029_));
 sg13g2_xnor2_1 _22806_ (.Y(_01030_),
    .A(_00988_),
    .B(_01029_));
 sg13g2_xnor2_1 _22807_ (.Y(_01031_),
    .A(net210),
    .B(_01030_));
 sg13g2_nand2_1 _22808_ (.Y(_01032_),
    .A(net215),
    .B(_04875_));
 sg13g2_o21ai_1 _22809_ (.B1(_01032_),
    .Y(_01033_),
    .A1(_12978_),
    .A2(_01030_));
 sg13g2_a21oi_1 _22810_ (.A1(_01028_),
    .A2(_01031_),
    .Y(_01034_),
    .B1(_01033_));
 sg13g2_xnor2_1 _22811_ (.Y(_01035_),
    .A(_01027_),
    .B(_01034_));
 sg13g2_nor2_1 _22812_ (.A(_12978_),
    .B(_01030_),
    .Y(_01036_));
 sg13g2_and2_1 _22813_ (.A(_04875_),
    .B(_12895_),
    .X(_01037_));
 sg13g2_nand2_1 _22814_ (.Y(_01038_),
    .A(_04174_),
    .B(net1084));
 sg13g2_xor2_1 _22815_ (.B(net789),
    .A(_12569_),
    .X(_01039_));
 sg13g2_and2_1 _22816_ (.A(net698),
    .B(_01039_),
    .X(_01040_));
 sg13g2_nor3_1 _22817_ (.A(_04264_),
    .B(_00988_),
    .C(_13021_),
    .Y(_01041_));
 sg13g2_o21ai_1 _22818_ (.B1(_12646_),
    .Y(_01042_),
    .A1(_01040_),
    .A2(_01041_));
 sg13g2_o21ai_1 _22819_ (.B1(_01042_),
    .Y(_01044_),
    .A1(_12658_),
    .A2(_01038_));
 sg13g2_nand2_1 _22820_ (.Y(_01045_),
    .A(net365),
    .B(net457));
 sg13g2_nor3_1 _22821_ (.A(net363),
    .B(_12990_),
    .C(_01045_),
    .Y(_01046_));
 sg13g2_a221oi_1 _22822_ (.B2(net363),
    .C1(_01046_),
    .B1(_01044_),
    .A1(_01036_),
    .Y(_01047_),
    .A2(_01037_));
 sg13g2_a21oi_1 _22823_ (.A1(_01035_),
    .A2(_01047_),
    .Y(_01048_),
    .B1(net96));
 sg13g2_xnor2_1 _22824_ (.Y(_01049_),
    .A(_04109_),
    .B(_12895_));
 sg13g2_xnor2_1 _22825_ (.Y(_01050_),
    .A(_01030_),
    .B(_01049_));
 sg13g2_a21oi_1 _22826_ (.A1(net66),
    .A2(_01050_),
    .Y(_01051_),
    .B1(net449));
 sg13g2_or3_1 _22827_ (.A(_01017_),
    .B(_01048_),
    .C(_01051_),
    .X(_01052_));
 sg13g2_o21ai_1 _22828_ (.B1(_01052_),
    .Y(_00464_),
    .A1(net32),
    .A2(_00980_));
 sg13g2_nand2_1 _22829_ (.Y(_01054_),
    .A(net363),
    .B(_13076_));
 sg13g2_o21ai_1 _22830_ (.B1(_01054_),
    .Y(_01055_),
    .A1(_13019_),
    .A2(_01021_));
 sg13g2_nand2_1 _22831_ (.Y(_01056_),
    .A(_04789_),
    .B(net788));
 sg13g2_nor2_1 _22832_ (.A(_12697_),
    .B(_01056_),
    .Y(_01057_));
 sg13g2_a21o_1 _22833_ (.A2(_01055_),
    .A1(net213),
    .B1(_01057_),
    .X(_01058_));
 sg13g2_nand2_1 _22834_ (.Y(_01059_),
    .A(net363),
    .B(net456));
 sg13g2_nor2_1 _22835_ (.A(net361),
    .B(_01059_),
    .Y(_01060_));
 sg13g2_nand2b_1 _22836_ (.Y(_01061_),
    .B(_12653_),
    .A_N(net788));
 sg13g2_o21ai_1 _22837_ (.B1(net788),
    .Y(_01062_),
    .A1(net1024),
    .A2(net1027));
 sg13g2_o21ai_1 _22838_ (.B1(_01062_),
    .Y(_01063_),
    .A1(_04977_),
    .A2(_01061_));
 sg13g2_nand2b_1 _22839_ (.Y(_01065_),
    .B(_12653_),
    .A_N(net1088));
 sg13g2_nand3_1 _22840_ (.B(_04949_),
    .C(_01065_),
    .A(net1087),
    .Y(_01066_));
 sg13g2_nand2_1 _22841_ (.Y(_01067_),
    .A(net798),
    .B(net455));
 sg13g2_nor3_1 _22842_ (.A(net687),
    .B(net694),
    .C(_13016_),
    .Y(_01068_));
 sg13g2_nand2_1 _22843_ (.Y(_01069_),
    .A(_01067_),
    .B(_01068_));
 sg13g2_o21ai_1 _22844_ (.B1(_01069_),
    .Y(_01070_),
    .A1(_01063_),
    .A2(_01066_));
 sg13g2_xnor2_1 _22845_ (.Y(_01071_),
    .A(_04947_),
    .B(_12652_));
 sg13g2_xor2_1 _22846_ (.B(_01071_),
    .A(_13076_),
    .X(_01072_));
 sg13g2_xnor2_1 _22847_ (.Y(_01073_),
    .A(net694),
    .B(_01072_));
 sg13g2_nand2_1 _22848_ (.Y(_01074_),
    .A(_13052_),
    .B(_01073_));
 sg13g2_xnor2_1 _22849_ (.Y(_01076_),
    .A(_12937_),
    .B(net1088));
 sg13g2_xnor2_1 _22850_ (.Y(_01077_),
    .A(_13015_),
    .B(_01076_));
 sg13g2_xnor2_1 _22851_ (.Y(_01078_),
    .A(_04952_),
    .B(_01077_));
 sg13g2_buf_1 _22852_ (.A(_01078_),
    .X(_01079_));
 sg13g2_a21oi_1 _22853_ (.A1(_00988_),
    .A2(_01079_),
    .Y(_01080_),
    .B1(_04962_));
 sg13g2_nand2b_1 _22854_ (.Y(_01081_),
    .B(_12616_),
    .A_N(_01079_));
 sg13g2_o21ai_1 _22855_ (.B1(_01081_),
    .Y(_01082_),
    .A1(_01074_),
    .A2(_01080_));
 sg13g2_a21o_1 _22856_ (.A2(_01079_),
    .A1(_00988_),
    .B1(_04962_),
    .X(_01083_));
 sg13g2_o21ai_1 _22857_ (.B1(_04962_),
    .Y(_01084_),
    .A1(_00988_),
    .A2(_01079_));
 sg13g2_a21oi_1 _22858_ (.A1(_00988_),
    .A2(_01079_),
    .Y(_01085_),
    .B1(_01070_));
 sg13g2_a22oi_1 _22859_ (.Y(_01087_),
    .B1(_01084_),
    .B2(_01085_),
    .A2(_01083_),
    .A1(_01070_));
 sg13g2_a22oi_1 _22860_ (.Y(_01088_),
    .B1(_01087_),
    .B2(_01074_),
    .A2(_01082_),
    .A1(_01070_));
 sg13g2_a221oi_1 _22861_ (.B2(_13045_),
    .C1(_01088_),
    .B1(_01060_),
    .A1(net361),
    .Y(_01089_),
    .A2(_01058_));
 sg13g2_xnor2_1 _22862_ (.Y(_01090_),
    .A(_00994_),
    .B(_01079_));
 sg13g2_a21oi_1 _22863_ (.A1(net114),
    .A2(_01090_),
    .Y(_01091_),
    .B1(net789));
 sg13g2_nor2_1 _22864_ (.A(_01017_),
    .B(_01091_),
    .Y(_01092_));
 sg13g2_o21ai_1 _22865_ (.B1(_01092_),
    .Y(_01093_),
    .A1(net81),
    .A2(_01089_));
 sg13g2_o21ai_1 _22866_ (.B1(_01093_),
    .Y(_00465_),
    .A1(net29),
    .A2(_00980_));
 sg13g2_nand2_1 _22867_ (.Y(_01094_),
    .A(net1024),
    .B(net797));
 sg13g2_a21oi_1 _22868_ (.A1(net454),
    .A2(_01094_),
    .Y(_01095_),
    .B1(_13112_));
 sg13g2_nand2_1 _22869_ (.Y(_01097_),
    .A(net797),
    .B(net787));
 sg13g2_a21oi_1 _22870_ (.A1(net454),
    .A2(_01097_),
    .Y(_01098_),
    .B1(net687));
 sg13g2_nor2_1 _22871_ (.A(_01095_),
    .B(_01098_),
    .Y(_01099_));
 sg13g2_nand2_1 _22872_ (.Y(_01100_),
    .A(net688),
    .B(net455));
 sg13g2_or2_1 _22873_ (.X(_01101_),
    .B(net787),
    .A(net1024));
 sg13g2_buf_1 _22874_ (.A(_01101_),
    .X(_01102_));
 sg13g2_a21o_1 _22875_ (.A2(_01100_),
    .A1(_12721_),
    .B1(_01102_),
    .X(_01103_));
 sg13g2_o21ai_1 _22876_ (.B1(_01103_),
    .Y(_01104_),
    .A1(net358),
    .A2(_01099_));
 sg13g2_a21oi_1 _22877_ (.A1(net213),
    .A2(net136),
    .Y(_01105_),
    .B1(_05043_));
 sg13g2_a22oi_1 _22878_ (.Y(_01106_),
    .B1(_01105_),
    .B2(_13109_),
    .A2(_01104_),
    .A1(_12756_));
 sg13g2_nand2b_1 _22879_ (.Y(_01108_),
    .B(_05030_),
    .A_N(_12618_));
 sg13g2_xnor2_1 _22880_ (.Y(_01109_),
    .A(_13061_),
    .B(_01071_));
 sg13g2_xnor2_1 _22881_ (.Y(_01110_),
    .A(net688),
    .B(_01109_));
 sg13g2_xnor2_1 _22882_ (.Y(_01111_),
    .A(net789),
    .B(_01110_));
 sg13g2_nand2b_1 _22883_ (.Y(_01112_),
    .B(_12618_),
    .A_N(_05030_));
 sg13g2_o21ai_1 _22884_ (.B1(_01112_),
    .Y(_01113_),
    .A1(_13087_),
    .A2(_01110_));
 sg13g2_a21oi_1 _22885_ (.A1(_01108_),
    .A2(_01111_),
    .Y(_01114_),
    .B1(_01113_));
 sg13g2_xnor2_1 _22886_ (.Y(_01115_),
    .A(_01106_),
    .B(_01114_));
 sg13g2_and2_1 _22887_ (.A(net361),
    .B(net213),
    .X(_01116_));
 sg13g2_nor2_1 _22888_ (.A(net164),
    .B(_13065_),
    .Y(_01117_));
 sg13g2_nand2_1 _22889_ (.Y(_01119_),
    .A(net687),
    .B(_13108_));
 sg13g2_xor2_1 _22890_ (.B(net447),
    .A(net797),
    .X(_01120_));
 sg13g2_nand2_1 _22891_ (.Y(_01121_),
    .A(net687),
    .B(_01120_));
 sg13g2_o21ai_1 _22892_ (.B1(_01121_),
    .Y(_01122_),
    .A1(net361),
    .A2(_01097_));
 sg13g2_nand2_1 _22893_ (.Y(_01123_),
    .A(net136),
    .B(_01122_));
 sg13g2_o21ai_1 _22894_ (.B1(_01123_),
    .Y(_01124_),
    .A1(_12756_),
    .A2(_01119_));
 sg13g2_nand2b_1 _22895_ (.Y(_01125_),
    .B(_12983_),
    .A_N(_05030_));
 sg13g2_nor3_1 _22896_ (.A(_13087_),
    .B(_01110_),
    .C(_01125_),
    .Y(_01126_));
 sg13g2_a221oi_1 _22897_ (.B2(net164),
    .C1(_01126_),
    .B1(_01124_),
    .A1(_01116_),
    .Y(_01127_),
    .A2(_01117_));
 sg13g2_a21oi_1 _22898_ (.A1(_01115_),
    .A2(_01127_),
    .Y(_01128_),
    .B1(net96));
 sg13g2_xnor2_1 _22899_ (.Y(_01130_),
    .A(net363),
    .B(_12983_));
 sg13g2_xnor2_1 _22900_ (.Y(_01131_),
    .A(_01110_),
    .B(_01130_));
 sg13g2_a21oi_1 _22901_ (.A1(net66),
    .A2(_01131_),
    .Y(_01132_),
    .B1(net448));
 sg13g2_or3_1 _22902_ (.A(_01017_),
    .B(_01128_),
    .C(_01132_),
    .X(_01133_));
 sg13g2_o21ai_1 _22903_ (.B1(_01133_),
    .Y(_00466_),
    .A1(net43),
    .A2(_00980_));
 sg13g2_xnor2_1 _22904_ (.Y(_01134_),
    .A(_12716_),
    .B(net452));
 sg13g2_nand3_1 _22905_ (.B(_12716_),
    .C(_12837_),
    .A(_02604_),
    .Y(_01135_));
 sg13g2_o21ai_1 _22906_ (.B1(_01135_),
    .Y(_01136_),
    .A1(net175),
    .A2(_01134_));
 sg13g2_buf_2 _22907_ (.A(_00156_),
    .X(_01137_));
 sg13g2_inv_1 _22908_ (.Y(_01138_),
    .A(_01137_));
 sg13g2_and2_1 _22909_ (.A(_01138_),
    .B(_00877_),
    .X(_01140_));
 sg13g2_a21oi_1 _22910_ (.A1(net137),
    .A2(_01136_),
    .Y(_01141_),
    .B1(_01140_));
 sg13g2_a21oi_1 _22911_ (.A1(net136),
    .A2(_00884_),
    .Y(_01142_),
    .B1(net164));
 sg13g2_a21o_1 _22912_ (.A2(_01141_),
    .A1(net164),
    .B1(_01142_),
    .X(_01143_));
 sg13g2_xnor2_1 _22913_ (.Y(_01144_),
    .A(_05065_),
    .B(_12751_));
 sg13g2_xnor2_1 _22914_ (.Y(_01145_),
    .A(_12837_),
    .B(_01144_));
 sg13g2_nor2_1 _22915_ (.A(_05096_),
    .B(_13015_),
    .Y(_01146_));
 sg13g2_nand3_1 _22916_ (.B(_01145_),
    .C(_01146_),
    .A(_13130_),
    .Y(_01147_));
 sg13g2_xnor2_1 _22917_ (.Y(_01148_),
    .A(_13014_),
    .B(_12700_));
 sg13g2_xnor2_1 _22918_ (.Y(_01149_),
    .A(_12870_),
    .B(_01148_));
 sg13g2_xnor2_1 _22919_ (.Y(_01151_),
    .A(_05058_),
    .B(_01149_));
 sg13g2_nand2b_1 _22920_ (.Y(_01152_),
    .B(_05096_),
    .A_N(net455));
 sg13g2_nor2b_1 _22921_ (.A(_05096_),
    .B_N(_12661_),
    .Y(_01153_));
 sg13g2_a221oi_1 _22922_ (.B2(_01152_),
    .C1(_01153_),
    .B1(_01151_),
    .A1(_13130_),
    .Y(_01154_),
    .A2(_01145_));
 sg13g2_nand2b_1 _22923_ (.Y(_01155_),
    .B(_00924_),
    .A_N(net688));
 sg13g2_a21oi_1 _22924_ (.A1(net707),
    .A2(net794),
    .Y(_01156_),
    .B1(net1020));
 sg13g2_o21ai_1 _22925_ (.B1(_01137_),
    .Y(_01157_),
    .A1(_00924_),
    .A2(_01156_));
 sg13g2_a21o_1 _22926_ (.A2(_01157_),
    .A1(_01155_),
    .B1(_12469_),
    .X(_01158_));
 sg13g2_nor3_1 _22927_ (.A(_01137_),
    .B(net707),
    .C(_12834_),
    .Y(_01159_));
 sg13g2_nor3_1 _22928_ (.A(_12791_),
    .B(_00877_),
    .C(_01159_),
    .Y(_01160_));
 sg13g2_o21ai_1 _22929_ (.B1(net358),
    .Y(_01162_),
    .A1(_01140_),
    .A2(_01160_));
 sg13g2_nor2b_1 _22930_ (.A(net1020),
    .B_N(_01137_),
    .Y(_01163_));
 sg13g2_mux2_1 _22931_ (.A0(_12833_),
    .A1(_12455_),
    .S(net1039),
    .X(_01164_));
 sg13g2_a22oi_1 _22932_ (.Y(_01165_),
    .B1(_01163_),
    .B2(_01164_),
    .A2(_00884_),
    .A1(_01138_));
 sg13g2_nand2b_1 _22933_ (.Y(_01166_),
    .B(net212),
    .A_N(_01165_));
 sg13g2_nand3_1 _22934_ (.B(_12834_),
    .C(net165),
    .A(_12456_),
    .Y(_01167_));
 sg13g2_a21o_1 _22935_ (.A2(_01167_),
    .A1(_01155_),
    .B1(_12721_),
    .X(_01168_));
 sg13g2_nand4_1 _22936_ (.B(_01162_),
    .C(_01166_),
    .A(_01158_),
    .Y(_01169_),
    .D(_01168_));
 sg13g2_xor2_1 _22937_ (.B(_01169_),
    .A(_01154_),
    .X(_01170_));
 sg13g2_nand4_1 _22938_ (.B(_01143_),
    .C(_01147_),
    .A(net167),
    .Y(_01171_),
    .D(_01170_));
 sg13g2_xor2_1 _22939_ (.B(_01151_),
    .A(_01071_),
    .X(_01173_));
 sg13g2_nor2_1 _22940_ (.A(_01171_),
    .B(_01173_),
    .Y(_01174_));
 sg13g2_nand2_1 _22941_ (.Y(_01175_),
    .A(net85),
    .B(_01171_));
 sg13g2_o21ai_1 _22942_ (.B1(_01175_),
    .Y(_01176_),
    .A1(net208),
    .A2(_01174_));
 sg13g2_o21ai_1 _22943_ (.B1(net435),
    .Y(_01177_),
    .A1(net45),
    .A2(_00873_));
 sg13g2_a21oi_1 _22944_ (.A1(_00873_),
    .A2(_01176_),
    .Y(_00467_),
    .B1(_01177_));
 sg13g2_nor2_1 _22945_ (.A(net707),
    .B(net787),
    .Y(_01178_));
 sg13g2_nand2b_1 _22946_ (.Y(_01179_),
    .B(_01178_),
    .A_N(net688));
 sg13g2_and2_1 _22947_ (.A(_02583_),
    .B(_13062_),
    .X(_01180_));
 sg13g2_buf_1 _22948_ (.A(_01180_),
    .X(_01181_));
 sg13g2_nor2_1 _22949_ (.A(net688),
    .B(_01181_),
    .Y(_01183_));
 sg13g2_o21ai_1 _22950_ (.B1(_01137_),
    .Y(_01184_),
    .A1(_01178_),
    .A2(_01183_));
 sg13g2_a21oi_1 _22951_ (.A1(_01179_),
    .A2(_01184_),
    .Y(_01185_),
    .B1(net137));
 sg13g2_nand2_1 _22952_ (.Y(_01186_),
    .A(_02593_),
    .B(_13108_));
 sg13g2_nor2_1 _22953_ (.A(_01137_),
    .B(_01186_),
    .Y(_01187_));
 sg13g2_nor3_1 _22954_ (.A(_01137_),
    .B(net372),
    .C(net447),
    .Y(_01188_));
 sg13g2_nor3_1 _22955_ (.A(_12791_),
    .B(_01181_),
    .C(_01188_),
    .Y(_01189_));
 sg13g2_o21ai_1 _22956_ (.B1(net164),
    .Y(_01190_),
    .A1(_01187_),
    .A2(_01189_));
 sg13g2_nand2_1 _22957_ (.Y(_01191_),
    .A(_01138_),
    .B(net459));
 sg13g2_and2_1 _22958_ (.A(net707),
    .B(_12456_),
    .X(_01192_));
 sg13g2_nor2b_1 _22959_ (.A(net707),
    .B_N(net447),
    .Y(_01194_));
 sg13g2_o21ai_1 _22960_ (.B1(_01163_),
    .Y(_01195_),
    .A1(_01192_),
    .A2(_01194_));
 sg13g2_o21ai_1 _22961_ (.B1(_01195_),
    .Y(_01196_),
    .A1(_01186_),
    .A2(_01191_));
 sg13g2_nand3_1 _22962_ (.B(_12469_),
    .C(net165),
    .A(net208),
    .Y(_01197_));
 sg13g2_a21oi_1 _22963_ (.A1(_01179_),
    .A2(_01197_),
    .Y(_01198_),
    .B1(_12776_));
 sg13g2_a21oi_1 _22964_ (.A1(_12776_),
    .A2(_01196_),
    .Y(_01199_),
    .B1(_01198_));
 sg13g2_nand3b_1 _22965_ (.B(_01190_),
    .C(_01199_),
    .Y(_01200_),
    .A_N(_01185_));
 sg13g2_xnor2_1 _22966_ (.Y(_01201_),
    .A(_05065_),
    .B(_13077_));
 sg13g2_xor2_1 _22967_ (.B(_01201_),
    .A(net460),
    .X(_01202_));
 sg13g2_xnor2_1 _22968_ (.Y(_01203_),
    .A(net1085),
    .B(_01202_));
 sg13g2_o21ai_1 _22969_ (.B1(_00957_),
    .Y(_01205_),
    .A1(_12864_),
    .A2(_01202_));
 sg13g2_a21oi_1 _22970_ (.A1(_00953_),
    .A2(_01203_),
    .Y(_01206_),
    .B1(_01205_));
 sg13g2_xnor2_1 _22971_ (.Y(_01207_),
    .A(_01200_),
    .B(_01206_));
 sg13g2_nand2_1 _22972_ (.Y(_01208_),
    .A(net173),
    .B(_13061_));
 sg13g2_o21ai_1 _22973_ (.B1(_01208_),
    .Y(_01209_),
    .A1(net173),
    .A2(_13065_));
 sg13g2_a21oi_1 _22974_ (.A1(_12459_),
    .A2(_01209_),
    .Y(_01210_),
    .B1(_01187_));
 sg13g2_nor2b_1 _22975_ (.A(_01210_),
    .B_N(net164),
    .Y(_01211_));
 sg13g2_xnor2_1 _22976_ (.Y(_01212_),
    .A(_00972_),
    .B(_01202_));
 sg13g2_xnor2_1 _22977_ (.Y(_01213_),
    .A(_12459_),
    .B(_01201_));
 sg13g2_a221oi_1 _22978_ (.B2(_00967_),
    .C1(net170),
    .B1(_01213_),
    .A1(_01117_),
    .Y(_01214_),
    .A2(_01192_));
 sg13g2_o21ai_1 _22979_ (.B1(_01214_),
    .Y(_01216_),
    .A1(net209),
    .A2(_01212_));
 sg13g2_nor3_1 _22980_ (.A(_01207_),
    .B(_01211_),
    .C(_01216_),
    .Y(_01217_));
 sg13g2_a221oi_1 _22981_ (.B2(_00870_),
    .C1(_01217_),
    .B1(_06467_),
    .A1(_13111_),
    .Y(_01218_),
    .A2(net103));
 sg13g2_nor2b_1 _22982_ (.A(_11347_),
    .B_N(_00870_),
    .Y(_01219_));
 sg13g2_nor3_1 _22983_ (.A(net557),
    .B(_01218_),
    .C(_01219_),
    .Y(_00468_));
 sg13g2_nor2_1 _22984_ (.A(_08817_),
    .B(_12448_),
    .Y(_01220_));
 sg13g2_nand2_1 _22985_ (.Y(_01221_),
    .A(net44),
    .B(_01220_));
 sg13g2_xnor2_1 _22986_ (.Y(_01222_),
    .A(net1186),
    .B(_12829_));
 sg13g2_xor2_1 _22987_ (.B(_01222_),
    .A(_02226_),
    .X(_01223_));
 sg13g2_xnor2_1 _22988_ (.Y(_01224_),
    .A(net1018),
    .B(_01223_));
 sg13g2_xor2_1 _22989_ (.B(_01224_),
    .A(net1085),
    .X(_01226_));
 sg13g2_a22oi_1 _22990_ (.Y(_01227_),
    .B1(_01226_),
    .B2(net1183),
    .A2(_01224_),
    .A1(_12866_));
 sg13g2_nand2_1 _22991_ (.Y(_01228_),
    .A(net1018),
    .B(_00917_));
 sg13g2_nand4_1 _22992_ (.B(net1038),
    .C(net894),
    .A(net795),
    .Y(_01229_),
    .D(net372));
 sg13g2_o21ai_1 _22993_ (.B1(_01229_),
    .Y(_01230_),
    .A1(net451),
    .A2(_01228_));
 sg13g2_nand2b_1 _22994_ (.Y(_01231_),
    .B(_02593_),
    .A_N(_09178_));
 sg13g2_nor2_1 _22995_ (.A(net1038),
    .B(_02604_),
    .Y(_01232_));
 sg13g2_a21oi_1 _22996_ (.A1(net1038),
    .A2(_01231_),
    .Y(_01233_),
    .B1(_01232_));
 sg13g2_mux2_1 _22997_ (.A0(net1018),
    .A1(_02604_),
    .S(net1038),
    .X(_01234_));
 sg13g2_a22oi_1 _22998_ (.Y(_01235_),
    .B1(_01234_),
    .B2(_04352_),
    .A2(_00917_),
    .A1(net893));
 sg13g2_o21ai_1 _22999_ (.B1(_01235_),
    .Y(_01237_),
    .A1(net684),
    .A2(_01233_));
 sg13g2_nand2_1 _23000_ (.Y(_01238_),
    .A(net1018),
    .B(net372));
 sg13g2_nand2_1 _23001_ (.Y(_01239_),
    .A(net894),
    .B(net175));
 sg13g2_nand3_1 _23002_ (.B(_01238_),
    .C(_01239_),
    .A(net706),
    .Y(_01240_));
 sg13g2_inv_1 _23003_ (.Y(_01241_),
    .A(_00917_));
 sg13g2_nor2_1 _23004_ (.A(net1038),
    .B(_01231_),
    .Y(_01242_));
 sg13g2_a21oi_1 _23005_ (.A1(_09199_),
    .A2(_01241_),
    .Y(_01243_),
    .B1(_01242_));
 sg13g2_a21oi_1 _23006_ (.A1(_01240_),
    .A2(_01243_),
    .Y(_01244_),
    .B1(net211));
 sg13g2_a221oi_1 _23007_ (.B2(net211),
    .C1(_01244_),
    .B1(_01237_),
    .A1(net1042),
    .Y(_01245_),
    .A2(_01230_));
 sg13g2_buf_2 _23008_ (.A(_00191_),
    .X(_01246_));
 sg13g2_xnor2_1 _23009_ (.Y(_01248_),
    .A(net1183),
    .B(net1085));
 sg13g2_xor2_1 _23010_ (.B(_01248_),
    .A(_01224_),
    .X(_01249_));
 sg13g2_nor2_1 _23011_ (.A(_01246_),
    .B(_01249_),
    .Y(_01250_));
 sg13g2_nor2_1 _23012_ (.A(_01245_),
    .B(_01250_),
    .Y(_01251_));
 sg13g2_a21oi_1 _23013_ (.A1(net1038),
    .A2(net372),
    .Y(_01252_),
    .B1(net1018));
 sg13g2_a21o_1 _23014_ (.A2(_02226_),
    .A1(net1046),
    .B1(_01252_),
    .X(_01253_));
 sg13g2_nand2_1 _23015_ (.Y(_01254_),
    .A(net1042),
    .B(net684));
 sg13g2_a22oi_1 _23016_ (.Y(_01255_),
    .B1(_01254_),
    .B2(_00917_),
    .A2(_01253_),
    .A1(net894));
 sg13g2_o21ai_1 _23017_ (.B1(net684),
    .Y(_01256_),
    .A1(_04352_),
    .A2(_12831_));
 sg13g2_nand3_1 _23018_ (.B(_00917_),
    .C(_01256_),
    .A(net894),
    .Y(_01257_));
 sg13g2_o21ai_1 _23019_ (.B1(_01257_),
    .Y(_01259_),
    .A1(_12890_),
    .A2(_01255_));
 sg13g2_xnor2_1 _23020_ (.Y(_01260_),
    .A(_01227_),
    .B(_01250_));
 sg13g2_a221oi_1 _23021_ (.B2(_01260_),
    .C1(net100),
    .B1(_01259_),
    .A1(_01227_),
    .Y(_01261_),
    .A2(_01251_));
 sg13g2_xnor2_1 _23022_ (.Y(_01262_),
    .A(net209),
    .B(_01248_));
 sg13g2_xor2_1 _23023_ (.B(_01262_),
    .A(_01224_),
    .X(_01263_));
 sg13g2_a21oi_1 _23024_ (.A1(net113),
    .A2(_01263_),
    .Y(_01264_),
    .B1(net1035));
 sg13g2_or3_1 _23025_ (.A(_01220_),
    .B(_01261_),
    .C(_01264_),
    .X(_01265_));
 sg13g2_a21oi_1 _23026_ (.A1(_01221_),
    .A2(_01265_),
    .Y(_00469_),
    .B1(net440));
 sg13g2_nor2_1 _23027_ (.A(net795),
    .B(_03606_),
    .Y(_01266_));
 sg13g2_nand2_1 _23028_ (.Y(_01267_),
    .A(net364),
    .B(_01266_));
 sg13g2_nand4_1 _23029_ (.B(_12890_),
    .C(_04099_),
    .A(net1035),
    .Y(_01269_),
    .D(net894));
 sg13g2_o21ai_1 _23030_ (.B1(_01269_),
    .Y(_01270_),
    .A1(net1035),
    .A2(_01267_));
 sg13g2_nand2_1 _23031_ (.Y(_01271_),
    .A(net1036),
    .B(net893));
 sg13g2_mux2_1 _23032_ (.A0(net703),
    .A1(_01271_),
    .S(net451),
    .X(_01272_));
 sg13g2_mux2_1 _23033_ (.A0(_03530_),
    .A1(_03541_),
    .S(_12830_),
    .X(_01273_));
 sg13g2_nor2_1 _23034_ (.A(net1046),
    .B(_01273_),
    .Y(_01274_));
 sg13g2_a221oi_1 _23035_ (.B2(_03530_),
    .C1(_01274_),
    .B1(_01272_),
    .A1(net893),
    .Y(_01275_),
    .A2(_01266_));
 sg13g2_nand2_1 _23036_ (.Y(_01276_),
    .A(net1035),
    .B(_01275_));
 sg13g2_inv_2 _23037_ (.Y(_01277_),
    .A(net1184));
 sg13g2_or3_1 _23038_ (.A(net1046),
    .B(_03530_),
    .C(_01266_),
    .X(_01278_));
 sg13g2_nand2_1 _23039_ (.Y(_01280_),
    .A(net1034),
    .B(_03541_));
 sg13g2_o21ai_1 _23040_ (.B1(_01280_),
    .Y(_01281_),
    .A1(net703),
    .A2(net893));
 sg13g2_mux2_1 _23041_ (.A0(_01271_),
    .A1(_01281_),
    .S(net451),
    .X(_01282_));
 sg13g2_nand3_1 _23042_ (.B(_01278_),
    .C(_01282_),
    .A(_01277_),
    .Y(_01283_));
 sg13g2_a22oi_1 _23043_ (.Y(_01284_),
    .B1(_01276_),
    .B2(_01283_),
    .A2(_01270_),
    .A1(net710));
 sg13g2_xnor2_1 _23044_ (.Y(_01285_),
    .A(_12830_),
    .B(net1036));
 sg13g2_xnor2_1 _23045_ (.Y(_01286_),
    .A(_02841_),
    .B(_01285_));
 sg13g2_xnor2_1 _23046_ (.Y(_01287_),
    .A(net1034),
    .B(_01286_));
 sg13g2_xor2_1 _23047_ (.B(_01287_),
    .A(net1085),
    .X(_01288_));
 sg13g2_o21ai_1 _23048_ (.B1(_01288_),
    .Y(_01289_),
    .A1(net1037),
    .A2(_12979_));
 sg13g2_and2_1 _23049_ (.A(_12866_),
    .B(_01287_),
    .X(_01291_));
 sg13g2_a21oi_1 _23050_ (.A1(net1037),
    .A2(_12979_),
    .Y(_01292_),
    .B1(_01291_));
 sg13g2_nand2_1 _23051_ (.Y(_01293_),
    .A(_01289_),
    .B(_01292_));
 sg13g2_xnor2_1 _23052_ (.Y(_01294_),
    .A(_01284_),
    .B(_01293_));
 sg13g2_and2_1 _23053_ (.A(_12979_),
    .B(_01248_),
    .X(_01295_));
 sg13g2_nor2_1 _23054_ (.A(_04352_),
    .B(_01285_),
    .Y(_01296_));
 sg13g2_nand2_1 _23055_ (.Y(_01297_),
    .A(_12849_),
    .B(net367));
 sg13g2_nor2_1 _23056_ (.A(net1042),
    .B(_01297_),
    .Y(_01298_));
 sg13g2_o21ai_1 _23057_ (.B1(net364),
    .Y(_01299_),
    .A1(_01296_),
    .A2(_01298_));
 sg13g2_o21ai_1 _23058_ (.B1(_01299_),
    .Y(_01300_),
    .A1(_12831_),
    .A2(_01271_));
 sg13g2_nor3_1 _23059_ (.A(net1035),
    .B(_09240_),
    .C(_01297_),
    .Y(_01302_));
 sg13g2_a221oi_1 _23060_ (.B2(net1035),
    .C1(_01302_),
    .B1(_01300_),
    .A1(_01291_),
    .Y(_01303_),
    .A2(_01295_));
 sg13g2_a21oi_1 _23061_ (.A1(_01294_),
    .A2(_01303_),
    .Y(_01304_),
    .B1(net79));
 sg13g2_xnor2_1 _23062_ (.Y(_01305_),
    .A(_12893_),
    .B(_01248_));
 sg13g2_xnor2_1 _23063_ (.Y(_01306_),
    .A(_01287_),
    .B(_01305_));
 sg13g2_a21oi_1 _23064_ (.A1(net112),
    .A2(_01306_),
    .Y(_01307_),
    .B1(net135));
 sg13g2_nor2b_1 _23065_ (.A(_12448_),
    .B_N(_05748_),
    .Y(_01308_));
 sg13g2_nand2_1 _23066_ (.Y(_01309_),
    .A(net327),
    .B(_01308_));
 sg13g2_nand2_1 _23067_ (.Y(_01310_),
    .A(net1197),
    .B(_01309_));
 sg13g2_buf_2 _23068_ (.A(_01310_),
    .X(_01311_));
 sg13g2_or2_1 _23069_ (.X(_01313_),
    .B(_01311_),
    .A(_01307_));
 sg13g2_nand2_1 _23070_ (.Y(_01314_),
    .A(net1002),
    .B(_01220_));
 sg13g2_nand2b_1 _23071_ (.Y(_01315_),
    .B(net42),
    .A_N(_01314_));
 sg13g2_o21ai_1 _23072_ (.B1(_01315_),
    .Y(_00470_),
    .A1(_01304_),
    .A2(_01313_));
 sg13g2_nor2_1 _23073_ (.A(_12908_),
    .B(net698),
    .Y(_01316_));
 sg13g2_and2_1 _23074_ (.A(_12892_),
    .B(net1030),
    .X(_01317_));
 sg13g2_xor2_1 _23075_ (.B(net1030),
    .A(net791),
    .X(_01318_));
 sg13g2_nand2_1 _23076_ (.Y(_01319_),
    .A(net1034),
    .B(_01318_));
 sg13g2_o21ai_1 _23077_ (.B1(_01319_),
    .Y(_01320_),
    .A1(net1031),
    .A2(_01317_));
 sg13g2_a22oi_1 _23078_ (.Y(_01321_),
    .B1(_01320_),
    .B2(net1182),
    .A2(_01316_),
    .A1(_09310_));
 sg13g2_a21oi_1 _23079_ (.A1(_02669_),
    .A2(net705),
    .Y(_01323_),
    .B1(net700));
 sg13g2_nand3b_1 _23080_ (.B(_01316_),
    .C(net1182),
    .Y(_01324_),
    .A_N(_01323_));
 sg13g2_o21ai_1 _23081_ (.B1(_01324_),
    .Y(_01325_),
    .A1(net135),
    .A2(_01321_));
 sg13g2_nor2_1 _23082_ (.A(net1042),
    .B(_13052_),
    .Y(_01326_));
 sg13g2_xnor2_1 _23083_ (.Y(_01327_),
    .A(_03174_),
    .B(_12891_));
 sg13g2_xnor2_1 _23084_ (.Y(_01328_),
    .A(_04506_),
    .B(_01327_));
 sg13g2_xor2_1 _23085_ (.B(_01328_),
    .A(_02658_),
    .X(_01329_));
 sg13g2_xnor2_1 _23086_ (.Y(_01330_),
    .A(_12849_),
    .B(_01329_));
 sg13g2_a22oi_1 _23087_ (.Y(_01331_),
    .B1(_12949_),
    .B2(_01329_),
    .A2(_13052_),
    .A1(net1042));
 sg13g2_o21ai_1 _23088_ (.B1(_01331_),
    .Y(_01332_),
    .A1(_01326_),
    .A2(_01330_));
 sg13g2_xnor2_1 _23089_ (.Y(_01334_),
    .A(_01325_),
    .B(_01332_));
 sg13g2_and2_1 _23090_ (.A(_12949_),
    .B(_01329_),
    .X(_01335_));
 sg13g2_and2_1 _23091_ (.A(_13052_),
    .B(_01222_),
    .X(_01336_));
 sg13g2_nand2_1 _23092_ (.Y(_01337_),
    .A(net791),
    .B(net698));
 sg13g2_o21ai_1 _23093_ (.B1(_01319_),
    .Y(_01338_),
    .A1(net705),
    .A2(_01337_));
 sg13g2_nand2_1 _23094_ (.Y(_01339_),
    .A(net697),
    .B(_01338_));
 sg13g2_o21ai_1 _23095_ (.B1(_01339_),
    .Y(_01340_),
    .A1(net1182),
    .A2(_01337_));
 sg13g2_nor4_1 _23096_ (.A(_00875_),
    .B(_03530_),
    .C(_12893_),
    .D(_04516_),
    .Y(_01341_));
 sg13g2_a221oi_1 _23097_ (.B2(_00875_),
    .C1(_01341_),
    .B1(_01340_),
    .A1(_01335_),
    .Y(_01342_),
    .A2(_01336_));
 sg13g2_a21oi_1 _23098_ (.A1(_01334_),
    .A2(_01342_),
    .Y(_01343_),
    .B1(net97));
 sg13g2_xor2_1 _23099_ (.B(_01222_),
    .A(net449),
    .X(_01345_));
 sg13g2_xnor2_1 _23100_ (.Y(_01346_),
    .A(_01329_),
    .B(_01345_));
 sg13g2_a21oi_1 _23101_ (.A1(net66),
    .A2(_01346_),
    .Y(_01347_),
    .B1(net169));
 sg13g2_or3_1 _23102_ (.A(_01311_),
    .B(_01343_),
    .C(_01347_),
    .X(_01348_));
 sg13g2_o21ai_1 _23103_ (.B1(_01348_),
    .Y(_00471_),
    .A1(net35),
    .A2(_01314_));
 sg13g2_nor2_1 _23104_ (.A(net694),
    .B(_12962_),
    .Y(_01349_));
 sg13g2_nand2_1 _23105_ (.Y(_01350_),
    .A(net1027),
    .B(net790));
 sg13g2_inv_1 _23106_ (.Y(_01351_),
    .A(_01350_));
 sg13g2_xor2_1 _23107_ (.B(_12938_),
    .A(net1027),
    .X(_01352_));
 sg13g2_nand2_1 _23108_ (.Y(_01353_),
    .A(net1031),
    .B(_01352_));
 sg13g2_o21ai_1 _23109_ (.B1(_01353_),
    .Y(_01355_),
    .A1(net1028),
    .A2(_01351_));
 sg13g2_a22oi_1 _23110_ (.Y(_01356_),
    .B1(_01355_),
    .B2(net1181),
    .A2(_01349_),
    .A1(_09350_));
 sg13g2_nand2_1 _23111_ (.Y(_01357_),
    .A(net1028),
    .B(_04313_));
 sg13g2_nand3_1 _23112_ (.B(_01349_),
    .C(_01357_),
    .A(net1181),
    .Y(_01358_));
 sg13g2_o21ai_1 _23113_ (.B1(_01358_),
    .Y(_01359_),
    .A1(net169),
    .A2(_01356_));
 sg13g2_nor2_1 _23114_ (.A(net364),
    .B(_13088_),
    .Y(_01360_));
 sg13g2_xnor2_1 _23115_ (.Y(_01361_),
    .A(_04131_),
    .B(_12937_));
 sg13g2_xnor2_1 _23116_ (.Y(_01362_),
    .A(_04748_),
    .B(_01361_));
 sg13g2_xnor2_1 _23117_ (.Y(_01363_),
    .A(net1036),
    .B(_01362_));
 sg13g2_xnor2_1 _23118_ (.Y(_01364_),
    .A(_12908_),
    .B(_01363_));
 sg13g2_a22oi_1 _23119_ (.Y(_01366_),
    .B1(_12979_),
    .B2(_01363_),
    .A2(_13088_),
    .A1(net364));
 sg13g2_o21ai_1 _23120_ (.B1(_01366_),
    .Y(_01367_),
    .A1(_01360_),
    .A2(_01364_));
 sg13g2_xnor2_1 _23121_ (.Y(_01368_),
    .A(_01359_),
    .B(_01367_));
 sg13g2_o21ai_1 _23122_ (.B1(_01353_),
    .Y(_01369_),
    .A1(net697),
    .A2(_01350_));
 sg13g2_nand2_1 _23123_ (.Y(_01370_),
    .A(net695),
    .B(_01369_));
 sg13g2_o21ai_1 _23124_ (.B1(_01370_),
    .Y(_01371_),
    .A1(net1181),
    .A2(_01350_));
 sg13g2_and2_1 _23125_ (.A(_13088_),
    .B(_01327_),
    .X(_01372_));
 sg13g2_and2_1 _23126_ (.A(_12979_),
    .B(_01363_),
    .X(_01373_));
 sg13g2_nor3_1 _23127_ (.A(_04109_),
    .B(_09350_),
    .C(_01350_),
    .Y(_01374_));
 sg13g2_a221oi_1 _23128_ (.B2(_01373_),
    .C1(_01374_),
    .B1(_01372_),
    .A1(net169),
    .Y(_01375_),
    .A2(_01371_));
 sg13g2_a21oi_1 _23129_ (.A1(_01368_),
    .A2(_01375_),
    .Y(_01377_),
    .B1(net97));
 sg13g2_xnor2_1 _23130_ (.Y(_01378_),
    .A(_13021_),
    .B(_01327_));
 sg13g2_xnor2_1 _23131_ (.Y(_01379_),
    .A(_01363_),
    .B(_01378_));
 sg13g2_a21oi_1 _23132_ (.A1(net66),
    .A2(_01379_),
    .Y(_01380_),
    .B1(net365));
 sg13g2_or3_1 _23133_ (.A(_01311_),
    .B(_01377_),
    .C(_01380_),
    .X(_01381_));
 sg13g2_o21ai_1 _23134_ (.B1(_01381_),
    .Y(_00472_),
    .A1(net26),
    .A2(_01309_));
 sg13g2_nand3_1 _23135_ (.B(net698),
    .C(_12993_),
    .A(_05064_),
    .Y(_01382_));
 sg13g2_xor2_1 _23136_ (.B(_12981_),
    .A(_04163_),
    .X(_01383_));
 sg13g2_nand2_1 _23137_ (.Y(_01384_),
    .A(net687),
    .B(_01383_));
 sg13g2_o21ai_1 _23138_ (.B1(_01384_),
    .Y(_01385_),
    .A1(net687),
    .A2(_01038_));
 sg13g2_nand2_1 _23139_ (.Y(_01387_),
    .A(net695),
    .B(_01385_));
 sg13g2_o21ai_1 _23140_ (.B1(_01387_),
    .Y(_01388_),
    .A1(net695),
    .A2(_01382_));
 sg13g2_xnor2_1 _23141_ (.Y(_01389_),
    .A(net1180),
    .B(_12981_));
 sg13g2_xor2_1 _23142_ (.B(_04163_),
    .A(_04948_),
    .X(_01390_));
 sg13g2_xnor2_1 _23143_ (.Y(_01391_),
    .A(_01389_),
    .B(_01390_));
 sg13g2_xnor2_1 _23144_ (.Y(_01392_),
    .A(net1179),
    .B(_01391_));
 sg13g2_nor2_1 _23145_ (.A(_13029_),
    .B(_01392_),
    .Y(_01393_));
 sg13g2_and2_1 _23146_ (.A(_13130_),
    .B(_01361_),
    .X(_01394_));
 sg13g2_nor2_1 _23147_ (.A(_04857_),
    .B(_01382_),
    .Y(_01395_));
 sg13g2_a221oi_1 _23148_ (.B2(_01394_),
    .C1(_01395_),
    .B1(_01393_),
    .A1(net685),
    .Y(_01396_),
    .A2(_01388_));
 sg13g2_nand2_1 _23149_ (.Y(_01398_),
    .A(_13129_),
    .B(net700));
 sg13g2_xnor2_1 _23150_ (.Y(_01399_),
    .A(_12962_),
    .B(_01392_));
 sg13g2_nand2_1 _23151_ (.Y(_01400_),
    .A(_13130_),
    .B(net697));
 sg13g2_o21ai_1 _23152_ (.B1(_01400_),
    .Y(_01401_),
    .A1(_13029_),
    .A2(_01392_));
 sg13g2_a21oi_1 _23153_ (.A1(_01398_),
    .A2(_01399_),
    .Y(_01402_),
    .B1(_01401_));
 sg13g2_a21oi_1 _23154_ (.A1(net1028),
    .A2(_05014_),
    .Y(_01403_),
    .B1(_05101_));
 sg13g2_a22oi_1 _23155_ (.Y(_01404_),
    .B1(_01383_),
    .B2(net1180),
    .A2(_01038_),
    .A1(_05101_));
 sg13g2_or2_1 _23156_ (.X(_01405_),
    .B(_01404_),
    .A(_05014_));
 sg13g2_o21ai_1 _23157_ (.B1(_01405_),
    .Y(_01406_),
    .A1(_01020_),
    .A2(_01403_));
 sg13g2_nor2_1 _23158_ (.A(net361),
    .B(_01020_),
    .Y(_01407_));
 sg13g2_a22oi_1 _23159_ (.Y(_01409_),
    .B1(_01407_),
    .B2(_09392_),
    .A2(_01406_),
    .A1(_04857_));
 sg13g2_xnor2_1 _23160_ (.Y(_01410_),
    .A(_01402_),
    .B(_01409_));
 sg13g2_a21oi_1 _23161_ (.A1(_01396_),
    .A2(_01410_),
    .Y(_01411_),
    .B1(net97));
 sg13g2_xnor2_1 _23162_ (.Y(_01412_),
    .A(net448),
    .B(_01361_));
 sg13g2_xnor2_1 _23163_ (.Y(_01413_),
    .A(_01392_),
    .B(_01412_));
 sg13g2_a21oi_1 _23164_ (.A1(net66),
    .A2(_01413_),
    .Y(_01414_),
    .B1(net363));
 sg13g2_or3_1 _23165_ (.A(_01311_),
    .B(_01411_),
    .C(_01414_),
    .X(_01415_));
 sg13g2_o21ai_1 _23166_ (.B1(_01415_),
    .Y(_00473_),
    .A1(net29),
    .A2(_01314_));
 sg13g2_nand3_1 _23167_ (.B(net694),
    .C(net448),
    .A(net358),
    .Y(_01416_));
 sg13g2_xor2_1 _23168_ (.B(_13016_),
    .A(_04779_),
    .X(_01417_));
 sg13g2_nand2_1 _23169_ (.Y(_01419_),
    .A(net358),
    .B(_01417_));
 sg13g2_o21ai_1 _23170_ (.B1(_01419_),
    .Y(_01420_),
    .A1(net358),
    .A2(_01056_));
 sg13g2_nand2_1 _23171_ (.Y(_01421_),
    .A(net685),
    .B(_01420_));
 sg13g2_o21ai_1 _23172_ (.B1(_01421_),
    .Y(_01422_),
    .A1(net685),
    .A2(_01416_));
 sg13g2_xnor2_1 _23173_ (.Y(_01423_),
    .A(net1179),
    .B(_13014_));
 sg13g2_xor2_1 _23174_ (.B(net1027),
    .A(net1020),
    .X(_01424_));
 sg13g2_xnor2_1 _23175_ (.Y(_01425_),
    .A(_01423_),
    .B(_01424_));
 sg13g2_xnor2_1 _23176_ (.Y(_01426_),
    .A(net1019),
    .B(_01425_));
 sg13g2_nor2_1 _23177_ (.A(_13087_),
    .B(_01426_),
    .Y(_01427_));
 sg13g2_buf_1 _23178_ (.A(_00159_),
    .X(_01428_));
 sg13g2_nor2b_1 _23179_ (.A(_01428_),
    .B_N(_01389_),
    .Y(_01430_));
 sg13g2_nor2_1 _23180_ (.A(_04946_),
    .B(_01416_),
    .Y(_01431_));
 sg13g2_a221oi_1 _23181_ (.B2(_01430_),
    .C1(_01431_),
    .B1(_01427_),
    .A1(net360),
    .Y(_01432_),
    .A2(_01422_));
 sg13g2_nand2_1 _23182_ (.Y(_01433_),
    .A(_01428_),
    .B(_04830_));
 sg13g2_xnor2_1 _23183_ (.Y(_01434_),
    .A(_12993_),
    .B(_01426_));
 sg13g2_nand2b_1 _23184_ (.Y(_01435_),
    .B(net1028),
    .A_N(_01428_));
 sg13g2_o21ai_1 _23185_ (.B1(_01435_),
    .Y(_01436_),
    .A1(_13087_),
    .A2(_01426_));
 sg13g2_a21oi_1 _23186_ (.A1(_01433_),
    .A2(_01434_),
    .Y(_01437_),
    .B1(_01436_));
 sg13g2_a22oi_1 _23187_ (.Y(_01438_),
    .B1(_01417_),
    .B2(net1023),
    .A2(_01056_),
    .A1(net683));
 sg13g2_a21oi_1 _23188_ (.A1(net1023),
    .A2(_05013_),
    .Y(_01439_),
    .B1(net683));
 sg13g2_or3_1 _23189_ (.A(net694),
    .B(_13025_),
    .C(_01439_),
    .X(_01441_));
 sg13g2_o21ai_1 _23190_ (.B1(_01441_),
    .Y(_01442_),
    .A1(_05074_),
    .A2(_01438_));
 sg13g2_nor3_1 _23191_ (.A(net358),
    .B(_04789_),
    .C(_13025_),
    .Y(_01443_));
 sg13g2_a22oi_1 _23192_ (.Y(_01444_),
    .B1(_01443_),
    .B2(_09406_),
    .A2(_01442_),
    .A1(_04946_));
 sg13g2_xnor2_1 _23193_ (.Y(_01445_),
    .A(_01437_),
    .B(_01444_));
 sg13g2_a21oi_1 _23194_ (.A1(_01432_),
    .A2(_01445_),
    .Y(_01446_),
    .B1(net97));
 sg13g2_xnor2_1 _23195_ (.Y(_01447_),
    .A(_13112_),
    .B(_01389_));
 sg13g2_xnor2_1 _23196_ (.Y(_01448_),
    .A(_01426_),
    .B(_01447_));
 sg13g2_a21oi_1 _23197_ (.A1(net66),
    .A2(_01448_),
    .Y(_01449_),
    .B1(_05064_));
 sg13g2_or3_1 _23198_ (.A(_01311_),
    .B(_01446_),
    .C(_01449_),
    .X(_01450_));
 sg13g2_o21ai_1 _23199_ (.B1(_01450_),
    .Y(_00474_),
    .A1(net43),
    .A2(_01314_));
 sg13g2_nor2_1 _23200_ (.A(net1021),
    .B(_02615_),
    .Y(_01452_));
 sg13g2_and2_1 _23201_ (.A(net1024),
    .B(_13062_),
    .X(_01453_));
 sg13g2_buf_1 _23202_ (.A(_01453_),
    .X(_01454_));
 sg13g2_nand2_1 _23203_ (.Y(_01455_),
    .A(_02647_),
    .B(net361));
 sg13g2_xnor2_1 _23204_ (.Y(_01456_),
    .A(net1039),
    .B(net1024));
 sg13g2_mux2_1 _23205_ (.A0(_01455_),
    .A1(_01456_),
    .S(net208),
    .X(_01457_));
 sg13g2_nand3_1 _23206_ (.B(net361),
    .C(_01181_),
    .A(net683),
    .Y(_01458_));
 sg13g2_o21ai_1 _23207_ (.B1(_01458_),
    .Y(_01459_),
    .A1(net683),
    .A2(_01457_));
 sg13g2_a221oi_1 _23208_ (.B2(net359),
    .C1(net102),
    .B1(_01459_),
    .A1(_01452_),
    .Y(_01460_),
    .A2(_01454_));
 sg13g2_inv_1 _23209_ (.Y(_01461_),
    .A(_01246_));
 sg13g2_xnor2_1 _23210_ (.Y(_01462_),
    .A(_09463_),
    .B(_01456_));
 sg13g2_xnor2_1 _23211_ (.Y(_01463_),
    .A(net447),
    .B(_01462_));
 sg13g2_and2_1 _23212_ (.A(_13130_),
    .B(_01463_),
    .X(_01464_));
 sg13g2_nand3_1 _23213_ (.B(_01423_),
    .C(_01464_),
    .A(_01461_),
    .Y(_01465_));
 sg13g2_xnor2_1 _23214_ (.Y(_01466_),
    .A(_13111_),
    .B(_01423_));
 sg13g2_xnor2_1 _23215_ (.Y(_01467_),
    .A(_01463_),
    .B(_01466_));
 sg13g2_nand2b_1 _23216_ (.Y(_01468_),
    .B(_01467_),
    .A_N(net164));
 sg13g2_xor2_1 _23217_ (.B(net173),
    .A(net1021),
    .X(_01469_));
 sg13g2_nand3_1 _23218_ (.B(_02636_),
    .C(_01119_),
    .A(net1021),
    .Y(_01470_));
 sg13g2_o21ai_1 _23219_ (.B1(_01470_),
    .Y(_01472_),
    .A1(net1021),
    .A2(_01119_));
 sg13g2_a21oi_1 _23220_ (.A1(_01102_),
    .A2(_01469_),
    .Y(_01473_),
    .B1(_01472_));
 sg13g2_nand2b_1 _23221_ (.Y(_01474_),
    .B(net175),
    .A_N(_01102_));
 sg13g2_o21ai_1 _23222_ (.B1(_01474_),
    .Y(_01475_),
    .A1(_01238_),
    .A2(_01119_));
 sg13g2_o21ai_1 _23223_ (.B1(_01102_),
    .Y(_01476_),
    .A1(_02636_),
    .A2(_01454_));
 sg13g2_nand2_1 _23224_ (.Y(_01477_),
    .A(net1021),
    .B(_01476_));
 sg13g2_a21oi_1 _23225_ (.A1(_01474_),
    .A2(_01477_),
    .Y(_01478_),
    .B1(net684));
 sg13g2_a221oi_1 _23226_ (.B2(net683),
    .C1(_01478_),
    .B1(_01475_),
    .A1(_01452_),
    .Y(_01479_),
    .A2(_01454_));
 sg13g2_o21ai_1 _23227_ (.B1(_01479_),
    .Y(_01480_),
    .A1(_09449_),
    .A2(_01473_));
 sg13g2_xnor2_1 _23228_ (.Y(_01481_),
    .A(_13019_),
    .B(_01463_));
 sg13g2_o21ai_1 _23229_ (.B1(_01481_),
    .Y(_01483_),
    .A1(_01461_),
    .A2(net685));
 sg13g2_a21oi_1 _23230_ (.A1(_01461_),
    .A2(net685),
    .Y(_01484_),
    .B1(_01464_));
 sg13g2_nand2_1 _23231_ (.Y(_01485_),
    .A(_01483_),
    .B(_01484_));
 sg13g2_xnor2_1 _23232_ (.Y(_01486_),
    .A(_01480_),
    .B(_01485_));
 sg13g2_nand4_1 _23233_ (.B(_01465_),
    .C(_01468_),
    .A(_01460_),
    .Y(_01487_),
    .D(_01486_));
 sg13g2_a22oi_1 _23234_ (.Y(_01488_),
    .B1(net25),
    .B2(_01308_),
    .A2(net72),
    .A1(net164));
 sg13g2_a221oi_1 _23235_ (.B2(_01488_),
    .C1(_09818_),
    .B1(_01487_),
    .A1(net24),
    .Y(_00475_),
    .A2(_01308_));
 sg13g2_nand2_1 _23236_ (.Y(_01489_),
    .A(_05012_),
    .B(_13060_));
 sg13g2_buf_2 _23237_ (.A(_01489_),
    .X(_01490_));
 sg13g2_nor2_1 _23238_ (.A(net1184),
    .B(_01490_),
    .Y(_01491_));
 sg13g2_nor2_1 _23239_ (.A(net1020),
    .B(_13060_),
    .Y(_01493_));
 sg13g2_xnor2_1 _23240_ (.Y(_01494_),
    .A(net1184),
    .B(net1178));
 sg13g2_nand3_1 _23241_ (.B(net1178),
    .C(_01490_),
    .A(_02830_),
    .Y(_01495_));
 sg13g2_o21ai_1 _23242_ (.B1(_01495_),
    .Y(_01496_),
    .A1(_01493_),
    .A2(_01494_));
 sg13g2_nor2_1 _23243_ (.A(_01491_),
    .B(_01496_),
    .Y(_01497_));
 sg13g2_nor3_1 _23244_ (.A(_01277_),
    .B(_09198_),
    .C(_01490_),
    .Y(_01498_));
 sg13g2_a21o_1 _23245_ (.A2(_01493_),
    .A1(_01277_),
    .B1(_01498_),
    .X(_01499_));
 sg13g2_a21oi_1 _23246_ (.A1(net1178),
    .A2(_01490_),
    .Y(_01500_),
    .B1(_01493_));
 sg13g2_nand2_1 _23247_ (.Y(_01501_),
    .A(net1178),
    .B(_01493_));
 sg13g2_o21ai_1 _23248_ (.B1(_01501_),
    .Y(_01502_),
    .A1(_02830_),
    .A2(_01500_));
 sg13g2_nor3_1 _23249_ (.A(_01277_),
    .B(net1178),
    .C(_01490_),
    .Y(_01504_));
 sg13g2_a221oi_1 _23250_ (.B2(_09198_),
    .C1(_01504_),
    .B1(_01502_),
    .A1(net683),
    .Y(_01505_),
    .A2(_01499_));
 sg13g2_o21ai_1 _23251_ (.B1(_01505_),
    .Y(_01506_),
    .A1(_09449_),
    .A2(_01497_));
 sg13g2_buf_1 _23252_ (.A(_01506_),
    .X(_01507_));
 sg13g2_nor2_1 _23253_ (.A(net1183),
    .B(_01461_),
    .Y(_01508_));
 sg13g2_nor2b_1 _23254_ (.A(_01246_),
    .B_N(net1085),
    .Y(_01509_));
 sg13g2_nand2b_1 _23255_ (.Y(_01510_),
    .B(_01246_),
    .A_N(net792));
 sg13g2_o21ai_1 _23256_ (.B1(_01510_),
    .Y(_01511_),
    .A1(net1037),
    .A2(_01509_));
 sg13g2_xnor2_1 _23257_ (.Y(_01512_),
    .A(_05012_),
    .B(_13060_));
 sg13g2_xnor2_1 _23258_ (.Y(_01513_),
    .A(_09463_),
    .B(_01512_));
 sg13g2_xnor2_1 _23259_ (.Y(_01515_),
    .A(_01277_),
    .B(_01513_));
 sg13g2_buf_2 _23260_ (.A(_01515_),
    .X(_01516_));
 sg13g2_a22oi_1 _23261_ (.Y(_01517_),
    .B1(_01511_),
    .B2(_01516_),
    .A2(_01508_),
    .A1(net793));
 sg13g2_a21o_1 _23262_ (.A2(_01516_),
    .A1(net792),
    .B1(_01461_),
    .X(_01518_));
 sg13g2_a221oi_1 _23263_ (.B2(_01516_),
    .C1(_01507_),
    .B1(_01509_),
    .A1(net1037),
    .Y(_01519_),
    .A2(_01518_));
 sg13g2_a21o_1 _23264_ (.A2(_01517_),
    .A1(_01507_),
    .B1(_01519_),
    .X(_01520_));
 sg13g2_xor2_1 _23265_ (.B(_01516_),
    .A(_01262_),
    .X(_01521_));
 sg13g2_o21ai_1 _23266_ (.B1(net175),
    .Y(_01522_),
    .A1(net105),
    .A2(_01521_));
 sg13g2_nand2b_1 _23267_ (.Y(_01523_),
    .B(net686),
    .A_N(_01512_));
 sg13g2_o21ai_1 _23268_ (.B1(_01523_),
    .Y(_01524_),
    .A1(net686),
    .A2(_01490_));
 sg13g2_nor2_1 _23269_ (.A(net689),
    .B(_01490_),
    .Y(_01526_));
 sg13g2_a21oi_1 _23270_ (.A1(net359),
    .A2(_01524_),
    .Y(_01527_),
    .B1(_01526_));
 sg13g2_nor2_1 _23271_ (.A(_01277_),
    .B(_01527_),
    .Y(_01528_));
 sg13g2_nand3_1 _23272_ (.B(_12866_),
    .C(_01509_),
    .A(net1037),
    .Y(_01529_));
 sg13g2_nor2_1 _23273_ (.A(_01516_),
    .B(_01529_),
    .Y(_01530_));
 sg13g2_nor3_1 _23274_ (.A(net1035),
    .B(_09449_),
    .C(_01490_),
    .Y(_01531_));
 sg13g2_nor4_1 _23275_ (.A(_01311_),
    .B(_01528_),
    .C(_01530_),
    .D(_01531_),
    .Y(_01532_));
 sg13g2_nand3_1 _23276_ (.B(_01522_),
    .C(_01532_),
    .A(_01520_),
    .Y(_01533_));
 sg13g2_and2_1 _23277_ (.A(net792),
    .B(net793),
    .X(_01534_));
 sg13g2_nor2_1 _23278_ (.A(net792),
    .B(_01246_),
    .Y(_01535_));
 sg13g2_a22oi_1 _23279_ (.Y(_01537_),
    .B1(_01535_),
    .B2(_12866_),
    .A2(_01534_),
    .A1(_01507_));
 sg13g2_o21ai_1 _23280_ (.B1(net793),
    .Y(_01538_),
    .A1(_12884_),
    .A2(_01508_));
 sg13g2_inv_1 _23281_ (.Y(_01539_),
    .A(_01538_));
 sg13g2_nand3_1 _23282_ (.B(_01246_),
    .C(net793),
    .A(net792),
    .Y(_01540_));
 sg13g2_mux2_1 _23283_ (.A0(_01539_),
    .A1(_01540_),
    .S(_01507_),
    .X(_01541_));
 sg13g2_o21ai_1 _23284_ (.B1(_01541_),
    .Y(_01542_),
    .A1(net1037),
    .A2(_01537_));
 sg13g2_nor2b_1 _23285_ (.A(_01516_),
    .B_N(_01542_),
    .Y(_01543_));
 sg13g2_nand3_1 _23286_ (.B(net110),
    .C(_01309_),
    .A(net173),
    .Y(_01544_));
 sg13g2_o21ai_1 _23287_ (.B1(_01544_),
    .Y(_01545_),
    .A1(net121),
    .A2(_01309_));
 sg13g2_nand2_1 _23288_ (.Y(_01546_),
    .A(net356),
    .B(_01545_));
 sg13g2_o21ai_1 _23289_ (.B1(_01546_),
    .Y(_00476_),
    .A1(_01533_),
    .A2(_01543_));
 sg13g2_or2_1 _23290_ (.X(_01548_),
    .B(_13185_),
    .A(_08817_));
 sg13g2_buf_1 _23291_ (.A(_01548_),
    .X(_01549_));
 sg13g2_buf_1 _23292_ (.A(_01549_),
    .X(_01550_));
 sg13g2_buf_1 _23293_ (.A(_13229_),
    .X(_01551_));
 sg13g2_buf_1 _23294_ (.A(\grid.cell_3_0.se ),
    .X(_01552_));
 sg13g2_buf_1 _23295_ (.A(net1081),
    .X(_01553_));
 sg13g2_buf_1 _23296_ (.A(net776),
    .X(_01554_));
 sg13g2_buf_2 _23297_ (.A(\grid.cell_3_0.sw ),
    .X(_01555_));
 sg13g2_buf_1 _23298_ (.A(_01555_),
    .X(_01556_));
 sg13g2_nor2_1 _23299_ (.A(net785),
    .B(net775),
    .Y(_01558_));
 sg13g2_buf_2 _23300_ (.A(_01558_),
    .X(_01559_));
 sg13g2_inv_1 _23301_ (.Y(_01560_),
    .A(_01559_));
 sg13g2_and2_1 _23302_ (.A(_13192_),
    .B(_01555_),
    .X(_01561_));
 sg13g2_buf_1 _23303_ (.A(_01561_),
    .X(_01562_));
 sg13g2_nand3_1 _23304_ (.B(_09185_),
    .C(_01562_),
    .A(net776),
    .Y(_01563_));
 sg13g2_o21ai_1 _23305_ (.B1(_01563_),
    .Y(_01564_),
    .A1(net434),
    .A2(_01560_));
 sg13g2_nand2_1 _23306_ (.Y(_01565_),
    .A(net274),
    .B(_01564_));
 sg13g2_buf_1 _23307_ (.A(_01554_),
    .X(_01566_));
 sg13g2_nand3_1 _23308_ (.B(_09289_),
    .C(_01562_),
    .A(net204),
    .Y(_01567_));
 sg13g2_nand2_1 _23309_ (.Y(_01569_),
    .A(net785),
    .B(net775));
 sg13g2_buf_2 _23310_ (.A(_01569_),
    .X(_01570_));
 sg13g2_nor2_1 _23311_ (.A(net434),
    .B(_01570_),
    .Y(_01571_));
 sg13g2_xnor2_1 _23312_ (.Y(_01572_),
    .A(net776),
    .B(net1125));
 sg13g2_nand3_1 _23313_ (.B(net1125),
    .C(_01570_),
    .A(net776),
    .Y(_01573_));
 sg13g2_o21ai_1 _23314_ (.B1(_01573_),
    .Y(_01574_),
    .A1(_01559_),
    .A2(_01572_));
 sg13g2_o21ai_1 _23315_ (.B1(_09181_),
    .Y(_01575_),
    .A1(_01571_),
    .A2(_01574_));
 sg13g2_a21oi_1 _23316_ (.A1(net1125),
    .A2(_01570_),
    .Y(_01576_),
    .B1(_01559_));
 sg13g2_nand2_1 _23317_ (.Y(_01577_),
    .A(net1125),
    .B(_01559_));
 sg13g2_o21ai_1 _23318_ (.B1(_01577_),
    .Y(_01578_),
    .A1(net434),
    .A2(_01576_));
 sg13g2_nand2_1 _23319_ (.Y(_01580_),
    .A(net272),
    .B(_01578_));
 sg13g2_nand4_1 _23320_ (.B(_01567_),
    .C(_01575_),
    .A(_01565_),
    .Y(_01581_),
    .D(_01580_));
 sg13g2_buf_1 _23321_ (.A(_00268_),
    .X(_01582_));
 sg13g2_nand2_1 _23322_ (.Y(_01583_),
    .A(net892),
    .B(net1080));
 sg13g2_inv_2 _23323_ (.Y(_01584_),
    .A(_01556_));
 sg13g2_xnor2_1 _23324_ (.Y(_01585_),
    .A(_09173_),
    .B(net1081));
 sg13g2_xnor2_1 _23325_ (.Y(_01586_),
    .A(_13220_),
    .B(_01585_));
 sg13g2_xnor2_1 _23326_ (.Y(_01587_),
    .A(_01584_),
    .B(_01586_));
 sg13g2_xnor2_1 _23327_ (.Y(_01588_),
    .A(net446),
    .B(_01587_));
 sg13g2_inv_2 _23328_ (.Y(_01589_),
    .A(_01582_));
 sg13g2_nand2_1 _23329_ (.Y(_01591_),
    .A(net890),
    .B(_01589_));
 sg13g2_o21ai_1 _23330_ (.B1(_01591_),
    .Y(_01592_),
    .A1(net781),
    .A2(_01587_));
 sg13g2_a21oi_1 _23331_ (.A1(_01583_),
    .A2(_01588_),
    .Y(_01593_),
    .B1(_01592_));
 sg13g2_xor2_1 _23332_ (.B(_01593_),
    .A(_01581_),
    .X(_01594_));
 sg13g2_buf_2 _23333_ (.A(\grid.cell_3_0.s ),
    .X(_01595_));
 sg13g2_buf_1 _23334_ (.A(_01595_),
    .X(_01596_));
 sg13g2_xor2_1 _23335_ (.B(net786),
    .A(_09216_),
    .X(_01597_));
 sg13g2_xnor2_1 _23336_ (.Y(_01598_),
    .A(net774),
    .B(_01597_));
 sg13g2_xnor2_1 _23337_ (.Y(_01599_),
    .A(_01587_),
    .B(_01598_));
 sg13g2_buf_1 _23338_ (.A(_01556_),
    .X(_01600_));
 sg13g2_buf_1 _23339_ (.A(_01600_),
    .X(_01602_));
 sg13g2_nor2_1 _23340_ (.A(net274),
    .B(net776),
    .Y(_01603_));
 sg13g2_nand4_1 _23341_ (.B(net207),
    .C(net203),
    .A(net270),
    .Y(_01604_),
    .D(_01603_));
 sg13g2_xnor2_1 _23342_ (.Y(_01605_),
    .A(_13192_),
    .B(_01555_));
 sg13g2_nor2_1 _23343_ (.A(net274),
    .B(_01605_),
    .Y(_01606_));
 sg13g2_nor2_1 _23344_ (.A(net895),
    .B(_01570_),
    .Y(_01607_));
 sg13g2_o21ai_1 _23345_ (.B1(net270),
    .Y(_01608_),
    .A1(_01606_),
    .A2(_01607_));
 sg13g2_o21ai_1 _23346_ (.B1(_01608_),
    .Y(_01609_),
    .A1(_09288_),
    .A2(_01570_));
 sg13g2_nand2_1 _23347_ (.Y(_01610_),
    .A(net204),
    .B(_01609_));
 sg13g2_or4_1 _23348_ (.A(net1080),
    .B(net781),
    .C(_01587_),
    .D(_01597_),
    .X(_01611_));
 sg13g2_nand4_1 _23349_ (.B(_01604_),
    .C(_01610_),
    .A(net119),
    .Y(_01613_),
    .D(_01611_));
 sg13g2_a21oi_1 _23350_ (.A1(_13230_),
    .A2(_01599_),
    .Y(_01614_),
    .B1(_01613_));
 sg13g2_a22oi_1 _23351_ (.Y(_01615_),
    .B1(_01594_),
    .B2(_01614_),
    .A2(net67),
    .A1(net777));
 sg13g2_o21ai_1 _23352_ (.B1(_00977_),
    .Y(_01616_),
    .A1(_09235_),
    .A2(net36));
 sg13g2_a21oi_1 _23353_ (.A1(net36),
    .A2(_01615_),
    .Y(_00477_),
    .B1(_01616_));
 sg13g2_buf_8 _23354_ (.A(\grid.cell_3_1.se ),
    .X(_01617_));
 sg13g2_buf_1 _23355_ (.A(_01617_),
    .X(_01618_));
 sg13g2_buf_1 _23356_ (.A(net773),
    .X(_01619_));
 sg13g2_nand2_1 _23357_ (.Y(_01620_),
    .A(net443),
    .B(net432));
 sg13g2_xor2_1 _23358_ (.B(_01617_),
    .A(_13252_),
    .X(_01621_));
 sg13g2_and2_1 _23359_ (.A(net895),
    .B(_01621_),
    .X(_01623_));
 sg13g2_nor2_1 _23360_ (.A(net552),
    .B(_01620_),
    .Y(_01624_));
 sg13g2_o21ai_1 _23361_ (.B1(net268),
    .Y(_01625_),
    .A1(_01623_),
    .A2(_01624_));
 sg13g2_o21ai_1 _23362_ (.B1(_01625_),
    .Y(_01626_),
    .A1(net1125),
    .A2(_01620_));
 sg13g2_inv_2 _23363_ (.Y(_01627_),
    .A(_01617_));
 sg13g2_xnor2_1 _23364_ (.Y(_01628_),
    .A(_01627_),
    .B(_13304_));
 sg13g2_xnor2_1 _23365_ (.Y(_01629_),
    .A(_01585_),
    .B(_01628_));
 sg13g2_buf_1 _23366_ (.A(_01629_),
    .X(_01630_));
 sg13g2_xnor2_1 _23367_ (.Y(_01631_),
    .A(_13229_),
    .B(_01630_));
 sg13g2_o21ai_1 _23368_ (.B1(net892),
    .Y(_01632_),
    .A1(net1080),
    .A2(_01631_));
 sg13g2_nand2_1 _23369_ (.Y(_01634_),
    .A(net1080),
    .B(_01631_));
 sg13g2_nand2_1 _23370_ (.Y(_01635_),
    .A(net268),
    .B(_01603_));
 sg13g2_nor2_1 _23371_ (.A(net783),
    .B(net773),
    .Y(_01636_));
 sg13g2_nand3_1 _23372_ (.B(_01603_),
    .C(_01636_),
    .A(net268),
    .Y(_01637_));
 sg13g2_xor2_1 _23373_ (.B(net891),
    .A(net1081),
    .X(_01638_));
 sg13g2_nand3_1 _23374_ (.B(net776),
    .C(_09279_),
    .A(_09174_),
    .Y(_01639_));
 sg13g2_o21ai_1 _23375_ (.B1(_01639_),
    .Y(_01640_),
    .A1(net552),
    .A2(_01638_));
 sg13g2_xnor2_1 _23376_ (.Y(_01641_),
    .A(_09279_),
    .B(_01585_));
 sg13g2_nand2_1 _23377_ (.Y(_01642_),
    .A(_01621_),
    .B(_01641_));
 sg13g2_o21ai_1 _23378_ (.B1(_01642_),
    .Y(_01643_),
    .A1(_01621_),
    .A2(_01640_));
 sg13g2_nand3b_1 _23379_ (.B(_01637_),
    .C(_01643_),
    .Y(_01645_),
    .A_N(_13217_));
 sg13g2_o21ai_1 _23380_ (.B1(_01645_),
    .Y(_01646_),
    .A1(_01620_),
    .A2(_01635_));
 sg13g2_a221oi_1 _23381_ (.B2(_01634_),
    .C1(_01646_),
    .B1(_01632_),
    .A1(net204),
    .Y(_01647_),
    .A2(_01626_));
 sg13g2_a21oi_1 _23382_ (.A1(_09174_),
    .A2(net776),
    .Y(_01648_),
    .B1(net550));
 sg13g2_nor4_1 _23383_ (.A(net443),
    .B(net432),
    .C(_09289_),
    .D(_01648_),
    .Y(_01649_));
 sg13g2_a21oi_1 _23384_ (.A1(net443),
    .A2(net773),
    .Y(_01650_),
    .B1(net891));
 sg13g2_o21ai_1 _23385_ (.B1(_09288_),
    .Y(_01651_),
    .A1(_01623_),
    .A2(_01650_));
 sg13g2_o21ai_1 _23386_ (.B1(_01636_),
    .Y(_01652_),
    .A1(net274),
    .A2(_09279_));
 sg13g2_a21oi_1 _23387_ (.A1(_01651_),
    .A2(_01652_),
    .Y(_01653_),
    .B1(net434));
 sg13g2_nor2_1 _23388_ (.A(_01649_),
    .B(_01653_),
    .Y(_01654_));
 sg13g2_nand2_1 _23389_ (.Y(_01656_),
    .A(net83),
    .B(_01654_));
 sg13g2_xnor2_1 _23390_ (.Y(_01657_),
    .A(_01595_),
    .B(_13308_));
 sg13g2_xor2_1 _23391_ (.B(_01657_),
    .A(_01630_),
    .X(_01658_));
 sg13g2_a21oi_1 _23392_ (.A1(net119),
    .A2(_01658_),
    .Y(_01659_),
    .B1(_13190_));
 sg13g2_or2_1 _23393_ (.X(_01660_),
    .B(_13216_),
    .A(_09216_));
 sg13g2_a21o_1 _23394_ (.A2(_01660_),
    .A1(_01630_),
    .B1(_13230_),
    .X(_01661_));
 sg13g2_nand2b_1 _23395_ (.Y(_01662_),
    .B(_13229_),
    .A_N(_13216_));
 sg13g2_nor2b_1 _23396_ (.A(net777),
    .B_N(net784),
    .Y(_01663_));
 sg13g2_a22oi_1 _23397_ (.Y(_01664_),
    .B1(_01663_),
    .B2(_01630_),
    .A2(_01662_),
    .A1(net890));
 sg13g2_a21oi_1 _23398_ (.A1(_01661_),
    .A2(_01664_),
    .Y(_01665_),
    .B1(net1080));
 sg13g2_nand3b_1 _23399_ (.B(_01630_),
    .C(net1080),
    .Y(_01667_),
    .A_N(net784));
 sg13g2_o21ai_1 _23400_ (.B1(_01667_),
    .Y(_01668_),
    .A1(_09217_),
    .A2(_01631_));
 sg13g2_nor4_1 _23401_ (.A(net168),
    .B(_01654_),
    .C(_01665_),
    .D(_01668_),
    .Y(_01669_));
 sg13g2_nor2_1 _23402_ (.A(_01659_),
    .B(_01669_),
    .Y(_01670_));
 sg13g2_o21ai_1 _23403_ (.B1(_01670_),
    .Y(_01671_),
    .A1(_01647_),
    .A2(_01656_));
 sg13g2_nand2_1 _23404_ (.Y(_01672_),
    .A(_12977_),
    .B(net36));
 sg13g2_nor2_2 _23405_ (.A(_08817_),
    .B(_13185_),
    .Y(_01673_));
 sg13g2_nand2_1 _23406_ (.Y(_01674_),
    .A(net1060),
    .B(_01673_));
 sg13g2_nand2b_1 _23407_ (.Y(_01675_),
    .B(net42),
    .A_N(_01674_));
 sg13g2_o21ai_1 _23408_ (.B1(_01675_),
    .Y(_00478_),
    .A1(_01671_),
    .A2(_01672_));
 sg13g2_buf_2 _23409_ (.A(\grid.cell_3_2.se ),
    .X(_01677_));
 sg13g2_xor2_1 _23410_ (.B(_01677_),
    .A(_00613_),
    .X(_01678_));
 sg13g2_buf_1 _23411_ (.A(_01677_),
    .X(_01679_));
 sg13g2_nand2_1 _23412_ (.Y(_01680_),
    .A(_00614_),
    .B(net772));
 sg13g2_a22oi_1 _23413_ (.Y(_01681_),
    .B1(_01680_),
    .B2(_09308_),
    .A2(_01678_),
    .A1(_09238_));
 sg13g2_nor2_1 _23414_ (.A(_00614_),
    .B(net772),
    .Y(_01682_));
 sg13g2_o21ai_1 _23415_ (.B1(_01682_),
    .Y(_01683_),
    .A1(_09279_),
    .A2(_09308_));
 sg13g2_o21ai_1 _23416_ (.B1(_01683_),
    .Y(_01684_),
    .A1(net1124),
    .A2(_01681_));
 sg13g2_buf_1 _23417_ (.A(net772),
    .X(_01685_));
 sg13g2_a21oi_1 _23418_ (.A1(net891),
    .A2(net773),
    .Y(_01686_),
    .B1(net269));
 sg13g2_nor4_1 _23419_ (.A(net1124),
    .B(net441),
    .C(net431),
    .D(_01686_),
    .Y(_01688_));
 sg13g2_a21oi_2 _23420_ (.B1(_01688_),
    .Y(_01689_),
    .A2(_01684_),
    .A1(_01627_));
 sg13g2_nand3_1 _23421_ (.B(net446),
    .C(net781),
    .A(net274),
    .Y(_01690_));
 sg13g2_buf_2 _23422_ (.A(_00267_),
    .X(_01691_));
 sg13g2_inv_2 _23423_ (.Y(_01692_),
    .A(_01691_));
 sg13g2_inv_2 _23424_ (.Y(_01693_),
    .A(net1082));
 sg13g2_nand4_1 _23425_ (.B(net444),
    .C(_01692_),
    .A(_09176_),
    .Y(_01694_),
    .D(_01693_));
 sg13g2_o21ai_1 _23426_ (.B1(_01694_),
    .Y(_01695_),
    .A1(_01689_),
    .A2(_01690_));
 sg13g2_buf_1 _23427_ (.A(_01691_),
    .X(_01696_));
 sg13g2_nand3_1 _23428_ (.B(net771),
    .C(net781),
    .A(net446),
    .Y(_01697_));
 sg13g2_a21oi_1 _23429_ (.A1(_09176_),
    .A2(net771),
    .Y(_01699_),
    .B1(net786));
 sg13g2_o21ai_1 _23430_ (.B1(_01689_),
    .Y(_01700_),
    .A1(_01693_),
    .A2(_01699_));
 sg13g2_o21ai_1 _23431_ (.B1(_01700_),
    .Y(_01701_),
    .A1(_01689_),
    .A2(_01697_));
 sg13g2_xnor2_1 _23432_ (.Y(_01702_),
    .A(net1126),
    .B(_01617_));
 sg13g2_xnor2_1 _23433_ (.Y(_01703_),
    .A(_01677_),
    .B(_00620_));
 sg13g2_xor2_1 _23434_ (.B(_01703_),
    .A(_01702_),
    .X(_01704_));
 sg13g2_inv_1 _23435_ (.Y(_01705_),
    .A(_01704_));
 sg13g2_o21ai_1 _23436_ (.B1(_01705_),
    .Y(_01706_),
    .A1(_01695_),
    .A2(_01701_));
 sg13g2_xnor2_1 _23437_ (.Y(_01707_),
    .A(net444),
    .B(_01585_));
 sg13g2_xnor2_1 _23438_ (.Y(_01708_),
    .A(_01704_),
    .B(_01707_));
 sg13g2_o21ai_1 _23439_ (.B1(_13264_),
    .Y(_01710_),
    .A1(net105),
    .A2(_01708_));
 sg13g2_buf_1 _23440_ (.A(net773),
    .X(_01711_));
 sg13g2_nand2_1 _23441_ (.Y(_01712_),
    .A(_09239_),
    .B(_01678_));
 sg13g2_o21ai_1 _23442_ (.B1(_01712_),
    .Y(_01713_),
    .A1(net268),
    .A2(_01680_));
 sg13g2_nand2_1 _23443_ (.Y(_01714_),
    .A(net549),
    .B(_01713_));
 sg13g2_o21ai_1 _23444_ (.B1(_01714_),
    .Y(_01715_),
    .A1(_00215_),
    .A2(_01680_));
 sg13g2_nor2_1 _23445_ (.A(net444),
    .B(net771),
    .Y(_01716_));
 sg13g2_nor2_1 _23446_ (.A(net550),
    .B(net432),
    .Y(_01717_));
 sg13g2_nand3_1 _23447_ (.B(_01717_),
    .C(_01682_),
    .A(net549),
    .Y(_01718_));
 sg13g2_and4_1 _23448_ (.A(net271),
    .B(_01693_),
    .C(_01716_),
    .D(_01718_),
    .X(_01719_));
 sg13g2_xor2_1 _23449_ (.B(net549),
    .A(net432),
    .X(_01721_));
 sg13g2_nand3_1 _23450_ (.B(net430),
    .C(net269),
    .A(net268),
    .Y(_01722_));
 sg13g2_o21ai_1 _23451_ (.B1(_01722_),
    .Y(_01723_),
    .A1(_09319_),
    .A2(_01721_));
 sg13g2_xnor2_1 _23452_ (.Y(_01724_),
    .A(net269),
    .B(_01702_));
 sg13g2_nand2_1 _23453_ (.Y(_01725_),
    .A(_01678_),
    .B(_01724_));
 sg13g2_o21ai_1 _23454_ (.B1(_01725_),
    .Y(_01726_),
    .A1(_01678_),
    .A2(_01723_));
 sg13g2_buf_1 _23455_ (.A(_01685_),
    .X(_01727_));
 sg13g2_nand2_1 _23456_ (.Y(_01728_),
    .A(net202),
    .B(_01717_));
 sg13g2_o21ai_1 _23457_ (.B1(_01550_),
    .Y(_01729_),
    .A1(_00633_),
    .A2(_01728_));
 sg13g2_a221oi_1 _23458_ (.B2(_01726_),
    .C1(_01729_),
    .B1(_01719_),
    .A1(net430),
    .Y(_01730_),
    .A2(_01715_));
 sg13g2_nand2_1 _23459_ (.Y(_01732_),
    .A(net444),
    .B(net771));
 sg13g2_o21ai_1 _23460_ (.B1(_01732_),
    .Y(_01733_),
    .A1(net552),
    .A2(_01716_));
 sg13g2_nor3_1 _23461_ (.A(_09196_),
    .B(_01692_),
    .C(_01693_),
    .Y(_01734_));
 sg13g2_a21oi_1 _23462_ (.A1(_01704_),
    .A2(_01733_),
    .Y(_01735_),
    .B1(_01734_));
 sg13g2_o21ai_1 _23463_ (.B1(net771),
    .Y(_01736_),
    .A1(net444),
    .A2(_01705_));
 sg13g2_a22oi_1 _23464_ (.Y(_01737_),
    .B1(_01736_),
    .B2(_09197_),
    .A2(_01716_),
    .A1(_01704_));
 sg13g2_mux2_1 _23465_ (.A0(_01735_),
    .A1(_01737_),
    .S(_01689_),
    .X(_01738_));
 sg13g2_nand4_1 _23466_ (.B(_01710_),
    .C(_01730_),
    .A(_01706_),
    .Y(_01739_),
    .D(_01738_));
 sg13g2_o21ai_1 _23467_ (.B1(net36),
    .Y(_01740_),
    .A1(_13264_),
    .A2(net83));
 sg13g2_o21ai_1 _23468_ (.B1(_01740_),
    .Y(_01741_),
    .A1(_05811_),
    .A2(_01550_));
 sg13g2_a21oi_1 _23469_ (.A1(_01739_),
    .A2(_01741_),
    .Y(_00479_),
    .B1(net440));
 sg13g2_buf_2 _23470_ (.A(\grid.cell_3_3.se ),
    .X(_01743_));
 sg13g2_xor2_1 _23471_ (.B(_01743_),
    .A(_00664_),
    .X(_01744_));
 sg13g2_xor2_1 _23472_ (.B(_01744_),
    .A(_09344_),
    .X(_01745_));
 sg13g2_xnor2_1 _23473_ (.Y(_01746_),
    .A(net431),
    .B(_01745_));
 sg13g2_xor2_1 _23474_ (.B(_01746_),
    .A(_01628_),
    .X(_01747_));
 sg13g2_a21oi_1 _23475_ (.A1(net78),
    .A2(_01747_),
    .Y(_01748_),
    .B1(net442));
 sg13g2_inv_1 _23476_ (.Y(_01749_),
    .A(_01743_));
 sg13g2_buf_1 _23477_ (.A(_01749_),
    .X(_01750_));
 sg13g2_xor2_1 _23478_ (.B(net438),
    .A(net431),
    .X(_01751_));
 sg13g2_inv_1 _23479_ (.Y(_01753_),
    .A(net772));
 sg13g2_o21ai_1 _23480_ (.B1(net269),
    .Y(_01754_),
    .A1(_01753_),
    .A2(net439));
 sg13g2_o21ai_1 _23481_ (.B1(_01754_),
    .Y(_01755_),
    .A1(net269),
    .A2(_01751_));
 sg13g2_nand4_1 _23482_ (.B(net202),
    .C(net438),
    .A(net549),
    .Y(_01756_),
    .D(net429));
 sg13g2_o21ai_1 _23483_ (.B1(_01756_),
    .Y(_01757_),
    .A1(net429),
    .A2(_01755_));
 sg13g2_nor2b_1 _23484_ (.A(_00678_),
    .B_N(_01746_),
    .Y(_01758_));
 sg13g2_buf_2 _23485_ (.A(_00266_),
    .X(_01759_));
 sg13g2_nor2_1 _23486_ (.A(_01759_),
    .B(_13304_),
    .Y(_01760_));
 sg13g2_or4_1 _23487_ (.A(_09382_),
    .B(_01753_),
    .C(net439),
    .D(net429),
    .X(_01761_));
 sg13g2_nand3_1 _23488_ (.B(_01549_),
    .C(_01761_),
    .A(net1054),
    .Y(_01762_));
 sg13g2_a221oi_1 _23489_ (.B2(_01760_),
    .C1(_01762_),
    .B1(_01758_),
    .A1(net548),
    .Y(_01764_),
    .A2(_01757_));
 sg13g2_xnor2_1 _23490_ (.Y(_01765_),
    .A(net206),
    .B(_01746_));
 sg13g2_a21oi_1 _23491_ (.A1(_09280_),
    .A2(_01759_),
    .Y(_01766_),
    .B1(_01765_));
 sg13g2_nor2_1 _23492_ (.A(net550),
    .B(_01759_),
    .Y(_01767_));
 sg13g2_nor3_1 _23493_ (.A(_01758_),
    .B(_01766_),
    .C(_01767_),
    .Y(_01768_));
 sg13g2_buf_1 _23494_ (.A(_01743_),
    .X(_01769_));
 sg13g2_buf_1 _23495_ (.A(_01769_),
    .X(_01770_));
 sg13g2_nand2_1 _23496_ (.Y(_01771_),
    .A(net438),
    .B(net428));
 sg13g2_a22oi_1 _23497_ (.Y(_01772_),
    .B1(_01771_),
    .B2(_09336_),
    .A2(_01744_),
    .A1(net549));
 sg13g2_a21oi_1 _23498_ (.A1(_09303_),
    .A2(net431),
    .Y(_01773_),
    .B1(_09336_));
 sg13g2_or3_1 _23499_ (.A(net438),
    .B(net428),
    .C(_01773_),
    .X(_01775_));
 sg13g2_o21ai_1 _23500_ (.B1(_01775_),
    .Y(_01776_),
    .A1(net202),
    .A2(_01772_));
 sg13g2_nor3_1 _23501_ (.A(net202),
    .B(net438),
    .C(net428),
    .Y(_01777_));
 sg13g2_a22oi_1 _23502_ (.Y(_01778_),
    .B1(_01777_),
    .B2(_09335_),
    .A2(_01776_),
    .A1(_09382_));
 sg13g2_xnor2_1 _23503_ (.Y(_01779_),
    .A(_01768_),
    .B(_01778_));
 sg13g2_a22oi_1 _23504_ (.Y(_01780_),
    .B1(_01764_),
    .B2(_01779_),
    .A2(net36),
    .A1(_08877_));
 sg13g2_nand2b_1 _23505_ (.Y(_01781_),
    .B(_01673_),
    .A_N(net26));
 sg13g2_o21ai_1 _23506_ (.B1(_01781_),
    .Y(_00480_),
    .A1(_01748_),
    .A2(_01780_));
 sg13g2_buf_1 _23507_ (.A(\grid.cell_3_4.se ),
    .X(_01782_));
 sg13g2_xor2_1 _23508_ (.B(net1079),
    .A(_00709_),
    .X(_01783_));
 sg13g2_xnor2_1 _23509_ (.Y(_01785_),
    .A(_09387_),
    .B(_01783_));
 sg13g2_xnor2_1 _23510_ (.Y(_01786_),
    .A(net770),
    .B(_01785_));
 sg13g2_nand2_1 _23511_ (.Y(_01787_),
    .A(_00741_),
    .B(_01786_));
 sg13g2_buf_1 _23512_ (.A(_00037_),
    .X(_01788_));
 sg13g2_nand2b_1 _23513_ (.Y(_01789_),
    .B(_00620_),
    .A_N(net1078));
 sg13g2_buf_1 _23514_ (.A(net1079),
    .X(_01790_));
 sg13g2_nand3_1 _23515_ (.B(net779),
    .C(net769),
    .A(net770),
    .Y(_01791_));
 sg13g2_xnor2_1 _23516_ (.Y(_01792_),
    .A(_00709_),
    .B(net1079));
 sg13g2_nor2_1 _23517_ (.A(net429),
    .B(_01792_),
    .Y(_01793_));
 sg13g2_nand2_1 _23518_ (.Y(_01794_),
    .A(net779),
    .B(net769));
 sg13g2_nor2_1 _23519_ (.A(net770),
    .B(_01794_),
    .Y(_01796_));
 sg13g2_o21ai_1 _23520_ (.B1(_09358_),
    .Y(_01797_),
    .A1(_01793_),
    .A2(_01796_));
 sg13g2_o21ai_1 _23521_ (.B1(_01797_),
    .Y(_01798_),
    .A1(net548),
    .A2(_01791_));
 sg13g2_nor2_1 _23522_ (.A(_09419_),
    .B(_01791_),
    .Y(_01799_));
 sg13g2_a21oi_1 _23523_ (.A1(net267),
    .A2(_01798_),
    .Y(_01800_),
    .B1(_01799_));
 sg13g2_o21ai_1 _23524_ (.B1(_01800_),
    .Y(_01801_),
    .A1(_01787_),
    .A2(_01789_));
 sg13g2_nand2_1 _23525_ (.Y(_01802_),
    .A(net1078),
    .B(_09309_));
 sg13g2_xor2_1 _23526_ (.B(_01786_),
    .A(net442),
    .X(_01803_));
 sg13g2_nor2_1 _23527_ (.A(net1078),
    .B(_09309_),
    .Y(_01804_));
 sg13g2_a221oi_1 _23528_ (.B2(_01803_),
    .C1(_01804_),
    .B1(_01802_),
    .A1(_00741_),
    .Y(_01805_),
    .A2(_01786_));
 sg13g2_a22oi_1 _23529_ (.Y(_01807_),
    .B1(_01783_),
    .B2(_09339_),
    .A2(_01794_),
    .A1(_09413_));
 sg13g2_inv_2 _23530_ (.Y(_01808_),
    .A(_01782_));
 sg13g2_o21ai_1 _23531_ (.B1(net887),
    .Y(_01809_),
    .A1(_09336_),
    .A2(net429));
 sg13g2_nand3_1 _23532_ (.B(_01808_),
    .C(_01809_),
    .A(_00718_),
    .Y(_01810_));
 sg13g2_o21ai_1 _23533_ (.B1(_01810_),
    .Y(_01811_),
    .A1(net428),
    .A2(_01807_));
 sg13g2_buf_1 _23534_ (.A(net769),
    .X(_01812_));
 sg13g2_nor3_1 _23535_ (.A(net428),
    .B(net437),
    .C(net427),
    .Y(_01813_));
 sg13g2_a22oi_1 _23536_ (.Y(_01814_),
    .B1(_01813_),
    .B2(_09372_),
    .A2(_01811_),
    .A1(_09419_));
 sg13g2_xor2_1 _23537_ (.B(_01814_),
    .A(_01805_),
    .X(_01815_));
 sg13g2_o21ai_1 _23538_ (.B1(net83),
    .Y(_01816_),
    .A1(_01801_),
    .A2(_01815_));
 sg13g2_xnor2_1 _23539_ (.Y(_01818_),
    .A(_01703_),
    .B(_01786_));
 sg13g2_o21ai_1 _23540_ (.B1(net439),
    .Y(_01819_),
    .A1(_04624_),
    .A2(_01818_));
 sg13g2_nand4_1 _23541_ (.B(net36),
    .C(_01816_),
    .A(_05355_),
    .Y(_01820_),
    .D(_01819_));
 sg13g2_o21ai_1 _23542_ (.B1(_01820_),
    .Y(_00481_),
    .A1(net29),
    .A2(_01674_));
 sg13g2_buf_2 _23543_ (.A(\grid.cell_3_5.se ),
    .X(_01821_));
 sg13g2_buf_1 _23544_ (.A(_01821_),
    .X(_01822_));
 sg13g2_nand2_1 _23545_ (.Y(_01823_),
    .A(_00753_),
    .B(net768));
 sg13g2_xor2_1 _23546_ (.B(_01821_),
    .A(_00752_),
    .X(_01824_));
 sg13g2_buf_2 _23547_ (.A(_01824_),
    .X(_01825_));
 sg13g2_nand2_1 _23548_ (.Y(_01826_),
    .A(net427),
    .B(_01825_));
 sg13g2_o21ai_1 _23549_ (.B1(_01826_),
    .Y(_01828_),
    .A1(net427),
    .A2(_01823_));
 sg13g2_buf_1 _23550_ (.A(_01822_),
    .X(_01829_));
 sg13g2_nand3_1 _23551_ (.B(net205),
    .C(net426),
    .A(net769),
    .Y(_01830_));
 sg13g2_nor2_1 _23552_ (.A(net267),
    .B(_01830_),
    .Y(_01831_));
 sg13g2_a21oi_1 _23553_ (.A1(_09381_),
    .A2(_01828_),
    .Y(_01832_),
    .B1(_01831_));
 sg13g2_nand2b_1 _23554_ (.Y(_01833_),
    .B(_09461_),
    .A_N(_01830_));
 sg13g2_o21ai_1 _23555_ (.B1(_01833_),
    .Y(_01834_),
    .A1(_09412_),
    .A2(_01832_));
 sg13g2_o21ai_1 _23556_ (.B1(_00763_),
    .Y(_01835_),
    .A1(_09336_),
    .A2(_00665_));
 sg13g2_nor2_1 _23557_ (.A(_09336_),
    .B(net439),
    .Y(_01836_));
 sg13g2_xnor2_1 _23558_ (.Y(_01837_),
    .A(_09407_),
    .B(net1079));
 sg13g2_xnor2_1 _23559_ (.Y(_01839_),
    .A(_01825_),
    .B(_01837_));
 sg13g2_xnor2_1 _23560_ (.Y(_01840_),
    .A(net887),
    .B(_01839_));
 sg13g2_mux2_1 _23561_ (.A0(_01835_),
    .A1(_01836_),
    .S(_01840_),
    .X(_01841_));
 sg13g2_a22oi_1 _23562_ (.Y(_01842_),
    .B1(_01825_),
    .B2(_09371_),
    .A2(_01823_),
    .A1(_09411_));
 sg13g2_nand2_1 _23563_ (.Y(_01843_),
    .A(_09371_),
    .B(net1079));
 sg13g2_or2_1 _23564_ (.X(_01844_),
    .B(net768),
    .A(_00753_));
 sg13g2_a21o_1 _23565_ (.A2(_01843_),
    .A1(_09407_),
    .B1(_01844_),
    .X(_01845_));
 sg13g2_o21ai_1 _23566_ (.B1(_01845_),
    .Y(_01846_),
    .A1(net769),
    .A2(_01842_));
 sg13g2_a21oi_1 _23567_ (.A1(_09408_),
    .A2(net547),
    .Y(_01847_),
    .B1(_01844_));
 sg13g2_a22oi_1 _23568_ (.Y(_01848_),
    .B1(_01847_),
    .B2(_01808_),
    .A2(_01846_),
    .A1(_00099_));
 sg13g2_or2_1 _23569_ (.X(_01850_),
    .B(_01848_),
    .A(_01841_));
 sg13g2_xnor2_1 _23570_ (.Y(_01851_),
    .A(_01841_),
    .B(_01848_));
 sg13g2_buf_1 _23571_ (.A(_00069_),
    .X(_01852_));
 sg13g2_inv_1 _23572_ (.Y(_01853_),
    .A(_01852_));
 sg13g2_xnor2_1 _23573_ (.Y(_01854_),
    .A(_09387_),
    .B(_01839_));
 sg13g2_xnor2_1 _23574_ (.Y(_01855_),
    .A(net438),
    .B(_01854_));
 sg13g2_nand2_1 _23575_ (.Y(_01856_),
    .A(_01853_),
    .B(_01855_));
 sg13g2_mux2_1 _23576_ (.A0(_01850_),
    .A1(_01851_),
    .S(_01856_),
    .X(_01857_));
 sg13g2_o21ai_1 _23577_ (.B1(net82),
    .Y(_01858_),
    .A1(_01834_),
    .A2(_01857_));
 sg13g2_xnor2_1 _23578_ (.Y(_01859_),
    .A(_01744_),
    .B(_01854_));
 sg13g2_a21oi_1 _23579_ (.A1(net98),
    .A2(_01859_),
    .Y(_01861_),
    .B1(net437));
 sg13g2_nor2_1 _23580_ (.A(_01673_),
    .B(_01861_),
    .Y(_01862_));
 sg13g2_a22oi_1 _23581_ (.Y(_01863_),
    .B1(_01858_),
    .B2(_01862_),
    .A2(_01673_),
    .A1(_06330_));
 sg13g2_nor2_1 _23582_ (.A(net214),
    .B(_01863_),
    .Y(_00482_));
 sg13g2_nand2_1 _23583_ (.Y(_01864_),
    .A(net426),
    .B(_01562_));
 sg13g2_buf_1 _23584_ (.A(_01829_),
    .X(_01865_));
 sg13g2_nor2_1 _23585_ (.A(net768),
    .B(_01562_),
    .Y(_01866_));
 sg13g2_a21oi_1 _23586_ (.A1(net201),
    .A2(_01605_),
    .Y(_01867_),
    .B1(_01866_));
 sg13g2_nand2_1 _23587_ (.Y(_01868_),
    .A(_09471_),
    .B(_01867_));
 sg13g2_o21ai_1 _23588_ (.B1(_01868_),
    .Y(_01869_),
    .A1(_09471_),
    .A2(_01864_));
 sg13g2_xnor2_1 _23589_ (.Y(_01871_),
    .A(_01555_),
    .B(_09462_));
 sg13g2_xor2_1 _23590_ (.B(net785),
    .A(net768),
    .X(_01872_));
 sg13g2_xnor2_1 _23591_ (.Y(_01873_),
    .A(_01871_),
    .B(_01872_));
 sg13g2_nor2_1 _23592_ (.A(_00827_),
    .B(_01873_),
    .Y(_01874_));
 sg13g2_buf_2 _23593_ (.A(_00101_),
    .X(_01875_));
 sg13g2_xor2_1 _23594_ (.B(_00736_),
    .A(net267),
    .X(_01876_));
 sg13g2_nor2_1 _23595_ (.A(_01875_),
    .B(_01876_),
    .Y(_01877_));
 sg13g2_buf_1 _23596_ (.A(_00131_),
    .X(_01878_));
 sg13g2_nor2_1 _23597_ (.A(net1077),
    .B(_01864_),
    .Y(_01879_));
 sg13g2_a221oi_1 _23598_ (.B2(_01877_),
    .C1(_01879_),
    .B1(_01874_),
    .A1(net270),
    .Y(_01880_),
    .A2(_01869_));
 sg13g2_nand2_1 _23599_ (.Y(_01882_),
    .A(net546),
    .B(net270));
 sg13g2_xor2_1 _23600_ (.B(net426),
    .A(net1077),
    .X(_01883_));
 sg13g2_nand3_1 _23601_ (.B(net426),
    .C(_01570_),
    .A(net1077),
    .Y(_01884_));
 sg13g2_o21ai_1 _23602_ (.B1(_01884_),
    .Y(_01885_),
    .A1(net1077),
    .A2(_01570_));
 sg13g2_a21oi_1 _23603_ (.A1(_01560_),
    .A2(_01883_),
    .Y(_01886_),
    .B1(_01885_));
 sg13g2_inv_2 _23604_ (.Y(_01887_),
    .A(_01821_));
 sg13g2_nand2_1 _23605_ (.Y(_01888_),
    .A(_01887_),
    .B(_01559_));
 sg13g2_o21ai_1 _23606_ (.B1(_01888_),
    .Y(_01889_),
    .A1(net272),
    .A2(_01864_));
 sg13g2_o21ai_1 _23607_ (.B1(_00131_),
    .Y(_01890_),
    .A1(_01559_),
    .A2(_01866_));
 sg13g2_nand2_1 _23608_ (.Y(_01891_),
    .A(_01888_),
    .B(_01890_));
 sg13g2_a221oi_1 _23609_ (.B2(net272),
    .C1(_01879_),
    .B1(_01891_),
    .A1(_09412_),
    .Y(_01893_),
    .A2(_01889_));
 sg13g2_o21ai_1 _23610_ (.B1(_01893_),
    .Y(_01894_),
    .A1(_01882_),
    .A2(_01886_));
 sg13g2_xnor2_1 _23611_ (.Y(_01895_),
    .A(_00718_),
    .B(_01873_));
 sg13g2_a21oi_1 _23612_ (.A1(_01875_),
    .A2(_09413_),
    .Y(_01896_),
    .B1(_01895_));
 sg13g2_nor2_1 _23613_ (.A(_01875_),
    .B(_09413_),
    .Y(_01897_));
 sg13g2_nor3_1 _23614_ (.A(_01874_),
    .B(_01896_),
    .C(_01897_),
    .Y(_01898_));
 sg13g2_xor2_1 _23615_ (.B(_01898_),
    .A(_01894_),
    .X(_01899_));
 sg13g2_a21oi_1 _23616_ (.A1(_01880_),
    .A2(_01899_),
    .Y(_01900_),
    .B1(_05737_));
 sg13g2_xnor2_1 _23617_ (.Y(_01901_),
    .A(_09413_),
    .B(_01792_));
 sg13g2_xnor2_1 _23618_ (.Y(_01902_),
    .A(_01873_),
    .B(_01901_));
 sg13g2_o21ai_1 _23619_ (.B1(_00771_),
    .Y(_01904_),
    .A1(_06466_),
    .A2(_01902_));
 sg13g2_nand2b_1 _23620_ (.Y(_01905_),
    .B(_01904_),
    .A_N(_01672_));
 sg13g2_nand2b_1 _23621_ (.Y(_01906_),
    .B(net31),
    .A_N(_01674_));
 sg13g2_o21ai_1 _23622_ (.B1(_01906_),
    .Y(_00483_),
    .A1(_01900_),
    .A2(_01905_));
 sg13g2_xnor2_1 _23623_ (.Y(_01907_),
    .A(_01825_),
    .B(_01871_));
 sg13g2_xnor2_1 _23624_ (.Y(_01908_),
    .A(net777),
    .B(_01907_));
 sg13g2_nand2_1 _23625_ (.Y(_01909_),
    .A(_01583_),
    .B(_01908_));
 sg13g2_nor2_1 _23626_ (.A(_13217_),
    .B(_01907_),
    .Y(_01910_));
 sg13g2_a21oi_1 _23627_ (.A1(net890),
    .A2(_01589_),
    .Y(_01911_),
    .B1(_01910_));
 sg13g2_nand2_1 _23628_ (.Y(_01912_),
    .A(_01909_),
    .B(_01911_));
 sg13g2_nand2_2 _23629_ (.Y(_01914_),
    .A(net768),
    .B(net775));
 sg13g2_nand3_1 _23630_ (.B(net436),
    .C(_01914_),
    .A(_01878_),
    .Y(_01915_));
 sg13g2_o21ai_1 _23631_ (.B1(_01915_),
    .Y(_01916_),
    .A1(net1077),
    .A2(_01914_));
 sg13g2_inv_1 _23632_ (.Y(_01917_),
    .A(_01916_));
 sg13g2_nor2_1 _23633_ (.A(net426),
    .B(net433),
    .Y(_01918_));
 sg13g2_xor2_1 _23634_ (.B(net205),
    .A(net1077),
    .X(_01919_));
 sg13g2_nand2b_1 _23635_ (.Y(_01920_),
    .B(_01919_),
    .A_N(_01918_));
 sg13g2_a21oi_1 _23636_ (.A1(_01917_),
    .A2(_01920_),
    .Y(_01921_),
    .B1(_01882_));
 sg13g2_nand3_1 _23637_ (.B(net426),
    .C(net775),
    .A(net436),
    .Y(_01922_));
 sg13g2_buf_1 _23638_ (.A(_01922_),
    .X(_01923_));
 sg13g2_nand2_1 _23639_ (.Y(_01925_),
    .A(_00771_),
    .B(_01918_));
 sg13g2_o21ai_1 _23640_ (.B1(_01925_),
    .Y(_01926_),
    .A1(_09191_),
    .A2(_01923_));
 sg13g2_and2_1 _23641_ (.A(net545),
    .B(_01926_),
    .X(_01927_));
 sg13g2_nor2_1 _23642_ (.A(net1077),
    .B(_01923_),
    .Y(_01928_));
 sg13g2_a21oi_1 _23643_ (.A1(net201),
    .A2(net203),
    .Y(_01929_),
    .B1(net205));
 sg13g2_o21ai_1 _23644_ (.B1(net1077),
    .Y(_01930_),
    .A1(_01918_),
    .A2(_01929_));
 sg13g2_a21oi_1 _23645_ (.A1(_01925_),
    .A2(_01930_),
    .Y(_01931_),
    .B1(_09201_));
 sg13g2_nor4_1 _23646_ (.A(_01921_),
    .B(_01927_),
    .C(_01928_),
    .D(_01931_),
    .Y(_01932_));
 sg13g2_xnor2_1 _23647_ (.Y(_01933_),
    .A(_01912_),
    .B(_01932_));
 sg13g2_xnor2_1 _23648_ (.Y(_01934_),
    .A(_01657_),
    .B(_01907_));
 sg13g2_and2_1 _23649_ (.A(_01589_),
    .B(_13308_),
    .X(_01936_));
 sg13g2_and2_1 _23650_ (.A(net433),
    .B(_01825_),
    .X(_01937_));
 sg13g2_nor2_1 _23651_ (.A(net433),
    .B(_01823_),
    .Y(_01938_));
 sg13g2_o21ai_1 _23652_ (.B1(_09409_),
    .Y(_01939_),
    .A1(_01937_),
    .A2(_01938_));
 sg13g2_o21ai_1 _23653_ (.B1(_01939_),
    .Y(_01940_),
    .A1(_09409_),
    .A2(_01923_));
 sg13g2_nand2_1 _23654_ (.Y(_01941_),
    .A(net270),
    .B(_01940_));
 sg13g2_nor3_1 _23655_ (.A(_00648_),
    .B(net170),
    .C(_01928_),
    .Y(_01942_));
 sg13g2_nand2_1 _23656_ (.Y(_01943_),
    .A(_01941_),
    .B(_01942_));
 sg13g2_a221oi_1 _23657_ (.B2(_01936_),
    .C1(_01943_),
    .B1(_01910_),
    .A1(_05748_),
    .Y(_01944_),
    .A2(_00839_));
 sg13g2_o21ai_1 _23658_ (.B1(_01944_),
    .Y(_01945_),
    .A1(net207),
    .A2(_01934_));
 sg13g2_nand3_1 _23659_ (.B(net110),
    .C(net36),
    .A(net207),
    .Y(_01947_));
 sg13g2_o21ai_1 _23660_ (.B1(_01947_),
    .Y(_01948_),
    .A1(_05129_),
    .A2(net36));
 sg13g2_nand2_1 _23661_ (.Y(_01949_),
    .A(net356),
    .B(_01948_));
 sg13g2_o21ai_1 _23662_ (.B1(_01949_),
    .Y(_00484_),
    .A1(_01933_),
    .A2(_01945_));
 sg13g2_nor2_1 _23663_ (.A(_01989_),
    .B(_09520_),
    .Y(_01950_));
 sg13g2_nand2_2 _23664_ (.Y(_01951_),
    .A(_06113_),
    .B(_01950_));
 sg13g2_buf_1 _23665_ (.A(\grid.cell_4_0.se ),
    .X(_01952_));
 sg13g2_buf_1 _23666_ (.A(net1076),
    .X(_01953_));
 sg13g2_buf_1 _23667_ (.A(net767),
    .X(_01954_));
 sg13g2_buf_2 _23668_ (.A(\grid.cell_4_0.sw ),
    .X(_01955_));
 sg13g2_buf_1 _23669_ (.A(_01955_),
    .X(_01957_));
 sg13g2_buf_1 _23670_ (.A(net766),
    .X(_01958_));
 sg13g2_buf_1 _23671_ (.A(net424),
    .X(_01959_));
 sg13g2_buf_1 _23672_ (.A(net200),
    .X(_01960_));
 sg13g2_nand2_1 _23673_ (.Y(_01961_),
    .A(net424),
    .B(_01693_));
 sg13g2_o21ai_1 _23674_ (.B1(_01961_),
    .Y(_01962_),
    .A1(net134),
    .A2(_13209_));
 sg13g2_nor2_1 _23675_ (.A(net134),
    .B(net1082),
    .Y(_01963_));
 sg13g2_nor3_1 _23676_ (.A(net203),
    .B(_13209_),
    .C(_01963_),
    .Y(_01964_));
 sg13g2_a21o_1 _23677_ (.A2(_01962_),
    .A1(net203),
    .B1(_01964_),
    .X(_01965_));
 sg13g2_nor2_1 _23678_ (.A(net200),
    .B(_01693_),
    .Y(_01966_));
 sg13g2_a21o_1 _23679_ (.A2(_01961_),
    .A1(_01584_),
    .B1(_01966_),
    .X(_01968_));
 sg13g2_nand2_1 _23680_ (.Y(_01969_),
    .A(net200),
    .B(net1082));
 sg13g2_o21ai_1 _23681_ (.B1(net433),
    .Y(_01970_),
    .A1(net200),
    .A2(net1082));
 sg13g2_a21oi_1 _23682_ (.A1(_01969_),
    .A2(_01970_),
    .Y(_01971_),
    .B1(_13209_));
 sg13g2_a21oi_1 _23683_ (.A1(_13194_),
    .A2(_01968_),
    .Y(_01972_),
    .B1(_01971_));
 sg13g2_inv_1 _23684_ (.Y(_01973_),
    .A(net1076));
 sg13g2_nor2_1 _23685_ (.A(net775),
    .B(net424),
    .Y(_01974_));
 sg13g2_nand2_1 _23686_ (.Y(_01975_),
    .A(_01973_),
    .B(_01974_));
 sg13g2_and2_1 _23687_ (.A(_01555_),
    .B(net766),
    .X(_01976_));
 sg13g2_buf_1 _23688_ (.A(_01976_),
    .X(_01977_));
 sg13g2_nand3_1 _23689_ (.B(net445),
    .C(_01977_),
    .A(net767),
    .Y(_01979_));
 sg13g2_a21oi_1 _23690_ (.A1(_01975_),
    .A2(_01979_),
    .Y(_01980_),
    .B1(net786));
 sg13g2_a21oi_1 _23691_ (.A1(_01559_),
    .A2(_01966_),
    .Y(_01981_),
    .B1(_01980_));
 sg13g2_o21ai_1 _23692_ (.B1(_01981_),
    .Y(_01982_),
    .A1(net425),
    .A2(_01972_));
 sg13g2_a21oi_1 _23693_ (.A1(net425),
    .A2(_01965_),
    .Y(_01983_),
    .B1(_01982_));
 sg13g2_xnor2_1 _23694_ (.Y(_01984_),
    .A(_13188_),
    .B(net1076));
 sg13g2_xnor2_1 _23695_ (.Y(_01985_),
    .A(_01605_),
    .B(_01984_));
 sg13g2_xnor2_1 _23696_ (.Y(_01986_),
    .A(net424),
    .B(_01985_));
 sg13g2_xor2_1 _23697_ (.B(_01986_),
    .A(_01553_),
    .X(_01987_));
 sg13g2_buf_1 _23698_ (.A(_00265_),
    .X(_01988_));
 sg13g2_nand2_1 _23699_ (.Y(_01990_),
    .A(_13230_),
    .B(_01988_));
 sg13g2_buf_1 _23700_ (.A(_01988_),
    .X(_01991_));
 sg13g2_nor2_1 _23701_ (.A(_13230_),
    .B(net765),
    .Y(_01992_));
 sg13g2_a221oi_1 _23702_ (.B2(_01990_),
    .C1(_01992_),
    .B1(_01987_),
    .A1(_01692_),
    .Y(_01993_),
    .A2(_01986_));
 sg13g2_xnor2_1 _23703_ (.Y(_01994_),
    .A(_01983_),
    .B(_01993_));
 sg13g2_buf_2 _23704_ (.A(\grid.cell_4_0.s ),
    .X(_01995_));
 sg13g2_xor2_1 _23705_ (.B(_01995_),
    .A(_13229_),
    .X(_01996_));
 sg13g2_xor2_1 _23706_ (.B(_01996_),
    .A(_01987_),
    .X(_01997_));
 sg13g2_nor2_1 _23707_ (.A(net774),
    .B(_01997_),
    .Y(_01998_));
 sg13g2_nand2_1 _23708_ (.Y(_01999_),
    .A(_01692_),
    .B(_01986_));
 sg13g2_xor2_1 _23709_ (.B(net204),
    .A(net777),
    .X(_02001_));
 sg13g2_nor3_1 _23710_ (.A(net765),
    .B(_01999_),
    .C(_02001_),
    .Y(_02002_));
 sg13g2_inv_1 _23711_ (.Y(_02003_),
    .A(net766));
 sg13g2_nor2_1 _23712_ (.A(_02003_),
    .B(net781),
    .Y(_02004_));
 sg13g2_nand2_1 _23713_ (.Y(_02005_),
    .A(net775),
    .B(net766));
 sg13g2_buf_2 _23714_ (.A(_02005_),
    .X(_02006_));
 sg13g2_xor2_1 _23715_ (.B(_01955_),
    .A(_01555_),
    .X(_02007_));
 sg13g2_nand2_1 _23716_ (.Y(_02008_),
    .A(net786),
    .B(_02007_));
 sg13g2_o21ai_1 _23717_ (.B1(_02008_),
    .Y(_02009_),
    .A1(net786),
    .A2(_02006_));
 sg13g2_buf_1 _23718_ (.A(_01973_),
    .X(_02010_));
 sg13g2_a221oi_1 _23719_ (.B2(net207),
    .C1(net423),
    .B1(_02009_),
    .A1(net203),
    .Y(_02012_),
    .A2(_02004_));
 sg13g2_o21ai_1 _23720_ (.B1(net423),
    .Y(_02013_),
    .A1(_13209_),
    .A2(_02006_));
 sg13g2_nor2b_1 _23721_ (.A(_02012_),
    .B_N(_02013_),
    .Y(_02014_));
 sg13g2_nor4_1 _23722_ (.A(net106),
    .B(_01998_),
    .C(_02002_),
    .D(_02014_),
    .Y(_02015_));
 sg13g2_a22oi_1 _23723_ (.Y(_02016_),
    .B1(_01994_),
    .B2(_02015_),
    .A2(_11411_),
    .A1(net774));
 sg13g2_o21ai_1 _23724_ (.B1(_00977_),
    .Y(_02017_),
    .A1(_09235_),
    .A2(_01951_));
 sg13g2_a21oi_1 _23725_ (.A1(_01951_),
    .A2(_02016_),
    .Y(_00485_),
    .B1(_02017_));
 sg13g2_inv_1 _23726_ (.Y(_02018_),
    .A(_01595_));
 sg13g2_o21ai_1 _23727_ (.B1(net777),
    .Y(_02019_),
    .A1(net764),
    .A2(_01582_));
 sg13g2_nor2_1 _23728_ (.A(_13229_),
    .B(_00268_),
    .Y(_02020_));
 sg13g2_buf_2 _23729_ (.A(\grid.cell_4_1.se ),
    .X(_02022_));
 sg13g2_inv_1 _23730_ (.Y(_02023_),
    .A(_02022_));
 sg13g2_xnor2_1 _23731_ (.Y(_02024_),
    .A(net763),
    .B(_01621_));
 sg13g2_xnor2_1 _23732_ (.Y(_02025_),
    .A(_01984_),
    .B(_02024_));
 sg13g2_nand2b_1 _23733_ (.Y(_02026_),
    .B(_02025_),
    .A_N(_02020_));
 sg13g2_nor2_1 _23734_ (.A(net774),
    .B(_01589_),
    .Y(_02027_));
 sg13g2_a22oi_1 _23735_ (.Y(_02028_),
    .B1(_02027_),
    .B2(_02025_),
    .A2(_02026_),
    .A1(net774));
 sg13g2_a21oi_1 _23736_ (.A1(_02019_),
    .A2(_02028_),
    .Y(_02029_),
    .B1(net765));
 sg13g2_xnor2_1 _23737_ (.Y(_02030_),
    .A(_01595_),
    .B(_02025_));
 sg13g2_nand3_1 _23738_ (.B(_01589_),
    .C(_02025_),
    .A(_01988_),
    .Y(_02031_));
 sg13g2_o21ai_1 _23739_ (.B1(_02031_),
    .Y(_02033_),
    .A1(_13230_),
    .A2(_02030_));
 sg13g2_or2_1 _23740_ (.X(_02034_),
    .B(_02033_),
    .A(_02029_));
 sg13g2_buf_1 _23741_ (.A(_02022_),
    .X(_02035_));
 sg13g2_nor2_1 _23742_ (.A(net773),
    .B(net762),
    .Y(_02036_));
 sg13g2_xor2_1 _23743_ (.B(_02022_),
    .A(_01617_),
    .X(_02037_));
 sg13g2_buf_1 _23744_ (.A(net762),
    .X(_02038_));
 sg13g2_a21oi_1 _23745_ (.A1(_01619_),
    .A2(net422),
    .Y(_02039_),
    .B1(net443));
 sg13g2_a21o_1 _23746_ (.A2(_02037_),
    .A1(_13189_),
    .B1(_02039_),
    .X(_02040_));
 sg13g2_a22oi_1 _23747_ (.Y(_02041_),
    .B1(_02040_),
    .B2(_00626_),
    .A2(_02036_),
    .A1(_13276_));
 sg13g2_o21ai_1 _23748_ (.B1(net206),
    .Y(_02042_),
    .A1(_13238_),
    .A2(net423));
 sg13g2_nand3_1 _23749_ (.B(_02042_),
    .C(_02036_),
    .A(_00626_),
    .Y(_02044_));
 sg13g2_o21ai_1 _23750_ (.B1(_02044_),
    .Y(_02045_),
    .A1(net425),
    .A2(_02041_));
 sg13g2_nand2_1 _23751_ (.Y(_02046_),
    .A(net762),
    .B(_01693_));
 sg13g2_o21ai_1 _23752_ (.B1(_02046_),
    .Y(_02047_),
    .A1(net422),
    .A2(_13276_));
 sg13g2_nor2_1 _23753_ (.A(net762),
    .B(net1082),
    .Y(_02048_));
 sg13g2_nor3_1 _23754_ (.A(_01619_),
    .B(_13276_),
    .C(_02048_),
    .Y(_02049_));
 sg13g2_a21oi_1 _23755_ (.A1(net430),
    .A2(_02047_),
    .Y(_02050_),
    .B1(_02049_));
 sg13g2_nand2_1 _23756_ (.Y(_02051_),
    .A(net763),
    .B(_00619_));
 sg13g2_nand2_1 _23757_ (.Y(_02052_),
    .A(_01627_),
    .B(_02046_));
 sg13g2_a21oi_1 _23758_ (.A1(_02051_),
    .A2(_02052_),
    .Y(_02053_),
    .B1(_13299_));
 sg13g2_nor2_1 _23759_ (.A(_01627_),
    .B(_02048_),
    .Y(_02055_));
 sg13g2_a21oi_1 _23760_ (.A1(net422),
    .A2(net1082),
    .Y(_02056_),
    .B1(_02055_));
 sg13g2_nor2_1 _23761_ (.A(_13276_),
    .B(_02056_),
    .Y(_02057_));
 sg13g2_nor3_1 _23762_ (.A(net767),
    .B(_02053_),
    .C(_02057_),
    .Y(_02058_));
 sg13g2_a21oi_1 _23763_ (.A1(net425),
    .A2(_02050_),
    .Y(_02059_),
    .B1(_02058_));
 sg13g2_nand2_1 _23764_ (.Y(_02060_),
    .A(_01973_),
    .B(_02036_));
 sg13g2_nor2_1 _23765_ (.A(_13276_),
    .B(_02060_),
    .Y(_02061_));
 sg13g2_xnor2_1 _23766_ (.Y(_02062_),
    .A(net1076),
    .B(net783));
 sg13g2_nand2_1 _23767_ (.Y(_02063_),
    .A(_13237_),
    .B(_02062_));
 sg13g2_nand2b_1 _23768_ (.Y(_02064_),
    .B(net786),
    .A_N(_02062_));
 sg13g2_and3_1 _23769_ (.X(_02066_),
    .A(_02037_),
    .B(_02063_),
    .C(_02064_));
 sg13g2_nand3_1 _23770_ (.B(net767),
    .C(_13264_),
    .A(net786),
    .Y(_02067_));
 sg13g2_a21oi_1 _23771_ (.A1(_02063_),
    .A2(_02067_),
    .Y(_02068_),
    .B1(_02037_));
 sg13g2_nor4_1 _23772_ (.A(net1080),
    .B(_02061_),
    .C(_02066_),
    .D(_02068_),
    .Y(_02069_));
 sg13g2_buf_1 _23773_ (.A(net762),
    .X(_02070_));
 sg13g2_nand4_1 _23774_ (.B(net206),
    .C(net430),
    .A(net767),
    .Y(_02071_),
    .D(net421));
 sg13g2_a21oi_1 _23775_ (.A1(_02060_),
    .A2(_02071_),
    .Y(_02072_),
    .B1(net446));
 sg13g2_nor3_1 _23776_ (.A(_13299_),
    .B(net430),
    .C(_02051_),
    .Y(_02073_));
 sg13g2_nor4_1 _23777_ (.A(_02059_),
    .B(_02069_),
    .C(_02072_),
    .D(_02073_),
    .Y(_02074_));
 sg13g2_o21ai_1 _23778_ (.B1(_13230_),
    .Y(_02075_),
    .A1(net765),
    .A2(_02030_));
 sg13g2_nand2_1 _23779_ (.Y(_02077_),
    .A(net765),
    .B(_02030_));
 sg13g2_nand2_1 _23780_ (.Y(_02078_),
    .A(_02075_),
    .B(_02077_));
 sg13g2_a221oi_1 _23781_ (.B2(_02078_),
    .C1(_08737_),
    .B1(_02074_),
    .A1(_02034_),
    .Y(_02079_),
    .A2(_02045_));
 sg13g2_xnor2_1 _23782_ (.Y(_02080_),
    .A(_01996_),
    .B(_02030_));
 sg13g2_a21oi_1 _23783_ (.A1(_05739_),
    .A2(_02080_),
    .Y(_02081_),
    .B1(net204));
 sg13g2_nand2_1 _23784_ (.Y(_02082_),
    .A(_13074_),
    .B(_01951_));
 sg13g2_or2_1 _23785_ (.X(_02083_),
    .B(_02082_),
    .A(_02081_));
 sg13g2_nor3_1 _23786_ (.A(_01989_),
    .B(net375),
    .C(_09520_),
    .Y(_02084_));
 sg13g2_buf_2 _23787_ (.A(_02084_),
    .X(_02085_));
 sg13g2_nand2_1 _23788_ (.Y(_02086_),
    .A(net1002),
    .B(_02085_));
 sg13g2_nand2b_1 _23789_ (.Y(_02088_),
    .B(_07276_),
    .A_N(_02086_));
 sg13g2_o21ai_1 _23790_ (.B1(_02088_),
    .Y(_00486_),
    .A1(_02079_),
    .A2(_02083_));
 sg13g2_nand2_1 _23791_ (.Y(_02089_),
    .A(_05812_),
    .B(_02085_));
 sg13g2_xnor2_1 _23792_ (.Y(_02090_),
    .A(_13252_),
    .B(_02022_));
 sg13g2_buf_1 _23793_ (.A(\grid.cell_4_2.se ),
    .X(_02091_));
 sg13g2_buf_1 _23794_ (.A(_02091_),
    .X(_02092_));
 sg13g2_xor2_1 _23795_ (.B(_01678_),
    .A(net761),
    .X(_02093_));
 sg13g2_xnor2_1 _23796_ (.Y(_02094_),
    .A(_02090_),
    .B(_02093_));
 sg13g2_nand2_1 _23797_ (.Y(_02095_),
    .A(_01692_),
    .B(_02094_));
 sg13g2_nand2_1 _23798_ (.Y(_02096_),
    .A(net772),
    .B(net761));
 sg13g2_xnor2_1 _23799_ (.Y(_02098_),
    .A(_01677_),
    .B(_02091_));
 sg13g2_nor2b_1 _23800_ (.A(_02098_),
    .B_N(net783),
    .Y(_02099_));
 sg13g2_nor2_1 _23801_ (.A(net443),
    .B(_02096_),
    .Y(_02100_));
 sg13g2_o21ai_1 _23802_ (.B1(_00644_),
    .Y(_02101_),
    .A1(_02099_),
    .A2(_02100_));
 sg13g2_o21ai_1 _23803_ (.B1(_02101_),
    .Y(_02102_),
    .A1(_00678_),
    .A2(_02096_));
 sg13g2_nand2_1 _23804_ (.Y(_02103_),
    .A(_13298_),
    .B(net441));
 sg13g2_nor2_1 _23805_ (.A(net421),
    .B(_02103_),
    .Y(_02104_));
 sg13g2_and2_1 _23806_ (.A(net772),
    .B(net761),
    .X(_02105_));
 sg13g2_a22oi_1 _23807_ (.Y(_02106_),
    .B1(_02104_),
    .B2(_02105_),
    .A2(_02102_),
    .A1(net421));
 sg13g2_buf_1 _23808_ (.A(_00264_),
    .X(_02107_));
 sg13g2_buf_1 _23809_ (.A(net1075),
    .X(_02109_));
 sg13g2_xnor2_1 _23810_ (.Y(_02110_),
    .A(net1081),
    .B(_00613_));
 sg13g2_xnor2_1 _23811_ (.Y(_02111_),
    .A(_02090_),
    .B(_02110_));
 sg13g2_xnor2_1 _23812_ (.Y(_02112_),
    .A(_02098_),
    .B(_02111_));
 sg13g2_buf_1 _23813_ (.A(_02112_),
    .X(_02113_));
 sg13g2_nor2_1 _23814_ (.A(net760),
    .B(_02113_),
    .Y(_02114_));
 sg13g2_nand2_1 _23815_ (.Y(_02115_),
    .A(net760),
    .B(_02113_));
 sg13g2_o21ai_1 _23816_ (.B1(_02115_),
    .Y(_02116_),
    .A1(_13190_),
    .A2(_02114_));
 sg13g2_nand3_1 _23817_ (.B(_02106_),
    .C(_02116_),
    .A(_02095_),
    .Y(_02117_));
 sg13g2_and2_1 _23818_ (.A(_01692_),
    .B(_02094_),
    .X(_02118_));
 sg13g2_o21ai_1 _23819_ (.B1(_02113_),
    .Y(_02120_),
    .A1(net760),
    .A2(_02118_));
 sg13g2_a21oi_1 _23820_ (.A1(_13238_),
    .A2(_02113_),
    .Y(_02121_),
    .B1(net760));
 sg13g2_nor2_1 _23821_ (.A(_02095_),
    .B(_02121_),
    .Y(_02122_));
 sg13g2_a221oi_1 _23822_ (.B2(net446),
    .C1(_02122_),
    .B1(_02120_),
    .A1(_02095_),
    .Y(_02123_),
    .A2(_02114_));
 sg13g2_buf_1 _23823_ (.A(net761),
    .X(_02124_));
 sg13g2_nor2_1 _23824_ (.A(net431),
    .B(net420),
    .Y(_02125_));
 sg13g2_nor2_1 _23825_ (.A(net782),
    .B(_02105_),
    .Y(_02126_));
 sg13g2_or2_1 _23826_ (.X(_02127_),
    .B(_02126_),
    .A(_02099_));
 sg13g2_a22oi_1 _23827_ (.Y(_02128_),
    .B1(_02127_),
    .B2(_00678_),
    .A2(_02103_),
    .A1(_02125_));
 sg13g2_o21ai_1 _23828_ (.B1(_00644_),
    .Y(_02129_),
    .A1(_13264_),
    .A2(net763));
 sg13g2_nand3_1 _23829_ (.B(_02129_),
    .C(_02125_),
    .A(_00678_),
    .Y(_02131_));
 sg13g2_o21ai_1 _23830_ (.B1(_02131_),
    .Y(_02132_),
    .A1(net421),
    .A2(_02128_));
 sg13g2_mux2_1 _23831_ (.A0(_02117_),
    .A1(_02123_),
    .S(_02132_),
    .X(_02133_));
 sg13g2_xnor2_1 _23832_ (.Y(_02134_),
    .A(_01984_),
    .B(_02113_));
 sg13g2_o21ai_1 _23833_ (.B1(_01627_),
    .Y(_02135_),
    .A1(net168),
    .A2(_02134_));
 sg13g2_nand2_1 _23834_ (.Y(_02136_),
    .A(_01951_),
    .B(_02135_));
 sg13g2_a21o_1 _23835_ (.A2(_02133_),
    .A1(_05815_),
    .B1(_02136_),
    .X(_02137_));
 sg13g2_a21oi_1 _23836_ (.A1(_02089_),
    .A2(_02137_),
    .Y(_00487_),
    .B1(net440));
 sg13g2_buf_1 _23837_ (.A(_00263_),
    .X(_02138_));
 sg13g2_inv_1 _23838_ (.Y(_02139_),
    .A(_02138_));
 sg13g2_nor2_1 _23839_ (.A(net443),
    .B(_02139_),
    .Y(_02141_));
 sg13g2_buf_2 _23840_ (.A(\grid.cell_4_3.se ),
    .X(_02142_));
 sg13g2_xor2_1 _23841_ (.B(_02142_),
    .A(_01743_),
    .X(_02143_));
 sg13g2_buf_2 _23842_ (.A(_02143_),
    .X(_02144_));
 sg13g2_xnor2_1 _23843_ (.Y(_02145_),
    .A(_00670_),
    .B(_02144_));
 sg13g2_xnor2_1 _23844_ (.Y(_02146_),
    .A(net761),
    .B(_02145_));
 sg13g2_xnor2_1 _23845_ (.Y(_02147_),
    .A(net432),
    .B(_02146_));
 sg13g2_inv_1 _23846_ (.Y(_02148_),
    .A(_01759_));
 sg13g2_a22oi_1 _23847_ (.Y(_02149_),
    .B1(_02148_),
    .B2(_02146_),
    .A2(_02139_),
    .A1(_13298_));
 sg13g2_o21ai_1 _23848_ (.B1(_02149_),
    .Y(_02150_),
    .A1(_02141_),
    .A2(_02147_));
 sg13g2_buf_1 _23849_ (.A(net420),
    .X(_02152_));
 sg13g2_buf_1 _23850_ (.A(_02142_),
    .X(_02153_));
 sg13g2_nand2_1 _23851_ (.Y(_02154_),
    .A(net770),
    .B(net759));
 sg13g2_a22oi_1 _23852_ (.Y(_02155_),
    .B1(_02154_),
    .B2(_00717_),
    .A2(_02144_),
    .A1(net441));
 sg13g2_a21oi_1 _23853_ (.A1(net782),
    .A2(net420),
    .Y(_02156_),
    .B1(net439));
 sg13g2_or3_1 _23854_ (.A(net770),
    .B(net759),
    .C(_02156_),
    .X(_02157_));
 sg13g2_o21ai_1 _23855_ (.B1(_02157_),
    .Y(_02158_),
    .A1(net199),
    .A2(_02155_));
 sg13g2_buf_1 _23856_ (.A(net759),
    .X(_02159_));
 sg13g2_nor3_1 _23857_ (.A(net199),
    .B(net428),
    .C(net419),
    .Y(_02160_));
 sg13g2_a22oi_1 _23858_ (.Y(_02161_),
    .B1(_02160_),
    .B2(_00673_),
    .A2(_02158_),
    .A1(_00724_));
 sg13g2_xor2_1 _23859_ (.B(_02161_),
    .A(_02150_),
    .X(_02163_));
 sg13g2_nand2_1 _23860_ (.Y(_02164_),
    .A(net441),
    .B(_02144_));
 sg13g2_o21ai_1 _23861_ (.B1(_02164_),
    .Y(_02165_),
    .A1(_00647_),
    .A2(_02154_));
 sg13g2_nand2_1 _23862_ (.Y(_02166_),
    .A(_00735_),
    .B(_02165_));
 sg13g2_o21ai_1 _23863_ (.B1(_02166_),
    .Y(_02167_),
    .A1(_00724_),
    .A2(_02154_));
 sg13g2_nor2_1 _23864_ (.A(_02138_),
    .B(_01621_),
    .Y(_02168_));
 sg13g2_and2_1 _23865_ (.A(_02148_),
    .B(_02146_),
    .X(_02169_));
 sg13g2_nor3_1 _23866_ (.A(net199),
    .B(_00673_),
    .C(_02154_),
    .Y(_02170_));
 sg13g2_a221oi_1 _23867_ (.B2(_02169_),
    .C1(_02170_),
    .B1(_02168_),
    .A1(net199),
    .Y(_02171_),
    .A2(_02167_));
 sg13g2_a21oi_1 _23868_ (.A1(_02163_),
    .A2(_02171_),
    .Y(_02172_),
    .B1(net97));
 sg13g2_xor2_1 _23869_ (.B(_02146_),
    .A(_02024_),
    .X(_02174_));
 sg13g2_a21oi_1 _23870_ (.A1(_13104_),
    .A2(_02174_),
    .Y(_02175_),
    .B1(net202));
 sg13g2_or3_1 _23871_ (.A(_02082_),
    .B(_02172_),
    .C(_02175_),
    .X(_02176_));
 sg13g2_o21ai_1 _23872_ (.B1(_02176_),
    .Y(_00488_),
    .A1(net26),
    .A2(_01951_));
 sg13g2_buf_1 _23873_ (.A(\grid.cell_4_4.se ),
    .X(_02177_));
 sg13g2_buf_1 _23874_ (.A(_02177_),
    .X(_02178_));
 sg13g2_nand2_1 _23875_ (.Y(_02179_),
    .A(net1079),
    .B(net758));
 sg13g2_xor2_1 _23876_ (.B(_02177_),
    .A(net1079),
    .X(_02180_));
 sg13g2_and2_1 _23877_ (.A(net780),
    .B(_02180_),
    .X(_02181_));
 sg13g2_a21oi_1 _23878_ (.A1(_00718_),
    .A2(_02179_),
    .Y(_02182_),
    .B1(_02181_));
 sg13g2_inv_1 _23879_ (.Y(_02184_),
    .A(net758));
 sg13g2_buf_1 _23880_ (.A(_02184_),
    .X(_02185_));
 sg13g2_inv_1 _23881_ (.Y(_02186_),
    .A(_02142_));
 sg13g2_o21ai_1 _23882_ (.B1(net779),
    .Y(_02187_),
    .A1(net439),
    .A2(_02186_));
 sg13g2_nand3_1 _23883_ (.B(net198),
    .C(_02187_),
    .A(_01808_),
    .Y(_02188_));
 sg13g2_o21ai_1 _23884_ (.B1(_02188_),
    .Y(_02189_),
    .A1(net419),
    .A2(_02182_));
 sg13g2_buf_1 _23885_ (.A(net758),
    .X(_02190_));
 sg13g2_nor4_1 _23886_ (.A(net759),
    .B(net769),
    .C(net418),
    .D(_00719_),
    .Y(_02191_));
 sg13g2_a21o_1 _23887_ (.A2(_02189_),
    .A1(_00763_),
    .B1(_02191_),
    .X(_02192_));
 sg13g2_buf_1 _23888_ (.A(_00036_),
    .X(_02193_));
 sg13g2_xnor2_1 _23889_ (.Y(_02195_),
    .A(_02177_),
    .B(_01792_));
 sg13g2_xnor2_1 _23890_ (.Y(_02196_),
    .A(_00664_),
    .B(_02142_));
 sg13g2_xnor2_1 _23891_ (.Y(_02197_),
    .A(_02195_),
    .B(_02196_));
 sg13g2_buf_1 _23892_ (.A(_02197_),
    .X(_02198_));
 sg13g2_a21o_1 _23893_ (.A2(_02198_),
    .A1(_01753_),
    .B1(_00647_),
    .X(_02199_));
 sg13g2_o21ai_1 _23894_ (.B1(_02198_),
    .Y(_02200_),
    .A1(net1078),
    .A2(net442));
 sg13g2_nor2b_1 _23895_ (.A(_01727_),
    .B_N(net442),
    .Y(_02201_));
 sg13g2_a221oi_1 _23896_ (.B2(net202),
    .C1(_02201_),
    .B1(_02200_),
    .A1(_01788_),
    .Y(_02202_),
    .A2(_02199_));
 sg13g2_xnor2_1 _23897_ (.Y(_02203_),
    .A(_01753_),
    .B(_02198_));
 sg13g2_nor2b_1 _23898_ (.A(net1078),
    .B_N(_02198_),
    .Y(_02204_));
 sg13g2_a22oi_1 _23899_ (.Y(_02206_),
    .B1(_02204_),
    .B2(_02193_),
    .A2(_02203_),
    .A1(net442));
 sg13g2_o21ai_1 _23900_ (.B1(_02206_),
    .Y(_02207_),
    .A1(_02193_),
    .A2(_02202_));
 sg13g2_nor3_1 _23901_ (.A(net419),
    .B(_00711_),
    .C(_02179_),
    .Y(_02208_));
 sg13g2_nor2_1 _23902_ (.A(net780),
    .B(_02179_),
    .Y(_02209_));
 sg13g2_o21ai_1 _23903_ (.B1(net437),
    .Y(_02210_),
    .A1(_02181_),
    .A2(_02209_));
 sg13g2_or2_1 _23904_ (.X(_02211_),
    .B(_02179_),
    .A(_00763_));
 sg13g2_a21oi_1 _23905_ (.A1(_02210_),
    .A2(_02211_),
    .Y(_02212_),
    .B1(_02186_));
 sg13g2_nor4_1 _23906_ (.A(_02192_),
    .B(_02204_),
    .C(_02208_),
    .D(_02212_),
    .Y(_02213_));
 sg13g2_nor2_1 _23907_ (.A(net442),
    .B(_02203_),
    .Y(_02214_));
 sg13g2_inv_1 _23908_ (.Y(_02215_),
    .A(_02193_));
 sg13g2_a21oi_1 _23909_ (.A1(net442),
    .A2(_02203_),
    .Y(_02217_),
    .B1(_02215_));
 sg13g2_or2_1 _23910_ (.X(_02218_),
    .B(_02217_),
    .A(_02214_));
 sg13g2_a221oi_1 _23911_ (.B2(_02218_),
    .C1(net106),
    .B1(_02213_),
    .A1(_02192_),
    .Y(_02219_),
    .A2(_02207_));
 sg13g2_xor2_1 _23912_ (.B(_02198_),
    .A(_02093_),
    .X(_02220_));
 sg13g2_a21oi_1 _23913_ (.A1(_13104_),
    .A2(_02220_),
    .Y(_02221_),
    .B1(_01770_));
 sg13g2_or3_1 _23914_ (.A(_02082_),
    .B(_02219_),
    .C(_02221_),
    .X(_02222_));
 sg13g2_o21ai_1 _23915_ (.B1(_02222_),
    .Y(_00489_),
    .A1(net29),
    .A2(_02086_));
 sg13g2_buf_2 _23916_ (.A(\grid.cell_4_5.se ),
    .X(_02223_));
 sg13g2_nand2_2 _23917_ (.Y(_02224_),
    .A(net768),
    .B(_02223_));
 sg13g2_xor2_1 _23918_ (.B(_02223_),
    .A(_01821_),
    .X(_02225_));
 sg13g2_buf_2 _23919_ (.A(_02225_),
    .X(_02227_));
 sg13g2_nand2_1 _23920_ (.Y(_02228_),
    .A(net437),
    .B(_02227_));
 sg13g2_o21ai_1 _23921_ (.B1(_02228_),
    .Y(_02229_),
    .A1(_00736_),
    .A2(_02224_));
 sg13g2_nor2_1 _23922_ (.A(_00827_),
    .B(_02224_),
    .Y(_02230_));
 sg13g2_a21oi_1 _23923_ (.A1(net205),
    .A2(_02229_),
    .Y(_02231_),
    .B1(_02230_));
 sg13g2_nor2_1 _23924_ (.A(net198),
    .B(_02231_),
    .Y(_02232_));
 sg13g2_nor3_1 _23925_ (.A(net418),
    .B(_00756_),
    .C(_02224_),
    .Y(_02233_));
 sg13g2_a22oi_1 _23926_ (.Y(_02234_),
    .B1(_02224_),
    .B2(_00771_),
    .A2(_02227_),
    .A1(net779));
 sg13g2_buf_1 _23927_ (.A(_02223_),
    .X(_02235_));
 sg13g2_nor2_1 _23928_ (.A(net768),
    .B(net757),
    .Y(_02236_));
 sg13g2_o21ai_1 _23929_ (.B1(net436),
    .Y(_02238_),
    .A1(_00718_),
    .A2(net198));
 sg13g2_nand2_1 _23930_ (.Y(_02239_),
    .A(_02236_),
    .B(_02238_));
 sg13g2_o21ai_1 _23931_ (.B1(_02239_),
    .Y(_02240_),
    .A1(net418),
    .A2(_02234_));
 sg13g2_and2_1 _23932_ (.A(_00756_),
    .B(_02236_),
    .X(_02241_));
 sg13g2_a22oi_1 _23933_ (.Y(_02242_),
    .B1(_02241_),
    .B2(net198),
    .A2(_02240_),
    .A1(_00827_));
 sg13g2_buf_1 _23934_ (.A(_00068_),
    .X(_02243_));
 sg13g2_xnor2_1 _23935_ (.Y(_02244_),
    .A(net758),
    .B(net778));
 sg13g2_xnor2_1 _23936_ (.Y(_02245_),
    .A(_00713_),
    .B(_02244_));
 sg13g2_xnor2_1 _23937_ (.Y(_02246_),
    .A(_02227_),
    .B(_02245_));
 sg13g2_xnor2_1 _23938_ (.Y(_02247_),
    .A(net429),
    .B(_02246_));
 sg13g2_nor2_1 _23939_ (.A(_02243_),
    .B(_02247_),
    .Y(_02249_));
 sg13g2_xnor2_1 _23940_ (.Y(_02250_),
    .A(_02144_),
    .B(_02246_));
 sg13g2_a21oi_1 _23941_ (.A1(net172),
    .A2(_02250_),
    .Y(_02251_),
    .B1(net427));
 sg13g2_a21o_1 _23942_ (.A2(_02249_),
    .A1(_02242_),
    .B1(_02251_),
    .X(_02252_));
 sg13g2_nor4_1 _23943_ (.A(_02085_),
    .B(_02232_),
    .C(_02233_),
    .D(_02252_),
    .Y(_02253_));
 sg13g2_xnor2_1 _23944_ (.Y(_02254_),
    .A(net758),
    .B(net757));
 sg13g2_xor2_1 _23945_ (.B(_02254_),
    .A(_01825_),
    .X(_02255_));
 sg13g2_xnor2_1 _23946_ (.Y(_02256_),
    .A(_00710_),
    .B(_02255_));
 sg13g2_xnor2_1 _23947_ (.Y(_02257_),
    .A(net429),
    .B(_02256_));
 sg13g2_a22oi_1 _23948_ (.Y(_02258_),
    .B1(_02257_),
    .B2(_00735_),
    .A2(_02256_),
    .A1(_01853_));
 sg13g2_nor2_1 _23949_ (.A(_02242_),
    .B(_02249_),
    .Y(_02260_));
 sg13g2_xor2_1 _23950_ (.B(_02260_),
    .A(_02258_),
    .X(_02261_));
 sg13g2_a21oi_1 _23951_ (.A1(net427),
    .A2(net120),
    .Y(_02262_),
    .B1(_02085_));
 sg13g2_a21oi_1 _23952_ (.A1(_05002_),
    .A2(_02085_),
    .Y(_02263_),
    .B1(_02262_));
 sg13g2_a21oi_1 _23953_ (.A1(_02253_),
    .A2(_02261_),
    .Y(_02264_),
    .B1(_02263_));
 sg13g2_nor2_1 _23954_ (.A(net214),
    .B(_02264_),
    .Y(_00490_));
 sg13g2_buf_1 _23955_ (.A(_00130_),
    .X(_02265_));
 sg13g2_nor2_1 _23956_ (.A(net1074),
    .B(_02006_),
    .Y(_02266_));
 sg13g2_buf_1 _23957_ (.A(net757),
    .X(_02267_));
 sg13g2_nand3_1 _23958_ (.B(net417),
    .C(_02006_),
    .A(net1074),
    .Y(_02268_));
 sg13g2_nor2b_1 _23959_ (.A(_02266_),
    .B_N(_02268_),
    .Y(_02270_));
 sg13g2_xor2_1 _23960_ (.B(net417),
    .A(net1074),
    .X(_02271_));
 sg13g2_nand2b_1 _23961_ (.Y(_02272_),
    .B(_02271_),
    .A_N(_01974_));
 sg13g2_a21oi_1 _23962_ (.A1(_02270_),
    .A2(_02272_),
    .Y(_02273_),
    .B1(_00799_));
 sg13g2_inv_1 _23963_ (.Y(_02274_),
    .A(_02223_));
 sg13g2_nand2_1 _23964_ (.Y(_02275_),
    .A(net756),
    .B(_01974_));
 sg13g2_nor2_1 _23965_ (.A(net417),
    .B(_01977_),
    .Y(_02276_));
 sg13g2_o21ai_1 _23966_ (.B1(net1074),
    .Y(_02277_),
    .A1(_01974_),
    .A2(_02276_));
 sg13g2_a21oi_1 _23967_ (.A1(_02275_),
    .A2(_02277_),
    .Y(_02278_),
    .B1(net207));
 sg13g2_nand3_1 _23968_ (.B(net445),
    .C(_01977_),
    .A(net417),
    .Y(_02279_));
 sg13g2_a21oi_1 _23969_ (.A1(_02275_),
    .A2(_02279_),
    .Y(_02281_),
    .B1(_00778_));
 sg13g2_nor3_1 _23970_ (.A(net1074),
    .B(net756),
    .C(_02006_),
    .Y(_02282_));
 sg13g2_nor4_1 _23971_ (.A(_02273_),
    .B(_02278_),
    .C(_02281_),
    .D(_02282_),
    .Y(_02283_));
 sg13g2_buf_1 _23972_ (.A(_00100_),
    .X(_02284_));
 sg13g2_inv_1 _23973_ (.Y(_02285_),
    .A(_02284_));
 sg13g2_xnor2_1 _23974_ (.Y(_02286_),
    .A(_02223_),
    .B(_01955_));
 sg13g2_xnor2_1 _23975_ (.Y(_02287_),
    .A(_01605_),
    .B(_02286_));
 sg13g2_xnor2_1 _23976_ (.Y(_02288_),
    .A(net436),
    .B(_02287_));
 sg13g2_xnor2_1 _23977_ (.Y(_02289_),
    .A(_01808_),
    .B(_02288_));
 sg13g2_o21ai_1 _23978_ (.B1(_02289_),
    .Y(_02290_),
    .A1(_02285_),
    .A2(net437));
 sg13g2_nand2b_1 _23979_ (.Y(_02292_),
    .B(_02288_),
    .A_N(_01875_));
 sg13g2_nand2_1 _23980_ (.Y(_02293_),
    .A(_02285_),
    .B(net437));
 sg13g2_nand3_1 _23981_ (.B(_02292_),
    .C(_02293_),
    .A(_02290_),
    .Y(_02294_));
 sg13g2_xnor2_1 _23982_ (.Y(_02295_),
    .A(_02283_),
    .B(_02294_));
 sg13g2_xor2_1 _23983_ (.B(_02288_),
    .A(_02195_),
    .X(_02296_));
 sg13g2_nor3_1 _23984_ (.A(_02284_),
    .B(_01783_),
    .C(_02292_),
    .Y(_02297_));
 sg13g2_nand2_1 _23985_ (.Y(_02298_),
    .A(net436),
    .B(_02007_));
 sg13g2_o21ai_1 _23986_ (.B1(_02298_),
    .Y(_02299_),
    .A1(net436),
    .A2(_02006_));
 sg13g2_a21oi_1 _23987_ (.A1(_13244_),
    .A2(_02299_),
    .Y(_02300_),
    .B1(_02266_));
 sg13g2_nor2_1 _23988_ (.A(net756),
    .B(_02300_),
    .Y(_02301_));
 sg13g2_buf_1 _23989_ (.A(net417),
    .X(_02303_));
 sg13g2_nor3_1 _23990_ (.A(net197),
    .B(_00799_),
    .C(_02006_),
    .Y(_02304_));
 sg13g2_nor4_1 _23991_ (.A(_03821_),
    .B(_02297_),
    .C(_02301_),
    .D(_02304_),
    .Y(_02305_));
 sg13g2_o21ai_1 _23992_ (.B1(_02305_),
    .Y(_02306_),
    .A1(net201),
    .A2(_02296_));
 sg13g2_or2_1 _23993_ (.X(_02307_),
    .B(_02306_),
    .A(_02295_));
 sg13g2_a22oi_1 _23994_ (.Y(_02308_),
    .B1(net25),
    .B2(_01950_),
    .A2(net72),
    .A1(_01865_));
 sg13g2_a221oi_1 _23995_ (.B2(_02308_),
    .C1(net557),
    .B1(_02307_),
    .A1(_06813_),
    .Y(_00491_),
    .A2(_01950_));
 sg13g2_nand2_1 _23996_ (.Y(_02309_),
    .A(_02223_),
    .B(_01955_));
 sg13g2_buf_2 _23997_ (.A(_02309_),
    .X(_02310_));
 sg13g2_o21ai_1 _23998_ (.B1(_01821_),
    .Y(_02311_),
    .A1(_02223_),
    .A2(net766));
 sg13g2_a21o_1 _23999_ (.A2(_02311_),
    .A1(_02310_),
    .B1(_13194_),
    .X(_02313_));
 sg13g2_mux2_1 _24000_ (.A0(net757),
    .A1(_02310_),
    .S(_01821_),
    .X(_02314_));
 sg13g2_a22oi_1 _24001_ (.Y(_02315_),
    .B1(_02314_),
    .B2(net785),
    .A2(_02236_),
    .A1(net424));
 sg13g2_mux2_1 _24002_ (.A0(_02313_),
    .A1(_02315_),
    .S(net1074),
    .X(_02316_));
 sg13g2_nand2_1 _24003_ (.Y(_02317_),
    .A(net785),
    .B(net766));
 sg13g2_nand3_1 _24004_ (.B(net756),
    .C(_02003_),
    .A(_01887_),
    .Y(_02318_));
 sg13g2_o21ai_1 _24005_ (.B1(_02318_),
    .Y(_02319_),
    .A1(_02224_),
    .A2(_02317_));
 sg13g2_nor2_1 _24006_ (.A(net1074),
    .B(_02310_),
    .Y(_02320_));
 sg13g2_nand3_1 _24007_ (.B(_02310_),
    .C(_02311_),
    .A(_02265_),
    .Y(_02321_));
 sg13g2_a21oi_1 _24008_ (.A1(_02318_),
    .A2(_02321_),
    .Y(_02322_),
    .B1(_13195_));
 sg13g2_a221oi_1 _24009_ (.B2(net426),
    .C1(_02322_),
    .B1(_02320_),
    .A1(_00771_),
    .Y(_02324_),
    .A2(_02319_));
 sg13g2_o21ai_1 _24010_ (.B1(_02324_),
    .Y(_02325_),
    .A1(_00771_),
    .A2(_02316_));
 sg13g2_buf_1 _24011_ (.A(_02325_),
    .X(_02326_));
 sg13g2_nor3_1 _24012_ (.A(net777),
    .B(net764),
    .C(_01589_),
    .Y(_02327_));
 sg13g2_nor2_1 _24013_ (.A(net774),
    .B(net765),
    .Y(_02328_));
 sg13g2_a22oi_1 _24014_ (.Y(_02329_),
    .B1(_02328_),
    .B2(_02020_),
    .A2(_02327_),
    .A1(_02326_));
 sg13g2_a21oi_1 _24015_ (.A1(net764),
    .A2(_01990_),
    .Y(_02330_),
    .B1(_01589_));
 sg13g2_and2_1 _24016_ (.A(_01988_),
    .B(net1080),
    .X(_02331_));
 sg13g2_nand2_1 _24017_ (.Y(_02332_),
    .A(net774),
    .B(_02331_));
 sg13g2_mux2_1 _24018_ (.A0(_02330_),
    .A1(_02332_),
    .S(_02326_),
    .X(_02333_));
 sg13g2_xor2_1 _24019_ (.B(_02286_),
    .A(_01825_),
    .X(_02335_));
 sg13g2_xnor2_1 _24020_ (.Y(_02336_),
    .A(_13194_),
    .B(_02335_));
 sg13g2_a21oi_1 _24021_ (.A1(_02329_),
    .A2(_02333_),
    .Y(_02337_),
    .B1(_02336_));
 sg13g2_xnor2_1 _24022_ (.Y(_02338_),
    .A(net764),
    .B(_01996_));
 sg13g2_xnor2_1 _24023_ (.Y(_02339_),
    .A(_02336_),
    .B(_02338_));
 sg13g2_nor2_1 _24024_ (.A(net203),
    .B(_02339_),
    .Y(_02340_));
 sg13g2_nor3_1 _24025_ (.A(net201),
    .B(_00799_),
    .C(_02310_),
    .Y(_02341_));
 sg13g2_nand2b_1 _24026_ (.Y(_02342_),
    .B(_00776_),
    .A_N(_02286_));
 sg13g2_o21ai_1 _24027_ (.B1(_02342_),
    .Y(_02343_),
    .A1(_00778_),
    .A2(_02310_));
 sg13g2_a21oi_1 _24028_ (.A1(_13244_),
    .A2(_02343_),
    .Y(_02344_),
    .B1(_02320_));
 sg13g2_xnor2_1 _24029_ (.Y(_02346_),
    .A(_13195_),
    .B(_02335_));
 sg13g2_nor2_1 _24030_ (.A(net764),
    .B(_01988_),
    .Y(_02347_));
 sg13g2_nand4_1 _24031_ (.B(_01589_),
    .C(_02346_),
    .A(net777),
    .Y(_02348_),
    .D(_02347_));
 sg13g2_o21ai_1 _24032_ (.B1(_02348_),
    .Y(_02349_),
    .A1(_01887_),
    .A2(_02344_));
 sg13g2_nor4_1 _24033_ (.A(net125),
    .B(_02340_),
    .C(_02341_),
    .D(_02349_),
    .Y(_02350_));
 sg13g2_nand2_1 _24034_ (.Y(_02351_),
    .A(net764),
    .B(_01988_));
 sg13g2_o21ai_1 _24035_ (.B1(_02351_),
    .Y(_02352_),
    .A1(_01551_),
    .A2(_02347_));
 sg13g2_a22oi_1 _24036_ (.Y(_02353_),
    .B1(_02352_),
    .B2(_02336_),
    .A2(_02331_),
    .A1(_13230_));
 sg13g2_o21ai_1 _24037_ (.B1(_01988_),
    .Y(_02354_),
    .A1(net764),
    .A2(_02346_));
 sg13g2_a221oi_1 _24038_ (.B2(net777),
    .C1(_02326_),
    .B1(_02354_),
    .A1(_02336_),
    .Y(_02355_),
    .A2(_02347_));
 sg13g2_a21o_1 _24039_ (.A2(_02353_),
    .A1(_02326_),
    .B1(_02355_),
    .X(_02357_));
 sg13g2_nand3b_1 _24040_ (.B(_02350_),
    .C(_02357_),
    .Y(_02358_),
    .A_N(_02337_));
 sg13g2_a21oi_1 _24041_ (.A1(net203),
    .A2(_07561_),
    .Y(_02359_),
    .B1(_02085_));
 sg13g2_a221oi_1 _24042_ (.B2(_02359_),
    .C1(net557),
    .B1(_02358_),
    .A1(_05129_),
    .Y(_00492_),
    .A2(_02085_));
 sg13g2_nor2_2 _24043_ (.A(_06474_),
    .B(_09520_),
    .Y(_02360_));
 sg13g2_inv_1 _24044_ (.Y(_02361_),
    .A(_02360_));
 sg13g2_nor2_2 _24045_ (.A(net176),
    .B(_02361_),
    .Y(_02362_));
 sg13g2_nand2_1 _24046_ (.Y(_02363_),
    .A(_05757_),
    .B(_02362_));
 sg13g2_buf_1 _24047_ (.A(\grid.cell_5_0.se ),
    .X(_02364_));
 sg13g2_xnor2_1 _24048_ (.Y(_02365_),
    .A(net1081),
    .B(net1073));
 sg13g2_xnor2_1 _24049_ (.Y(_02367_),
    .A(net1076),
    .B(_02365_));
 sg13g2_buf_2 _24050_ (.A(\grid.cell_5_0.sw ),
    .X(_02368_));
 sg13g2_inv_2 _24051_ (.Y(_02369_),
    .A(_02368_));
 sg13g2_xnor2_1 _24052_ (.Y(_02370_),
    .A(_02369_),
    .B(_02007_));
 sg13g2_xnor2_1 _24053_ (.Y(_02371_),
    .A(net764),
    .B(_02370_));
 sg13g2_xnor2_1 _24054_ (.Y(_02372_),
    .A(_02367_),
    .B(_02371_));
 sg13g2_buf_1 _24055_ (.A(_00262_),
    .X(_02373_));
 sg13g2_inv_2 _24056_ (.Y(_02374_),
    .A(_02373_));
 sg13g2_nand2b_1 _24057_ (.Y(_02375_),
    .B(_02374_),
    .A_N(_02372_));
 sg13g2_buf_1 _24058_ (.A(net1073),
    .X(_02376_));
 sg13g2_inv_1 _24059_ (.Y(_02378_),
    .A(net755));
 sg13g2_buf_1 _24060_ (.A(_02368_),
    .X(_02379_));
 sg13g2_nand2_1 _24061_ (.Y(_02380_),
    .A(net766),
    .B(net754));
 sg13g2_buf_1 _24062_ (.A(_02380_),
    .X(_02381_));
 sg13g2_xor2_1 _24063_ (.B(_02368_),
    .A(_01955_),
    .X(_02382_));
 sg13g2_a22oi_1 _24064_ (.Y(_02383_),
    .B1(_02382_),
    .B2(net1081),
    .A2(_02381_),
    .A1(_01584_));
 sg13g2_nor2_2 _24065_ (.A(net424),
    .B(net754),
    .Y(_02384_));
 sg13g2_nand2_1 _24066_ (.Y(_02385_),
    .A(net1081),
    .B(net775));
 sg13g2_nand2_1 _24067_ (.Y(_02386_),
    .A(_02384_),
    .B(_02385_));
 sg13g2_o21ai_1 _24068_ (.B1(_02386_),
    .Y(_02387_),
    .A1(_01692_),
    .A2(_02383_));
 sg13g2_buf_1 _24069_ (.A(net754),
    .X(_02389_));
 sg13g2_nand2b_1 _24070_ (.Y(_02390_),
    .B(_01691_),
    .A_N(net415));
 sg13g2_a21oi_1 _24071_ (.A1(_01553_),
    .A2(_02376_),
    .Y(_02391_),
    .B1(_01584_));
 sg13g2_nor3_1 _24072_ (.A(net134),
    .B(_02390_),
    .C(_02391_),
    .Y(_02392_));
 sg13g2_a21oi_1 _24073_ (.A1(net416),
    .A2(_02387_),
    .Y(_02393_),
    .B1(_02392_));
 sg13g2_inv_1 _24074_ (.Y(_02394_),
    .A(net760));
 sg13g2_xnor2_1 _24075_ (.Y(_02395_),
    .A(_02365_),
    .B(_02370_));
 sg13g2_xor2_1 _24076_ (.B(_02367_),
    .A(_02370_),
    .X(_02396_));
 sg13g2_a22oi_1 _24077_ (.Y(_02397_),
    .B1(_02396_),
    .B2(net774),
    .A2(_02395_),
    .A1(_02394_));
 sg13g2_nand2b_1 _24078_ (.Y(_02398_),
    .B(_02397_),
    .A_N(_02393_));
 sg13g2_buf_1 _24079_ (.A(net754),
    .X(_02400_));
 sg13g2_nand2b_1 _24080_ (.Y(_02401_),
    .B(net414),
    .A_N(_01691_));
 sg13g2_o21ai_1 _24081_ (.B1(_02401_),
    .Y(_02402_),
    .A1(net414),
    .A2(_02385_));
 sg13g2_nor2_1 _24082_ (.A(net414),
    .B(net771),
    .Y(_02403_));
 sg13g2_nor3_1 _24083_ (.A(net200),
    .B(_02385_),
    .C(_02403_),
    .Y(_02404_));
 sg13g2_a21oi_1 _24084_ (.A1(net134),
    .A2(_02402_),
    .Y(_02405_),
    .B1(_02404_));
 sg13g2_nor2_1 _24085_ (.A(net416),
    .B(_02405_),
    .Y(_02406_));
 sg13g2_buf_1 _24086_ (.A(net755),
    .X(_02407_));
 sg13g2_nor2b_1 _24087_ (.A(_01691_),
    .B_N(net415),
    .Y(_02408_));
 sg13g2_o21ai_1 _24088_ (.B1(_02390_),
    .Y(_02409_),
    .A1(_01959_),
    .A2(_02408_));
 sg13g2_nand2_1 _24089_ (.Y(_02411_),
    .A(net414),
    .B(net771));
 sg13g2_o21ai_1 _24090_ (.B1(net424),
    .Y(_02412_),
    .A1(net415),
    .A2(_01691_));
 sg13g2_a21oi_1 _24091_ (.A1(_02411_),
    .A2(_02412_),
    .Y(_02413_),
    .B1(_02385_));
 sg13g2_a21oi_1 _24092_ (.A1(_01584_),
    .A2(_02409_),
    .Y(_02414_),
    .B1(_02413_));
 sg13g2_or3_1 _24093_ (.A(net1073),
    .B(net424),
    .C(net415),
    .X(_02415_));
 sg13g2_nand4_1 _24094_ (.B(net775),
    .C(_01958_),
    .A(net1073),
    .Y(_02416_),
    .D(net415));
 sg13g2_a21oi_1 _24095_ (.A1(_02415_),
    .A2(_02416_),
    .Y(_02417_),
    .B1(net776));
 sg13g2_nor3_1 _24096_ (.A(net433),
    .B(_01959_),
    .C(_02390_),
    .Y(_02418_));
 sg13g2_nor2_1 _24097_ (.A(_02417_),
    .B(_02418_),
    .Y(_02419_));
 sg13g2_o21ai_1 _24098_ (.B1(_02419_),
    .Y(_02420_),
    .A1(net413),
    .A2(_02414_));
 sg13g2_o21ai_1 _24099_ (.B1(_02397_),
    .Y(_02422_),
    .A1(_02406_),
    .A2(_02420_));
 sg13g2_nand2b_1 _24100_ (.Y(_02423_),
    .B(_02393_),
    .A_N(_02397_));
 sg13g2_nand3_1 _24101_ (.B(_02423_),
    .C(_02375_),
    .A(_02422_),
    .Y(_02424_));
 sg13g2_o21ai_1 _24102_ (.B1(_02424_),
    .Y(_02425_),
    .A1(_02375_),
    .A2(_02398_));
 sg13g2_buf_2 _24103_ (.A(\grid.cell_5_0.s ),
    .X(_02426_));
 sg13g2_buf_1 _24104_ (.A(_02426_),
    .X(_02427_));
 sg13g2_xnor2_1 _24105_ (.Y(_02428_),
    .A(net753),
    .B(_02372_));
 sg13g2_buf_1 _24106_ (.A(_01995_),
    .X(_02429_));
 sg13g2_a21oi_1 _24107_ (.A1(_05415_),
    .A2(_02428_),
    .Y(_02430_),
    .B1(net752));
 sg13g2_nor2_1 _24108_ (.A(_02362_),
    .B(_02430_),
    .Y(_02431_));
 sg13g2_o21ai_1 _24109_ (.B1(_02431_),
    .Y(_02433_),
    .A1(_06817_),
    .A2(_02425_));
 sg13g2_a21oi_1 _24110_ (.A1(_02363_),
    .A2(_02433_),
    .Y(_00493_),
    .B1(_00661_));
 sg13g2_nand2_1 _24111_ (.Y(_02434_),
    .A(_06112_),
    .B(_02360_));
 sg13g2_buf_1 _24112_ (.A(_02434_),
    .X(_02435_));
 sg13g2_buf_1 _24113_ (.A(\grid.cell_5_1.se ),
    .X(_02436_));
 sg13g2_buf_8 _24114_ (.A(_02436_),
    .X(_02437_));
 sg13g2_buf_1 _24115_ (.A(net751),
    .X(_02438_));
 sg13g2_nor2_1 _24116_ (.A(net412),
    .B(_01692_),
    .Y(_02439_));
 sg13g2_nor2b_1 _24117_ (.A(_01691_),
    .B_N(net751),
    .Y(_02440_));
 sg13g2_buf_1 _24118_ (.A(net751),
    .X(_02441_));
 sg13g2_nand2_1 _24119_ (.Y(_02443_),
    .A(net1081),
    .B(net773));
 sg13g2_nor2_1 _24120_ (.A(net411),
    .B(_02443_),
    .Y(_02444_));
 sg13g2_o21ai_1 _24121_ (.B1(net421),
    .Y(_02445_),
    .A1(_02440_),
    .A2(_02444_));
 sg13g2_nor2_1 _24122_ (.A(net422),
    .B(_02443_),
    .Y(_02446_));
 sg13g2_o21ai_1 _24123_ (.B1(_02446_),
    .Y(_02447_),
    .A1(net411),
    .A2(net771));
 sg13g2_nand3_1 _24124_ (.B(_02445_),
    .C(_02447_),
    .A(net413),
    .Y(_02448_));
 sg13g2_nor2_1 _24125_ (.A(net762),
    .B(_02440_),
    .Y(_02449_));
 sg13g2_or2_1 _24126_ (.X(_02450_),
    .B(_02449_),
    .A(_02439_));
 sg13g2_nand2_1 _24127_ (.Y(_02451_),
    .A(net412),
    .B(_01696_));
 sg13g2_o21ai_1 _24128_ (.B1(net762),
    .Y(_02452_),
    .A1(net412),
    .A2(_01696_));
 sg13g2_a21oi_1 _24129_ (.A1(_02451_),
    .A2(_02452_),
    .Y(_02454_),
    .B1(_02443_));
 sg13g2_a21oi_1 _24130_ (.A1(_01627_),
    .A2(_02450_),
    .Y(_02455_),
    .B1(_02454_));
 sg13g2_nand2_1 _24131_ (.Y(_02456_),
    .A(net416),
    .B(_02455_));
 sg13g2_inv_2 _24132_ (.Y(_02457_),
    .A(_02437_));
 sg13g2_nand3_1 _24133_ (.B(net763),
    .C(_02457_),
    .A(net416),
    .Y(_02458_));
 sg13g2_buf_1 _24134_ (.A(net411),
    .X(_02459_));
 sg13g2_nand4_1 _24135_ (.B(net430),
    .C(net422),
    .A(net413),
    .Y(_02460_),
    .D(net196));
 sg13g2_a21oi_1 _24136_ (.A1(_02458_),
    .A2(_02460_),
    .Y(_02461_),
    .B1(net204));
 sg13g2_a221oi_1 _24137_ (.B2(_02456_),
    .C1(_02461_),
    .B1(_02448_),
    .A1(_02036_),
    .Y(_02462_),
    .A2(_02439_));
 sg13g2_nand2_1 _24138_ (.Y(_02463_),
    .A(_02018_),
    .B(_02373_));
 sg13g2_xnor2_1 _24139_ (.Y(_02465_),
    .A(_02457_),
    .B(_02037_));
 sg13g2_xor2_1 _24140_ (.B(_02465_),
    .A(_02365_),
    .X(_02466_));
 sg13g2_xnor2_1 _24141_ (.Y(_02467_),
    .A(net752),
    .B(_02466_));
 sg13g2_nand2_1 _24142_ (.Y(_02468_),
    .A(_01596_),
    .B(_02374_));
 sg13g2_o21ai_1 _24143_ (.B1(_02468_),
    .Y(_02469_),
    .A1(net765),
    .A2(_02466_));
 sg13g2_a21oi_1 _24144_ (.A1(_02463_),
    .A2(_02467_),
    .Y(_02470_),
    .B1(_02469_));
 sg13g2_xnor2_1 _24145_ (.Y(_02471_),
    .A(_02462_),
    .B(_02470_));
 sg13g2_nand2_1 _24146_ (.Y(_02472_),
    .A(net422),
    .B(net411));
 sg13g2_xor2_1 _24147_ (.B(net751),
    .A(_02022_),
    .X(_02473_));
 sg13g2_nand2_1 _24148_ (.Y(_02474_),
    .A(net434),
    .B(_02473_));
 sg13g2_o21ai_1 _24149_ (.B1(_02474_),
    .Y(_02476_),
    .A1(net434),
    .A2(_02472_));
 sg13g2_a22oi_1 _24150_ (.Y(_02477_),
    .B1(_02476_),
    .B2(net430),
    .A2(_02440_),
    .A1(_02070_));
 sg13g2_nor2_1 _24151_ (.A(net416),
    .B(_02477_),
    .Y(_02478_));
 sg13g2_xor2_1 _24152_ (.B(_01995_),
    .A(_01595_),
    .X(_02479_));
 sg13g2_nor4_1 _24153_ (.A(_02373_),
    .B(net765),
    .C(_02479_),
    .D(_02466_),
    .Y(_02480_));
 sg13g2_nand4_1 _24154_ (.B(net416),
    .C(_01711_),
    .A(net204),
    .Y(_02481_),
    .D(net421));
 sg13g2_o21ai_1 _24155_ (.B1(net118),
    .Y(_02482_),
    .A1(_02457_),
    .A2(_02481_));
 sg13g2_inv_2 _24156_ (.Y(_02483_),
    .A(_02426_));
 sg13g2_xnor2_1 _24157_ (.Y(_02484_),
    .A(_02483_),
    .B(_02479_));
 sg13g2_xnor2_1 _24158_ (.Y(_02485_),
    .A(_02466_),
    .B(_02484_));
 sg13g2_nor2_1 _24159_ (.A(net425),
    .B(_02485_),
    .Y(_02487_));
 sg13g2_nor4_1 _24160_ (.A(_02478_),
    .B(_02480_),
    .C(_02482_),
    .D(_02487_),
    .Y(_02488_));
 sg13g2_a22oi_1 _24161_ (.Y(_02489_),
    .B1(_02471_),
    .B2(_02488_),
    .A2(_11411_),
    .A1(net425));
 sg13g2_o21ai_1 _24162_ (.B1(net435),
    .Y(_02490_),
    .A1(net38),
    .A2(_02435_));
 sg13g2_a21oi_1 _24163_ (.A1(_02435_),
    .A2(_02489_),
    .Y(_00494_),
    .B1(_02490_));
 sg13g2_buf_1 _24164_ (.A(\grid.cell_5_2.se ),
    .X(_02491_));
 sg13g2_buf_2 _24165_ (.A(_02491_),
    .X(_02492_));
 sg13g2_xnor2_1 _24166_ (.Y(_02493_),
    .A(net750),
    .B(_02098_));
 sg13g2_xnor2_1 _24167_ (.Y(_02494_),
    .A(net773),
    .B(net751));
 sg13g2_xnor2_1 _24168_ (.Y(_02495_),
    .A(_02493_),
    .B(_02494_));
 sg13g2_buf_1 _24169_ (.A(_02495_),
    .X(_02497_));
 sg13g2_xnor2_1 _24170_ (.Y(_02498_),
    .A(_02367_),
    .B(_02497_));
 sg13g2_o21ai_1 _24171_ (.B1(net763),
    .Y(_02499_),
    .A1(_06244_),
    .A2(_02498_));
 sg13g2_nand2_1 _24172_ (.Y(_02500_),
    .A(_04067_),
    .B(_02362_));
 sg13g2_buf_1 _24173_ (.A(net750),
    .X(_02501_));
 sg13g2_nand2_1 _24174_ (.Y(_02502_),
    .A(net420),
    .B(net410));
 sg13g2_xor2_1 _24175_ (.B(_02491_),
    .A(_02091_),
    .X(_02503_));
 sg13g2_nand2_1 _24176_ (.Y(_02504_),
    .A(net432),
    .B(_02503_));
 sg13g2_o21ai_1 _24177_ (.B1(_02504_),
    .Y(_02505_),
    .A1(_01711_),
    .A2(_02502_));
 sg13g2_nand2_1 _24178_ (.Y(_02506_),
    .A(_01727_),
    .B(_02505_));
 sg13g2_nand2b_1 _24179_ (.Y(_02508_),
    .B(_02148_),
    .A_N(_02502_));
 sg13g2_a21oi_1 _24180_ (.A1(_02506_),
    .A2(_02508_),
    .Y(_02509_),
    .B1(_02457_));
 sg13g2_nand2_1 _24181_ (.Y(_02510_),
    .A(_01618_),
    .B(net772));
 sg13g2_nor3_1 _24182_ (.A(net196),
    .B(_02502_),
    .C(_02510_),
    .Y(_02511_));
 sg13g2_buf_2 _24183_ (.A(_00261_),
    .X(_02512_));
 sg13g2_buf_1 _24184_ (.A(_02512_),
    .X(_02513_));
 sg13g2_nor2_1 _24185_ (.A(net423),
    .B(net749),
    .Y(_02514_));
 sg13g2_and4_1 _24186_ (.A(net204),
    .B(_02394_),
    .C(_02497_),
    .D(_02514_),
    .X(_02515_));
 sg13g2_nor4_1 _24187_ (.A(_00648_),
    .B(_02509_),
    .C(_02511_),
    .D(_02515_),
    .Y(_02516_));
 sg13g2_inv_1 _24188_ (.Y(_02517_),
    .A(_02497_));
 sg13g2_o21ai_1 _24189_ (.B1(net749),
    .Y(_02519_),
    .A1(net423),
    .A2(_02497_));
 sg13g2_a22oi_1 _24190_ (.Y(_02520_),
    .B1(_02519_),
    .B2(_01566_),
    .A2(_02514_),
    .A1(_02517_));
 sg13g2_inv_2 _24191_ (.Y(_02521_),
    .A(_02512_));
 sg13g2_nor2_1 _24192_ (.A(net434),
    .B(_02521_),
    .Y(_02522_));
 sg13g2_nand2_1 _24193_ (.Y(_02523_),
    .A(net423),
    .B(net749));
 sg13g2_o21ai_1 _24194_ (.B1(_02523_),
    .Y(_02524_),
    .A1(_01554_),
    .A2(_02514_));
 sg13g2_a22oi_1 _24195_ (.Y(_02525_),
    .B1(_02524_),
    .B2(_02517_),
    .A2(_02522_),
    .A1(net760));
 sg13g2_nor2_1 _24196_ (.A(_02092_),
    .B(net750),
    .Y(_02526_));
 sg13g2_a21oi_1 _24197_ (.A1(net761),
    .A2(net750),
    .Y(_02527_),
    .B1(_01679_));
 sg13g2_a21o_1 _24198_ (.A2(_02503_),
    .A1(_01618_),
    .B1(_02527_),
    .X(_02528_));
 sg13g2_a22oi_1 _24199_ (.Y(_02530_),
    .B1(_02528_),
    .B2(_01759_),
    .A2(_02526_),
    .A1(_02510_));
 sg13g2_o21ai_1 _24200_ (.B1(_01679_),
    .Y(_02531_),
    .A1(_01627_),
    .A2(_02457_));
 sg13g2_nand3_1 _24201_ (.B(_02531_),
    .C(_02526_),
    .A(_01759_),
    .Y(_02532_));
 sg13g2_o21ai_1 _24202_ (.B1(_02532_),
    .Y(_02533_),
    .A1(net411),
    .A2(_02530_));
 sg13g2_buf_1 _24203_ (.A(_02533_),
    .X(_02534_));
 sg13g2_mux2_1 _24204_ (.A0(_02520_),
    .A1(_02525_),
    .S(_02534_),
    .X(_02535_));
 sg13g2_nand4_1 _24205_ (.B(_02500_),
    .C(_02516_),
    .A(_02499_),
    .Y(_02536_),
    .D(_02535_));
 sg13g2_nand3_1 _24206_ (.B(net760),
    .C(_02534_),
    .A(net425),
    .Y(_02537_));
 sg13g2_nand3_1 _24207_ (.B(_02521_),
    .C(_02394_),
    .A(net423),
    .Y(_02538_));
 sg13g2_a21oi_1 _24208_ (.A1(_02537_),
    .A2(_02538_),
    .Y(_02539_),
    .B1(_01566_));
 sg13g2_nand3_1 _24209_ (.B(net749),
    .C(_02109_),
    .A(net425),
    .Y(_02541_));
 sg13g2_o21ai_1 _24210_ (.B1(_02109_),
    .Y(_02542_),
    .A1(_01954_),
    .A2(_02522_));
 sg13g2_nor2_1 _24211_ (.A(_02534_),
    .B(_02542_),
    .Y(_02543_));
 sg13g2_a21oi_1 _24212_ (.A1(_02534_),
    .A2(_02541_),
    .Y(_02544_),
    .B1(_02543_));
 sg13g2_o21ai_1 _24213_ (.B1(_02497_),
    .Y(_02545_),
    .A1(_02539_),
    .A2(_02544_));
 sg13g2_inv_1 _24214_ (.Y(_02546_),
    .A(_02545_));
 sg13g2_nand3_1 _24215_ (.B(_06055_),
    .C(_02435_),
    .A(_02070_),
    .Y(_02547_));
 sg13g2_o21ai_1 _24216_ (.B1(_02547_),
    .Y(_02548_),
    .A1(_04067_),
    .A2(_02435_));
 sg13g2_nand2_1 _24217_ (.Y(_02549_),
    .A(_05124_),
    .B(_02548_));
 sg13g2_o21ai_1 _24218_ (.B1(_02549_),
    .Y(_00495_),
    .A1(_02536_),
    .A2(_02546_));
 sg13g2_buf_1 _24219_ (.A(_00260_),
    .X(_02551_));
 sg13g2_inv_1 _24220_ (.Y(_02552_),
    .A(_02551_));
 sg13g2_nor2_1 _24221_ (.A(net432),
    .B(_02552_),
    .Y(_02553_));
 sg13g2_buf_2 _24222_ (.A(\grid.cell_5_3.se ),
    .X(_02554_));
 sg13g2_inv_2 _24223_ (.Y(_02555_),
    .A(_02554_));
 sg13g2_xnor2_1 _24224_ (.Y(_02556_),
    .A(_02555_),
    .B(_02144_));
 sg13g2_xnor2_1 _24225_ (.Y(_02557_),
    .A(_01677_),
    .B(net750));
 sg13g2_xnor2_1 _24226_ (.Y(_02558_),
    .A(_02556_),
    .B(_02557_));
 sg13g2_xnor2_1 _24227_ (.Y(_02559_),
    .A(net422),
    .B(_02558_));
 sg13g2_a22oi_1 _24228_ (.Y(_02560_),
    .B1(_02139_),
    .B2(_02558_),
    .A2(_02552_),
    .A1(net432));
 sg13g2_o21ai_1 _24229_ (.B1(_02560_),
    .Y(_02562_),
    .A1(_02553_),
    .A2(_02559_));
 sg13g2_buf_1 _24230_ (.A(net410),
    .X(_02563_));
 sg13g2_buf_1 _24231_ (.A(_02554_),
    .X(_02564_));
 sg13g2_xor2_1 _24232_ (.B(net748),
    .A(_02142_),
    .X(_02565_));
 sg13g2_nand2_1 _24233_ (.Y(_02566_),
    .A(net759),
    .B(net748));
 sg13g2_a22oi_1 _24234_ (.Y(_02567_),
    .B1(_02566_),
    .B2(net429),
    .A2(_02565_),
    .A1(net431));
 sg13g2_a21oi_1 _24235_ (.A1(net772),
    .A2(net750),
    .Y(_02568_),
    .B1(_01749_));
 sg13g2_or3_1 _24236_ (.A(net759),
    .B(net748),
    .C(_02568_),
    .X(_02569_));
 sg13g2_o21ai_1 _24237_ (.B1(_02569_),
    .Y(_02570_),
    .A1(net195),
    .A2(_02567_));
 sg13g2_nand2_1 _24238_ (.Y(_02571_),
    .A(net431),
    .B(_01770_));
 sg13g2_buf_1 _24239_ (.A(net748),
    .X(_02573_));
 sg13g2_nor3_1 _24240_ (.A(net195),
    .B(net419),
    .C(net409),
    .Y(_02574_));
 sg13g2_a22oi_1 _24241_ (.Y(_02575_),
    .B1(_02571_),
    .B2(_02574_),
    .A2(_02570_),
    .A1(net1078));
 sg13g2_xor2_1 _24242_ (.B(_02575_),
    .A(_02562_),
    .X(_02576_));
 sg13g2_nand2_1 _24243_ (.Y(_02577_),
    .A(net431),
    .B(_02565_));
 sg13g2_o21ai_1 _24244_ (.B1(_02577_),
    .Y(_02578_),
    .A1(_01685_),
    .A2(_02566_));
 sg13g2_nand2_1 _24245_ (.Y(_02579_),
    .A(net428),
    .B(_02578_));
 sg13g2_o21ai_1 _24246_ (.B1(_02579_),
    .Y(_02580_),
    .A1(net1078),
    .A2(_02566_));
 sg13g2_nor2_1 _24247_ (.A(_02551_),
    .B(_02037_),
    .Y(_02581_));
 sg13g2_and2_1 _24248_ (.A(_02139_),
    .B(_02558_),
    .X(_02582_));
 sg13g2_nor3_1 _24249_ (.A(net195),
    .B(_02566_),
    .C(_02571_),
    .Y(_02584_));
 sg13g2_a221oi_1 _24250_ (.B2(_02582_),
    .C1(_02584_),
    .B1(_02581_),
    .A1(net195),
    .Y(_02585_),
    .A2(_02580_));
 sg13g2_a21oi_1 _24251_ (.A1(_02576_),
    .A2(_02585_),
    .Y(_02586_),
    .B1(_05408_));
 sg13g2_xor2_1 _24252_ (.B(_02558_),
    .A(_02465_),
    .X(_02587_));
 sg13g2_a21oi_1 _24253_ (.A1(_04860_),
    .A2(_02587_),
    .Y(_02588_),
    .B1(net199));
 sg13g2_nand2_1 _24254_ (.Y(_02589_),
    .A(net1054),
    .B(_02435_));
 sg13g2_or3_1 _24255_ (.A(_02586_),
    .B(_02588_),
    .C(_02589_),
    .X(_02590_));
 sg13g2_o21ai_1 _24256_ (.B1(_02590_),
    .Y(_00496_),
    .A1(_06249_),
    .A2(_02435_));
 sg13g2_nand2_1 _24257_ (.Y(_02591_),
    .A(_01064_),
    .B(_02362_));
 sg13g2_buf_1 _24258_ (.A(_00039_),
    .X(_02592_));
 sg13g2_inv_1 _24259_ (.Y(_02594_),
    .A(_02592_));
 sg13g2_nor2_1 _24260_ (.A(_02594_),
    .B(net202),
    .Y(_02595_));
 sg13g2_buf_2 _24261_ (.A(\grid.cell_5_4.se ),
    .X(_02596_));
 sg13g2_inv_2 _24262_ (.Y(_02597_),
    .A(_02596_));
 sg13g2_xnor2_1 _24263_ (.Y(_02598_),
    .A(_02597_),
    .B(_02180_));
 sg13g2_xnor2_1 _24264_ (.Y(_02599_),
    .A(_01743_),
    .B(_02554_));
 sg13g2_xnor2_1 _24265_ (.Y(_02600_),
    .A(_02598_),
    .B(_02599_));
 sg13g2_xnor2_1 _24266_ (.Y(_02601_),
    .A(net420),
    .B(_02600_));
 sg13g2_a22oi_1 _24267_ (.Y(_02602_),
    .B1(_02600_),
    .B2(_02215_),
    .A2(net202),
    .A1(_02594_));
 sg13g2_o21ai_1 _24268_ (.B1(_02602_),
    .Y(_02603_),
    .A1(_02595_),
    .A2(_02601_));
 sg13g2_xor2_1 _24269_ (.B(_02596_),
    .A(_02177_),
    .X(_02605_));
 sg13g2_buf_1 _24270_ (.A(_02596_),
    .X(_02606_));
 sg13g2_nand2_1 _24271_ (.Y(_02607_),
    .A(net758),
    .B(net747));
 sg13g2_a22oi_1 _24272_ (.Y(_02608_),
    .B1(_02607_),
    .B2(_01808_),
    .A2(_02605_),
    .A1(net770));
 sg13g2_o21ai_1 _24273_ (.B1(net769),
    .Y(_02609_),
    .A1(_01750_),
    .A2(_02555_));
 sg13g2_nand3_1 _24274_ (.B(_02597_),
    .C(_02609_),
    .A(net198),
    .Y(_02610_));
 sg13g2_o21ai_1 _24275_ (.B1(_02610_),
    .Y(_02611_),
    .A1(net409),
    .A2(_02608_));
 sg13g2_nand2_1 _24276_ (.Y(_02612_),
    .A(net428),
    .B(_01812_));
 sg13g2_buf_1 _24277_ (.A(net747),
    .X(_02613_));
 sg13g2_nor3_1 _24278_ (.A(net409),
    .B(net418),
    .C(net408),
    .Y(_02614_));
 sg13g2_a22oi_1 _24279_ (.Y(_02616_),
    .B1(_02612_),
    .B2(_02614_),
    .A2(_02611_),
    .A1(_01852_));
 sg13g2_xor2_1 _24280_ (.B(_02616_),
    .A(_02603_),
    .X(_02617_));
 sg13g2_nand2_1 _24281_ (.Y(_02618_),
    .A(net770),
    .B(_02605_));
 sg13g2_o21ai_1 _24282_ (.B1(_02618_),
    .Y(_02619_),
    .A1(net770),
    .A2(_02607_));
 sg13g2_nand2_1 _24283_ (.Y(_02620_),
    .A(_01812_),
    .B(_02619_));
 sg13g2_o21ai_1 _24284_ (.B1(_02620_),
    .Y(_02621_),
    .A1(_01852_),
    .A2(_02607_));
 sg13g2_and2_1 _24285_ (.A(_02594_),
    .B(_02098_),
    .X(_02622_));
 sg13g2_and2_1 _24286_ (.A(_02215_),
    .B(_02600_),
    .X(_02623_));
 sg13g2_nor3_1 _24287_ (.A(net409),
    .B(_02607_),
    .C(_02612_),
    .Y(_02624_));
 sg13g2_a221oi_1 _24288_ (.B2(_02623_),
    .C1(_02624_),
    .B1(_02622_),
    .A1(net409),
    .Y(_02625_),
    .A2(_02621_));
 sg13g2_a21oi_1 _24289_ (.A1(_02617_),
    .A2(_02625_),
    .Y(_02627_),
    .B1(net97));
 sg13g2_xor2_1 _24290_ (.B(_02600_),
    .A(_02493_),
    .X(_02628_));
 sg13g2_a21oi_1 _24291_ (.A1(net70),
    .A2(_02628_),
    .Y(_02629_),
    .B1(net419));
 sg13g2_or3_1 _24292_ (.A(_02589_),
    .B(_02627_),
    .C(_02629_),
    .X(_02630_));
 sg13g2_o21ai_1 _24293_ (.B1(_02630_),
    .Y(_00497_),
    .A1(_12298_),
    .A2(_02591_));
 sg13g2_buf_1 _24294_ (.A(_00071_),
    .X(_02631_));
 sg13g2_nand2_1 _24295_ (.Y(_02632_),
    .A(_02631_),
    .B(_01750_));
 sg13g2_buf_2 _24296_ (.A(\grid.cell_5_5.se ),
    .X(_02633_));
 sg13g2_xnor2_1 _24297_ (.Y(_02634_),
    .A(_02596_),
    .B(_02633_));
 sg13g2_xnor2_1 _24298_ (.Y(_02635_),
    .A(_02227_),
    .B(_02634_));
 sg13g2_xnor2_1 _24299_ (.Y(_02637_),
    .A(net769),
    .B(_02635_));
 sg13g2_xnor2_1 _24300_ (.Y(_02638_),
    .A(net419),
    .B(_02637_));
 sg13g2_inv_1 _24301_ (.Y(_02639_),
    .A(_02631_));
 sg13g2_nand2_1 _24302_ (.Y(_02640_),
    .A(_02639_),
    .B(_01769_));
 sg13g2_o21ai_1 _24303_ (.B1(_02640_),
    .Y(_02641_),
    .A1(_02243_),
    .A2(_02637_));
 sg13g2_a21oi_1 _24304_ (.A1(_02632_),
    .A2(_02638_),
    .Y(_02642_),
    .B1(_02641_));
 sg13g2_xor2_1 _24305_ (.B(_02633_),
    .A(_02223_),
    .X(_02643_));
 sg13g2_buf_1 _24306_ (.A(_02633_),
    .X(_02644_));
 sg13g2_nand2_1 _24307_ (.Y(_02645_),
    .A(net757),
    .B(net746));
 sg13g2_a22oi_1 _24308_ (.Y(_02646_),
    .B1(_02645_),
    .B2(_01887_),
    .A2(_02643_),
    .A1(_01790_));
 sg13g2_nor2_1 _24309_ (.A(_02235_),
    .B(net746),
    .Y(_02648_));
 sg13g2_o21ai_1 _24310_ (.B1(net426),
    .Y(_02649_),
    .A1(_01808_),
    .A2(_02597_));
 sg13g2_nand2_1 _24311_ (.Y(_02650_),
    .A(_02648_),
    .B(_02649_));
 sg13g2_o21ai_1 _24312_ (.B1(_02650_),
    .Y(_02651_),
    .A1(net747),
    .A2(_02646_));
 sg13g2_nand2_1 _24313_ (.Y(_02652_),
    .A(net427),
    .B(net201));
 sg13g2_buf_1 _24314_ (.A(net746),
    .X(_02653_));
 sg13g2_buf_1 _24315_ (.A(net407),
    .X(_02654_));
 sg13g2_nor3_1 _24316_ (.A(net408),
    .B(net197),
    .C(net194),
    .Y(_02655_));
 sg13g2_a22oi_1 _24317_ (.Y(_02656_),
    .B1(_02652_),
    .B2(_02655_),
    .A2(_02651_),
    .A1(_01875_));
 sg13g2_xor2_1 _24318_ (.B(_02656_),
    .A(_02642_),
    .X(_02657_));
 sg13g2_nand2_1 _24319_ (.Y(_02659_),
    .A(_01790_),
    .B(_02643_));
 sg13g2_o21ai_1 _24320_ (.B1(_02659_),
    .Y(_02660_),
    .A1(net427),
    .A2(_02645_));
 sg13g2_nor2_1 _24321_ (.A(_01875_),
    .B(_02645_),
    .Y(_02661_));
 sg13g2_a21oi_1 _24322_ (.A1(net201),
    .A2(_02660_),
    .Y(_02662_),
    .B1(_02661_));
 sg13g2_nor2_1 _24323_ (.A(_02597_),
    .B(_02662_),
    .Y(_02663_));
 sg13g2_nor3_1 _24324_ (.A(net408),
    .B(_02645_),
    .C(_02652_),
    .Y(_02664_));
 sg13g2_nor4_1 _24325_ (.A(_02243_),
    .B(_02631_),
    .C(_02144_),
    .D(_02637_),
    .Y(_02665_));
 sg13g2_nor4_1 _24326_ (.A(_02657_),
    .B(_02663_),
    .C(_02664_),
    .D(_02665_),
    .Y(_02666_));
 sg13g2_xnor2_1 _24327_ (.Y(_02667_),
    .A(_02556_),
    .B(_02637_));
 sg13g2_a21oi_1 _24328_ (.A1(net114),
    .A2(_02667_),
    .Y(_02668_),
    .B1(net418));
 sg13g2_nor2_1 _24329_ (.A(_02589_),
    .B(_02668_),
    .Y(_02670_));
 sg13g2_o21ai_1 _24330_ (.B1(_02670_),
    .Y(_02671_),
    .A1(net81),
    .A2(_02666_));
 sg13g2_o21ai_1 _24331_ (.B1(_02671_),
    .Y(_00498_),
    .A1(net43),
    .A2(_02591_));
 sg13g2_buf_1 _24332_ (.A(_00133_),
    .X(_02672_));
 sg13g2_nor2_1 _24333_ (.A(net1072),
    .B(_02381_),
    .Y(_02673_));
 sg13g2_and3_1 _24334_ (.X(_02674_),
    .A(net1072),
    .B(net407),
    .C(_02381_));
 sg13g2_xnor2_1 _24335_ (.Y(_02675_),
    .A(net1072),
    .B(net407));
 sg13g2_nor2_1 _24336_ (.A(_02384_),
    .B(_02675_),
    .Y(_02676_));
 sg13g2_nor3_1 _24337_ (.A(_02673_),
    .B(_02674_),
    .C(_02676_),
    .Y(_02677_));
 sg13g2_inv_1 _24338_ (.Y(_02678_),
    .A(net746));
 sg13g2_buf_1 _24339_ (.A(_02678_),
    .X(_02680_));
 sg13g2_nand2_1 _24340_ (.Y(_02681_),
    .A(net193),
    .B(_02384_));
 sg13g2_a21oi_1 _24341_ (.A1(net200),
    .A2(net414),
    .Y(_02682_),
    .B1(net407));
 sg13g2_o21ai_1 _24342_ (.B1(net1072),
    .Y(_02683_),
    .A1(_02384_),
    .A2(_02682_));
 sg13g2_a21oi_1 _24343_ (.A1(_02681_),
    .A2(_02683_),
    .Y(_02684_),
    .B1(_01602_));
 sg13g2_buf_1 _24344_ (.A(net415),
    .X(_02685_));
 sg13g2_nand4_1 _24345_ (.B(net433),
    .C(net200),
    .A(net407),
    .Y(_02686_),
    .D(net192));
 sg13g2_a21oi_1 _24346_ (.A1(_02681_),
    .A2(_02686_),
    .Y(_02687_),
    .B1(net201));
 sg13g2_nor3_1 _24347_ (.A(_02672_),
    .B(net193),
    .C(_02381_),
    .Y(_02688_));
 sg13g2_nor3_1 _24348_ (.A(_02684_),
    .B(_02687_),
    .C(_02688_),
    .Y(_02689_));
 sg13g2_o21ai_1 _24349_ (.B1(_02689_),
    .Y(_02691_),
    .A1(_01914_),
    .A2(_02677_));
 sg13g2_buf_1 _24350_ (.A(_00103_),
    .X(_02692_));
 sg13g2_inv_1 _24351_ (.Y(_02693_),
    .A(_02692_));
 sg13g2_xnor2_1 _24352_ (.Y(_02694_),
    .A(_02633_),
    .B(_02368_));
 sg13g2_xor2_1 _24353_ (.B(_02694_),
    .A(_02007_),
    .X(_02695_));
 sg13g2_xnor2_1 _24354_ (.Y(_02696_),
    .A(_01822_),
    .B(_02695_));
 sg13g2_xnor2_1 _24355_ (.Y(_02697_),
    .A(net418),
    .B(_02696_));
 sg13g2_a21oi_1 _24356_ (.A1(_02692_),
    .A2(_01808_),
    .Y(_02698_),
    .B1(_02697_));
 sg13g2_a221oi_1 _24357_ (.B2(_02285_),
    .C1(_02698_),
    .B1(_02696_),
    .A1(_02693_),
    .Y(_02699_),
    .A2(net427));
 sg13g2_xor2_1 _24358_ (.B(_02699_),
    .A(_02691_),
    .X(_02700_));
 sg13g2_nand2_1 _24359_ (.Y(_02702_),
    .A(_01829_),
    .B(_02382_));
 sg13g2_o21ai_1 _24360_ (.B1(_02702_),
    .Y(_02703_),
    .A1(net201),
    .A2(_02381_));
 sg13g2_a21oi_1 _24361_ (.A1(net203),
    .A2(_02703_),
    .Y(_02704_),
    .B1(_02673_));
 sg13g2_nor2_1 _24362_ (.A(net193),
    .B(_02704_),
    .Y(_02705_));
 sg13g2_nor3_1 _24363_ (.A(net194),
    .B(_01914_),
    .C(_02381_),
    .Y(_02706_));
 sg13g2_nand2_1 _24364_ (.Y(_02707_),
    .A(_02285_),
    .B(_02696_));
 sg13g2_nor3_1 _24365_ (.A(_02692_),
    .B(_02180_),
    .C(_02707_),
    .Y(_02708_));
 sg13g2_nor4_1 _24366_ (.A(net125),
    .B(_02705_),
    .C(_02706_),
    .D(_02708_),
    .Y(_02709_));
 sg13g2_xnor2_1 _24367_ (.Y(_02710_),
    .A(_02598_),
    .B(_02696_));
 sg13g2_nand2_1 _24368_ (.Y(_02711_),
    .A(net756),
    .B(_02710_));
 sg13g2_nand3_1 _24369_ (.B(_02709_),
    .C(_02711_),
    .A(_02700_),
    .Y(_02713_));
 sg13g2_a22oi_1 _24370_ (.Y(_02714_),
    .B1(net25),
    .B2(_02360_),
    .A2(_07199_),
    .A1(net197));
 sg13g2_a221oi_1 _24371_ (.B2(_02714_),
    .C1(net557),
    .B1(_02713_),
    .A1(_06813_),
    .Y(_00499_),
    .A2(_02360_));
 sg13g2_nand2_1 _24372_ (.Y(_02715_),
    .A(_02633_),
    .B(net754));
 sg13g2_buf_2 _24373_ (.A(_02715_),
    .X(_02716_));
 sg13g2_o21ai_1 _24374_ (.B1(net757),
    .Y(_02717_),
    .A1(net746),
    .A2(net415));
 sg13g2_a21oi_1 _24375_ (.A1(_02716_),
    .A2(_02717_),
    .Y(_02718_),
    .B1(_01584_));
 sg13g2_nand2b_1 _24376_ (.Y(_02719_),
    .B(_02718_),
    .A_N(net1072));
 sg13g2_mux2_1 _24377_ (.A0(net407),
    .A1(_02716_),
    .S(_02235_),
    .X(_02720_));
 sg13g2_a22oi_1 _24378_ (.Y(_02721_),
    .B1(_02720_),
    .B2(net433),
    .A2(_02648_),
    .A1(net192));
 sg13g2_nand2b_1 _24379_ (.Y(_02723_),
    .B(net1072),
    .A_N(_02721_));
 sg13g2_nand3_1 _24380_ (.B(_02719_),
    .C(_02723_),
    .A(_01865_),
    .Y(_02724_));
 sg13g2_nand3_1 _24381_ (.B(net193),
    .C(_02369_),
    .A(net756),
    .Y(_02725_));
 sg13g2_nand4_1 _24382_ (.B(net194),
    .C(net433),
    .A(net197),
    .Y(_02726_),
    .D(net192));
 sg13g2_nand3_1 _24383_ (.B(_02725_),
    .C(_02726_),
    .A(_01887_),
    .Y(_02727_));
 sg13g2_nor2_1 _24384_ (.A(net1072),
    .B(_02716_),
    .Y(_02728_));
 sg13g2_nand3_1 _24385_ (.B(_02716_),
    .C(_02717_),
    .A(net1072),
    .Y(_02729_));
 sg13g2_a21oi_1 _24386_ (.A1(_02725_),
    .A2(_02729_),
    .Y(_02730_),
    .B1(_01602_));
 sg13g2_a221oi_1 _24387_ (.B2(net197),
    .C1(_02730_),
    .B1(_02728_),
    .A1(_02724_),
    .Y(_02731_),
    .A2(_02727_));
 sg13g2_inv_1 _24388_ (.Y(_02732_),
    .A(_01995_));
 sg13g2_xor2_1 _24389_ (.B(_02694_),
    .A(_02227_),
    .X(_02734_));
 sg13g2_xnor2_1 _24390_ (.Y(_02735_),
    .A(_01600_),
    .B(_02734_));
 sg13g2_xnor2_1 _24391_ (.Y(_02736_),
    .A(_02732_),
    .B(_02735_));
 sg13g2_inv_1 _24392_ (.Y(_02737_),
    .A(_02735_));
 sg13g2_o21ai_1 _24393_ (.B1(_02468_),
    .Y(_02738_),
    .A1(_01991_),
    .A2(_02737_));
 sg13g2_a21oi_1 _24394_ (.A1(_02463_),
    .A2(_02736_),
    .Y(_02739_),
    .B1(_02738_));
 sg13g2_xnor2_1 _24395_ (.Y(_02740_),
    .A(_02731_),
    .B(_02739_));
 sg13g2_nor2_1 _24396_ (.A(_02680_),
    .B(_02369_),
    .Y(_02741_));
 sg13g2_nor2_1 _24397_ (.A(_01887_),
    .B(_02694_),
    .Y(_02742_));
 sg13g2_a21oi_1 _24398_ (.A1(_01887_),
    .A2(_02741_),
    .Y(_02743_),
    .B1(_02742_));
 sg13g2_nor2_1 _24399_ (.A(_01584_),
    .B(_02743_),
    .Y(_02745_));
 sg13g2_o21ai_1 _24400_ (.B1(net197),
    .Y(_02746_),
    .A1(_02728_),
    .A2(_02745_));
 sg13g2_xor2_1 _24401_ (.B(_02735_),
    .A(_02484_),
    .X(_02747_));
 sg13g2_nor2_1 _24402_ (.A(net134),
    .B(_02747_),
    .Y(_02748_));
 sg13g2_nor4_1 _24403_ (.A(_02373_),
    .B(_01991_),
    .C(_02479_),
    .D(_02737_),
    .Y(_02749_));
 sg13g2_nor3_1 _24404_ (.A(net197),
    .B(_01914_),
    .C(_02716_),
    .Y(_02750_));
 sg13g2_nor4_1 _24405_ (.A(_06897_),
    .B(_02748_),
    .C(_02749_),
    .D(_02750_),
    .Y(_02751_));
 sg13g2_nand3_1 _24406_ (.B(_02746_),
    .C(_02751_),
    .A(_02740_),
    .Y(_02752_));
 sg13g2_a22oi_1 _24407_ (.Y(_02753_),
    .B1(net76),
    .B2(_02360_),
    .A2(_06817_),
    .A1(net134));
 sg13g2_o21ai_1 _24408_ (.B1(net435),
    .Y(_02754_),
    .A1(_11347_),
    .A2(_02361_));
 sg13g2_a21oi_1 _24409_ (.A1(_02752_),
    .A2(_02753_),
    .Y(_00500_),
    .B1(_02754_));
 sg13g2_nor3_1 _24410_ (.A(_02032_),
    .B(_05185_),
    .C(_09520_),
    .Y(_02756_));
 sg13g2_buf_1 _24411_ (.A(_02756_),
    .X(_02757_));
 sg13g2_buf_2 _24412_ (.A(\grid.cell_6_0.sw ),
    .X(_02758_));
 sg13g2_buf_1 _24413_ (.A(_02758_),
    .X(_02759_));
 sg13g2_buf_1 _24414_ (.A(_02759_),
    .X(_02760_));
 sg13g2_buf_1 _24415_ (.A(\grid.cell_6_0.se ),
    .X(_02761_));
 sg13g2_xnor2_1 _24416_ (.Y(_02762_),
    .A(_01952_),
    .B(_02761_));
 sg13g2_xor2_1 _24417_ (.B(_02762_),
    .A(_02382_),
    .X(_02763_));
 sg13g2_xnor2_1 _24418_ (.Y(_02764_),
    .A(net406),
    .B(_02763_));
 sg13g2_buf_1 _24419_ (.A(_02764_),
    .X(_02766_));
 sg13g2_xnor2_1 _24420_ (.Y(_02767_),
    .A(net416),
    .B(_02766_));
 sg13g2_nand2_1 _24421_ (.Y(_02768_),
    .A(net752),
    .B(_02767_));
 sg13g2_buf_2 _24422_ (.A(_00259_),
    .X(_02769_));
 sg13g2_inv_2 _24423_ (.Y(_02770_),
    .A(_02769_));
 sg13g2_a21oi_1 _24424_ (.A1(net755),
    .A2(_02521_),
    .Y(_02771_),
    .B1(_02732_));
 sg13g2_nor2_1 _24425_ (.A(net755),
    .B(_02521_),
    .Y(_02772_));
 sg13g2_mux2_1 _24426_ (.A0(net755),
    .A1(_02772_),
    .S(_02766_),
    .X(_02773_));
 sg13g2_nand2_1 _24427_ (.Y(_02774_),
    .A(net1076),
    .B(_01957_));
 sg13g2_nand2b_1 _24428_ (.Y(_02775_),
    .B(net745),
    .A_N(net1075));
 sg13g2_o21ai_1 _24429_ (.B1(_02775_),
    .Y(_02777_),
    .A1(net406),
    .A2(_02774_));
 sg13g2_or2_1 _24430_ (.X(_02778_),
    .B(net1075),
    .A(net745));
 sg13g2_nor2_1 _24431_ (.A(net754),
    .B(_02774_),
    .Y(_02779_));
 sg13g2_buf_1 _24432_ (.A(_02761_),
    .X(_02780_));
 sg13g2_inv_1 _24433_ (.Y(_02781_),
    .A(_02780_));
 sg13g2_buf_1 _24434_ (.A(_02781_),
    .X(_02782_));
 sg13g2_a221oi_1 _24435_ (.B2(_02779_),
    .C1(net191),
    .B1(_02778_),
    .A1(_02389_),
    .Y(_02783_),
    .A2(_02777_));
 sg13g2_nor2b_1 _24436_ (.A(net745),
    .B_N(_02107_),
    .Y(_02784_));
 sg13g2_a21o_1 _24437_ (.A2(_02775_),
    .A1(_02369_),
    .B1(_02784_),
    .X(_02785_));
 sg13g2_and2_1 _24438_ (.A(net745),
    .B(_02107_),
    .X(_02786_));
 sg13g2_a21o_1 _24439_ (.A2(_02778_),
    .A1(net754),
    .B1(_02786_),
    .X(_02788_));
 sg13g2_inv_1 _24440_ (.Y(_02789_),
    .A(_02774_));
 sg13g2_a221oi_1 _24441_ (.B2(_02789_),
    .C1(net744),
    .B1(_02788_),
    .A1(_02003_),
    .Y(_02790_),
    .A2(_02785_));
 sg13g2_nor2_1 _24442_ (.A(_02368_),
    .B(net745),
    .Y(_02791_));
 sg13g2_buf_2 _24443_ (.A(_02791_),
    .X(_02792_));
 sg13g2_and3_1 _24444_ (.X(_02793_),
    .A(_01955_),
    .B(_02368_),
    .C(_02758_));
 sg13g2_buf_1 _24445_ (.A(_02793_),
    .X(_02794_));
 sg13g2_mux2_1 _24446_ (.A0(_02792_),
    .A1(_02794_),
    .S(net744),
    .X(_02795_));
 sg13g2_a22oi_1 _24447_ (.Y(_02796_),
    .B1(_02784_),
    .B2(_02384_),
    .A2(_02795_),
    .A1(_01973_));
 sg13g2_o21ai_1 _24448_ (.B1(_02796_),
    .Y(_02797_),
    .A1(_02783_),
    .A2(_02790_));
 sg13g2_buf_1 _24449_ (.A(_02797_),
    .X(_02799_));
 sg13g2_o21ai_1 _24450_ (.B1(_02799_),
    .Y(_02800_),
    .A1(_02771_),
    .A2(_02773_));
 sg13g2_nand2_1 _24451_ (.Y(_02801_),
    .A(_02521_),
    .B(_02766_));
 sg13g2_and3_1 _24452_ (.X(_02802_),
    .A(_02769_),
    .B(_02799_),
    .C(_02801_));
 sg13g2_a21o_1 _24453_ (.A2(_02800_),
    .A1(_02770_),
    .B1(_02802_),
    .X(_02803_));
 sg13g2_nand2_1 _24454_ (.Y(_02804_),
    .A(net413),
    .B(_02766_));
 sg13g2_a21oi_1 _24455_ (.A1(net749),
    .A2(_02799_),
    .Y(_02805_),
    .B1(_02804_));
 sg13g2_nor3_1 _24456_ (.A(net413),
    .B(_02766_),
    .C(_02799_),
    .Y(_02806_));
 sg13g2_o21ai_1 _24457_ (.B1(_02732_),
    .Y(_02807_),
    .A1(_02805_),
    .A2(_02806_));
 sg13g2_nand3_1 _24458_ (.B(_02803_),
    .C(_02807_),
    .A(_02768_),
    .Y(_02808_));
 sg13g2_buf_1 _24459_ (.A(net744),
    .X(_02810_));
 sg13g2_nor2_1 _24460_ (.A(net423),
    .B(net405),
    .Y(_02811_));
 sg13g2_nand2_2 _24461_ (.Y(_02812_),
    .A(net415),
    .B(net406));
 sg13g2_xor2_1 _24462_ (.B(net745),
    .A(_02368_),
    .X(_02813_));
 sg13g2_and2_1 _24463_ (.A(net767),
    .B(_02813_),
    .X(_02814_));
 sg13g2_nor2_1 _24464_ (.A(net767),
    .B(_02812_),
    .Y(_02815_));
 sg13g2_o21ai_1 _24465_ (.B1(_01960_),
    .Y(_02816_),
    .A1(_02814_),
    .A2(_02815_));
 sg13g2_o21ai_1 _24466_ (.B1(_02816_),
    .Y(_02817_),
    .A1(net760),
    .A2(_02812_));
 sg13g2_a221oi_1 _24467_ (.B2(net405),
    .C1(_06244_),
    .B1(_02817_),
    .A1(_02811_),
    .Y(_02818_),
    .A2(_02794_));
 sg13g2_buf_1 _24468_ (.A(\grid.cell_6_0.s ),
    .X(_02819_));
 sg13g2_buf_1 _24469_ (.A(net1071),
    .X(_02821_));
 sg13g2_xor2_1 _24470_ (.B(net743),
    .A(net752),
    .X(_02822_));
 sg13g2_xnor2_1 _24471_ (.Y(_02823_),
    .A(_02767_),
    .B(_02822_));
 sg13g2_a21oi_1 _24472_ (.A1(_02768_),
    .A2(_02801_),
    .Y(_02824_),
    .B1(_02799_));
 sg13g2_a21oi_1 _24473_ (.A1(_02483_),
    .A2(_02823_),
    .Y(_02825_),
    .B1(_02824_));
 sg13g2_nand3_1 _24474_ (.B(_02818_),
    .C(_02825_),
    .A(_02808_),
    .Y(_02826_));
 sg13g2_a21oi_1 _24475_ (.A1(net753),
    .A2(_07561_),
    .Y(_02827_),
    .B1(net52));
 sg13g2_a221oi_1 _24476_ (.B2(_02827_),
    .C1(net557),
    .B1(_02826_),
    .A1(net50),
    .Y(_00501_),
    .A2(net52));
 sg13g2_nor2_1 _24477_ (.A(_05185_),
    .B(_09520_),
    .Y(_02828_));
 sg13g2_nand2_2 _24478_ (.Y(_02829_),
    .A(net108),
    .B(_02828_));
 sg13g2_buf_1 _24479_ (.A(\grid.cell_6_1.se ),
    .X(_02831_));
 sg13g2_buf_1 _24480_ (.A(net1070),
    .X(_02832_));
 sg13g2_nand2_1 _24481_ (.Y(_02833_),
    .A(net412),
    .B(net742));
 sg13g2_nand2_1 _24482_ (.Y(_02834_),
    .A(net1076),
    .B(_02022_));
 sg13g2_nor3_1 _24483_ (.A(net405),
    .B(_02833_),
    .C(_02834_),
    .Y(_02835_));
 sg13g2_xor2_1 _24484_ (.B(net742),
    .A(net751),
    .X(_02836_));
 sg13g2_nand2_1 _24485_ (.Y(_02837_),
    .A(net1076),
    .B(_02836_));
 sg13g2_o21ai_1 _24486_ (.B1(_02837_),
    .Y(_02838_),
    .A1(_01953_),
    .A2(_02833_));
 sg13g2_nor2b_1 _24487_ (.A(net1075),
    .B_N(net1070),
    .Y(_02839_));
 sg13g2_a22oi_1 _24488_ (.Y(_02840_),
    .B1(_02839_),
    .B2(_02459_),
    .A2(_02838_),
    .A1(net422));
 sg13g2_nor2_1 _24489_ (.A(net191),
    .B(_02840_),
    .Y(_02842_));
 sg13g2_xnor2_1 _24490_ (.Y(_02843_),
    .A(_01995_),
    .B(_02426_));
 sg13g2_inv_1 _24491_ (.Y(_02844_),
    .A(net1070));
 sg13g2_xnor2_1 _24492_ (.Y(_02845_),
    .A(_02844_),
    .B(_02473_));
 sg13g2_xnor2_1 _24493_ (.Y(_02846_),
    .A(_02762_),
    .B(_02845_));
 sg13g2_and4_1 _24494_ (.A(_02770_),
    .B(_02374_),
    .C(_02843_),
    .D(_02846_),
    .X(_02847_));
 sg13g2_or4_1 _24495_ (.A(_03821_),
    .B(_02835_),
    .C(_02842_),
    .D(_02847_),
    .X(_02848_));
 sg13g2_nor2_1 _24496_ (.A(_01995_),
    .B(_02770_),
    .Y(_02849_));
 sg13g2_xnor2_1 _24497_ (.Y(_02850_),
    .A(_02426_),
    .B(_02846_));
 sg13g2_a22oi_1 _24498_ (.Y(_02851_),
    .B1(_02374_),
    .B2(_02846_),
    .A2(_02770_),
    .A1(net752));
 sg13g2_o21ai_1 _24499_ (.B1(_02851_),
    .Y(_02853_),
    .A1(_02849_),
    .A2(_02850_));
 sg13g2_buf_1 _24500_ (.A(net742),
    .X(_02854_));
 sg13g2_nor2_1 _24501_ (.A(net412),
    .B(net404),
    .Y(_02855_));
 sg13g2_nor2_1 _24502_ (.A(_02038_),
    .B(_02394_),
    .Y(_02856_));
 sg13g2_nor2_1 _24503_ (.A(net742),
    .B(_02834_),
    .Y(_02857_));
 sg13g2_o21ai_1 _24504_ (.B1(net412),
    .Y(_02858_),
    .A1(_02839_),
    .A2(_02857_));
 sg13g2_nor2_1 _24505_ (.A(net412),
    .B(_02834_),
    .Y(_02859_));
 sg13g2_o21ai_1 _24506_ (.B1(_02859_),
    .Y(_02860_),
    .A1(net404),
    .A2(net1075));
 sg13g2_nand3_1 _24507_ (.B(_02858_),
    .C(_02860_),
    .A(net744),
    .Y(_02861_));
 sg13g2_nand2b_1 _24508_ (.Y(_02862_),
    .B(net1075),
    .A_N(net742));
 sg13g2_o21ai_1 _24509_ (.B1(_02862_),
    .Y(_02864_),
    .A1(net751),
    .A2(_02839_));
 sg13g2_nand2_1 _24510_ (.Y(_02865_),
    .A(net742),
    .B(net1075));
 sg13g2_o21ai_1 _24511_ (.B1(net751),
    .Y(_02866_),
    .A1(net1070),
    .A2(net1075));
 sg13g2_a21oi_1 _24512_ (.A1(_02865_),
    .A2(_02866_),
    .Y(_02867_),
    .B1(_02834_));
 sg13g2_a21oi_1 _24513_ (.A1(net763),
    .A2(_02864_),
    .Y(_02868_),
    .B1(_02867_));
 sg13g2_nand2_1 _24514_ (.Y(_02869_),
    .A(net191),
    .B(_02868_));
 sg13g2_nand2_1 _24515_ (.Y(_02870_),
    .A(net191),
    .B(_02855_));
 sg13g2_nand4_1 _24516_ (.B(net762),
    .C(net412),
    .A(net744),
    .Y(_02871_),
    .D(net404));
 sg13g2_a21oi_1 _24517_ (.A1(_02870_),
    .A2(_02871_),
    .Y(_02872_),
    .B1(_01953_));
 sg13g2_a221oi_1 _24518_ (.B2(_02869_),
    .C1(_02872_),
    .B1(_02861_),
    .A1(_02855_),
    .Y(_02873_),
    .A2(_02856_));
 sg13g2_xnor2_1 _24519_ (.Y(_02875_),
    .A(_02853_),
    .B(_02873_));
 sg13g2_xnor2_1 _24520_ (.Y(_02876_),
    .A(_02426_),
    .B(net1071));
 sg13g2_xnor2_1 _24521_ (.Y(_02877_),
    .A(_01995_),
    .B(_02876_));
 sg13g2_xnor2_1 _24522_ (.Y(_02878_),
    .A(_02846_),
    .B(_02877_));
 sg13g2_nor3_1 _24523_ (.A(_02848_),
    .B(_02875_),
    .C(_02878_),
    .Y(_02879_));
 sg13g2_o21ai_1 _24524_ (.B1(_02787_),
    .Y(_02880_),
    .A1(_02848_),
    .A2(_02875_));
 sg13g2_o21ai_1 _24525_ (.B1(_02880_),
    .Y(_02881_),
    .A1(net413),
    .A2(_02879_));
 sg13g2_o21ai_1 _24526_ (.B1(net435),
    .Y(_02882_),
    .A1(_11113_),
    .A2(_02829_));
 sg13g2_a21oi_1 _24527_ (.A1(_02829_),
    .A2(_02881_),
    .Y(_00502_),
    .B1(_02882_));
 sg13g2_nand2_1 _24528_ (.Y(_02883_),
    .A(_05812_),
    .B(net52));
 sg13g2_buf_1 _24529_ (.A(_00258_),
    .X(_02885_));
 sg13g2_buf_1 _24530_ (.A(_02885_),
    .X(_02886_));
 sg13g2_xor2_1 _24531_ (.B(net742),
    .A(_02022_),
    .X(_02887_));
 sg13g2_buf_2 _24532_ (.A(\grid.cell_6_2.se ),
    .X(_02888_));
 sg13g2_inv_1 _24533_ (.Y(_02889_),
    .A(_02888_));
 sg13g2_xnor2_1 _24534_ (.Y(_02890_),
    .A(net740),
    .B(_02503_));
 sg13g2_xnor2_1 _24535_ (.Y(_02891_),
    .A(_02887_),
    .B(_02890_));
 sg13g2_nor2_1 _24536_ (.A(net749),
    .B(_02891_),
    .Y(_02892_));
 sg13g2_xnor2_1 _24537_ (.Y(_02893_),
    .A(_02491_),
    .B(_02888_));
 sg13g2_xnor2_1 _24538_ (.Y(_02894_),
    .A(_02022_),
    .B(_02092_));
 sg13g2_xnor2_1 _24539_ (.Y(_02896_),
    .A(net1073),
    .B(net1070));
 sg13g2_xnor2_1 _24540_ (.Y(_02897_),
    .A(_02894_),
    .B(_02896_));
 sg13g2_xnor2_1 _24541_ (.Y(_02898_),
    .A(_02893_),
    .B(_02897_));
 sg13g2_buf_1 _24542_ (.A(_02898_),
    .X(_02899_));
 sg13g2_o21ai_1 _24543_ (.B1(_02899_),
    .Y(_02900_),
    .A1(net741),
    .A2(_02892_));
 sg13g2_nor2_1 _24544_ (.A(net741),
    .B(_02899_),
    .Y(_02901_));
 sg13g2_a21o_1 _24545_ (.A2(_02899_),
    .A1(_02010_),
    .B1(net741),
    .X(_02902_));
 sg13g2_mux2_1 _24546_ (.A0(_02901_),
    .A1(_02902_),
    .S(_02892_),
    .X(_02903_));
 sg13g2_a21o_1 _24547_ (.A2(_02900_),
    .A1(_01954_),
    .B1(_02903_),
    .X(_02904_));
 sg13g2_buf_1 _24548_ (.A(net404),
    .X(_02905_));
 sg13g2_nor2_1 _24549_ (.A(net763),
    .B(_02893_),
    .Y(_02907_));
 sg13g2_nand2_1 _24550_ (.Y(_02908_),
    .A(net750),
    .B(_02888_));
 sg13g2_nor2_1 _24551_ (.A(_02035_),
    .B(_02908_),
    .Y(_02909_));
 sg13g2_or2_1 _24552_ (.X(_02910_),
    .B(_02909_),
    .A(_02907_));
 sg13g2_nor2_1 _24553_ (.A(_02138_),
    .B(_02908_),
    .Y(_02911_));
 sg13g2_a21oi_1 _24554_ (.A1(_02152_),
    .A2(_02910_),
    .Y(_02912_),
    .B1(_02911_));
 sg13g2_nand2_1 _24555_ (.Y(_02913_),
    .A(net190),
    .B(_02912_));
 sg13g2_nand2_1 _24556_ (.Y(_02914_),
    .A(_02035_),
    .B(_02124_));
 sg13g2_buf_1 _24557_ (.A(_02844_),
    .X(_02915_));
 sg13g2_o21ai_1 _24558_ (.B1(_02915_),
    .Y(_02916_),
    .A1(_02914_),
    .A2(_02908_));
 sg13g2_nand2_1 _24559_ (.Y(_02918_),
    .A(net741),
    .B(_02899_));
 sg13g2_o21ai_1 _24560_ (.B1(_02010_),
    .Y(_02919_),
    .A1(net741),
    .A2(_02899_));
 sg13g2_a221oi_1 _24561_ (.B2(_02919_),
    .C1(_02892_),
    .B1(_02918_),
    .A1(_02913_),
    .Y(_02920_),
    .A2(_02916_));
 sg13g2_nand2_1 _24562_ (.Y(_02921_),
    .A(net421),
    .B(net190));
 sg13g2_buf_1 _24563_ (.A(_02888_),
    .X(_02922_));
 sg13g2_nor2_1 _24564_ (.A(net410),
    .B(net739),
    .Y(_02923_));
 sg13g2_nand2_1 _24565_ (.Y(_02924_),
    .A(_02138_),
    .B(_02923_));
 sg13g2_a21oi_1 _24566_ (.A1(_02152_),
    .A2(_02921_),
    .Y(_02925_),
    .B1(_02924_));
 sg13g2_nand2_1 _24567_ (.Y(_02926_),
    .A(_02923_),
    .B(_02914_));
 sg13g2_a21oi_1 _24568_ (.A1(net410),
    .A2(net739),
    .Y(_02927_),
    .B1(_02124_));
 sg13g2_o21ai_1 _24569_ (.B1(_02138_),
    .Y(_02929_),
    .A1(_02907_),
    .A2(_02927_));
 sg13g2_a21oi_1 _24570_ (.A1(_02926_),
    .A2(_02929_),
    .Y(_02930_),
    .B1(net190));
 sg13g2_nor2_1 _24571_ (.A(_02925_),
    .B(_02930_),
    .Y(_02931_));
 sg13g2_mux2_1 _24572_ (.A0(_02904_),
    .A1(_02920_),
    .S(_02931_),
    .X(_02932_));
 sg13g2_xor2_1 _24573_ (.B(_02899_),
    .A(_02762_),
    .X(_02933_));
 sg13g2_a21oi_1 _24574_ (.A1(_05415_),
    .A2(_02933_),
    .Y(_02934_),
    .B1(_02459_));
 sg13g2_nor2_1 _24575_ (.A(_02757_),
    .B(_02934_),
    .Y(_02935_));
 sg13g2_o21ai_1 _24576_ (.B1(_02935_),
    .Y(_02936_),
    .A1(net74),
    .A2(_02932_));
 sg13g2_a21oi_1 _24577_ (.A1(_02883_),
    .A2(_02936_),
    .Y(_00503_),
    .B1(_00661_));
 sg13g2_buf_1 _24578_ (.A(_00257_),
    .X(_02937_));
 sg13g2_buf_1 _24579_ (.A(\grid.cell_6_3.se ),
    .X(_02939_));
 sg13g2_xor2_1 _24580_ (.B(net1068),
    .A(_02142_),
    .X(_02940_));
 sg13g2_xnor2_1 _24581_ (.Y(_02941_),
    .A(_02888_),
    .B(_02554_));
 sg13g2_xnor2_1 _24582_ (.Y(_02942_),
    .A(_02940_),
    .B(_02941_));
 sg13g2_xnor2_1 _24583_ (.Y(_02943_),
    .A(net761),
    .B(_02942_));
 sg13g2_nor4_1 _24584_ (.A(net1069),
    .B(_02551_),
    .C(_02473_),
    .D(_02943_),
    .Y(_02944_));
 sg13g2_buf_1 _24585_ (.A(net739),
    .X(_02945_));
 sg13g2_nand2_2 _24586_ (.Y(_02946_),
    .A(_02564_),
    .B(net1068));
 sg13g2_xor2_1 _24587_ (.B(net1068),
    .A(_02554_),
    .X(_02947_));
 sg13g2_and2_1 _24588_ (.A(net420),
    .B(_02947_),
    .X(_02948_));
 sg13g2_a21oi_1 _24589_ (.A1(_02186_),
    .A2(_02946_),
    .Y(_02950_),
    .B1(_02948_));
 sg13g2_buf_1 _24590_ (.A(net1068),
    .X(_02951_));
 sg13g2_a21oi_1 _24591_ (.A1(net420),
    .A2(net739),
    .Y(_02952_),
    .B1(_02186_));
 sg13g2_or3_1 _24592_ (.A(_02564_),
    .B(net738),
    .C(_02952_),
    .X(_02953_));
 sg13g2_o21ai_1 _24593_ (.B1(_02953_),
    .Y(_02954_),
    .A1(net402),
    .A2(_02950_));
 sg13g2_nand2_1 _24594_ (.Y(_02955_),
    .A(net199),
    .B(_02159_));
 sg13g2_buf_1 _24595_ (.A(_02951_),
    .X(_02956_));
 sg13g2_nor3_1 _24596_ (.A(net402),
    .B(net409),
    .C(net401),
    .Y(_02957_));
 sg13g2_a22oi_1 _24597_ (.Y(_02958_),
    .B1(_02955_),
    .B2(_02957_),
    .A2(_02954_),
    .A1(_02193_));
 sg13g2_nand2_1 _24598_ (.Y(_02959_),
    .A(_02023_),
    .B(net1069));
 sg13g2_xnor2_1 _24599_ (.Y(_02960_),
    .A(net411),
    .B(_02943_));
 sg13g2_nand2b_1 _24600_ (.Y(_02961_),
    .B(_02038_),
    .A_N(net1069));
 sg13g2_o21ai_1 _24601_ (.B1(_02961_),
    .Y(_02962_),
    .A1(_02551_),
    .A2(_02943_));
 sg13g2_a21oi_1 _24602_ (.A1(_02959_),
    .A2(_02960_),
    .Y(_02963_),
    .B1(_02962_));
 sg13g2_xor2_1 _24603_ (.B(_02963_),
    .A(_02958_),
    .X(_02964_));
 sg13g2_nor2_1 _24604_ (.A(net199),
    .B(_02946_),
    .Y(_02965_));
 sg13g2_o21ai_1 _24605_ (.B1(_02159_),
    .Y(_02966_),
    .A1(_02948_),
    .A2(_02965_));
 sg13g2_nand2b_1 _24606_ (.Y(_02967_),
    .B(_02215_),
    .A_N(_02946_));
 sg13g2_a21oi_1 _24607_ (.A1(_02966_),
    .A2(_02967_),
    .Y(_02968_),
    .B1(net740));
 sg13g2_nor3_1 _24608_ (.A(net402),
    .B(_02946_),
    .C(_02955_),
    .Y(_02969_));
 sg13g2_nand2b_1 _24609_ (.Y(_02971_),
    .B(_01053_),
    .A_N(_02969_));
 sg13g2_nor4_1 _24610_ (.A(_02944_),
    .B(_02964_),
    .C(_02968_),
    .D(_02971_),
    .Y(_02972_));
 sg13g2_xnor2_1 _24611_ (.Y(_02973_),
    .A(_02845_),
    .B(_02943_));
 sg13g2_a21oi_1 _24612_ (.A1(_05517_),
    .A2(_02973_),
    .Y(_02974_),
    .B1(net195));
 sg13g2_nor2_1 _24613_ (.A(_02757_),
    .B(_02974_),
    .Y(_02975_));
 sg13g2_o21ai_1 _24614_ (.B1(_02975_),
    .Y(_02976_),
    .A1(_08877_),
    .A2(_02972_));
 sg13g2_o21ai_1 _24615_ (.B1(_02976_),
    .Y(_00504_),
    .A1(_06249_),
    .A2(_02829_));
 sg13g2_nand2_1 _24616_ (.Y(_02977_),
    .A(_07426_),
    .B(net52));
 sg13g2_buf_1 _24617_ (.A(\grid.cell_6_4.se ),
    .X(_02978_));
 sg13g2_inv_2 _24618_ (.Y(_02979_),
    .A(_02978_));
 sg13g2_xnor2_1 _24619_ (.Y(_02981_),
    .A(_02979_),
    .B(_02605_));
 sg13g2_xor2_1 _24620_ (.B(_02981_),
    .A(_02940_),
    .X(_02982_));
 sg13g2_inv_2 _24621_ (.Y(_02983_),
    .A(net750));
 sg13g2_xnor2_1 _24622_ (.Y(_02984_),
    .A(_02983_),
    .B(_02982_));
 sg13g2_buf_1 _24623_ (.A(_00038_),
    .X(_02985_));
 sg13g2_nand2b_1 _24624_ (.Y(_02986_),
    .B(net1066),
    .A_N(net420));
 sg13g2_nor2b_1 _24625_ (.A(net1066),
    .B_N(net199),
    .Y(_02987_));
 sg13g2_a221oi_1 _24626_ (.B2(_02986_),
    .C1(_02987_),
    .B1(_02984_),
    .A1(_02594_),
    .Y(_02988_),
    .A2(_02982_));
 sg13g2_xor2_1 _24627_ (.B(net1067),
    .A(_02596_),
    .X(_02989_));
 sg13g2_buf_1 _24628_ (.A(net1067),
    .X(_02990_));
 sg13g2_nand2_1 _24629_ (.Y(_02992_),
    .A(net747),
    .B(net737));
 sg13g2_a22oi_1 _24630_ (.Y(_02993_),
    .B1(_02992_),
    .B2(net198),
    .A2(_02989_),
    .A1(net759));
 sg13g2_a21oi_1 _24631_ (.A1(net759),
    .A2(net1068),
    .Y(_02994_),
    .B1(net198));
 sg13g2_or3_1 _24632_ (.A(net747),
    .B(net737),
    .C(_02994_),
    .X(_02995_));
 sg13g2_o21ai_1 _24633_ (.B1(_02995_),
    .Y(_02996_),
    .A1(net401),
    .A2(_02993_));
 sg13g2_nand2_1 _24634_ (.Y(_02997_),
    .A(net419),
    .B(net418));
 sg13g2_buf_1 _24635_ (.A(net737),
    .X(_02998_));
 sg13g2_nor3_1 _24636_ (.A(net401),
    .B(net747),
    .C(net400),
    .Y(_02999_));
 sg13g2_a22oi_1 _24637_ (.Y(_03000_),
    .B1(_02997_),
    .B2(_02999_),
    .A2(_02996_),
    .A1(_02243_));
 sg13g2_xnor2_1 _24638_ (.Y(_03001_),
    .A(_02988_),
    .B(_03000_));
 sg13g2_nand2_1 _24639_ (.Y(_03003_),
    .A(_02153_),
    .B(_02989_));
 sg13g2_o21ai_1 _24640_ (.B1(_03003_),
    .Y(_03004_),
    .A1(_02153_),
    .A2(_02992_));
 sg13g2_nand2_1 _24641_ (.Y(_03005_),
    .A(net418),
    .B(_03004_));
 sg13g2_o21ai_1 _24642_ (.B1(_03005_),
    .Y(_03006_),
    .A1(_02243_),
    .A2(_02992_));
 sg13g2_nor2_1 _24643_ (.A(net1066),
    .B(_02503_),
    .Y(_03007_));
 sg13g2_and2_1 _24644_ (.A(_02594_),
    .B(_02982_),
    .X(_03008_));
 sg13g2_nor3_1 _24645_ (.A(net401),
    .B(_02992_),
    .C(_02997_),
    .Y(_03009_));
 sg13g2_a221oi_1 _24646_ (.B2(_03008_),
    .C1(_03009_),
    .B1(_03007_),
    .A1(net401),
    .Y(_03010_),
    .A2(_03006_));
 sg13g2_a21oi_1 _24647_ (.A1(_03001_),
    .A2(_03010_),
    .Y(_03011_),
    .B1(_06897_));
 sg13g2_xor2_1 _24648_ (.B(_02982_),
    .A(_02890_),
    .X(_03012_));
 sg13g2_a21oi_1 _24649_ (.A1(_05619_),
    .A2(_03012_),
    .Y(_03014_),
    .B1(net409));
 sg13g2_or3_1 _24650_ (.A(net52),
    .B(_03011_),
    .C(_03014_),
    .X(_03015_));
 sg13g2_a21oi_1 _24651_ (.A1(_02977_),
    .A2(_03015_),
    .Y(_00505_),
    .B1(net440));
 sg13g2_buf_2 _24652_ (.A(\grid.cell_6_5.se ),
    .X(_03016_));
 sg13g2_buf_1 _24653_ (.A(_03016_),
    .X(_03017_));
 sg13g2_buf_1 _24654_ (.A(net736),
    .X(_03018_));
 sg13g2_nand2_2 _24655_ (.Y(_03019_),
    .A(net746),
    .B(net399));
 sg13g2_xor2_1 _24656_ (.B(_03016_),
    .A(_02633_),
    .X(_03020_));
 sg13g2_buf_2 _24657_ (.A(_03020_),
    .X(_03021_));
 sg13g2_nand2_1 _24658_ (.Y(_03022_),
    .A(_02190_),
    .B(_03021_));
 sg13g2_o21ai_1 _24659_ (.B1(_03022_),
    .Y(_03024_),
    .A1(_02190_),
    .A2(_03019_));
 sg13g2_nor2_1 _24660_ (.A(_02284_),
    .B(_03019_),
    .Y(_03025_));
 sg13g2_a21oi_1 _24661_ (.A1(net197),
    .A2(_03024_),
    .Y(_03026_),
    .B1(_03025_));
 sg13g2_nor2_1 _24662_ (.A(_02979_),
    .B(_03026_),
    .Y(_03027_));
 sg13g2_nand2_1 _24663_ (.Y(_03028_),
    .A(_02178_),
    .B(net417));
 sg13g2_nor3_1 _24664_ (.A(net400),
    .B(_03019_),
    .C(_03028_),
    .Y(_03029_));
 sg13g2_xor2_1 _24665_ (.B(net1067),
    .A(_02142_),
    .X(_03030_));
 sg13g2_xnor2_1 _24666_ (.Y(_03031_),
    .A(_02254_),
    .B(_03030_));
 sg13g2_xnor2_1 _24667_ (.Y(_03032_),
    .A(_03021_),
    .B(_03031_));
 sg13g2_xnor2_1 _24668_ (.Y(_03033_),
    .A(_02947_),
    .B(_03032_));
 sg13g2_a21oi_1 _24669_ (.A1(net127),
    .A2(_03033_),
    .Y(_03035_),
    .B1(net408));
 sg13g2_nor4_1 _24670_ (.A(net52),
    .B(_03027_),
    .C(_03029_),
    .D(_03035_),
    .Y(_03036_));
 sg13g2_buf_2 _24671_ (.A(_00070_),
    .X(_03037_));
 sg13g2_xnor2_1 _24672_ (.Y(_03038_),
    .A(_02555_),
    .B(_03032_));
 sg13g2_nor2_1 _24673_ (.A(_03037_),
    .B(_03038_),
    .Y(_03039_));
 sg13g2_xnor2_1 _24674_ (.Y(_03040_),
    .A(net1067),
    .B(_03016_));
 sg13g2_xor2_1 _24675_ (.B(_03040_),
    .A(_02643_),
    .X(_03041_));
 sg13g2_xnor2_1 _24676_ (.Y(_03042_),
    .A(net758),
    .B(_03041_));
 sg13g2_xnor2_1 _24677_ (.Y(_03043_),
    .A(_02555_),
    .B(_03042_));
 sg13g2_a22oi_1 _24678_ (.Y(_03044_),
    .B1(_03043_),
    .B2(net419),
    .A2(_03042_),
    .A1(_02639_));
 sg13g2_a22oi_1 _24679_ (.Y(_03046_),
    .B1(_03019_),
    .B2(net756),
    .A2(_03021_),
    .A1(_02178_));
 sg13g2_nor2_1 _24680_ (.A(_02633_),
    .B(net736),
    .Y(_03047_));
 sg13g2_o21ai_1 _24681_ (.B1(net417),
    .Y(_03048_),
    .A1(net198),
    .A2(_02979_));
 sg13g2_nand2_1 _24682_ (.Y(_03049_),
    .A(_03047_),
    .B(_03048_));
 sg13g2_o21ai_1 _24683_ (.B1(_03049_),
    .Y(_03050_),
    .A1(net400),
    .A2(_03046_));
 sg13g2_and2_1 _24684_ (.A(_03028_),
    .B(_03047_),
    .X(_03051_));
 sg13g2_a22oi_1 _24685_ (.Y(_03052_),
    .B1(_03051_),
    .B2(_02979_),
    .A2(_03050_),
    .A1(_02284_));
 sg13g2_xor2_1 _24686_ (.B(_03052_),
    .A(_03044_),
    .X(_03053_));
 sg13g2_nand3b_1 _24687_ (.B(_03044_),
    .C(_03039_),
    .Y(_03054_),
    .A_N(_03052_));
 sg13g2_o21ai_1 _24688_ (.B1(_03054_),
    .Y(_03055_),
    .A1(_03039_),
    .A2(_03053_));
 sg13g2_a21oi_1 _24689_ (.A1(net408),
    .A2(_05131_),
    .Y(_03057_),
    .B1(_02756_));
 sg13g2_a21oi_1 _24690_ (.A1(_05002_),
    .A2(net52),
    .Y(_03058_),
    .B1(_03057_));
 sg13g2_a21oi_1 _24691_ (.A1(_03036_),
    .A2(_03055_),
    .Y(_03059_),
    .B1(_03058_));
 sg13g2_nor2_1 _24692_ (.A(net214),
    .B(_03059_),
    .Y(_00506_));
 sg13g2_nand2_1 _24693_ (.Y(_03060_),
    .A(net194),
    .B(_07117_));
 sg13g2_inv_1 _24694_ (.Y(_03061_),
    .A(_03018_));
 sg13g2_nand2_1 _24695_ (.Y(_03062_),
    .A(_03061_),
    .B(_02792_));
 sg13g2_buf_1 _24696_ (.A(net406),
    .X(_03063_));
 sg13g2_buf_1 _24697_ (.A(_03018_),
    .X(_03064_));
 sg13g2_a21oi_1 _24698_ (.A1(net192),
    .A2(net189),
    .Y(_03065_),
    .B1(net188));
 sg13g2_buf_1 _24699_ (.A(_00132_),
    .X(_03067_));
 sg13g2_o21ai_1 _24700_ (.B1(net1065),
    .Y(_03068_),
    .A1(_02792_),
    .A2(_03065_));
 sg13g2_a21oi_1 _24701_ (.A1(_03062_),
    .A2(_03068_),
    .Y(_03069_),
    .B1(net134));
 sg13g2_nor2_1 _24702_ (.A(net1065),
    .B(_02812_),
    .Y(_03070_));
 sg13g2_and3_1 _24703_ (.X(_03071_),
    .A(net1065),
    .B(net399),
    .C(_02812_));
 sg13g2_xnor2_1 _24704_ (.Y(_03072_),
    .A(net1065),
    .B(net399));
 sg13g2_nor2_1 _24705_ (.A(_02792_),
    .B(_03072_),
    .Y(_03073_));
 sg13g2_nor3_1 _24706_ (.A(_03070_),
    .B(_03071_),
    .C(_03073_),
    .Y(_03074_));
 sg13g2_mux2_1 _24707_ (.A0(_02792_),
    .A1(_02794_),
    .S(net188),
    .X(_03075_));
 sg13g2_a22oi_1 _24708_ (.Y(_03076_),
    .B1(_03075_),
    .B2(net756),
    .A2(_03070_),
    .A1(net188));
 sg13g2_o21ai_1 _24709_ (.B1(_03076_),
    .Y(_03078_),
    .A1(_02310_),
    .A2(_03074_));
 sg13g2_nor2_1 _24710_ (.A(_03069_),
    .B(_03078_),
    .Y(_03079_));
 sg13g2_buf_2 _24711_ (.A(_00102_),
    .X(_03080_));
 sg13g2_xnor2_1 _24712_ (.Y(_03081_),
    .A(_03016_),
    .B(_02758_));
 sg13g2_xor2_1 _24713_ (.B(_03081_),
    .A(_02382_),
    .X(_03082_));
 sg13g2_xnor2_1 _24714_ (.Y(_03083_),
    .A(net757),
    .B(_03082_));
 sg13g2_xnor2_1 _24715_ (.Y(_03084_),
    .A(net408),
    .B(_03083_));
 sg13g2_a21oi_1 _24716_ (.A1(_03080_),
    .A2(_02185_),
    .Y(_03085_),
    .B1(_03084_));
 sg13g2_nand2_1 _24717_ (.Y(_03086_),
    .A(_02693_),
    .B(_03083_));
 sg13g2_o21ai_1 _24718_ (.B1(_03086_),
    .Y(_03087_),
    .A1(_03080_),
    .A2(_02185_));
 sg13g2_nor2_1 _24719_ (.A(_03085_),
    .B(_03087_),
    .Y(_03089_));
 sg13g2_xnor2_1 _24720_ (.Y(_03090_),
    .A(_03079_),
    .B(_03089_));
 sg13g2_buf_1 _24721_ (.A(_03064_),
    .X(_03091_));
 sg13g2_nand2_1 _24722_ (.Y(_03092_),
    .A(net417),
    .B(_02813_));
 sg13g2_o21ai_1 _24723_ (.B1(_03092_),
    .Y(_03093_),
    .A1(_02303_),
    .A2(_02812_));
 sg13g2_a21oi_1 _24724_ (.A1(net134),
    .A2(_03093_),
    .Y(_03094_),
    .B1(_03070_));
 sg13g2_a21oi_1 _24725_ (.A1(_02303_),
    .A2(_02794_),
    .Y(_03095_),
    .B1(net133));
 sg13g2_a21oi_1 _24726_ (.A1(net133),
    .A2(_03094_),
    .Y(_03096_),
    .B1(_03095_));
 sg13g2_nor3_1 _24727_ (.A(_03080_),
    .B(_02605_),
    .C(_03086_),
    .Y(_03097_));
 sg13g2_xor2_1 _24728_ (.B(_03083_),
    .A(_02981_),
    .X(_03098_));
 sg13g2_nor2_1 _24729_ (.A(net194),
    .B(_03098_),
    .Y(_03100_));
 sg13g2_nor4_1 _24730_ (.A(_03831_),
    .B(_03096_),
    .C(_03097_),
    .D(_03100_),
    .Y(_03101_));
 sg13g2_a22oi_1 _24731_ (.Y(_03102_),
    .B1(_03090_),
    .B2(_03101_),
    .A2(_02828_),
    .A1(_06810_));
 sg13g2_a221oi_1 _24732_ (.B2(_03102_),
    .C1(_08965_),
    .B1(_03060_),
    .A1(_06813_),
    .Y(_00507_),
    .A2(_02828_));
 sg13g2_xor2_1 _24733_ (.B(_03081_),
    .A(_02643_),
    .X(_03103_));
 sg13g2_xnor2_1 _24734_ (.Y(_03104_),
    .A(_01957_),
    .B(_03103_));
 sg13g2_buf_2 _24735_ (.A(_03104_),
    .X(_03105_));
 sg13g2_and2_1 _24736_ (.A(_02374_),
    .B(_03105_),
    .X(_03106_));
 sg13g2_buf_1 _24737_ (.A(_03106_),
    .X(_03107_));
 sg13g2_nand2_1 _24738_ (.Y(_03108_),
    .A(_03016_),
    .B(net745));
 sg13g2_buf_2 _24739_ (.A(_03108_),
    .X(_03110_));
 sg13g2_o21ai_1 _24740_ (.B1(net746),
    .Y(_03111_),
    .A1(net736),
    .A2(net406));
 sg13g2_a21o_1 _24741_ (.A2(_03111_),
    .A1(_03110_),
    .B1(_02003_),
    .X(_03112_));
 sg13g2_mux2_1 _24742_ (.A0(net399),
    .A1(_03110_),
    .S(_02644_),
    .X(_03113_));
 sg13g2_a22oi_1 _24743_ (.Y(_03114_),
    .B1(_03113_),
    .B2(net200),
    .A2(_03047_),
    .A1(net189));
 sg13g2_mux2_1 _24744_ (.A0(_03112_),
    .A1(_03114_),
    .S(net1065),
    .X(_03115_));
 sg13g2_nand2b_1 _24745_ (.Y(_03116_),
    .B(_03047_),
    .A_N(net189));
 sg13g2_nand4_1 _24746_ (.B(net399),
    .C(_01958_),
    .A(_02644_),
    .Y(_03117_),
    .D(net189));
 sg13g2_a21oi_1 _24747_ (.A1(_03116_),
    .A2(_03117_),
    .Y(_03118_),
    .B1(_02267_));
 sg13g2_nor3_1 _24748_ (.A(net1065),
    .B(net193),
    .C(_03110_),
    .Y(_03119_));
 sg13g2_nand3_1 _24749_ (.B(_03110_),
    .C(_03111_),
    .A(net1065),
    .Y(_03121_));
 sg13g2_a21oi_1 _24750_ (.A1(_03116_),
    .A2(_03121_),
    .Y(_03122_),
    .B1(_01960_));
 sg13g2_nor3_1 _24751_ (.A(_03118_),
    .B(_03119_),
    .C(_03122_),
    .Y(_03123_));
 sg13g2_o21ai_1 _24752_ (.B1(_03123_),
    .Y(_03124_),
    .A1(_02274_),
    .A2(_03115_));
 sg13g2_inv_1 _24753_ (.Y(_03125_),
    .A(_03124_));
 sg13g2_o21ai_1 _24754_ (.B1(_02769_),
    .Y(_03126_),
    .A1(_03107_),
    .A2(_03125_));
 sg13g2_nor2_1 _24755_ (.A(net753),
    .B(_02374_),
    .Y(_03127_));
 sg13g2_o21ai_1 _24756_ (.B1(_03105_),
    .Y(_03128_),
    .A1(net752),
    .A2(_02373_));
 sg13g2_a21oi_1 _24757_ (.A1(net753),
    .A2(_02374_),
    .Y(_03129_),
    .B1(_02732_));
 sg13g2_a221oi_1 _24758_ (.B2(net753),
    .C1(_03129_),
    .B1(_03128_),
    .A1(_03105_),
    .Y(_03130_),
    .A2(_03127_));
 sg13g2_or3_1 _24759_ (.A(_02769_),
    .B(_03125_),
    .C(_03130_),
    .X(_03132_));
 sg13g2_xnor2_1 _24760_ (.Y(_03133_),
    .A(_02483_),
    .B(_03105_));
 sg13g2_and2_1 _24761_ (.A(net752),
    .B(_03133_),
    .X(_03134_));
 sg13g2_buf_1 _24762_ (.A(_03134_),
    .X(_03135_));
 sg13g2_nor3_1 _24763_ (.A(net752),
    .B(_03133_),
    .C(_03124_),
    .Y(_03136_));
 sg13g2_nor2_1 _24764_ (.A(_03135_),
    .B(_03136_),
    .Y(_03137_));
 sg13g2_nand3_1 _24765_ (.B(_03132_),
    .C(_03137_),
    .A(_03126_),
    .Y(_03138_));
 sg13g2_buf_1 _24766_ (.A(_03063_),
    .X(_03139_));
 sg13g2_buf_1 _24767_ (.A(net132),
    .X(_03140_));
 sg13g2_nor3_1 _24768_ (.A(net194),
    .B(net133),
    .C(net95),
    .Y(_03141_));
 sg13g2_o21ai_1 _24769_ (.B1(_03141_),
    .Y(_03143_),
    .A1(_03135_),
    .A2(_03107_));
 sg13g2_nor2_1 _24770_ (.A(net95),
    .B(_03019_),
    .Y(_03144_));
 sg13g2_a21oi_1 _24771_ (.A1(net95),
    .A2(_03021_),
    .Y(_03145_),
    .B1(_03144_));
 sg13g2_a21oi_1 _24772_ (.A1(_03143_),
    .A2(_03145_),
    .Y(_03146_),
    .B1(_02310_));
 sg13g2_nor2_1 _24773_ (.A(_03135_),
    .B(_03107_),
    .Y(_03147_));
 sg13g2_o21ai_1 _24774_ (.B1(_03067_),
    .Y(_03148_),
    .A1(_02267_),
    .A2(_02003_));
 sg13g2_or2_1 _24775_ (.X(_03149_),
    .B(_03148_),
    .A(net132));
 sg13g2_and2_1 _24776_ (.A(net132),
    .B(_03148_),
    .X(_03150_));
 sg13g2_a21oi_1 _24777_ (.A1(net133),
    .A2(_03149_),
    .Y(_03151_),
    .B1(_03150_));
 sg13g2_xor2_1 _24778_ (.B(_03105_),
    .A(_02877_),
    .X(_03152_));
 sg13g2_a21oi_1 _24779_ (.A1(net172),
    .A2(_03152_),
    .Y(_03154_),
    .B1(net192));
 sg13g2_nor3_1 _24780_ (.A(_00648_),
    .B(_02756_),
    .C(_03154_),
    .Y(_03155_));
 sg13g2_o21ai_1 _24781_ (.B1(_03155_),
    .Y(_03156_),
    .A1(_03147_),
    .A2(_03151_));
 sg13g2_nor2_1 _24782_ (.A(_03091_),
    .B(_03149_),
    .Y(_03157_));
 sg13g2_a221oi_1 _24783_ (.B2(net133),
    .C1(_03107_),
    .B1(_03150_),
    .A1(_02429_),
    .Y(_03158_),
    .A2(_03133_));
 sg13g2_nor3_1 _24784_ (.A(net193),
    .B(_03157_),
    .C(_03158_),
    .Y(_03159_));
 sg13g2_nor3_1 _24785_ (.A(_03146_),
    .B(_03156_),
    .C(_03159_),
    .Y(_03160_));
 sg13g2_nand2_1 _24786_ (.Y(_03161_),
    .A(net80),
    .B(net52));
 sg13g2_nand3_1 _24787_ (.B(_05471_),
    .C(_02829_),
    .A(net192),
    .Y(_03162_));
 sg13g2_a21oi_1 _24788_ (.A1(_03161_),
    .A2(_03162_),
    .Y(_03163_),
    .B1(_00669_));
 sg13g2_a21o_1 _24789_ (.A2(_03160_),
    .A1(_03138_),
    .B1(_03163_),
    .X(_00508_));
 sg13g2_xnor2_1 _24790_ (.Y(_03165_),
    .A(net1073),
    .B(_02379_));
 sg13g2_buf_1 _24791_ (.A(\grid.cell_7_0.sw ),
    .X(_03166_));
 sg13g2_xor2_1 _24792_ (.B(_03166_),
    .A(_02758_),
    .X(_03167_));
 sg13g2_buf_2 _24793_ (.A(\grid.cell_7_0.se ),
    .X(_03168_));
 sg13g2_xnor2_1 _24794_ (.Y(_03169_),
    .A(_02761_),
    .B(_03168_));
 sg13g2_xor2_1 _24795_ (.B(_03169_),
    .A(_03167_),
    .X(_03170_));
 sg13g2_xnor2_1 _24796_ (.Y(_03171_),
    .A(_03165_),
    .B(_03170_));
 sg13g2_buf_2 _24797_ (.A(_03171_),
    .X(_03172_));
 sg13g2_buf_1 _24798_ (.A(\grid.cell_7_0.s ),
    .X(_03173_));
 sg13g2_buf_1 _24799_ (.A(_03173_),
    .X(_03175_));
 sg13g2_buf_1 _24800_ (.A(net735),
    .X(_03176_));
 sg13g2_xor2_1 _24801_ (.B(net398),
    .A(_02427_),
    .X(_03177_));
 sg13g2_xnor2_1 _24802_ (.Y(_03178_),
    .A(_03172_),
    .B(_03177_));
 sg13g2_a21oi_1 _24803_ (.A1(net78),
    .A2(_03178_),
    .Y(_03179_),
    .B1(net743));
 sg13g2_nor2_2 _24804_ (.A(_05750_),
    .B(_09520_),
    .Y(_03180_));
 sg13g2_nand2_1 _24805_ (.Y(_03181_),
    .A(net327),
    .B(_03180_));
 sg13g2_buf_2 _24806_ (.A(_03181_),
    .X(_03182_));
 sg13g2_buf_1 _24807_ (.A(_00254_),
    .X(_03183_));
 sg13g2_buf_1 _24808_ (.A(_03183_),
    .X(_03184_));
 sg13g2_buf_1 _24809_ (.A(_03166_),
    .X(_03186_));
 sg13g2_buf_1 _24810_ (.A(_03186_),
    .X(_03187_));
 sg13g2_xnor2_1 _24811_ (.Y(_03188_),
    .A(net1073),
    .B(_03168_));
 sg13g2_xnor2_1 _24812_ (.Y(_03189_),
    .A(net397),
    .B(_03188_));
 sg13g2_xnor2_1 _24813_ (.Y(_03190_),
    .A(_02813_),
    .B(_03189_));
 sg13g2_nor2_1 _24814_ (.A(net741),
    .B(_03190_),
    .Y(_03191_));
 sg13g2_o21ai_1 _24815_ (.B1(_03172_),
    .Y(_03192_),
    .A1(net734),
    .A2(_03191_));
 sg13g2_nor2_1 _24816_ (.A(net734),
    .B(_03172_),
    .Y(_03193_));
 sg13g2_a21o_1 _24817_ (.A2(_03172_),
    .A1(_02483_),
    .B1(_03183_),
    .X(_03194_));
 sg13g2_mux2_1 _24818_ (.A0(_03193_),
    .A1(_03194_),
    .S(_03191_),
    .X(_03195_));
 sg13g2_a21o_1 _24819_ (.A2(_03192_),
    .A1(net753),
    .B1(_03195_),
    .X(_03197_));
 sg13g2_nand2_1 _24820_ (.Y(_03198_),
    .A(net734),
    .B(_03172_));
 sg13g2_o21ai_1 _24821_ (.B1(_02483_),
    .Y(_03199_),
    .A1(net734),
    .A2(_03172_));
 sg13g2_a21oi_1 _24822_ (.A1(_03198_),
    .A2(_03199_),
    .Y(_03200_),
    .B1(_03191_));
 sg13g2_buf_1 _24823_ (.A(_03168_),
    .X(_03201_));
 sg13g2_buf_1 _24824_ (.A(net732),
    .X(_03202_));
 sg13g2_inv_1 _24825_ (.Y(_03203_),
    .A(net397));
 sg13g2_nand2_1 _24826_ (.Y(_03204_),
    .A(net755),
    .B(_02400_));
 sg13g2_a21o_1 _24827_ (.A2(_02521_),
    .A1(_03203_),
    .B1(_03204_),
    .X(_03205_));
 sg13g2_nor2b_1 _24828_ (.A(_02512_),
    .B_N(net397),
    .Y(_03206_));
 sg13g2_buf_1 _24829_ (.A(net397),
    .X(_03208_));
 sg13g2_nor2_1 _24830_ (.A(net187),
    .B(_03204_),
    .Y(_03209_));
 sg13g2_o21ai_1 _24831_ (.B1(net132),
    .Y(_03210_),
    .A1(_03206_),
    .A2(_03209_));
 sg13g2_o21ai_1 _24832_ (.B1(_03210_),
    .Y(_03211_),
    .A1(net132),
    .A2(_03205_));
 sg13g2_nor2_1 _24833_ (.A(net397),
    .B(_02521_),
    .Y(_03212_));
 sg13g2_nor2_1 _24834_ (.A(net189),
    .B(_03206_),
    .Y(_03213_));
 sg13g2_or2_1 _24835_ (.X(_03214_),
    .B(_03213_),
    .A(_03212_));
 sg13g2_nand2_1 _24836_ (.Y(_03215_),
    .A(net187),
    .B(net749));
 sg13g2_o21ai_1 _24837_ (.B1(net189),
    .Y(_03216_),
    .A1(net187),
    .A2(net749));
 sg13g2_a21oi_1 _24838_ (.A1(_03215_),
    .A2(_03216_),
    .Y(_03217_),
    .B1(_03204_));
 sg13g2_a21oi_1 _24839_ (.A1(_02369_),
    .A2(_03214_),
    .Y(_03219_),
    .B1(_03217_));
 sg13g2_or2_1 _24840_ (.X(_03220_),
    .B(net733),
    .A(net406));
 sg13g2_buf_1 _24841_ (.A(_03220_),
    .X(_03221_));
 sg13g2_and2_1 _24842_ (.A(net406),
    .B(_03186_),
    .X(_03222_));
 sg13g2_buf_1 _24843_ (.A(_03222_),
    .X(_03223_));
 sg13g2_nand3_1 _24844_ (.B(net414),
    .C(_03223_),
    .A(net732),
    .Y(_03224_));
 sg13g2_o21ai_1 _24845_ (.B1(_03224_),
    .Y(_03225_),
    .A1(net732),
    .A2(_03221_));
 sg13g2_a22oi_1 _24846_ (.Y(_03226_),
    .B1(_03225_),
    .B2(net416),
    .A2(_03212_),
    .A1(_02792_));
 sg13g2_o21ai_1 _24847_ (.B1(_03226_),
    .Y(_03227_),
    .A1(net396),
    .A2(_03219_));
 sg13g2_a21oi_1 _24848_ (.A1(net396),
    .A2(_03211_),
    .Y(_03228_),
    .B1(_03227_));
 sg13g2_mux2_1 _24849_ (.A0(_03197_),
    .A1(_03200_),
    .S(_03228_),
    .X(_03230_));
 sg13g2_inv_1 _24850_ (.Y(_03231_),
    .A(_03168_));
 sg13g2_buf_1 _24851_ (.A(_03231_),
    .X(_03232_));
 sg13g2_nand2_2 _24852_ (.Y(_03233_),
    .A(net406),
    .B(net397));
 sg13g2_nand2_1 _24853_ (.Y(_03234_),
    .A(_02407_),
    .B(_03167_));
 sg13g2_o21ai_1 _24854_ (.B1(_03234_),
    .Y(_03235_),
    .A1(net413),
    .A2(_03233_));
 sg13g2_a22oi_1 _24855_ (.Y(_03236_),
    .B1(_03235_),
    .B2(net192),
    .A2(_03206_),
    .A1(net95));
 sg13g2_nor2_1 _24856_ (.A(net395),
    .B(_03236_),
    .Y(_03237_));
 sg13g2_nor3_1 _24857_ (.A(net396),
    .B(_03233_),
    .C(_03204_),
    .Y(_03238_));
 sg13g2_nand2_1 _24858_ (.Y(_03239_),
    .A(net1194),
    .B(_03182_));
 sg13g2_nor3_1 _24859_ (.A(_03237_),
    .B(_03238_),
    .C(_03239_),
    .Y(_03241_));
 sg13g2_a22oi_1 _24860_ (.Y(_03242_),
    .B1(_03230_),
    .B2(_03241_),
    .A2(_03182_),
    .A1(_08877_));
 sg13g2_inv_1 _24861_ (.Y(_03243_),
    .A(_03180_));
 sg13g2_nor2_1 _24862_ (.A(_02043_),
    .B(_03243_),
    .Y(_03244_));
 sg13g2_nand3_1 _24863_ (.B(net44),
    .C(_03244_),
    .A(_06118_),
    .Y(_03245_));
 sg13g2_o21ai_1 _24864_ (.B1(_03245_),
    .Y(_00509_),
    .A1(_03179_),
    .A2(_03242_));
 sg13g2_buf_2 _24865_ (.A(\grid.cell_7_1.se ),
    .X(_03246_));
 sg13g2_xnor2_1 _24866_ (.Y(_03247_),
    .A(net1070),
    .B(_03246_));
 sg13g2_buf_1 _24867_ (.A(_03246_),
    .X(_03248_));
 sg13g2_buf_1 _24868_ (.A(net731),
    .X(_03249_));
 sg13g2_a21oi_1 _24869_ (.A1(net404),
    .A2(net394),
    .Y(_03251_),
    .B1(net755));
 sg13g2_a21oi_1 _24870_ (.A1(net755),
    .A2(_03247_),
    .Y(_03252_),
    .B1(_03251_));
 sg13g2_nor2b_1 _24871_ (.A(_02512_),
    .B_N(_03246_),
    .Y(_03253_));
 sg13g2_a22oi_1 _24872_ (.Y(_03254_),
    .B1(_03253_),
    .B2(_02905_),
    .A2(_03252_),
    .A1(net411));
 sg13g2_nor2_1 _24873_ (.A(net395),
    .B(_03254_),
    .Y(_03255_));
 sg13g2_inv_1 _24874_ (.Y(_03256_),
    .A(net394));
 sg13g2_nor4_1 _24875_ (.A(_02378_),
    .B(net396),
    .C(_03256_),
    .D(_02833_),
    .Y(_03257_));
 sg13g2_xnor2_1 _24876_ (.Y(_03258_),
    .A(_02436_),
    .B(_03246_));
 sg13g2_xnor2_1 _24877_ (.Y(_03259_),
    .A(_02896_),
    .B(_03258_));
 sg13g2_xnor2_1 _24878_ (.Y(_03260_),
    .A(_03231_),
    .B(_03259_));
 sg13g2_inv_1 _24879_ (.Y(_03262_),
    .A(_03183_));
 sg13g2_nand2_1 _24880_ (.Y(_03263_),
    .A(net730),
    .B(_02876_));
 sg13g2_nor3_1 _24881_ (.A(_02769_),
    .B(_03260_),
    .C(_03263_),
    .Y(_03264_));
 sg13g2_or4_1 _24882_ (.A(net368),
    .B(_03255_),
    .C(_03257_),
    .D(_03264_),
    .X(_03265_));
 sg13g2_nand2_1 _24883_ (.Y(_03266_),
    .A(_02483_),
    .B(net734));
 sg13g2_xnor2_1 _24884_ (.Y(_03267_),
    .A(net1071),
    .B(_03260_));
 sg13g2_nand2_1 _24885_ (.Y(_03268_),
    .A(_02426_),
    .B(net730));
 sg13g2_o21ai_1 _24886_ (.B1(_03268_),
    .Y(_03269_),
    .A1(_02769_),
    .A2(_03260_));
 sg13g2_a21oi_1 _24887_ (.A1(_03266_),
    .A2(_03267_),
    .Y(_03270_),
    .B1(_03269_));
 sg13g2_buf_1 _24888_ (.A(_03249_),
    .X(_03271_));
 sg13g2_nor2_1 _24889_ (.A(net186),
    .B(_02521_),
    .Y(_03273_));
 sg13g2_nand2_1 _24890_ (.Y(_03274_),
    .A(_02364_),
    .B(_02437_));
 sg13g2_nor2_1 _24891_ (.A(net731),
    .B(_03274_),
    .Y(_03275_));
 sg13g2_o21ai_1 _24892_ (.B1(_02854_),
    .Y(_03276_),
    .A1(_03253_),
    .A2(_03275_));
 sg13g2_nor2_1 _24893_ (.A(_02854_),
    .B(_03274_),
    .Y(_03277_));
 sg13g2_o21ai_1 _24894_ (.B1(_03277_),
    .Y(_03278_),
    .A1(net394),
    .A2(_02513_));
 sg13g2_nand3_1 _24895_ (.B(_03276_),
    .C(_03278_),
    .A(net732),
    .Y(_03279_));
 sg13g2_nand2b_1 _24896_ (.Y(_03280_),
    .B(_02512_),
    .A_N(net731));
 sg13g2_o21ai_1 _24897_ (.B1(_03280_),
    .Y(_03281_),
    .A1(_02832_),
    .A2(_03253_));
 sg13g2_nand2_1 _24898_ (.Y(_03282_),
    .A(net731),
    .B(_02513_));
 sg13g2_o21ai_1 _24899_ (.B1(_02832_),
    .Y(_03284_),
    .A1(net731),
    .A2(_02512_));
 sg13g2_a21oi_1 _24900_ (.A1(_03282_),
    .A2(_03284_),
    .Y(_03285_),
    .B1(_03274_));
 sg13g2_a21oi_1 _24901_ (.A1(_02457_),
    .A2(_03281_),
    .Y(_03286_),
    .B1(_03285_));
 sg13g2_nand2_1 _24902_ (.Y(_03287_),
    .A(net395),
    .B(_03286_));
 sg13g2_nand3_1 _24903_ (.B(net403),
    .C(_03256_),
    .A(net395),
    .Y(_03288_));
 sg13g2_nand4_1 _24904_ (.B(_02438_),
    .C(net404),
    .A(net732),
    .Y(_03289_),
    .D(net394));
 sg13g2_a21oi_1 _24905_ (.A1(_03288_),
    .A2(_03289_),
    .Y(_03290_),
    .B1(_02376_));
 sg13g2_a221oi_1 _24906_ (.B2(_03287_),
    .C1(_03290_),
    .B1(_03279_),
    .A1(_02855_),
    .Y(_03291_),
    .A2(_03273_));
 sg13g2_xor2_1 _24907_ (.B(_03291_),
    .A(_03270_),
    .X(_03292_));
 sg13g2_xnor2_1 _24908_ (.Y(_03293_),
    .A(net735),
    .B(_02876_));
 sg13g2_xor2_1 _24909_ (.B(_03293_),
    .A(_03260_),
    .X(_03295_));
 sg13g2_nor3_1 _24910_ (.A(_03265_),
    .B(_03292_),
    .C(_03295_),
    .Y(_03296_));
 sg13g2_o21ai_1 _24911_ (.B1(net85),
    .Y(_03297_),
    .A1(_03265_),
    .A2(_03292_));
 sg13g2_o21ai_1 _24912_ (.B1(_03297_),
    .Y(_03298_),
    .A1(net405),
    .A2(_03296_));
 sg13g2_o21ai_1 _24913_ (.B1(net435),
    .Y(_03299_),
    .A1(net38),
    .A2(_03182_));
 sg13g2_a21oi_1 _24914_ (.A1(_03182_),
    .A2(_03298_),
    .Y(_00510_),
    .B1(_03299_));
 sg13g2_buf_2 _24915_ (.A(\grid.cell_7_2.se ),
    .X(_03300_));
 sg13g2_buf_1 _24916_ (.A(_03300_),
    .X(_03301_));
 sg13g2_nand2_2 _24917_ (.Y(_03302_),
    .A(net739),
    .B(net729));
 sg13g2_xor2_1 _24918_ (.B(net729),
    .A(_02888_),
    .X(_03303_));
 sg13g2_nand2_1 _24919_ (.Y(_03305_),
    .A(net196),
    .B(_03303_));
 sg13g2_o21ai_1 _24920_ (.B1(_03305_),
    .Y(_03306_),
    .A1(net196),
    .A2(_03302_));
 sg13g2_nor2_1 _24921_ (.A(_02551_),
    .B(_03302_),
    .Y(_03307_));
 sg13g2_a21oi_1 _24922_ (.A1(_02563_),
    .A2(_03306_),
    .Y(_03308_),
    .B1(_03307_));
 sg13g2_nor2_1 _24923_ (.A(_03256_),
    .B(_03308_),
    .Y(_03309_));
 sg13g2_nand2_1 _24924_ (.Y(_03310_),
    .A(_02438_),
    .B(_02501_));
 sg13g2_nor3_1 _24925_ (.A(net186),
    .B(_03302_),
    .C(_03310_),
    .Y(_03311_));
 sg13g2_xnor2_1 _24926_ (.Y(_03312_),
    .A(_02888_),
    .B(_03300_));
 sg13g2_xnor2_1 _24927_ (.Y(_03313_),
    .A(_02364_),
    .B(_02492_));
 sg13g2_xnor2_1 _24928_ (.Y(_03314_),
    .A(_03258_),
    .B(_03313_));
 sg13g2_xnor2_1 _24929_ (.Y(_03316_),
    .A(_03312_),
    .B(_03314_));
 sg13g2_xor2_1 _24930_ (.B(_03316_),
    .A(_03169_),
    .X(_03317_));
 sg13g2_a21oi_1 _24931_ (.A1(_02776_),
    .A2(_03317_),
    .Y(_03318_),
    .B1(net190));
 sg13g2_nor4_1 _24932_ (.A(_03244_),
    .B(_03309_),
    .C(_03311_),
    .D(_03318_),
    .Y(_03319_));
 sg13g2_a22oi_1 _24933_ (.Y(_03320_),
    .B1(_03302_),
    .B2(_02983_),
    .A2(_03303_),
    .A1(net411));
 sg13g2_nor2_1 _24934_ (.A(_02922_),
    .B(net729),
    .Y(_03321_));
 sg13g2_nand2_1 _24935_ (.Y(_03322_),
    .A(_03310_),
    .B(_03321_));
 sg13g2_o21ai_1 _24936_ (.B1(_03322_),
    .Y(_03323_),
    .A1(_02552_),
    .A2(_03320_));
 sg13g2_buf_1 _24937_ (.A(net729),
    .X(_03324_));
 sg13g2_a21oi_1 _24938_ (.A1(_02441_),
    .A2(net394),
    .Y(_03325_),
    .B1(_02983_));
 sg13g2_nor4_1 _24939_ (.A(net402),
    .B(net393),
    .C(_02552_),
    .D(_03325_),
    .Y(_03327_));
 sg13g2_a21oi_1 _24940_ (.A1(_03256_),
    .A2(_03323_),
    .Y(_03328_),
    .B1(_03327_));
 sg13g2_inv_2 _24941_ (.Y(_03329_),
    .A(_02885_));
 sg13g2_xnor2_1 _24942_ (.Y(_03330_),
    .A(_03300_),
    .B(_02893_));
 sg13g2_xnor2_1 _24943_ (.Y(_03331_),
    .A(_03258_),
    .B(_03330_));
 sg13g2_xnor2_1 _24944_ (.Y(_03332_),
    .A(net191),
    .B(_03331_));
 sg13g2_a22oi_1 _24945_ (.Y(_03333_),
    .B1(_03332_),
    .B2(_02407_),
    .A2(_03331_),
    .A1(_03329_));
 sg13g2_nor2b_1 _24946_ (.A(_03328_),
    .B_N(_03333_),
    .Y(_03334_));
 sg13g2_xnor2_1 _24947_ (.Y(_03335_),
    .A(_03333_),
    .B(_03328_));
 sg13g2_buf_1 _24948_ (.A(_00256_),
    .X(_03336_));
 sg13g2_inv_1 _24949_ (.Y(_03338_),
    .A(_03336_));
 sg13g2_xnor2_1 _24950_ (.Y(_03339_),
    .A(net405),
    .B(_03316_));
 sg13g2_nand2_1 _24951_ (.Y(_03340_),
    .A(_03338_),
    .B(_03339_));
 sg13g2_mux2_1 _24952_ (.A0(_03334_),
    .A1(_03335_),
    .S(_03340_),
    .X(_03341_));
 sg13g2_nand3_1 _24953_ (.B(_07553_),
    .C(_03182_),
    .A(net190),
    .Y(_03342_));
 sg13g2_o21ai_1 _24954_ (.B1(_03342_),
    .Y(_03343_),
    .A1(_04077_),
    .A2(_03182_));
 sg13g2_a21oi_1 _24955_ (.A1(_03319_),
    .A2(_03341_),
    .Y(_03344_),
    .B1(_03343_));
 sg13g2_nor2_1 _24956_ (.A(net214),
    .B(_03344_),
    .Y(_00511_));
 sg13g2_buf_1 _24957_ (.A(_00255_),
    .X(_03345_));
 sg13g2_nand2b_1 _24958_ (.Y(_03346_),
    .B(net190),
    .A_N(_02937_));
 sg13g2_buf_2 _24959_ (.A(\grid.cell_7_3.se ),
    .X(_03348_));
 sg13g2_xor2_1 _24960_ (.B(_02947_),
    .A(_03348_),
    .X(_03349_));
 sg13g2_xnor2_1 _24961_ (.Y(_03350_),
    .A(_02492_),
    .B(_03300_));
 sg13g2_xnor2_1 _24962_ (.Y(_03351_),
    .A(_03349_),
    .B(_03350_));
 sg13g2_and2_1 _24963_ (.A(net1069),
    .B(_03351_),
    .X(_03352_));
 sg13g2_or2_1 _24964_ (.X(_03353_),
    .B(_02937_),
    .A(_02441_));
 sg13g2_a21oi_1 _24965_ (.A1(_03351_),
    .A2(_03353_),
    .Y(_03354_),
    .B1(net403));
 sg13g2_a221oi_1 _24966_ (.B2(net403),
    .C1(_03354_),
    .B1(_03352_),
    .A1(net196),
    .Y(_03355_),
    .A2(_03346_));
 sg13g2_nor2b_1 _24967_ (.A(net1069),
    .B_N(_03351_),
    .Y(_03356_));
 sg13g2_xnor2_1 _24968_ (.Y(_03357_),
    .A(net403),
    .B(_03351_));
 sg13g2_a22oi_1 _24969_ (.Y(_03359_),
    .B1(_03357_),
    .B2(net196),
    .A2(_03356_),
    .A1(_03345_));
 sg13g2_o21ai_1 _24970_ (.B1(_03359_),
    .Y(_03360_),
    .A1(_03345_),
    .A2(_03355_));
 sg13g2_buf_1 _24971_ (.A(_03348_),
    .X(_03361_));
 sg13g2_nand2_1 _24972_ (.Y(_03362_),
    .A(_02951_),
    .B(net728));
 sg13g2_xor2_1 _24973_ (.B(_03348_),
    .A(net1068),
    .X(_03363_));
 sg13g2_and2_1 _24974_ (.A(net410),
    .B(_03363_),
    .X(_03364_));
 sg13g2_nor2_1 _24975_ (.A(net410),
    .B(_03362_),
    .Y(_03365_));
 sg13g2_o21ai_1 _24976_ (.B1(_02573_),
    .Y(_03366_),
    .A1(_03364_),
    .A2(_03365_));
 sg13g2_o21ai_1 _24977_ (.B1(_03366_),
    .Y(_03367_),
    .A1(_02592_),
    .A2(_03362_));
 sg13g2_nand2_1 _24978_ (.Y(_03368_),
    .A(_02457_),
    .B(_03345_));
 sg13g2_inv_1 _24979_ (.Y(_03370_),
    .A(_03345_));
 sg13g2_nor3_1 _24980_ (.A(_02983_),
    .B(net729),
    .C(_02946_),
    .Y(_03371_));
 sg13g2_buf_1 _24981_ (.A(net728),
    .X(_03372_));
 sg13g2_a22oi_1 _24982_ (.Y(_03373_),
    .B1(_03371_),
    .B2(net392),
    .A2(_03370_),
    .A1(net196));
 sg13g2_nand2b_1 _24983_ (.Y(_03374_),
    .B(_03373_),
    .A_N(_03356_));
 sg13g2_a221oi_1 _24984_ (.B2(_03368_),
    .C1(_03374_),
    .B1(_03357_),
    .A1(net393),
    .Y(_03375_),
    .A2(_03367_));
 sg13g2_a21oi_1 _24985_ (.A1(_02555_),
    .A2(_03362_),
    .Y(_03376_),
    .B1(_03364_));
 sg13g2_a21oi_1 _24986_ (.A1(net410),
    .A2(net729),
    .Y(_03377_),
    .B1(_02555_));
 sg13g2_or3_1 _24987_ (.A(net738),
    .B(_03361_),
    .C(_03377_),
    .X(_03378_));
 sg13g2_o21ai_1 _24988_ (.B1(_03378_),
    .Y(_03379_),
    .A1(net393),
    .A2(_03376_));
 sg13g2_nand2_1 _24989_ (.Y(_03381_),
    .A(net195),
    .B(net409));
 sg13g2_nor3_1 _24990_ (.A(net393),
    .B(_02956_),
    .C(net392),
    .Y(_03382_));
 sg13g2_a22oi_1 _24991_ (.Y(_03383_),
    .B1(_03381_),
    .B2(_03382_),
    .A2(_03379_),
    .A1(_02592_));
 sg13g2_mux2_1 _24992_ (.A0(_03360_),
    .A1(_03375_),
    .S(_03383_),
    .X(_03384_));
 sg13g2_xor2_1 _24993_ (.B(_03357_),
    .A(_03258_),
    .X(_03385_));
 sg13g2_o21ai_1 _24994_ (.B1(net740),
    .Y(_03386_),
    .A1(_05471_),
    .A2(_03385_));
 sg13g2_o21ai_1 _24995_ (.B1(_03386_),
    .Y(_03387_),
    .A1(_08737_),
    .A2(_03384_));
 sg13g2_nand2_1 _24996_ (.Y(_03388_),
    .A(_00788_),
    .B(_03244_));
 sg13g2_nand2b_1 _24997_ (.Y(_03389_),
    .B(_06621_),
    .A_N(_03388_));
 sg13g2_o21ai_1 _24998_ (.B1(_03389_),
    .Y(_00512_),
    .A1(_03239_),
    .A2(_03387_));
 sg13g2_buf_1 _24999_ (.A(\grid.cell_7_4.se ),
    .X(_03391_));
 sg13g2_xor2_1 _25000_ (.B(net1064),
    .A(net1067),
    .X(_03392_));
 sg13g2_nand2_1 _25001_ (.Y(_03393_),
    .A(net737),
    .B(net1064));
 sg13g2_a22oi_1 _25002_ (.Y(_03394_),
    .B1(_03393_),
    .B2(_02597_),
    .A2(_03392_),
    .A1(net748));
 sg13g2_buf_1 _25003_ (.A(net1064),
    .X(_03395_));
 sg13g2_a21oi_1 _25004_ (.A1(net748),
    .A2(_03348_),
    .Y(_03396_),
    .B1(_02597_));
 sg13g2_or3_1 _25005_ (.A(net737),
    .B(net727),
    .C(_03396_),
    .X(_03397_));
 sg13g2_o21ai_1 _25006_ (.B1(_03397_),
    .Y(_03398_),
    .A1(net728),
    .A2(_03394_));
 sg13g2_nor2_1 _25007_ (.A(_02555_),
    .B(_02597_),
    .Y(_03399_));
 sg13g2_nor4_1 _25008_ (.A(_03361_),
    .B(_02990_),
    .C(net727),
    .D(_03399_),
    .Y(_03400_));
 sg13g2_a21o_1 _25009_ (.A2(_03398_),
    .A1(_02631_),
    .B1(_03400_),
    .X(_03402_));
 sg13g2_buf_1 _25010_ (.A(_00041_),
    .X(_03403_));
 sg13g2_xor2_1 _25011_ (.B(_02989_),
    .A(net1064),
    .X(_03404_));
 sg13g2_xnor2_1 _25012_ (.Y(_03405_),
    .A(_02554_),
    .B(_03348_));
 sg13g2_xnor2_1 _25013_ (.Y(_03406_),
    .A(_03404_),
    .B(_03405_));
 sg13g2_buf_2 _25014_ (.A(_03406_),
    .X(_03407_));
 sg13g2_a21o_1 _25015_ (.A2(_03407_),
    .A1(net740),
    .B1(_02501_),
    .X(_03408_));
 sg13g2_o21ai_1 _25016_ (.B1(_03407_),
    .Y(_03409_),
    .A1(net1066),
    .A2(net410));
 sg13g2_nor2_1 _25017_ (.A(_02983_),
    .B(net402),
    .Y(_03410_));
 sg13g2_a221oi_1 _25018_ (.B2(net402),
    .C1(_03410_),
    .B1(_03409_),
    .A1(_02985_),
    .Y(_03411_),
    .A2(_03408_));
 sg13g2_xnor2_1 _25019_ (.Y(_03413_),
    .A(net740),
    .B(_03407_));
 sg13g2_nor2b_1 _25020_ (.A(net1066),
    .B_N(_03407_),
    .Y(_03414_));
 sg13g2_a22oi_1 _25021_ (.Y(_03415_),
    .B1(_03414_),
    .B2(net1063),
    .A2(_03413_),
    .A1(net195));
 sg13g2_o21ai_1 _25022_ (.B1(_03415_),
    .Y(_03416_),
    .A1(net1063),
    .A2(_03411_));
 sg13g2_and2_1 _25023_ (.A(net737),
    .B(net1064),
    .X(_03417_));
 sg13g2_buf_1 _25024_ (.A(_03417_),
    .X(_03418_));
 sg13g2_nand2_1 _25025_ (.Y(_03419_),
    .A(net748),
    .B(_03392_));
 sg13g2_o21ai_1 _25026_ (.B1(_03419_),
    .Y(_03420_),
    .A1(net748),
    .A2(_03393_));
 sg13g2_a22oi_1 _25027_ (.Y(_03421_),
    .B1(_03420_),
    .B2(net408),
    .A2(_03418_),
    .A1(_02639_));
 sg13g2_a21oi_1 _25028_ (.A1(_03418_),
    .A2(_03399_),
    .Y(_03422_),
    .B1(net392));
 sg13g2_a21oi_1 _25029_ (.A1(net392),
    .A2(_03421_),
    .Y(_03424_),
    .B1(_03422_));
 sg13g2_nor3_1 _25030_ (.A(_03402_),
    .B(_03414_),
    .C(_03424_),
    .Y(_03425_));
 sg13g2_nand2_1 _25031_ (.Y(_03426_),
    .A(net195),
    .B(_03413_));
 sg13g2_nor2_1 _25032_ (.A(_02563_),
    .B(_03413_),
    .Y(_03427_));
 sg13g2_a21o_1 _25033_ (.A2(_03426_),
    .A1(net1063),
    .B1(_03427_),
    .X(_03428_));
 sg13g2_a221oi_1 _25034_ (.B2(_03428_),
    .C1(_06285_),
    .B1(_03425_),
    .A1(_03402_),
    .Y(_03429_),
    .A2(_03416_));
 sg13g2_xor2_1 _25035_ (.B(_03407_),
    .A(_03330_),
    .X(_03430_));
 sg13g2_a21oi_1 _25036_ (.A1(net70),
    .A2(_03430_),
    .Y(_03431_),
    .B1(_02956_));
 sg13g2_or3_1 _25037_ (.A(_03239_),
    .B(_03429_),
    .C(_03431_),
    .X(_03432_));
 sg13g2_o21ai_1 _25038_ (.B1(_03432_),
    .Y(_00513_),
    .A1(_12298_),
    .A2(_03388_));
 sg13g2_buf_2 _25039_ (.A(_00073_),
    .X(_03434_));
 sg13g2_nand2_1 _25040_ (.Y(_03435_),
    .A(_03434_),
    .B(_02555_));
 sg13g2_buf_1 _25041_ (.A(\grid.cell_7_5.se ),
    .X(_03436_));
 sg13g2_buf_1 _25042_ (.A(_03436_),
    .X(_03437_));
 sg13g2_xnor2_1 _25043_ (.Y(_03438_),
    .A(net1064),
    .B(net726));
 sg13g2_xnor2_1 _25044_ (.Y(_03439_),
    .A(_03021_),
    .B(_03438_));
 sg13g2_xnor2_1 _25045_ (.Y(_03440_),
    .A(_02596_),
    .B(_03439_));
 sg13g2_xnor2_1 _25046_ (.Y(_03441_),
    .A(net738),
    .B(_03440_));
 sg13g2_inv_1 _25047_ (.Y(_03442_),
    .A(_03434_));
 sg13g2_nand2_1 _25048_ (.Y(_03443_),
    .A(_03442_),
    .B(_02573_));
 sg13g2_o21ai_1 _25049_ (.B1(_03443_),
    .Y(_03445_),
    .A1(_03037_),
    .A2(_03440_));
 sg13g2_a21oi_1 _25050_ (.A1(_03435_),
    .A2(_03441_),
    .Y(_03446_),
    .B1(_03445_));
 sg13g2_buf_1 _25051_ (.A(_03395_),
    .X(_03447_));
 sg13g2_xor2_1 _25052_ (.B(_03437_),
    .A(_03017_),
    .X(_03448_));
 sg13g2_nand2_1 _25053_ (.Y(_03449_),
    .A(_03016_),
    .B(net726));
 sg13g2_buf_2 _25054_ (.A(_03449_),
    .X(_03450_));
 sg13g2_a22oi_1 _25055_ (.Y(_03451_),
    .B1(_03450_),
    .B2(net193),
    .A2(_03448_),
    .A1(net747));
 sg13g2_and2_1 _25056_ (.A(net747),
    .B(net727),
    .X(_03452_));
 sg13g2_buf_1 _25057_ (.A(net726),
    .X(_03453_));
 sg13g2_nor2_1 _25058_ (.A(net736),
    .B(net390),
    .Y(_03454_));
 sg13g2_o21ai_1 _25059_ (.B1(_03454_),
    .Y(_03456_),
    .A1(net193),
    .A2(_03452_));
 sg13g2_o21ai_1 _25060_ (.B1(_03456_),
    .Y(_03457_),
    .A1(net391),
    .A2(_03451_));
 sg13g2_nand2_1 _25061_ (.Y(_03458_),
    .A(_02606_),
    .B(net194));
 sg13g2_buf_1 _25062_ (.A(_03437_),
    .X(_03459_));
 sg13g2_buf_1 _25063_ (.A(net389),
    .X(_03460_));
 sg13g2_nor3_1 _25064_ (.A(net391),
    .B(net188),
    .C(net185),
    .Y(_03461_));
 sg13g2_a22oi_1 _25065_ (.Y(_03462_),
    .B1(_03458_),
    .B2(_03461_),
    .A2(_03457_),
    .A1(_02692_));
 sg13g2_xor2_1 _25066_ (.B(_03462_),
    .A(_03446_),
    .X(_03463_));
 sg13g2_nand2_1 _25067_ (.Y(_03464_),
    .A(_02606_),
    .B(_03448_));
 sg13g2_o21ai_1 _25068_ (.B1(_03464_),
    .Y(_03465_),
    .A1(net408),
    .A2(_03450_));
 sg13g2_nor2_1 _25069_ (.A(_02692_),
    .B(_03450_),
    .Y(_03467_));
 sg13g2_a21oi_1 _25070_ (.A1(net194),
    .A2(_03465_),
    .Y(_03468_),
    .B1(_03467_));
 sg13g2_nor2b_1 _25071_ (.A(_03468_),
    .B_N(net391),
    .Y(_03469_));
 sg13g2_nor3_1 _25072_ (.A(net391),
    .B(_03450_),
    .C(_03458_),
    .Y(_03470_));
 sg13g2_nor4_1 _25073_ (.A(_03037_),
    .B(_03434_),
    .C(_02947_),
    .D(_03440_),
    .Y(_03471_));
 sg13g2_nor4_1 _25074_ (.A(_03463_),
    .B(_03469_),
    .C(_03470_),
    .D(_03471_),
    .Y(_03472_));
 sg13g2_xnor2_1 _25075_ (.Y(_03473_),
    .A(_03349_),
    .B(_03440_));
 sg13g2_a21oi_1 _25076_ (.A1(net114),
    .A2(_03473_),
    .Y(_03474_),
    .B1(net400));
 sg13g2_nor2_1 _25077_ (.A(_03239_),
    .B(_03474_),
    .Y(_03475_));
 sg13g2_o21ai_1 _25078_ (.B1(_03475_),
    .Y(_03476_),
    .A1(_05472_),
    .A2(_03472_));
 sg13g2_o21ai_1 _25079_ (.B1(_03476_),
    .Y(_00514_),
    .A1(net43),
    .A2(_03388_));
 sg13g2_buf_1 _25080_ (.A(_00105_),
    .X(_03478_));
 sg13g2_inv_1 _25081_ (.Y(_03479_),
    .A(_03478_));
 sg13g2_xnor2_1 _25082_ (.Y(_03480_),
    .A(_03436_),
    .B(_03166_));
 sg13g2_xor2_1 _25083_ (.B(_03480_),
    .A(_02813_),
    .X(_03481_));
 sg13g2_xnor2_1 _25084_ (.Y(_03482_),
    .A(net407),
    .B(_03481_));
 sg13g2_xnor2_1 _25085_ (.Y(_03483_),
    .A(_02979_),
    .B(_03482_));
 sg13g2_o21ai_1 _25086_ (.B1(_03483_),
    .Y(_03484_),
    .A1(_03479_),
    .A2(_02613_));
 sg13g2_nand2b_1 _25087_ (.Y(_03485_),
    .B(_03482_),
    .A_N(_03080_));
 sg13g2_nand2_1 _25088_ (.Y(_03486_),
    .A(_03479_),
    .B(_02613_));
 sg13g2_nand3_1 _25089_ (.B(_03485_),
    .C(_03486_),
    .A(_03484_),
    .Y(_03488_));
 sg13g2_or2_1 _25090_ (.X(_03489_),
    .B(_03221_),
    .A(net389));
 sg13g2_buf_2 _25091_ (.A(_00135_),
    .X(_03490_));
 sg13g2_o21ai_1 _25092_ (.B1(_03221_),
    .Y(_03491_),
    .A1(net185),
    .A2(_03223_));
 sg13g2_nand2_1 _25093_ (.Y(_03492_),
    .A(_03490_),
    .B(_03491_));
 sg13g2_a21oi_1 _25094_ (.A1(_03489_),
    .A2(_03492_),
    .Y(_03493_),
    .B1(net192));
 sg13g2_and2_1 _25095_ (.A(_03490_),
    .B(net389),
    .X(_03494_));
 sg13g2_xor2_1 _25096_ (.B(net389),
    .A(_03490_),
    .X(_03495_));
 sg13g2_nor2_1 _25097_ (.A(_03490_),
    .B(_03233_),
    .Y(_03496_));
 sg13g2_a221oi_1 _25098_ (.B2(_03221_),
    .C1(_03496_),
    .B1(_03495_),
    .A1(_03233_),
    .Y(_03497_),
    .A2(_03494_));
 sg13g2_nand3_1 _25099_ (.B(net414),
    .C(_03223_),
    .A(net185),
    .Y(_03499_));
 sg13g2_nand2_1 _25100_ (.Y(_03500_),
    .A(_03489_),
    .B(_03499_));
 sg13g2_a22oi_1 _25101_ (.Y(_03501_),
    .B1(_03500_),
    .B2(_02680_),
    .A2(_03496_),
    .A1(net185));
 sg13g2_o21ai_1 _25102_ (.B1(_03501_),
    .Y(_03502_),
    .A1(_02716_),
    .A2(_03497_));
 sg13g2_nor2_1 _25103_ (.A(_03493_),
    .B(_03502_),
    .Y(_03503_));
 sg13g2_xor2_1 _25104_ (.B(_03503_),
    .A(_03488_),
    .X(_03504_));
 sg13g2_nor3_1 _25105_ (.A(_03478_),
    .B(_02989_),
    .C(_03485_),
    .Y(_03505_));
 sg13g2_nand2_1 _25106_ (.Y(_03506_),
    .A(_02653_),
    .B(_03167_));
 sg13g2_o21ai_1 _25107_ (.B1(_03506_),
    .Y(_03507_),
    .A1(_02654_),
    .A2(_03233_));
 sg13g2_a21oi_1 _25108_ (.A1(_02685_),
    .A2(_03507_),
    .Y(_03508_),
    .B1(_03496_));
 sg13g2_a21oi_1 _25109_ (.A1(_02741_),
    .A2(_03223_),
    .Y(_03510_),
    .B1(net185));
 sg13g2_a21oi_1 _25110_ (.A1(net185),
    .A2(_03508_),
    .Y(_03511_),
    .B1(_03510_));
 sg13g2_xor2_1 _25111_ (.B(_03482_),
    .A(_03404_),
    .X(_03512_));
 sg13g2_nor2_1 _25112_ (.A(net133),
    .B(_03512_),
    .Y(_03513_));
 sg13g2_nor4_1 _25113_ (.A(_07553_),
    .B(_03505_),
    .C(_03511_),
    .D(_03513_),
    .Y(_03514_));
 sg13g2_nand2_1 _25114_ (.Y(_03515_),
    .A(_03504_),
    .B(_03514_));
 sg13g2_a22oi_1 _25115_ (.Y(_03516_),
    .B1(_07562_),
    .B2(_03180_),
    .A2(_07199_),
    .A1(net133));
 sg13g2_a221oi_1 _25116_ (.B2(_03516_),
    .C1(_08965_),
    .B1(_03515_),
    .A1(_06813_),
    .Y(_00515_),
    .A2(_03180_));
 sg13g2_a22oi_1 _25117_ (.Y(_03517_),
    .B1(_06468_),
    .B2(_03180_),
    .A2(_07117_),
    .A1(net95));
 sg13g2_xor2_1 _25118_ (.B(_03480_),
    .A(_03021_),
    .X(_03518_));
 sg13g2_xnor2_1 _25119_ (.Y(_03520_),
    .A(_02389_),
    .B(_03518_));
 sg13g2_buf_2 _25120_ (.A(_03520_),
    .X(_03521_));
 sg13g2_xnor2_1 _25121_ (.Y(_03522_),
    .A(net1071),
    .B(_03521_));
 sg13g2_nor2_1 _25122_ (.A(_02483_),
    .B(_03522_),
    .Y(_03523_));
 sg13g2_inv_1 _25123_ (.Y(_03524_),
    .A(_03490_));
 sg13g2_nand2_1 _25124_ (.Y(_03525_),
    .A(net726),
    .B(net733));
 sg13g2_buf_1 _25125_ (.A(_03525_),
    .X(_03526_));
 sg13g2_mux2_1 _25126_ (.A0(net390),
    .A1(_03526_),
    .S(net736),
    .X(_03527_));
 sg13g2_a22oi_1 _25127_ (.Y(_03528_),
    .B1(_03527_),
    .B2(net414),
    .A2(_03454_),
    .A1(net187));
 sg13g2_o21ai_1 _25128_ (.B1(net736),
    .Y(_03529_),
    .A1(net726),
    .A2(net733));
 sg13g2_a21oi_1 _25129_ (.A1(_03526_),
    .A2(_03529_),
    .Y(_03531_),
    .B1(_02369_));
 sg13g2_nand2_1 _25130_ (.Y(_03532_),
    .A(_03524_),
    .B(_03531_));
 sg13g2_o21ai_1 _25131_ (.B1(_03532_),
    .Y(_03533_),
    .A1(_03524_),
    .A2(_03528_));
 sg13g2_or3_1 _25132_ (.A(_03017_),
    .B(net726),
    .C(net733),
    .X(_03534_));
 sg13g2_nand3_1 _25133_ (.B(_03526_),
    .C(_03529_),
    .A(_03490_),
    .Y(_03535_));
 sg13g2_a21oi_1 _25134_ (.A1(_03534_),
    .A2(_03535_),
    .Y(_03536_),
    .B1(_02400_));
 sg13g2_nand2_1 _25135_ (.Y(_03537_),
    .A(_02379_),
    .B(net397));
 sg13g2_o21ai_1 _25136_ (.B1(_03534_),
    .Y(_03538_),
    .A1(_03450_),
    .A2(_03537_));
 sg13g2_nor2_1 _25137_ (.A(_03490_),
    .B(_03526_),
    .Y(_03539_));
 sg13g2_a22oi_1 _25138_ (.Y(_03540_),
    .B1(_03539_),
    .B2(net399),
    .A2(_03538_),
    .A1(_02678_));
 sg13g2_nand2b_1 _25139_ (.Y(_03542_),
    .B(_03540_),
    .A_N(_03536_));
 sg13g2_a21oi_2 _25140_ (.B1(_03542_),
    .Y(_03543_),
    .A2(_03533_),
    .A1(_02654_));
 sg13g2_nand2_1 _25141_ (.Y(_03544_),
    .A(net1071),
    .B(_02770_));
 sg13g2_nor2_1 _25142_ (.A(net1071),
    .B(_02770_),
    .Y(_03545_));
 sg13g2_inv_1 _25143_ (.Y(_03546_),
    .A(_02819_));
 sg13g2_nor2_1 _25144_ (.A(_03546_),
    .B(_03521_),
    .Y(_03547_));
 sg13g2_a221oi_1 _25145_ (.B2(_03521_),
    .C1(_03547_),
    .B1(_03545_),
    .A1(_02427_),
    .Y(_03548_),
    .A2(_03544_));
 sg13g2_or3_1 _25146_ (.A(net734),
    .B(_03543_),
    .C(_03548_),
    .X(_03549_));
 sg13g2_and2_1 _25147_ (.A(_02770_),
    .B(_03521_),
    .X(_03550_));
 sg13g2_o21ai_1 _25148_ (.B1(net734),
    .Y(_03551_),
    .A1(_03543_),
    .A2(_03550_));
 sg13g2_nand3b_1 _25149_ (.B(_03549_),
    .C(_03551_),
    .Y(_03553_),
    .A_N(_03523_));
 sg13g2_and2_1 _25150_ (.A(net743),
    .B(_03521_),
    .X(_03554_));
 sg13g2_o21ai_1 _25151_ (.B1(_03554_),
    .Y(_03555_),
    .A1(_02770_),
    .A2(_03543_));
 sg13g2_nand3b_1 _25152_ (.B(_03543_),
    .C(_03546_),
    .Y(_03556_),
    .A_N(_03521_));
 sg13g2_a21oi_1 _25153_ (.A1(_03555_),
    .A2(_03556_),
    .Y(_03557_),
    .B1(net753));
 sg13g2_nand2b_1 _25154_ (.Y(_03558_),
    .B(net407),
    .A_N(_03480_));
 sg13g2_o21ai_1 _25155_ (.B1(_03558_),
    .Y(_03559_),
    .A1(_02653_),
    .A2(_03526_));
 sg13g2_a21oi_1 _25156_ (.A1(_02685_),
    .A2(_03559_),
    .Y(_03560_),
    .B1(_03539_));
 sg13g2_nor2_1 _25157_ (.A(_03061_),
    .B(_03560_),
    .Y(_03561_));
 sg13g2_nor3_1 _25158_ (.A(net133),
    .B(_02716_),
    .C(_03526_),
    .Y(_03562_));
 sg13g2_xor2_1 _25159_ (.B(_03521_),
    .A(_03293_),
    .X(_03564_));
 sg13g2_o21ai_1 _25160_ (.B1(_02809_),
    .Y(_03565_),
    .A1(net95),
    .A2(_03564_));
 sg13g2_nor3_1 _25161_ (.A(_03561_),
    .B(_03562_),
    .C(_03565_),
    .Y(_03566_));
 sg13g2_o21ai_1 _25162_ (.B1(_03543_),
    .Y(_03567_),
    .A1(_03523_),
    .A2(_03550_));
 sg13g2_and2_1 _25163_ (.A(_03566_),
    .B(_03567_),
    .X(_03568_));
 sg13g2_o21ai_1 _25164_ (.B1(_03568_),
    .Y(_03569_),
    .A1(_03553_),
    .A2(_03557_));
 sg13g2_o21ai_1 _25165_ (.B1(net435),
    .Y(_03570_),
    .A1(_11347_),
    .A2(_03243_));
 sg13g2_a21oi_1 _25166_ (.A1(_03517_),
    .A2(_03569_),
    .Y(_00516_),
    .B1(_03570_));
 sg13g2_nand3_1 _25167_ (.B(_01967_),
    .C(_05180_),
    .A(_01913_),
    .Y(_03571_));
 sg13g2_nor2_2 _25168_ (.A(_02043_),
    .B(_03571_),
    .Y(_03572_));
 sg13g2_nand2_1 _25169_ (.Y(_03574_),
    .A(net44),
    .B(_03572_));
 sg13g2_xnor2_1 _25170_ (.Y(_03575_),
    .A(net1016),
    .B(_05202_));
 sg13g2_xor2_1 _25171_ (.B(_03575_),
    .A(_03167_),
    .X(_03576_));
 sg13g2_xnor2_1 _25172_ (.Y(_03577_),
    .A(net191),
    .B(_03576_));
 sg13g2_nor2_1 _25173_ (.A(_03336_),
    .B(_03577_),
    .Y(_03578_));
 sg13g2_or2_1 _25174_ (.X(_03579_),
    .B(net733),
    .A(net1013));
 sg13g2_buf_1 _25175_ (.A(_03579_),
    .X(_03580_));
 sg13g2_nand2_1 _25176_ (.Y(_03581_),
    .A(net351),
    .B(net189));
 sg13g2_nand4_1 _25177_ (.B(net336),
    .C(net187),
    .A(net682),
    .Y(_03582_),
    .D(_02886_));
 sg13g2_o21ai_1 _25178_ (.B1(_03582_),
    .Y(_03583_),
    .A1(_03580_),
    .A2(_03581_));
 sg13g2_nand2b_1 _25179_ (.Y(_03585_),
    .B(net397),
    .A_N(_02885_));
 sg13g2_nor2_1 _25180_ (.A(net677),
    .B(_03203_),
    .Y(_03586_));
 sg13g2_a21oi_1 _25181_ (.A1(net336),
    .A2(_03585_),
    .Y(_03587_),
    .B1(_03586_));
 sg13g2_nor2_1 _25182_ (.A(net677),
    .B(net187),
    .Y(_03588_));
 sg13g2_inv_1 _25183_ (.Y(_03589_),
    .A(net676));
 sg13g2_nor2b_1 _25184_ (.A(_03187_),
    .B_N(net676),
    .Y(_03590_));
 sg13g2_a21o_1 _25185_ (.A2(net189),
    .A1(_03589_),
    .B1(_03590_),
    .X(_03591_));
 sg13g2_a22oi_1 _25186_ (.Y(_03592_),
    .B1(_03591_),
    .B2(net191),
    .A2(_03588_),
    .A1(_03329_));
 sg13g2_o21ai_1 _25187_ (.B1(_03592_),
    .Y(_03593_),
    .A1(net132),
    .A2(_03587_));
 sg13g2_buf_1 _25188_ (.A(_05190_),
    .X(_03594_));
 sg13g2_nand3_1 _25189_ (.B(net132),
    .C(_03580_),
    .A(net191),
    .Y(_03596_));
 sg13g2_nand2b_1 _25190_ (.Y(_03597_),
    .B(_03187_),
    .A_N(_02760_));
 sg13g2_o21ai_1 _25191_ (.B1(_03597_),
    .Y(_03598_),
    .A1(_03208_),
    .A2(net741));
 sg13g2_nor2_1 _25192_ (.A(net677),
    .B(_03585_),
    .Y(_03599_));
 sg13g2_a21oi_1 _25193_ (.A1(net336),
    .A2(_03598_),
    .Y(_03600_),
    .B1(_03599_));
 sg13g2_a21oi_1 _25194_ (.A1(_03596_),
    .A2(_03600_),
    .Y(_03601_),
    .B1(net682));
 sg13g2_a221oi_1 _25195_ (.B2(net184),
    .C1(_03601_),
    .B1(_03593_),
    .A1(net405),
    .Y(_03602_),
    .A2(_03583_));
 sg13g2_nor2_1 _25196_ (.A(_03578_),
    .B(_03602_),
    .Y(_03603_));
 sg13g2_xnor2_1 _25197_ (.Y(_03604_),
    .A(_03170_),
    .B(_03575_));
 sg13g2_nor2_1 _25198_ (.A(_05220_),
    .B(_03604_),
    .Y(_03605_));
 sg13g2_nand2_1 _25199_ (.Y(_03607_),
    .A(_05221_),
    .B(_03604_));
 sg13g2_o21ai_1 _25200_ (.B1(_03607_),
    .Y(_03608_),
    .A1(net743),
    .A2(_03605_));
 sg13g2_and2_1 _25201_ (.A(_05209_),
    .B(net733),
    .X(_03609_));
 sg13g2_buf_1 _25202_ (.A(_03609_),
    .X(_03610_));
 sg13g2_o21ai_1 _25203_ (.B1(_02780_),
    .Y(_03611_),
    .A1(_03586_),
    .A2(_03590_));
 sg13g2_o21ai_1 _25204_ (.B1(_03611_),
    .Y(_03612_),
    .A1(net132),
    .A2(_03610_));
 sg13g2_nand2_1 _25205_ (.Y(_03613_),
    .A(net405),
    .B(_03139_));
 sg13g2_a22oi_1 _25206_ (.Y(_03614_),
    .B1(_03613_),
    .B2(_03588_),
    .A2(_03612_),
    .A1(net741));
 sg13g2_o21ai_1 _25207_ (.B1(_03139_),
    .Y(_03615_),
    .A1(_02782_),
    .A2(net351));
 sg13g2_nand3_1 _25208_ (.B(_03588_),
    .C(_03615_),
    .A(_02886_),
    .Y(_03616_));
 sg13g2_o21ai_1 _25209_ (.B1(_03616_),
    .Y(_03618_),
    .A1(net184),
    .A2(_03614_));
 sg13g2_o21ai_1 _25210_ (.B1(_03604_),
    .Y(_03619_),
    .A1(_05221_),
    .A2(_03578_));
 sg13g2_xor2_1 _25211_ (.B(_03575_),
    .A(_03170_),
    .X(_03620_));
 sg13g2_o21ai_1 _25212_ (.B1(_05243_),
    .Y(_03621_),
    .A1(net1071),
    .A2(_03620_));
 sg13g2_mux2_1 _25213_ (.A0(_03605_),
    .A1(_03621_),
    .S(_03578_),
    .X(_03622_));
 sg13g2_a21o_1 _25214_ (.A2(_03619_),
    .A1(net743),
    .B1(_03622_),
    .X(_03623_));
 sg13g2_a221oi_1 _25215_ (.B2(_03623_),
    .C1(_05131_),
    .B1(_03618_),
    .A1(_03603_),
    .Y(_03624_),
    .A2(_03608_));
 sg13g2_xnor2_1 _25216_ (.Y(_03625_),
    .A(_02819_),
    .B(net1006));
 sg13g2_xnor2_1 _25217_ (.Y(_03626_),
    .A(_03620_),
    .B(_03625_));
 sg13g2_a21oi_1 _25218_ (.A1(net113),
    .A2(_03626_),
    .Y(_03627_),
    .B1(net398));
 sg13g2_or3_1 _25219_ (.A(_03572_),
    .B(_03624_),
    .C(_03627_),
    .X(_03629_));
 sg13g2_a21oi_1 _25220_ (.A1(_03574_),
    .A2(_03629_),
    .Y(_00517_),
    .B1(net440));
 sg13g2_nor2b_1 _25221_ (.A(_01989_),
    .B_N(_05180_),
    .Y(_03630_));
 sg13g2_nand2_2 _25222_ (.Y(_03631_),
    .A(net158),
    .B(_03630_));
 sg13g2_xnor2_1 _25223_ (.Y(_03632_),
    .A(net744),
    .B(net1016));
 sg13g2_xnor2_1 _25224_ (.Y(_03633_),
    .A(net1005),
    .B(_03247_));
 sg13g2_xnor2_1 _25225_ (.Y(_03634_),
    .A(_03632_),
    .B(_03633_));
 sg13g2_buf_1 _25226_ (.A(_03634_),
    .X(_03635_));
 sg13g2_xnor2_1 _25227_ (.Y(_03636_),
    .A(net735),
    .B(_03635_));
 sg13g2_nand2b_1 _25228_ (.Y(_03637_),
    .B(net743),
    .A_N(_03636_));
 sg13g2_a21oi_1 _25229_ (.A1(net398),
    .A2(net730),
    .Y(_03639_),
    .B1(_03546_));
 sg13g2_nor2_1 _25230_ (.A(_03175_),
    .B(net730),
    .Y(_03640_));
 sg13g2_mux2_1 _25231_ (.A0(net398),
    .A1(_03640_),
    .S(_03635_),
    .X(_03641_));
 sg13g2_and2_1 _25232_ (.A(_02761_),
    .B(net1070),
    .X(_03642_));
 sg13g2_buf_1 _25233_ (.A(_03642_),
    .X(_03643_));
 sg13g2_nor2b_1 _25234_ (.A(_02885_),
    .B_N(net1005),
    .Y(_03644_));
 sg13g2_a21o_1 _25235_ (.A2(_03643_),
    .A1(_05318_),
    .B1(_03644_),
    .X(_03645_));
 sg13g2_nand2_1 _25236_ (.Y(_03646_),
    .A(_05319_),
    .B(_03329_));
 sg13g2_nor2b_1 _25237_ (.A(net731),
    .B_N(_03643_),
    .Y(_03647_));
 sg13g2_a221oi_1 _25238_ (.B2(_03647_),
    .C1(net351),
    .B1(_03646_),
    .A1(_03248_),
    .Y(_03648_),
    .A2(_03645_));
 sg13g2_nand2b_1 _25239_ (.Y(_03650_),
    .B(_02885_),
    .A_N(net1005));
 sg13g2_o21ai_1 _25240_ (.B1(_03650_),
    .Y(_03651_),
    .A1(_03248_),
    .A2(_03644_));
 sg13g2_o21ai_1 _25241_ (.B1(_03246_),
    .Y(_03652_),
    .A1(net1005),
    .A2(_02885_));
 sg13g2_o21ai_1 _25242_ (.B1(_03652_),
    .Y(_03653_),
    .A1(_05318_),
    .A2(_03329_));
 sg13g2_a221oi_1 _25243_ (.B2(_03643_),
    .C1(net682),
    .B1(_03653_),
    .A1(net403),
    .Y(_03654_),
    .A2(_03651_));
 sg13g2_or2_1 _25244_ (.X(_03655_),
    .B(_05305_),
    .A(_03246_));
 sg13g2_nand4_1 _25245_ (.B(net1070),
    .C(net731),
    .A(net1016),
    .Y(_03656_),
    .D(net669));
 sg13g2_o21ai_1 _25246_ (.B1(_03656_),
    .Y(_03657_),
    .A1(net675),
    .A2(_03655_));
 sg13g2_nor3_1 _25247_ (.A(net742),
    .B(_03329_),
    .C(_03655_),
    .Y(_03658_));
 sg13g2_a21oi_1 _25248_ (.A1(_02782_),
    .A2(_03657_),
    .Y(_03659_),
    .B1(_03658_));
 sg13g2_o21ai_1 _25249_ (.B1(_03659_),
    .Y(_03661_),
    .A1(_03648_),
    .A2(_03654_));
 sg13g2_buf_1 _25250_ (.A(_03661_),
    .X(_03662_));
 sg13g2_and2_1 _25251_ (.A(_05243_),
    .B(_03662_),
    .X(_03663_));
 sg13g2_o21ai_1 _25252_ (.B1(_03663_),
    .Y(_03664_),
    .A1(_03639_),
    .A2(_03641_));
 sg13g2_nand2_1 _25253_ (.Y(_03665_),
    .A(_03262_),
    .B(_03635_));
 sg13g2_a21o_1 _25254_ (.A2(_03665_),
    .A1(_03662_),
    .B1(_05243_),
    .X(_03666_));
 sg13g2_nand2_1 _25255_ (.Y(_03667_),
    .A(net398),
    .B(_03635_));
 sg13g2_a21oi_1 _25256_ (.A1(net734),
    .A2(_03662_),
    .Y(_03668_),
    .B1(_03667_));
 sg13g2_nor3_1 _25257_ (.A(net398),
    .B(_03635_),
    .C(_03662_),
    .Y(_03669_));
 sg13g2_o21ai_1 _25258_ (.B1(_03546_),
    .Y(_03670_),
    .A1(_03668_),
    .A2(_03669_));
 sg13g2_nand4_1 _25259_ (.B(_03664_),
    .C(_03666_),
    .A(_03637_),
    .Y(_03672_),
    .D(_03670_));
 sg13g2_xor2_1 _25260_ (.B(_03636_),
    .A(_03625_),
    .X(_03673_));
 sg13g2_nor2_1 _25261_ (.A(_03202_),
    .B(_03673_),
    .Y(_03674_));
 sg13g2_a21oi_1 _25262_ (.A1(_03637_),
    .A2(_03665_),
    .Y(_03675_),
    .B1(_03662_));
 sg13g2_and2_1 _25263_ (.A(net394),
    .B(_05306_),
    .X(_03676_));
 sg13g2_buf_1 _25264_ (.A(_03676_),
    .X(_03677_));
 sg13g2_xor2_1 _25265_ (.B(_05306_),
    .A(_03249_),
    .X(_03678_));
 sg13g2_mux2_1 _25266_ (.A0(_03677_),
    .A1(_03678_),
    .S(net744),
    .X(_03679_));
 sg13g2_a22oi_1 _25267_ (.Y(_03680_),
    .B1(_03679_),
    .B2(_02905_),
    .A2(_03677_),
    .A1(_03329_));
 sg13g2_a21oi_1 _25268_ (.A1(_03677_),
    .A2(_03643_),
    .Y(_03681_),
    .B1(_03594_));
 sg13g2_a21oi_1 _25269_ (.A1(net184),
    .A2(_03680_),
    .Y(_03683_),
    .B1(_03681_));
 sg13g2_nor4_1 _25270_ (.A(_06285_),
    .B(_03674_),
    .C(_03675_),
    .D(_03683_),
    .Y(_03684_));
 sg13g2_a22oi_1 _25271_ (.Y(_03685_),
    .B1(_03672_),
    .B2(_03684_),
    .A2(net74),
    .A1(_03202_));
 sg13g2_o21ai_1 _25272_ (.B1(net435),
    .Y(_03686_),
    .A1(net38),
    .A2(_03631_));
 sg13g2_a21oi_1 _25273_ (.A1(_03631_),
    .A2(_03685_),
    .Y(_00518_),
    .B1(_03686_));
 sg13g2_nand2_1 _25274_ (.Y(_03687_),
    .A(_12988_),
    .B(_03572_));
 sg13g2_and2_1 _25275_ (.A(net999),
    .B(_03301_),
    .X(_03688_));
 sg13g2_xor2_1 _25276_ (.B(_03300_),
    .A(net999),
    .X(_03689_));
 sg13g2_nand2_1 _25277_ (.Y(_03690_),
    .A(net404),
    .B(_03689_));
 sg13g2_o21ai_1 _25278_ (.B1(_03690_),
    .Y(_03691_),
    .A1(_02922_),
    .A2(_03688_));
 sg13g2_nand2_1 _25279_ (.Y(_03693_),
    .A(net190),
    .B(_02945_));
 sg13g2_nor2_1 _25280_ (.A(net665),
    .B(net729),
    .Y(_03694_));
 sg13g2_a22oi_1 _25281_ (.Y(_03695_),
    .B1(_03693_),
    .B2(_03694_),
    .A2(_03691_),
    .A1(net1069));
 sg13g2_o21ai_1 _25282_ (.B1(net402),
    .Y(_03696_),
    .A1(net403),
    .A2(_05319_));
 sg13g2_nand3_1 _25283_ (.B(_03696_),
    .C(_03694_),
    .A(net1069),
    .Y(_03697_));
 sg13g2_o21ai_1 _25284_ (.B1(_03697_),
    .Y(_03698_),
    .A1(_05357_),
    .A2(_03695_));
 sg13g2_nor2_1 _25285_ (.A(_02810_),
    .B(_05382_),
    .Y(_03699_));
 sg13g2_xnor2_1 _25286_ (.Y(_03700_),
    .A(net999),
    .B(_03312_));
 sg13g2_xnor2_1 _25287_ (.Y(_03701_),
    .A(_02831_),
    .B(_05305_));
 sg13g2_xnor2_1 _25288_ (.Y(_03702_),
    .A(_03700_),
    .B(_03701_));
 sg13g2_xnor2_1 _25289_ (.Y(_03704_),
    .A(_03201_),
    .B(_03702_));
 sg13g2_a22oi_1 _25290_ (.Y(_03705_),
    .B1(_03338_),
    .B2(_03702_),
    .A2(_05382_),
    .A1(_02810_));
 sg13g2_o21ai_1 _25291_ (.B1(_03705_),
    .Y(_03706_),
    .A1(_03699_),
    .A2(_03704_));
 sg13g2_xnor2_1 _25292_ (.Y(_03707_),
    .A(_03698_),
    .B(_03706_));
 sg13g2_nand2_1 _25293_ (.Y(_03708_),
    .A(_05366_),
    .B(_03301_));
 sg13g2_o21ai_1 _25294_ (.B1(_03690_),
    .Y(_03709_),
    .A1(net404),
    .A2(_03708_));
 sg13g2_nand2_1 _25295_ (.Y(_03710_),
    .A(_02945_),
    .B(_03709_));
 sg13g2_o21ai_1 _25296_ (.B1(_03710_),
    .Y(_03711_),
    .A1(net1069),
    .A2(_03708_));
 sg13g2_nor3_1 _25297_ (.A(_02915_),
    .B(net348),
    .C(_03302_),
    .Y(_03712_));
 sg13g2_and4_1 _25298_ (.A(_05382_),
    .B(_03338_),
    .C(_03169_),
    .D(_03702_),
    .X(_03713_));
 sg13g2_a221oi_1 _25299_ (.B2(net347),
    .C1(_03713_),
    .B1(_03712_),
    .A1(_05357_),
    .Y(_03715_),
    .A2(_03711_));
 sg13g2_a21oi_1 _25300_ (.A1(_03707_),
    .A2(_03715_),
    .Y(_03716_),
    .B1(net117));
 sg13g2_xnor2_1 _25301_ (.Y(_03717_),
    .A(net351),
    .B(_03169_));
 sg13g2_xnor2_1 _25302_ (.Y(_03718_),
    .A(_03702_),
    .B(_03717_));
 sg13g2_a21oi_1 _25303_ (.A1(net122),
    .A2(_03718_),
    .Y(_03719_),
    .B1(net186));
 sg13g2_nand2_1 _25304_ (.Y(_03720_),
    .A(_00777_),
    .B(_03631_));
 sg13g2_or3_1 _25305_ (.A(_03716_),
    .B(_03719_),
    .C(_03720_),
    .X(_03721_));
 sg13g2_o21ai_1 _25306_ (.B1(_03721_),
    .Y(_00519_),
    .A1(_04077_),
    .A2(_03687_));
 sg13g2_xnor2_1 _25307_ (.Y(_03722_),
    .A(_05439_),
    .B(_03363_));
 sg13g2_xnor2_1 _25308_ (.Y(_03723_),
    .A(net739),
    .B(_03722_));
 sg13g2_nand2_1 _25309_ (.Y(_03725_),
    .A(_03370_),
    .B(_03723_));
 sg13g2_nand2b_1 _25310_ (.Y(_03726_),
    .B(_03247_),
    .A_N(_05429_));
 sg13g2_nand2_1 _25311_ (.Y(_03727_),
    .A(net999),
    .B(net728));
 sg13g2_xnor2_1 _25312_ (.Y(_03728_),
    .A(net739),
    .B(net728));
 sg13g2_a21oi_1 _25313_ (.A1(net739),
    .A2(net728),
    .Y(_03729_),
    .B1(_05366_));
 sg13g2_a21oi_1 _25314_ (.A1(net347),
    .A2(_03728_),
    .Y(_03730_),
    .B1(_03729_));
 sg13g2_nand2_1 _25315_ (.Y(_03731_),
    .A(net401),
    .B(_03730_));
 sg13g2_o21ai_1 _25316_ (.B1(_03731_),
    .Y(_03732_),
    .A1(net1066),
    .A2(_03727_));
 sg13g2_nor4_1 _25317_ (.A(net339),
    .B(_05377_),
    .C(net740),
    .D(_03362_),
    .Y(_03733_));
 sg13g2_a21oi_1 _25318_ (.A1(net339),
    .A2(_03732_),
    .Y(_03734_),
    .B1(_03733_));
 sg13g2_o21ai_1 _25319_ (.B1(_03734_),
    .Y(_03736_),
    .A1(_03725_),
    .A2(_03726_));
 sg13g2_nand2_1 _25320_ (.Y(_03737_),
    .A(net403),
    .B(_05429_));
 sg13g2_xor2_1 _25321_ (.B(_03723_),
    .A(_03271_),
    .X(_03738_));
 sg13g2_nor2_1 _25322_ (.A(net403),
    .B(_05429_),
    .Y(_03739_));
 sg13g2_a221oi_1 _25323_ (.B2(_03738_),
    .C1(_03739_),
    .B1(_03737_),
    .A1(_03370_),
    .Y(_03740_),
    .A2(_03723_));
 sg13g2_inv_1 _25324_ (.Y(_03741_),
    .A(net738));
 sg13g2_nor2_1 _25325_ (.A(net665),
    .B(net728),
    .Y(_03742_));
 sg13g2_o21ai_1 _25326_ (.B1(_03742_),
    .Y(_03743_),
    .A1(net740),
    .A2(_03741_));
 sg13g2_nand3b_1 _25327_ (.B(net738),
    .C(_03742_),
    .Y(_03744_),
    .A_N(net657));
 sg13g2_o21ai_1 _25328_ (.B1(net392),
    .Y(_03745_),
    .A1(net657),
    .A2(_05367_));
 sg13g2_a22oi_1 _25329_ (.Y(_03747_),
    .B1(net740),
    .B2(net738),
    .A2(_05367_),
    .A1(net657));
 sg13g2_nand4_1 _25330_ (.B(_03744_),
    .C(_03745_),
    .A(net1066),
    .Y(_03748_),
    .D(_03747_));
 sg13g2_o21ai_1 _25331_ (.B1(_03748_),
    .Y(_03749_),
    .A1(net339),
    .A2(_03743_));
 sg13g2_xnor2_1 _25332_ (.Y(_03750_),
    .A(_03740_),
    .B(_03749_));
 sg13g2_o21ai_1 _25333_ (.B1(_05416_),
    .Y(_03751_),
    .A1(_03736_),
    .A2(_03750_));
 sg13g2_xor2_1 _25334_ (.B(_03723_),
    .A(_03633_),
    .X(_03752_));
 sg13g2_a21oi_1 _25335_ (.A1(net98),
    .A2(_03752_),
    .Y(_03753_),
    .B1(_03324_));
 sg13g2_nor2_1 _25336_ (.A(_03572_),
    .B(_03753_),
    .Y(_03754_));
 sg13g2_a22oi_1 _25337_ (.Y(_03755_),
    .B1(_03751_),
    .B2(_03754_),
    .A2(_03572_),
    .A1(_06621_));
 sg13g2_nor2_1 _25338_ (.A(net214),
    .B(_03755_),
    .Y(_00520_));
 sg13g2_xor2_1 _25339_ (.B(_03392_),
    .A(_05478_),
    .X(_03757_));
 sg13g2_xor2_1 _25340_ (.B(net1068),
    .A(_05418_),
    .X(_03758_));
 sg13g2_xnor2_1 _25341_ (.Y(_03759_),
    .A(_03757_),
    .B(_03758_));
 sg13g2_nor4_1 _25342_ (.A(_03403_),
    .B(_05473_),
    .C(_03303_),
    .D(_03759_),
    .Y(_03760_));
 sg13g2_nor2_1 _25343_ (.A(net996),
    .B(net727),
    .Y(_03761_));
 sg13g2_o21ai_1 _25344_ (.B1(_03761_),
    .Y(_03762_),
    .A1(_03741_),
    .A2(_02979_));
 sg13g2_nand3b_1 _25345_ (.B(_02990_),
    .C(_03761_),
    .Y(_03763_),
    .A_N(net654));
 sg13g2_o21ai_1 _25346_ (.B1(net391),
    .Y(_03764_),
    .A1(net654),
    .A2(net657));
 sg13g2_a22oi_1 _25347_ (.Y(_03765_),
    .B1(_03741_),
    .B2(net400),
    .A2(_05451_),
    .A1(net654));
 sg13g2_nand4_1 _25348_ (.B(_03763_),
    .C(_03764_),
    .A(_03037_),
    .Y(_03766_),
    .D(_03765_));
 sg13g2_o21ai_1 _25349_ (.B1(_03766_),
    .Y(_03768_),
    .A1(net343),
    .A2(_03762_));
 sg13g2_nand2_1 _25350_ (.Y(_03769_),
    .A(_05473_),
    .B(_02889_));
 sg13g2_xnor2_1 _25351_ (.Y(_03770_),
    .A(_03324_),
    .B(_03759_));
 sg13g2_nand2b_1 _25352_ (.Y(_03771_),
    .B(net402),
    .A_N(_05473_));
 sg13g2_o21ai_1 _25353_ (.B1(_03771_),
    .Y(_03772_),
    .A1(net1063),
    .A2(_03759_));
 sg13g2_a21oi_1 _25354_ (.A1(_03769_),
    .A2(_03770_),
    .Y(_03773_),
    .B1(_03772_));
 sg13g2_xnor2_1 _25355_ (.Y(_03774_),
    .A(_03768_),
    .B(_03773_));
 sg13g2_nand3_1 _25356_ (.B(net401),
    .C(_03418_),
    .A(net339),
    .Y(_03775_));
 sg13g2_nand2_1 _25357_ (.Y(_03776_),
    .A(net996),
    .B(net727));
 sg13g2_xor2_1 _25358_ (.B(net727),
    .A(_02939_),
    .X(_03777_));
 sg13g2_and2_1 _25359_ (.A(net996),
    .B(_03777_),
    .X(_03779_));
 sg13g2_nand2_1 _25360_ (.Y(_03780_),
    .A(net738),
    .B(net727));
 sg13g2_nor2_1 _25361_ (.A(_05451_),
    .B(_03780_),
    .Y(_03781_));
 sg13g2_o21ai_1 _25362_ (.B1(net400),
    .Y(_03782_),
    .A1(_03779_),
    .A2(_03781_));
 sg13g2_o21ai_1 _25363_ (.B1(_03782_),
    .Y(_03783_),
    .A1(_03037_),
    .A2(_03776_));
 sg13g2_nand2_1 _25364_ (.Y(_03784_),
    .A(net343),
    .B(_03783_));
 sg13g2_o21ai_1 _25365_ (.B1(_03784_),
    .Y(_03785_),
    .A1(net343),
    .A2(_03775_));
 sg13g2_nor3_1 _25366_ (.A(_03760_),
    .B(_03774_),
    .C(_03785_),
    .Y(_03786_));
 sg13g2_xnor2_1 _25367_ (.Y(_03787_),
    .A(_03700_),
    .B(_03759_));
 sg13g2_a21oi_1 _25368_ (.A1(_02820_),
    .A2(_03787_),
    .Y(_03788_),
    .B1(net392));
 sg13g2_nor2_1 _25369_ (.A(_03720_),
    .B(_03788_),
    .Y(_03790_));
 sg13g2_o21ai_1 _25370_ (.B1(_03790_),
    .Y(_03791_),
    .A1(_05472_),
    .A2(_03786_));
 sg13g2_o21ai_1 _25371_ (.B1(_03791_),
    .Y(_00521_),
    .A1(net29),
    .A2(_03687_));
 sg13g2_or2_1 _25372_ (.X(_03792_),
    .B(net726),
    .A(_05478_));
 sg13g2_buf_2 _25373_ (.A(_03792_),
    .X(_03793_));
 sg13g2_a21oi_1 _25374_ (.A1(net650),
    .A2(net737),
    .Y(_03794_),
    .B1(_03061_));
 sg13g2_nand2_1 _25375_ (.Y(_03795_),
    .A(net993),
    .B(net1067));
 sg13g2_a21oi_1 _25376_ (.A1(net399),
    .A2(_03795_),
    .Y(_03796_),
    .B1(net389));
 sg13g2_nand2_1 _25377_ (.Y(_03797_),
    .A(net1067),
    .B(net390));
 sg13g2_a21oi_1 _25378_ (.A1(net399),
    .A2(_03797_),
    .Y(_03798_),
    .B1(net654));
 sg13g2_o21ai_1 _25379_ (.B1(_05648_),
    .Y(_03800_),
    .A1(_03796_),
    .A2(_03798_));
 sg13g2_o21ai_1 _25380_ (.B1(_03800_),
    .Y(_03801_),
    .A1(_03793_),
    .A2(_03794_));
 sg13g2_a21oi_1 _25381_ (.A1(net400),
    .A2(_03064_),
    .Y(_03802_),
    .B1(_03793_));
 sg13g2_a22oi_1 _25382_ (.Y(_03803_),
    .B1(_03802_),
    .B2(_05648_),
    .A2(_03801_),
    .A1(_03080_));
 sg13g2_xor2_1 _25383_ (.B(_03040_),
    .A(_05538_),
    .X(_03804_));
 sg13g2_xnor2_1 _25384_ (.Y(_03805_),
    .A(net390),
    .B(_03804_));
 sg13g2_xor2_1 _25385_ (.B(_03805_),
    .A(net392),
    .X(_03806_));
 sg13g2_nand2b_1 _25386_ (.Y(_03807_),
    .B(_05546_),
    .A_N(net738));
 sg13g2_nor2b_1 _25387_ (.A(_05546_),
    .B_N(net401),
    .Y(_03808_));
 sg13g2_a221oi_1 _25388_ (.B2(_03807_),
    .C1(_03808_),
    .B1(_03806_),
    .A1(_03442_),
    .Y(_03809_),
    .A2(_03805_));
 sg13g2_xnor2_1 _25389_ (.Y(_03811_),
    .A(_03803_),
    .B(_03809_));
 sg13g2_and2_1 _25390_ (.A(_05502_),
    .B(net400),
    .X(_03812_));
 sg13g2_buf_1 _25391_ (.A(net337),
    .X(_03813_));
 sg13g2_nor2_1 _25392_ (.A(net131),
    .B(_03450_),
    .Y(_03814_));
 sg13g2_nand2_2 _25393_ (.Y(_03815_),
    .A(_05493_),
    .B(net389));
 sg13g2_xor2_1 _25394_ (.B(net390),
    .A(net737),
    .X(_03816_));
 sg13g2_nand2_1 _25395_ (.Y(_03817_),
    .A(_05497_),
    .B(_03816_));
 sg13g2_o21ai_1 _25396_ (.B1(_03817_),
    .Y(_03818_),
    .A1(_05502_),
    .A2(_03797_));
 sg13g2_nand2_1 _25397_ (.Y(_03819_),
    .A(net188),
    .B(_03818_));
 sg13g2_o21ai_1 _25398_ (.B1(_03819_),
    .Y(_03820_),
    .A1(_03080_),
    .A2(_03815_));
 sg13g2_nand2_1 _25399_ (.Y(_03822_),
    .A(_03442_),
    .B(_03805_));
 sg13g2_nor3_1 _25400_ (.A(_05546_),
    .B(_03363_),
    .C(_03822_),
    .Y(_03823_));
 sg13g2_a221oi_1 _25401_ (.B2(net131),
    .C1(_03823_),
    .B1(_03820_),
    .A1(_03812_),
    .Y(_03824_),
    .A2(_03814_));
 sg13g2_a21oi_1 _25402_ (.A1(_03811_),
    .A2(_03824_),
    .Y(_03825_),
    .B1(_10150_));
 sg13g2_xnor2_1 _25403_ (.Y(_03826_),
    .A(net339),
    .B(_03363_));
 sg13g2_xnor2_1 _25404_ (.Y(_03827_),
    .A(_03805_),
    .B(_03826_));
 sg13g2_a21oi_1 _25405_ (.A1(_08586_),
    .A2(_03827_),
    .Y(_03828_),
    .B1(net391));
 sg13g2_or3_1 _25406_ (.A(_03720_),
    .B(_03825_),
    .C(_03828_),
    .X(_03829_));
 sg13g2_o21ai_1 _25407_ (.B1(_03829_),
    .Y(_00522_),
    .A1(net43),
    .A2(_03687_));
 sg13g2_buf_1 _25408_ (.A(_00134_),
    .X(_03830_));
 sg13g2_o21ai_1 _25409_ (.B1(_03580_),
    .Y(_03832_),
    .A1(net337),
    .A2(_03610_));
 sg13g2_nor2_1 _25410_ (.A(net650),
    .B(_03580_),
    .Y(_03833_));
 sg13g2_a21oi_1 _25411_ (.A1(net1062),
    .A2(_03832_),
    .Y(_03834_),
    .B1(_03833_));
 sg13g2_nor2b_1 _25412_ (.A(net1062),
    .B_N(_03610_),
    .Y(_03835_));
 sg13g2_nor2_1 _25413_ (.A(_03110_),
    .B(_03610_),
    .Y(_03836_));
 sg13g2_o21ai_1 _25414_ (.B1(_03836_),
    .Y(_03837_),
    .A1(net1062),
    .A2(_03580_));
 sg13g2_nand2b_1 _25415_ (.Y(_03838_),
    .B(_03837_),
    .A_N(_03835_));
 sg13g2_nand2_1 _25416_ (.Y(_03839_),
    .A(net354),
    .B(_03223_));
 sg13g2_and2_1 _25417_ (.A(_05209_),
    .B(_02760_),
    .X(_03840_));
 sg13g2_buf_1 _25418_ (.A(_03840_),
    .X(_03841_));
 sg13g2_nor2b_1 _25419_ (.A(net650),
    .B_N(net1062),
    .Y(_03843_));
 sg13g2_o21ai_1 _25420_ (.B1(_03843_),
    .Y(_03844_),
    .A1(_03586_),
    .A2(_03841_));
 sg13g2_o21ai_1 _25421_ (.B1(_03844_),
    .Y(_03845_),
    .A1(net1062),
    .A2(_03839_));
 sg13g2_a21oi_1 _25422_ (.A1(_05580_),
    .A2(_03223_),
    .Y(_03846_),
    .B1(_03833_));
 sg13g2_nor2_1 _25423_ (.A(net188),
    .B(_03846_),
    .Y(_03847_));
 sg13g2_a221oi_1 _25424_ (.B2(_03091_),
    .C1(_03847_),
    .B1(_03845_),
    .A1(net131),
    .Y(_03848_),
    .A2(_03838_));
 sg13g2_o21ai_1 _25425_ (.B1(_03848_),
    .Y(_03849_),
    .A1(net95),
    .A2(_03834_));
 sg13g2_xor2_1 _25426_ (.B(net733),
    .A(net736),
    .X(_03850_));
 sg13g2_xnor2_1 _25427_ (.Y(_03851_),
    .A(_05202_),
    .B(_02759_));
 sg13g2_xnor2_1 _25428_ (.Y(_03852_),
    .A(net990),
    .B(_03851_));
 sg13g2_xnor2_1 _25429_ (.Y(_03854_),
    .A(_03850_),
    .B(_03852_));
 sg13g2_xnor2_1 _25430_ (.Y(_03855_),
    .A(net391),
    .B(_03854_));
 sg13g2_o21ai_1 _25431_ (.B1(_03855_),
    .Y(_03856_),
    .A1(_05576_),
    .A2(_02998_));
 sg13g2_nor2_1 _25432_ (.A(_03478_),
    .B(_03854_),
    .Y(_03857_));
 sg13g2_a21oi_1 _25433_ (.A1(_05576_),
    .A2(_02998_),
    .Y(_03858_),
    .B1(_03857_));
 sg13g2_nand2_1 _25434_ (.Y(_03859_),
    .A(_03856_),
    .B(_03858_));
 sg13g2_xnor2_1 _25435_ (.Y(_03860_),
    .A(_03849_),
    .B(_03859_));
 sg13g2_xnor2_1 _25436_ (.Y(_03861_),
    .A(_03757_),
    .B(_03854_));
 sg13g2_nor2_1 _25437_ (.A(_03460_),
    .B(_03861_),
    .Y(_03862_));
 sg13g2_nor4_1 _25438_ (.A(_03478_),
    .B(_05575_),
    .C(_03392_),
    .D(_03854_),
    .Y(_03863_));
 sg13g2_nand2_1 _25439_ (.Y(_03865_),
    .A(net188),
    .B(_03208_));
 sg13g2_nand2_1 _25440_ (.Y(_03866_),
    .A(net354),
    .B(_03850_));
 sg13g2_o21ai_1 _25441_ (.B1(_03866_),
    .Y(_03867_),
    .A1(net354),
    .A2(_03865_));
 sg13g2_a21oi_1 _25442_ (.A1(_03140_),
    .A2(_03867_),
    .Y(_03868_),
    .B1(_03835_));
 sg13g2_nor2b_1 _25443_ (.A(_03868_),
    .B_N(net131),
    .Y(_03869_));
 sg13g2_nand2b_1 _25444_ (.Y(_03870_),
    .B(_03610_),
    .A_N(_03110_));
 sg13g2_o21ai_1 _25445_ (.B1(_02776_),
    .Y(_03871_),
    .A1(net131),
    .A2(_03870_));
 sg13g2_nor4_1 _25446_ (.A(_03862_),
    .B(_03863_),
    .C(_03869_),
    .D(_03871_),
    .Y(_03872_));
 sg13g2_a22oi_1 _25447_ (.Y(_03873_),
    .B1(_03860_),
    .B2(_03872_),
    .A2(net74),
    .A1(_03460_));
 sg13g2_o21ai_1 _25448_ (.B1(net637),
    .Y(_03874_),
    .A1(net45),
    .A2(_03631_));
 sg13g2_a21oi_1 _25449_ (.A1(_03631_),
    .A2(_03873_),
    .Y(_00523_),
    .B1(_03874_));
 sg13g2_and2_1 _25450_ (.A(net676),
    .B(net390),
    .X(_03875_));
 sg13g2_buf_1 _25451_ (.A(_03875_),
    .X(_03876_));
 sg13g2_or2_1 _25452_ (.X(_03877_),
    .B(net726),
    .A(net676));
 sg13g2_buf_1 _25453_ (.A(_03877_),
    .X(_03878_));
 sg13g2_o21ai_1 _25454_ (.B1(_03878_),
    .Y(_03879_),
    .A1(net337),
    .A2(_03876_));
 sg13g2_nor2_1 _25455_ (.A(net337),
    .B(_03878_),
    .Y(_03880_));
 sg13g2_a21oi_1 _25456_ (.A1(net1062),
    .A2(_03879_),
    .Y(_03881_),
    .B1(_03880_));
 sg13g2_or2_1 _25457_ (.X(_03882_),
    .B(_03881_),
    .A(net95));
 sg13g2_nor2b_1 _25458_ (.A(net1062),
    .B_N(_03876_),
    .Y(_03883_));
 sg13g2_nor2_1 _25459_ (.A(_03830_),
    .B(_03878_),
    .Y(_03885_));
 sg13g2_nor3_1 _25460_ (.A(_03110_),
    .B(_03876_),
    .C(_03885_),
    .Y(_03886_));
 sg13g2_o21ai_1 _25461_ (.B1(_03813_),
    .Y(_03887_),
    .A1(_03883_),
    .A2(_03886_));
 sg13g2_and2_1 _25462_ (.A(_03459_),
    .B(_03063_),
    .X(_03888_));
 sg13g2_a21oi_1 _25463_ (.A1(_05580_),
    .A2(_03888_),
    .Y(_03889_),
    .B1(_03880_));
 sg13g2_a21o_1 _25464_ (.A2(_03459_),
    .A1(_03589_),
    .B1(_03841_),
    .X(_03890_));
 sg13g2_nor2_1 _25465_ (.A(net1062),
    .B(_03589_),
    .Y(_03891_));
 sg13g2_a22oi_1 _25466_ (.Y(_03892_),
    .B1(_03888_),
    .B2(_03891_),
    .A2(_03890_),
    .A1(_03843_));
 sg13g2_mux2_1 _25467_ (.A0(_03889_),
    .A1(_03892_),
    .S(net188),
    .X(_03893_));
 sg13g2_nand3_1 _25468_ (.B(_03887_),
    .C(_03893_),
    .A(_03882_),
    .Y(_03894_));
 sg13g2_xnor2_1 _25469_ (.Y(_03896_),
    .A(_03448_),
    .B(_03852_));
 sg13g2_xor2_1 _25470_ (.B(_03896_),
    .A(_03176_),
    .X(_03897_));
 sg13g2_nor2_1 _25471_ (.A(net743),
    .B(_05243_),
    .Y(_03898_));
 sg13g2_nor2_1 _25472_ (.A(_03184_),
    .B(_03896_),
    .Y(_03899_));
 sg13g2_a21oi_1 _25473_ (.A1(_02821_),
    .A2(_05243_),
    .Y(_03900_),
    .B1(_03899_));
 sg13g2_o21ai_1 _25474_ (.B1(_03900_),
    .Y(_03901_),
    .A1(_03897_),
    .A2(_03898_));
 sg13g2_xnor2_1 _25475_ (.Y(_03902_),
    .A(_03894_),
    .B(_03901_));
 sg13g2_nand2_1 _25476_ (.Y(_03903_),
    .A(net354),
    .B(_03448_));
 sg13g2_o21ai_1 _25477_ (.B1(_03903_),
    .Y(_03904_),
    .A1(net354),
    .A2(_03450_));
 sg13g2_a21o_1 _25478_ (.A2(_03904_),
    .A1(_03140_),
    .B1(_03883_),
    .X(_03905_));
 sg13g2_a221oi_1 _25479_ (.B2(_03813_),
    .C1(net115),
    .B1(_03905_),
    .A1(_03814_),
    .Y(_03907_),
    .A2(_03841_));
 sg13g2_xnor2_1 _25480_ (.Y(_03908_),
    .A(_02821_),
    .B(_03176_));
 sg13g2_nand3_1 _25481_ (.B(_03908_),
    .C(_03899_),
    .A(_05243_),
    .Y(_03909_));
 sg13g2_xnor2_1 _25482_ (.Y(_03910_),
    .A(_03625_),
    .B(_03897_));
 sg13g2_nand2_1 _25483_ (.Y(_03911_),
    .A(_03203_),
    .B(_03910_));
 sg13g2_nand4_1 _25484_ (.B(_03907_),
    .C(_03909_),
    .A(_03902_),
    .Y(_03912_),
    .D(_03911_));
 sg13g2_a22oi_1 _25485_ (.Y(_03913_),
    .B1(_06468_),
    .B2(_03630_),
    .A2(net74),
    .A1(net187));
 sg13g2_o21ai_1 _25486_ (.B1(_06118_),
    .Y(_03914_),
    .A1(_11347_),
    .A2(_03571_));
 sg13g2_a21oi_1 _25487_ (.A1(_03912_),
    .A2(_03913_),
    .Y(_00524_),
    .B1(_03914_));
 sg13g2_nor2_1 _25488_ (.A(net983),
    .B(_03589_),
    .Y(_03915_));
 sg13g2_nor3_1 _25489_ (.A(net351),
    .B(_05238_),
    .C(net336),
    .Y(_03917_));
 sg13g2_a21o_1 _25490_ (.A2(_05276_),
    .A1(net354),
    .B1(_03917_),
    .X(_03918_));
 sg13g2_a22oi_1 _25491_ (.Y(_03919_),
    .B1(_03918_),
    .B2(_05624_),
    .A2(_03915_),
    .A1(net184));
 sg13g2_nor2_1 _25492_ (.A(net395),
    .B(_03919_),
    .Y(_03920_));
 sg13g2_nand4_1 _25493_ (.B(net184),
    .C(_05624_),
    .A(net395),
    .Y(_03921_),
    .D(_05205_));
 sg13g2_o21ai_1 _25494_ (.B1(_02809_),
    .Y(_03922_),
    .A1(net352),
    .A2(_03921_));
 sg13g2_buf_2 _25495_ (.A(_00169_),
    .X(_03923_));
 sg13g2_inv_1 _25496_ (.Y(_03924_),
    .A(_03923_));
 sg13g2_xnor2_1 _25497_ (.Y(_03925_),
    .A(_03168_),
    .B(_05226_));
 sg13g2_xnor2_1 _25498_ (.Y(_03926_),
    .A(_05222_),
    .B(_03925_));
 sg13g2_xnor2_1 _25499_ (.Y(_03928_),
    .A(_05189_),
    .B(_03926_));
 sg13g2_xnor2_1 _25500_ (.Y(_03929_),
    .A(net735),
    .B(_05172_));
 sg13g2_and4_1 _25501_ (.A(_03924_),
    .B(net730),
    .C(_03928_),
    .D(_03929_),
    .X(_03930_));
 sg13g2_nand2_1 _25502_ (.Y(_03931_),
    .A(net671),
    .B(_03923_));
 sg13g2_xor2_1 _25503_ (.B(_03928_),
    .A(net735),
    .X(_03932_));
 sg13g2_nor2_1 _25504_ (.A(net671),
    .B(_03923_),
    .Y(_03933_));
 sg13g2_a221oi_1 _25505_ (.B2(_03932_),
    .C1(_03933_),
    .B1(_03931_),
    .A1(net730),
    .Y(_03934_),
    .A2(_03928_));
 sg13g2_nor2_1 _25506_ (.A(net675),
    .B(net676),
    .Y(_03935_));
 sg13g2_nand3_1 _25507_ (.B(net1014),
    .C(_03935_),
    .A(net395),
    .Y(_03936_));
 sg13g2_nand4_1 _25508_ (.B(_05190_),
    .C(net983),
    .A(net732),
    .Y(_03937_),
    .D(net677));
 sg13g2_nand2_1 _25509_ (.Y(_03939_),
    .A(_03936_),
    .B(_03937_));
 sg13g2_mux2_1 _25510_ (.A0(_05703_),
    .A1(_05195_),
    .S(net1013),
    .X(_03940_));
 sg13g2_nor2_1 _25511_ (.A(_05249_),
    .B(_03940_),
    .Y(_03941_));
 sg13g2_a21oi_1 _25512_ (.A1(_05250_),
    .A2(_03915_),
    .Y(_03942_),
    .B1(_03941_));
 sg13g2_o21ai_1 _25513_ (.B1(_03942_),
    .Y(_03943_),
    .A1(_05720_),
    .A2(_03935_));
 sg13g2_nand2b_1 _25514_ (.Y(_03944_),
    .B(net676),
    .A_N(_05703_));
 sg13g2_mux2_1 _25515_ (.A0(net677),
    .A1(_03944_),
    .S(net675),
    .X(_03945_));
 sg13g2_nand2b_1 _25516_ (.Y(_03946_),
    .B(net1014),
    .A_N(_05210_));
 sg13g2_a21oi_1 _25517_ (.A1(_05211_),
    .A2(_03946_),
    .Y(_03947_),
    .B1(net1009));
 sg13g2_a221oi_1 _25518_ (.B2(net678),
    .C1(_03947_),
    .B1(_03945_),
    .A1(_05711_),
    .Y(_03948_),
    .A2(_03935_));
 sg13g2_nor2_1 _25519_ (.A(net395),
    .B(_03948_),
    .Y(_03950_));
 sg13g2_a221oi_1 _25520_ (.B2(_03232_),
    .C1(_03950_),
    .B1(_03943_),
    .A1(net662),
    .Y(_03951_),
    .A2(_03939_));
 sg13g2_xnor2_1 _25521_ (.Y(_03952_),
    .A(_03934_),
    .B(_03951_));
 sg13g2_nor4_1 _25522_ (.A(_03920_),
    .B(_03922_),
    .C(_03930_),
    .D(_03952_),
    .Y(_03953_));
 sg13g2_nor2_1 _25523_ (.A(_05182_),
    .B(_06474_),
    .Y(_03954_));
 sg13g2_buf_1 _25524_ (.A(_03954_),
    .X(_03955_));
 sg13g2_nor2b_1 _25525_ (.A(net51),
    .B_N(net672),
    .Y(_03956_));
 sg13g2_o21ai_1 _25526_ (.B1(_03956_),
    .Y(_03957_),
    .A1(net75),
    .A2(_03953_));
 sg13g2_xnor2_1 _25527_ (.Y(_03958_),
    .A(net187),
    .B(_03929_));
 sg13g2_xnor2_1 _25528_ (.Y(_03959_),
    .A(_03928_),
    .B(_03958_));
 sg13g2_nor2_1 _25529_ (.A(net51),
    .B(_03959_),
    .Y(_03961_));
 sg13g2_a22oi_1 _25530_ (.Y(_03962_),
    .B1(_03953_),
    .B2(_03961_),
    .A2(_03955_),
    .A1(_01806_));
 sg13g2_a21oi_1 _25531_ (.A1(_03957_),
    .A2(_03962_),
    .Y(_00525_),
    .B1(net440));
 sg13g2_xor2_1 _25532_ (.B(net348),
    .A(net1009),
    .X(_03963_));
 sg13g2_nor3_1 _25533_ (.A(net396),
    .B(_05239_),
    .C(net349),
    .Y(_03964_));
 sg13g2_a21oi_1 _25534_ (.A1(net396),
    .A2(_03963_),
    .Y(_03965_),
    .B1(_03964_));
 sg13g2_nand3_1 _25535_ (.B(net669),
    .C(_05711_),
    .A(_03168_),
    .Y(_03966_));
 sg13g2_o21ai_1 _25536_ (.B1(_03966_),
    .Y(_03967_),
    .A1(net345),
    .A2(_03965_));
 sg13g2_nor3_1 _25537_ (.A(net672),
    .B(_03232_),
    .C(_05303_),
    .Y(_03968_));
 sg13g2_a22oi_1 _25538_ (.Y(_03969_),
    .B1(_03968_),
    .B2(net662),
    .A2(_03967_),
    .A1(net672));
 sg13g2_xor2_1 _25539_ (.B(_03925_),
    .A(_05298_),
    .X(_03971_));
 sg13g2_xnor2_1 _25540_ (.Y(_03972_),
    .A(_03173_),
    .B(_05349_));
 sg13g2_xnor2_1 _25541_ (.Y(_03973_),
    .A(_03971_),
    .B(_03972_));
 sg13g2_nor2_1 _25542_ (.A(_03345_),
    .B(_03973_),
    .Y(_03974_));
 sg13g2_nand2_1 _25543_ (.Y(_03975_),
    .A(_03231_),
    .B(net349));
 sg13g2_nand2b_1 _25544_ (.Y(_03976_),
    .B(net1004),
    .A_N(net1006));
 sg13g2_nand4_1 _25545_ (.B(net732),
    .C(net669),
    .A(net1006),
    .Y(_03977_),
    .D(net983));
 sg13g2_o21ai_1 _25546_ (.B1(_03977_),
    .Y(_03978_),
    .A1(_03975_),
    .A2(_03976_));
 sg13g2_mux2_1 _25547_ (.A0(net349),
    .A1(_05307_),
    .S(_03231_),
    .X(_03979_));
 sg13g2_nand2_1 _25548_ (.Y(_03980_),
    .A(_05238_),
    .B(_03979_));
 sg13g2_nand3_1 _25549_ (.B(_03966_),
    .C(_03975_),
    .A(_05426_),
    .Y(_03982_));
 sg13g2_nand2b_1 _25550_ (.Y(_03983_),
    .B(_05711_),
    .A_N(_03975_));
 sg13g2_nand3_1 _25551_ (.B(_03982_),
    .C(_03983_),
    .A(_03980_),
    .Y(_03984_));
 sg13g2_nand2_1 _25552_ (.Y(_03985_),
    .A(net349),
    .B(_05704_));
 sg13g2_nand3_1 _25553_ (.B(_05303_),
    .C(_03985_),
    .A(net732),
    .Y(_03986_));
 sg13g2_nor2_1 _25554_ (.A(_05227_),
    .B(_05321_),
    .Y(_03987_));
 sg13g2_nor3_1 _25555_ (.A(_03201_),
    .B(net349),
    .C(_05704_),
    .Y(_03988_));
 sg13g2_a21oi_1 _25556_ (.A1(_03975_),
    .A2(_03987_),
    .Y(_03989_),
    .B1(_03988_));
 sg13g2_a21oi_1 _25557_ (.A1(_03986_),
    .A2(_03989_),
    .Y(_03990_),
    .B1(net1006));
 sg13g2_a221oi_1 _25558_ (.B2(net672),
    .C1(_03990_),
    .B1(_03984_),
    .A1(net662),
    .Y(_03991_),
    .A2(_03978_));
 sg13g2_xnor2_1 _25559_ (.Y(_03993_),
    .A(net1006),
    .B(_03971_));
 sg13g2_nand2_1 _25560_ (.Y(_03994_),
    .A(net735),
    .B(net1017));
 sg13g2_o21ai_1 _25561_ (.B1(_03183_),
    .Y(_03995_),
    .A1(net735),
    .A2(net671));
 sg13g2_nor2_1 _25562_ (.A(_03995_),
    .B(_03993_),
    .Y(_03996_));
 sg13g2_a21oi_1 _25563_ (.A1(_03993_),
    .A2(_03994_),
    .Y(_03997_),
    .B1(_03996_));
 sg13g2_xor2_1 _25564_ (.B(_03997_),
    .A(_03991_),
    .X(_03998_));
 sg13g2_nand3b_1 _25565_ (.B(_03991_),
    .C(_03974_),
    .Y(_03999_),
    .A_N(_03997_));
 sg13g2_o21ai_1 _25566_ (.B1(_03999_),
    .Y(_04000_),
    .A1(_03974_),
    .A2(_03998_));
 sg13g2_a21oi_1 _25567_ (.A1(_03969_),
    .A2(_04000_),
    .Y(_04001_),
    .B1(net79));
 sg13g2_xnor2_1 _25568_ (.Y(_04002_),
    .A(net186),
    .B(_03973_));
 sg13g2_a21oi_1 _25569_ (.A1(net112),
    .A2(_04002_),
    .Y(_04004_),
    .B1(net184));
 sg13g2_o21ai_1 _25570_ (.B1(net1197),
    .Y(_04005_),
    .A1(_05182_),
    .A2(_06474_));
 sg13g2_buf_1 _25571_ (.A(_04005_),
    .X(_04006_));
 sg13g2_or2_1 _25572_ (.X(_04007_),
    .B(_04006_),
    .A(_04004_));
 sg13g2_nand2_1 _25573_ (.Y(_04008_),
    .A(net1060),
    .B(net51));
 sg13g2_nand2b_1 _25574_ (.Y(_04009_),
    .B(_07276_),
    .A_N(_04008_));
 sg13g2_o21ai_1 _25575_ (.B1(_04009_),
    .Y(_00526_),
    .A1(_04001_),
    .A2(_04007_));
 sg13g2_nor2_1 _25576_ (.A(net731),
    .B(_05365_),
    .Y(_04010_));
 sg13g2_nand2_1 _25577_ (.Y(_04011_),
    .A(_05362_),
    .B(_04010_));
 sg13g2_a22oi_1 _25578_ (.Y(_04012_),
    .B1(net665),
    .B2(net394),
    .A2(_05362_),
    .A1(_05321_));
 sg13g2_and2_1 _25579_ (.A(_04011_),
    .B(_04012_),
    .X(_04014_));
 sg13g2_a22oi_1 _25580_ (.Y(_04015_),
    .B1(_04014_),
    .B2(net1176),
    .A2(_04010_),
    .A1(_05842_));
 sg13g2_o21ai_1 _25581_ (.B1(_05363_),
    .Y(_04016_),
    .A1(net351),
    .A2(_05426_));
 sg13g2_nand3_1 _25582_ (.B(_04016_),
    .C(_04010_),
    .A(_05310_),
    .Y(_04017_));
 sg13g2_o21ai_1 _25583_ (.B1(_04017_),
    .Y(_04018_),
    .A1(net184),
    .A2(_04015_));
 sg13g2_nand2_1 _25584_ (.Y(_04019_),
    .A(net352),
    .B(net1063));
 sg13g2_xnor2_1 _25585_ (.Y(_04020_),
    .A(_03246_),
    .B(_05284_));
 sg13g2_xor2_1 _25586_ (.B(_04020_),
    .A(_05369_),
    .X(_04021_));
 sg13g2_xnor2_1 _25587_ (.Y(_04022_),
    .A(_05249_),
    .B(_04021_));
 sg13g2_xnor2_1 _25588_ (.Y(_04023_),
    .A(net396),
    .B(_04022_));
 sg13g2_nand2b_1 _25589_ (.Y(_04025_),
    .B(net1009),
    .A_N(_00041_));
 sg13g2_o21ai_1 _25590_ (.B1(_04025_),
    .Y(_04026_),
    .A1(_03336_),
    .A2(_04022_));
 sg13g2_a21oi_1 _25591_ (.A1(_04019_),
    .A2(_04023_),
    .Y(_04027_),
    .B1(_04026_));
 sg13g2_xnor2_1 _25592_ (.Y(_04028_),
    .A(_04018_),
    .B(_04027_));
 sg13g2_nand2_1 _25593_ (.Y(_04029_),
    .A(net661),
    .B(net347));
 sg13g2_xor2_1 _25594_ (.B(net665),
    .A(_05411_),
    .X(_04030_));
 sg13g2_nand2_1 _25595_ (.Y(_04031_),
    .A(net186),
    .B(_04030_));
 sg13g2_o21ai_1 _25596_ (.B1(_04031_),
    .Y(_04032_),
    .A1(net186),
    .A2(_04029_));
 sg13g2_nor2b_1 _25597_ (.A(_05310_),
    .B_N(net186),
    .Y(_04033_));
 sg13g2_a22oi_1 _25598_ (.Y(_04034_),
    .B1(_04033_),
    .B2(net347),
    .A2(_04032_),
    .A1(_05363_));
 sg13g2_nor2_1 _25599_ (.A(net351),
    .B(_04034_),
    .Y(_04036_));
 sg13g2_nand2_1 _25600_ (.Y(_04037_),
    .A(_03271_),
    .B(_05411_));
 sg13g2_nor3_1 _25601_ (.A(net184),
    .B(_05371_),
    .C(_04037_),
    .Y(_04038_));
 sg13g2_nand2b_1 _25602_ (.Y(_04039_),
    .B(_03925_),
    .A_N(net1063));
 sg13g2_nor3_1 _25603_ (.A(_03336_),
    .B(_04022_),
    .C(_04039_),
    .Y(_04040_));
 sg13g2_nor4_1 _25604_ (.A(_04028_),
    .B(_04036_),
    .C(_04038_),
    .D(_04040_),
    .Y(_04041_));
 sg13g2_xnor2_1 _25605_ (.Y(_04042_),
    .A(net393),
    .B(_03925_));
 sg13g2_xnor2_1 _25606_ (.Y(_04043_),
    .A(_04022_),
    .B(_04042_));
 sg13g2_a21oi_1 _25607_ (.A1(net126),
    .A2(_04043_),
    .Y(_04044_),
    .B1(net348));
 sg13g2_nor2_1 _25608_ (.A(_04006_),
    .B(_04044_),
    .Y(_04045_));
 sg13g2_o21ai_1 _25609_ (.B1(_04045_),
    .Y(_04047_),
    .A1(_05737_),
    .A2(_04041_));
 sg13g2_o21ai_1 _25610_ (.B1(_04047_),
    .Y(_00527_),
    .A1(net35),
    .A2(_04008_));
 sg13g2_xnor2_1 _25611_ (.Y(_04048_),
    .A(_05287_),
    .B(_05418_));
 sg13g2_xor2_1 _25612_ (.B(_04048_),
    .A(net729),
    .X(_04049_));
 sg13g2_o21ai_1 _25613_ (.B1(_05379_),
    .Y(_04050_),
    .A1(_05445_),
    .A2(net666));
 sg13g2_nand2_1 _25614_ (.Y(_04051_),
    .A(_05879_),
    .B(_04049_));
 sg13g2_o21ai_1 _25615_ (.B1(_04051_),
    .Y(_04052_),
    .A1(_04049_),
    .A2(_04050_));
 sg13g2_xnor2_1 _25616_ (.Y(_04053_),
    .A(_05361_),
    .B(_03300_));
 sg13g2_xnor2_1 _25617_ (.Y(_04054_),
    .A(_04048_),
    .B(_04053_));
 sg13g2_xnor2_1 _25618_ (.Y(_04055_),
    .A(net997),
    .B(_04054_));
 sg13g2_nand2_1 _25619_ (.Y(_04057_),
    .A(net345),
    .B(_03434_));
 sg13g2_xor2_1 _25620_ (.B(_04055_),
    .A(net394),
    .X(_04058_));
 sg13g2_nor2_1 _25621_ (.A(net345),
    .B(_03434_),
    .Y(_04059_));
 sg13g2_a221oi_1 _25622_ (.B2(_04058_),
    .C1(_04059_),
    .B1(_04057_),
    .A1(_03370_),
    .Y(_04060_),
    .A2(_04055_));
 sg13g2_and2_1 _25623_ (.A(_04052_),
    .B(_04060_),
    .X(_04061_));
 sg13g2_nand4_1 _25624_ (.B(_03370_),
    .C(_04020_),
    .A(_03442_),
    .Y(_04062_),
    .D(_04055_));
 sg13g2_o21ai_1 _25625_ (.B1(_04062_),
    .Y(_04063_),
    .A1(_04052_),
    .A2(_04060_));
 sg13g2_nor2_1 _25626_ (.A(net339),
    .B(net393),
    .Y(_04064_));
 sg13g2_a21oi_1 _25627_ (.A1(net339),
    .A2(net393),
    .Y(_04065_),
    .B1(net348));
 sg13g2_nor2_1 _25628_ (.A(_04064_),
    .B(_04065_),
    .Y(_04066_));
 sg13g2_nor2_1 _25629_ (.A(_03831_),
    .B(_04066_),
    .Y(_04068_));
 sg13g2_o21ai_1 _25630_ (.B1(_04068_),
    .Y(_04069_),
    .A1(_04061_),
    .A2(_04063_));
 sg13g2_xnor2_1 _25631_ (.Y(_04070_),
    .A(net392),
    .B(_04020_));
 sg13g2_xnor2_1 _25632_ (.Y(_04071_),
    .A(_04055_),
    .B(_04070_));
 sg13g2_o21ai_1 _25633_ (.B1(_05377_),
    .Y(_04072_),
    .A1(_05408_),
    .A2(_04071_));
 sg13g2_nand3b_1 _25634_ (.B(_04066_),
    .C(_04650_),
    .Y(_04073_),
    .A_N(_04061_));
 sg13g2_nand3_1 _25635_ (.B(_04072_),
    .C(_04073_),
    .A(_04069_),
    .Y(_04074_));
 sg13g2_or2_1 _25636_ (.X(_04075_),
    .B(_04008_),
    .A(_05863_));
 sg13g2_o21ai_1 _25637_ (.B1(_04075_),
    .Y(_00528_),
    .A1(_04006_),
    .A2(_04074_));
 sg13g2_nand3_1 _25638_ (.B(net347),
    .C(net728),
    .A(net343),
    .Y(_04076_));
 sg13g2_xor2_1 _25639_ (.B(_03348_),
    .A(net999),
    .X(_04078_));
 sg13g2_nand2_1 _25640_ (.Y(_04079_),
    .A(net654),
    .B(_04078_));
 sg13g2_o21ai_1 _25641_ (.B1(_04079_),
    .Y(_04080_),
    .A1(net654),
    .A2(_03727_));
 sg13g2_nand2_1 _25642_ (.Y(_04081_),
    .A(net658),
    .B(_04080_));
 sg13g2_o21ai_1 _25643_ (.B1(_04081_),
    .Y(_04082_),
    .A1(net658),
    .A2(_04076_));
 sg13g2_xnor2_1 _25644_ (.Y(_04083_),
    .A(_05420_),
    .B(_03348_));
 sg13g2_xor2_1 _25645_ (.B(_04083_),
    .A(_05479_),
    .X(_04084_));
 sg13g2_xnor2_1 _25646_ (.Y(_04085_),
    .A(_05377_),
    .B(_04084_));
 sg13g2_nor2_1 _25647_ (.A(_03403_),
    .B(_04085_),
    .Y(_04086_));
 sg13g2_and2_1 _25648_ (.A(_03479_),
    .B(_04053_),
    .X(_04087_));
 sg13g2_nor2_1 _25649_ (.A(_05434_),
    .B(_04076_),
    .Y(_04089_));
 sg13g2_a221oi_1 _25650_ (.B2(_04087_),
    .C1(_04089_),
    .B1(_04086_),
    .A1(net342),
    .Y(_04090_),
    .A2(_04082_));
 sg13g2_nand2_1 _25651_ (.Y(_04091_),
    .A(_03478_),
    .B(_05391_));
 sg13g2_xnor2_1 _25652_ (.Y(_04092_),
    .A(net393),
    .B(_04085_));
 sg13g2_nand2_1 _25653_ (.Y(_04093_),
    .A(_03479_),
    .B(net666));
 sg13g2_o21ai_1 _25654_ (.B1(_04093_),
    .Y(_04094_),
    .A1(net1063),
    .A2(_04085_));
 sg13g2_a21oi_1 _25655_ (.A1(_04091_),
    .A2(_04092_),
    .Y(_04095_),
    .B1(_04094_));
 sg13g2_a22oi_1 _25656_ (.Y(_04096_),
    .B1(_04078_),
    .B2(_05438_),
    .A2(_03727_),
    .A1(_05604_));
 sg13g2_and2_1 _25657_ (.A(_05438_),
    .B(_05497_),
    .X(_04097_));
 sg13g2_o21ai_1 _25658_ (.B1(_03742_),
    .Y(_04098_),
    .A1(_05604_),
    .A2(_04097_));
 sg13g2_o21ai_1 _25659_ (.B1(_04098_),
    .Y(_04100_),
    .A1(net343),
    .A2(_04096_));
 sg13g2_nor3_1 _25660_ (.A(net343),
    .B(net347),
    .C(_03372_),
    .Y(_04101_));
 sg13g2_a22oi_1 _25661_ (.Y(_04102_),
    .B1(_04101_),
    .B2(_05918_),
    .A2(_04100_),
    .A1(_05434_));
 sg13g2_xnor2_1 _25662_ (.Y(_04103_),
    .A(_04095_),
    .B(_04102_));
 sg13g2_a21oi_1 _25663_ (.A1(_04090_),
    .A2(_04103_),
    .Y(_04104_),
    .B1(_10150_));
 sg13g2_xnor2_1 _25664_ (.Y(_04105_),
    .A(net391),
    .B(_04053_));
 sg13g2_xnor2_1 _25665_ (.Y(_04106_),
    .A(_04085_),
    .B(_04105_));
 sg13g2_a21oi_1 _25666_ (.A1(_08586_),
    .A2(_04106_),
    .Y(_04107_),
    .B1(net339));
 sg13g2_or3_1 _25667_ (.A(_04006_),
    .B(_04104_),
    .C(_04107_),
    .X(_04108_));
 sg13g2_o21ai_1 _25668_ (.B1(_04108_),
    .Y(_00529_),
    .A1(_04941_),
    .A2(_04008_));
 sg13g2_nand3_1 _25669_ (.B(net657),
    .C(_03447_),
    .A(net337),
    .Y(_04110_));
 sg13g2_xor2_1 _25670_ (.B(_03391_),
    .A(_05442_),
    .X(_04111_));
 sg13g2_and2_1 _25671_ (.A(net337),
    .B(_04111_),
    .X(_04112_));
 sg13g2_nor2_1 _25672_ (.A(net337),
    .B(_03776_),
    .Y(_04113_));
 sg13g2_o21ai_1 _25673_ (.B1(net342),
    .Y(_04114_),
    .A1(_04112_),
    .A2(_04113_));
 sg13g2_o21ai_1 _25674_ (.B1(_04114_),
    .Y(_04115_),
    .A1(net342),
    .A2(_04110_));
 sg13g2_xnor2_1 _25675_ (.Y(_04116_),
    .A(_05477_),
    .B(net1064));
 sg13g2_xnor2_1 _25676_ (.Y(_04117_),
    .A(_05638_),
    .B(_04116_));
 sg13g2_xnor2_1 _25677_ (.Y(_04118_),
    .A(_05442_),
    .B(_04117_));
 sg13g2_nor2_1 _25678_ (.A(_03434_),
    .B(_04118_),
    .Y(_04119_));
 sg13g2_buf_1 _25679_ (.A(_00137_),
    .X(_04121_));
 sg13g2_nor2b_1 _25680_ (.A(_04121_),
    .B_N(_04083_),
    .Y(_04122_));
 sg13g2_nor2_1 _25681_ (.A(_05488_),
    .B(_04110_),
    .Y(_04123_));
 sg13g2_a221oi_1 _25682_ (.B2(_04122_),
    .C1(_04123_),
    .B1(_04119_),
    .A1(net340),
    .Y(_04124_),
    .A2(_04115_));
 sg13g2_nand2_1 _25683_ (.Y(_04125_),
    .A(_04121_),
    .B(_05445_));
 sg13g2_xnor2_1 _25684_ (.Y(_04126_),
    .A(_03372_),
    .B(_04118_));
 sg13g2_nand2b_1 _25685_ (.Y(_04127_),
    .B(net658),
    .A_N(_04121_));
 sg13g2_o21ai_1 _25686_ (.B1(_04127_),
    .Y(_04128_),
    .A1(_03434_),
    .A2(_04118_));
 sg13g2_a21oi_1 _25687_ (.A1(_04125_),
    .A2(_04126_),
    .Y(_04129_),
    .B1(_04128_));
 sg13g2_a22oi_1 _25688_ (.Y(_04130_),
    .B1(_04111_),
    .B2(_05492_),
    .A2(_03776_),
    .A1(net649));
 sg13g2_and2_1 _25689_ (.A(_05491_),
    .B(net650),
    .X(_04132_));
 sg13g2_o21ai_1 _25690_ (.B1(_03761_),
    .Y(_04133_),
    .A1(net649),
    .A2(_04132_));
 sg13g2_o21ai_1 _25691_ (.B1(_04133_),
    .Y(_04134_),
    .A1(net131),
    .A2(_04130_));
 sg13g2_nor3_1 _25692_ (.A(net131),
    .B(_05568_),
    .C(_03447_),
    .Y(_04135_));
 sg13g2_a22oi_1 _25693_ (.Y(_04136_),
    .B1(_04135_),
    .B2(_05954_),
    .A2(_04134_),
    .A1(_05488_));
 sg13g2_xnor2_1 _25694_ (.Y(_04137_),
    .A(_04129_),
    .B(_04136_));
 sg13g2_a21o_1 _25695_ (.A2(_04137_),
    .A1(_04124_),
    .B1(net103),
    .X(_04138_));
 sg13g2_xnor2_1 _25696_ (.Y(_04139_),
    .A(net185),
    .B(_04083_));
 sg13g2_xnor2_1 _25697_ (.Y(_04140_),
    .A(_04118_),
    .B(_04139_));
 sg13g2_a21oi_1 _25698_ (.A1(_08549_),
    .A2(_04140_),
    .Y(_04141_),
    .B1(net343));
 sg13g2_nor2_1 _25699_ (.A(net51),
    .B(_04141_),
    .Y(_04143_));
 sg13g2_a22oi_1 _25700_ (.Y(_04144_),
    .B1(_04138_),
    .B2(_04143_),
    .A2(net51),
    .A1(_06330_));
 sg13g2_nor2_1 _25701_ (.A(_12651_),
    .B(_04144_),
    .Y(_00530_));
 sg13g2_nor2_1 _25702_ (.A(net677),
    .B(_03793_),
    .Y(_04145_));
 sg13g2_xnor2_1 _25703_ (.Y(_04146_),
    .A(_05478_),
    .B(_03436_));
 sg13g2_a21o_1 _25704_ (.A2(net390),
    .A1(net993),
    .B1(net1014),
    .X(_04147_));
 sg13g2_o21ai_1 _25705_ (.B1(_04147_),
    .Y(_04148_),
    .A1(net649),
    .A2(_04146_));
 sg13g2_nand2_1 _25706_ (.Y(_04149_),
    .A(_05536_),
    .B(net677));
 sg13g2_a21oi_1 _25707_ (.A1(_05196_),
    .A2(_04149_),
    .Y(_04150_),
    .B1(_03793_));
 sg13g2_a21o_1 _25708_ (.A2(_04148_),
    .A1(_03589_),
    .B1(_04150_),
    .X(_04151_));
 sg13g2_a22oi_1 _25709_ (.Y(_04153_),
    .B1(_04151_),
    .B2(net652),
    .A2(_04145_),
    .A1(_05989_));
 sg13g2_xor2_1 _25710_ (.B(net336),
    .A(net991),
    .X(_04154_));
 sg13g2_nand3_1 _25711_ (.B(net336),
    .C(_03815_),
    .A(net991),
    .Y(_04155_));
 sg13g2_o21ai_1 _25712_ (.B1(_04155_),
    .Y(_04156_),
    .A1(net652),
    .A2(_03815_));
 sg13g2_a21oi_1 _25713_ (.A1(_03793_),
    .A2(_04154_),
    .Y(_04157_),
    .B1(_04156_));
 sg13g2_and2_1 _25714_ (.A(_05493_),
    .B(_03453_),
    .X(_04158_));
 sg13g2_nand3_1 _25715_ (.B(_05627_),
    .C(_04158_),
    .A(_05196_),
    .Y(_04159_));
 sg13g2_o21ai_1 _25716_ (.B1(_04159_),
    .Y(_04160_),
    .A1(_05627_),
    .A2(_03793_));
 sg13g2_o21ai_1 _25717_ (.B1(_03793_),
    .Y(_04161_),
    .A1(net677),
    .A2(_04158_));
 sg13g2_a21o_1 _25718_ (.A2(_04161_),
    .A1(net991),
    .B1(_04145_),
    .X(_04162_));
 sg13g2_nor3_1 _25719_ (.A(net652),
    .B(_03589_),
    .C(_03815_),
    .Y(_04164_));
 sg13g2_a221oi_1 _25720_ (.B2(net678),
    .C1(_04164_),
    .B1(_04162_),
    .A1(net649),
    .Y(_04165_),
    .A2(_04160_));
 sg13g2_o21ai_1 _25721_ (.B1(_04165_),
    .Y(_04166_),
    .A1(_05989_),
    .A2(_04157_));
 sg13g2_and2_1 _25722_ (.A(net994),
    .B(net727),
    .X(_04167_));
 sg13g2_nor2_1 _25723_ (.A(_05604_),
    .B(_03395_),
    .Y(_04168_));
 sg13g2_xnor2_1 _25724_ (.Y(_04169_),
    .A(_05222_),
    .B(_04146_));
 sg13g2_xnor2_1 _25725_ (.Y(_04170_),
    .A(net989),
    .B(_04169_));
 sg13g2_mux2_1 _25726_ (.A0(_04167_),
    .A1(_04168_),
    .S(_04170_),
    .X(_04171_));
 sg13g2_and2_1 _25727_ (.A(_03479_),
    .B(_04170_),
    .X(_04172_));
 sg13g2_nor2_1 _25728_ (.A(_04171_),
    .B(_04172_),
    .Y(_04173_));
 sg13g2_mux2_1 _25729_ (.A0(_04153_),
    .A1(_04166_),
    .S(_04173_),
    .X(_04175_));
 sg13g2_xnor2_1 _25730_ (.Y(_04176_),
    .A(_04116_),
    .B(_04170_));
 sg13g2_and2_1 _25731_ (.A(_03924_),
    .B(_04176_),
    .X(_04177_));
 sg13g2_nor3_1 _25732_ (.A(_04171_),
    .B(_04172_),
    .C(_04153_),
    .Y(_04178_));
 sg13g2_a21oi_1 _25733_ (.A1(_04177_),
    .A2(_04178_),
    .Y(_04179_),
    .B1(net99));
 sg13g2_o21ai_1 _25734_ (.B1(_04179_),
    .Y(_04180_),
    .A1(_04175_),
    .A2(_04177_));
 sg13g2_xnor2_1 _25735_ (.Y(_04181_),
    .A(_03203_),
    .B(_04176_));
 sg13g2_a21oi_1 _25736_ (.A1(_08549_),
    .A2(_04181_),
    .Y(_04182_),
    .B1(net131));
 sg13g2_nor2_1 _25737_ (.A(net51),
    .B(_04182_),
    .Y(_04183_));
 sg13g2_a22oi_1 _25738_ (.Y(_04184_),
    .B1(_04180_),
    .B2(_04183_),
    .A2(net51),
    .A1(_06019_));
 sg13g2_nor2_1 _25739_ (.A(_12651_),
    .B(_04184_),
    .Y(_00531_));
 sg13g2_xnor2_1 _25740_ (.Y(_04186_),
    .A(_05195_),
    .B(_03436_));
 sg13g2_xnor2_1 _25741_ (.Y(_04187_),
    .A(_05638_),
    .B(_04186_));
 sg13g2_xnor2_1 _25742_ (.Y(_04188_),
    .A(_05273_),
    .B(_04187_));
 sg13g2_buf_1 _25743_ (.A(_04188_),
    .X(_04189_));
 sg13g2_a21oi_1 _25744_ (.A1(net671),
    .A2(net730),
    .Y(_04190_),
    .B1(_04189_));
 sg13g2_nand2_1 _25745_ (.Y(_04191_),
    .A(net398),
    .B(_04190_));
 sg13g2_o21ai_1 _25746_ (.B1(net671),
    .Y(_04192_),
    .A1(net730),
    .A2(_04189_));
 sg13g2_or2_1 _25747_ (.X(_04193_),
    .B(_04192_),
    .A(net398));
 sg13g2_a22oi_1 _25748_ (.Y(_04194_),
    .B1(_04191_),
    .B2(_04193_),
    .A2(_03184_),
    .A1(_05173_));
 sg13g2_nor2_1 _25749_ (.A(_03183_),
    .B(_04189_),
    .Y(_04196_));
 sg13g2_nand2_1 _25750_ (.Y(_04197_),
    .A(net650),
    .B(net389));
 sg13g2_nor2_1 _25751_ (.A(net672),
    .B(_04197_),
    .Y(_04198_));
 sg13g2_nor2_2 _25752_ (.A(_05625_),
    .B(_03453_),
    .Y(_04199_));
 sg13g2_xnor2_1 _25753_ (.Y(_04200_),
    .A(net1006),
    .B(net991));
 sg13g2_nand3_1 _25754_ (.B(net991),
    .C(_04197_),
    .A(net1006),
    .Y(_04201_));
 sg13g2_o21ai_1 _25755_ (.B1(_04201_),
    .Y(_04202_),
    .A1(_04199_),
    .A2(_04200_));
 sg13g2_o21ai_1 _25756_ (.B1(_06048_),
    .Y(_04203_),
    .A1(_04198_),
    .A2(_04202_));
 sg13g2_and3_1 _25757_ (.X(_04204_),
    .A(_05274_),
    .B(_05625_),
    .C(net389));
 sg13g2_a21oi_1 _25758_ (.A1(_05529_),
    .A2(_04197_),
    .Y(_04205_),
    .B1(_04199_));
 sg13g2_nand2_1 _25759_ (.Y(_04207_),
    .A(_05529_),
    .B(_04199_));
 sg13g2_o21ai_1 _25760_ (.B1(_04207_),
    .Y(_04208_),
    .A1(net672),
    .A2(_04205_));
 sg13g2_nand2b_1 _25761_ (.Y(_04209_),
    .B(_04199_),
    .A_N(net1006));
 sg13g2_nand2_1 _25762_ (.Y(_04210_),
    .A(_05197_),
    .B(_04204_));
 sg13g2_a21oi_1 _25763_ (.A1(_04209_),
    .A2(_04210_),
    .Y(_04211_),
    .B1(_05537_));
 sg13g2_a221oi_1 _25764_ (.B2(net678),
    .C1(_04211_),
    .B1(_04208_),
    .A1(net987),
    .Y(_04212_),
    .A2(_04204_));
 sg13g2_xnor2_1 _25765_ (.Y(_04213_),
    .A(net735),
    .B(_04189_));
 sg13g2_and2_1 _25766_ (.A(net1017),
    .B(_04213_),
    .X(_04214_));
 sg13g2_a221oi_1 _25767_ (.B2(_04212_),
    .C1(_04214_),
    .B1(_04203_),
    .A1(_03923_),
    .Y(_04215_),
    .A2(_04196_));
 sg13g2_o21ai_1 _25768_ (.B1(_04215_),
    .Y(_04216_),
    .A1(_03923_),
    .A2(_04194_));
 sg13g2_or2_1 _25769_ (.X(_04218_),
    .B(_04196_),
    .A(_03933_));
 sg13g2_a21oi_1 _25770_ (.A1(_03931_),
    .A2(_04213_),
    .Y(_04219_),
    .B1(_04218_));
 sg13g2_inv_1 _25771_ (.Y(_04220_),
    .A(_04197_));
 sg13g2_nor3_1 _25772_ (.A(_05200_),
    .B(net337),
    .C(net185),
    .Y(_04221_));
 sg13g2_nor3_1 _25773_ (.A(_06050_),
    .B(_04220_),
    .C(_04221_),
    .Y(_04222_));
 sg13g2_a22oi_1 _25774_ (.Y(_04223_),
    .B1(_04222_),
    .B2(_05530_),
    .A2(_04199_),
    .A1(_05989_));
 sg13g2_nor2_1 _25775_ (.A(_05275_),
    .B(_04223_),
    .Y(_04224_));
 sg13g2_a21oi_1 _25776_ (.A1(net672),
    .A2(net340),
    .Y(_04225_),
    .B1(_05200_));
 sg13g2_nor2_1 _25777_ (.A(_04207_),
    .B(_04225_),
    .Y(_04226_));
 sg13g2_or3_1 _25778_ (.A(_04219_),
    .B(_04224_),
    .C(_04226_),
    .X(_04227_));
 sg13g2_a21oi_1 _25779_ (.A1(_04216_),
    .A2(_04227_),
    .Y(_04229_),
    .B1(net79));
 sg13g2_xnor2_1 _25780_ (.Y(_04230_),
    .A(_03958_),
    .B(_04189_));
 sg13g2_a21oi_1 _25781_ (.A1(net112),
    .A2(_04230_),
    .Y(_04231_),
    .B1(_05205_));
 sg13g2_or2_1 _25782_ (.X(_04232_),
    .B(_04231_),
    .A(_04006_));
 sg13g2_nand3_1 _25783_ (.B(net80),
    .C(net51),
    .A(net637),
    .Y(_04233_));
 sg13g2_o21ai_1 _25784_ (.B1(_04233_),
    .Y(_00532_),
    .A1(_04229_),
    .A2(_04232_));
 sg13g2_xnor2_1 _25785_ (.Y(_04234_),
    .A(_13020_),
    .B(_00969_));
 sg13g2_nor2_1 _25786_ (.A(_00926_),
    .B(_04234_),
    .Y(_00559_));
 sg13g2_a21oi_1 _25787_ (.A1(_13020_),
    .A2(_00969_),
    .Y(_04235_),
    .B1(_00926_));
 sg13g2_and2_1 _25788_ (.A(_00904_),
    .B(_04235_),
    .X(_00560_));
 sg13g2_nor2_1 _25789_ (.A(_13031_),
    .B(_00926_),
    .Y(_00562_));
 sg13g2_inv_1 _25790_ (.Y(_04237_),
    .A(_00969_));
 sg13g2_buf_1 _25791_ (.A(_00022_),
    .X(_04238_));
 sg13g2_nor3_1 _25792_ (.A(_04237_),
    .B(_00904_),
    .C(_04238_),
    .Y(_04239_));
 sg13g2_mux2_1 _25793_ (.A0(\max7219.o_sck ),
    .A1(_00004_),
    .S(_04239_),
    .X(_04240_));
 sg13g2_nor2b_1 _25794_ (.A(_00926_),
    .B_N(_04240_),
    .Y(_00564_));
 sg13g2_inv_1 _25795_ (.Y(_04241_),
    .A(_01043_));
 sg13g2_nand2b_1 _25796_ (.Y(_04242_),
    .B(net7),
    .A_N(prev_rst_n));
 sg13g2_a21oi_1 _25797_ (.A1(_04241_),
    .A2(_04242_),
    .Y(_00276_),
    .B1(_06111_));
 sg13g2_buf_4 _25798_ (.X(_04243_),
    .A(\grid.row_select2[0] ));
 sg13g2_buf_2 _25799_ (.A(_04243_),
    .X(_04245_));
 sg13g2_buf_2 _25800_ (.A(_04245_),
    .X(_04246_));
 sg13g2_buf_2 _25801_ (.A(net388),
    .X(_04247_));
 sg13g2_buf_1 _25802_ (.A(\max7219.load_row ),
    .X(_04248_));
 sg13g2_xor2_1 _25803_ (.B(net1061),
    .A(net183),
    .X(_04249_));
 sg13g2_and3_1 _25804_ (.X(_00533_),
    .A(net317),
    .B(_00680_),
    .C(_04249_));
 sg13g2_nand2_1 _25805_ (.Y(_04250_),
    .A(_13063_),
    .B(net377));
 sg13g2_nand2_1 _25806_ (.Y(_04251_),
    .A(net668),
    .B(_04250_));
 sg13g2_buf_2 _25807_ (.A(\grid.row_select2[1] ),
    .X(_04252_));
 sg13g2_buf_2 _25808_ (.A(_04252_),
    .X(_04253_));
 sg13g2_inv_2 _25809_ (.Y(_04255_),
    .A(net724));
 sg13g2_nand2_1 _25810_ (.Y(_04256_),
    .A(net183),
    .B(net1061));
 sg13g2_xnor2_1 _25811_ (.Y(_04257_),
    .A(_04255_),
    .B(_04256_));
 sg13g2_nor2_1 _25812_ (.A(_04251_),
    .B(_04257_),
    .Y(_00534_));
 sg13g2_buf_2 _25813_ (.A(net724),
    .X(_04258_));
 sg13g2_buf_2 _25814_ (.A(net387),
    .X(_04259_));
 sg13g2_nand2_2 _25815_ (.Y(_04260_),
    .A(net182),
    .B(net183));
 sg13g2_xor2_1 _25816_ (.B(_04260_),
    .A(_00026_),
    .X(_04261_));
 sg13g2_buf_2 _25817_ (.A(\grid.row_select2[2] ),
    .X(_04262_));
 sg13g2_buf_2 _25818_ (.A(_04262_),
    .X(_04263_));
 sg13g2_buf_2 _25819_ (.A(net723),
    .X(_04265_));
 sg13g2_buf_1 _25820_ (.A(net386),
    .X(_04266_));
 sg13g2_nor2b_1 _25821_ (.A(net1061),
    .B_N(net181),
    .Y(_04267_));
 sg13g2_a21oi_1 _25822_ (.A1(_04248_),
    .A2(_04261_),
    .Y(_04268_),
    .B1(_04267_));
 sg13g2_nor2_1 _25823_ (.A(_04251_),
    .B(_04268_),
    .Y(_00535_));
 sg13g2_nor2b_1 _25824_ (.A(_00723_),
    .B_N(net1193),
    .Y(_04269_));
 sg13g2_nor2_1 _25825_ (.A(_00712_),
    .B(_13159_),
    .Y(_04270_));
 sg13g2_mux2_1 _25826_ (.A0(_13063_),
    .A1(_04270_),
    .S(net1193),
    .X(_04271_));
 sg13g2_nand2_1 _25827_ (.Y(_04272_),
    .A(net377),
    .B(_04271_));
 sg13g2_mux2_1 _25828_ (.A0(_04269_),
    .A1(_00723_),
    .S(_04272_),
    .X(_04273_));
 sg13g2_and2_1 _25829_ (.A(net378),
    .B(_04273_),
    .X(_00536_));
 sg13g2_nand2b_1 _25830_ (.Y(_04275_),
    .B(_00723_),
    .A_N(_00734_));
 sg13g2_nand2b_1 _25831_ (.Y(_04276_),
    .B(_00734_),
    .A_N(_00723_));
 sg13g2_o21ai_1 _25832_ (.B1(_04276_),
    .Y(_04277_),
    .A1(_04272_),
    .A2(_04275_));
 sg13g2_a22oi_1 _25833_ (.Y(_04278_),
    .B1(_04277_),
    .B2(net1193),
    .A2(_04272_),
    .A1(_00734_));
 sg13g2_nor2_1 _25834_ (.A(net214),
    .B(_04278_),
    .Y(_00537_));
 sg13g2_inv_1 _25835_ (.Y(_04279_),
    .A(_13289_));
 sg13g2_nor2_1 _25836_ (.A(net1193),
    .B(net1058),
    .Y(_04280_));
 sg13g2_nand2_1 _25837_ (.Y(_04281_),
    .A(_04279_),
    .B(_04280_));
 sg13g2_or3_1 _25838_ (.A(_04279_),
    .B(_00691_),
    .C(_13159_),
    .X(_04282_));
 sg13g2_o21ai_1 _25839_ (.B1(_04282_),
    .Y(_04284_),
    .A1(_13063_),
    .A2(_04281_));
 sg13g2_inv_2 _25840_ (.Y(_04285_),
    .A(net1196));
 sg13g2_inv_1 _25841_ (.Y(_04286_),
    .A(_13138_));
 sg13g2_nor2_2 _25842_ (.A(_04285_),
    .B(_04286_),
    .Y(_04287_));
 sg13g2_a21oi_1 _25843_ (.A1(_04287_),
    .A2(_00840_),
    .Y(_04288_),
    .B1(_13202_));
 sg13g2_nor2_1 _25844_ (.A(_13300_),
    .B(_04288_),
    .Y(_04289_));
 sg13g2_o21ai_1 _25845_ (.B1(net377),
    .Y(_04290_),
    .A1(_04284_),
    .A2(_04289_));
 sg13g2_nand2_2 _25846_ (.Y(_04291_),
    .A(_13010_),
    .B(_13031_));
 sg13g2_nor2_1 _25847_ (.A(net1193),
    .B(_04291_),
    .Y(_04292_));
 sg13g2_nand3_1 _25848_ (.B(net183),
    .C(_04266_),
    .A(net182),
    .Y(_04293_));
 sg13g2_nand2_1 _25849_ (.Y(_04295_),
    .A(_04248_),
    .B(_04293_));
 sg13g2_a21o_1 _25850_ (.A2(_04292_),
    .A1(_04279_),
    .B1(_04295_),
    .X(_04296_));
 sg13g2_a21oi_1 _25851_ (.A1(_04290_),
    .A2(_04296_),
    .Y(_00538_),
    .B1(net638));
 sg13g2_nand2_1 _25852_ (.Y(_04297_),
    .A(_00028_),
    .B(_04280_));
 sg13g2_nand3_1 _25853_ (.B(net377),
    .C(_04297_),
    .A(_04285_),
    .Y(_04298_));
 sg13g2_buf_1 _25854_ (.A(net1196),
    .X(_04299_));
 sg13g2_buf_1 _25855_ (.A(_04299_),
    .X(_04300_));
 sg13g2_a22oi_1 _25856_ (.Y(_04301_),
    .B1(_13300_),
    .B2(_04281_),
    .A2(_04291_),
    .A1(net385));
 sg13g2_a21oi_1 _25857_ (.A1(_04298_),
    .A2(_04301_),
    .Y(_00539_),
    .B1(net638));
 sg13g2_buf_2 _25858_ (.A(_04286_),
    .X(_04302_));
 sg13g2_nor3_1 _25859_ (.A(_04302_),
    .B(_04279_),
    .C(_13116_),
    .Y(_04304_));
 sg13g2_buf_1 _25860_ (.A(_13138_),
    .X(_04305_));
 sg13g2_nor3_1 _25861_ (.A(_04279_),
    .B(_00028_),
    .C(_04287_),
    .Y(_04306_));
 sg13g2_nor2b_1 _25862_ (.A(_04306_),
    .B_N(_04280_),
    .Y(_04307_));
 sg13g2_nor3_1 _25863_ (.A(net721),
    .B(_04291_),
    .C(_04307_),
    .Y(_04308_));
 sg13g2_o21ai_1 _25864_ (.B1(net385),
    .Y(_04309_),
    .A1(_04304_),
    .A2(_04308_));
 sg13g2_a21oi_1 _25865_ (.A1(net385),
    .A2(_13116_),
    .Y(_04310_),
    .B1(_04307_));
 sg13g2_o21ai_1 _25866_ (.B1(net721),
    .Y(_04311_),
    .A1(_04291_),
    .A2(_04310_));
 sg13g2_a21oi_1 _25867_ (.A1(_04309_),
    .A2(_04311_),
    .Y(_00540_),
    .B1(net638));
 sg13g2_buf_1 _25868_ (.A(net715),
    .X(_04312_));
 sg13g2_a21o_1 _25869_ (.A2(_13300_),
    .A1(net377),
    .B1(\max7219.max7219_enabled ),
    .X(_04314_));
 sg13g2_a22oi_1 _25870_ (.Y(_04315_),
    .B1(_04314_),
    .B2(_13289_),
    .A2(_04250_),
    .A1(\max7219.max7219_enabled ));
 sg13g2_nor2_1 _25871_ (.A(net180),
    .B(_04315_),
    .Y(_00541_));
 sg13g2_nor2b_1 _25872_ (.A(net1195),
    .B_N(_13191_),
    .Y(_04316_));
 sg13g2_nor2_1 _25873_ (.A(net1058),
    .B(_13289_),
    .Y(_04317_));
 sg13g2_o21ai_1 _25874_ (.B1(_04292_),
    .Y(_04318_),
    .A1(_04270_),
    .A2(_04317_));
 sg13g2_buf_1 _25875_ (.A(_04318_),
    .X(_04319_));
 sg13g2_mux2_1 _25876_ (.A0(_04316_),
    .A1(net1195),
    .S(_04319_),
    .X(_04320_));
 sg13g2_and2_1 _25877_ (.A(net378),
    .B(_04320_),
    .X(_00542_));
 sg13g2_inv_1 _25878_ (.Y(_04321_),
    .A(_13235_));
 sg13g2_nand2_1 _25879_ (.Y(_04323_),
    .A(_04321_),
    .B(net1195));
 sg13g2_nand2b_1 _25880_ (.Y(_04324_),
    .B(_13235_),
    .A_N(net1195));
 sg13g2_o21ai_1 _25881_ (.B1(_04324_),
    .Y(_04325_),
    .A1(_04319_),
    .A2(_04323_));
 sg13g2_a22oi_1 _25882_ (.Y(_04326_),
    .B1(_04325_),
    .B2(net1058),
    .A2(_04319_),
    .A1(_13235_));
 sg13g2_nor2_1 _25883_ (.A(net180),
    .B(_04326_),
    .Y(_00543_));
 sg13g2_and2_1 _25884_ (.A(_13235_),
    .B(net1195),
    .X(_04327_));
 sg13g2_xnor2_1 _25885_ (.Y(_04328_),
    .A(_00027_),
    .B(_04327_));
 sg13g2_nand2_1 _25886_ (.Y(_04329_),
    .A(_13202_),
    .B(_04328_));
 sg13g2_nor2_1 _25887_ (.A(_04319_),
    .B(_04329_),
    .Y(_04330_));
 sg13g2_a21oi_1 _25888_ (.A1(_13213_),
    .A2(_04319_),
    .Y(_04331_),
    .B1(_04330_));
 sg13g2_nor2_1 _25889_ (.A(net180),
    .B(_04331_),
    .Y(_00544_));
 sg13g2_a21oi_1 _25890_ (.A1(_13159_),
    .A2(_04281_),
    .Y(_04333_),
    .B1(_04291_));
 sg13g2_nor2_1 _25891_ (.A(_00712_),
    .B(_04333_),
    .Y(_04334_));
 sg13g2_nand3_1 _25892_ (.B(_04297_),
    .C(_04333_),
    .A(_00691_),
    .Y(_04335_));
 sg13g2_nand3b_1 _25893_ (.B(_04335_),
    .C(net378),
    .Y(_00545_),
    .A_N(_04334_));
 sg13g2_nor2b_1 _25894_ (.A(net181),
    .B_N(\max7219.load_row ),
    .Y(_04336_));
 sg13g2_nor2_1 _25895_ (.A(net182),
    .B(net183),
    .Y(_04337_));
 sg13g2_nand2_1 _25896_ (.Y(_04338_),
    .A(_04336_),
    .B(_04337_));
 sg13g2_mux4_1 _25897_ (.S0(net725),
    .A0(_10820_),
    .A1(_11195_),
    .A2(_11574_),
    .A3(net1096),
    .S1(net724),
    .X(_04339_));
 sg13g2_mux4_1 _25898_ (.S0(_04243_),
    .A0(_12300_),
    .A1(_12652_),
    .A2(_13014_),
    .A3(_04947_),
    .S1(net724),
    .X(_04340_));
 sg13g2_mux2_1 _25899_ (.A0(_04339_),
    .A1(_04340_),
    .S(_04262_),
    .X(_04342_));
 sg13g2_nor2_2 _25900_ (.A(net1196),
    .B(net384),
    .Y(_04343_));
 sg13g2_mux4_1 _25901_ (.S0(net725),
    .A0(net936),
    .A1(net1147),
    .A2(_08193_),
    .A3(net1136),
    .S1(net724),
    .X(_04344_));
 sg13g2_mux4_1 _25902_ (.S0(_04245_),
    .A0(net1129),
    .A1(_09696_),
    .A2(net871),
    .A3(_10431_),
    .S1(net724),
    .X(_04345_));
 sg13g2_mux2_1 _25903_ (.A0(_04344_),
    .A1(_04345_),
    .S(net723),
    .X(_04346_));
 sg13g2_a22oi_1 _25904_ (.Y(_04347_),
    .B1(_04343_),
    .B2(_04346_),
    .A2(_04342_),
    .A1(_04287_));
 sg13g2_nand2_1 _25905_ (.Y(_04348_),
    .A(net1195),
    .B(_04347_));
 sg13g2_buf_2 _25906_ (.A(_04243_),
    .X(_04349_));
 sg13g2_mux4_1 _25907_ (.S0(net720),
    .A0(_10784_),
    .A1(_11154_),
    .A2(_12266_),
    .A3(net1088),
    .S1(_04262_),
    .X(_04350_));
 sg13g2_buf_2 _25908_ (.A(_04252_),
    .X(_04351_));
 sg13g2_mux4_1 _25909_ (.S0(_04243_),
    .A0(_11521_),
    .A1(_11878_),
    .A2(net1084),
    .A3(net1027),
    .S1(_04262_),
    .X(_04353_));
 sg13g2_and2_1 _25910_ (.A(net719),
    .B(_04353_),
    .X(_04354_));
 sg13g2_a21oi_1 _25911_ (.A1(_04255_),
    .A2(_04350_),
    .Y(_04355_),
    .B1(_04354_));
 sg13g2_mux4_1 _25912_ (.S0(_04243_),
    .A0(_07389_),
    .A1(net1148),
    .A2(net1141),
    .A3(_08505_),
    .S1(_04252_),
    .X(_04356_));
 sg13g2_mux4_1 _25913_ (.S0(_04243_),
    .A0(_08924_),
    .A1(_09659_),
    .A2(_10021_),
    .A3(_10398_),
    .S1(_04252_),
    .X(_04357_));
 sg13g2_mux2_1 _25914_ (.A0(_04356_),
    .A1(_04357_),
    .S(_04262_),
    .X(_04358_));
 sg13g2_a21oi_1 _25915_ (.A1(_04343_),
    .A2(_04358_),
    .Y(_04359_),
    .B1(\max7219.max7219_row[0] ));
 sg13g2_o21ai_1 _25916_ (.B1(_04359_),
    .Y(_04360_),
    .A1(_13159_),
    .A2(_04355_));
 sg13g2_a21o_1 _25917_ (.A2(_04360_),
    .A1(_04348_),
    .B1(net384),
    .X(_04361_));
 sg13g2_buf_2 _25918_ (.A(_04243_),
    .X(_04362_));
 sg13g2_buf_2 _25919_ (.A(net718),
    .X(_04364_));
 sg13g2_mux4_1 _25920_ (.S0(net719),
    .A0(net1179),
    .A1(net887),
    .A2(_04943_),
    .A3(_00709_),
    .S1(net383),
    .X(_04365_));
 sg13g2_buf_2 _25921_ (.A(net725),
    .X(_04366_));
 sg13g2_buf_2 _25922_ (.A(net724),
    .X(_04367_));
 sg13g2_mux4_1 _25923_ (.S0(net382),
    .A0(net1064),
    .A1(net993),
    .A2(_05491_),
    .A3(_05475_),
    .S1(net381),
    .X(_04368_));
 sg13g2_mux4_1 _25924_ (.S0(net382),
    .A0(net1079),
    .A1(net758),
    .A2(_02596_),
    .A3(net1067),
    .S1(net381),
    .X(_04369_));
 sg13g2_mux4_1 _25925_ (.S0(net382),
    .A0(_05901_),
    .A1(net965),
    .A2(net957),
    .A3(net1161),
    .S1(net381),
    .X(_04370_));
 sg13g2_mux4_1 _25926_ (.S0(net722),
    .A0(_04365_),
    .A1(_04368_),
    .A2(_04369_),
    .A3(_04370_),
    .S1(_04265_),
    .X(_04371_));
 sg13g2_or2_1 _25927_ (.X(_04372_),
    .B(_04371_),
    .A(_04348_));
 sg13g2_mux4_1 _25928_ (.S0(net719),
    .A0(net1180),
    .A1(_09334_),
    .A2(_04705_),
    .A3(net780),
    .S1(net383),
    .X(_04373_));
 sg13g2_mux4_1 _25929_ (.S0(_04366_),
    .A0(_03348_),
    .A1(_05418_),
    .A2(net997),
    .A3(net1175),
    .S1(net381),
    .X(_04375_));
 sg13g2_mux4_1 _25930_ (.S0(net388),
    .A0(_01743_),
    .A1(_02142_),
    .A2(_02554_),
    .A3(net1068),
    .S1(net387),
    .X(_04376_));
 sg13g2_mux4_1 _25931_ (.S0(_04246_),
    .A0(net1172),
    .A1(net1169),
    .A2(net1166),
    .A3(net1163),
    .S1(_04258_),
    .X(_04377_));
 sg13g2_mux4_1 _25932_ (.S0(net722),
    .A0(_04373_),
    .A1(_04375_),
    .A2(_04376_),
    .A3(_04377_),
    .S1(net386),
    .X(_04378_));
 sg13g2_or2_1 _25933_ (.X(_04379_),
    .B(_04378_),
    .A(_04360_));
 sg13g2_nand4_1 _25934_ (.B(_04361_),
    .C(_04372_),
    .A(_04321_),
    .Y(_04380_),
    .D(_04379_));
 sg13g2_mux4_1 _25935_ (.S0(net388),
    .A0(_07207_),
    .A1(_07608_),
    .A2(net923),
    .A3(net915),
    .S1(net387),
    .X(_04381_));
 sg13g2_buf_2 _25936_ (.A(_04252_),
    .X(_04382_));
 sg13g2_buf_2 _25937_ (.A(net720),
    .X(_04383_));
 sg13g2_mux4_1 _25938_ (.S0(net717),
    .A0(_10609_),
    .A1(net1102),
    .A2(_11002_),
    .A3(net825),
    .S1(net380),
    .X(_04384_));
 sg13g2_mux4_1 _25939_ (.S0(net718),
    .A0(net907),
    .A1(_09525_),
    .A2(_09857_),
    .A3(_10572_),
    .S1(net719),
    .X(_04386_));
 sg13g2_mux4_1 _25940_ (.S0(net718),
    .A0(_12100_),
    .A1(net1090),
    .A2(net794),
    .A3(net1039),
    .S1(net719),
    .X(_04387_));
 sg13g2_mux4_1 _25941_ (.S0(net722),
    .A0(_04381_),
    .A1(_04384_),
    .A2(_04386_),
    .A3(_04387_),
    .S1(net386),
    .X(_04388_));
 sg13g2_mux4_1 _25942_ (.S0(net718),
    .A0(net1018),
    .A1(_02421_),
    .A2(net896),
    .A3(_13192_),
    .S1(net719),
    .X(_04389_));
 sg13g2_mux4_1 _25943_ (.S0(_04246_),
    .A0(net733),
    .A1(net1013),
    .A2(_05195_),
    .A3(_05192_),
    .S1(_04258_),
    .X(_04390_));
 sg13g2_mux4_1 _25944_ (.S0(_04362_),
    .A0(_01555_),
    .A1(net766),
    .A2(net754),
    .A3(net745),
    .S1(_04351_),
    .X(_04391_));
 sg13g2_mux4_1 _25945_ (.S0(net718),
    .A0(net984),
    .A1(net972),
    .A2(net962),
    .A3(net955),
    .S1(_04351_),
    .X(_04392_));
 sg13g2_mux4_1 _25946_ (.S0(net722),
    .A0(_04389_),
    .A1(_04390_),
    .A2(_04391_),
    .A3(_04392_),
    .S1(_04263_),
    .X(_04393_));
 sg13g2_mux2_1 _25947_ (.A0(_04388_),
    .A1(_04393_),
    .S(net384),
    .X(_04394_));
 sg13g2_buf_2 _25948_ (.A(net719),
    .X(_04395_));
 sg13g2_mux4_1 _25949_ (.S0(net383),
    .A0(_12341_),
    .A1(net454),
    .A2(net787),
    .A3(net688),
    .S1(net379),
    .X(_04397_));
 sg13g2_nand2_1 _25950_ (.Y(_04398_),
    .A(_04287_),
    .B(_04397_));
 sg13g2_mux4_1 _25951_ (.S0(_04247_),
    .A0(net975),
    .A1(net964),
    .A2(net956),
    .A3(_07076_),
    .S1(_04259_),
    .X(_04399_));
 sg13g2_nor2_1 _25952_ (.A(_04285_),
    .B(net721),
    .Y(_04400_));
 sg13g2_nand2_1 _25953_ (.Y(_04401_),
    .A(_04399_),
    .B(_04400_));
 sg13g2_mux4_1 _25954_ (.S0(net380),
    .A0(net897),
    .A1(_09732_),
    .A2(net870),
    .A3(_10469_),
    .S1(net379),
    .X(_04402_));
 sg13g2_mux4_1 _25955_ (.S0(net383),
    .A0(net768),
    .A1(net757),
    .A2(net746),
    .A3(net736),
    .S1(_04395_),
    .X(_04403_));
 sg13g2_nor2_1 _25956_ (.A(net722),
    .B(net721),
    .Y(_04404_));
 sg13g2_a22oi_1 _25957_ (.Y(_04405_),
    .B1(_04403_),
    .B2(_04404_),
    .A2(_04402_),
    .A1(_04343_));
 sg13g2_nand4_1 _25958_ (.B(_04398_),
    .C(_04401_),
    .A(net386),
    .Y(_04406_),
    .D(_04405_));
 sg13g2_mux4_1 _25959_ (.S0(net380),
    .A0(net935),
    .A1(_07856_),
    .A2(_08230_),
    .A3(net908),
    .S1(net379),
    .X(_04408_));
 sg13g2_mux4_1 _25960_ (.S0(net380),
    .A0(_05016_),
    .A1(net1022),
    .A2(net1123),
    .A3(net778),
    .S1(net379),
    .X(_04409_));
 sg13g2_a221oi_1 _25961_ (.B2(_04404_),
    .C1(net386),
    .B1(_04409_),
    .A1(_04343_),
    .Y(_04410_),
    .A2(_04408_));
 sg13g2_mux4_1 _25962_ (.S0(net381),
    .A0(net849),
    .A1(net828),
    .A2(_11235_),
    .A3(_11973_),
    .S1(net183),
    .X(_04411_));
 sg13g2_mux4_1 _25963_ (.S0(net383),
    .A0(net390),
    .A1(net650),
    .A2(_05535_),
    .A3(_05524_),
    .S1(_04395_),
    .X(_04412_));
 sg13g2_a22oi_1 _25964_ (.Y(_04413_),
    .B1(_04412_),
    .B2(_04400_),
    .A2(_04411_),
    .A1(_04287_));
 sg13g2_a21oi_1 _25965_ (.A1(_04410_),
    .A2(_04413_),
    .Y(_04414_),
    .B1(_04324_));
 sg13g2_a221oi_1 _25966_ (.B2(_04414_),
    .C1(_13224_),
    .B1(_04406_),
    .A1(_04327_),
    .Y(_04415_),
    .A2(_04394_));
 sg13g2_mux2_1 _25967_ (.A0(_03300_),
    .A1(_05365_),
    .S(_04383_),
    .X(_04416_));
 sg13g2_nor2_1 _25968_ (.A(_04366_),
    .B(_05361_),
    .Y(_04417_));
 sg13g2_a21oi_1 _25969_ (.A1(net383),
    .A2(_05375_),
    .Y(_04419_),
    .B1(_04417_));
 sg13g2_nor2_1 _25970_ (.A(net382),
    .B(_10737_),
    .Y(_04420_));
 sg13g2_a21oi_1 _25971_ (.A1(net383),
    .A2(_11162_),
    .Y(_04421_),
    .B1(_04420_));
 sg13g2_mux2_1 _25972_ (.A0(_11481_),
    .A1(_11843_),
    .S(net382),
    .X(_04422_));
 sg13g2_mux4_1 _25973_ (.S0(net379),
    .A0(_04416_),
    .A1(_04419_),
    .A2(_04421_),
    .A3(_04422_),
    .S1(net721),
    .X(_04423_));
 sg13g2_nand2_1 _25974_ (.Y(_04424_),
    .A(net385),
    .B(_04423_));
 sg13g2_mux4_1 _25975_ (.S0(net388),
    .A0(net1156),
    .A1(net1150),
    .A2(net920),
    .A3(_08469_),
    .S1(net387),
    .X(_04425_));
 sg13g2_mux4_1 _25976_ (.S0(net717),
    .A0(_04131_),
    .A1(net889),
    .A2(net1029),
    .A3(net782),
    .S1(_04383_),
    .X(_04426_));
 sg13g2_mux2_1 _25977_ (.A0(_04425_),
    .A1(_04426_),
    .S(net384),
    .X(_04427_));
 sg13g2_a21oi_1 _25978_ (.A1(_04285_),
    .A2(_04427_),
    .Y(_04428_),
    .B1(net386));
 sg13g2_a21oi_1 _25979_ (.A1(_04424_),
    .A2(_04428_),
    .Y(_04430_),
    .B1(_13256_));
 sg13g2_mux4_1 _25980_ (.S0(net383),
    .A0(_12229_),
    .A1(net1089),
    .A2(_12938_),
    .A3(net1030),
    .S1(net379),
    .X(_04431_));
 sg13g2_mux4_1 _25981_ (.S0(_04364_),
    .A0(net979),
    .A1(net968),
    .A2(net959),
    .A3(net950),
    .S1(net379),
    .X(_04432_));
 sg13g2_mux2_1 _25982_ (.A0(_04431_),
    .A1(_04432_),
    .S(net384),
    .X(_04433_));
 sg13g2_mux4_1 _25983_ (.S0(net382),
    .A0(net902),
    .A1(net881),
    .A2(_09980_),
    .A3(_10353_),
    .S1(net381),
    .X(_04434_));
 sg13g2_mux4_1 _25984_ (.S0(net720),
    .A0(_01677_),
    .A1(net761),
    .A2(_02491_),
    .A3(_02888_),
    .S1(_04253_),
    .X(_04435_));
 sg13g2_and2_1 _25985_ (.A(net384),
    .B(_04435_),
    .X(_04436_));
 sg13g2_a21oi_1 _25986_ (.A1(net721),
    .A2(_04434_),
    .Y(_04437_),
    .B1(_04436_));
 sg13g2_o21ai_1 _25987_ (.B1(net386),
    .Y(_04438_),
    .A1(net385),
    .A2(_04437_));
 sg13g2_a21o_1 _25988_ (.A2(_04433_),
    .A1(net385),
    .B1(_04438_),
    .X(_04439_));
 sg13g2_a21oi_1 _25989_ (.A1(_04430_),
    .A2(_04439_),
    .Y(_04441_),
    .B1(_13213_));
 sg13g2_nor2_1 _25990_ (.A(_04321_),
    .B(net1195),
    .Y(_04442_));
 sg13g2_mux4_1 _25991_ (.S0(net380),
    .A0(_07302_),
    .A1(_07749_),
    .A2(_08051_),
    .A3(_08422_),
    .S1(net379),
    .X(_04443_));
 sg13g2_mux4_1 _25992_ (.S0(net388),
    .A0(_10685_),
    .A1(net844),
    .A2(net834),
    .A3(net1098),
    .S1(net387),
    .X(_04444_));
 sg13g2_nand2_1 _25993_ (.Y(_04445_),
    .A(net722),
    .B(_04444_));
 sg13g2_o21ai_1 _25994_ (.B1(_04445_),
    .Y(_04446_),
    .A1(net385),
    .A2(_04443_));
 sg13g2_mux4_1 _25995_ (.S0(net380),
    .A0(_08844_),
    .A1(_09587_),
    .A2(_12176_),
    .A3(_12533_),
    .S1(net722),
    .X(_04447_));
 sg13g2_mux4_1 _25996_ (.S0(net388),
    .A0(_09936_),
    .A1(net865),
    .A2(_12891_),
    .A3(net1036),
    .S1(net1196),
    .X(_04448_));
 sg13g2_nand2_1 _25997_ (.Y(_04449_),
    .A(net182),
    .B(_04448_));
 sg13g2_o21ai_1 _25998_ (.B1(_04449_),
    .Y(_04450_),
    .A1(net182),
    .A2(_04447_));
 sg13g2_mux4_1 _25999_ (.S0(net382),
    .A0(_03326_),
    .A1(_03185_),
    .A2(net1126),
    .A3(net783),
    .S1(net381),
    .X(_04452_));
 sg13g2_mux4_1 _26000_ (.S0(net382),
    .A0(_03246_),
    .A1(net669),
    .A2(net1004),
    .A3(_05311_),
    .S1(_04367_),
    .X(_04453_));
 sg13g2_mux2_1 _26001_ (.A0(_04452_),
    .A1(_04453_),
    .S(net722),
    .X(_04454_));
 sg13g2_mux4_1 _26002_ (.S0(net380),
    .A0(_01627_),
    .A1(net763),
    .A2(_02457_),
    .A3(_02844_),
    .S1(_04367_),
    .X(_04455_));
 sg13g2_mux4_1 _26003_ (.S0(net718),
    .A0(net981),
    .A1(net969),
    .A2(_06539_),
    .A3(net1164),
    .S1(net719),
    .X(_04456_));
 sg13g2_nand2_1 _26004_ (.Y(_04457_),
    .A(_04299_),
    .B(_04456_));
 sg13g2_o21ai_1 _26005_ (.B1(_04457_),
    .Y(_04458_),
    .A1(_04300_),
    .A2(_04455_));
 sg13g2_mux4_1 _26006_ (.S0(_04265_),
    .A0(_04446_),
    .A1(_04450_),
    .A2(_04454_),
    .A3(_04458_),
    .S1(_04302_),
    .X(_04459_));
 sg13g2_mux4_1 _26007_ (.S0(_04349_),
    .A0(_07268_),
    .A1(_07614_),
    .A2(_08034_),
    .A3(_08413_),
    .S1(net717),
    .X(_04460_));
 sg13g2_mux4_1 _26008_ (.S0(net720),
    .A0(_08811_),
    .A1(_09579_),
    .A2(_09865_),
    .A3(_10252_),
    .S1(net717),
    .X(_04461_));
 sg13g2_mux2_1 _26009_ (.A0(_04460_),
    .A1(_04461_),
    .S(net723),
    .X(_04463_));
 sg13g2_mux4_1 _26010_ (.S0(net720),
    .A0(net1107),
    .A1(_11056_),
    .A2(_11399_),
    .A3(_11754_),
    .S1(net717),
    .X(_04464_));
 sg13g2_mux4_1 _26011_ (.S0(net720),
    .A0(_12163_),
    .A1(_12491_),
    .A2(net1085),
    .A3(net1184),
    .S1(net717),
    .X(_04465_));
 sg13g2_mux2_1 _26012_ (.A0(_04464_),
    .A1(_04465_),
    .S(net723),
    .X(_04466_));
 sg13g2_mux2_1 _26013_ (.A0(_04463_),
    .A1(_04466_),
    .S(net385),
    .X(_04467_));
 sg13g2_nand2_1 _26014_ (.Y(_04468_),
    .A(net721),
    .B(_04467_));
 sg13g2_nor2b_1 _26015_ (.A(net380),
    .B_N(\grid.cell_13_0.s ),
    .Y(_04469_));
 sg13g2_a21oi_1 _26016_ (.A1(_04364_),
    .A2(_06856_),
    .Y(_04470_),
    .B1(_04469_));
 sg13g2_nand3_1 _26017_ (.B(_04259_),
    .C(_04470_),
    .A(_04300_),
    .Y(_04471_));
 sg13g2_mux2_1 _26018_ (.A0(net1174),
    .A1(_06095_),
    .S(net725),
    .X(_04472_));
 sg13g2_nor3_1 _26019_ (.A(_04285_),
    .B(net387),
    .C(_04472_),
    .Y(_04474_));
 sg13g2_mux2_1 _26020_ (.A0(_02426_),
    .A1(net1071),
    .S(net720),
    .X(_04475_));
 sg13g2_nor3_1 _26021_ (.A(net1196),
    .B(_04255_),
    .C(_04475_),
    .Y(_04476_));
 sg13g2_nand2_1 _26022_ (.Y(_04477_),
    .A(net384),
    .B(net723));
 sg13g2_mux2_1 _26023_ (.A0(_01595_),
    .A1(_01995_),
    .S(net718),
    .X(_04478_));
 sg13g2_nor3_1 _26024_ (.A(_13127_),
    .B(net381),
    .C(_04478_),
    .Y(_04479_));
 sg13g2_nor4_1 _26025_ (.A(_04474_),
    .B(_04476_),
    .C(_04477_),
    .D(_04479_),
    .Y(_04480_));
 sg13g2_mux4_1 _26026_ (.S0(net388),
    .A0(_03173_),
    .A1(_05273_),
    .A2(_05172_),
    .A3(_05214_),
    .S1(net387),
    .X(_04481_));
 sg13g2_mux4_1 _26027_ (.S0(net388),
    .A0(_02863_),
    .A1(_02173_),
    .A2(_09216_),
    .A3(_13229_),
    .S1(net387),
    .X(_04482_));
 sg13g2_mux2_1 _26028_ (.A0(_04481_),
    .A1(_04482_),
    .S(_04285_),
    .X(_04483_));
 sg13g2_nor2_1 _26029_ (.A(net721),
    .B(net723),
    .Y(_04485_));
 sg13g2_a221oi_1 _26030_ (.B2(_04485_),
    .C1(_13246_),
    .B1(_04483_),
    .A1(_04471_),
    .Y(_04486_),
    .A2(_04480_));
 sg13g2_mux4_1 _26031_ (.S0(net725),
    .A0(_09860_),
    .A1(_10248_),
    .A2(net795),
    .A3(_02658_),
    .S1(net1196),
    .X(_04487_));
 sg13g2_mux4_1 _26032_ (.S0(net725),
    .A0(_08739_),
    .A1(_09539_),
    .A2(_12098_),
    .A3(_12452_),
    .S1(net1196),
    .X(_04488_));
 sg13g2_mux2_1 _26033_ (.A0(_04487_),
    .A1(_04488_),
    .S(_04255_),
    .X(_04489_));
 sg13g2_nand3_1 _26034_ (.B(net386),
    .C(_04489_),
    .A(_04305_),
    .Y(_04490_));
 sg13g2_mux4_1 _26035_ (.S0(net725),
    .A0(_10607_),
    .A1(_10998_),
    .A2(_11352_),
    .A3(_11716_),
    .S1(net724),
    .X(_04491_));
 sg13g2_mux4_1 _26036_ (.S0(net725),
    .A0(_07203_),
    .A1(net1152),
    .A2(net1143),
    .A3(net914),
    .S1(_04253_),
    .X(_04492_));
 sg13g2_mux2_1 _26037_ (.A0(_04491_),
    .A1(_04492_),
    .S(_04285_),
    .X(_04493_));
 sg13g2_nand3b_1 _26038_ (.B(_04493_),
    .C(_04305_),
    .Y(_04494_),
    .A_N(net723));
 sg13g2_and3_1 _26039_ (.X(_04496_),
    .A(_13246_),
    .B(_04490_),
    .C(_04494_));
 sg13g2_mux4_1 _26040_ (.S0(_04362_),
    .A0(_03168_),
    .A1(net1016),
    .A2(_05226_),
    .A3(_05228_),
    .S1(net717),
    .X(_04497_));
 sg13g2_mux4_1 _26041_ (.S0(net718),
    .A0(net986),
    .A1(net973),
    .A2(_06478_),
    .A3(_06837_),
    .S1(_04382_),
    .X(_04498_));
 sg13g2_mux2_1 _26042_ (.A0(_04497_),
    .A1(_04498_),
    .S(_04263_),
    .X(_04499_));
 sg13g2_mux4_1 _26043_ (.S0(net720),
    .A0(net1186),
    .A1(_02076_),
    .A2(net895),
    .A3(net1083),
    .S1(_04382_),
    .X(_04500_));
 sg13g2_mux4_1 _26044_ (.S0(_04349_),
    .A0(_01552_),
    .A1(_01952_),
    .A2(net1073),
    .A3(net744),
    .S1(net717),
    .X(_04501_));
 sg13g2_mux2_1 _26045_ (.A0(_04500_),
    .A1(_04501_),
    .S(net723),
    .X(_04502_));
 sg13g2_mux2_1 _26046_ (.A0(_04499_),
    .A1(_04502_),
    .S(_04285_),
    .X(_04503_));
 sg13g2_nand2_1 _26047_ (.Y(_04504_),
    .A(net384),
    .B(_04503_));
 sg13g2_a22oi_1 _26048_ (.Y(_04505_),
    .B1(_04496_),
    .B2(_04504_),
    .A2(_04486_),
    .A1(_04468_));
 sg13g2_a22oi_1 _26049_ (.Y(_04507_),
    .B1(_04505_),
    .B2(_04321_),
    .A2(_04459_),
    .A1(_04442_));
 sg13g2_a22oi_1 _26050_ (.Y(_04508_),
    .B1(_04441_),
    .B2(_04507_),
    .A2(_04415_),
    .A1(_04380_));
 sg13g2_buf_1 _26051_ (.A(_04508_),
    .X(_04509_));
 sg13g2_inv_1 _26052_ (.Y(_04510_),
    .A(_00253_));
 sg13g2_nor3_1 _26053_ (.A(net181),
    .B(_04510_),
    .C(_04338_),
    .Y(_04511_));
 sg13g2_a22oi_1 _26054_ (.Y(_04512_),
    .B1(net28),
    .B2(_04511_),
    .A2(_04338_),
    .A1(\max7219.row_data[0] ));
 sg13g2_nor2_1 _26055_ (.A(net180),
    .B(_04512_),
    .Y(_00546_));
 sg13g2_or2_1 _26056_ (.X(_04513_),
    .B(net183),
    .A(net182));
 sg13g2_buf_1 _26057_ (.A(_04513_),
    .X(_04514_));
 sg13g2_nor2b_1 _26058_ (.A(net182),
    .B_N(net183),
    .Y(_04515_));
 sg13g2_nand3_1 _26059_ (.B(_04336_),
    .C(_04515_),
    .A(_00253_),
    .Y(_04517_));
 sg13g2_o21ai_1 _26060_ (.B1(_04517_),
    .Y(_04518_),
    .A1(\max7219.row_data[1] ),
    .A2(_04514_));
 sg13g2_nand2_1 _26061_ (.Y(_04519_),
    .A(_04336_),
    .B(_04515_));
 sg13g2_nor2_1 _26062_ (.A(_04509_),
    .B(_04519_),
    .Y(_04520_));
 sg13g2_nand2b_1 _26063_ (.Y(_04521_),
    .B(net1061),
    .A_N(net181));
 sg13g2_buf_1 _26064_ (.A(_04521_),
    .X(_04522_));
 sg13g2_nand3_1 _26065_ (.B(_04510_),
    .C(_04260_),
    .A(net1194),
    .Y(_04523_));
 sg13g2_nor2_1 _26066_ (.A(_04522_),
    .B(_04523_),
    .Y(_04524_));
 sg13g2_a22oi_1 _26067_ (.Y(_04525_),
    .B1(net28),
    .B2(_04524_),
    .A2(\max7219.row_data[1] ),
    .A1(net668));
 sg13g2_nor3_1 _26068_ (.A(_04518_),
    .B(_04520_),
    .C(_04525_),
    .Y(_00547_));
 sg13g2_nand2b_1 _26069_ (.Y(_04527_),
    .B(net182),
    .A_N(_04247_));
 sg13g2_buf_1 _26070_ (.A(_04527_),
    .X(_04528_));
 sg13g2_nor2_1 _26071_ (.A(_04522_),
    .B(_04528_),
    .Y(_04529_));
 sg13g2_nand2_1 _26072_ (.Y(_04530_),
    .A(net28),
    .B(_04529_));
 sg13g2_o21ai_1 _26073_ (.B1(\max7219.row_data[2] ),
    .Y(_04531_),
    .A1(_04522_),
    .A2(_04528_));
 sg13g2_a21oi_1 _26074_ (.A1(_04530_),
    .A2(_04531_),
    .Y(_00548_),
    .B1(net638));
 sg13g2_o21ai_1 _26075_ (.B1(\max7219.row_data[3] ),
    .Y(_04532_),
    .A1(_04260_),
    .A2(_04522_));
 sg13g2_nand2_1 _26076_ (.Y(_04533_),
    .A(net181),
    .B(_04337_));
 sg13g2_o21ai_1 _26077_ (.B1(_04533_),
    .Y(_04534_),
    .A1(net181),
    .A2(_04260_));
 sg13g2_and2_1 _26078_ (.A(net1061),
    .B(_04534_),
    .X(_04535_));
 sg13g2_nand3_1 _26079_ (.B(net28),
    .C(_04535_),
    .A(_04510_),
    .Y(_04537_));
 sg13g2_a21oi_1 _26080_ (.A1(_04532_),
    .A2(_04537_),
    .Y(_00549_),
    .B1(net638));
 sg13g2_nand2_1 _26081_ (.Y(_04538_),
    .A(_00253_),
    .B(_04535_));
 sg13g2_nand2_2 _26082_ (.Y(_04539_),
    .A(net181),
    .B(net1061));
 sg13g2_nor2_1 _26083_ (.A(_04514_),
    .B(_04539_),
    .Y(_04540_));
 sg13g2_a22oi_1 _26084_ (.Y(_04541_),
    .B1(_04540_),
    .B2(_04509_),
    .A2(_04538_),
    .A1(\max7219.row_data[4] ));
 sg13g2_nor2_1 _26085_ (.A(net180),
    .B(_04541_),
    .Y(_00550_));
 sg13g2_nand3_1 _26086_ (.B(net1061),
    .C(_04515_),
    .A(_04266_),
    .Y(_04542_));
 sg13g2_nand2b_1 _26087_ (.Y(_04543_),
    .B(_04337_),
    .A_N(\max7219.row_data[5] ));
 sg13g2_o21ai_1 _26088_ (.B1(_04543_),
    .Y(_04544_),
    .A1(_04510_),
    .A2(_04542_));
 sg13g2_nor2_1 _26089_ (.A(net28),
    .B(_04542_),
    .Y(_04546_));
 sg13g2_nor2_1 _26090_ (.A(_04523_),
    .B(_04539_),
    .Y(_04547_));
 sg13g2_a22oi_1 _26091_ (.Y(_04548_),
    .B1(net28),
    .B2(_04547_),
    .A2(\max7219.row_data[5] ),
    .A1(net668));
 sg13g2_nor3_1 _26092_ (.A(_04544_),
    .B(_04546_),
    .C(_04548_),
    .Y(_00551_));
 sg13g2_nor2_1 _26093_ (.A(_04528_),
    .B(_04539_),
    .Y(_04549_));
 sg13g2_nand2_1 _26094_ (.Y(_04550_),
    .A(net28),
    .B(_04549_));
 sg13g2_o21ai_1 _26095_ (.B1(\max7219.row_data[6] ),
    .Y(_04551_),
    .A1(_04528_),
    .A2(_04539_));
 sg13g2_a21oi_1 _26096_ (.A1(_04550_),
    .A2(_04551_),
    .Y(_00552_),
    .B1(net638));
 sg13g2_nand2_1 _26097_ (.Y(_04552_),
    .A(_04510_),
    .B(net28));
 sg13g2_and2_1 _26098_ (.A(net1002),
    .B(\max7219.row_data[7] ),
    .X(_04553_));
 sg13g2_o21ai_1 _26099_ (.B1(_04553_),
    .Y(_04555_),
    .A1(_04260_),
    .A2(_04539_));
 sg13g2_o21ai_1 _26100_ (.B1(_04293_),
    .Y(_04556_),
    .A1(net181),
    .A2(_04514_));
 sg13g2_a21oi_1 _26101_ (.A1(net1061),
    .A2(_04556_),
    .Y(_04557_),
    .B1(\max7219.row_data[7] ));
 sg13g2_nand2b_1 _26102_ (.Y(_04558_),
    .B(net356),
    .A_N(_04557_));
 sg13g2_a21oi_1 _26103_ (.A1(_04552_),
    .A2(_04555_),
    .Y(_00553_),
    .B1(_04558_));
 sg13g2_nand2b_1 _26104_ (.Y(_04559_),
    .B(_04281_),
    .A_N(_13300_));
 sg13g2_nand2_1 _26105_ (.Y(_04560_),
    .A(net312),
    .B(_13053_));
 sg13g2_a21oi_1 _26106_ (.A1(_04297_),
    .A2(_04559_),
    .Y(_00554_),
    .B1(_04560_));
 sg13g2_nor2_1 _26107_ (.A(_00969_),
    .B(_00904_),
    .Y(_04561_));
 sg13g2_nand4_1 _26108_ (.B(_00004_),
    .C(_00023_),
    .A(_13020_),
    .Y(_04562_),
    .D(_04561_));
 sg13g2_buf_1 _26109_ (.A(_04562_),
    .X(_04564_));
 sg13g2_a21oi_1 _26110_ (.A1(net1055),
    .A2(_04564_),
    .Y(_04565_),
    .B1(net715));
 sg13g2_inv_1 _26111_ (.Y(_04566_),
    .A(_13020_));
 sg13g2_inv_1 _26112_ (.Y(_04567_),
    .A(net1055));
 sg13g2_nand3_1 _26113_ (.B(_04566_),
    .C(_00023_),
    .A(\max7219.spi_start ),
    .Y(_04568_));
 sg13g2_nand2_1 _26114_ (.Y(_04569_),
    .A(_04564_),
    .B(_04568_));
 sg13g2_buf_2 _26115_ (.A(_04569_),
    .X(_04570_));
 sg13g2_o21ai_1 _26116_ (.B1(_04570_),
    .Y(_04571_),
    .A1(_04566_),
    .A2(_04567_));
 sg13g2_nand2_1 _26117_ (.Y(_00555_),
    .A(_04565_),
    .B(_04571_));
 sg13g2_nor2b_1 _26118_ (.A(_00990_),
    .B_N(_01001_),
    .Y(_04572_));
 sg13g2_nor2_1 _26119_ (.A(_04567_),
    .B(net1192),
    .Y(_04574_));
 sg13g2_a21oi_1 _26120_ (.A1(_04570_),
    .A2(_04572_),
    .Y(_04575_),
    .B1(_04574_));
 sg13g2_nor2_1 _26121_ (.A(_04238_),
    .B(_04575_),
    .Y(_04576_));
 sg13g2_nor2_1 _26122_ (.A(net1192),
    .B(_04570_),
    .Y(_04577_));
 sg13g2_o21ai_1 _26123_ (.B1(net378),
    .Y(_00556_),
    .A1(_04576_),
    .A2(_04577_));
 sg13g2_nor2_1 _26124_ (.A(net1055),
    .B(net1192),
    .Y(_04578_));
 sg13g2_nand3_1 _26125_ (.B(_04570_),
    .C(_04578_),
    .A(_00936_),
    .Y(_04579_));
 sg13g2_or2_1 _26126_ (.X(_04580_),
    .B(_04578_),
    .A(_00936_));
 sg13g2_a21oi_1 _26127_ (.A1(_04579_),
    .A2(_04580_),
    .Y(_04581_),
    .B1(_04238_));
 sg13g2_nor2_1 _26128_ (.A(_00936_),
    .B(_04570_),
    .Y(_04582_));
 sg13g2_o21ai_1 _26129_ (.B1(net378),
    .Y(_00557_),
    .A1(_04581_),
    .A2(_04582_));
 sg13g2_nor3_1 _26130_ (.A(net1055),
    .B(net1192),
    .C(_00936_),
    .Y(_04584_));
 sg13g2_nand3_1 _26131_ (.B(_04570_),
    .C(_04584_),
    .A(_00947_),
    .Y(_04585_));
 sg13g2_or2_1 _26132_ (.X(_04586_),
    .B(_04584_),
    .A(_00947_));
 sg13g2_a21oi_1 _26133_ (.A1(_04585_),
    .A2(_04586_),
    .Y(_04587_),
    .B1(_04238_));
 sg13g2_nor2_1 _26134_ (.A(_00947_),
    .B(_04570_),
    .Y(_04588_));
 sg13g2_o21ai_1 _26135_ (.B1(net378),
    .Y(_00558_),
    .A1(_04587_),
    .A2(_04588_));
 sg13g2_nand2_1 _26136_ (.Y(_04589_),
    .A(_04279_),
    .B(_00030_));
 sg13g2_inv_1 _26137_ (.Y(_04590_),
    .A(_00030_));
 sg13g2_a221oi_1 _26138_ (.B2(_04590_),
    .C1(_04567_),
    .B1(_00755_),
    .A1(_13191_),
    .Y(_04591_),
    .A2(\max7219.row_data[4] ));
 sg13g2_a221oi_1 _26139_ (.B2(_13191_),
    .C1(_00990_),
    .B1(\max7219.row_data[5] ),
    .A1(net1193),
    .Y(_04593_),
    .A2(_00723_));
 sg13g2_o21ai_1 _26140_ (.B1(_01001_),
    .Y(_04594_),
    .A1(_04591_),
    .A2(_04593_));
 sg13g2_a221oi_1 _26141_ (.B2(_13289_),
    .C1(\max7219.spim.bit_index[1] ),
    .B1(_04567_),
    .A1(net1193),
    .Y(_04595_),
    .A2(_00723_));
 sg13g2_mux2_1 _26142_ (.A0(\max7219.row_data[7] ),
    .A1(\max7219.row_data[6] ),
    .S(_00979_),
    .X(_04596_));
 sg13g2_nand2_1 _26143_ (.Y(_04597_),
    .A(_13191_),
    .B(_04596_));
 sg13g2_a21oi_1 _26144_ (.A1(_04595_),
    .A2(_04597_),
    .Y(_04598_),
    .B1(_00936_));
 sg13g2_nand3_1 _26145_ (.B(_04594_),
    .C(_04598_),
    .A(_04589_),
    .Y(_04599_));
 sg13g2_nand2b_1 _26146_ (.Y(_04600_),
    .B(_04599_),
    .A_N(net1058));
 sg13g2_mux4_1 _26147_ (.S0(net1055),
    .A0(\max7219.row_data[3] ),
    .A1(\max7219.row_data[2] ),
    .A2(\max7219.row_data[1] ),
    .A3(\max7219.row_data[0] ),
    .S1(net1192),
    .X(_04601_));
 sg13g2_a22oi_1 _26148_ (.Y(_04602_),
    .B1(_04601_),
    .B2(_00936_),
    .A2(_04598_),
    .A1(_04594_));
 sg13g2_nor2_1 _26149_ (.A(_00947_),
    .B(_04602_),
    .Y(_04604_));
 sg13g2_nand2b_1 _26150_ (.Y(_04605_),
    .B(_04269_),
    .A_N(_00734_));
 sg13g2_nand4_1 _26151_ (.B(_04329_),
    .C(_04572_),
    .A(_00028_),
    .Y(_04606_),
    .D(_04605_));
 sg13g2_nand2_1 _26152_ (.Y(_04607_),
    .A(_04324_),
    .B(_04323_));
 sg13g2_a22oi_1 _26153_ (.Y(_04608_),
    .B1(_04607_),
    .B2(net1058),
    .A2(_04276_),
    .A1(_04590_));
 sg13g2_and2_1 _26154_ (.A(_04574_),
    .B(_04608_),
    .X(_04609_));
 sg13g2_nand3b_1 _26155_ (.B(_13213_),
    .C(_13235_),
    .Y(_04610_),
    .A_N(_00031_));
 sg13g2_nand3_1 _26156_ (.B(net1192),
    .C(_04610_),
    .A(net1055),
    .Y(_04611_));
 sg13g2_a21oi_1 _26157_ (.A1(net1058),
    .A2(_04611_),
    .Y(_04612_),
    .B1(_04589_));
 sg13g2_nand2_1 _26158_ (.Y(_04613_),
    .A(_00947_),
    .B(_00029_));
 sg13g2_nor2_1 _26159_ (.A(_00030_),
    .B(_00755_),
    .Y(_04615_));
 sg13g2_nor4_1 _26160_ (.A(net1055),
    .B(net1192),
    .C(_04316_),
    .D(_04615_),
    .Y(_04616_));
 sg13g2_nor4_1 _26161_ (.A(_04609_),
    .B(_04612_),
    .C(_04613_),
    .D(_04616_),
    .Y(_04617_));
 sg13g2_a22oi_1 _26162_ (.Y(_04618_),
    .B1(_04606_),
    .B2(_04617_),
    .A2(_04604_),
    .A1(_04600_));
 sg13g2_nand2_1 _26163_ (.Y(_04619_),
    .A(\max7219.o_mosi ),
    .B(_04564_));
 sg13g2_o21ai_1 _26164_ (.B1(_04619_),
    .Y(_04620_),
    .A1(_04564_),
    .A2(_04618_));
 sg13g2_and2_1 _26165_ (.A(net378),
    .B(_04620_),
    .X(_00563_));
 sg13g2_o21ai_1 _26166_ (.B1(_00777_),
    .Y(_04621_),
    .A1(_04241_),
    .A2(_01440_));
 sg13g2_buf_1 _26167_ (.A(_04621_),
    .X(_04622_));
 sg13g2_buf_1 _26168_ (.A(_04622_),
    .X(_04623_));
 sg13g2_xnor2_1 _26169_ (.Y(_04625_),
    .A(net1191),
    .B(_01408_));
 sg13g2_nor2_1 _26170_ (.A(net64),
    .B(_04625_),
    .Y(_00565_));
 sg13g2_inv_1 _26171_ (.Y(_04626_),
    .A(\silife_demo_inst.counter[9] ));
 sg13g2_and3_1 _26172_ (.X(_04627_),
    .A(_01365_),
    .B(\silife_demo_inst.counter[7] ),
    .C(_01215_));
 sg13g2_and4_1 _26173_ (.A(net1191),
    .B(_01204_),
    .C(_01408_),
    .D(\silife_demo_inst.counter[2] ),
    .X(_04628_));
 sg13g2_buf_1 _26174_ (.A(_04628_),
    .X(_04629_));
 sg13g2_nand4_1 _26175_ (.B(_01386_),
    .C(_04627_),
    .A(\silife_demo_inst.counter[8] ),
    .Y(_04630_),
    .D(_04629_));
 sg13g2_buf_1 _26176_ (.A(_04630_),
    .X(_04631_));
 sg13g2_nor2_2 _26177_ (.A(_04626_),
    .B(_04631_),
    .Y(_04632_));
 sg13g2_xnor2_1 _26178_ (.Y(_04633_),
    .A(_01118_),
    .B(_04632_));
 sg13g2_nor2_1 _26179_ (.A(net64),
    .B(_04633_),
    .Y(_00566_));
 sg13g2_nand2_1 _26180_ (.Y(_04635_),
    .A(_01118_),
    .B(_04632_));
 sg13g2_xnor2_1 _26181_ (.Y(_04636_),
    .A(_01290_),
    .B(_04635_));
 sg13g2_nor2_1 _26182_ (.A(net64),
    .B(_04636_),
    .Y(_00567_));
 sg13g2_and3_1 _26183_ (.X(_04637_),
    .A(_01118_),
    .B(\silife_demo_inst.counter[11] ),
    .C(_04632_));
 sg13g2_buf_1 _26184_ (.A(_04637_),
    .X(_04638_));
 sg13g2_xnor2_1 _26185_ (.Y(_04639_),
    .A(_01312_),
    .B(_04638_));
 sg13g2_nor2_1 _26186_ (.A(net64),
    .B(_04639_),
    .Y(_00568_));
 sg13g2_nand2_1 _26187_ (.Y(_04640_),
    .A(_01312_),
    .B(_04638_));
 sg13g2_xor2_1 _26188_ (.B(_04640_),
    .A(_01301_),
    .X(_04641_));
 sg13g2_nor2_1 _26189_ (.A(net64),
    .B(_04641_),
    .Y(_00569_));
 sg13g2_nand3_1 _26190_ (.B(_01312_),
    .C(_04638_),
    .A(_01301_),
    .Y(_04643_));
 sg13g2_xor2_1 _26191_ (.B(_04643_),
    .A(_01344_),
    .X(_04644_));
 sg13g2_nor2_1 _26192_ (.A(net64),
    .B(_04644_),
    .Y(_00570_));
 sg13g2_and4_1 _26193_ (.A(_01118_),
    .B(\silife_demo_inst.counter[11] ),
    .C(_01301_),
    .D(_01312_),
    .X(_04645_));
 sg13g2_nand3_1 _26194_ (.B(_04632_),
    .C(_04645_),
    .A(_01344_),
    .Y(_04646_));
 sg13g2_xor2_1 _26195_ (.B(_04646_),
    .A(\silife_demo_inst.counter[15] ),
    .X(_04647_));
 sg13g2_nor2_1 _26196_ (.A(net64),
    .B(_04647_),
    .Y(_00571_));
 sg13g2_nand3_1 _26197_ (.B(_01344_),
    .C(_04645_),
    .A(\silife_demo_inst.counter[15] ),
    .Y(_04648_));
 sg13g2_nor3_2 _26198_ (.A(_04626_),
    .B(_04631_),
    .C(_04648_),
    .Y(_04649_));
 sg13g2_xnor2_1 _26199_ (.Y(_04651_),
    .A(_01268_),
    .B(_04649_));
 sg13g2_nor2_1 _26200_ (.A(_04623_),
    .B(_04651_),
    .Y(_00572_));
 sg13g2_nand2_1 _26201_ (.Y(_04652_),
    .A(_01268_),
    .B(_04649_));
 sg13g2_xor2_1 _26202_ (.B(_04652_),
    .A(_01258_),
    .X(_04653_));
 sg13g2_nor2_1 _26203_ (.A(_04623_),
    .B(_04653_),
    .Y(_00573_));
 sg13g2_buf_1 _26204_ (.A(_04622_),
    .X(_04654_));
 sg13g2_and3_1 _26205_ (.X(_04655_),
    .A(_01258_),
    .B(_01268_),
    .C(_04649_));
 sg13g2_buf_1 _26206_ (.A(_04655_),
    .X(_04656_));
 sg13g2_xnor2_1 _26207_ (.Y(_04657_),
    .A(_01096_),
    .B(_04656_));
 sg13g2_nor2_1 _26208_ (.A(net63),
    .B(_04657_),
    .Y(_00574_));
 sg13g2_nand2_1 _26209_ (.Y(_04659_),
    .A(_01096_),
    .B(_04656_));
 sg13g2_xor2_1 _26210_ (.B(_04659_),
    .A(_01086_),
    .X(_04660_));
 sg13g2_nor2_1 _26211_ (.A(net63),
    .B(_04660_),
    .Y(_00575_));
 sg13g2_nand2_1 _26212_ (.Y(_04661_),
    .A(net1191),
    .B(_01408_));
 sg13g2_xor2_1 _26213_ (.B(_04661_),
    .A(_01204_),
    .X(_04662_));
 sg13g2_nor2_1 _26214_ (.A(_04654_),
    .B(_04662_),
    .Y(_00576_));
 sg13g2_nand3_1 _26215_ (.B(_01096_),
    .C(_04656_),
    .A(_01086_),
    .Y(_04663_));
 sg13g2_xor2_1 _26216_ (.B(_04663_),
    .A(\silife_demo_inst.counter[20] ),
    .X(_04664_));
 sg13g2_nor2_1 _26217_ (.A(net63),
    .B(_04664_),
    .Y(_00577_));
 sg13g2_nand4_1 _26218_ (.B(_01096_),
    .C(\silife_demo_inst.counter[20] ),
    .A(_01086_),
    .Y(_04665_),
    .D(_04656_));
 sg13g2_xor2_1 _26219_ (.B(_04665_),
    .A(\silife_demo_inst.counter[21] ),
    .X(_04667_));
 sg13g2_nor2_1 _26220_ (.A(net63),
    .B(_04667_),
    .Y(_00578_));
 sg13g2_and4_1 _26221_ (.A(_01258_),
    .B(_01268_),
    .C(_01107_),
    .D(_04649_),
    .X(_04668_));
 sg13g2_buf_1 _26222_ (.A(_04668_),
    .X(_04669_));
 sg13g2_xnor2_1 _26223_ (.Y(_04670_),
    .A(_01354_),
    .B(_04669_));
 sg13g2_nor2_1 _26224_ (.A(net63),
    .B(_04670_),
    .Y(_00579_));
 sg13g2_nand2_1 _26225_ (.Y(_04671_),
    .A(_01354_),
    .B(_04669_));
 sg13g2_xor2_1 _26226_ (.B(_04671_),
    .A(_01247_),
    .X(_04672_));
 sg13g2_nor2_1 _26227_ (.A(net63),
    .B(_04672_),
    .Y(_00580_));
 sg13g2_nand3_1 _26228_ (.B(_01354_),
    .C(_04669_),
    .A(_01247_),
    .Y(_04673_));
 sg13g2_xor2_1 _26229_ (.B(_04673_),
    .A(_01129_),
    .X(_04675_));
 sg13g2_nor2_1 _26230_ (.A(net63),
    .B(_04675_),
    .Y(_00581_));
 sg13g2_nand4_1 _26231_ (.B(_01354_),
    .C(_01129_),
    .A(_01247_),
    .Y(_04676_),
    .D(_04669_));
 sg13g2_xor2_1 _26232_ (.B(_04676_),
    .A(\silife_demo_inst.counter[25] ),
    .X(_04677_));
 sg13g2_nor2_1 _26233_ (.A(net63),
    .B(_04677_),
    .Y(_00582_));
 sg13g2_and4_1 _26234_ (.A(_01247_),
    .B(_01354_),
    .C(\silife_demo_inst.counter[25] ),
    .D(_01129_),
    .X(_04678_));
 sg13g2_and2_1 _26235_ (.A(_04669_),
    .B(_04678_),
    .X(_04679_));
 sg13g2_buf_1 _26236_ (.A(_04679_),
    .X(_04680_));
 sg13g2_xnor2_1 _26237_ (.Y(_04681_),
    .A(_01161_),
    .B(_04680_));
 sg13g2_nor2_1 _26238_ (.A(_04654_),
    .B(_04681_),
    .Y(_00583_));
 sg13g2_buf_1 _26239_ (.A(_04622_),
    .X(_04683_));
 sg13g2_nand2_1 _26240_ (.Y(_04684_),
    .A(_01161_),
    .B(_04680_));
 sg13g2_xor2_1 _26241_ (.B(_04684_),
    .A(_01139_),
    .X(_04685_));
 sg13g2_nor2_1 _26242_ (.A(net62),
    .B(_04685_),
    .Y(_00584_));
 sg13g2_nand3_1 _26243_ (.B(_01161_),
    .C(_04680_),
    .A(_01139_),
    .Y(_04686_));
 sg13g2_xor2_1 _26244_ (.B(_04686_),
    .A(\silife_demo_inst.counter[28] ),
    .X(_04687_));
 sg13g2_nor2_1 _26245_ (.A(net62),
    .B(_04687_),
    .Y(_00585_));
 sg13g2_and4_1 _26246_ (.A(_01139_),
    .B(_01161_),
    .C(\silife_demo_inst.counter[28] ),
    .D(_04680_),
    .X(_04688_));
 sg13g2_buf_1 _26247_ (.A(_04688_),
    .X(_04689_));
 sg13g2_xnor2_1 _26248_ (.Y(_04690_),
    .A(_01172_),
    .B(_04689_));
 sg13g2_nor2_1 _26249_ (.A(net62),
    .B(_04690_),
    .Y(_00586_));
 sg13g2_nand3_1 _26250_ (.B(_01204_),
    .C(_01408_),
    .A(net1191),
    .Y(_04692_));
 sg13g2_xor2_1 _26251_ (.B(_04692_),
    .A(\silife_demo_inst.counter[2] ),
    .X(_04693_));
 sg13g2_nor2_1 _26252_ (.A(net62),
    .B(_04693_),
    .Y(_00587_));
 sg13g2_nand2_1 _26253_ (.Y(_04694_),
    .A(_01172_),
    .B(_04689_));
 sg13g2_xor2_1 _26254_ (.B(_04694_),
    .A(\silife_demo_inst.counter[30] ),
    .X(_04695_));
 sg13g2_nor2_1 _26255_ (.A(_04683_),
    .B(_04695_),
    .Y(_00588_));
 sg13g2_nand3_1 _26256_ (.B(\silife_demo_inst.counter[30] ),
    .C(_04689_),
    .A(_01172_),
    .Y(_04696_));
 sg13g2_xor2_1 _26257_ (.B(_04696_),
    .A(\silife_demo_inst.counter[31] ),
    .X(_04697_));
 sg13g2_nor2_1 _26258_ (.A(_04683_),
    .B(_04697_),
    .Y(_00589_));
 sg13g2_xnor2_1 _26259_ (.Y(_04698_),
    .A(\silife_demo_inst.counter[3] ),
    .B(_04629_));
 sg13g2_nor2_1 _26260_ (.A(net62),
    .B(_04698_),
    .Y(_00590_));
 sg13g2_nand2_1 _26261_ (.Y(_04699_),
    .A(\silife_demo_inst.counter[3] ),
    .B(_04629_));
 sg13g2_xor2_1 _26262_ (.B(_04699_),
    .A(\silife_demo_inst.counter[4] ),
    .X(_04700_));
 sg13g2_nor2_1 _26263_ (.A(net62),
    .B(_04700_),
    .Y(_00591_));
 sg13g2_and2_1 _26264_ (.A(_01386_),
    .B(_04629_),
    .X(_04701_));
 sg13g2_buf_1 _26265_ (.A(_04701_),
    .X(_04702_));
 sg13g2_xnor2_1 _26266_ (.Y(_04703_),
    .A(_01365_),
    .B(_04702_));
 sg13g2_nor2_1 _26267_ (.A(net62),
    .B(_04703_),
    .Y(_00592_));
 sg13g2_nand2_1 _26268_ (.Y(_04704_),
    .A(_01365_),
    .B(_04702_));
 sg13g2_xor2_1 _26269_ (.B(_04704_),
    .A(_01215_),
    .X(_04706_));
 sg13g2_nor2_1 _26270_ (.A(net62),
    .B(_04706_),
    .Y(_00593_));
 sg13g2_nand3_1 _26271_ (.B(_01215_),
    .C(_04702_),
    .A(_01365_),
    .Y(_04707_));
 sg13g2_xor2_1 _26272_ (.B(_04707_),
    .A(\silife_demo_inst.counter[7] ),
    .X(_04708_));
 sg13g2_nor2_1 _26273_ (.A(_04622_),
    .B(_04708_),
    .Y(_00594_));
 sg13g2_nand2_1 _26274_ (.Y(_04709_),
    .A(_04627_),
    .B(_04702_));
 sg13g2_xnor2_1 _26275_ (.Y(_04710_),
    .A(\silife_demo_inst.counter[8] ),
    .B(_04709_));
 sg13g2_nor2b_1 _26276_ (.A(net64),
    .B_N(_04710_),
    .Y(_00595_));
 sg13g2_xnor2_1 _26277_ (.Y(_04711_),
    .A(_04626_),
    .B(_04631_));
 sg13g2_nor2_1 _26278_ (.A(_04622_),
    .B(_04711_),
    .Y(_00596_));
 sg13g2_nor2b_1 _26279_ (.A(_03970_),
    .B_N(_04907_),
    .Y(_04713_));
 sg13g2_and2_1 _26280_ (.A(_01742_),
    .B(_04713_),
    .X(_04714_));
 sg13g2_buf_1 _26281_ (.A(\silife_demo_inst.init_done ),
    .X(_04715_));
 sg13g2_a21oi_1 _26282_ (.A1(net1191),
    .A2(_04714_),
    .Y(_04716_),
    .B1(_04715_));
 sg13g2_nor2_1 _26283_ (.A(_04312_),
    .B(_04716_),
    .Y(_00597_));
 sg13g2_nand3b_1 _26284_ (.B(net1191),
    .C(_01503_),
    .Y(_04717_),
    .A_N(_04715_));
 sg13g2_buf_1 _26285_ (.A(_04717_),
    .X(_04718_));
 sg13g2_mux2_1 _26286_ (.A0(_00275_),
    .A1(_01612_),
    .S(_04718_),
    .X(_04719_));
 sg13g2_and2_1 _26287_ (.A(_12999_),
    .B(_04719_),
    .X(_00598_));
 sg13g2_nor2_1 _26288_ (.A(_03002_),
    .B(_04718_),
    .Y(_04720_));
 sg13g2_xnor2_1 _26289_ (.Y(_04722_),
    .A(net1032),
    .B(_04720_));
 sg13g2_nor2_1 _26290_ (.A(net180),
    .B(_04722_),
    .Y(_00599_));
 sg13g2_nor2_1 _26291_ (.A(_03970_),
    .B(_04718_),
    .Y(_04723_));
 sg13g2_xnor2_1 _26292_ (.Y(_04724_),
    .A(_01676_),
    .B(_04723_));
 sg13g2_nor2_1 _26293_ (.A(net180),
    .B(_04724_),
    .Y(_00600_));
 sg13g2_nand2_1 _26294_ (.Y(_04725_),
    .A(net712),
    .B(_04723_));
 sg13g2_xor2_1 _26295_ (.B(_04725_),
    .A(net1052),
    .X(_04726_));
 sg13g2_nor2_1 _26296_ (.A(net180),
    .B(_04726_),
    .Y(_00601_));
 sg13g2_xor2_1 _26297_ (.B(_04713_),
    .A(_00017_),
    .X(_04727_));
 sg13g2_nor2_1 _26298_ (.A(_04718_),
    .B(_04727_),
    .Y(_04728_));
 sg13g2_a21oi_1 _26299_ (.A1(_01742_),
    .A2(_04718_),
    .Y(_04730_),
    .B1(_04728_));
 sg13g2_nor2_1 _26300_ (.A(_04312_),
    .B(_04730_),
    .Y(_00602_));
 sg13g2_nor2_1 _26301_ (.A(_04715_),
    .B(_04714_),
    .Y(_04731_));
 sg13g2_a21oi_1 _26302_ (.A1(_01503_),
    .A2(_04715_),
    .Y(_04732_),
    .B1(_04731_));
 sg13g2_nor2_1 _26303_ (.A(_01075_),
    .B(_04732_),
    .Y(_00604_));
 sg13g2_inv_1 _26304_ (.Y(_04733_),
    .A(wr_available));
 sg13g2_a21oi_1 _26305_ (.A1(_04733_),
    .A2(net7),
    .Y(_00605_),
    .B1(net638));
 sg13g2_buf_2 _26306_ (.A(_13010_),
    .X(_04734_));
 sg13g2_buf_2 _26307_ (.A(_01935_),
    .X(_04735_));
 sg13g2_mux4_1 _26308_ (.S0(net130),
    .A0(net941),
    .A1(net933),
    .A2(net582),
    .A3(net572),
    .S1(net143),
    .X(_04736_));
 sg13g2_mux4_1 _26309_ (.S0(net130),
    .A0(net904),
    .A1(net883),
    .A2(_10244_),
    .A3(net855),
    .S1(net139),
    .X(_04738_));
 sg13g2_buf_2 _26310_ (.A(_01935_),
    .X(_04739_));
 sg13g2_mux4_1 _26311_ (.S0(net129),
    .A0(_11060_),
    .A1(_11057_),
    .A2(_11715_),
    .A3(_11755_),
    .S1(net143),
    .X(_04740_));
 sg13g2_mux4_1 _26312_ (.S0(net129),
    .A0(_12451_),
    .A1(_12492_),
    .A2(_12883_),
    .A3(_03272_),
    .S1(net143),
    .X(_04741_));
 sg13g2_mux4_1 _26313_ (.S0(_05177_),
    .A0(_04736_),
    .A1(_04738_),
    .A2(_04740_),
    .A3(_04741_),
    .S1(_05179_),
    .X(_04742_));
 sg13g2_mux4_1 _26314_ (.S0(net129),
    .A0(net1183),
    .A1(_02475_),
    .A2(_09266_),
    .A3(_01551_),
    .S1(net143),
    .X(_04743_));
 sg13g2_mux4_1 _26315_ (.S0(net129),
    .A0(_01596_),
    .A1(_02429_),
    .A2(net753),
    .A3(net743),
    .S1(net143),
    .X(_04744_));
 sg13g2_mux4_1 _26316_ (.S0(net129),
    .A0(_03175_),
    .A1(_05275_),
    .A2(_05173_),
    .A3(_05215_),
    .S1(_09916_),
    .X(_04745_));
 sg13g2_mux4_1 _26317_ (.S0(net129),
    .A0(net1174),
    .A1(net971),
    .A2(net1167),
    .A3(net953),
    .S1(_09916_),
    .X(_04746_));
 sg13g2_mux4_1 _26318_ (.S0(_05177_),
    .A0(_04743_),
    .A1(_04744_),
    .A2(_04745_),
    .A3(_04746_),
    .S1(_05179_),
    .X(_04747_));
 sg13g2_buf_1 _26319_ (.A(net177),
    .X(_04749_));
 sg13g2_mux2_1 _26320_ (.A0(_04742_),
    .A1(_04747_),
    .S(net94),
    .X(_04750_));
 sg13g2_nor2_1 _26321_ (.A(_13010_),
    .B(_04750_),
    .Y(_04751_));
 sg13g2_a21oi_1 _26322_ (.A1(_04734_),
    .A2(_00712_),
    .Y(net16),
    .B1(_04751_));
 sg13g2_mux4_1 _26323_ (.S0(_04735_),
    .A0(net1042),
    .A1(net711),
    .A2(_09196_),
    .A3(net446),
    .S1(_11407_),
    .X(_04752_));
 sg13g2_mux4_1 _26324_ (.S0(net130),
    .A0(net434),
    .A1(net767),
    .A2(net413),
    .A3(net405),
    .S1(net139),
    .X(_04753_));
 sg13g2_mux4_1 _26325_ (.S0(net130),
    .A0(net396),
    .A1(_03594_),
    .A2(_05401_),
    .A3(net673),
    .S1(net139),
    .X(_04754_));
 sg13g2_mux4_1 _26326_ (.S0(net130),
    .A0(_05698_),
    .A1(net640),
    .A2(net624),
    .A3(net612),
    .S1(net139),
    .X(_04755_));
 sg13g2_mux4_1 _26327_ (.S0(_05177_),
    .A0(_04752_),
    .A1(_04753_),
    .A2(_04754_),
    .A3(_04755_),
    .S1(_05179_),
    .X(_04756_));
 sg13g2_buf_1 _26328_ (.A(net320),
    .X(_04757_));
 sg13g2_mux4_1 _26329_ (.S0(_04739_),
    .A0(net605),
    .A1(net932),
    .A2(net584),
    .A3(net287),
    .S1(net128),
    .X(_04759_));
 sg13g2_mux4_1 _26330_ (.S0(net129),
    .A0(net906),
    .A1(net541),
    .A2(net529),
    .A3(net521),
    .S1(net143),
    .X(_04760_));
 sg13g2_buf_4 _26331_ (.X(_04761_),
    .A(_01935_));
 sg13g2_mux4_1 _26332_ (.S0(_04761_),
    .A0(_10656_),
    .A1(_10999_),
    .A2(_11362_),
    .A3(_11729_),
    .S1(net128),
    .X(_04762_));
 sg13g2_mux4_1 _26333_ (.S0(_04761_),
    .A0(_12154_),
    .A1(net806),
    .A2(net211),
    .A3(net371),
    .S1(net128),
    .X(_04763_));
 sg13g2_mux4_1 _26334_ (.S0(_05177_),
    .A0(_04759_),
    .A1(_04760_),
    .A2(_04762_),
    .A3(_04763_),
    .S1(_05179_),
    .X(_04764_));
 sg13g2_nor2b_1 _26335_ (.A(net94),
    .B_N(_04764_),
    .Y(_04765_));
 sg13g2_a21oi_1 _26336_ (.A1(net94),
    .A2(_04756_),
    .Y(_04766_),
    .B1(_04765_));
 sg13g2_nand2_1 _26337_ (.Y(_04767_),
    .A(net1549),
    .B(\max7219.o_sck ));
 sg13g2_o21ai_1 _26338_ (.B1(_04767_),
    .Y(net17),
    .A1(net1549),
    .A2(_04766_));
 sg13g2_mux4_1 _26339_ (.S0(net130),
    .A0(_04674_),
    .A1(_03756_),
    .A2(net268),
    .A3(net206),
    .S1(net139),
    .X(_04769_));
 sg13g2_mux4_1 _26340_ (.S0(_04735_),
    .A0(net430),
    .A1(net421),
    .A2(net196),
    .A3(net190),
    .S1(net139),
    .X(_04770_));
 sg13g2_mux4_1 _26341_ (.S0(net130),
    .A0(net186),
    .A1(net348),
    .A2(net661),
    .A3(net346),
    .S1(_11407_),
    .X(_04771_));
 sg13g2_mux4_1 _26342_ (.S0(net130),
    .A0(net160),
    .A1(net157),
    .A2(net626),
    .A3(_06905_),
    .S1(net139),
    .X(_04772_));
 sg13g2_mux4_1 _26343_ (.S0(_05177_),
    .A0(_04769_),
    .A1(_04770_),
    .A2(_04771_),
    .A3(_04772_),
    .S1(_05179_),
    .X(_04773_));
 sg13g2_mux4_1 _26344_ (.S0(_04739_),
    .A0(_07335_),
    .A1(net590),
    .A2(net294),
    .A3(net571),
    .S1(net128),
    .X(_04774_));
 sg13g2_mux4_1 _26345_ (.S0(net129),
    .A0(net560),
    .A1(net542),
    .A2(_09976_),
    .A3(_10307_),
    .S1(net143),
    .X(_04775_));
 sg13g2_mux4_1 _26346_ (.S0(_04761_),
    .A0(_10716_),
    .A1(_11100_),
    .A2(_11415_),
    .A3(_11851_),
    .S1(net128),
    .X(_04776_));
 sg13g2_mux4_1 _26347_ (.S0(_04761_),
    .A0(_12212_),
    .A1(net215),
    .A2(_12936_),
    .A3(_04099_),
    .S1(net128),
    .X(_04777_));
 sg13g2_mux4_1 _26348_ (.S0(_05177_),
    .A0(_04774_),
    .A1(_04775_),
    .A2(_04776_),
    .A3(_04777_),
    .S1(_05179_),
    .X(_04778_));
 sg13g2_nor2b_1 _26349_ (.A(net94),
    .B_N(_04778_),
    .Y(_04780_));
 sg13g2_a21oi_1 _26350_ (.A1(net94),
    .A2(_04773_),
    .Y(_04781_),
    .B1(_04780_));
 sg13g2_nand2_1 _26351_ (.Y(_04782_),
    .A(net1549),
    .B(\max7219.o_mosi ));
 sg13g2_o21ai_1 _26352_ (.B1(_04782_),
    .Y(net18),
    .A1(net1549),
    .A2(_04781_));
 sg13g2_buf_2 _26353_ (.A(_04761_),
    .X(_04783_));
 sg13g2_buf_1 _26354_ (.A(net128),
    .X(_04784_));
 sg13g2_mux4_1 _26355_ (.S0(net93),
    .A0(_07428_),
    .A1(net1146),
    .A2(_08178_),
    .A3(net1135),
    .S1(net92),
    .X(_04785_));
 sg13g2_mux4_1 _26356_ (.S0(net93),
    .A0(_08975_),
    .A1(_09706_),
    .A2(_10075_),
    .A3(net1111),
    .S1(net92),
    .X(_04786_));
 sg13g2_buf_2 _26357_ (.A(_04761_),
    .X(_04787_));
 sg13g2_buf_1 _26358_ (.A(net128),
    .X(_04788_));
 sg13g2_mux4_1 _26359_ (.S0(net91),
    .A0(_10844_),
    .A1(_11207_),
    .A2(_11584_),
    .A3(_11928_),
    .S1(net90),
    .X(_04790_));
 sg13g2_mux4_1 _26360_ (.S0(_04787_),
    .A0(_12305_),
    .A1(_12658_),
    .A2(_13029_),
    .A3(_04962_),
    .S1(_04788_),
    .X(_04791_));
 sg13g2_buf_2 _26361_ (.A(_05177_),
    .X(_04792_));
 sg13g2_buf_1 _26362_ (.A(_05179_),
    .X(_04793_));
 sg13g2_mux4_1 _26363_ (.S0(net179),
    .A0(_04785_),
    .A1(_04786_),
    .A2(_04790_),
    .A3(_04791_),
    .S1(net178),
    .X(_04794_));
 sg13g2_buf_2 _26364_ (.A(_04761_),
    .X(_04795_));
 sg13g2_buf_1 _26365_ (.A(_04757_),
    .X(_04796_));
 sg13g2_mux4_1 _26366_ (.S0(net89),
    .A0(net1181),
    .A1(_04870_),
    .A2(_09382_),
    .A3(_00724_),
    .S1(net88),
    .X(_04797_));
 sg13g2_mux4_1 _26367_ (.S0(net89),
    .A0(net1078),
    .A1(_02193_),
    .A2(_02592_),
    .A3(net1066),
    .S1(net88),
    .X(_04798_));
 sg13g2_buf_2 _26368_ (.A(_04761_),
    .X(_04799_));
 sg13g2_buf_1 _26369_ (.A(_04757_),
    .X(_04801_));
 sg13g2_mux4_1 _26370_ (.S0(net87),
    .A0(net1063),
    .A1(_05473_),
    .A2(_05379_),
    .A3(_00042_),
    .S1(net86),
    .X(_04802_));
 sg13g2_mux4_1 _26371_ (.S0(net87),
    .A0(_05916_),
    .A1(_06304_),
    .A2(_06691_),
    .A3(net1160),
    .S1(net86),
    .X(_04803_));
 sg13g2_mux4_1 _26372_ (.S0(net179),
    .A0(_04797_),
    .A1(_04798_),
    .A2(_04802_),
    .A3(_04803_),
    .S1(net178),
    .X(_04804_));
 sg13g2_mux2_1 _26373_ (.A0(_04794_),
    .A1(_04804_),
    .S(net94),
    .X(_04805_));
 sg13g2_nor2_1 _26374_ (.A(_04734_),
    .B(_04805_),
    .Y(net19));
 sg13g2_mux4_1 _26375_ (.S0(net93),
    .A0(_07495_),
    .A1(_07853_),
    .A2(net1140),
    .A3(net1133),
    .S1(net92),
    .X(_04806_));
 sg13g2_mux4_1 _26376_ (.S0(_04783_),
    .A0(_09019_),
    .A1(_09746_),
    .A2(_10131_),
    .A3(_10467_),
    .S1(_04784_),
    .X(_04807_));
 sg13g2_mux4_1 _26377_ (.S0(net91),
    .A0(_10884_),
    .A1(_11232_),
    .A2(_11624_),
    .A3(_11984_),
    .S1(net90),
    .X(_04808_));
 sg13g2_mux4_1 _26378_ (.S0(net91),
    .A0(_12357_),
    .A1(net1087),
    .A2(_13087_),
    .A3(_05030_),
    .S1(net90),
    .X(_04809_));
 sg13g2_mux4_1 _26379_ (.S0(net179),
    .A0(_04806_),
    .A1(_04807_),
    .A2(_04808_),
    .A3(_04809_),
    .S1(net178),
    .X(_04811_));
 sg13g2_mux4_1 _26380_ (.S0(net89),
    .A0(_04857_),
    .A1(_04970_),
    .A2(_09419_),
    .A3(_00763_),
    .S1(net88),
    .X(_04812_));
 sg13g2_mux4_1 _26381_ (.S0(net89),
    .A0(_01852_),
    .A1(_02243_),
    .A2(_02631_),
    .A3(_03037_),
    .S1(net88),
    .X(_04813_));
 sg13g2_mux4_1 _26382_ (.S0(net87),
    .A0(_03434_),
    .A1(_05546_),
    .A2(_05434_),
    .A3(_05484_),
    .S1(net86),
    .X(_04814_));
 sg13g2_mux4_1 _26383_ (.S0(net87),
    .A0(_05951_),
    .A1(net1168),
    .A2(_06721_),
    .A3(_07082_),
    .S1(net86),
    .X(_04815_));
 sg13g2_mux4_1 _26384_ (.S0(net179),
    .A0(_04812_),
    .A1(_04813_),
    .A2(_04814_),
    .A3(_04815_),
    .S1(net178),
    .X(_04816_));
 sg13g2_mux2_1 _26385_ (.A0(_04811_),
    .A1(_04816_),
    .S(net94),
    .X(_04817_));
 sg13g2_nor2_1 _26386_ (.A(net1549),
    .B(_04817_),
    .Y(net20));
 sg13g2_mux4_1 _26387_ (.S0(net93),
    .A0(_07538_),
    .A1(net1144),
    .A2(_08292_),
    .A3(net1131),
    .S1(net92),
    .X(_04818_));
 sg13g2_mux4_1 _26388_ (.S0(_04783_),
    .A0(_09077_),
    .A1(net1119),
    .A2(net869),
    .A3(_10520_),
    .S1(_04784_),
    .X(_04819_));
 sg13g2_mux4_1 _26389_ (.S0(net91),
    .A0(_10944_),
    .A1(_11280_),
    .A2(_11662_),
    .A3(_12021_),
    .S1(net90),
    .X(_04821_));
 sg13g2_mux4_1 _26390_ (.S0(net91),
    .A0(_12392_),
    .A1(_12756_),
    .A2(_13129_),
    .A3(_05096_),
    .S1(net90),
    .X(_04822_));
 sg13g2_mux4_1 _26391_ (.S0(net179),
    .A0(_04818_),
    .A1(_04819_),
    .A2(_04821_),
    .A3(_04822_),
    .S1(net178),
    .X(_04823_));
 sg13g2_mux4_1 _26392_ (.S0(net89),
    .A0(_04946_),
    .A1(_05024_),
    .A2(_00099_),
    .A3(_00827_),
    .S1(net88),
    .X(_04824_));
 sg13g2_mux4_1 _26393_ (.S0(_04795_),
    .A0(_01875_),
    .A1(_02284_),
    .A2(_02692_),
    .A3(_03080_),
    .S1(_04796_),
    .X(_04825_));
 sg13g2_mux4_1 _26394_ (.S0(net87),
    .A0(_03478_),
    .A1(_05575_),
    .A2(_05488_),
    .A3(_05553_),
    .S1(net86),
    .X(_04826_));
 sg13g2_mux4_1 _26395_ (.S0(net87),
    .A0(net974),
    .A1(_06392_),
    .A2(_06784_),
    .A3(_07137_),
    .S1(net86),
    .X(_04827_));
 sg13g2_mux4_1 _26396_ (.S0(net179),
    .A0(_04824_),
    .A1(_04825_),
    .A2(_04826_),
    .A3(_04827_),
    .S1(net178),
    .X(_04828_));
 sg13g2_mux2_1 _26397_ (.A0(_04823_),
    .A1(_04828_),
    .S(_04749_),
    .X(_04829_));
 sg13g2_nor2_1 _26398_ (.A(net1549),
    .B(_04829_),
    .Y(net21));
 sg13g2_mux4_1 _26399_ (.S0(net93),
    .A0(_08270_),
    .A1(_08648_),
    .A2(net1128),
    .A3(_09774_),
    .S1(net92),
    .X(_04831_));
 sg13g2_mux4_1 _26400_ (.S0(net93),
    .A0(net1113),
    .A1(_10533_),
    .A2(_10924_),
    .A3(_11272_),
    .S1(net92),
    .X(_04832_));
 sg13g2_mux4_1 _26401_ (.S0(net91),
    .A0(_11644_),
    .A1(_12003_),
    .A2(_12374_),
    .A3(_12759_),
    .S1(net90),
    .X(_04833_));
 sg13g2_mux4_1 _26402_ (.S0(_04787_),
    .A0(_13114_),
    .A1(_01137_),
    .A2(_01428_),
    .A3(_00158_),
    .S1(_04788_),
    .X(_04834_));
 sg13g2_mux4_1 _26403_ (.S0(net179),
    .A0(_04831_),
    .A1(_04832_),
    .A2(_04833_),
    .A3(_04834_),
    .S1(net178),
    .X(_04835_));
 sg13g2_mux4_1 _26404_ (.S0(net89),
    .A0(_05010_),
    .A1(_05102_),
    .A2(_01878_),
    .A3(net1074),
    .S1(net88),
    .X(_04836_));
 sg13g2_mux4_1 _26405_ (.S0(net89),
    .A0(_02672_),
    .A1(net1065),
    .A2(_03490_),
    .A3(_03830_),
    .S1(net88),
    .X(_04837_));
 sg13g2_mux4_1 _26406_ (.S0(_04799_),
    .A0(_04121_),
    .A1(_00136_),
    .A2(_05530_),
    .A3(_05601_),
    .S1(_04801_),
    .X(_04838_));
 sg13g2_mux4_1 _26407_ (.S0(net87),
    .A0(_06767_),
    .A1(_07119_),
    .A2(_07520_),
    .A3(_07894_),
    .S1(net86),
    .X(_04839_));
 sg13g2_mux4_1 _26408_ (.S0(_04792_),
    .A0(_04836_),
    .A1(_04837_),
    .A2(_04838_),
    .A3(_04839_),
    .S1(_04793_),
    .X(_04840_));
 sg13g2_mux2_1 _26409_ (.A0(_04835_),
    .A1(_04840_),
    .S(_04749_),
    .X(_04842_));
 sg13g2_nor2_1 _26410_ (.A(net1549),
    .B(_04842_),
    .Y(net22));
 sg13g2_mux4_1 _26411_ (.S0(net93),
    .A0(_00177_),
    .A1(_00176_),
    .A2(_00179_),
    .A3(_00178_),
    .S1(net92),
    .X(_04843_));
 sg13g2_mux4_1 _26412_ (.S0(net93),
    .A0(_00181_),
    .A1(_00180_),
    .A2(_00183_),
    .A3(_00182_),
    .S1(net92),
    .X(_04844_));
 sg13g2_mux4_1 _26413_ (.S0(net91),
    .A0(_00185_),
    .A1(_00184_),
    .A2(_00187_),
    .A3(_00186_),
    .S1(net90),
    .X(_04845_));
 sg13g2_mux4_1 _26414_ (.S0(net91),
    .A0(_00189_),
    .A1(_00188_),
    .A2(_01246_),
    .A3(_00190_),
    .S1(net90),
    .X(_04846_));
 sg13g2_mux4_1 _26415_ (.S0(net179),
    .A0(_04843_),
    .A1(_04844_),
    .A2(_04845_),
    .A3(_04846_),
    .S1(net178),
    .X(_04847_));
 sg13g2_mux4_1 _26416_ (.S0(net89),
    .A0(_02410_),
    .A1(_00160_),
    .A2(_00163_),
    .A3(_00162_),
    .S1(net88),
    .X(_04848_));
 sg13g2_mux4_1 _26417_ (.S0(_04795_),
    .A0(_00165_),
    .A1(_00164_),
    .A2(_00167_),
    .A3(_00166_),
    .S1(_04796_),
    .X(_04849_));
 sg13g2_mux4_1 _26418_ (.S0(_04799_),
    .A0(_03923_),
    .A1(_00168_),
    .A2(_05233_),
    .A3(_00170_),
    .S1(_04801_),
    .X(_04850_));
 sg13g2_mux4_1 _26419_ (.S0(net87),
    .A0(_00173_),
    .A1(_00172_),
    .A2(_00175_),
    .A3(_00174_),
    .S1(net86),
    .X(_04852_));
 sg13g2_mux4_1 _26420_ (.S0(_04792_),
    .A0(_04848_),
    .A1(_04849_),
    .A2(_04850_),
    .A3(_04852_),
    .S1(_04793_),
    .X(_04853_));
 sg13g2_mux2_1 _26421_ (.A0(_04847_),
    .A1(_04853_),
    .S(net94),
    .X(_04854_));
 sg13g2_nor2_1 _26422_ (.A(net1549),
    .B(_04854_),
    .Y(net23));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi \demo_mode$_SDFFE_PN0P__1214  (.L_HI(net1214));
 sg13g2_buf_1 _26425_ (.A(net1198),
    .X(uio_oe[0]));
 sg13g2_buf_1 _26426_ (.A(net1199),
    .X(uio_oe[1]));
 sg13g2_buf_1 _26427_ (.A(net1200),
    .X(uio_oe[2]));
 sg13g2_buf_1 _26428_ (.A(net1201),
    .X(uio_oe[3]));
 sg13g2_buf_1 _26429_ (.A(net1202),
    .X(uio_oe[4]));
 sg13g2_buf_1 _26430_ (.A(net1203),
    .X(uio_oe[5]));
 sg13g2_buf_1 _26431_ (.A(net1204),
    .X(uio_oe[6]));
 sg13g2_buf_1 _26432_ (.A(net1205),
    .X(uio_oe[7]));
 sg13g2_buf_1 _26433_ (.A(net1206),
    .X(uio_out[0]));
 sg13g2_buf_1 _26434_ (.A(net1207),
    .X(uio_out[1]));
 sg13g2_buf_1 _26435_ (.A(net1208),
    .X(uio_out[2]));
 sg13g2_buf_1 _26436_ (.A(net1209),
    .X(uio_out[3]));
 sg13g2_buf_1 _26437_ (.A(net1210),
    .X(uio_out[4]));
 sg13g2_buf_1 _26438_ (.A(net1211),
    .X(uio_out[5]));
 sg13g2_buf_1 _26439_ (.A(net1212),
    .X(uio_out[6]));
 sg13g2_buf_1 _26440_ (.A(net1213),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \demo_mode$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1214),
    .D(_00276_),
    .Q_N(_13372_),
    .Q(demo_mode));
 sg13g2_dfrbp_1 \grid.cell_0_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1215),
    .D(_00277_),
    .Q_N(_13371_),
    .Q(\grid.cell_0_0.out ));
 sg13g2_dfrbp_1 \grid.cell_0_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1216),
    .D(_00278_),
    .Q_N(_00219_),
    .Q(\grid.cell_0_0.e ));
 sg13g2_dfrbp_1 \grid.cell_0_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1217),
    .D(_00279_),
    .Q_N(_00216_),
    .Q(\grid.cell_0_1.e ));
 sg13g2_dfrbp_1 \grid.cell_0_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1218),
    .D(_00280_),
    .Q_N(_00033_),
    .Q(\grid.cell_0_2.e ));
 sg13g2_dfrbp_1 \grid.cell_0_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1219),
    .D(_00281_),
    .Q_N(_00065_),
    .Q(\grid.cell_0_3.e ));
 sg13g2_dfrbp_1 \grid.cell_0_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1220),
    .D(_00282_),
    .Q_N(_00097_),
    .Q(\grid.cell_0_4.e ));
 sg13g2_dfrbp_1 \grid.cell_0_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1221),
    .D(_00283_),
    .Q_N(_00129_),
    .Q(\grid.cell_0_5.e ));
 sg13g2_dfrbp_1 \grid.cell_0_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1222),
    .D(_00284_),
    .Q_N(_00161_),
    .Q(\grid.cell_0_0.w ));
 sg13g2_dfrbp_1 \grid.cell_10_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1223),
    .D(_00285_),
    .Q_N(_13370_),
    .Q(\grid.cell_10_0.out ));
 sg13g2_dfrbp_1 \grid.cell_10_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1224),
    .D(_00286_),
    .Q_N(_00246_),
    .Q(\grid.cell_10_0.e ));
 sg13g2_dfrbp_1 \grid.cell_10_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1225),
    .D(_00287_),
    .Q_N(_00245_),
    .Q(\grid.cell_10_1.e ));
 sg13g2_dfrbp_1 \grid.cell_10_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1226),
    .D(_00288_),
    .Q_N(_00043_),
    .Q(\grid.cell_10_2.e ));
 sg13g2_dfrbp_1 \grid.cell_10_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1227),
    .D(_00289_),
    .Q_N(_00075_),
    .Q(\grid.cell_10_3.e ));
 sg13g2_dfrbp_1 \grid.cell_10_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1228),
    .D(_00290_),
    .Q_N(_00107_),
    .Q(\grid.cell_10_4.e ));
 sg13g2_dfrbp_1 \grid.cell_10_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1229),
    .D(_00291_),
    .Q_N(_00139_),
    .Q(\grid.cell_10_5.e ));
 sg13g2_dfrbp_1 \grid.cell_10_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1230),
    .D(_00292_),
    .Q_N(_00171_),
    .Q(\grid.cell_10_0.w ));
 sg13g2_dfrbp_1 \grid.cell_11_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1231),
    .D(_00293_),
    .Q_N(_00244_),
    .Q(\grid.cell_10_0.s ));
 sg13g2_dfrbp_1 \grid.cell_11_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1232),
    .D(_00294_),
    .Q_N(_00243_),
    .Q(\grid.cell_10_0.se ));
 sg13g2_dfrbp_1 \grid.cell_11_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1233),
    .D(_00295_),
    .Q_N(_00242_),
    .Q(\grid.cell_10_1.se ));
 sg13g2_dfrbp_1 \grid.cell_11_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1234),
    .D(_00296_),
    .Q_N(_00042_),
    .Q(\grid.cell_10_2.se ));
 sg13g2_dfrbp_1 \grid.cell_11_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1235),
    .D(_00297_),
    .Q_N(_00074_),
    .Q(\grid.cell_10_3.se ));
 sg13g2_dfrbp_1 \grid.cell_11_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1236),
    .D(_00298_),
    .Q_N(_00106_),
    .Q(\grid.cell_10_4.se ));
 sg13g2_dfrbp_1 \grid.cell_11_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1237),
    .D(_00299_),
    .Q_N(_00138_),
    .Q(\grid.cell_10_5.se ));
 sg13g2_dfrbp_1 \grid.cell_11_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1238),
    .D(_00300_),
    .Q_N(_00170_),
    .Q(\grid.cell_10_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_12_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1239),
    .D(_00301_),
    .Q_N(_00241_),
    .Q(\grid.cell_11_0.s ));
 sg13g2_dfrbp_1 \grid.cell_12_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1240),
    .D(_00302_),
    .Q_N(_00240_),
    .Q(\grid.cell_11_0.se ));
 sg13g2_dfrbp_1 \grid.cell_12_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1241),
    .D(_00303_),
    .Q_N(_00239_),
    .Q(\grid.cell_11_1.se ));
 sg13g2_dfrbp_1 \grid.cell_12_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1242),
    .D(_00304_),
    .Q_N(_00045_),
    .Q(\grid.cell_11_2.se ));
 sg13g2_dfrbp_1 \grid.cell_12_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1243),
    .D(_00305_),
    .Q_N(_00077_),
    .Q(\grid.cell_11_3.se ));
 sg13g2_dfrbp_1 \grid.cell_12_5.state$_SDFFE_PP0P_  (.CLK(clknet_4_11__leaf_clk),
    .RESET_B(net1244),
    .D(_00306_),
    .Q_N(_00109_),
    .Q(\grid.cell_11_4.se ));
 sg13g2_dfrbp_1 \grid.cell_12_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1245),
    .D(_00307_),
    .Q_N(_00141_),
    .Q(\grid.cell_11_5.se ));
 sg13g2_dfrbp_1 \grid.cell_12_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1246),
    .D(_00308_),
    .Q_N(_00173_),
    .Q(\grid.cell_11_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_13_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1247),
    .D(_00309_),
    .Q_N(_00238_),
    .Q(\grid.cell_12_0.s ));
 sg13g2_dfrbp_1 \grid.cell_13_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1248),
    .D(_00310_),
    .Q_N(_00237_),
    .Q(\grid.cell_12_0.se ));
 sg13g2_dfrbp_1 \grid.cell_13_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1249),
    .D(_00311_),
    .Q_N(_00236_),
    .Q(\grid.cell_12_1.se ));
 sg13g2_dfrbp_1 \grid.cell_13_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1250),
    .D(_00312_),
    .Q_N(_00044_),
    .Q(\grid.cell_12_2.se ));
 sg13g2_dfrbp_1 \grid.cell_13_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1251),
    .D(_00313_),
    .Q_N(_00076_),
    .Q(\grid.cell_12_3.se ));
 sg13g2_dfrbp_1 \grid.cell_13_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1252),
    .D(_00314_),
    .Q_N(_00108_),
    .Q(\grid.cell_12_4.se ));
 sg13g2_dfrbp_1 \grid.cell_13_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1253),
    .D(_00315_),
    .Q_N(_00140_),
    .Q(\grid.cell_12_5.se ));
 sg13g2_dfrbp_1 \grid.cell_13_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1254),
    .D(_00316_),
    .Q_N(_00172_),
    .Q(\grid.cell_12_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_14_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1255),
    .D(_00317_),
    .Q_N(_00235_),
    .Q(\grid.cell_13_0.s ));
 sg13g2_dfrbp_1 \grid.cell_14_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1256),
    .D(_00318_),
    .Q_N(_00234_),
    .Q(\grid.cell_13_0.se ));
 sg13g2_dfrbp_1 \grid.cell_14_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1257),
    .D(_00319_),
    .Q_N(_00233_),
    .Q(\grid.cell_13_1.se ));
 sg13g2_dfrbp_1 \grid.cell_14_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1258),
    .D(_00320_),
    .Q_N(_00047_),
    .Q(\grid.cell_13_2.se ));
 sg13g2_dfrbp_1 \grid.cell_14_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1259),
    .D(_00321_),
    .Q_N(_00079_),
    .Q(\grid.cell_13_3.se ));
 sg13g2_dfrbp_1 \grid.cell_14_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1260),
    .D(_00322_),
    .Q_N(_00111_),
    .Q(\grid.cell_13_4.se ));
 sg13g2_dfrbp_1 \grid.cell_14_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1261),
    .D(_00323_),
    .Q_N(_00143_),
    .Q(\grid.cell_13_5.se ));
 sg13g2_dfrbp_1 \grid.cell_14_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1262),
    .D(_00324_),
    .Q_N(_00175_),
    .Q(\grid.cell_13_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_15_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1263),
    .D(_00325_),
    .Q_N(_00232_),
    .Q(\grid.cell_14_0.s ));
 sg13g2_dfrbp_1 \grid.cell_15_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1264),
    .D(_00326_),
    .Q_N(_00231_),
    .Q(\grid.cell_14_0.se ));
 sg13g2_dfrbp_1 \grid.cell_15_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1265),
    .D(_00327_),
    .Q_N(_00230_),
    .Q(\grid.cell_14_1.se ));
 sg13g2_dfrbp_1 \grid.cell_15_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1266),
    .D(_00328_),
    .Q_N(_00046_),
    .Q(\grid.cell_14_2.se ));
 sg13g2_dfrbp_1 \grid.cell_15_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1267),
    .D(_00329_),
    .Q_N(_00078_),
    .Q(\grid.cell_14_3.se ));
 sg13g2_dfrbp_1 \grid.cell_15_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1268),
    .D(_00330_),
    .Q_N(_00110_),
    .Q(\grid.cell_14_4.se ));
 sg13g2_dfrbp_1 \grid.cell_15_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1269),
    .D(_00331_),
    .Q_N(_00142_),
    .Q(\grid.cell_14_5.se ));
 sg13g2_dfrbp_1 \grid.cell_15_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1270),
    .D(_00332_),
    .Q_N(_00174_),
    .Q(\grid.cell_14_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_16_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1271),
    .D(_00333_),
    .Q_N(_00229_),
    .Q(\grid.cell_15_0.s ));
 sg13g2_dfrbp_1 \grid.cell_16_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1272),
    .D(_00334_),
    .Q_N(_00228_),
    .Q(\grid.cell_15_0.se ));
 sg13g2_dfrbp_1 \grid.cell_16_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1273),
    .D(_00335_),
    .Q_N(_00227_),
    .Q(\grid.cell_15_1.se ));
 sg13g2_dfrbp_1 \grid.cell_16_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1274),
    .D(_00336_),
    .Q_N(_00049_),
    .Q(\grid.cell_15_2.se ));
 sg13g2_dfrbp_1 \grid.cell_16_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1275),
    .D(_00337_),
    .Q_N(_00081_),
    .Q(\grid.cell_15_3.se ));
 sg13g2_dfrbp_1 \grid.cell_16_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1276),
    .D(_00338_),
    .Q_N(_00113_),
    .Q(\grid.cell_15_4.se ));
 sg13g2_dfrbp_1 \grid.cell_16_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1277),
    .D(_00339_),
    .Q_N(_00145_),
    .Q(\grid.cell_15_5.se ));
 sg13g2_dfrbp_1 \grid.cell_16_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1278),
    .D(_00340_),
    .Q_N(_00177_),
    .Q(\grid.cell_15_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_17_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1279),
    .D(_00341_),
    .Q_N(_00226_),
    .Q(\grid.cell_16_0.s ));
 sg13g2_dfrbp_1 \grid.cell_17_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1280),
    .D(_00342_),
    .Q_N(_00225_),
    .Q(\grid.cell_16_0.se ));
 sg13g2_dfrbp_1 \grid.cell_17_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1281),
    .D(_00343_),
    .Q_N(_00224_),
    .Q(\grid.cell_16_1.se ));
 sg13g2_dfrbp_1 \grid.cell_17_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1282),
    .D(_00344_),
    .Q_N(_00048_),
    .Q(\grid.cell_16_2.se ));
 sg13g2_dfrbp_1 \grid.cell_17_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1283),
    .D(_00345_),
    .Q_N(_00080_),
    .Q(\grid.cell_16_3.se ));
 sg13g2_dfrbp_1 \grid.cell_17_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1284),
    .D(_00346_),
    .Q_N(_00112_),
    .Q(\grid.cell_16_4.se ));
 sg13g2_dfrbp_1 \grid.cell_17_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1285),
    .D(_00347_),
    .Q_N(_00144_),
    .Q(\grid.cell_16_5.se ));
 sg13g2_dfrbp_1 \grid.cell_17_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1286),
    .D(_00348_),
    .Q_N(_00176_),
    .Q(\grid.cell_16_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_18_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1287),
    .D(_00349_),
    .Q_N(_00223_),
    .Q(\grid.cell_17_0.s ));
 sg13g2_dfrbp_1 \grid.cell_18_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1288),
    .D(_00350_),
    .Q_N(_00222_),
    .Q(\grid.cell_17_0.se ));
 sg13g2_dfrbp_1 \grid.cell_18_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1289),
    .D(_00351_),
    .Q_N(_00221_),
    .Q(\grid.cell_17_1.se ));
 sg13g2_dfrbp_1 \grid.cell_18_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1290),
    .D(_00352_),
    .Q_N(_00051_),
    .Q(\grid.cell_17_2.se ));
 sg13g2_dfrbp_1 \grid.cell_18_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1291),
    .D(_00353_),
    .Q_N(_00083_),
    .Q(\grid.cell_17_3.se ));
 sg13g2_dfrbp_1 \grid.cell_18_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1292),
    .D(_00354_),
    .Q_N(_00115_),
    .Q(\grid.cell_17_4.se ));
 sg13g2_dfrbp_1 \grid.cell_18_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1293),
    .D(_00355_),
    .Q_N(_00147_),
    .Q(\grid.cell_17_5.se ));
 sg13g2_dfrbp_1 \grid.cell_18_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1294),
    .D(_00356_),
    .Q_N(_00179_),
    .Q(\grid.cell_17_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_19_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1295),
    .D(_00357_),
    .Q_N(_00220_),
    .Q(\grid.cell_18_0.s ));
 sg13g2_dfrbp_1 \grid.cell_19_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1296),
    .D(_00358_),
    .Q_N(_00211_),
    .Q(\grid.cell_18_0.se ));
 sg13g2_dfrbp_1 \grid.cell_19_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1297),
    .D(_00359_),
    .Q_N(_00210_),
    .Q(\grid.cell_18_1.se ));
 sg13g2_dfrbp_1 \grid.cell_19_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1298),
    .D(_00360_),
    .Q_N(_00050_),
    .Q(\grid.cell_18_2.se ));
 sg13g2_dfrbp_1 \grid.cell_19_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1299),
    .D(_00361_),
    .Q_N(_00082_),
    .Q(\grid.cell_18_3.se ));
 sg13g2_dfrbp_1 \grid.cell_19_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1300),
    .D(_00362_),
    .Q_N(_00114_),
    .Q(\grid.cell_18_4.se ));
 sg13g2_dfrbp_1 \grid.cell_19_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1301),
    .D(_00363_),
    .Q_N(_00146_),
    .Q(\grid.cell_18_5.se ));
 sg13g2_dfrbp_1 \grid.cell_19_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1302),
    .D(_00364_),
    .Q_N(_00178_),
    .Q(\grid.cell_18_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_1_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1303),
    .D(_00365_),
    .Q_N(_00212_),
    .Q(\grid.cell_0_0.s ));
 sg13g2_dfrbp_1 \grid.cell_1_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1304),
    .D(_00366_),
    .Q_N(_00217_),
    .Q(\grid.cell_0_0.se ));
 sg13g2_dfrbp_1 \grid.cell_1_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1305),
    .D(_00367_),
    .Q_N(_00214_),
    .Q(\grid.cell_0_1.se ));
 sg13g2_dfrbp_1 \grid.cell_1_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1306),
    .D(_00368_),
    .Q_N(_00032_),
    .Q(\grid.cell_0_2.se ));
 sg13g2_dfrbp_1 \grid.cell_1_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1307),
    .D(_00369_),
    .Q_N(_00064_),
    .Q(\grid.cell_0_3.se ));
 sg13g2_dfrbp_1 \grid.cell_1_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1308),
    .D(_00370_),
    .Q_N(_00096_),
    .Q(\grid.cell_0_4.se ));
 sg13g2_dfrbp_1 \grid.cell_1_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1309),
    .D(_00371_),
    .Q_N(_00128_),
    .Q(\grid.cell_0_5.se ));
 sg13g2_dfrbp_1 \grid.cell_1_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1310),
    .D(_00372_),
    .Q_N(_00160_),
    .Q(\grid.cell_0_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_20_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1311),
    .D(_00373_),
    .Q_N(_00209_),
    .Q(\grid.cell_19_0.s ));
 sg13g2_dfrbp_1 \grid.cell_20_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1312),
    .D(_00374_),
    .Q_N(_00208_),
    .Q(\grid.cell_19_0.se ));
 sg13g2_dfrbp_1 \grid.cell_20_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1313),
    .D(_00375_),
    .Q_N(_00207_),
    .Q(\grid.cell_19_1.se ));
 sg13g2_dfrbp_1 \grid.cell_20_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1314),
    .D(_00376_),
    .Q_N(_00053_),
    .Q(\grid.cell_19_2.se ));
 sg13g2_dfrbp_1 \grid.cell_20_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1315),
    .D(_00377_),
    .Q_N(_00085_),
    .Q(\grid.cell_19_3.se ));
 sg13g2_dfrbp_1 \grid.cell_20_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1316),
    .D(_00378_),
    .Q_N(_00117_),
    .Q(\grid.cell_19_4.se ));
 sg13g2_dfrbp_1 \grid.cell_20_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1317),
    .D(_00379_),
    .Q_N(_00149_),
    .Q(\grid.cell_19_5.se ));
 sg13g2_dfrbp_1 \grid.cell_20_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1318),
    .D(_00380_),
    .Q_N(_00181_),
    .Q(\grid.cell_19_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_21_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1319),
    .D(_00381_),
    .Q_N(_00206_),
    .Q(\grid.cell_20_0.s ));
 sg13g2_dfrbp_1 \grid.cell_21_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1320),
    .D(_00382_),
    .Q_N(_00205_),
    .Q(\grid.cell_20_0.se ));
 sg13g2_dfrbp_1 \grid.cell_21_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1321),
    .D(_00383_),
    .Q_N(_00204_),
    .Q(\grid.cell_20_1.se ));
 sg13g2_dfrbp_1 \grid.cell_21_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1322),
    .D(_00384_),
    .Q_N(_00052_),
    .Q(\grid.cell_20_2.se ));
 sg13g2_dfrbp_1 \grid.cell_21_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1323),
    .D(_00385_),
    .Q_N(_00084_),
    .Q(\grid.cell_20_3.se ));
 sg13g2_dfrbp_1 \grid.cell_21_5.state$_SDFFE_PP0P_  (.CLK(clknet_4_3__leaf_clk),
    .RESET_B(net1324),
    .D(_00386_),
    .Q_N(_00116_),
    .Q(\grid.cell_20_4.se ));
 sg13g2_dfrbp_1 \grid.cell_21_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1325),
    .D(_00387_),
    .Q_N(_00148_),
    .Q(\grid.cell_20_5.se ));
 sg13g2_dfrbp_1 \grid.cell_21_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1326),
    .D(_00388_),
    .Q_N(_00180_),
    .Q(\grid.cell_20_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_22_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1327),
    .D(_00389_),
    .Q_N(_00203_),
    .Q(\grid.cell_21_0.s ));
 sg13g2_dfrbp_1 \grid.cell_22_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1328),
    .D(_00390_),
    .Q_N(_00202_),
    .Q(\grid.cell_21_0.se ));
 sg13g2_dfrbp_1 \grid.cell_22_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1329),
    .D(_00391_),
    .Q_N(_00201_),
    .Q(\grid.cell_21_1.se ));
 sg13g2_dfrbp_1 \grid.cell_22_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1330),
    .D(_00392_),
    .Q_N(_00055_),
    .Q(\grid.cell_21_2.se ));
 sg13g2_dfrbp_1 \grid.cell_22_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1331),
    .D(_00393_),
    .Q_N(_00087_),
    .Q(\grid.cell_21_3.se ));
 sg13g2_dfrbp_1 \grid.cell_22_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1332),
    .D(_00394_),
    .Q_N(_00119_),
    .Q(\grid.cell_21_4.se ));
 sg13g2_dfrbp_1 \grid.cell_22_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1333),
    .D(_00395_),
    .Q_N(_00151_),
    .Q(\grid.cell_21_5.se ));
 sg13g2_dfrbp_1 \grid.cell_22_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1334),
    .D(_00396_),
    .Q_N(_00183_),
    .Q(\grid.cell_21_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_23_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1335),
    .D(_00397_),
    .Q_N(_00200_),
    .Q(\grid.cell_22_0.s ));
 sg13g2_dfrbp_1 \grid.cell_23_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1336),
    .D(_00398_),
    .Q_N(_00197_),
    .Q(\grid.cell_22_0.se ));
 sg13g2_dfrbp_1 \grid.cell_23_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1337),
    .D(_00399_),
    .Q_N(_00194_),
    .Q(\grid.cell_22_1.se ));
 sg13g2_dfrbp_1 \grid.cell_23_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1338),
    .D(_00400_),
    .Q_N(_00054_),
    .Q(\grid.cell_22_2.se ));
 sg13g2_dfrbp_1 \grid.cell_23_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1339),
    .D(_00401_),
    .Q_N(_00086_),
    .Q(\grid.cell_22_3.se ));
 sg13g2_dfrbp_1 \grid.cell_23_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1340),
    .D(_00402_),
    .Q_N(_00118_),
    .Q(\grid.cell_22_4.se ));
 sg13g2_dfrbp_1 \grid.cell_23_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1341),
    .D(_00403_),
    .Q_N(_00150_),
    .Q(\grid.cell_22_5.se ));
 sg13g2_dfrbp_1 \grid.cell_23_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1342),
    .D(_00404_),
    .Q_N(_00182_),
    .Q(\grid.cell_22_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_24_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1343),
    .D(_00405_),
    .Q_N(_00198_),
    .Q(\grid.cell_23_0.s ));
 sg13g2_dfrbp_1 \grid.cell_24_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1344),
    .D(_00406_),
    .Q_N(_00195_),
    .Q(\grid.cell_23_0.se ));
 sg13g2_dfrbp_1 \grid.cell_24_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1345),
    .D(_00407_),
    .Q_N(_00192_),
    .Q(\grid.cell_23_1.se ));
 sg13g2_dfrbp_1 \grid.cell_24_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1346),
    .D(_00408_),
    .Q_N(_00056_),
    .Q(\grid.cell_23_2.se ));
 sg13g2_dfrbp_1 \grid.cell_24_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1347),
    .D(_00409_),
    .Q_N(_00088_),
    .Q(\grid.cell_23_3.se ));
 sg13g2_dfrbp_1 \grid.cell_24_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1348),
    .D(_00410_),
    .Q_N(_00120_),
    .Q(\grid.cell_23_4.se ));
 sg13g2_dfrbp_1 \grid.cell_24_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1349),
    .D(_00411_),
    .Q_N(_00152_),
    .Q(\grid.cell_23_5.se ));
 sg13g2_dfrbp_1 \grid.cell_24_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1350),
    .D(_00412_),
    .Q_N(_00185_),
    .Q(\grid.cell_23_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_25_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1351),
    .D(_00413_),
    .Q_N(_00199_),
    .Q(\grid.cell_24_0.s ));
 sg13g2_dfrbp_1 \grid.cell_25_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1352),
    .D(_00414_),
    .Q_N(_00196_),
    .Q(\grid.cell_24_0.se ));
 sg13g2_dfrbp_1 \grid.cell_25_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1353),
    .D(_00415_),
    .Q_N(_00193_),
    .Q(\grid.cell_24_1.se ));
 sg13g2_dfrbp_1 \grid.cell_25_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1354),
    .D(_00416_),
    .Q_N(_00057_),
    .Q(\grid.cell_24_2.se ));
 sg13g2_dfrbp_1 \grid.cell_25_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1355),
    .D(_00417_),
    .Q_N(_00089_),
    .Q(\grid.cell_24_3.se ));
 sg13g2_dfrbp_1 \grid.cell_25_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1356),
    .D(_00418_),
    .Q_N(_00121_),
    .Q(\grid.cell_24_4.se ));
 sg13g2_dfrbp_1 \grid.cell_25_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1357),
    .D(_00419_),
    .Q_N(_00153_),
    .Q(\grid.cell_24_5.se ));
 sg13g2_dfrbp_1 \grid.cell_25_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1358),
    .D(_00420_),
    .Q_N(_00184_),
    .Q(\grid.cell_24_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_26_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1359),
    .D(_00421_),
    .Q_N(_00016_),
    .Q(\grid.cell_25_0.s ));
 sg13g2_dfrbp_1 \grid.cell_26_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1360),
    .D(_00422_),
    .Q_N(_00015_),
    .Q(\grid.cell_25_0.se ));
 sg13g2_dfrbp_1 \grid.cell_26_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1361),
    .D(_00423_),
    .Q_N(_00014_),
    .Q(\grid.cell_25_1.se ));
 sg13g2_dfrbp_1 \grid.cell_26_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1362),
    .D(_00424_),
    .Q_N(_00059_),
    .Q(\grid.cell_25_2.se ));
 sg13g2_dfrbp_1 \grid.cell_26_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1363),
    .D(_00425_),
    .Q_N(_00091_),
    .Q(\grid.cell_25_3.se ));
 sg13g2_dfrbp_1 \grid.cell_26_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1364),
    .D(_00426_),
    .Q_N(_00123_),
    .Q(\grid.cell_25_4.se ));
 sg13g2_dfrbp_1 \grid.cell_26_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1365),
    .D(_00427_),
    .Q_N(_00155_),
    .Q(\grid.cell_25_5.se ));
 sg13g2_dfrbp_1 \grid.cell_26_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1366),
    .D(_00428_),
    .Q_N(_00187_),
    .Q(\grid.cell_25_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_27_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1367),
    .D(_00429_),
    .Q_N(_00013_),
    .Q(\grid.cell_26_0.s ));
 sg13g2_dfrbp_1 \grid.cell_27_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1368),
    .D(_00430_),
    .Q_N(_00012_),
    .Q(\grid.cell_26_0.se ));
 sg13g2_dfrbp_1 \grid.cell_27_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1369),
    .D(_00431_),
    .Q_N(_00011_),
    .Q(\grid.cell_26_1.se ));
 sg13g2_dfrbp_1 \grid.cell_27_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1370),
    .D(_00432_),
    .Q_N(_00058_),
    .Q(\grid.cell_26_2.se ));
 sg13g2_dfrbp_1 \grid.cell_27_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1371),
    .D(_00433_),
    .Q_N(_00090_),
    .Q(\grid.cell_26_3.se ));
 sg13g2_dfrbp_1 \grid.cell_27_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1372),
    .D(_00434_),
    .Q_N(_00122_),
    .Q(\grid.cell_26_4.se ));
 sg13g2_dfrbp_1 \grid.cell_27_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1373),
    .D(_00435_),
    .Q_N(_00154_),
    .Q(\grid.cell_26_5.se ));
 sg13g2_dfrbp_1 \grid.cell_27_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1374),
    .D(_00436_),
    .Q_N(_00186_),
    .Q(\grid.cell_26_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_28_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1375),
    .D(_00437_),
    .Q_N(_00010_),
    .Q(\grid.cell_27_0.s ));
 sg13g2_dfrbp_1 \grid.cell_28_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1376),
    .D(_00438_),
    .Q_N(_00009_),
    .Q(\grid.cell_27_0.se ));
 sg13g2_dfrbp_1 \grid.cell_28_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1377),
    .D(_00439_),
    .Q_N(_00008_),
    .Q(\grid.cell_27_1.se ));
 sg13g2_dfrbp_1 \grid.cell_28_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1378),
    .D(_00440_),
    .Q_N(_00061_),
    .Q(\grid.cell_27_2.se ));
 sg13g2_dfrbp_1 \grid.cell_28_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1379),
    .D(_00441_),
    .Q_N(_00093_),
    .Q(\grid.cell_27_3.se ));
 sg13g2_dfrbp_1 \grid.cell_28_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1380),
    .D(_00442_),
    .Q_N(_00125_),
    .Q(\grid.cell_27_4.se ));
 sg13g2_dfrbp_1 \grid.cell_28_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1381),
    .D(_00443_),
    .Q_N(_00157_),
    .Q(\grid.cell_27_5.se ));
 sg13g2_dfrbp_1 \grid.cell_28_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1382),
    .D(_00444_),
    .Q_N(_00189_),
    .Q(\grid.cell_27_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_29_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1383),
    .D(_00445_),
    .Q_N(_00007_),
    .Q(\grid.cell_28_0.s ));
 sg13g2_dfrbp_1 \grid.cell_29_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1384),
    .D(_00446_),
    .Q_N(_00006_),
    .Q(\grid.cell_28_0.se ));
 sg13g2_dfrbp_1 \grid.cell_29_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1385),
    .D(_00447_),
    .Q_N(_00005_),
    .Q(\grid.cell_28_1.se ));
 sg13g2_dfrbp_1 \grid.cell_29_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1386),
    .D(_00448_),
    .Q_N(_00060_),
    .Q(\grid.cell_28_2.se ));
 sg13g2_dfrbp_1 \grid.cell_29_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1387),
    .D(_00449_),
    .Q_N(_00092_),
    .Q(\grid.cell_28_3.se ));
 sg13g2_dfrbp_1 \grid.cell_29_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1388),
    .D(_00450_),
    .Q_N(_00124_),
    .Q(\grid.cell_28_4.se ));
 sg13g2_dfrbp_1 \grid.cell_29_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1389),
    .D(_00451_),
    .Q_N(_00156_),
    .Q(\grid.cell_28_5.se ));
 sg13g2_dfrbp_1 \grid.cell_29_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1390),
    .D(_00452_),
    .Q_N(_00188_),
    .Q(\grid.cell_28_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_2_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1391),
    .D(_00453_),
    .Q_N(_00213_),
    .Q(\grid.cell_1_0.s ));
 sg13g2_dfrbp_1 \grid.cell_2_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1392),
    .D(_00454_),
    .Q_N(_00218_),
    .Q(\grid.cell_1_0.se ));
 sg13g2_dfrbp_1 \grid.cell_2_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1393),
    .D(_00455_),
    .Q_N(_00215_),
    .Q(\grid.cell_1_1.se ));
 sg13g2_dfrbp_1 \grid.cell_2_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1394),
    .D(_00456_),
    .Q_N(_00035_),
    .Q(\grid.cell_1_2.se ));
 sg13g2_dfrbp_1 \grid.cell_2_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1395),
    .D(_00457_),
    .Q_N(_00067_),
    .Q(\grid.cell_1_3.se ));
 sg13g2_dfrbp_1 \grid.cell_2_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1396),
    .D(_00458_),
    .Q_N(_00099_),
    .Q(\grid.cell_1_4.se ));
 sg13g2_dfrbp_1 \grid.cell_2_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1397),
    .D(_00459_),
    .Q_N(_00131_),
    .Q(\grid.cell_1_5.se ));
 sg13g2_dfrbp_1 \grid.cell_2_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1398),
    .D(_00460_),
    .Q_N(_00163_),
    .Q(\grid.cell_1_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_30_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1399),
    .D(_00461_),
    .Q_N(_00272_),
    .Q(\grid.cell_29_0.s ));
 sg13g2_dfrbp_1 \grid.cell_30_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1400),
    .D(_00462_),
    .Q_N(_00274_),
    .Q(\grid.cell_29_0.se ));
 sg13g2_dfrbp_1 \grid.cell_30_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1401),
    .D(_00463_),
    .Q_N(_00273_),
    .Q(\grid.cell_29_1.se ));
 sg13g2_dfrbp_1 \grid.cell_30_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1402),
    .D(_00464_),
    .Q_N(_00063_),
    .Q(\grid.cell_29_2.se ));
 sg13g2_dfrbp_1 \grid.cell_30_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1403),
    .D(_00465_),
    .Q_N(_00095_),
    .Q(\grid.cell_29_3.se ));
 sg13g2_dfrbp_1 \grid.cell_30_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1404),
    .D(_00466_),
    .Q_N(_00127_),
    .Q(\grid.cell_29_4.se ));
 sg13g2_dfrbp_1 \grid.cell_30_6.state$_SDFFE_PP0P_  (.CLK(clknet_4_6__leaf_clk),
    .RESET_B(net1405),
    .D(_00467_),
    .Q_N(_00159_),
    .Q(\grid.cell_29_5.se ));
 sg13g2_dfrbp_1 \grid.cell_30_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1406),
    .D(_00468_),
    .Q_N(_00191_),
    .Q(\grid.cell_29_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_31_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1407),
    .D(_00469_),
    .Q_N(_00250_),
    .Q(\grid.cell_0_0.n ));
 sg13g2_dfrbp_1 \grid.cell_31_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1408),
    .D(_00470_),
    .Q_N(_00252_),
    .Q(\grid.cell_0_0.ne ));
 sg13g2_dfrbp_1 \grid.cell_31_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1409),
    .D(_00471_),
    .Q_N(_00251_),
    .Q(\grid.cell_0_1.ne ));
 sg13g2_dfrbp_1 \grid.cell_31_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1410),
    .D(_00472_),
    .Q_N(_00062_),
    .Q(\grid.cell_0_2.ne ));
 sg13g2_dfrbp_1 \grid.cell_31_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1411),
    .D(_00473_),
    .Q_N(_00094_),
    .Q(\grid.cell_0_3.ne ));
 sg13g2_dfrbp_1 \grid.cell_31_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1412),
    .D(_00474_),
    .Q_N(_00126_),
    .Q(\grid.cell_0_4.ne ));
 sg13g2_dfrbp_1 \grid.cell_31_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1413),
    .D(_00475_),
    .Q_N(_00158_),
    .Q(\grid.cell_0_5.ne ));
 sg13g2_dfrbp_1 \grid.cell_31_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1414),
    .D(_00476_),
    .Q_N(_00190_),
    .Q(\grid.cell_0_0.nw ));
 sg13g2_dfrbp_1 \grid.cell_3_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1415),
    .D(_00477_),
    .Q_N(_00271_),
    .Q(\grid.cell_2_0.s ));
 sg13g2_dfrbp_1 \grid.cell_3_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1416),
    .D(_00478_),
    .Q_N(_00270_),
    .Q(\grid.cell_2_0.se ));
 sg13g2_dfrbp_1 \grid.cell_3_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1417),
    .D(_00479_),
    .Q_N(_00269_),
    .Q(\grid.cell_2_1.se ));
 sg13g2_dfrbp_1 \grid.cell_3_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1418),
    .D(_00480_),
    .Q_N(_00034_),
    .Q(\grid.cell_2_2.se ));
 sg13g2_dfrbp_1 \grid.cell_3_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1419),
    .D(_00481_),
    .Q_N(_00066_),
    .Q(\grid.cell_2_3.se ));
 sg13g2_dfrbp_1 \grid.cell_3_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1420),
    .D(_00482_),
    .Q_N(_00098_),
    .Q(\grid.cell_2_4.se ));
 sg13g2_dfrbp_1 \grid.cell_3_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1421),
    .D(_00483_),
    .Q_N(_00130_),
    .Q(\grid.cell_2_5.se ));
 sg13g2_dfrbp_1 \grid.cell_3_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1422),
    .D(_00484_),
    .Q_N(_00162_),
    .Q(\grid.cell_2_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_4_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1423),
    .D(_00485_),
    .Q_N(_00268_),
    .Q(\grid.cell_3_0.s ));
 sg13g2_dfrbp_1 \grid.cell_4_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1424),
    .D(_00486_),
    .Q_N(_00267_),
    .Q(\grid.cell_3_0.se ));
 sg13g2_dfrbp_1 \grid.cell_4_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1425),
    .D(_00487_),
    .Q_N(_00266_),
    .Q(\grid.cell_3_1.se ));
 sg13g2_dfrbp_1 \grid.cell_4_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1426),
    .D(_00488_),
    .Q_N(_00037_),
    .Q(\grid.cell_3_2.se ));
 sg13g2_dfrbp_1 \grid.cell_4_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1427),
    .D(_00489_),
    .Q_N(_00069_),
    .Q(\grid.cell_3_3.se ));
 sg13g2_dfrbp_1 \grid.cell_4_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1428),
    .D(_00490_),
    .Q_N(_00101_),
    .Q(\grid.cell_3_4.se ));
 sg13g2_dfrbp_1 \grid.cell_4_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1429),
    .D(_00491_),
    .Q_N(_00133_),
    .Q(\grid.cell_3_5.se ));
 sg13g2_dfrbp_1 \grid.cell_4_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1430),
    .D(_00492_),
    .Q_N(_00165_),
    .Q(\grid.cell_3_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_5_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1431),
    .D(_00493_),
    .Q_N(_00265_),
    .Q(\grid.cell_4_0.s ));
 sg13g2_dfrbp_1 \grid.cell_5_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1432),
    .D(_00494_),
    .Q_N(_00264_),
    .Q(\grid.cell_4_0.se ));
 sg13g2_dfrbp_1 \grid.cell_5_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1433),
    .D(_00495_),
    .Q_N(_00263_),
    .Q(\grid.cell_4_1.se ));
 sg13g2_dfrbp_1 \grid.cell_5_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1434),
    .D(_00496_),
    .Q_N(_00036_),
    .Q(\grid.cell_4_2.se ));
 sg13g2_dfrbp_1 \grid.cell_5_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1435),
    .D(_00497_),
    .Q_N(_00068_),
    .Q(\grid.cell_4_3.se ));
 sg13g2_dfrbp_1 \grid.cell_5_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1436),
    .D(_00498_),
    .Q_N(_00100_),
    .Q(\grid.cell_4_4.se ));
 sg13g2_dfrbp_1 \grid.cell_5_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1437),
    .D(_00499_),
    .Q_N(_00132_),
    .Q(\grid.cell_4_5.se ));
 sg13g2_dfrbp_1 \grid.cell_5_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1438),
    .D(_00500_),
    .Q_N(_00164_),
    .Q(\grid.cell_4_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_6_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1439),
    .D(_00501_),
    .Q_N(_00262_),
    .Q(\grid.cell_5_0.s ));
 sg13g2_dfrbp_1 \grid.cell_6_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1440),
    .D(_00502_),
    .Q_N(_00261_),
    .Q(\grid.cell_5_0.se ));
 sg13g2_dfrbp_1 \grid.cell_6_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1441),
    .D(_00503_),
    .Q_N(_00260_),
    .Q(\grid.cell_5_1.se ));
 sg13g2_dfrbp_1 \grid.cell_6_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1442),
    .D(_00504_),
    .Q_N(_00039_),
    .Q(\grid.cell_5_2.se ));
 sg13g2_dfrbp_1 \grid.cell_6_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1443),
    .D(_00505_),
    .Q_N(_00071_),
    .Q(\grid.cell_5_3.se ));
 sg13g2_dfrbp_1 \grid.cell_6_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1444),
    .D(_00506_),
    .Q_N(_00103_),
    .Q(\grid.cell_5_4.se ));
 sg13g2_dfrbp_1 \grid.cell_6_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1445),
    .D(_00507_),
    .Q_N(_00135_),
    .Q(\grid.cell_5_5.se ));
 sg13g2_dfrbp_1 \grid.cell_6_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1446),
    .D(_00508_),
    .Q_N(_00167_),
    .Q(\grid.cell_5_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_7_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1447),
    .D(_00509_),
    .Q_N(_00259_),
    .Q(\grid.cell_6_0.s ));
 sg13g2_dfrbp_1 \grid.cell_7_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1448),
    .D(_00510_),
    .Q_N(_00258_),
    .Q(\grid.cell_6_0.se ));
 sg13g2_dfrbp_1 \grid.cell_7_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1449),
    .D(_00511_),
    .Q_N(_00257_),
    .Q(\grid.cell_6_1.se ));
 sg13g2_dfrbp_1 \grid.cell_7_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1450),
    .D(_00512_),
    .Q_N(_00038_),
    .Q(\grid.cell_6_2.se ));
 sg13g2_dfrbp_1 \grid.cell_7_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1451),
    .D(_00513_),
    .Q_N(_00070_),
    .Q(\grid.cell_6_3.se ));
 sg13g2_dfrbp_1 \grid.cell_7_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1452),
    .D(_00514_),
    .Q_N(_00102_),
    .Q(\grid.cell_6_4.se ));
 sg13g2_dfrbp_1 \grid.cell_7_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1453),
    .D(_00515_),
    .Q_N(_00134_),
    .Q(\grid.cell_6_5.se ));
 sg13g2_dfrbp_1 \grid.cell_7_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1454),
    .D(_00516_),
    .Q_N(_00166_),
    .Q(\grid.cell_6_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_8_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1455),
    .D(_00517_),
    .Q_N(_00254_),
    .Q(\grid.cell_7_0.s ));
 sg13g2_dfrbp_1 \grid.cell_8_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1456),
    .D(_00518_),
    .Q_N(_00256_),
    .Q(\grid.cell_7_0.se ));
 sg13g2_dfrbp_1 \grid.cell_8_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1457),
    .D(_00519_),
    .Q_N(_00255_),
    .Q(\grid.cell_7_1.se ));
 sg13g2_dfrbp_1 \grid.cell_8_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1458),
    .D(_00520_),
    .Q_N(_00041_),
    .Q(\grid.cell_7_2.se ));
 sg13g2_dfrbp_1 \grid.cell_8_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1459),
    .D(_00521_),
    .Q_N(_00073_),
    .Q(\grid.cell_7_3.se ));
 sg13g2_dfrbp_1 \grid.cell_8_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1460),
    .D(_00522_),
    .Q_N(_00105_),
    .Q(\grid.cell_7_4.se ));
 sg13g2_dfrbp_1 \grid.cell_8_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1461),
    .D(_00523_),
    .Q_N(_00137_),
    .Q(\grid.cell_7_5.se ));
 sg13g2_dfrbp_1 \grid.cell_8_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1462),
    .D(_00524_),
    .Q_N(_00169_),
    .Q(\grid.cell_7_0.sw ));
 sg13g2_dfrbp_1 \grid.cell_9_0.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1463),
    .D(_00525_),
    .Q_N(_00247_),
    .Q(\grid.cell_10_0.n ));
 sg13g2_dfrbp_1 \grid.cell_9_1.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1464),
    .D(_00526_),
    .Q_N(_00249_),
    .Q(\grid.cell_10_0.ne ));
 sg13g2_dfrbp_1 \grid.cell_9_2.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1465),
    .D(_00527_),
    .Q_N(_00248_),
    .Q(\grid.cell_10_1.ne ));
 sg13g2_dfrbp_1 \grid.cell_9_3.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1466),
    .D(_00528_),
    .Q_N(_00040_),
    .Q(\grid.cell_10_2.ne ));
 sg13g2_dfrbp_1 \grid.cell_9_4.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1467),
    .D(_00529_),
    .Q_N(_00072_),
    .Q(\grid.cell_10_3.ne ));
 sg13g2_dfrbp_1 \grid.cell_9_5.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1468),
    .D(_00530_),
    .Q_N(_00104_),
    .Q(\grid.cell_10_4.ne ));
 sg13g2_dfrbp_1 \grid.cell_9_6.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1469),
    .D(_00531_),
    .Q_N(_00136_),
    .Q(\grid.cell_10_5.ne ));
 sg13g2_dfrbp_1 \grid.cell_9_7.state$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1470),
    .D(_00532_),
    .Q_N(_00168_),
    .Q(\grid.cell_10_0.nw ));
 sg13g2_dfrbp_1 \max7219.col_index[0]$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1471),
    .D(_00533_),
    .Q_N(_00253_),
    .Q(\grid.row_select2[0] ));
 sg13g2_dfrbp_1 \max7219.col_index[1]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1472),
    .D(_00534_),
    .Q_N(_13369_),
    .Q(\grid.row_select2[1] ));
 sg13g2_dfrbp_1 \max7219.col_index[2]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1473),
    .D(_00535_),
    .Q_N(_00026_),
    .Q(\grid.row_select2[2] ));
 sg13g2_dfrbp_1 \max7219.init_index[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1474),
    .D(_00536_),
    .Q_N(_13368_),
    .Q(\max7219.init_index[0] ));
 sg13g2_dfrbp_1 \max7219.init_index[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1475),
    .D(_00537_),
    .Q_N(_13367_),
    .Q(\max7219.init_index[1] ));
 sg13g2_dfrbp_1 \max7219.load_row$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1476),
    .D(_00538_),
    .Q_N(_13366_),
    .Q(\max7219.load_row ));
 sg13g2_dfrbp_1 \max7219.matrix_index[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1477),
    .D(_00539_),
    .Q_N(_13365_),
    .Q(\grid.row_select2[3] ));
 sg13g2_dfrbp_1 \max7219.matrix_index[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1478),
    .D(_00540_),
    .Q_N(_13364_),
    .Q(\grid.row_select2[4] ));
 sg13g2_dfrbp_1 \max7219.max7219_enabled$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1479),
    .D(_00541_),
    .Q_N(_13363_),
    .Q(\max7219.max7219_enabled ));
 sg13g2_dfrbp_1 \max7219.max7219_row[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1480),
    .D(_00542_),
    .Q_N(_00031_),
    .Q(\max7219.max7219_row[0] ));
 sg13g2_dfrbp_1 \max7219.max7219_row[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1481),
    .D(_00543_),
    .Q_N(_13362_),
    .Q(\max7219.max7219_row[1] ));
 sg13g2_dfrbp_1 \max7219.max7219_row[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1482),
    .D(_00544_),
    .Q_N(_00027_),
    .Q(\max7219.max7219_row[2] ));
 sg13g2_dfrbp_1 \max7219.o_cs$_SDFFE_PN1P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1483),
    .D(_00545_),
    .Q_N(_00025_),
    .Q(\max7219.o_cs ));
 sg13g2_dfrbp_1 \max7219.row_data[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1484),
    .D(_00546_),
    .Q_N(_13361_),
    .Q(\max7219.row_data[0] ));
 sg13g2_dfrbp_1 \max7219.row_data[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1485),
    .D(_00547_),
    .Q_N(_13360_),
    .Q(\max7219.row_data[1] ));
 sg13g2_dfrbp_1 \max7219.row_data[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1486),
    .D(_00548_),
    .Q_N(_13359_),
    .Q(\max7219.row_data[2] ));
 sg13g2_dfrbp_1 \max7219.row_data[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1487),
    .D(_00549_),
    .Q_N(_13358_),
    .Q(\max7219.row_data[3] ));
 sg13g2_dfrbp_1 \max7219.row_data[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1488),
    .D(_00550_),
    .Q_N(_13357_),
    .Q(\max7219.row_data[4] ));
 sg13g2_dfrbp_1 \max7219.row_data[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1489),
    .D(_00551_),
    .Q_N(_13356_),
    .Q(\max7219.row_data[5] ));
 sg13g2_dfrbp_1 \max7219.row_data[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1490),
    .D(_00552_),
    .Q_N(_13355_),
    .Q(\max7219.row_data[6] ));
 sg13g2_dfrbp_1 \max7219.row_data[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1491),
    .D(_00553_),
    .Q_N(_13354_),
    .Q(\max7219.row_data[7] ));
 sg13g2_dfrbp_1 \max7219.spi_start$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1492),
    .D(_00554_),
    .Q_N(_13353_),
    .Q(\max7219.spi_start ));
 sg13g2_dfrbp_1 \max7219.spim.bit_index[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1493),
    .D(_00555_),
    .Q_N(_13352_),
    .Q(\max7219.spim.bit_index[0] ));
 sg13g2_dfrbp_1 \max7219.spim.bit_index[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1494),
    .D(_00556_),
    .Q_N(_13351_),
    .Q(\max7219.spim.bit_index[1] ));
 sg13g2_dfrbp_1 \max7219.spim.bit_index[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1495),
    .D(_00557_),
    .Q_N(_00029_),
    .Q(\max7219.spim.bit_index[2] ));
 sg13g2_dfrbp_1 \max7219.spim.bit_index[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1496),
    .D(_00558_),
    .Q_N(_13350_),
    .Q(\max7219.spim.bit_index[3] ));
 sg13g2_dfrbp_1 \max7219.spim.clk_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1497),
    .D(_00559_),
    .Q_N(_13349_),
    .Q(\max7219.spim.clk_count[0] ));
 sg13g2_dfrbp_1 \max7219.spim.clk_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1498),
    .D(_00560_),
    .Q_N(_13348_),
    .Q(\max7219.spim.clk_count[1] ));
 sg13g2_dfrbp_1 \max7219.spim.finish$_SDFFCE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1499),
    .D(_00561_),
    .Q_N(_00023_),
    .Q(\max7219.spim.finish ));
 sg13g2_dfrbp_1 \max7219.spim.o_busy$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1500),
    .D(_00562_),
    .Q_N(_00022_),
    .Q(\max7219.spi_busy ));
 sg13g2_dfrbp_1 \max7219.spim.o_mosi$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1501),
    .D(_00563_),
    .Q_N(_13347_),
    .Q(\max7219.o_mosi ));
 sg13g2_dfrbp_1 \max7219.spim.o_sck$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1502),
    .D(_00564_),
    .Q_N(_00004_),
    .Q(\max7219.o_sck ));
 sg13g2_dfrbp_1 \max7219.state[0]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1503),
    .D(_00000_),
    .Q_N(_00024_),
    .Q(\max7219.state[0] ));
 sg13g2_dfrbp_1 \max7219.state[1]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1504),
    .D(_00001_),
    .Q_N(_13373_),
    .Q(\max7219.state[1] ));
 sg13g2_dfrbp_1 \max7219.state[2]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1505),
    .D(_00002_),
    .Q_N(_00030_),
    .Q(\max7219.state[2] ));
 sg13g2_dfrbp_1 \max7219.state[3]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1506),
    .D(_00003_),
    .Q_N(_00028_),
    .Q(\max7219.state[3] ));
 sg13g2_dfrbp_1 \prev_rst_n$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1507),
    .D(net1),
    .Q_N(_13346_),
    .Q(prev_rst_n));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1508),
    .D(_00565_),
    .Q_N(_13345_),
    .Q(\silife_demo_inst.counter[0] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1509),
    .D(_00566_),
    .Q_N(_13344_),
    .Q(\silife_demo_inst.counter[10] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1510),
    .D(_00567_),
    .Q_N(_13343_),
    .Q(\silife_demo_inst.counter[11] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1511),
    .D(_00568_),
    .Q_N(_13342_),
    .Q(\silife_demo_inst.counter[12] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1512),
    .D(_00569_),
    .Q_N(_13341_),
    .Q(\silife_demo_inst.counter[13] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1513),
    .D(_00570_),
    .Q_N(_13340_),
    .Q(\silife_demo_inst.counter[14] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1514),
    .D(_00571_),
    .Q_N(_13339_),
    .Q(\silife_demo_inst.counter[15] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1515),
    .D(_00572_),
    .Q_N(_13338_),
    .Q(\silife_demo_inst.counter[16] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1516),
    .D(_00573_),
    .Q_N(_13337_),
    .Q(\silife_demo_inst.counter[17] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1517),
    .D(_00574_),
    .Q_N(_13336_),
    .Q(\silife_demo_inst.counter[18] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1518),
    .D(_00575_),
    .Q_N(_13335_),
    .Q(\silife_demo_inst.counter[19] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1519),
    .D(_00576_),
    .Q_N(_13334_),
    .Q(\silife_demo_inst.counter[1] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1520),
    .D(_00577_),
    .Q_N(_13333_),
    .Q(\silife_demo_inst.counter[20] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1521),
    .D(_00578_),
    .Q_N(_13332_),
    .Q(\silife_demo_inst.counter[21] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1522),
    .D(_00579_),
    .Q_N(_13331_),
    .Q(\silife_demo_inst.counter[22] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1523),
    .D(_00580_),
    .Q_N(_13330_),
    .Q(\silife_demo_inst.counter[23] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1524),
    .D(_00581_),
    .Q_N(_13329_),
    .Q(\silife_demo_inst.counter[24] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1525),
    .D(_00582_),
    .Q_N(_13328_),
    .Q(\silife_demo_inst.counter[25] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1526),
    .D(_00583_),
    .Q_N(_13327_),
    .Q(\silife_demo_inst.counter[26] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1527),
    .D(_00584_),
    .Q_N(_13326_),
    .Q(\silife_demo_inst.counter[27] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1528),
    .D(_00585_),
    .Q_N(_13325_),
    .Q(\silife_demo_inst.counter[28] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1529),
    .D(_00586_),
    .Q_N(_13324_),
    .Q(\silife_demo_inst.counter[29] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1530),
    .D(_00587_),
    .Q_N(_13323_),
    .Q(\silife_demo_inst.counter[2] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1531),
    .D(_00588_),
    .Q_N(_13322_),
    .Q(\silife_demo_inst.counter[30] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1532),
    .D(_00589_),
    .Q_N(_13321_),
    .Q(\silife_demo_inst.counter[31] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1533),
    .D(_00590_),
    .Q_N(_13320_),
    .Q(\silife_demo_inst.counter[3] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1534),
    .D(_00591_),
    .Q_N(_13319_),
    .Q(\silife_demo_inst.counter[4] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1535),
    .D(_00592_),
    .Q_N(_13318_),
    .Q(\silife_demo_inst.counter[5] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1536),
    .D(_00593_),
    .Q_N(_13317_),
    .Q(\silife_demo_inst.counter[6] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1537),
    .D(_00594_),
    .Q_N(_13316_),
    .Q(\silife_demo_inst.counter[7] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1538),
    .D(_00595_),
    .Q_N(_13315_),
    .Q(\silife_demo_inst.counter[8] ));
 sg13g2_dfrbp_1 \silife_demo_inst.counter[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1539),
    .D(_00596_),
    .Q_N(_13314_),
    .Q(\silife_demo_inst.counter[9] ));
 sg13g2_dfrbp_1 \silife_demo_inst.init_done$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1540),
    .D(_00597_),
    .Q_N(_13313_),
    .Q(\silife_demo_inst.init_done ));
 sg13g2_dfrbp_1 \silife_demo_inst.row_select[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1541),
    .D(_00598_),
    .Q_N(_00275_),
    .Q(\demo_row_select[0] ));
 sg13g2_dfrbp_1 \silife_demo_inst.row_select[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1542),
    .D(_00599_),
    .Q_N(_00020_),
    .Q(\demo_row_select[1] ));
 sg13g2_dfrbp_1 \silife_demo_inst.row_select[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1543),
    .D(_00600_),
    .Q_N(_00021_),
    .Q(\demo_row_select[2] ));
 sg13g2_dfrbp_1 \silife_demo_inst.row_select[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1544),
    .D(_00601_),
    .Q_N(_00019_),
    .Q(\demo_row_select[3] ));
 sg13g2_dfrbp_1 \silife_demo_inst.row_select[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1545),
    .D(_00602_),
    .Q_N(_00017_),
    .Q(\demo_row_select[4] ));
 sg13g2_dfrbp_1 \silife_demo_inst.step$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1546),
    .D(_00603_),
    .Q_N(_13312_),
    .Q(demo_step));
 sg13g2_dfrbp_1 \silife_demo_inst.wr_en$_SDFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1547),
    .D(_00604_),
    .Q_N(_00018_),
    .Q(demo_wr_en));
 sg13g2_dfrbp_1 \wr_available$_SDFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1548),
    .D(_00605_),
    .Q_N(_13311_),
    .Q(wr_available));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[6]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[7]),
    .X(net15));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[0]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[1]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[2]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[3]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[4]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[5]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[6]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout24 (.A(_06814_),
    .X(net24));
 sg13g2_buf_4 fanout25 (.X(net25),
    .A(_07562_));
 sg13g2_buf_2 fanout26 (.A(_06249_),
    .X(net26));
 sg13g2_buf_4 fanout27 (.X(net27),
    .A(_04088_));
 sg13g2_buf_2 fanout28 (.A(_04509_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_12298_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_10243_),
    .X(net30));
 sg13g2_buf_4 fanout31 (.X(net31),
    .A(_06019_));
 sg13g2_buf_2 fanout32 (.A(_05863_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_05812_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_04942_),
    .X(net34));
 sg13g2_buf_4 fanout35 (.X(net35),
    .A(_04077_));
 sg13g2_buf_2 fanout36 (.A(_01550_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_12828_),
    .X(net37));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(_11113_));
 sg13g2_buf_2 fanout39 (.A(_10684_),
    .X(net39));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(_09235_));
 sg13g2_buf_2 fanout41 (.A(_08352_),
    .X(net41));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(_07276_));
 sg13g2_buf_2 fanout43 (.A(_06762_),
    .X(net43));
 sg13g2_buf_4 fanout44 (.X(net44),
    .A(_05757_));
 sg13g2_buf_4 fanout45 (.X(net45),
    .A(_05119_));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(_05003_));
 sg13g2_buf_2 fanout47 (.A(_04941_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_04914_),
    .X(net48));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(_03164_));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(_01817_));
 sg13g2_buf_2 fanout51 (.A(_03955_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_02757_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_13187_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12514_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12450_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_09918_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_09856_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_08821_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_07201_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_06476_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_06065_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_04683_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_04654_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_04623_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_11714_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_13104_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_11411_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_09402_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_08737_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_08586_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_07561_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_07199_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_07117_),
    .X(net73));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(_06817_));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(_06538_));
 sg13g2_buf_4 fanout76 (.X(net76),
    .A(_06468_));
 sg13g2_buf_2 fanout77 (.A(_05897_),
    .X(net77));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(_05815_));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(_05737_));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_05678_));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(_05472_));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_05416_));
 sg13g2_buf_2 fanout83 (.A(_05268_),
    .X(net83));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(_04650_));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_02787_));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(_04801_));
 sg13g2_buf_8 fanout87 (.A(_04799_),
    .X(net87));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(_04796_));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(_04795_));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(_04788_));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(_04787_));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(_04784_));
 sg13g2_buf_8 fanout93 (.A(_04783_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_04749_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_03140_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_11608_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_10150_),
    .X(net97));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(_08549_));
 sg13g2_buf_2 fanout99 (.A(_07553_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_07194_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_06993_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_06897_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_06466_),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(_06425_));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(_06331_));
 sg13g2_buf_2 fanout106 (.A(_06285_),
    .X(net106));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(_06244_));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(_06114_));
 sg13g2_buf_2 fanout109 (.A(_06057_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_06055_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_05814_),
    .X(net111));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(_05739_));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(_05619_));
 sg13g2_buf_2 fanout114 (.A(_05517_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_05471_),
    .X(net115));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_05415_));
 sg13g2_buf_2 fanout117 (.A(_05408_),
    .X(net117));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(_05267_));
 sg13g2_buf_2 fanout119 (.A(_05136_),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(_05131_));
 sg13g2_buf_2 fanout121 (.A(_05129_),
    .X(net121));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(_04860_));
 sg13g2_buf_2 fanout123 (.A(_04642_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_04624_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_03831_),
    .X(net125));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_02820_));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_02776_));
 sg13g2_buf_2 fanout128 (.A(_04757_),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(_04739_),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(_04735_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_03813_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_03139_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_03091_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_01960_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_00875_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_12776_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_12459_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_11416_),
    .X(net138));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(_11407_));
 sg13g2_buf_2 fanout140 (.A(_11367_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_11116_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_10146_),
    .X(net142));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(_09916_));
 sg13g2_buf_2 fanout144 (.A(_09765_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_09083_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_08395_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_08299_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_08262_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_07887_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_07641_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_07505_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_07455_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_07211_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_07147_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_06844_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_06797_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_06179_),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(_06113_));
 sg13g2_buf_2 fanout159 (.A(_06063_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_05767_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_05710_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_05527_),
    .X(net162));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(_05130_));
 sg13g2_buf_2 fanout164 (.A(_05075_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_05057_),
    .X(net165));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(_04915_));
 sg13g2_buf_2 fanout167 (.A(_04859_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_04614_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_04109_),
    .X(net169));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(_03821_));
 sg13g2_buf_2 fanout171 (.A(_02809_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_02765_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_02647_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_02626_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_02615_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_02043_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_01913_),
    .X(net177));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(_04793_));
 sg13g2_buf_8 fanout179 (.A(_04792_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_04312_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_04266_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_04259_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_04247_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_03594_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_03460_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_03271_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_03208_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_03064_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_03063_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_02905_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_02782_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_02685_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_02680_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_02654_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_02563_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_02459_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_02303_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_02185_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_02152_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_01959_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_01865_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_01727_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_01602_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_01566_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_00778_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_13299_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_13244_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_13112_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_13111_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_12936_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_12890_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_12721_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_12678_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_12651_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_12567_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_12458_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_12423_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_12387_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_12286_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_12212_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_12154_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_12034_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_12013_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_11990_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_11886_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_11854_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_11795_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_11744_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_11741_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_11686_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_11490_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_11415_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_11364_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_11255_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_11161_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_11100_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_11085_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_11068_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_11048_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_10767_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_10658_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_10657_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_10534_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_10514_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_10496_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_10460_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_10401_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_10363_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_10307_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_10298_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_10257_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_10156_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_10116_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_10097_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_10083_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_09987_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_09976_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_09938_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_09799_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_09743_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_09717_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_09662_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_09634_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_09545_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_09542_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_09471_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_09381_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_09319_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_09309_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_09201_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_09197_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_09191_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_09185_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_09176_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_09041_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_08928_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_08927_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_08891_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_08768_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_08615_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_08607_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_08530_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_08507_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_08496_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_08402_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_08392_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_08373_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_08239_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_08234_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_08205_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_08195_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_08171_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_08124_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_08066_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_07993_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_07991_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_07886_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_07867_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_07836_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_07798_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_07673_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_07640_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_07624_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_07491_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_07480_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_07448_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_07396_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_07336_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_07210_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_06989_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_06905_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_06900_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_06888_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_06796_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_06729_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_06673_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_06667_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_06633_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_06542_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_06472_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_06457_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_06368_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_06323_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_06195_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_06178_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_06168_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_06112_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_05939_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_05904_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_05781_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_05764_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_05709_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_05698_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_05679_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_05646_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_05627_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_05626_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_05624_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_05568_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_05537_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_05526_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_05507_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_05502_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_05490_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_05426_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_05387_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_05367_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_05357_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_05319_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_05283_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_05250_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_05239_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_05216_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_05205_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_05194_),
    .X(net355));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(_05124_));
 sg13g2_buf_2 fanout357 (.A(_05105_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_05074_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_05073_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_05071_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_05064_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_05007_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_04800_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_04674_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_04545_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_04495_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_04099_),
    .X(net367));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(_03810_));
 sg13g2_buf_2 fanout369 (.A(_03756_),
    .X(net369));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(_02970_));
 sg13g2_buf_2 fanout371 (.A(_02679_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_02636_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_02572_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_02442_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_02032_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_01503_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_13053_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_12999_),
    .X(net378));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(_04395_));
 sg13g2_buf_8 fanout380 (.A(_04383_),
    .X(net380));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(_04367_));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(_04366_));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(_04364_));
 sg13g2_buf_2 fanout384 (.A(_04302_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_04300_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_04265_),
    .X(net386));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(_04258_));
 sg13g2_buf_8 fanout388 (.A(_04246_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_03459_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_03453_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_03447_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_03372_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_03324_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_03249_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_03232_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_03202_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_03187_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_03176_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_03018_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_02998_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_02956_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_02945_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_02915_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_02854_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_02810_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_02760_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_02653_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_02613_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_02573_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_02501_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_02441_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_02438_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_02407_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_02400_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_02389_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_02378_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_02267_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_02190_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_02159_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_02124_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_02070_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_02038_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_02010_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_01958_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_01954_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_01829_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_01812_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_01770_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_01750_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_01711_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_01685_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_01619_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_01600_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_01554_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_00977_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_00776_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_00736_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_00735_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_00717_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_00661_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_00647_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_00644_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_13298_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_13238_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_13195_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_13190_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_13108_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_13025_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_12962_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_12908_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_12849_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_12837_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_12834_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_12716_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_12661_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_12646_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_12616_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_12518_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_12469_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_12457_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_12454_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_12376_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_12318_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_12282_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_12264_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_12180_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_12118_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_12101_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_12099_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_12033_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_11989_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_11950_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_11885_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_11853_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_11851_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_11785_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_11729_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_11646_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_11629_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_11597_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_11593_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_11531_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_11489_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_11476_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_11414_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_11375_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_11363_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_11243_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_11218_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_11210_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_11180_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_11179_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_11067_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_11035_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_11019_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_11013_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_11000_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_10878_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_10872_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_10840_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_10831_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_10806_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_10785_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_10746_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_10716_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_10665_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_10656_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_10635_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_10615_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_10502_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_10487_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_10482_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_10439_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_10400_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_10392_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_10362_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_10311_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_10306_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_10267_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_10263_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_10256_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_10237_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_10200_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_10115_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_10096_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_10082_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_09986_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_09943_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_09889_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_09880_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_09872_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_09870_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_09818_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_09759_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_09742_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_09733_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_09698_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_09661_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_09642_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_09633_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_09602_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_09600_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_09544_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_09527_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_09412_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_09409_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_09373_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_09358_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_09313_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_09280_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_09239_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_09196_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_09184_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_09040_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_09035_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_08990_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_08965_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_08926_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_08892_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_08855_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_08843_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_08803_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_08763_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_08750_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_08741_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_08613_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_08606_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_08575_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_08506_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_08476_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_08442_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_08415_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_08378_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_08372_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_08231_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_08199_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_08164_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_08156_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_08123_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_08052_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_08047_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_08036_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_07990_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_07988_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_07869_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_07835_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_07797_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_07789_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_07744_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_07669_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_07632_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_07620_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_07484_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_07462_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_07447_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_07391_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_07381_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_07364_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_07362_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_07335_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_07334_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_07301_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_07244_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_07209_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_07205_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_07102_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_07092_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_07049_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_07044_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_07033_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_06965_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_06912_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_06904_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_06870_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_06859_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_06839_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_06815_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_06732_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_06728_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_06700_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_06672_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_06632_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_06597_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_06556_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_06548_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_06544_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_06507_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_06488_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_06383_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_06367_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_06362_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_06293_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_06282_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_06254_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_06194_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_06170_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_06118_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_06111_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_06077_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_06075_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_05957_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_05938_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_05903_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_05866_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_05849_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_05763_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_05700_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_05697_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_05634_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_05625_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_05536_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_05530_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_05525_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_05497_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_05492_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_05489_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_05451_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_05449_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_05444_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_05436_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_05411_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_05401_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_05386_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_05376_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_05366_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_05363_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_05360_),
    .X(net667));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(_05355_));
 sg13g2_buf_2 fanout669 (.A(_05306_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_05297_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_05294_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_05275_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_05241_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_05215_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_05210_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_05209_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_05204_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_05200_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_05199_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_05197_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_05193_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_05190_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_05121_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_05060_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_05051_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_05018_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_05014_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_05013_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_05010_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_05006_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_04958_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_04945_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_04885_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_04789_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_04768_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_04721_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_04283_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_04264_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_04217_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_04152_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_03682_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_03606_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_03541_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_03380_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_03369_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_02669_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_02593_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_02475_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_02432_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_02377_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_02162_),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_01676_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_01492_),
    .X(net713));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(_01064_));
 sg13g2_buf_2 fanout715 (.A(_00669_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_12988_),
    .X(net716));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(_04382_));
 sg13g2_buf_8 fanout718 (.A(_04362_),
    .X(net718));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(_04351_));
 sg13g2_buf_8 fanout720 (.A(_04349_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_04305_),
    .X(net721));
 sg13g2_buf_4 fanout722 (.X(net722),
    .A(_04299_));
 sg13g2_buf_2 fanout723 (.A(_04263_),
    .X(net723));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(_04253_));
 sg13g2_buf_4 fanout725 (.X(net725),
    .A(_04245_));
 sg13g2_buf_2 fanout726 (.A(_03437_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_03395_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_03361_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_03301_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_03262_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_03248_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_03201_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_03186_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_03184_),
    .X(net734));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(_03175_));
 sg13g2_buf_2 fanout736 (.A(_03017_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_02990_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_02951_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_02922_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_02889_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_02886_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_02832_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_02821_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_02780_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_02759_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_02644_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_02606_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_02564_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_02513_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_02492_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_02437_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_02429_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_02427_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_02379_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_02376_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_02274_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_02235_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_02178_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_02153_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_02109_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_02092_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_02035_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_02023_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_02018_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_01991_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_01957_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_01953_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_01822_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_01790_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_01769_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_01696_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_01679_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_01618_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_01596_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_01556_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_01553_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_01551_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_00753_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_00710_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_00665_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_00626_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_00614_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_13260_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_13217_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_13193_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_13189_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_13062_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(_13016_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_12993_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_12938_),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_12892_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_12884_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_12864_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_12833_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_12830_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_12700_),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(_12653_),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(_12618_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_12594_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_12570_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_12517_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_12492_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_12486_),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_12473_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_12456_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_12453_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_12451_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_12341_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_12309_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_12266_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_12252_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_12240_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_12179_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_12125_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_12100_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_12098_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_12003_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_11973_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_11918_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_11878_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_11857_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_11843_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_11784_),
    .X(net823));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(_11755_));
 sg13g2_buf_2 fanout825 (.A(_11737_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_11728_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_11715_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_11614_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_11576_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_11536_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_11522_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_11481_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_11472_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_11413_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_11362_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_11360_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_11351_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_11349_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_11242_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_11196_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_11159_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_11139_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_11129_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_11066_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_11060_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_11057_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_11002_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_10999_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_10875_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_10830_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_10784_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_10759_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_10738_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_10686_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_10650_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_10642_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_10634_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_10619_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_10572_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_10486_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_10431_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_10399_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_10365_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_10353_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_10305_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_10248_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_10246_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_10244_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_10165_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_10114_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_10078_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_10022_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_09991_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_09980_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_09936_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_09871_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_09869_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_09732_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_09697_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_09660_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_09632_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_09599_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_09580_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_09540_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_09539_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_09408_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_09371_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_09339_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_09303_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_09266_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_09238_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_09217_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_09186_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_09179_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_09174_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_09170_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_09038_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_09005_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_08989_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_08925_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_08908_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_08881_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_08824_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_08812_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_08775_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(_08767_),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_08749_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_08593_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_08555_),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_08505_),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(_08469_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_08426_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_08414_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_08371_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_08359_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_08355_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(_08230_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_08193_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_08151_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_08096_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_08045_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_08035_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_07989_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_07987_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_07856_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_07824_),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(_07787_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_07732_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_07718_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_07668_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_07653_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_07631_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_07615_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_07609_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_07483_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_07430_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_07390_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_07347_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_07333_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_07291_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_07269_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_07208_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_07204_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_07097_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_07091_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_07041_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_07014_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_06978_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_06972_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_06956_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_06914_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_06903_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_06857_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_06849_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_06841_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_06714_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_06671_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_06625_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_06596_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_06540_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_06533_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_06496_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_06495_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_06340_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_06292_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_06251_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_06200_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_06186_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_06122_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_06099_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_06096_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_06076_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_06074_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_05985_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_05937_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_05902_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_05883_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_05865_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_05836_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_05829_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_05760_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_05741_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_05704_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_05699_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_05693_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_05685_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_05644_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_05601_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_05535_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_05532_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_05529_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_05524_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_05493_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_05491_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_05476_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_05442_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_05438_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_05435_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_05365_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_05362_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_05359_),
    .X(net1001));
 sg13g2_buf_4 fanout1002 (.X(net1002),
    .A(_05354_));
 sg13g2_buf_2 fanout1003 (.A(_05311_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_05307_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_05305_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_05274_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_05233_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_05229_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_05227_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_05221_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_05219_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_05214_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_05203_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_05196_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_05192_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_05189_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_05173_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_05059_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_05017_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_05012_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_05009_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_05005_),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_04951_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_04948_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_04944_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_04884_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_04779_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_04758_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_04206_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_04174_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_04142_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_03895_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_03337_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_03326_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_03272_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_03229_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_02874_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_02658_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_02583_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_02464_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_02421_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_02366_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_02345_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_02302_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_02151_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_02130_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_02108_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_01742_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_01666_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_01612_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_01590_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_01525_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_01482_),
    .X(net1053));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(_01053_));
 sg13g2_buf_2 fanout1055 (.A(_00990_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_00788_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_00659_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_13202_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_13074_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_12977_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_04248_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_03830_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_03403_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_03391_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_03067_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_02985_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_02978_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_02939_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_02937_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_02831_),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_02819_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_02672_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(_02364_),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_02265_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_02107_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_01952_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_01878_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_01788_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_01782_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_01582_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_01552_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_00619_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(_13188_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_12981_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(_12883_),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_12759_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_12697_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(_12617_),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_12569_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_12455_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_12374_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_12334_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_12305_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_12229_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_12021_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_11916_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(_11833_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_11770_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_11725_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_11613_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_11584_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_11350_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_11195_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_11153_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_11117_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_10998_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_10651_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_10641_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_10533_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_10520_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_10447_),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_10252_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_10154_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_10131_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_10046_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_10021_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_09899_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_09857_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_09783_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(_09672_),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(_09620_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_09586_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_09407_),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(_09348_),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_09288_),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(_09237_),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(_09206_),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(_09081_),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_08966_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(_08907_),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_08671_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(_08648_),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_08600_),
    .X(net1133));
 sg13g2_buf_2 fanout1134 (.A(_08592_),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(_08563_),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(_08554_),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(_08421_),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(_08354_),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(_08270_),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(_08242_),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(_08132_),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(_08025_),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(_07981_),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(_07913_),
    .X(net1144));
 sg13g2_buf_2 fanout1145 (.A(_07894_),
    .X(net1145));
 sg13g2_buf_2 fanout1146 (.A(_07829_),
    .X(net1146));
 sg13g2_buf_2 fanout1147 (.A(_07815_),
    .X(net1147));
 sg13g2_buf_2 fanout1148 (.A(_07761_),
    .X(net1148));
 sg13g2_buf_2 fanout1149 (.A(_07759_),
    .X(net1149));
 sg13g2_buf_2 fanout1150 (.A(_07717_),
    .X(net1150));
 sg13g2_buf_2 fanout1151 (.A(_07667_),
    .X(net1151));
 sg13g2_buf_2 fanout1152 (.A(_07610_),
    .X(net1152));
 sg13g2_buf_2 fanout1153 (.A(_07520_),
    .X(net1153));
 sg13g2_buf_2 fanout1154 (.A(_07495_),
    .X(net1154));
 sg13g2_buf_2 fanout1155 (.A(_07400_),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(_07332_),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(_07279_),
    .X(net1157));
 sg13g2_buf_2 fanout1158 (.A(_07233_),
    .X(net1158));
 sg13g2_buf_2 fanout1159 (.A(_07076_),
    .X(net1159));
 sg13g2_buf_2 fanout1160 (.A(_07052_),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(_07040_),
    .X(net1161));
 sg13g2_buf_2 fanout1162 (.A(_07018_),
    .X(net1162));
 sg13g2_buf_2 fanout1163 (.A(_06998_),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(_06902_),
    .X(net1164));
 sg13g2_buf_2 fanout1165 (.A(_06837_),
    .X(net1165));
 sg13g2_buf_2 fanout1166 (.A(_06624_),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(_06532_),
    .X(net1167));
 sg13g2_buf_2 fanout1168 (.A(_06332_),
    .X(net1168));
 sg13g2_buf_2 fanout1169 (.A(_06250_),
    .X(net1169));
 sg13g2_buf_2 fanout1170 (.A(_06067_),
    .X(net1170));
 sg13g2_buf_2 fanout1171 (.A(_05936_),
    .X(net1171));
 sg13g2_buf_2 fanout1172 (.A(_05864_),
    .X(net1172));
 sg13g2_buf_2 fanout1173 (.A(_05823_),
    .X(net1173));
 sg13g2_buf_2 fanout1174 (.A(_05740_),
    .X(net1174));
 sg13g2_buf_2 fanout1175 (.A(_05419_),
    .X(net1175));
 sg13g2_buf_2 fanout1176 (.A(_05310_),
    .X(net1176));
 sg13g2_buf_2 fanout1177 (.A(_05102_),
    .X(net1177));
 sg13g2_buf_2 fanout1178 (.A(_05008_),
    .X(net1178));
 sg13g2_buf_2 fanout1179 (.A(_04950_),
    .X(net1179));
 sg13g2_buf_2 fanout1180 (.A(_04729_),
    .X(net1180));
 sg13g2_buf_2 fanout1181 (.A(_04120_),
    .X(net1181));
 sg13g2_buf_2 fanout1182 (.A(_03433_),
    .X(net1182));
 sg13g2_buf_2 fanout1183 (.A(_02863_),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(_02830_),
    .X(net1184));
 sg13g2_buf_2 fanout1185 (.A(_02173_),
    .X(net1185));
 sg13g2_buf_2 fanout1186 (.A(_02119_),
    .X(net1186));
 sg13g2_buf_2 fanout1187 (.A(_01720_),
    .X(net1187));
 sg13g2_buf_2 fanout1188 (.A(_01601_),
    .X(net1188));
 sg13g2_buf_2 fanout1189 (.A(_01579_),
    .X(net1189));
 sg13g2_buf_2 fanout1190 (.A(_01514_),
    .X(net1190));
 sg13g2_buf_2 fanout1191 (.A(_01043_),
    .X(net1191));
 sg13g2_buf_2 fanout1192 (.A(_01001_),
    .X(net1192));
 sg13g2_buf_2 fanout1193 (.A(_00798_),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(_00777_),
    .X(net1194));
 sg13g2_buf_2 fanout1195 (.A(_13246_),
    .X(net1195));
 sg13g2_buf_2 fanout1196 (.A(_13127_),
    .X(net1196));
 sg13g2_buf_2 fanout1197 (.A(_12967_),
    .X(net1197));
 sg13g2_tielo _26425__1198 (.L_LO(net1198));
 sg13g2_tielo _26426__1199 (.L_LO(net1199));
 sg13g2_tielo _26427__1200 (.L_LO(net1200));
 sg13g2_tielo _26428__1201 (.L_LO(net1201));
 sg13g2_tielo _26429__1202 (.L_LO(net1202));
 sg13g2_tielo _26430__1203 (.L_LO(net1203));
 sg13g2_tielo _26431__1204 (.L_LO(net1204));
 sg13g2_tielo _26432__1205 (.L_LO(net1205));
 sg13g2_tielo _26433__1206 (.L_LO(net1206));
 sg13g2_tielo _26434__1207 (.L_LO(net1207));
 sg13g2_tielo _26435__1208 (.L_LO(net1208));
 sg13g2_tielo _26436__1209 (.L_LO(net1209));
 sg13g2_tielo _26437__1210 (.L_LO(net1210));
 sg13g2_tielo _26438__1211 (.L_LO(net1211));
 sg13g2_tielo _26439__1212 (.L_LO(net1212));
 sg13g2_tielo _26440__1213 (.L_LO(net1213));
 sg13g2_tiehi \grid.cell_0_0.state$_SDFFE_PP0P__1215  (.L_HI(net1215));
 sg13g2_tiehi \grid.cell_0_1.state$_SDFFE_PP0P__1216  (.L_HI(net1216));
 sg13g2_tiehi \grid.cell_0_2.state$_SDFFE_PP0P__1217  (.L_HI(net1217));
 sg13g2_tiehi \grid.cell_0_3.state$_SDFFE_PP0P__1218  (.L_HI(net1218));
 sg13g2_tiehi \grid.cell_0_4.state$_SDFFE_PP0P__1219  (.L_HI(net1219));
 sg13g2_tiehi \grid.cell_0_5.state$_SDFFE_PP0P__1220  (.L_HI(net1220));
 sg13g2_tiehi \grid.cell_0_6.state$_SDFFE_PP0P__1221  (.L_HI(net1221));
 sg13g2_tiehi \grid.cell_0_7.state$_SDFFE_PP0P__1222  (.L_HI(net1222));
 sg13g2_tiehi \grid.cell_10_0.state$_SDFFE_PP0P__1223  (.L_HI(net1223));
 sg13g2_tiehi \grid.cell_10_1.state$_SDFFE_PP0P__1224  (.L_HI(net1224));
 sg13g2_tiehi \grid.cell_10_2.state$_SDFFE_PP0P__1225  (.L_HI(net1225));
 sg13g2_tiehi \grid.cell_10_3.state$_SDFFE_PP0P__1226  (.L_HI(net1226));
 sg13g2_tiehi \grid.cell_10_4.state$_SDFFE_PP0P__1227  (.L_HI(net1227));
 sg13g2_tiehi \grid.cell_10_5.state$_SDFFE_PP0P__1228  (.L_HI(net1228));
 sg13g2_tiehi \grid.cell_10_6.state$_SDFFE_PP0P__1229  (.L_HI(net1229));
 sg13g2_tiehi \grid.cell_10_7.state$_SDFFE_PP0P__1230  (.L_HI(net1230));
 sg13g2_tiehi \grid.cell_11_0.state$_SDFFE_PP0P__1231  (.L_HI(net1231));
 sg13g2_tiehi \grid.cell_11_1.state$_SDFFE_PP0P__1232  (.L_HI(net1232));
 sg13g2_tiehi \grid.cell_11_2.state$_SDFFE_PP0P__1233  (.L_HI(net1233));
 sg13g2_tiehi \grid.cell_11_3.state$_SDFFE_PP0P__1234  (.L_HI(net1234));
 sg13g2_tiehi \grid.cell_11_4.state$_SDFFE_PP0P__1235  (.L_HI(net1235));
 sg13g2_tiehi \grid.cell_11_5.state$_SDFFE_PP0P__1236  (.L_HI(net1236));
 sg13g2_tiehi \grid.cell_11_6.state$_SDFFE_PP0P__1237  (.L_HI(net1237));
 sg13g2_tiehi \grid.cell_11_7.state$_SDFFE_PP0P__1238  (.L_HI(net1238));
 sg13g2_tiehi \grid.cell_12_0.state$_SDFFE_PP0P__1239  (.L_HI(net1239));
 sg13g2_tiehi \grid.cell_12_1.state$_SDFFE_PP0P__1240  (.L_HI(net1240));
 sg13g2_tiehi \grid.cell_12_2.state$_SDFFE_PP0P__1241  (.L_HI(net1241));
 sg13g2_tiehi \grid.cell_12_3.state$_SDFFE_PP0P__1242  (.L_HI(net1242));
 sg13g2_tiehi \grid.cell_12_4.state$_SDFFE_PP0P__1243  (.L_HI(net1243));
 sg13g2_tiehi \grid.cell_12_5.state$_SDFFE_PP0P__1244  (.L_HI(net1244));
 sg13g2_tiehi \grid.cell_12_6.state$_SDFFE_PP0P__1245  (.L_HI(net1245));
 sg13g2_tiehi \grid.cell_12_7.state$_SDFFE_PP0P__1246  (.L_HI(net1246));
 sg13g2_tiehi \grid.cell_13_0.state$_SDFFE_PP0P__1247  (.L_HI(net1247));
 sg13g2_tiehi \grid.cell_13_1.state$_SDFFE_PP0P__1248  (.L_HI(net1248));
 sg13g2_tiehi \grid.cell_13_2.state$_SDFFE_PP0P__1249  (.L_HI(net1249));
 sg13g2_tiehi \grid.cell_13_3.state$_SDFFE_PP0P__1250  (.L_HI(net1250));
 sg13g2_tiehi \grid.cell_13_4.state$_SDFFE_PP0P__1251  (.L_HI(net1251));
 sg13g2_tiehi \grid.cell_13_5.state$_SDFFE_PP0P__1252  (.L_HI(net1252));
 sg13g2_tiehi \grid.cell_13_6.state$_SDFFE_PP0P__1253  (.L_HI(net1253));
 sg13g2_tiehi \grid.cell_13_7.state$_SDFFE_PP0P__1254  (.L_HI(net1254));
 sg13g2_tiehi \grid.cell_14_0.state$_SDFFE_PP0P__1255  (.L_HI(net1255));
 sg13g2_tiehi \grid.cell_14_1.state$_SDFFE_PP0P__1256  (.L_HI(net1256));
 sg13g2_tiehi \grid.cell_14_2.state$_SDFFE_PP0P__1257  (.L_HI(net1257));
 sg13g2_tiehi \grid.cell_14_3.state$_SDFFE_PP0P__1258  (.L_HI(net1258));
 sg13g2_tiehi \grid.cell_14_4.state$_SDFFE_PP0P__1259  (.L_HI(net1259));
 sg13g2_tiehi \grid.cell_14_5.state$_SDFFE_PP0P__1260  (.L_HI(net1260));
 sg13g2_tiehi \grid.cell_14_6.state$_SDFFE_PP0P__1261  (.L_HI(net1261));
 sg13g2_tiehi \grid.cell_14_7.state$_SDFFE_PP0P__1262  (.L_HI(net1262));
 sg13g2_tiehi \grid.cell_15_0.state$_SDFFE_PP0P__1263  (.L_HI(net1263));
 sg13g2_tiehi \grid.cell_15_1.state$_SDFFE_PP0P__1264  (.L_HI(net1264));
 sg13g2_tiehi \grid.cell_15_2.state$_SDFFE_PP0P__1265  (.L_HI(net1265));
 sg13g2_tiehi \grid.cell_15_3.state$_SDFFE_PP0P__1266  (.L_HI(net1266));
 sg13g2_tiehi \grid.cell_15_4.state$_SDFFE_PP0P__1267  (.L_HI(net1267));
 sg13g2_tiehi \grid.cell_15_5.state$_SDFFE_PP0P__1268  (.L_HI(net1268));
 sg13g2_tiehi \grid.cell_15_6.state$_SDFFE_PP0P__1269  (.L_HI(net1269));
 sg13g2_tiehi \grid.cell_15_7.state$_SDFFE_PP0P__1270  (.L_HI(net1270));
 sg13g2_tiehi \grid.cell_16_0.state$_SDFFE_PP0P__1271  (.L_HI(net1271));
 sg13g2_tiehi \grid.cell_16_1.state$_SDFFE_PP0P__1272  (.L_HI(net1272));
 sg13g2_tiehi \grid.cell_16_2.state$_SDFFE_PP0P__1273  (.L_HI(net1273));
 sg13g2_tiehi \grid.cell_16_3.state$_SDFFE_PP0P__1274  (.L_HI(net1274));
 sg13g2_tiehi \grid.cell_16_4.state$_SDFFE_PP0P__1275  (.L_HI(net1275));
 sg13g2_tiehi \grid.cell_16_5.state$_SDFFE_PP0P__1276  (.L_HI(net1276));
 sg13g2_tiehi \grid.cell_16_6.state$_SDFFE_PP0P__1277  (.L_HI(net1277));
 sg13g2_tiehi \grid.cell_16_7.state$_SDFFE_PP0P__1278  (.L_HI(net1278));
 sg13g2_tiehi \grid.cell_17_0.state$_SDFFE_PP0P__1279  (.L_HI(net1279));
 sg13g2_tiehi \grid.cell_17_1.state$_SDFFE_PP0P__1280  (.L_HI(net1280));
 sg13g2_tiehi \grid.cell_17_2.state$_SDFFE_PP0P__1281  (.L_HI(net1281));
 sg13g2_tiehi \grid.cell_17_3.state$_SDFFE_PP0P__1282  (.L_HI(net1282));
 sg13g2_tiehi \grid.cell_17_4.state$_SDFFE_PP0P__1283  (.L_HI(net1283));
 sg13g2_tiehi \grid.cell_17_5.state$_SDFFE_PP0P__1284  (.L_HI(net1284));
 sg13g2_tiehi \grid.cell_17_6.state$_SDFFE_PP0P__1285  (.L_HI(net1285));
 sg13g2_tiehi \grid.cell_17_7.state$_SDFFE_PP0P__1286  (.L_HI(net1286));
 sg13g2_tiehi \grid.cell_18_0.state$_SDFFE_PP0P__1287  (.L_HI(net1287));
 sg13g2_tiehi \grid.cell_18_1.state$_SDFFE_PP0P__1288  (.L_HI(net1288));
 sg13g2_tiehi \grid.cell_18_2.state$_SDFFE_PP0P__1289  (.L_HI(net1289));
 sg13g2_tiehi \grid.cell_18_3.state$_SDFFE_PP0P__1290  (.L_HI(net1290));
 sg13g2_tiehi \grid.cell_18_4.state$_SDFFE_PP0P__1291  (.L_HI(net1291));
 sg13g2_tiehi \grid.cell_18_5.state$_SDFFE_PP0P__1292  (.L_HI(net1292));
 sg13g2_tiehi \grid.cell_18_6.state$_SDFFE_PP0P__1293  (.L_HI(net1293));
 sg13g2_tiehi \grid.cell_18_7.state$_SDFFE_PP0P__1294  (.L_HI(net1294));
 sg13g2_tiehi \grid.cell_19_0.state$_SDFFE_PP0P__1295  (.L_HI(net1295));
 sg13g2_tiehi \grid.cell_19_1.state$_SDFFE_PP0P__1296  (.L_HI(net1296));
 sg13g2_tiehi \grid.cell_19_2.state$_SDFFE_PP0P__1297  (.L_HI(net1297));
 sg13g2_tiehi \grid.cell_19_3.state$_SDFFE_PP0P__1298  (.L_HI(net1298));
 sg13g2_tiehi \grid.cell_19_4.state$_SDFFE_PP0P__1299  (.L_HI(net1299));
 sg13g2_tiehi \grid.cell_19_5.state$_SDFFE_PP0P__1300  (.L_HI(net1300));
 sg13g2_tiehi \grid.cell_19_6.state$_SDFFE_PP0P__1301  (.L_HI(net1301));
 sg13g2_tiehi \grid.cell_19_7.state$_SDFFE_PP0P__1302  (.L_HI(net1302));
 sg13g2_tiehi \grid.cell_1_0.state$_SDFFE_PP0P__1303  (.L_HI(net1303));
 sg13g2_tiehi \grid.cell_1_1.state$_SDFFE_PP0P__1304  (.L_HI(net1304));
 sg13g2_tiehi \grid.cell_1_2.state$_SDFFE_PP0P__1305  (.L_HI(net1305));
 sg13g2_tiehi \grid.cell_1_3.state$_SDFFE_PP0P__1306  (.L_HI(net1306));
 sg13g2_tiehi \grid.cell_1_4.state$_SDFFE_PP0P__1307  (.L_HI(net1307));
 sg13g2_tiehi \grid.cell_1_5.state$_SDFFE_PP0P__1308  (.L_HI(net1308));
 sg13g2_tiehi \grid.cell_1_6.state$_SDFFE_PP0P__1309  (.L_HI(net1309));
 sg13g2_tiehi \grid.cell_1_7.state$_SDFFE_PP0P__1310  (.L_HI(net1310));
 sg13g2_tiehi \grid.cell_20_0.state$_SDFFE_PP0P__1311  (.L_HI(net1311));
 sg13g2_tiehi \grid.cell_20_1.state$_SDFFE_PP0P__1312  (.L_HI(net1312));
 sg13g2_tiehi \grid.cell_20_2.state$_SDFFE_PP0P__1313  (.L_HI(net1313));
 sg13g2_tiehi \grid.cell_20_3.state$_SDFFE_PP0P__1314  (.L_HI(net1314));
 sg13g2_tiehi \grid.cell_20_4.state$_SDFFE_PP0P__1315  (.L_HI(net1315));
 sg13g2_tiehi \grid.cell_20_5.state$_SDFFE_PP0P__1316  (.L_HI(net1316));
 sg13g2_tiehi \grid.cell_20_6.state$_SDFFE_PP0P__1317  (.L_HI(net1317));
 sg13g2_tiehi \grid.cell_20_7.state$_SDFFE_PP0P__1318  (.L_HI(net1318));
 sg13g2_tiehi \grid.cell_21_0.state$_SDFFE_PP0P__1319  (.L_HI(net1319));
 sg13g2_tiehi \grid.cell_21_1.state$_SDFFE_PP0P__1320  (.L_HI(net1320));
 sg13g2_tiehi \grid.cell_21_2.state$_SDFFE_PP0P__1321  (.L_HI(net1321));
 sg13g2_tiehi \grid.cell_21_3.state$_SDFFE_PP0P__1322  (.L_HI(net1322));
 sg13g2_tiehi \grid.cell_21_4.state$_SDFFE_PP0P__1323  (.L_HI(net1323));
 sg13g2_tiehi \grid.cell_21_5.state$_SDFFE_PP0P__1324  (.L_HI(net1324));
 sg13g2_tiehi \grid.cell_21_6.state$_SDFFE_PP0P__1325  (.L_HI(net1325));
 sg13g2_tiehi \grid.cell_21_7.state$_SDFFE_PP0P__1326  (.L_HI(net1326));
 sg13g2_tiehi \grid.cell_22_0.state$_SDFFE_PP0P__1327  (.L_HI(net1327));
 sg13g2_tiehi \grid.cell_22_1.state$_SDFFE_PP0P__1328  (.L_HI(net1328));
 sg13g2_tiehi \grid.cell_22_2.state$_SDFFE_PP0P__1329  (.L_HI(net1329));
 sg13g2_tiehi \grid.cell_22_3.state$_SDFFE_PP0P__1330  (.L_HI(net1330));
 sg13g2_tiehi \grid.cell_22_4.state$_SDFFE_PP0P__1331  (.L_HI(net1331));
 sg13g2_tiehi \grid.cell_22_5.state$_SDFFE_PP0P__1332  (.L_HI(net1332));
 sg13g2_tiehi \grid.cell_22_6.state$_SDFFE_PP0P__1333  (.L_HI(net1333));
 sg13g2_tiehi \grid.cell_22_7.state$_SDFFE_PP0P__1334  (.L_HI(net1334));
 sg13g2_tiehi \grid.cell_23_0.state$_SDFFE_PP0P__1335  (.L_HI(net1335));
 sg13g2_tiehi \grid.cell_23_1.state$_SDFFE_PP0P__1336  (.L_HI(net1336));
 sg13g2_tiehi \grid.cell_23_2.state$_SDFFE_PP0P__1337  (.L_HI(net1337));
 sg13g2_tiehi \grid.cell_23_3.state$_SDFFE_PP0P__1338  (.L_HI(net1338));
 sg13g2_tiehi \grid.cell_23_4.state$_SDFFE_PP0P__1339  (.L_HI(net1339));
 sg13g2_tiehi \grid.cell_23_5.state$_SDFFE_PP0P__1340  (.L_HI(net1340));
 sg13g2_tiehi \grid.cell_23_6.state$_SDFFE_PP0P__1341  (.L_HI(net1341));
 sg13g2_tiehi \grid.cell_23_7.state$_SDFFE_PP0P__1342  (.L_HI(net1342));
 sg13g2_tiehi \grid.cell_24_0.state$_SDFFE_PP0P__1343  (.L_HI(net1343));
 sg13g2_tiehi \grid.cell_24_1.state$_SDFFE_PP0P__1344  (.L_HI(net1344));
 sg13g2_tiehi \grid.cell_24_2.state$_SDFFE_PP0P__1345  (.L_HI(net1345));
 sg13g2_tiehi \grid.cell_24_3.state$_SDFFE_PP0P__1346  (.L_HI(net1346));
 sg13g2_tiehi \grid.cell_24_4.state$_SDFFE_PP0P__1347  (.L_HI(net1347));
 sg13g2_tiehi \grid.cell_24_5.state$_SDFFE_PP0P__1348  (.L_HI(net1348));
 sg13g2_tiehi \grid.cell_24_6.state$_SDFFE_PP0P__1349  (.L_HI(net1349));
 sg13g2_tiehi \grid.cell_24_7.state$_SDFFE_PP0P__1350  (.L_HI(net1350));
 sg13g2_tiehi \grid.cell_25_0.state$_SDFFE_PP0P__1351  (.L_HI(net1351));
 sg13g2_tiehi \grid.cell_25_1.state$_SDFFE_PP0P__1352  (.L_HI(net1352));
 sg13g2_tiehi \grid.cell_25_2.state$_SDFFE_PP0P__1353  (.L_HI(net1353));
 sg13g2_tiehi \grid.cell_25_3.state$_SDFFE_PP0P__1354  (.L_HI(net1354));
 sg13g2_tiehi \grid.cell_25_4.state$_SDFFE_PP0P__1355  (.L_HI(net1355));
 sg13g2_tiehi \grid.cell_25_5.state$_SDFFE_PP0P__1356  (.L_HI(net1356));
 sg13g2_tiehi \grid.cell_25_6.state$_SDFFE_PP0P__1357  (.L_HI(net1357));
 sg13g2_tiehi \grid.cell_25_7.state$_SDFFE_PP0P__1358  (.L_HI(net1358));
 sg13g2_tiehi \grid.cell_26_0.state$_SDFFE_PP0P__1359  (.L_HI(net1359));
 sg13g2_tiehi \grid.cell_26_1.state$_SDFFE_PP0P__1360  (.L_HI(net1360));
 sg13g2_tiehi \grid.cell_26_2.state$_SDFFE_PP0P__1361  (.L_HI(net1361));
 sg13g2_tiehi \grid.cell_26_3.state$_SDFFE_PP0P__1362  (.L_HI(net1362));
 sg13g2_tiehi \grid.cell_26_4.state$_SDFFE_PP0P__1363  (.L_HI(net1363));
 sg13g2_tiehi \grid.cell_26_5.state$_SDFFE_PP0P__1364  (.L_HI(net1364));
 sg13g2_tiehi \grid.cell_26_6.state$_SDFFE_PP0P__1365  (.L_HI(net1365));
 sg13g2_tiehi \grid.cell_26_7.state$_SDFFE_PP0P__1366  (.L_HI(net1366));
 sg13g2_tiehi \grid.cell_27_0.state$_SDFFE_PP0P__1367  (.L_HI(net1367));
 sg13g2_tiehi \grid.cell_27_1.state$_SDFFE_PP0P__1368  (.L_HI(net1368));
 sg13g2_tiehi \grid.cell_27_2.state$_SDFFE_PP0P__1369  (.L_HI(net1369));
 sg13g2_tiehi \grid.cell_27_3.state$_SDFFE_PP0P__1370  (.L_HI(net1370));
 sg13g2_tiehi \grid.cell_27_4.state$_SDFFE_PP0P__1371  (.L_HI(net1371));
 sg13g2_tiehi \grid.cell_27_5.state$_SDFFE_PP0P__1372  (.L_HI(net1372));
 sg13g2_tiehi \grid.cell_27_6.state$_SDFFE_PP0P__1373  (.L_HI(net1373));
 sg13g2_tiehi \grid.cell_27_7.state$_SDFFE_PP0P__1374  (.L_HI(net1374));
 sg13g2_tiehi \grid.cell_28_0.state$_SDFFE_PP0P__1375  (.L_HI(net1375));
 sg13g2_tiehi \grid.cell_28_1.state$_SDFFE_PP0P__1376  (.L_HI(net1376));
 sg13g2_tiehi \grid.cell_28_2.state$_SDFFE_PP0P__1377  (.L_HI(net1377));
 sg13g2_tiehi \grid.cell_28_3.state$_SDFFE_PP0P__1378  (.L_HI(net1378));
 sg13g2_tiehi \grid.cell_28_4.state$_SDFFE_PP0P__1379  (.L_HI(net1379));
 sg13g2_tiehi \grid.cell_28_5.state$_SDFFE_PP0P__1380  (.L_HI(net1380));
 sg13g2_tiehi \grid.cell_28_6.state$_SDFFE_PP0P__1381  (.L_HI(net1381));
 sg13g2_tiehi \grid.cell_28_7.state$_SDFFE_PP0P__1382  (.L_HI(net1382));
 sg13g2_tiehi \grid.cell_29_0.state$_SDFFE_PP0P__1383  (.L_HI(net1383));
 sg13g2_tiehi \grid.cell_29_1.state$_SDFFE_PP0P__1384  (.L_HI(net1384));
 sg13g2_tiehi \grid.cell_29_2.state$_SDFFE_PP0P__1385  (.L_HI(net1385));
 sg13g2_tiehi \grid.cell_29_3.state$_SDFFE_PP0P__1386  (.L_HI(net1386));
 sg13g2_tiehi \grid.cell_29_4.state$_SDFFE_PP0P__1387  (.L_HI(net1387));
 sg13g2_tiehi \grid.cell_29_5.state$_SDFFE_PP0P__1388  (.L_HI(net1388));
 sg13g2_tiehi \grid.cell_29_6.state$_SDFFE_PP0P__1389  (.L_HI(net1389));
 sg13g2_tiehi \grid.cell_29_7.state$_SDFFE_PP0P__1390  (.L_HI(net1390));
 sg13g2_tiehi \grid.cell_2_0.state$_SDFFE_PP0P__1391  (.L_HI(net1391));
 sg13g2_tiehi \grid.cell_2_1.state$_SDFFE_PP0P__1392  (.L_HI(net1392));
 sg13g2_tiehi \grid.cell_2_2.state$_SDFFE_PP0P__1393  (.L_HI(net1393));
 sg13g2_tiehi \grid.cell_2_3.state$_SDFFE_PP0P__1394  (.L_HI(net1394));
 sg13g2_tiehi \grid.cell_2_4.state$_SDFFE_PP0P__1395  (.L_HI(net1395));
 sg13g2_tiehi \grid.cell_2_5.state$_SDFFE_PP0P__1396  (.L_HI(net1396));
 sg13g2_tiehi \grid.cell_2_6.state$_SDFFE_PP0P__1397  (.L_HI(net1397));
 sg13g2_tiehi \grid.cell_2_7.state$_SDFFE_PP0P__1398  (.L_HI(net1398));
 sg13g2_tiehi \grid.cell_30_0.state$_SDFFE_PP0P__1399  (.L_HI(net1399));
 sg13g2_tiehi \grid.cell_30_1.state$_SDFFE_PP0P__1400  (.L_HI(net1400));
 sg13g2_tiehi \grid.cell_30_2.state$_SDFFE_PP0P__1401  (.L_HI(net1401));
 sg13g2_tiehi \grid.cell_30_3.state$_SDFFE_PP0P__1402  (.L_HI(net1402));
 sg13g2_tiehi \grid.cell_30_4.state$_SDFFE_PP0P__1403  (.L_HI(net1403));
 sg13g2_tiehi \grid.cell_30_5.state$_SDFFE_PP0P__1404  (.L_HI(net1404));
 sg13g2_tiehi \grid.cell_30_6.state$_SDFFE_PP0P__1405  (.L_HI(net1405));
 sg13g2_tiehi \grid.cell_30_7.state$_SDFFE_PP0P__1406  (.L_HI(net1406));
 sg13g2_tiehi \grid.cell_31_0.state$_SDFFE_PP0P__1407  (.L_HI(net1407));
 sg13g2_tiehi \grid.cell_31_1.state$_SDFFE_PP0P__1408  (.L_HI(net1408));
 sg13g2_tiehi \grid.cell_31_2.state$_SDFFE_PP0P__1409  (.L_HI(net1409));
 sg13g2_tiehi \grid.cell_31_3.state$_SDFFE_PP0P__1410  (.L_HI(net1410));
 sg13g2_tiehi \grid.cell_31_4.state$_SDFFE_PP0P__1411  (.L_HI(net1411));
 sg13g2_tiehi \grid.cell_31_5.state$_SDFFE_PP0P__1412  (.L_HI(net1412));
 sg13g2_tiehi \grid.cell_31_6.state$_SDFFE_PP0P__1413  (.L_HI(net1413));
 sg13g2_tiehi \grid.cell_31_7.state$_SDFFE_PP0P__1414  (.L_HI(net1414));
 sg13g2_tiehi \grid.cell_3_0.state$_SDFFE_PP0P__1415  (.L_HI(net1415));
 sg13g2_tiehi \grid.cell_3_1.state$_SDFFE_PP0P__1416  (.L_HI(net1416));
 sg13g2_tiehi \grid.cell_3_2.state$_SDFFE_PP0P__1417  (.L_HI(net1417));
 sg13g2_tiehi \grid.cell_3_3.state$_SDFFE_PP0P__1418  (.L_HI(net1418));
 sg13g2_tiehi \grid.cell_3_4.state$_SDFFE_PP0P__1419  (.L_HI(net1419));
 sg13g2_tiehi \grid.cell_3_5.state$_SDFFE_PP0P__1420  (.L_HI(net1420));
 sg13g2_tiehi \grid.cell_3_6.state$_SDFFE_PP0P__1421  (.L_HI(net1421));
 sg13g2_tiehi \grid.cell_3_7.state$_SDFFE_PP0P__1422  (.L_HI(net1422));
 sg13g2_tiehi \grid.cell_4_0.state$_SDFFE_PP0P__1423  (.L_HI(net1423));
 sg13g2_tiehi \grid.cell_4_1.state$_SDFFE_PP0P__1424  (.L_HI(net1424));
 sg13g2_tiehi \grid.cell_4_2.state$_SDFFE_PP0P__1425  (.L_HI(net1425));
 sg13g2_tiehi \grid.cell_4_3.state$_SDFFE_PP0P__1426  (.L_HI(net1426));
 sg13g2_tiehi \grid.cell_4_4.state$_SDFFE_PP0P__1427  (.L_HI(net1427));
 sg13g2_tiehi \grid.cell_4_5.state$_SDFFE_PP0P__1428  (.L_HI(net1428));
 sg13g2_tiehi \grid.cell_4_6.state$_SDFFE_PP0P__1429  (.L_HI(net1429));
 sg13g2_tiehi \grid.cell_4_7.state$_SDFFE_PP0P__1430  (.L_HI(net1430));
 sg13g2_tiehi \grid.cell_5_0.state$_SDFFE_PP0P__1431  (.L_HI(net1431));
 sg13g2_tiehi \grid.cell_5_1.state$_SDFFE_PP0P__1432  (.L_HI(net1432));
 sg13g2_tiehi \grid.cell_5_2.state$_SDFFE_PP0P__1433  (.L_HI(net1433));
 sg13g2_tiehi \grid.cell_5_3.state$_SDFFE_PP0P__1434  (.L_HI(net1434));
 sg13g2_tiehi \grid.cell_5_4.state$_SDFFE_PP0P__1435  (.L_HI(net1435));
 sg13g2_tiehi \grid.cell_5_5.state$_SDFFE_PP0P__1436  (.L_HI(net1436));
 sg13g2_tiehi \grid.cell_5_6.state$_SDFFE_PP0P__1437  (.L_HI(net1437));
 sg13g2_tiehi \grid.cell_5_7.state$_SDFFE_PP0P__1438  (.L_HI(net1438));
 sg13g2_tiehi \grid.cell_6_0.state$_SDFFE_PP0P__1439  (.L_HI(net1439));
 sg13g2_tiehi \grid.cell_6_1.state$_SDFFE_PP0P__1440  (.L_HI(net1440));
 sg13g2_tiehi \grid.cell_6_2.state$_SDFFE_PP0P__1441  (.L_HI(net1441));
 sg13g2_tiehi \grid.cell_6_3.state$_SDFFE_PP0P__1442  (.L_HI(net1442));
 sg13g2_tiehi \grid.cell_6_4.state$_SDFFE_PP0P__1443  (.L_HI(net1443));
 sg13g2_tiehi \grid.cell_6_5.state$_SDFFE_PP0P__1444  (.L_HI(net1444));
 sg13g2_tiehi \grid.cell_6_6.state$_SDFFE_PP0P__1445  (.L_HI(net1445));
 sg13g2_tiehi \grid.cell_6_7.state$_SDFFE_PP0P__1446  (.L_HI(net1446));
 sg13g2_tiehi \grid.cell_7_0.state$_SDFFE_PP0P__1447  (.L_HI(net1447));
 sg13g2_tiehi \grid.cell_7_1.state$_SDFFE_PP0P__1448  (.L_HI(net1448));
 sg13g2_tiehi \grid.cell_7_2.state$_SDFFE_PP0P__1449  (.L_HI(net1449));
 sg13g2_tiehi \grid.cell_7_3.state$_SDFFE_PP0P__1450  (.L_HI(net1450));
 sg13g2_tiehi \grid.cell_7_4.state$_SDFFE_PP0P__1451  (.L_HI(net1451));
 sg13g2_tiehi \grid.cell_7_5.state$_SDFFE_PP0P__1452  (.L_HI(net1452));
 sg13g2_tiehi \grid.cell_7_6.state$_SDFFE_PP0P__1453  (.L_HI(net1453));
 sg13g2_tiehi \grid.cell_7_7.state$_SDFFE_PP0P__1454  (.L_HI(net1454));
 sg13g2_tiehi \grid.cell_8_0.state$_SDFFE_PP0P__1455  (.L_HI(net1455));
 sg13g2_tiehi \grid.cell_8_1.state$_SDFFE_PP0P__1456  (.L_HI(net1456));
 sg13g2_tiehi \grid.cell_8_2.state$_SDFFE_PP0P__1457  (.L_HI(net1457));
 sg13g2_tiehi \grid.cell_8_3.state$_SDFFE_PP0P__1458  (.L_HI(net1458));
 sg13g2_tiehi \grid.cell_8_4.state$_SDFFE_PP0P__1459  (.L_HI(net1459));
 sg13g2_tiehi \grid.cell_8_5.state$_SDFFE_PP0P__1460  (.L_HI(net1460));
 sg13g2_tiehi \grid.cell_8_6.state$_SDFFE_PP0P__1461  (.L_HI(net1461));
 sg13g2_tiehi \grid.cell_8_7.state$_SDFFE_PP0P__1462  (.L_HI(net1462));
 sg13g2_tiehi \grid.cell_9_0.state$_SDFFE_PP0P__1463  (.L_HI(net1463));
 sg13g2_tiehi \grid.cell_9_1.state$_SDFFE_PP0P__1464  (.L_HI(net1464));
 sg13g2_tiehi \grid.cell_9_2.state$_SDFFE_PP0P__1465  (.L_HI(net1465));
 sg13g2_tiehi \grid.cell_9_3.state$_SDFFE_PP0P__1466  (.L_HI(net1466));
 sg13g2_tiehi \grid.cell_9_4.state$_SDFFE_PP0P__1467  (.L_HI(net1467));
 sg13g2_tiehi \grid.cell_9_5.state$_SDFFE_PP0P__1468  (.L_HI(net1468));
 sg13g2_tiehi \grid.cell_9_6.state$_SDFFE_PP0P__1469  (.L_HI(net1469));
 sg13g2_tiehi \grid.cell_9_7.state$_SDFFE_PP0P__1470  (.L_HI(net1470));
 sg13g2_tiehi \max7219.col_index[0]$_SDFF_PN0__1471  (.L_HI(net1471));
 sg13g2_tiehi \max7219.col_index[1]$_SDFF_PN0__1472  (.L_HI(net1472));
 sg13g2_tiehi \max7219.col_index[2]$_SDFF_PN0__1473  (.L_HI(net1473));
 sg13g2_tiehi \max7219.init_index[0]$_SDFFE_PN0P__1474  (.L_HI(net1474));
 sg13g2_tiehi \max7219.init_index[1]$_SDFFE_PN0P__1475  (.L_HI(net1475));
 sg13g2_tiehi \max7219.load_row$_SDFF_PN0__1476  (.L_HI(net1476));
 sg13g2_tiehi \max7219.matrix_index[0]$_SDFFE_PN0P__1477  (.L_HI(net1477));
 sg13g2_tiehi \max7219.matrix_index[1]$_SDFFE_PN0P__1478  (.L_HI(net1478));
 sg13g2_tiehi \max7219.max7219_enabled$_SDFFE_PN0P__1479  (.L_HI(net1479));
 sg13g2_tiehi \max7219.max7219_row[0]$_SDFFE_PN0P__1480  (.L_HI(net1480));
 sg13g2_tiehi \max7219.max7219_row[1]$_SDFFE_PN0P__1481  (.L_HI(net1481));
 sg13g2_tiehi \max7219.max7219_row[2]$_SDFFE_PN0P__1482  (.L_HI(net1482));
 sg13g2_tiehi \max7219.o_cs$_SDFFE_PN1P__1483  (.L_HI(net1483));
 sg13g2_tiehi \max7219.row_data[0]$_SDFFE_PN0P__1484  (.L_HI(net1484));
 sg13g2_tiehi \max7219.row_data[1]$_SDFFE_PN0P__1485  (.L_HI(net1485));
 sg13g2_tiehi \max7219.row_data[2]$_SDFFE_PN0P__1486  (.L_HI(net1486));
 sg13g2_tiehi \max7219.row_data[3]$_SDFFE_PN0P__1487  (.L_HI(net1487));
 sg13g2_tiehi \max7219.row_data[4]$_SDFFE_PN0P__1488  (.L_HI(net1488));
 sg13g2_tiehi \max7219.row_data[5]$_SDFFE_PN0P__1489  (.L_HI(net1489));
 sg13g2_tiehi \max7219.row_data[6]$_SDFFE_PN0P__1490  (.L_HI(net1490));
 sg13g2_tiehi \max7219.row_data[7]$_SDFFE_PN0P__1491  (.L_HI(net1491));
 sg13g2_tiehi \max7219.spi_start$_SDFF_PN0__1492  (.L_HI(net1492));
 sg13g2_tiehi \max7219.spim.bit_index[0]$_SDFFE_PN1P__1493  (.L_HI(net1493));
 sg13g2_tiehi \max7219.spim.bit_index[1]$_SDFFE_PN1P__1494  (.L_HI(net1494));
 sg13g2_tiehi \max7219.spim.bit_index[2]$_SDFFE_PN1P__1495  (.L_HI(net1495));
 sg13g2_tiehi \max7219.spim.bit_index[3]$_SDFFE_PN1P__1496  (.L_HI(net1496));
 sg13g2_tiehi \max7219.spim.clk_count[0]$_SDFFE_PP0P__1497  (.L_HI(net1497));
 sg13g2_tiehi \max7219.spim.clk_count[1]$_SDFFE_PP0P__1498  (.L_HI(net1498));
 sg13g2_tiehi \max7219.spim.finish$_SDFFCE_PP0P__1499  (.L_HI(net1499));
 sg13g2_tiehi \max7219.spim.o_busy$_SDFF_PP0__1500  (.L_HI(net1500));
 sg13g2_tiehi \max7219.spim.o_mosi$_SDFFE_PN0P__1501  (.L_HI(net1501));
 sg13g2_tiehi \max7219.spim.o_sck$_SDFFE_PP0P__1502  (.L_HI(net1502));
 sg13g2_tiehi \max7219.state[0]$_DFF_P__1503  (.L_HI(net1503));
 sg13g2_tiehi \max7219.state[1]$_DFF_P__1504  (.L_HI(net1504));
 sg13g2_tiehi \max7219.state[2]$_DFF_P__1505  (.L_HI(net1505));
 sg13g2_tiehi \max7219.state[3]$_DFF_P__1506  (.L_HI(net1506));
 sg13g2_tiehi \prev_rst_n$_DFF_P__1507  (.L_HI(net1507));
 sg13g2_tiehi \silife_demo_inst.counter[0]$_SDFFE_PN0P__1508  (.L_HI(net1508));
 sg13g2_tiehi \silife_demo_inst.counter[10]$_SDFFE_PN0P__1509  (.L_HI(net1509));
 sg13g2_tiehi \silife_demo_inst.counter[11]$_SDFFE_PN0P__1510  (.L_HI(net1510));
 sg13g2_tiehi \silife_demo_inst.counter[12]$_SDFFE_PN0P__1511  (.L_HI(net1511));
 sg13g2_tiehi \silife_demo_inst.counter[13]$_SDFFE_PN0P__1512  (.L_HI(net1512));
 sg13g2_tiehi \silife_demo_inst.counter[14]$_SDFFE_PN0P__1513  (.L_HI(net1513));
 sg13g2_tiehi \silife_demo_inst.counter[15]$_SDFFE_PN0P__1514  (.L_HI(net1514));
 sg13g2_tiehi \silife_demo_inst.counter[16]$_SDFFE_PN0P__1515  (.L_HI(net1515));
 sg13g2_tiehi \silife_demo_inst.counter[17]$_SDFFE_PN0P__1516  (.L_HI(net1516));
 sg13g2_tiehi \silife_demo_inst.counter[18]$_SDFFE_PN0P__1517  (.L_HI(net1517));
 sg13g2_tiehi \silife_demo_inst.counter[19]$_SDFFE_PN0P__1518  (.L_HI(net1518));
 sg13g2_tiehi \silife_demo_inst.counter[1]$_SDFFE_PN0P__1519  (.L_HI(net1519));
 sg13g2_tiehi \silife_demo_inst.counter[20]$_SDFFE_PN0P__1520  (.L_HI(net1520));
 sg13g2_tiehi \silife_demo_inst.counter[21]$_SDFFE_PN0P__1521  (.L_HI(net1521));
 sg13g2_tiehi \silife_demo_inst.counter[22]$_SDFFE_PN0P__1522  (.L_HI(net1522));
 sg13g2_tiehi \silife_demo_inst.counter[23]$_SDFFE_PN0P__1523  (.L_HI(net1523));
 sg13g2_tiehi \silife_demo_inst.counter[24]$_SDFFE_PN0P__1524  (.L_HI(net1524));
 sg13g2_tiehi \silife_demo_inst.counter[25]$_SDFFE_PN0P__1525  (.L_HI(net1525));
 sg13g2_tiehi \silife_demo_inst.counter[26]$_SDFFE_PN0P__1526  (.L_HI(net1526));
 sg13g2_tiehi \silife_demo_inst.counter[27]$_SDFFE_PN0P__1527  (.L_HI(net1527));
 sg13g2_tiehi \silife_demo_inst.counter[28]$_SDFFE_PN0P__1528  (.L_HI(net1528));
 sg13g2_tiehi \silife_demo_inst.counter[29]$_SDFFE_PN0P__1529  (.L_HI(net1529));
 sg13g2_tiehi \silife_demo_inst.counter[2]$_SDFFE_PN0P__1530  (.L_HI(net1530));
 sg13g2_tiehi \silife_demo_inst.counter[30]$_SDFFE_PN0P__1531  (.L_HI(net1531));
 sg13g2_tiehi \silife_demo_inst.counter[31]$_SDFFE_PN0P__1532  (.L_HI(net1532));
 sg13g2_tiehi \silife_demo_inst.counter[3]$_SDFFE_PN0P__1533  (.L_HI(net1533));
 sg13g2_tiehi \silife_demo_inst.counter[4]$_SDFFE_PN0P__1534  (.L_HI(net1534));
 sg13g2_tiehi \silife_demo_inst.counter[5]$_SDFFE_PN0P__1535  (.L_HI(net1535));
 sg13g2_tiehi \silife_demo_inst.counter[6]$_SDFFE_PN0P__1536  (.L_HI(net1536));
 sg13g2_tiehi \silife_demo_inst.counter[7]$_SDFFE_PN0P__1537  (.L_HI(net1537));
 sg13g2_tiehi \silife_demo_inst.counter[8]$_SDFFE_PN0P__1538  (.L_HI(net1538));
 sg13g2_tiehi \silife_demo_inst.counter[9]$_SDFFE_PN0P__1539  (.L_HI(net1539));
 sg13g2_tiehi \silife_demo_inst.init_done$_SDFFE_PN0P__1540  (.L_HI(net1540));
 sg13g2_tiehi \silife_demo_inst.row_select[0]$_SDFFE_PN0P__1541  (.L_HI(net1541));
 sg13g2_tiehi \silife_demo_inst.row_select[1]$_SDFFE_PN0P__1542  (.L_HI(net1542));
 sg13g2_tiehi \silife_demo_inst.row_select[2]$_SDFFE_PN0P__1543  (.L_HI(net1543));
 sg13g2_tiehi \silife_demo_inst.row_select[3]$_SDFFE_PN0P__1544  (.L_HI(net1544));
 sg13g2_tiehi \silife_demo_inst.row_select[4]$_SDFFE_PN0P__1545  (.L_HI(net1545));
 sg13g2_tiehi \silife_demo_inst.step$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \silife_demo_inst.wr_en$_SDFFE_PN0N__1547  (.L_HI(net1547));
 sg13g2_tiehi \wr_available$_SDFFE_PN0N__1548  (.L_HI(net1548));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_4_0__f_clk (.X(clknet_4_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_4_1__f_clk (.X(clknet_4_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_4_2__f_clk (.X(clknet_4_2__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_4_3__f_clk (.X(clknet_4_3__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_4_4__f_clk (.X(clknet_4_4__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_4_5__f_clk (.X(clknet_4_5__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_4_6__f_clk (.X(clknet_4_6__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_4_7__f_clk (.X(clknet_4_7__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_4_8__f_clk (.X(clknet_4_8__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_4_9__f_clk (.X(clknet_4_9__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_4_10__f_clk (.X(clknet_4_10__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_4_11__f_clk (.X(clknet_4_11__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_4_12__f_clk (.X(clknet_4_12__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_4_13__f_clk (.X(clknet_4_13__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_4_14__f_clk (.X(clknet_4_14__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_4_15__f_clk (.X(clknet_4_15__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_16 clkload0 (.A(clknet_4_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_7__leaf_clk));
 sg13g2_buf_16 clkload2 (.A(clknet_4_11__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_4_13__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_4_15__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_72_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_73_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_74_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_2_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_3_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_67_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_leaf_69_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_70_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_leaf_71_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_65_clk));
 sg13g2_buf_16 clkload18 (.A(clknet_leaf_11_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_leaf_13_clk));
 sg13g2_buf_16 clkload20 (.A(clknet_leaf_14_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_15_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_17_clk));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_22_clk));
 sg13g2_buf_8 clkload24 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_23_clk));
 sg13g2_inv_2 clkload26 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_24_clk));
 sg13g2_buf_16 clkload28 (.A(clknet_leaf_26_clk));
 sg13g2_buf_16 clkload29 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_60_clk));
 sg13g2_buf_8 clkload31 (.A(clknet_leaf_62_clk));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_63_clk));
 sg13g2_buf_8 clkload33 (.A(clknet_leaf_64_clk));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_29_clk));
 sg13g2_buf_16 clkload35 (.A(clknet_leaf_46_clk));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_48_clk));
 sg13g2_inv_1 clkload37 (.A(clknet_leaf_55_clk));
 sg13g2_inv_2 clkload38 (.A(clknet_leaf_59_clk));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_49_clk));
 sg13g2_inv_2 clkload40 (.A(clknet_leaf_30_clk));
 sg13g2_buf_16 clkload41 (.A(clknet_leaf_31_clk));
 sg13g2_buf_16 clkload42 (.A(clknet_leaf_44_clk));
 sg13g2_buf_8 clkload43 (.A(clknet_leaf_45_clk));
 sg13g2_buf_16 clkload44 (.A(clknet_leaf_32_clk));
 sg13g2_buf_8 clkload45 (.A(clknet_leaf_34_clk));
 sg13g2_buf_8 clkload46 (.A(clknet_leaf_35_clk));
 sg13g2_inv_2 clkload47 (.A(clknet_leaf_41_clk));
 sg13g2_buf_8 clkload48 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload49 (.A(clknet_leaf_52_clk));
 sg13g2_inv_1 clkload50 (.A(clknet_leaf_53_clk));
 sg13g2_buf_8 clkload51 (.A(clknet_leaf_40_clk));
 sg13g2_buf_1 fanout1 (.A(_04734_),
    .X(net1549));
 sg13g2_antennanp ANTENNA_1 (.A(_00387_));
 sg13g2_antennanp ANTENNA_2 (.A(_00461_));
 sg13g2_antennanp ANTENNA_3 (.A(_01440_));
 sg13g2_antennanp ANTENNA_4 (.A(_01440_));
 sg13g2_antennanp ANTENNA_5 (.A(_01795_));
 sg13g2_antennanp ANTENNA_6 (.A(_01795_));
 sg13g2_antennanp ANTENNA_7 (.A(_02776_));
 sg13g2_antennanp ANTENNA_8 (.A(_02776_));
 sg13g2_antennanp ANTENNA_9 (.A(_02776_));
 sg13g2_antennanp ANTENNA_10 (.A(_02776_));
 sg13g2_antennanp ANTENNA_11 (.A(_02787_));
 sg13g2_antennanp ANTENNA_12 (.A(_02787_));
 sg13g2_antennanp ANTENNA_13 (.A(_02787_));
 sg13g2_antennanp ANTENNA_14 (.A(_02787_));
 sg13g2_antennanp ANTENNA_15 (.A(_02787_));
 sg13g2_antennanp ANTENNA_16 (.A(_02787_));
 sg13g2_antennanp ANTENNA_17 (.A(_03810_));
 sg13g2_antennanp ANTENNA_18 (.A(_03810_));
 sg13g2_antennanp ANTENNA_19 (.A(_03810_));
 sg13g2_antennanp ANTENNA_20 (.A(_03810_));
 sg13g2_antennanp ANTENNA_21 (.A(_03810_));
 sg13g2_antennanp ANTENNA_22 (.A(_03810_));
 sg13g2_antennanp ANTENNA_23 (.A(_03810_));
 sg13g2_antennanp ANTENNA_24 (.A(_03821_));
 sg13g2_antennanp ANTENNA_25 (.A(_03821_));
 sg13g2_antennanp ANTENNA_26 (.A(_03821_));
 sg13g2_antennanp ANTENNA_27 (.A(_03821_));
 sg13g2_antennanp ANTENNA_28 (.A(_04067_));
 sg13g2_antennanp ANTENNA_29 (.A(_04067_));
 sg13g2_antennanp ANTENNA_30 (.A(_04067_));
 sg13g2_antennanp ANTENNA_31 (.A(_04067_));
 sg13g2_antennanp ANTENNA_32 (.A(_04067_));
 sg13g2_antennanp ANTENNA_33 (.A(_04067_));
 sg13g2_antennanp ANTENNA_34 (.A(_04067_));
 sg13g2_antennanp ANTENNA_35 (.A(_04067_));
 sg13g2_antennanp ANTENNA_36 (.A(_04077_));
 sg13g2_antennanp ANTENNA_37 (.A(_04077_));
 sg13g2_antennanp ANTENNA_38 (.A(_04077_));
 sg13g2_antennanp ANTENNA_39 (.A(_04077_));
 sg13g2_antennanp ANTENNA_40 (.A(_04077_));
 sg13g2_antennanp ANTENNA_41 (.A(_04242_));
 sg13g2_antennanp ANTENNA_42 (.A(_04242_));
 sg13g2_antennanp ANTENNA_43 (.A(_04371_));
 sg13g2_antennanp ANTENNA_44 (.A(_04378_));
 sg13g2_antennanp ANTENNA_45 (.A(_04393_));
 sg13g2_antennanp ANTENNA_46 (.A(_04399_));
 sg13g2_antennanp ANTENNA_47 (.A(_04403_));
 sg13g2_antennanp ANTENNA_48 (.A(_04411_));
 sg13g2_antennanp ANTENNA_49 (.A(_04412_));
 sg13g2_antennanp ANTENNA_50 (.A(_04416_));
 sg13g2_antennanp ANTENNA_51 (.A(_04419_));
 sg13g2_antennanp ANTENNA_52 (.A(_04432_));
 sg13g2_antennanp ANTENNA_53 (.A(_04453_));
 sg13g2_antennanp ANTENNA_54 (.A(_04481_));
 sg13g2_antennanp ANTENNA_55 (.A(_04508_));
 sg13g2_antennanp ANTENNA_56 (.A(_04508_));
 sg13g2_antennanp ANTENNA_57 (.A(_04747_));
 sg13g2_antennanp ANTENNA_58 (.A(_04756_));
 sg13g2_antennanp ANTENNA_59 (.A(_04773_));
 sg13g2_antennanp ANTENNA_60 (.A(_04804_));
 sg13g2_antennanp ANTENNA_61 (.A(_04816_));
 sg13g2_antennanp ANTENNA_62 (.A(_04817_));
 sg13g2_antennanp ANTENNA_63 (.A(_04828_));
 sg13g2_antennanp ANTENNA_64 (.A(_04838_));
 sg13g2_antennanp ANTENNA_65 (.A(_04840_));
 sg13g2_antennanp ANTENNA_66 (.A(_04842_));
 sg13g2_antennanp ANTENNA_67 (.A(_04843_));
 sg13g2_antennanp ANTENNA_68 (.A(_04850_));
 sg13g2_antennanp ANTENNA_69 (.A(_04853_));
 sg13g2_antennanp ANTENNA_70 (.A(_04860_));
 sg13g2_antennanp ANTENNA_71 (.A(_04860_));
 sg13g2_antennanp ANTENNA_72 (.A(_04860_));
 sg13g2_antennanp ANTENNA_73 (.A(_04860_));
 sg13g2_antennanp ANTENNA_74 (.A(_04860_));
 sg13g2_antennanp ANTENNA_75 (.A(_04914_));
 sg13g2_antennanp ANTENNA_76 (.A(_04914_));
 sg13g2_antennanp ANTENNA_77 (.A(_04941_));
 sg13g2_antennanp ANTENNA_78 (.A(_04941_));
 sg13g2_antennanp ANTENNA_79 (.A(_04941_));
 sg13g2_antennanp ANTENNA_80 (.A(_04941_));
 sg13g2_antennanp ANTENNA_81 (.A(_04941_));
 sg13g2_antennanp ANTENNA_82 (.A(_04941_));
 sg13g2_antennanp ANTENNA_83 (.A(_05117_));
 sg13g2_antennanp ANTENNA_84 (.A(_05117_));
 sg13g2_antennanp ANTENNA_85 (.A(_05131_));
 sg13g2_antennanp ANTENNA_86 (.A(_05131_));
 sg13g2_antennanp ANTENNA_87 (.A(_05131_));
 sg13g2_antennanp ANTENNA_88 (.A(_05131_));
 sg13g2_antennanp ANTENNA_89 (.A(_05131_));
 sg13g2_antennanp ANTENNA_90 (.A(_05131_));
 sg13g2_antennanp ANTENNA_91 (.A(_05131_));
 sg13g2_antennanp ANTENNA_92 (.A(_05131_));
 sg13g2_antennanp ANTENNA_93 (.A(_05131_));
 sg13g2_antennanp ANTENNA_94 (.A(_05131_));
 sg13g2_antennanp ANTENNA_95 (.A(_05131_));
 sg13g2_antennanp ANTENNA_96 (.A(_05131_));
 sg13g2_antennanp ANTENNA_97 (.A(_05179_));
 sg13g2_antennanp ANTENNA_98 (.A(_05179_));
 sg13g2_antennanp ANTENNA_99 (.A(_05179_));
 sg13g2_antennanp ANTENNA_100 (.A(_05179_));
 sg13g2_antennanp ANTENNA_101 (.A(_05179_));
 sg13g2_antennanp ANTENNA_102 (.A(_05179_));
 sg13g2_antennanp ANTENNA_103 (.A(_05179_));
 sg13g2_antennanp ANTENNA_104 (.A(_05179_));
 sg13g2_antennanp ANTENNA_105 (.A(_05179_));
 sg13g2_antennanp ANTENNA_106 (.A(_05267_));
 sg13g2_antennanp ANTENNA_107 (.A(_05267_));
 sg13g2_antennanp ANTENNA_108 (.A(_05267_));
 sg13g2_antennanp ANTENNA_109 (.A(_05267_));
 sg13g2_antennanp ANTENNA_110 (.A(_05267_));
 sg13g2_antennanp ANTENNA_111 (.A(_05267_));
 sg13g2_antennanp ANTENNA_112 (.A(_05267_));
 sg13g2_antennanp ANTENNA_113 (.A(_05267_));
 sg13g2_antennanp ANTENNA_114 (.A(_05267_));
 sg13g2_antennanp ANTENNA_115 (.A(_05267_));
 sg13g2_antennanp ANTENNA_116 (.A(_05408_));
 sg13g2_antennanp ANTENNA_117 (.A(_05408_));
 sg13g2_antennanp ANTENNA_118 (.A(_05408_));
 sg13g2_antennanp ANTENNA_119 (.A(_05408_));
 sg13g2_antennanp ANTENNA_120 (.A(_05408_));
 sg13g2_antennanp ANTENNA_121 (.A(_05415_));
 sg13g2_antennanp ANTENNA_122 (.A(_05415_));
 sg13g2_antennanp ANTENNA_123 (.A(_05415_));
 sg13g2_antennanp ANTENNA_124 (.A(_05416_));
 sg13g2_antennanp ANTENNA_125 (.A(_05416_));
 sg13g2_antennanp ANTENNA_126 (.A(_05416_));
 sg13g2_antennanp ANTENNA_127 (.A(_05416_));
 sg13g2_antennanp ANTENNA_128 (.A(_05416_));
 sg13g2_antennanp ANTENNA_129 (.A(_05416_));
 sg13g2_antennanp ANTENNA_130 (.A(_05737_));
 sg13g2_antennanp ANTENNA_131 (.A(_05737_));
 sg13g2_antennanp ANTENNA_132 (.A(_05737_));
 sg13g2_antennanp ANTENNA_133 (.A(_05757_));
 sg13g2_antennanp ANTENNA_134 (.A(_05757_));
 sg13g2_antennanp ANTENNA_135 (.A(_05757_));
 sg13g2_antennanp ANTENNA_136 (.A(_05811_));
 sg13g2_antennanp ANTENNA_137 (.A(_05811_));
 sg13g2_antennanp ANTENNA_138 (.A(_05811_));
 sg13g2_antennanp ANTENNA_139 (.A(_05811_));
 sg13g2_antennanp ANTENNA_140 (.A(_05811_));
 sg13g2_antennanp ANTENNA_141 (.A(_05811_));
 sg13g2_antennanp ANTENNA_142 (.A(_05811_));
 sg13g2_antennanp ANTENNA_143 (.A(_05811_));
 sg13g2_antennanp ANTENNA_144 (.A(_05811_));
 sg13g2_antennanp ANTENNA_145 (.A(_05811_));
 sg13g2_antennanp ANTENNA_146 (.A(_05811_));
 sg13g2_antennanp ANTENNA_147 (.A(_05811_));
 sg13g2_antennanp ANTENNA_148 (.A(_05811_));
 sg13g2_antennanp ANTENNA_149 (.A(_06055_));
 sg13g2_antennanp ANTENNA_150 (.A(_06055_));
 sg13g2_antennanp ANTENNA_151 (.A(_06055_));
 sg13g2_antennanp ANTENNA_152 (.A(_06055_));
 sg13g2_antennanp ANTENNA_153 (.A(_06055_));
 sg13g2_antennanp ANTENNA_154 (.A(_06055_));
 sg13g2_antennanp ANTENNA_155 (.A(_06055_));
 sg13g2_antennanp ANTENNA_156 (.A(_06055_));
 sg13g2_antennanp ANTENNA_157 (.A(_06055_));
 sg13g2_antennanp ANTENNA_158 (.A(_06055_));
 sg13g2_antennanp ANTENNA_159 (.A(_06057_));
 sg13g2_antennanp ANTENNA_160 (.A(_06057_));
 sg13g2_antennanp ANTENNA_161 (.A(_06057_));
 sg13g2_antennanp ANTENNA_162 (.A(_06111_));
 sg13g2_antennanp ANTENNA_163 (.A(_06111_));
 sg13g2_antennanp ANTENNA_164 (.A(_06111_));
 sg13g2_antennanp ANTENNA_165 (.A(_06111_));
 sg13g2_antennanp ANTENNA_166 (.A(_06111_));
 sg13g2_antennanp ANTENNA_167 (.A(_06111_));
 sg13g2_antennanp ANTENNA_168 (.A(_06111_));
 sg13g2_antennanp ANTENNA_169 (.A(_06111_));
 sg13g2_antennanp ANTENNA_170 (.A(_06111_));
 sg13g2_antennanp ANTENNA_171 (.A(_06111_));
 sg13g2_antennanp ANTENNA_172 (.A(_06111_));
 sg13g2_antennanp ANTENNA_173 (.A(_06111_));
 sg13g2_antennanp ANTENNA_174 (.A(_06111_));
 sg13g2_antennanp ANTENNA_175 (.A(_06111_));
 sg13g2_antennanp ANTENNA_176 (.A(_06111_));
 sg13g2_antennanp ANTENNA_177 (.A(_06111_));
 sg13g2_antennanp ANTENNA_178 (.A(_06111_));
 sg13g2_antennanp ANTENNA_179 (.A(_06111_));
 sg13g2_antennanp ANTENNA_180 (.A(_06285_));
 sg13g2_antennanp ANTENNA_181 (.A(_06285_));
 sg13g2_antennanp ANTENNA_182 (.A(_06285_));
 sg13g2_antennanp ANTENNA_183 (.A(_06285_));
 sg13g2_antennanp ANTENNA_184 (.A(_06285_));
 sg13g2_antennanp ANTENNA_185 (.A(_06285_));
 sg13g2_antennanp ANTENNA_186 (.A(_06474_));
 sg13g2_antennanp ANTENNA_187 (.A(_06474_));
 sg13g2_antennanp ANTENNA_188 (.A(_06474_));
 sg13g2_antennanp ANTENNA_189 (.A(_06474_));
 sg13g2_antennanp ANTENNA_190 (.A(_06474_));
 sg13g2_antennanp ANTENNA_191 (.A(_06474_));
 sg13g2_antennanp ANTENNA_192 (.A(_06667_));
 sg13g2_antennanp ANTENNA_193 (.A(_06667_));
 sg13g2_antennanp ANTENNA_194 (.A(_06667_));
 sg13g2_antennanp ANTENNA_195 (.A(_06667_));
 sg13g2_antennanp ANTENNA_196 (.A(_06897_));
 sg13g2_antennanp ANTENNA_197 (.A(_06897_));
 sg13g2_antennanp ANTENNA_198 (.A(_06897_));
 sg13g2_antennanp ANTENNA_199 (.A(_06897_));
 sg13g2_antennanp ANTENNA_200 (.A(_06897_));
 sg13g2_antennanp ANTENNA_201 (.A(_06900_));
 sg13g2_antennanp ANTENNA_202 (.A(_06900_));
 sg13g2_antennanp ANTENNA_203 (.A(_06900_));
 sg13g2_antennanp ANTENNA_204 (.A(_07117_));
 sg13g2_antennanp ANTENNA_205 (.A(_07117_));
 sg13g2_antennanp ANTENNA_206 (.A(_07117_));
 sg13g2_antennanp ANTENNA_207 (.A(_07117_));
 sg13g2_antennanp ANTENNA_208 (.A(_07194_));
 sg13g2_antennanp ANTENNA_209 (.A(_07194_));
 sg13g2_antennanp ANTENNA_210 (.A(_07194_));
 sg13g2_antennanp ANTENNA_211 (.A(_07561_));
 sg13g2_antennanp ANTENNA_212 (.A(_07561_));
 sg13g2_antennanp ANTENNA_213 (.A(_07561_));
 sg13g2_antennanp ANTENNA_214 (.A(_08349_));
 sg13g2_antennanp ANTENNA_215 (.A(_08349_));
 sg13g2_antennanp ANTENNA_216 (.A(_08349_));
 sg13g2_antennanp ANTENNA_217 (.A(_08349_));
 sg13g2_antennanp ANTENNA_218 (.A(_08349_));
 sg13g2_antennanp ANTENNA_219 (.A(_08349_));
 sg13g2_antennanp ANTENNA_220 (.A(_08737_));
 sg13g2_antennanp ANTENNA_221 (.A(_08737_));
 sg13g2_antennanp ANTENNA_222 (.A(_08737_));
 sg13g2_antennanp ANTENNA_223 (.A(_08737_));
 sg13g2_antennanp ANTENNA_224 (.A(_08737_));
 sg13g2_antennanp ANTENNA_225 (.A(_08737_));
 sg13g2_antennanp ANTENNA_226 (.A(_08737_));
 sg13g2_antennanp ANTENNA_227 (.A(_08737_));
 sg13g2_antennanp ANTENNA_228 (.A(_08737_));
 sg13g2_antennanp ANTENNA_229 (.A(_08737_));
 sg13g2_antennanp ANTENNA_230 (.A(_10237_));
 sg13g2_antennanp ANTENNA_231 (.A(_10237_));
 sg13g2_antennanp ANTENNA_232 (.A(_10237_));
 sg13g2_antennanp ANTENNA_233 (.A(_10237_));
 sg13g2_antennanp ANTENNA_234 (.A(_10237_));
 sg13g2_antennanp ANTENNA_235 (.A(_10237_));
 sg13g2_antennanp ANTENNA_236 (.A(_10237_));
 sg13g2_antennanp ANTENNA_237 (.A(_10237_));
 sg13g2_antennanp ANTENNA_238 (.A(_11347_));
 sg13g2_antennanp ANTENNA_239 (.A(_11347_));
 sg13g2_antennanp ANTENNA_240 (.A(_11347_));
 sg13g2_antennanp ANTENNA_241 (.A(_11347_));
 sg13g2_antennanp ANTENNA_242 (.A(_11347_));
 sg13g2_antennanp ANTENNA_243 (.A(_11347_));
 sg13g2_antennanp ANTENNA_244 (.A(_11347_));
 sg13g2_antennanp ANTENNA_245 (.A(_11347_));
 sg13g2_antennanp ANTENNA_246 (.A(_11347_));
 sg13g2_antennanp ANTENNA_247 (.A(_11347_));
 sg13g2_antennanp ANTENNA_248 (.A(_11347_));
 sg13g2_antennanp ANTENNA_249 (.A(_11347_));
 sg13g2_antennanp ANTENNA_250 (.A(_11347_));
 sg13g2_antennanp ANTENNA_251 (.A(_11347_));
 sg13g2_antennanp ANTENNA_252 (.A(_11347_));
 sg13g2_antennanp ANTENNA_253 (.A(_11347_));
 sg13g2_antennanp ANTENNA_254 (.A(_11347_));
 sg13g2_antennanp ANTENNA_255 (.A(_12651_));
 sg13g2_antennanp ANTENNA_256 (.A(_12651_));
 sg13g2_antennanp ANTENNA_257 (.A(_12651_));
 sg13g2_antennanp ANTENNA_258 (.A(_12651_));
 sg13g2_antennanp ANTENNA_259 (.A(_12651_));
 sg13g2_antennanp ANTENNA_260 (.A(_12651_));
 sg13g2_antennanp ANTENNA_261 (.A(_12651_));
 sg13g2_antennanp ANTENNA_262 (.A(_12651_));
 sg13g2_antennanp ANTENNA_263 (.A(_12651_));
 sg13g2_antennanp ANTENNA_264 (.A(_12967_));
 sg13g2_antennanp ANTENNA_265 (.A(_12967_));
 sg13g2_antennanp ANTENNA_266 (.A(_12967_));
 sg13g2_antennanp ANTENNA_267 (.A(_12999_));
 sg13g2_antennanp ANTENNA_268 (.A(_12999_));
 sg13g2_antennanp ANTENNA_269 (.A(_12999_));
 sg13g2_antennanp ANTENNA_270 (.A(_13104_));
 sg13g2_antennanp ANTENNA_271 (.A(_13104_));
 sg13g2_antennanp ANTENNA_272 (.A(_13104_));
 sg13g2_antennanp ANTENNA_273 (.A(_13104_));
 sg13g2_antennanp ANTENNA_274 (.A(_13127_));
 sg13g2_antennanp ANTENNA_275 (.A(_13127_));
 sg13g2_antennanp ANTENNA_276 (.A(_13127_));
 sg13g2_antennanp ANTENNA_277 (.A(net27));
 sg13g2_antennanp ANTENNA_278 (.A(net27));
 sg13g2_antennanp ANTENNA_279 (.A(net27));
 sg13g2_antennanp ANTENNA_280 (.A(net27));
 sg13g2_antennanp ANTENNA_281 (.A(net27));
 sg13g2_antennanp ANTENNA_282 (.A(net27));
 sg13g2_antennanp ANTENNA_283 (.A(net27));
 sg13g2_antennanp ANTENNA_284 (.A(net27));
 sg13g2_antennanp ANTENNA_285 (.A(net27));
 sg13g2_antennanp ANTENNA_286 (.A(net27));
 sg13g2_antennanp ANTENNA_287 (.A(net27));
 sg13g2_antennanp ANTENNA_288 (.A(net27));
 sg13g2_antennanp ANTENNA_289 (.A(net27));
 sg13g2_antennanp ANTENNA_290 (.A(net27));
 sg13g2_antennanp ANTENNA_291 (.A(net31));
 sg13g2_antennanp ANTENNA_292 (.A(net31));
 sg13g2_antennanp ANTENNA_293 (.A(net31));
 sg13g2_antennanp ANTENNA_294 (.A(net31));
 sg13g2_antennanp ANTENNA_295 (.A(net31));
 sg13g2_antennanp ANTENNA_296 (.A(net31));
 sg13g2_antennanp ANTENNA_297 (.A(net31));
 sg13g2_antennanp ANTENNA_298 (.A(net31));
 sg13g2_antennanp ANTENNA_299 (.A(net31));
 sg13g2_antennanp ANTENNA_300 (.A(net31));
 sg13g2_antennanp ANTENNA_301 (.A(net31));
 sg13g2_antennanp ANTENNA_302 (.A(net31));
 sg13g2_antennanp ANTENNA_303 (.A(net31));
 sg13g2_antennanp ANTENNA_304 (.A(net31));
 sg13g2_antennanp ANTENNA_305 (.A(net31));
 sg13g2_antennanp ANTENNA_306 (.A(net31));
 sg13g2_antennanp ANTENNA_307 (.A(net31));
 sg13g2_antennanp ANTENNA_308 (.A(net31));
 sg13g2_antennanp ANTENNA_309 (.A(net31));
 sg13g2_antennanp ANTENNA_310 (.A(net31));
 sg13g2_antennanp ANTENNA_311 (.A(net31));
 sg13g2_antennanp ANTENNA_312 (.A(net31));
 sg13g2_antennanp ANTENNA_313 (.A(net31));
 sg13g2_antennanp ANTENNA_314 (.A(net31));
 sg13g2_antennanp ANTENNA_315 (.A(net31));
 sg13g2_antennanp ANTENNA_316 (.A(net31));
 sg13g2_antennanp ANTENNA_317 (.A(net31));
 sg13g2_antennanp ANTENNA_318 (.A(net31));
 sg13g2_antennanp ANTENNA_319 (.A(net33));
 sg13g2_antennanp ANTENNA_320 (.A(net33));
 sg13g2_antennanp ANTENNA_321 (.A(net33));
 sg13g2_antennanp ANTENNA_322 (.A(net33));
 sg13g2_antennanp ANTENNA_323 (.A(net33));
 sg13g2_antennanp ANTENNA_324 (.A(net33));
 sg13g2_antennanp ANTENNA_325 (.A(net33));
 sg13g2_antennanp ANTENNA_326 (.A(net33));
 sg13g2_antennanp ANTENNA_327 (.A(net33));
 sg13g2_antennanp ANTENNA_328 (.A(net38));
 sg13g2_antennanp ANTENNA_329 (.A(net38));
 sg13g2_antennanp ANTENNA_330 (.A(net38));
 sg13g2_antennanp ANTENNA_331 (.A(net38));
 sg13g2_antennanp ANTENNA_332 (.A(net38));
 sg13g2_antennanp ANTENNA_333 (.A(net38));
 sg13g2_antennanp ANTENNA_334 (.A(net38));
 sg13g2_antennanp ANTENNA_335 (.A(net38));
 sg13g2_antennanp ANTENNA_336 (.A(net38));
 sg13g2_antennanp ANTENNA_337 (.A(net38));
 sg13g2_antennanp ANTENNA_338 (.A(net38));
 sg13g2_antennanp ANTENNA_339 (.A(net38));
 sg13g2_antennanp ANTENNA_340 (.A(net38));
 sg13g2_antennanp ANTENNA_341 (.A(net38));
 sg13g2_antennanp ANTENNA_342 (.A(net38));
 sg13g2_antennanp ANTENNA_343 (.A(net38));
 sg13g2_antennanp ANTENNA_344 (.A(net38));
 sg13g2_antennanp ANTENNA_345 (.A(net38));
 sg13g2_antennanp ANTENNA_346 (.A(net43));
 sg13g2_antennanp ANTENNA_347 (.A(net43));
 sg13g2_antennanp ANTENNA_348 (.A(net43));
 sg13g2_antennanp ANTENNA_349 (.A(net43));
 sg13g2_antennanp ANTENNA_350 (.A(net43));
 sg13g2_antennanp ANTENNA_351 (.A(net43));
 sg13g2_antennanp ANTENNA_352 (.A(net43));
 sg13g2_antennanp ANTENNA_353 (.A(net43));
 sg13g2_antennanp ANTENNA_354 (.A(net43));
 sg13g2_antennanp ANTENNA_355 (.A(net43));
 sg13g2_antennanp ANTENNA_356 (.A(net43));
 sg13g2_antennanp ANTENNA_357 (.A(net43));
 sg13g2_antennanp ANTENNA_358 (.A(net43));
 sg13g2_antennanp ANTENNA_359 (.A(net43));
 sg13g2_antennanp ANTENNA_360 (.A(net44));
 sg13g2_antennanp ANTENNA_361 (.A(net44));
 sg13g2_antennanp ANTENNA_362 (.A(net44));
 sg13g2_antennanp ANTENNA_363 (.A(net44));
 sg13g2_antennanp ANTENNA_364 (.A(net44));
 sg13g2_antennanp ANTENNA_365 (.A(net44));
 sg13g2_antennanp ANTENNA_366 (.A(net44));
 sg13g2_antennanp ANTENNA_367 (.A(net44));
 sg13g2_antennanp ANTENNA_368 (.A(net44));
 sg13g2_antennanp ANTENNA_369 (.A(net44));
 sg13g2_antennanp ANTENNA_370 (.A(net44));
 sg13g2_antennanp ANTENNA_371 (.A(net44));
 sg13g2_antennanp ANTENNA_372 (.A(net44));
 sg13g2_antennanp ANTENNA_373 (.A(net44));
 sg13g2_antennanp ANTENNA_374 (.A(net44));
 sg13g2_antennanp ANTENNA_375 (.A(net73));
 sg13g2_antennanp ANTENNA_376 (.A(net73));
 sg13g2_antennanp ANTENNA_377 (.A(net73));
 sg13g2_antennanp ANTENNA_378 (.A(net73));
 sg13g2_antennanp ANTENNA_379 (.A(net73));
 sg13g2_antennanp ANTENNA_380 (.A(net73));
 sg13g2_antennanp ANTENNA_381 (.A(net73));
 sg13g2_antennanp ANTENNA_382 (.A(net73));
 sg13g2_antennanp ANTENNA_383 (.A(net73));
 sg13g2_antennanp ANTENNA_384 (.A(net73));
 sg13g2_antennanp ANTENNA_385 (.A(net73));
 sg13g2_antennanp ANTENNA_386 (.A(net73));
 sg13g2_antennanp ANTENNA_387 (.A(net73));
 sg13g2_antennanp ANTENNA_388 (.A(net73));
 sg13g2_antennanp ANTENNA_389 (.A(net73));
 sg13g2_antennanp ANTENNA_390 (.A(net73));
 sg13g2_antennanp ANTENNA_391 (.A(net73));
 sg13g2_antennanp ANTENNA_392 (.A(net73));
 sg13g2_antennanp ANTENNA_393 (.A(net73));
 sg13g2_antennanp ANTENNA_394 (.A(net73));
 sg13g2_antennanp ANTENNA_395 (.A(net73));
 sg13g2_antennanp ANTENNA_396 (.A(net73));
 sg13g2_antennanp ANTENNA_397 (.A(net78));
 sg13g2_antennanp ANTENNA_398 (.A(net78));
 sg13g2_antennanp ANTENNA_399 (.A(net78));
 sg13g2_antennanp ANTENNA_400 (.A(net78));
 sg13g2_antennanp ANTENNA_401 (.A(net78));
 sg13g2_antennanp ANTENNA_402 (.A(net78));
 sg13g2_antennanp ANTENNA_403 (.A(net78));
 sg13g2_antennanp ANTENNA_404 (.A(net78));
 sg13g2_antennanp ANTENNA_405 (.A(net78));
 sg13g2_antennanp ANTENNA_406 (.A(net78));
 sg13g2_antennanp ANTENNA_407 (.A(net78));
 sg13g2_antennanp ANTENNA_408 (.A(net79));
 sg13g2_antennanp ANTENNA_409 (.A(net79));
 sg13g2_antennanp ANTENNA_410 (.A(net79));
 sg13g2_antennanp ANTENNA_411 (.A(net79));
 sg13g2_antennanp ANTENNA_412 (.A(net79));
 sg13g2_antennanp ANTENNA_413 (.A(net79));
 sg13g2_antennanp ANTENNA_414 (.A(net79));
 sg13g2_antennanp ANTENNA_415 (.A(net79));
 sg13g2_antennanp ANTENNA_416 (.A(net79));
 sg13g2_antennanp ANTENNA_417 (.A(net79));
 sg13g2_antennanp ANTENNA_418 (.A(net79));
 sg13g2_antennanp ANTENNA_419 (.A(net79));
 sg13g2_antennanp ANTENNA_420 (.A(net79));
 sg13g2_antennanp ANTENNA_421 (.A(net79));
 sg13g2_antennanp ANTENNA_422 (.A(net79));
 sg13g2_antennanp ANTENNA_423 (.A(net79));
 sg13g2_antennanp ANTENNA_424 (.A(net79));
 sg13g2_antennanp ANTENNA_425 (.A(net79));
 sg13g2_antennanp ANTENNA_426 (.A(net79));
 sg13g2_antennanp ANTENNA_427 (.A(net79));
 sg13g2_antennanp ANTENNA_428 (.A(net79));
 sg13g2_antennanp ANTENNA_429 (.A(net79));
 sg13g2_antennanp ANTENNA_430 (.A(net79));
 sg13g2_antennanp ANTENNA_431 (.A(net79));
 sg13g2_antennanp ANTENNA_432 (.A(net79));
 sg13g2_antennanp ANTENNA_433 (.A(net79));
 sg13g2_antennanp ANTENNA_434 (.A(net79));
 sg13g2_antennanp ANTENNA_435 (.A(net79));
 sg13g2_antennanp ANTENNA_436 (.A(net79));
 sg13g2_antennanp ANTENNA_437 (.A(net79));
 sg13g2_antennanp ANTENNA_438 (.A(net79));
 sg13g2_antennanp ANTENNA_439 (.A(net79));
 sg13g2_antennanp ANTENNA_440 (.A(net79));
 sg13g2_antennanp ANTENNA_441 (.A(net80));
 sg13g2_antennanp ANTENNA_442 (.A(net80));
 sg13g2_antennanp ANTENNA_443 (.A(net80));
 sg13g2_antennanp ANTENNA_444 (.A(net80));
 sg13g2_antennanp ANTENNA_445 (.A(net80));
 sg13g2_antennanp ANTENNA_446 (.A(net80));
 sg13g2_antennanp ANTENNA_447 (.A(net80));
 sg13g2_antennanp ANTENNA_448 (.A(net80));
 sg13g2_antennanp ANTENNA_449 (.A(net107));
 sg13g2_antennanp ANTENNA_450 (.A(net107));
 sg13g2_antennanp ANTENNA_451 (.A(net107));
 sg13g2_antennanp ANTENNA_452 (.A(net107));
 sg13g2_antennanp ANTENNA_453 (.A(net107));
 sg13g2_antennanp ANTENNA_454 (.A(net107));
 sg13g2_antennanp ANTENNA_455 (.A(net107));
 sg13g2_antennanp ANTENNA_456 (.A(net107));
 sg13g2_antennanp ANTENNA_457 (.A(net108));
 sg13g2_antennanp ANTENNA_458 (.A(net108));
 sg13g2_antennanp ANTENNA_459 (.A(net108));
 sg13g2_antennanp ANTENNA_460 (.A(net108));
 sg13g2_antennanp ANTENNA_461 (.A(net108));
 sg13g2_antennanp ANTENNA_462 (.A(net108));
 sg13g2_antennanp ANTENNA_463 (.A(net108));
 sg13g2_antennanp ANTENNA_464 (.A(net108));
 sg13g2_antennanp ANTENNA_465 (.A(net108));
 sg13g2_antennanp ANTENNA_466 (.A(net108));
 sg13g2_antennanp ANTENNA_467 (.A(net108));
 sg13g2_antennanp ANTENNA_468 (.A(net108));
 sg13g2_antennanp ANTENNA_469 (.A(net108));
 sg13g2_antennanp ANTENNA_470 (.A(net108));
 sg13g2_antennanp ANTENNA_471 (.A(net108));
 sg13g2_antennanp ANTENNA_472 (.A(net108));
 sg13g2_antennanp ANTENNA_473 (.A(net108));
 sg13g2_antennanp ANTENNA_474 (.A(net108));
 sg13g2_antennanp ANTENNA_475 (.A(net108));
 sg13g2_antennanp ANTENNA_476 (.A(net108));
 sg13g2_antennanp ANTENNA_477 (.A(net108));
 sg13g2_antennanp ANTENNA_478 (.A(net108));
 sg13g2_antennanp ANTENNA_479 (.A(net108));
 sg13g2_antennanp ANTENNA_480 (.A(net108));
 sg13g2_antennanp ANTENNA_481 (.A(net108));
 sg13g2_antennanp ANTENNA_482 (.A(net108));
 sg13g2_antennanp ANTENNA_483 (.A(net108));
 sg13g2_antennanp ANTENNA_484 (.A(net108));
 sg13g2_antennanp ANTENNA_485 (.A(net108));
 sg13g2_antennanp ANTENNA_486 (.A(net108));
 sg13g2_antennanp ANTENNA_487 (.A(net108));
 sg13g2_antennanp ANTENNA_488 (.A(net108));
 sg13g2_antennanp ANTENNA_489 (.A(net108));
 sg13g2_antennanp ANTENNA_490 (.A(net108));
 sg13g2_antennanp ANTENNA_491 (.A(net108));
 sg13g2_antennanp ANTENNA_492 (.A(net108));
 sg13g2_antennanp ANTENNA_493 (.A(net113));
 sg13g2_antennanp ANTENNA_494 (.A(net113));
 sg13g2_antennanp ANTENNA_495 (.A(net113));
 sg13g2_antennanp ANTENNA_496 (.A(net113));
 sg13g2_antennanp ANTENNA_497 (.A(net113));
 sg13g2_antennanp ANTENNA_498 (.A(net113));
 sg13g2_antennanp ANTENNA_499 (.A(net113));
 sg13g2_antennanp ANTENNA_500 (.A(net113));
 sg13g2_antennanp ANTENNA_501 (.A(net113));
 sg13g2_antennanp ANTENNA_502 (.A(net113));
 sg13g2_antennanp ANTENNA_503 (.A(net113));
 sg13g2_antennanp ANTENNA_504 (.A(net113));
 sg13g2_antennanp ANTENNA_505 (.A(net113));
 sg13g2_antennanp ANTENNA_506 (.A(net113));
 sg13g2_antennanp ANTENNA_507 (.A(net118));
 sg13g2_antennanp ANTENNA_508 (.A(net118));
 sg13g2_antennanp ANTENNA_509 (.A(net118));
 sg13g2_antennanp ANTENNA_510 (.A(net118));
 sg13g2_antennanp ANTENNA_511 (.A(net118));
 sg13g2_antennanp ANTENNA_512 (.A(net118));
 sg13g2_antennanp ANTENNA_513 (.A(net118));
 sg13g2_antennanp ANTENNA_514 (.A(net118));
 sg13g2_antennanp ANTENNA_515 (.A(net118));
 sg13g2_antennanp ANTENNA_516 (.A(net118));
 sg13g2_antennanp ANTENNA_517 (.A(net118));
 sg13g2_antennanp ANTENNA_518 (.A(net118));
 sg13g2_antennanp ANTENNA_519 (.A(net118));
 sg13g2_antennanp ANTENNA_520 (.A(net119));
 sg13g2_antennanp ANTENNA_521 (.A(net119));
 sg13g2_antennanp ANTENNA_522 (.A(net119));
 sg13g2_antennanp ANTENNA_523 (.A(net119));
 sg13g2_antennanp ANTENNA_524 (.A(net119));
 sg13g2_antennanp ANTENNA_525 (.A(net119));
 sg13g2_antennanp ANTENNA_526 (.A(net119));
 sg13g2_antennanp ANTENNA_527 (.A(net119));
 sg13g2_antennanp ANTENNA_528 (.A(net119));
 sg13g2_antennanp ANTENNA_529 (.A(net119));
 sg13g2_antennanp ANTENNA_530 (.A(net119));
 sg13g2_antennanp ANTENNA_531 (.A(net119));
 sg13g2_antennanp ANTENNA_532 (.A(net119));
 sg13g2_antennanp ANTENNA_533 (.A(net119));
 sg13g2_antennanp ANTENNA_534 (.A(net119));
 sg13g2_antennanp ANTENNA_535 (.A(net124));
 sg13g2_antennanp ANTENNA_536 (.A(net124));
 sg13g2_antennanp ANTENNA_537 (.A(net124));
 sg13g2_antennanp ANTENNA_538 (.A(net124));
 sg13g2_antennanp ANTENNA_539 (.A(net124));
 sg13g2_antennanp ANTENNA_540 (.A(net124));
 sg13g2_antennanp ANTENNA_541 (.A(net124));
 sg13g2_antennanp ANTENNA_542 (.A(net124));
 sg13g2_antennanp ANTENNA_543 (.A(net124));
 sg13g2_antennanp ANTENNA_544 (.A(net124));
 sg13g2_antennanp ANTENNA_545 (.A(net124));
 sg13g2_antennanp ANTENNA_546 (.A(net124));
 sg13g2_antennanp ANTENNA_547 (.A(net125));
 sg13g2_antennanp ANTENNA_548 (.A(net125));
 sg13g2_antennanp ANTENNA_549 (.A(net125));
 sg13g2_antennanp ANTENNA_550 (.A(net125));
 sg13g2_antennanp ANTENNA_551 (.A(net125));
 sg13g2_antennanp ANTENNA_552 (.A(net125));
 sg13g2_antennanp ANTENNA_553 (.A(net125));
 sg13g2_antennanp ANTENNA_554 (.A(net125));
 sg13g2_antennanp ANTENNA_555 (.A(net126));
 sg13g2_antennanp ANTENNA_556 (.A(net126));
 sg13g2_antennanp ANTENNA_557 (.A(net126));
 sg13g2_antennanp ANTENNA_558 (.A(net126));
 sg13g2_antennanp ANTENNA_559 (.A(net126));
 sg13g2_antennanp ANTENNA_560 (.A(net126));
 sg13g2_antennanp ANTENNA_561 (.A(net126));
 sg13g2_antennanp ANTENNA_562 (.A(net126));
 sg13g2_antennanp ANTENNA_563 (.A(net126));
 sg13g2_antennanp ANTENNA_564 (.A(net126));
 sg13g2_antennanp ANTENNA_565 (.A(net126));
 sg13g2_antennanp ANTENNA_566 (.A(net126));
 sg13g2_antennanp ANTENNA_567 (.A(net126));
 sg13g2_antennanp ANTENNA_568 (.A(net126));
 sg13g2_antennanp ANTENNA_569 (.A(net126));
 sg13g2_antennanp ANTENNA_570 (.A(net127));
 sg13g2_antennanp ANTENNA_571 (.A(net127));
 sg13g2_antennanp ANTENNA_572 (.A(net127));
 sg13g2_antennanp ANTENNA_573 (.A(net127));
 sg13g2_antennanp ANTENNA_574 (.A(net127));
 sg13g2_antennanp ANTENNA_575 (.A(net127));
 sg13g2_antennanp ANTENNA_576 (.A(net127));
 sg13g2_antennanp ANTENNA_577 (.A(net127));
 sg13g2_antennanp ANTENNA_578 (.A(net127));
 sg13g2_antennanp ANTENNA_579 (.A(net127));
 sg13g2_antennanp ANTENNA_580 (.A(net127));
 sg13g2_antennanp ANTENNA_581 (.A(net127));
 sg13g2_antennanp ANTENNA_582 (.A(net127));
 sg13g2_antennanp ANTENNA_583 (.A(net127));
 sg13g2_antennanp ANTENNA_584 (.A(net127));
 sg13g2_antennanp ANTENNA_585 (.A(net127));
 sg13g2_antennanp ANTENNA_586 (.A(net127));
 sg13g2_antennanp ANTENNA_587 (.A(net127));
 sg13g2_antennanp ANTENNA_588 (.A(net127));
 sg13g2_antennanp ANTENNA_589 (.A(net127));
 sg13g2_antennanp ANTENNA_590 (.A(net127));
 sg13g2_antennanp ANTENNA_591 (.A(net127));
 sg13g2_antennanp ANTENNA_592 (.A(net166));
 sg13g2_antennanp ANTENNA_593 (.A(net166));
 sg13g2_antennanp ANTENNA_594 (.A(net166));
 sg13g2_antennanp ANTENNA_595 (.A(net166));
 sg13g2_antennanp ANTENNA_596 (.A(net166));
 sg13g2_antennanp ANTENNA_597 (.A(net166));
 sg13g2_antennanp ANTENNA_598 (.A(net166));
 sg13g2_antennanp ANTENNA_599 (.A(net166));
 sg13g2_antennanp ANTENNA_600 (.A(net166));
 sg13g2_antennanp ANTENNA_601 (.A(net166));
 sg13g2_antennanp ANTENNA_602 (.A(net166));
 sg13g2_antennanp ANTENNA_603 (.A(net166));
 sg13g2_antennanp ANTENNA_604 (.A(net166));
 sg13g2_antennanp ANTENNA_605 (.A(net166));
 sg13g2_antennanp ANTENNA_606 (.A(net166));
 sg13g2_antennanp ANTENNA_607 (.A(net166));
 sg13g2_antennanp ANTENNA_608 (.A(net166));
 sg13g2_antennanp ANTENNA_609 (.A(net166));
 sg13g2_antennanp ANTENNA_610 (.A(net166));
 sg13g2_antennanp ANTENNA_611 (.A(net166));
 sg13g2_antennanp ANTENNA_612 (.A(net166));
 sg13g2_antennanp ANTENNA_613 (.A(net166));
 sg13g2_antennanp ANTENNA_614 (.A(net167));
 sg13g2_antennanp ANTENNA_615 (.A(net167));
 sg13g2_antennanp ANTENNA_616 (.A(net167));
 sg13g2_antennanp ANTENNA_617 (.A(net167));
 sg13g2_antennanp ANTENNA_618 (.A(net167));
 sg13g2_antennanp ANTENNA_619 (.A(net167));
 sg13g2_antennanp ANTENNA_620 (.A(net167));
 sg13g2_antennanp ANTENNA_621 (.A(net167));
 sg13g2_antennanp ANTENNA_622 (.A(net167));
 sg13g2_antennanp ANTENNA_623 (.A(net167));
 sg13g2_antennanp ANTENNA_624 (.A(net170));
 sg13g2_antennanp ANTENNA_625 (.A(net170));
 sg13g2_antennanp ANTENNA_626 (.A(net170));
 sg13g2_antennanp ANTENNA_627 (.A(net170));
 sg13g2_antennanp ANTENNA_628 (.A(net170));
 sg13g2_antennanp ANTENNA_629 (.A(net170));
 sg13g2_antennanp ANTENNA_630 (.A(net170));
 sg13g2_antennanp ANTENNA_631 (.A(net170));
 sg13g2_antennanp ANTENNA_632 (.A(net170));
 sg13g2_antennanp ANTENNA_633 (.A(net170));
 sg13g2_antennanp ANTENNA_634 (.A(net170));
 sg13g2_antennanp ANTENNA_635 (.A(net170));
 sg13g2_antennanp ANTENNA_636 (.A(net170));
 sg13g2_antennanp ANTENNA_637 (.A(net170));
 sg13g2_antennanp ANTENNA_638 (.A(net170));
 sg13g2_antennanp ANTENNA_639 (.A(net176));
 sg13g2_antennanp ANTENNA_640 (.A(net176));
 sg13g2_antennanp ANTENNA_641 (.A(net176));
 sg13g2_antennanp ANTENNA_642 (.A(net176));
 sg13g2_antennanp ANTENNA_643 (.A(net176));
 sg13g2_antennanp ANTENNA_644 (.A(net176));
 sg13g2_antennanp ANTENNA_645 (.A(net176));
 sg13g2_antennanp ANTENNA_646 (.A(net176));
 sg13g2_antennanp ANTENNA_647 (.A(net176));
 sg13g2_antennanp ANTENNA_648 (.A(net176));
 sg13g2_antennanp ANTENNA_649 (.A(net176));
 sg13g2_antennanp ANTENNA_650 (.A(net176));
 sg13g2_antennanp ANTENNA_651 (.A(net176));
 sg13g2_antennanp ANTENNA_652 (.A(net176));
 sg13g2_antennanp ANTENNA_653 (.A(net176));
 sg13g2_antennanp ANTENNA_654 (.A(net176));
 sg13g2_antennanp ANTENNA_655 (.A(net176));
 sg13g2_antennanp ANTENNA_656 (.A(net176));
 sg13g2_antennanp ANTENNA_657 (.A(net176));
 sg13g2_antennanp ANTENNA_658 (.A(net176));
 sg13g2_antennanp ANTENNA_659 (.A(net176));
 sg13g2_antennanp ANTENNA_660 (.A(net317));
 sg13g2_antennanp ANTENNA_661 (.A(net317));
 sg13g2_antennanp ANTENNA_662 (.A(net317));
 sg13g2_antennanp ANTENNA_663 (.A(net317));
 sg13g2_antennanp ANTENNA_664 (.A(net317));
 sg13g2_antennanp ANTENNA_665 (.A(net317));
 sg13g2_antennanp ANTENNA_666 (.A(net317));
 sg13g2_antennanp ANTENNA_667 (.A(net317));
 sg13g2_antennanp ANTENNA_668 (.A(net327));
 sg13g2_antennanp ANTENNA_669 (.A(net327));
 sg13g2_antennanp ANTENNA_670 (.A(net327));
 sg13g2_antennanp ANTENNA_671 (.A(net327));
 sg13g2_antennanp ANTENNA_672 (.A(net327));
 sg13g2_antennanp ANTENNA_673 (.A(net327));
 sg13g2_antennanp ANTENNA_674 (.A(net327));
 sg13g2_antennanp ANTENNA_675 (.A(net327));
 sg13g2_antennanp ANTENNA_676 (.A(net327));
 sg13g2_antennanp ANTENNA_677 (.A(net327));
 sg13g2_antennanp ANTENNA_678 (.A(net327));
 sg13g2_antennanp ANTENNA_679 (.A(net327));
 sg13g2_antennanp ANTENNA_680 (.A(net368));
 sg13g2_antennanp ANTENNA_681 (.A(net368));
 sg13g2_antennanp ANTENNA_682 (.A(net368));
 sg13g2_antennanp ANTENNA_683 (.A(net368));
 sg13g2_antennanp ANTENNA_684 (.A(net368));
 sg13g2_antennanp ANTENNA_685 (.A(net368));
 sg13g2_antennanp ANTENNA_686 (.A(net368));
 sg13g2_antennanp ANTENNA_687 (.A(net368));
 sg13g2_antennanp ANTENNA_688 (.A(net368));
 sg13g2_antennanp ANTENNA_689 (.A(net368));
 sg13g2_antennanp ANTENNA_690 (.A(net368));
 sg13g2_antennanp ANTENNA_691 (.A(net368));
 sg13g2_antennanp ANTENNA_692 (.A(net368));
 sg13g2_antennanp ANTENNA_693 (.A(net368));
 sg13g2_antennanp ANTENNA_694 (.A(net368));
 sg13g2_antennanp ANTENNA_695 (.A(net368));
 sg13g2_antennanp ANTENNA_696 (.A(net386));
 sg13g2_antennanp ANTENNA_697 (.A(net386));
 sg13g2_antennanp ANTENNA_698 (.A(net386));
 sg13g2_antennanp ANTENNA_699 (.A(net386));
 sg13g2_antennanp ANTENNA_700 (.A(net386));
 sg13g2_antennanp ANTENNA_701 (.A(net386));
 sg13g2_antennanp ANTENNA_702 (.A(net386));
 sg13g2_antennanp ANTENNA_703 (.A(net386));
 sg13g2_antennanp ANTENNA_704 (.A(net386));
 sg13g2_antennanp ANTENNA_705 (.A(net386));
 sg13g2_antennanp ANTENNA_706 (.A(net386));
 sg13g2_antennanp ANTENNA_707 (.A(net386));
 sg13g2_antennanp ANTENNA_708 (.A(net386));
 sg13g2_antennanp ANTENNA_709 (.A(net386));
 sg13g2_antennanp ANTENNA_710 (.A(net386));
 sg13g2_antennanp ANTENNA_711 (.A(net386));
 sg13g2_antennanp ANTENNA_712 (.A(net386));
 sg13g2_antennanp ANTENNA_713 (.A(net435));
 sg13g2_antennanp ANTENNA_714 (.A(net435));
 sg13g2_antennanp ANTENNA_715 (.A(net435));
 sg13g2_antennanp ANTENNA_716 (.A(net435));
 sg13g2_antennanp ANTENNA_717 (.A(net435));
 sg13g2_antennanp ANTENNA_718 (.A(net435));
 sg13g2_antennanp ANTENNA_719 (.A(net435));
 sg13g2_antennanp ANTENNA_720 (.A(net435));
 sg13g2_antennanp ANTENNA_721 (.A(net435));
 sg13g2_antennanp ANTENNA_722 (.A(net435));
 sg13g2_antennanp ANTENNA_723 (.A(net435));
 sg13g2_antennanp ANTENNA_724 (.A(net435));
 sg13g2_antennanp ANTENNA_725 (.A(net435));
 sg13g2_antennanp ANTENNA_726 (.A(net435));
 sg13g2_antennanp ANTENNA_727 (.A(net435));
 sg13g2_antennanp ANTENNA_728 (.A(net435));
 sg13g2_antennanp ANTENNA_729 (.A(net435));
 sg13g2_antennanp ANTENNA_730 (.A(net435));
 sg13g2_antennanp ANTENNA_731 (.A(net435));
 sg13g2_antennanp ANTENNA_732 (.A(net714));
 sg13g2_antennanp ANTENNA_733 (.A(net714));
 sg13g2_antennanp ANTENNA_734 (.A(net714));
 sg13g2_antennanp ANTENNA_735 (.A(net714));
 sg13g2_antennanp ANTENNA_736 (.A(net714));
 sg13g2_antennanp ANTENNA_737 (.A(net714));
 sg13g2_antennanp ANTENNA_738 (.A(net714));
 sg13g2_antennanp ANTENNA_739 (.A(net714));
 sg13g2_antennanp ANTENNA_740 (.A(net714));
 sg13g2_antennanp ANTENNA_741 (.A(net714));
 sg13g2_antennanp ANTENNA_742 (.A(net714));
 sg13g2_antennanp ANTENNA_743 (.A(net714));
 sg13g2_antennanp ANTENNA_744 (.A(net714));
 sg13g2_antennanp ANTENNA_745 (.A(net714));
 sg13g2_antennanp ANTENNA_746 (.A(net714));
 sg13g2_antennanp ANTENNA_747 (.A(net715));
 sg13g2_antennanp ANTENNA_748 (.A(net715));
 sg13g2_antennanp ANTENNA_749 (.A(net715));
 sg13g2_antennanp ANTENNA_750 (.A(net715));
 sg13g2_antennanp ANTENNA_751 (.A(net715));
 sg13g2_antennanp ANTENNA_752 (.A(net715));
 sg13g2_antennanp ANTENNA_753 (.A(net715));
 sg13g2_antennanp ANTENNA_754 (.A(net715));
 sg13g2_antennanp ANTENNA_755 (.A(net715));
 sg13g2_antennanp ANTENNA_756 (.A(net715));
 sg13g2_antennanp ANTENNA_757 (.A(net715));
 sg13g2_antennanp ANTENNA_758 (.A(net715));
 sg13g2_antennanp ANTENNA_759 (.A(net715));
 sg13g2_antennanp ANTENNA_760 (.A(net715));
 sg13g2_antennanp ANTENNA_761 (.A(net715));
 sg13g2_antennanp ANTENNA_762 (.A(net715));
 sg13g2_antennanp ANTENNA_763 (.A(net716));
 sg13g2_antennanp ANTENNA_764 (.A(net716));
 sg13g2_antennanp ANTENNA_765 (.A(net716));
 sg13g2_antennanp ANTENNA_766 (.A(net716));
 sg13g2_antennanp ANTENNA_767 (.A(net716));
 sg13g2_antennanp ANTENNA_768 (.A(net716));
 sg13g2_antennanp ANTENNA_769 (.A(net716));
 sg13g2_antennanp ANTENNA_770 (.A(net716));
 sg13g2_antennanp ANTENNA_771 (.A(net716));
 sg13g2_antennanp ANTENNA_772 (.A(net716));
 sg13g2_antennanp ANTENNA_773 (.A(net716));
 sg13g2_antennanp ANTENNA_774 (.A(net716));
 sg13g2_antennanp ANTENNA_775 (.A(net716));
 sg13g2_antennanp ANTENNA_776 (.A(net716));
 sg13g2_antennanp ANTENNA_777 (.A(net1054));
 sg13g2_antennanp ANTENNA_778 (.A(net1054));
 sg13g2_antennanp ANTENNA_779 (.A(net1054));
 sg13g2_antennanp ANTENNA_780 (.A(net1054));
 sg13g2_antennanp ANTENNA_781 (.A(net1054));
 sg13g2_antennanp ANTENNA_782 (.A(net1054));
 sg13g2_antennanp ANTENNA_783 (.A(net1054));
 sg13g2_antennanp ANTENNA_784 (.A(net1054));
 sg13g2_antennanp ANTENNA_785 (.A(net1054));
 sg13g2_antennanp ANTENNA_786 (.A(net1054));
 sg13g2_antennanp ANTENNA_787 (.A(net1054));
 sg13g2_antennanp ANTENNA_788 (.A(_00461_));
 sg13g2_antennanp ANTENNA_789 (.A(_00534_));
 sg13g2_antennanp ANTENNA_790 (.A(_00534_));
 sg13g2_antennanp ANTENNA_791 (.A(_00788_));
 sg13g2_antennanp ANTENNA_792 (.A(_00788_));
 sg13g2_antennanp ANTENNA_793 (.A(_00788_));
 sg13g2_antennanp ANTENNA_794 (.A(_01440_));
 sg13g2_antennanp ANTENNA_795 (.A(_01440_));
 sg13g2_antennanp ANTENNA_796 (.A(_01795_));
 sg13g2_antennanp ANTENNA_797 (.A(_01795_));
 sg13g2_antennanp ANTENNA_798 (.A(_02787_));
 sg13g2_antennanp ANTENNA_799 (.A(_02787_));
 sg13g2_antennanp ANTENNA_800 (.A(_02787_));
 sg13g2_antennanp ANTENNA_801 (.A(_02787_));
 sg13g2_antennanp ANTENNA_802 (.A(_02787_));
 sg13g2_antennanp ANTENNA_803 (.A(_02787_));
 sg13g2_antennanp ANTENNA_804 (.A(_03810_));
 sg13g2_antennanp ANTENNA_805 (.A(_03810_));
 sg13g2_antennanp ANTENNA_806 (.A(_03810_));
 sg13g2_antennanp ANTENNA_807 (.A(_03810_));
 sg13g2_antennanp ANTENNA_808 (.A(_03821_));
 sg13g2_antennanp ANTENNA_809 (.A(_03821_));
 sg13g2_antennanp ANTENNA_810 (.A(_03821_));
 sg13g2_antennanp ANTENNA_811 (.A(_03821_));
 sg13g2_antennanp ANTENNA_812 (.A(_04067_));
 sg13g2_antennanp ANTENNA_813 (.A(_04067_));
 sg13g2_antennanp ANTENNA_814 (.A(_04067_));
 sg13g2_antennanp ANTENNA_815 (.A(_04067_));
 sg13g2_antennanp ANTENNA_816 (.A(_04067_));
 sg13g2_antennanp ANTENNA_817 (.A(_04067_));
 sg13g2_antennanp ANTENNA_818 (.A(_04067_));
 sg13g2_antennanp ANTENNA_819 (.A(_04067_));
 sg13g2_antennanp ANTENNA_820 (.A(_04077_));
 sg13g2_antennanp ANTENNA_821 (.A(_04077_));
 sg13g2_antennanp ANTENNA_822 (.A(_04077_));
 sg13g2_antennanp ANTENNA_823 (.A(_04077_));
 sg13g2_antennanp ANTENNA_824 (.A(_04077_));
 sg13g2_antennanp ANTENNA_825 (.A(_04077_));
 sg13g2_antennanp ANTENNA_826 (.A(_04242_));
 sg13g2_antennanp ANTENNA_827 (.A(_04242_));
 sg13g2_antennanp ANTENNA_828 (.A(_04371_));
 sg13g2_antennanp ANTENNA_829 (.A(_04378_));
 sg13g2_antennanp ANTENNA_830 (.A(_04393_));
 sg13g2_antennanp ANTENNA_831 (.A(_04403_));
 sg13g2_antennanp ANTENNA_832 (.A(_04411_));
 sg13g2_antennanp ANTENNA_833 (.A(_04412_));
 sg13g2_antennanp ANTENNA_834 (.A(_04416_));
 sg13g2_antennanp ANTENNA_835 (.A(_04419_));
 sg13g2_antennanp ANTENNA_836 (.A(_04432_));
 sg13g2_antennanp ANTENNA_837 (.A(_04453_));
 sg13g2_antennanp ANTENNA_838 (.A(_04475_));
 sg13g2_antennanp ANTENNA_839 (.A(_04481_));
 sg13g2_antennanp ANTENNA_840 (.A(_04481_));
 sg13g2_antennanp ANTENNA_841 (.A(_04508_));
 sg13g2_antennanp ANTENNA_842 (.A(_04756_));
 sg13g2_antennanp ANTENNA_843 (.A(_04773_));
 sg13g2_antennanp ANTENNA_844 (.A(_04804_));
 sg13g2_antennanp ANTENNA_845 (.A(_04816_));
 sg13g2_antennanp ANTENNA_846 (.A(_04817_));
 sg13g2_antennanp ANTENNA_847 (.A(_04828_));
 sg13g2_antennanp ANTENNA_848 (.A(_04838_));
 sg13g2_antennanp ANTENNA_849 (.A(_04840_));
 sg13g2_antennanp ANTENNA_850 (.A(_04842_));
 sg13g2_antennanp ANTENNA_851 (.A(_04850_));
 sg13g2_antennanp ANTENNA_852 (.A(_04853_));
 sg13g2_antennanp ANTENNA_853 (.A(_04860_));
 sg13g2_antennanp ANTENNA_854 (.A(_04860_));
 sg13g2_antennanp ANTENNA_855 (.A(_04860_));
 sg13g2_antennanp ANTENNA_856 (.A(_04914_));
 sg13g2_antennanp ANTENNA_857 (.A(_04914_));
 sg13g2_antennanp ANTENNA_858 (.A(_04941_));
 sg13g2_antennanp ANTENNA_859 (.A(_04941_));
 sg13g2_antennanp ANTENNA_860 (.A(_04941_));
 sg13g2_antennanp ANTENNA_861 (.A(_04941_));
 sg13g2_antennanp ANTENNA_862 (.A(_04941_));
 sg13g2_antennanp ANTENNA_863 (.A(_04941_));
 sg13g2_antennanp ANTENNA_864 (.A(_04941_));
 sg13g2_antennanp ANTENNA_865 (.A(_04941_));
 sg13g2_antennanp ANTENNA_866 (.A(_05117_));
 sg13g2_antennanp ANTENNA_867 (.A(_05131_));
 sg13g2_antennanp ANTENNA_868 (.A(_05131_));
 sg13g2_antennanp ANTENNA_869 (.A(_05131_));
 sg13g2_antennanp ANTENNA_870 (.A(_05131_));
 sg13g2_antennanp ANTENNA_871 (.A(_05131_));
 sg13g2_antennanp ANTENNA_872 (.A(_05131_));
 sg13g2_antennanp ANTENNA_873 (.A(_05131_));
 sg13g2_antennanp ANTENNA_874 (.A(_05131_));
 sg13g2_antennanp ANTENNA_875 (.A(_05131_));
 sg13g2_antennanp ANTENNA_876 (.A(_05131_));
 sg13g2_antennanp ANTENNA_877 (.A(_05131_));
 sg13g2_antennanp ANTENNA_878 (.A(_05131_));
 sg13g2_antennanp ANTENNA_879 (.A(_05131_));
 sg13g2_antennanp ANTENNA_880 (.A(_05131_));
 sg13g2_antennanp ANTENNA_881 (.A(_05131_));
 sg13g2_antennanp ANTENNA_882 (.A(_05267_));
 sg13g2_antennanp ANTENNA_883 (.A(_05267_));
 sg13g2_antennanp ANTENNA_884 (.A(_05267_));
 sg13g2_antennanp ANTENNA_885 (.A(_05267_));
 sg13g2_antennanp ANTENNA_886 (.A(_05267_));
 sg13g2_antennanp ANTENNA_887 (.A(_05267_));
 sg13g2_antennanp ANTENNA_888 (.A(_05408_));
 sg13g2_antennanp ANTENNA_889 (.A(_05408_));
 sg13g2_antennanp ANTENNA_890 (.A(_05408_));
 sg13g2_antennanp ANTENNA_891 (.A(_05416_));
 sg13g2_antennanp ANTENNA_892 (.A(_05416_));
 sg13g2_antennanp ANTENNA_893 (.A(_05416_));
 sg13g2_antennanp ANTENNA_894 (.A(_05416_));
 sg13g2_antennanp ANTENNA_895 (.A(_05416_));
 sg13g2_antennanp ANTENNA_896 (.A(_05416_));
 sg13g2_antennanp ANTENNA_897 (.A(_05737_));
 sg13g2_antennanp ANTENNA_898 (.A(_05737_));
 sg13g2_antennanp ANTENNA_899 (.A(_05737_));
 sg13g2_antennanp ANTENNA_900 (.A(_05757_));
 sg13g2_antennanp ANTENNA_901 (.A(_05757_));
 sg13g2_antennanp ANTENNA_902 (.A(_05757_));
 sg13g2_antennanp ANTENNA_903 (.A(_05757_));
 sg13g2_antennanp ANTENNA_904 (.A(_05757_));
 sg13g2_antennanp ANTENNA_905 (.A(_05757_));
 sg13g2_antennanp ANTENNA_906 (.A(_05757_));
 sg13g2_antennanp ANTENNA_907 (.A(_05811_));
 sg13g2_antennanp ANTENNA_908 (.A(_05811_));
 sg13g2_antennanp ANTENNA_909 (.A(_05811_));
 sg13g2_antennanp ANTENNA_910 (.A(_05811_));
 sg13g2_antennanp ANTENNA_911 (.A(_05811_));
 sg13g2_antennanp ANTENNA_912 (.A(_05811_));
 sg13g2_antennanp ANTENNA_913 (.A(_05811_));
 sg13g2_antennanp ANTENNA_914 (.A(_06111_));
 sg13g2_antennanp ANTENNA_915 (.A(_06111_));
 sg13g2_antennanp ANTENNA_916 (.A(_06111_));
 sg13g2_antennanp ANTENNA_917 (.A(_06111_));
 sg13g2_antennanp ANTENNA_918 (.A(_06111_));
 sg13g2_antennanp ANTENNA_919 (.A(_06111_));
 sg13g2_antennanp ANTENNA_920 (.A(_06285_));
 sg13g2_antennanp ANTENNA_921 (.A(_06285_));
 sg13g2_antennanp ANTENNA_922 (.A(_06285_));
 sg13g2_antennanp ANTENNA_923 (.A(_06285_));
 sg13g2_antennanp ANTENNA_924 (.A(_06285_));
 sg13g2_antennanp ANTENNA_925 (.A(_06285_));
 sg13g2_antennanp ANTENNA_926 (.A(_06468_));
 sg13g2_antennanp ANTENNA_927 (.A(_06468_));
 sg13g2_antennanp ANTENNA_928 (.A(_06468_));
 sg13g2_antennanp ANTENNA_929 (.A(_06468_));
 sg13g2_antennanp ANTENNA_930 (.A(_06468_));
 sg13g2_antennanp ANTENNA_931 (.A(_06468_));
 sg13g2_antennanp ANTENNA_932 (.A(_06468_));
 sg13g2_antennanp ANTENNA_933 (.A(_06468_));
 sg13g2_antennanp ANTENNA_934 (.A(_06474_));
 sg13g2_antennanp ANTENNA_935 (.A(_06474_));
 sg13g2_antennanp ANTENNA_936 (.A(_06474_));
 sg13g2_antennanp ANTENNA_937 (.A(_06474_));
 sg13g2_antennanp ANTENNA_938 (.A(_06474_));
 sg13g2_antennanp ANTENNA_939 (.A(_06474_));
 sg13g2_antennanp ANTENNA_940 (.A(_06667_));
 sg13g2_antennanp ANTENNA_941 (.A(_06667_));
 sg13g2_antennanp ANTENNA_942 (.A(_06667_));
 sg13g2_antennanp ANTENNA_943 (.A(_06667_));
 sg13g2_antennanp ANTENNA_944 (.A(_06897_));
 sg13g2_antennanp ANTENNA_945 (.A(_06897_));
 sg13g2_antennanp ANTENNA_946 (.A(_06897_));
 sg13g2_antennanp ANTENNA_947 (.A(_06897_));
 sg13g2_antennanp ANTENNA_948 (.A(_06900_));
 sg13g2_antennanp ANTENNA_949 (.A(_06900_));
 sg13g2_antennanp ANTENNA_950 (.A(_06900_));
 sg13g2_antennanp ANTENNA_951 (.A(_06900_));
 sg13g2_antennanp ANTENNA_952 (.A(_06900_));
 sg13g2_antennanp ANTENNA_953 (.A(_06900_));
 sg13g2_antennanp ANTENNA_954 (.A(_06900_));
 sg13g2_antennanp ANTENNA_955 (.A(_06900_));
 sg13g2_antennanp ANTENNA_956 (.A(_06900_));
 sg13g2_antennanp ANTENNA_957 (.A(_06900_));
 sg13g2_antennanp ANTENNA_958 (.A(_07117_));
 sg13g2_antennanp ANTENNA_959 (.A(_07117_));
 sg13g2_antennanp ANTENNA_960 (.A(_07117_));
 sg13g2_antennanp ANTENNA_961 (.A(_07117_));
 sg13g2_antennanp ANTENNA_962 (.A(_08349_));
 sg13g2_antennanp ANTENNA_963 (.A(_08349_));
 sg13g2_antennanp ANTENNA_964 (.A(_08349_));
 sg13g2_antennanp ANTENNA_965 (.A(_08349_));
 sg13g2_antennanp ANTENNA_966 (.A(_08349_));
 sg13g2_antennanp ANTENNA_967 (.A(_08349_));
 sg13g2_antennanp ANTENNA_968 (.A(_08737_));
 sg13g2_antennanp ANTENNA_969 (.A(_08737_));
 sg13g2_antennanp ANTENNA_970 (.A(_08737_));
 sg13g2_antennanp ANTENNA_971 (.A(_10237_));
 sg13g2_antennanp ANTENNA_972 (.A(_10237_));
 sg13g2_antennanp ANTENNA_973 (.A(_10237_));
 sg13g2_antennanp ANTENNA_974 (.A(_10237_));
 sg13g2_antennanp ANTENNA_975 (.A(_10237_));
 sg13g2_antennanp ANTENNA_976 (.A(_10237_));
 sg13g2_antennanp ANTENNA_977 (.A(_10237_));
 sg13g2_antennanp ANTENNA_978 (.A(_10237_));
 sg13g2_antennanp ANTENNA_979 (.A(_10237_));
 sg13g2_antennanp ANTENNA_980 (.A(_12651_));
 sg13g2_antennanp ANTENNA_981 (.A(_12651_));
 sg13g2_antennanp ANTENNA_982 (.A(_12651_));
 sg13g2_antennanp ANTENNA_983 (.A(_12651_));
 sg13g2_antennanp ANTENNA_984 (.A(_12651_));
 sg13g2_antennanp ANTENNA_985 (.A(_12651_));
 sg13g2_antennanp ANTENNA_986 (.A(_12651_));
 sg13g2_antennanp ANTENNA_987 (.A(_12651_));
 sg13g2_antennanp ANTENNA_988 (.A(_12651_));
 sg13g2_antennanp ANTENNA_989 (.A(_12999_));
 sg13g2_antennanp ANTENNA_990 (.A(_12999_));
 sg13g2_antennanp ANTENNA_991 (.A(_12999_));
 sg13g2_antennanp ANTENNA_992 (.A(_12999_));
 sg13g2_antennanp ANTENNA_993 (.A(_12999_));
 sg13g2_antennanp ANTENNA_994 (.A(_12999_));
 sg13g2_antennanp ANTENNA_995 (.A(_13104_));
 sg13g2_antennanp ANTENNA_996 (.A(_13104_));
 sg13g2_antennanp ANTENNA_997 (.A(_13104_));
 sg13g2_antennanp ANTENNA_998 (.A(_13104_));
 sg13g2_antennanp ANTENNA_999 (.A(_13127_));
 sg13g2_antennanp ANTENNA_1000 (.A(_13127_));
 sg13g2_antennanp ANTENNA_1001 (.A(_13127_));
 sg13g2_antennanp ANTENNA_1002 (.A(net43));
 sg13g2_antennanp ANTENNA_1003 (.A(net43));
 sg13g2_antennanp ANTENNA_1004 (.A(net43));
 sg13g2_antennanp ANTENNA_1005 (.A(net43));
 sg13g2_antennanp ANTENNA_1006 (.A(net43));
 sg13g2_antennanp ANTENNA_1007 (.A(net43));
 sg13g2_antennanp ANTENNA_1008 (.A(net43));
 sg13g2_antennanp ANTENNA_1009 (.A(net43));
 sg13g2_antennanp ANTENNA_1010 (.A(net43));
 sg13g2_antennanp ANTENNA_1011 (.A(net43));
 sg13g2_antennanp ANTENNA_1012 (.A(net43));
 sg13g2_antennanp ANTENNA_1013 (.A(net43));
 sg13g2_antennanp ANTENNA_1014 (.A(net43));
 sg13g2_antennanp ANTENNA_1015 (.A(net43));
 sg13g2_antennanp ANTENNA_1016 (.A(net44));
 sg13g2_antennanp ANTENNA_1017 (.A(net44));
 sg13g2_antennanp ANTENNA_1018 (.A(net44));
 sg13g2_antennanp ANTENNA_1019 (.A(net44));
 sg13g2_antennanp ANTENNA_1020 (.A(net44));
 sg13g2_antennanp ANTENNA_1021 (.A(net44));
 sg13g2_antennanp ANTENNA_1022 (.A(net44));
 sg13g2_antennanp ANTENNA_1023 (.A(net44));
 sg13g2_antennanp ANTENNA_1024 (.A(net44));
 sg13g2_antennanp ANTENNA_1025 (.A(net44));
 sg13g2_antennanp ANTENNA_1026 (.A(net44));
 sg13g2_antennanp ANTENNA_1027 (.A(net44));
 sg13g2_antennanp ANTENNA_1028 (.A(net44));
 sg13g2_antennanp ANTENNA_1029 (.A(net44));
 sg13g2_antennanp ANTENNA_1030 (.A(net73));
 sg13g2_antennanp ANTENNA_1031 (.A(net73));
 sg13g2_antennanp ANTENNA_1032 (.A(net73));
 sg13g2_antennanp ANTENNA_1033 (.A(net73));
 sg13g2_antennanp ANTENNA_1034 (.A(net73));
 sg13g2_antennanp ANTENNA_1035 (.A(net73));
 sg13g2_antennanp ANTENNA_1036 (.A(net73));
 sg13g2_antennanp ANTENNA_1037 (.A(net73));
 sg13g2_antennanp ANTENNA_1038 (.A(net73));
 sg13g2_antennanp ANTENNA_1039 (.A(net78));
 sg13g2_antennanp ANTENNA_1040 (.A(net78));
 sg13g2_antennanp ANTENNA_1041 (.A(net78));
 sg13g2_antennanp ANTENNA_1042 (.A(net78));
 sg13g2_antennanp ANTENNA_1043 (.A(net78));
 sg13g2_antennanp ANTENNA_1044 (.A(net78));
 sg13g2_antennanp ANTENNA_1045 (.A(net78));
 sg13g2_antennanp ANTENNA_1046 (.A(net78));
 sg13g2_antennanp ANTENNA_1047 (.A(net78));
 sg13g2_antennanp ANTENNA_1048 (.A(net78));
 sg13g2_antennanp ANTENNA_1049 (.A(net78));
 sg13g2_antennanp ANTENNA_1050 (.A(net78));
 sg13g2_antennanp ANTENNA_1051 (.A(net78));
 sg13g2_antennanp ANTENNA_1052 (.A(net78));
 sg13g2_antennanp ANTENNA_1053 (.A(net78));
 sg13g2_antennanp ANTENNA_1054 (.A(net78));
 sg13g2_antennanp ANTENNA_1055 (.A(net78));
 sg13g2_antennanp ANTENNA_1056 (.A(net78));
 sg13g2_antennanp ANTENNA_1057 (.A(net78));
 sg13g2_antennanp ANTENNA_1058 (.A(net78));
 sg13g2_antennanp ANTENNA_1059 (.A(net78));
 sg13g2_antennanp ANTENNA_1060 (.A(net78));
 sg13g2_antennanp ANTENNA_1061 (.A(net79));
 sg13g2_antennanp ANTENNA_1062 (.A(net79));
 sg13g2_antennanp ANTENNA_1063 (.A(net79));
 sg13g2_antennanp ANTENNA_1064 (.A(net79));
 sg13g2_antennanp ANTENNA_1065 (.A(net79));
 sg13g2_antennanp ANTENNA_1066 (.A(net79));
 sg13g2_antennanp ANTENNA_1067 (.A(net79));
 sg13g2_antennanp ANTENNA_1068 (.A(net79));
 sg13g2_antennanp ANTENNA_1069 (.A(net79));
 sg13g2_antennanp ANTENNA_1070 (.A(net79));
 sg13g2_antennanp ANTENNA_1071 (.A(net79));
 sg13g2_antennanp ANTENNA_1072 (.A(net79));
 sg13g2_antennanp ANTENNA_1073 (.A(net79));
 sg13g2_antennanp ANTENNA_1074 (.A(net79));
 sg13g2_antennanp ANTENNA_1075 (.A(net79));
 sg13g2_antennanp ANTENNA_1076 (.A(net79));
 sg13g2_antennanp ANTENNA_1077 (.A(net79));
 sg13g2_antennanp ANTENNA_1078 (.A(net79));
 sg13g2_antennanp ANTENNA_1079 (.A(net79));
 sg13g2_antennanp ANTENNA_1080 (.A(net79));
 sg13g2_antennanp ANTENNA_1081 (.A(net79));
 sg13g2_antennanp ANTENNA_1082 (.A(net79));
 sg13g2_antennanp ANTENNA_1083 (.A(net79));
 sg13g2_antennanp ANTENNA_1084 (.A(net79));
 sg13g2_antennanp ANTENNA_1085 (.A(net79));
 sg13g2_antennanp ANTENNA_1086 (.A(net79));
 sg13g2_antennanp ANTENNA_1087 (.A(net79));
 sg13g2_antennanp ANTENNA_1088 (.A(net79));
 sg13g2_antennanp ANTENNA_1089 (.A(net79));
 sg13g2_antennanp ANTENNA_1090 (.A(net79));
 sg13g2_antennanp ANTENNA_1091 (.A(net79));
 sg13g2_antennanp ANTENNA_1092 (.A(net79));
 sg13g2_antennanp ANTENNA_1093 (.A(net79));
 sg13g2_antennanp ANTENNA_1094 (.A(net79));
 sg13g2_antennanp ANTENNA_1095 (.A(net79));
 sg13g2_antennanp ANTENNA_1096 (.A(net79));
 sg13g2_antennanp ANTENNA_1097 (.A(net103));
 sg13g2_antennanp ANTENNA_1098 (.A(net103));
 sg13g2_antennanp ANTENNA_1099 (.A(net103));
 sg13g2_antennanp ANTENNA_1100 (.A(net103));
 sg13g2_antennanp ANTENNA_1101 (.A(net103));
 sg13g2_antennanp ANTENNA_1102 (.A(net103));
 sg13g2_antennanp ANTENNA_1103 (.A(net103));
 sg13g2_antennanp ANTENNA_1104 (.A(net103));
 sg13g2_antennanp ANTENNA_1105 (.A(net107));
 sg13g2_antennanp ANTENNA_1106 (.A(net107));
 sg13g2_antennanp ANTENNA_1107 (.A(net107));
 sg13g2_antennanp ANTENNA_1108 (.A(net107));
 sg13g2_antennanp ANTENNA_1109 (.A(net107));
 sg13g2_antennanp ANTENNA_1110 (.A(net107));
 sg13g2_antennanp ANTENNA_1111 (.A(net107));
 sg13g2_antennanp ANTENNA_1112 (.A(net107));
 sg13g2_antennanp ANTENNA_1113 (.A(net107));
 sg13g2_antennanp ANTENNA_1114 (.A(net107));
 sg13g2_antennanp ANTENNA_1115 (.A(net107));
 sg13g2_antennanp ANTENNA_1116 (.A(net107));
 sg13g2_antennanp ANTENNA_1117 (.A(net107));
 sg13g2_antennanp ANTENNA_1118 (.A(net107));
 sg13g2_antennanp ANTENNA_1119 (.A(net107));
 sg13g2_antennanp ANTENNA_1120 (.A(net107));
 sg13g2_antennanp ANTENNA_1121 (.A(net107));
 sg13g2_antennanp ANTENNA_1122 (.A(net107));
 sg13g2_antennanp ANTENNA_1123 (.A(net107));
 sg13g2_antennanp ANTENNA_1124 (.A(net107));
 sg13g2_antennanp ANTENNA_1125 (.A(net107));
 sg13g2_antennanp ANTENNA_1126 (.A(net107));
 sg13g2_antennanp ANTENNA_1127 (.A(net107));
 sg13g2_antennanp ANTENNA_1128 (.A(net107));
 sg13g2_antennanp ANTENNA_1129 (.A(net107));
 sg13g2_antennanp ANTENNA_1130 (.A(net107));
 sg13g2_antennanp ANTENNA_1131 (.A(net107));
 sg13g2_antennanp ANTENNA_1132 (.A(net113));
 sg13g2_antennanp ANTENNA_1133 (.A(net113));
 sg13g2_antennanp ANTENNA_1134 (.A(net113));
 sg13g2_antennanp ANTENNA_1135 (.A(net113));
 sg13g2_antennanp ANTENNA_1136 (.A(net113));
 sg13g2_antennanp ANTENNA_1137 (.A(net113));
 sg13g2_antennanp ANTENNA_1138 (.A(net113));
 sg13g2_antennanp ANTENNA_1139 (.A(net113));
 sg13g2_antennanp ANTENNA_1140 (.A(net113));
 sg13g2_antennanp ANTENNA_1141 (.A(net113));
 sg13g2_antennanp ANTENNA_1142 (.A(net113));
 sg13g2_antennanp ANTENNA_1143 (.A(net113));
 sg13g2_antennanp ANTENNA_1144 (.A(net113));
 sg13g2_antennanp ANTENNA_1145 (.A(net113));
 sg13g2_antennanp ANTENNA_1146 (.A(net113));
 sg13g2_antennanp ANTENNA_1147 (.A(net116));
 sg13g2_antennanp ANTENNA_1148 (.A(net116));
 sg13g2_antennanp ANTENNA_1149 (.A(net116));
 sg13g2_antennanp ANTENNA_1150 (.A(net116));
 sg13g2_antennanp ANTENNA_1151 (.A(net116));
 sg13g2_antennanp ANTENNA_1152 (.A(net116));
 sg13g2_antennanp ANTENNA_1153 (.A(net116));
 sg13g2_antennanp ANTENNA_1154 (.A(net116));
 sg13g2_antennanp ANTENNA_1155 (.A(net118));
 sg13g2_antennanp ANTENNA_1156 (.A(net118));
 sg13g2_antennanp ANTENNA_1157 (.A(net118));
 sg13g2_antennanp ANTENNA_1158 (.A(net118));
 sg13g2_antennanp ANTENNA_1159 (.A(net118));
 sg13g2_antennanp ANTENNA_1160 (.A(net118));
 sg13g2_antennanp ANTENNA_1161 (.A(net118));
 sg13g2_antennanp ANTENNA_1162 (.A(net118));
 sg13g2_antennanp ANTENNA_1163 (.A(net118));
 sg13g2_antennanp ANTENNA_1164 (.A(net118));
 sg13g2_antennanp ANTENNA_1165 (.A(net118));
 sg13g2_antennanp ANTENNA_1166 (.A(net118));
 sg13g2_antennanp ANTENNA_1167 (.A(net118));
 sg13g2_antennanp ANTENNA_1168 (.A(net118));
 sg13g2_antennanp ANTENNA_1169 (.A(net118));
 sg13g2_antennanp ANTENNA_1170 (.A(net118));
 sg13g2_antennanp ANTENNA_1171 (.A(net118));
 sg13g2_antennanp ANTENNA_1172 (.A(net118));
 sg13g2_antennanp ANTENNA_1173 (.A(net118));
 sg13g2_antennanp ANTENNA_1174 (.A(net118));
 sg13g2_antennanp ANTENNA_1175 (.A(net118));
 sg13g2_antennanp ANTENNA_1176 (.A(net118));
 sg13g2_antennanp ANTENNA_1177 (.A(net124));
 sg13g2_antennanp ANTENNA_1178 (.A(net124));
 sg13g2_antennanp ANTENNA_1179 (.A(net124));
 sg13g2_antennanp ANTENNA_1180 (.A(net124));
 sg13g2_antennanp ANTENNA_1181 (.A(net124));
 sg13g2_antennanp ANTENNA_1182 (.A(net124));
 sg13g2_antennanp ANTENNA_1183 (.A(net124));
 sg13g2_antennanp ANTENNA_1184 (.A(net124));
 sg13g2_antennanp ANTENNA_1185 (.A(net124));
 sg13g2_antennanp ANTENNA_1186 (.A(net124));
 sg13g2_antennanp ANTENNA_1187 (.A(net124));
 sg13g2_antennanp ANTENNA_1188 (.A(net124));
 sg13g2_antennanp ANTENNA_1189 (.A(net124));
 sg13g2_antennanp ANTENNA_1190 (.A(net125));
 sg13g2_antennanp ANTENNA_1191 (.A(net125));
 sg13g2_antennanp ANTENNA_1192 (.A(net125));
 sg13g2_antennanp ANTENNA_1193 (.A(net125));
 sg13g2_antennanp ANTENNA_1194 (.A(net125));
 sg13g2_antennanp ANTENNA_1195 (.A(net125));
 sg13g2_antennanp ANTENNA_1196 (.A(net125));
 sg13g2_antennanp ANTENNA_1197 (.A(net125));
 sg13g2_antennanp ANTENNA_1198 (.A(net125));
 sg13g2_antennanp ANTENNA_1199 (.A(net125));
 sg13g2_antennanp ANTENNA_1200 (.A(net125));
 sg13g2_antennanp ANTENNA_1201 (.A(net125));
 sg13g2_antennanp ANTENNA_1202 (.A(net125));
 sg13g2_antennanp ANTENNA_1203 (.A(net125));
 sg13g2_antennanp ANTENNA_1204 (.A(net125));
 sg13g2_antennanp ANTENNA_1205 (.A(net125));
 sg13g2_antennanp ANTENNA_1206 (.A(net125));
 sg13g2_antennanp ANTENNA_1207 (.A(net125));
 sg13g2_antennanp ANTENNA_1208 (.A(net125));
 sg13g2_antennanp ANTENNA_1209 (.A(net127));
 sg13g2_antennanp ANTENNA_1210 (.A(net127));
 sg13g2_antennanp ANTENNA_1211 (.A(net127));
 sg13g2_antennanp ANTENNA_1212 (.A(net127));
 sg13g2_antennanp ANTENNA_1213 (.A(net127));
 sg13g2_antennanp ANTENNA_1214 (.A(net127));
 sg13g2_antennanp ANTENNA_1215 (.A(net127));
 sg13g2_antennanp ANTENNA_1216 (.A(net127));
 sg13g2_antennanp ANTENNA_1217 (.A(net127));
 sg13g2_antennanp ANTENNA_1218 (.A(net127));
 sg13g2_antennanp ANTENNA_1219 (.A(net127));
 sg13g2_antennanp ANTENNA_1220 (.A(net127));
 sg13g2_antennanp ANTENNA_1221 (.A(net127));
 sg13g2_antennanp ANTENNA_1222 (.A(net127));
 sg13g2_antennanp ANTENNA_1223 (.A(net127));
 sg13g2_antennanp ANTENNA_1224 (.A(net127));
 sg13g2_antennanp ANTENNA_1225 (.A(net127));
 sg13g2_antennanp ANTENNA_1226 (.A(net127));
 sg13g2_antennanp ANTENNA_1227 (.A(net127));
 sg13g2_antennanp ANTENNA_1228 (.A(net127));
 sg13g2_antennanp ANTENNA_1229 (.A(net127));
 sg13g2_antennanp ANTENNA_1230 (.A(net127));
 sg13g2_antennanp ANTENNA_1231 (.A(net127));
 sg13g2_antennanp ANTENNA_1232 (.A(net127));
 sg13g2_antennanp ANTENNA_1233 (.A(net127));
 sg13g2_antennanp ANTENNA_1234 (.A(net127));
 sg13g2_antennanp ANTENNA_1235 (.A(net127));
 sg13g2_antennanp ANTENNA_1236 (.A(net127));
 sg13g2_antennanp ANTENNA_1237 (.A(net127));
 sg13g2_antennanp ANTENNA_1238 (.A(net127));
 sg13g2_antennanp ANTENNA_1239 (.A(net127));
 sg13g2_antennanp ANTENNA_1240 (.A(net127));
 sg13g2_antennanp ANTENNA_1241 (.A(net127));
 sg13g2_antennanp ANTENNA_1242 (.A(net127));
 sg13g2_antennanp ANTENNA_1243 (.A(net127));
 sg13g2_antennanp ANTENNA_1244 (.A(net127));
 sg13g2_antennanp ANTENNA_1245 (.A(net127));
 sg13g2_antennanp ANTENNA_1246 (.A(net127));
 sg13g2_antennanp ANTENNA_1247 (.A(net127));
 sg13g2_antennanp ANTENNA_1248 (.A(net127));
 sg13g2_antennanp ANTENNA_1249 (.A(net127));
 sg13g2_antennanp ANTENNA_1250 (.A(net127));
 sg13g2_antennanp ANTENNA_1251 (.A(net127));
 sg13g2_antennanp ANTENNA_1252 (.A(net127));
 sg13g2_antennanp ANTENNA_1253 (.A(net127));
 sg13g2_antennanp ANTENNA_1254 (.A(net166));
 sg13g2_antennanp ANTENNA_1255 (.A(net166));
 sg13g2_antennanp ANTENNA_1256 (.A(net166));
 sg13g2_antennanp ANTENNA_1257 (.A(net166));
 sg13g2_antennanp ANTENNA_1258 (.A(net166));
 sg13g2_antennanp ANTENNA_1259 (.A(net166));
 sg13g2_antennanp ANTENNA_1260 (.A(net166));
 sg13g2_antennanp ANTENNA_1261 (.A(net166));
 sg13g2_antennanp ANTENNA_1262 (.A(net166));
 sg13g2_antennanp ANTENNA_1263 (.A(net166));
 sg13g2_antennanp ANTENNA_1264 (.A(net166));
 sg13g2_antennanp ANTENNA_1265 (.A(net166));
 sg13g2_antennanp ANTENNA_1266 (.A(net166));
 sg13g2_antennanp ANTENNA_1267 (.A(net166));
 sg13g2_antennanp ANTENNA_1268 (.A(net166));
 sg13g2_antennanp ANTENNA_1269 (.A(net170));
 sg13g2_antennanp ANTENNA_1270 (.A(net170));
 sg13g2_antennanp ANTENNA_1271 (.A(net170));
 sg13g2_antennanp ANTENNA_1272 (.A(net170));
 sg13g2_antennanp ANTENNA_1273 (.A(net170));
 sg13g2_antennanp ANTENNA_1274 (.A(net170));
 sg13g2_antennanp ANTENNA_1275 (.A(net170));
 sg13g2_antennanp ANTENNA_1276 (.A(net170));
 sg13g2_antennanp ANTENNA_1277 (.A(net368));
 sg13g2_antennanp ANTENNA_1278 (.A(net368));
 sg13g2_antennanp ANTENNA_1279 (.A(net368));
 sg13g2_antennanp ANTENNA_1280 (.A(net368));
 sg13g2_antennanp ANTENNA_1281 (.A(net368));
 sg13g2_antennanp ANTENNA_1282 (.A(net368));
 sg13g2_antennanp ANTENNA_1283 (.A(net368));
 sg13g2_antennanp ANTENNA_1284 (.A(net368));
 sg13g2_antennanp ANTENNA_1285 (.A(net368));
 sg13g2_antennanp ANTENNA_1286 (.A(net368));
 sg13g2_antennanp ANTENNA_1287 (.A(net368));
 sg13g2_antennanp ANTENNA_1288 (.A(net368));
 sg13g2_antennanp ANTENNA_1289 (.A(net368));
 sg13g2_antennanp ANTENNA_1290 (.A(net368));
 sg13g2_antennanp ANTENNA_1291 (.A(net368));
 sg13g2_antennanp ANTENNA_1292 (.A(net368));
 sg13g2_antennanp ANTENNA_1293 (.A(net368));
 sg13g2_antennanp ANTENNA_1294 (.A(net368));
 sg13g2_antennanp ANTENNA_1295 (.A(net368));
 sg13g2_antennanp ANTENNA_1296 (.A(net368));
 sg13g2_antennanp ANTENNA_1297 (.A(net368));
 sg13g2_antennanp ANTENNA_1298 (.A(net368));
 sg13g2_antennanp ANTENNA_1299 (.A(net368));
 sg13g2_antennanp ANTENNA_1300 (.A(net368));
 sg13g2_antennanp ANTENNA_1301 (.A(net368));
 sg13g2_antennanp ANTENNA_1302 (.A(net368));
 sg13g2_antennanp ANTENNA_1303 (.A(net368));
 sg13g2_antennanp ANTENNA_1304 (.A(net368));
 sg13g2_antennanp ANTENNA_1305 (.A(net368));
 sg13g2_antennanp ANTENNA_1306 (.A(net368));
 sg13g2_antennanp ANTENNA_1307 (.A(net368));
 sg13g2_antennanp ANTENNA_1308 (.A(net368));
 sg13g2_antennanp ANTENNA_1309 (.A(net368));
 sg13g2_antennanp ANTENNA_1310 (.A(net368));
 sg13g2_antennanp ANTENNA_1311 (.A(net368));
 sg13g2_antennanp ANTENNA_1312 (.A(net368));
 sg13g2_antennanp ANTENNA_1313 (.A(net368));
 sg13g2_antennanp ANTENNA_1314 (.A(net368));
 sg13g2_antennanp ANTENNA_1315 (.A(net368));
 sg13g2_antennanp ANTENNA_1316 (.A(net368));
 sg13g2_antennanp ANTENNA_1317 (.A(net368));
 sg13g2_antennanp ANTENNA_1318 (.A(net368));
 sg13g2_antennanp ANTENNA_1319 (.A(net386));
 sg13g2_antennanp ANTENNA_1320 (.A(net386));
 sg13g2_antennanp ANTENNA_1321 (.A(net386));
 sg13g2_antennanp ANTENNA_1322 (.A(net386));
 sg13g2_antennanp ANTENNA_1323 (.A(net386));
 sg13g2_antennanp ANTENNA_1324 (.A(net386));
 sg13g2_antennanp ANTENNA_1325 (.A(net386));
 sg13g2_antennanp ANTENNA_1326 (.A(net386));
 sg13g2_antennanp ANTENNA_1327 (.A(net386));
 sg13g2_antennanp ANTENNA_1328 (.A(net386));
 sg13g2_antennanp ANTENNA_1329 (.A(net386));
 sg13g2_antennanp ANTENNA_1330 (.A(net386));
 sg13g2_antennanp ANTENNA_1331 (.A(net386));
 sg13g2_antennanp ANTENNA_1332 (.A(net386));
 sg13g2_antennanp ANTENNA_1333 (.A(net386));
 sg13g2_antennanp ANTENNA_1334 (.A(net386));
 sg13g2_antennanp ANTENNA_1335 (.A(net386));
 sg13g2_antennanp ANTENNA_1336 (.A(net716));
 sg13g2_antennanp ANTENNA_1337 (.A(net716));
 sg13g2_antennanp ANTENNA_1338 (.A(net716));
 sg13g2_antennanp ANTENNA_1339 (.A(net716));
 sg13g2_antennanp ANTENNA_1340 (.A(net716));
 sg13g2_antennanp ANTENNA_1341 (.A(net716));
 sg13g2_antennanp ANTENNA_1342 (.A(net716));
 sg13g2_antennanp ANTENNA_1343 (.A(net716));
 sg13g2_antennanp ANTENNA_1344 (.A(net1002));
 sg13g2_antennanp ANTENNA_1345 (.A(net1002));
 sg13g2_antennanp ANTENNA_1346 (.A(net1002));
 sg13g2_antennanp ANTENNA_1347 (.A(net1002));
 sg13g2_antennanp ANTENNA_1348 (.A(net1002));
 sg13g2_antennanp ANTENNA_1349 (.A(net1002));
 sg13g2_antennanp ANTENNA_1350 (.A(net1002));
 sg13g2_antennanp ANTENNA_1351 (.A(net1002));
 sg13g2_antennanp ANTENNA_1352 (.A(net1002));
 sg13g2_antennanp ANTENNA_1353 (.A(net1002));
 sg13g2_antennanp ANTENNA_1354 (.A(net1002));
 sg13g2_antennanp ANTENNA_1355 (.A(net1002));
 sg13g2_antennanp ANTENNA_1356 (.A(net1002));
 sg13g2_antennanp ANTENNA_1357 (.A(net1002));
 sg13g2_antennanp ANTENNA_1358 (.A(net1002));
 sg13g2_antennanp ANTENNA_1359 (.A(net1002));
 sg13g2_antennanp ANTENNA_1360 (.A(_00461_));
 sg13g2_antennanp ANTENNA_1361 (.A(_00534_));
 sg13g2_antennanp ANTENNA_1362 (.A(_00534_));
 sg13g2_antennanp ANTENNA_1363 (.A(_00788_));
 sg13g2_antennanp ANTENNA_1364 (.A(_00788_));
 sg13g2_antennanp ANTENNA_1365 (.A(_00788_));
 sg13g2_antennanp ANTENNA_1366 (.A(_01440_));
 sg13g2_antennanp ANTENNA_1367 (.A(_01440_));
 sg13g2_antennanp ANTENNA_1368 (.A(_01795_));
 sg13g2_antennanp ANTENNA_1369 (.A(_01795_));
 sg13g2_antennanp ANTENNA_1370 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1371 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1372 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1373 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1374 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1375 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1376 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1377 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1378 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1379 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1380 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1381 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1382 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1383 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1384 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1385 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1386 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1387 (.A(_03821_));
 sg13g2_antennanp ANTENNA_1388 (.A(_03821_));
 sg13g2_antennanp ANTENNA_1389 (.A(_03821_));
 sg13g2_antennanp ANTENNA_1390 (.A(_03821_));
 sg13g2_antennanp ANTENNA_1391 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1392 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1393 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1394 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1395 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1396 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1397 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1398 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1399 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1400 (.A(_04077_));
 sg13g2_antennanp ANTENNA_1401 (.A(_04077_));
 sg13g2_antennanp ANTENNA_1402 (.A(_04077_));
 sg13g2_antennanp ANTENNA_1403 (.A(_04242_));
 sg13g2_antennanp ANTENNA_1404 (.A(_04242_));
 sg13g2_antennanp ANTENNA_1405 (.A(_04371_));
 sg13g2_antennanp ANTENNA_1406 (.A(_04378_));
 sg13g2_antennanp ANTENNA_1407 (.A(_04393_));
 sg13g2_antennanp ANTENNA_1408 (.A(_04403_));
 sg13g2_antennanp ANTENNA_1409 (.A(_04411_));
 sg13g2_antennanp ANTENNA_1410 (.A(_04412_));
 sg13g2_antennanp ANTENNA_1411 (.A(_04416_));
 sg13g2_antennanp ANTENNA_1412 (.A(_04419_));
 sg13g2_antennanp ANTENNA_1413 (.A(_04432_));
 sg13g2_antennanp ANTENNA_1414 (.A(_04453_));
 sg13g2_antennanp ANTENNA_1415 (.A(_04481_));
 sg13g2_antennanp ANTENNA_1416 (.A(_04508_));
 sg13g2_antennanp ANTENNA_1417 (.A(_04756_));
 sg13g2_antennanp ANTENNA_1418 (.A(_04773_));
 sg13g2_antennanp ANTENNA_1419 (.A(_04804_));
 sg13g2_antennanp ANTENNA_1420 (.A(_04816_));
 sg13g2_antennanp ANTENNA_1421 (.A(_04817_));
 sg13g2_antennanp ANTENNA_1422 (.A(_04828_));
 sg13g2_antennanp ANTENNA_1423 (.A(_04838_));
 sg13g2_antennanp ANTENNA_1424 (.A(_04840_));
 sg13g2_antennanp ANTENNA_1425 (.A(_04842_));
 sg13g2_antennanp ANTENNA_1426 (.A(_04850_));
 sg13g2_antennanp ANTENNA_1427 (.A(_04853_));
 sg13g2_antennanp ANTENNA_1428 (.A(_04860_));
 sg13g2_antennanp ANTENNA_1429 (.A(_04860_));
 sg13g2_antennanp ANTENNA_1430 (.A(_04860_));
 sg13g2_antennanp ANTENNA_1431 (.A(_04914_));
 sg13g2_antennanp ANTENNA_1432 (.A(_04914_));
 sg13g2_antennanp ANTENNA_1433 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1434 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1435 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1436 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1437 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1438 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1439 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1440 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1441 (.A(_05117_));
 sg13g2_antennanp ANTENNA_1442 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1443 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1444 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1445 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1446 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1447 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1448 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1449 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1450 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1451 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1452 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1453 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1454 (.A(_05416_));
 sg13g2_antennanp ANTENNA_1455 (.A(_05416_));
 sg13g2_antennanp ANTENNA_1456 (.A(_05416_));
 sg13g2_antennanp ANTENNA_1457 (.A(_05737_));
 sg13g2_antennanp ANTENNA_1458 (.A(_05737_));
 sg13g2_antennanp ANTENNA_1459 (.A(_05737_));
 sg13g2_antennanp ANTENNA_1460 (.A(_05757_));
 sg13g2_antennanp ANTENNA_1461 (.A(_05757_));
 sg13g2_antennanp ANTENNA_1462 (.A(_05757_));
 sg13g2_antennanp ANTENNA_1463 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1464 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1465 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1466 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1467 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1468 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1469 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1470 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1471 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1472 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1473 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1474 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1475 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1476 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1477 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1478 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1479 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1480 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1481 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1482 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1483 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1484 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1485 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1486 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1487 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1488 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1489 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1490 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1491 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1492 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1493 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1494 (.A(_06468_));
 sg13g2_antennanp ANTENNA_1495 (.A(_06474_));
 sg13g2_antennanp ANTENNA_1496 (.A(_06474_));
 sg13g2_antennanp ANTENNA_1497 (.A(_06474_));
 sg13g2_antennanp ANTENNA_1498 (.A(_06474_));
 sg13g2_antennanp ANTENNA_1499 (.A(_06474_));
 sg13g2_antennanp ANTENNA_1500 (.A(_06474_));
 sg13g2_antennanp ANTENNA_1501 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1502 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1503 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1504 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1505 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1506 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1507 (.A(_06897_));
 sg13g2_antennanp ANTENNA_1508 (.A(_06897_));
 sg13g2_antennanp ANTENNA_1509 (.A(_06897_));
 sg13g2_antennanp ANTENNA_1510 (.A(_06897_));
 sg13g2_antennanp ANTENNA_1511 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1512 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1513 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1514 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1515 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1516 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1517 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1518 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1519 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1520 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1521 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1522 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1523 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1524 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1525 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1526 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1527 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1528 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1529 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1530 (.A(_08737_));
 sg13g2_antennanp ANTENNA_1531 (.A(_08737_));
 sg13g2_antennanp ANTENNA_1532 (.A(_08737_));
 sg13g2_antennanp ANTENNA_1533 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1534 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1535 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1536 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1537 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1538 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1539 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1540 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1541 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1542 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1543 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1544 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1545 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1546 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1547 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1548 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1549 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1550 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1551 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1552 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1553 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1554 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1555 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1556 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1557 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1558 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1559 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1560 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1561 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1562 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1563 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1564 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1565 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1566 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1567 (.A(_13104_));
 sg13g2_antennanp ANTENNA_1568 (.A(_13104_));
 sg13g2_antennanp ANTENNA_1569 (.A(_13104_));
 sg13g2_antennanp ANTENNA_1570 (.A(_13104_));
 sg13g2_antennanp ANTENNA_1571 (.A(net31));
 sg13g2_antennanp ANTENNA_1572 (.A(net31));
 sg13g2_antennanp ANTENNA_1573 (.A(net31));
 sg13g2_antennanp ANTENNA_1574 (.A(net31));
 sg13g2_antennanp ANTENNA_1575 (.A(net31));
 sg13g2_antennanp ANTENNA_1576 (.A(net31));
 sg13g2_antennanp ANTENNA_1577 (.A(net31));
 sg13g2_antennanp ANTENNA_1578 (.A(net31));
 sg13g2_antennanp ANTENNA_1579 (.A(net31));
 sg13g2_antennanp ANTENNA_1580 (.A(net31));
 sg13g2_antennanp ANTENNA_1581 (.A(net31));
 sg13g2_antennanp ANTENNA_1582 (.A(net31));
 sg13g2_antennanp ANTENNA_1583 (.A(net31));
 sg13g2_antennanp ANTENNA_1584 (.A(net31));
 sg13g2_antennanp ANTENNA_1585 (.A(net43));
 sg13g2_antennanp ANTENNA_1586 (.A(net43));
 sg13g2_antennanp ANTENNA_1587 (.A(net43));
 sg13g2_antennanp ANTENNA_1588 (.A(net43));
 sg13g2_antennanp ANTENNA_1589 (.A(net43));
 sg13g2_antennanp ANTENNA_1590 (.A(net43));
 sg13g2_antennanp ANTENNA_1591 (.A(net43));
 sg13g2_antennanp ANTENNA_1592 (.A(net43));
 sg13g2_antennanp ANTENNA_1593 (.A(net43));
 sg13g2_antennanp ANTENNA_1594 (.A(net43));
 sg13g2_antennanp ANTENNA_1595 (.A(net43));
 sg13g2_antennanp ANTENNA_1596 (.A(net43));
 sg13g2_antennanp ANTENNA_1597 (.A(net43));
 sg13g2_antennanp ANTENNA_1598 (.A(net43));
 sg13g2_antennanp ANTENNA_1599 (.A(net44));
 sg13g2_antennanp ANTENNA_1600 (.A(net44));
 sg13g2_antennanp ANTENNA_1601 (.A(net44));
 sg13g2_antennanp ANTENNA_1602 (.A(net44));
 sg13g2_antennanp ANTENNA_1603 (.A(net44));
 sg13g2_antennanp ANTENNA_1604 (.A(net44));
 sg13g2_antennanp ANTENNA_1605 (.A(net44));
 sg13g2_antennanp ANTENNA_1606 (.A(net44));
 sg13g2_antennanp ANTENNA_1607 (.A(net44));
 sg13g2_antennanp ANTENNA_1608 (.A(net44));
 sg13g2_antennanp ANTENNA_1609 (.A(net44));
 sg13g2_antennanp ANTENNA_1610 (.A(net73));
 sg13g2_antennanp ANTENNA_1611 (.A(net73));
 sg13g2_antennanp ANTENNA_1612 (.A(net73));
 sg13g2_antennanp ANTENNA_1613 (.A(net73));
 sg13g2_antennanp ANTENNA_1614 (.A(net73));
 sg13g2_antennanp ANTENNA_1615 (.A(net73));
 sg13g2_antennanp ANTENNA_1616 (.A(net73));
 sg13g2_antennanp ANTENNA_1617 (.A(net73));
 sg13g2_antennanp ANTENNA_1618 (.A(net73));
 sg13g2_antennanp ANTENNA_1619 (.A(net75));
 sg13g2_antennanp ANTENNA_1620 (.A(net75));
 sg13g2_antennanp ANTENNA_1621 (.A(net75));
 sg13g2_antennanp ANTENNA_1622 (.A(net75));
 sg13g2_antennanp ANTENNA_1623 (.A(net75));
 sg13g2_antennanp ANTENNA_1624 (.A(net75));
 sg13g2_antennanp ANTENNA_1625 (.A(net75));
 sg13g2_antennanp ANTENNA_1626 (.A(net75));
 sg13g2_antennanp ANTENNA_1627 (.A(net75));
 sg13g2_antennanp ANTENNA_1628 (.A(net75));
 sg13g2_antennanp ANTENNA_1629 (.A(net75));
 sg13g2_antennanp ANTENNA_1630 (.A(net75));
 sg13g2_antennanp ANTENNA_1631 (.A(net75));
 sg13g2_antennanp ANTENNA_1632 (.A(net75));
 sg13g2_antennanp ANTENNA_1633 (.A(net75));
 sg13g2_antennanp ANTENNA_1634 (.A(net75));
 sg13g2_antennanp ANTENNA_1635 (.A(net75));
 sg13g2_antennanp ANTENNA_1636 (.A(net75));
 sg13g2_antennanp ANTENNA_1637 (.A(net75));
 sg13g2_antennanp ANTENNA_1638 (.A(net75));
 sg13g2_antennanp ANTENNA_1639 (.A(net75));
 sg13g2_antennanp ANTENNA_1640 (.A(net75));
 sg13g2_antennanp ANTENNA_1641 (.A(net79));
 sg13g2_antennanp ANTENNA_1642 (.A(net79));
 sg13g2_antennanp ANTENNA_1643 (.A(net79));
 sg13g2_antennanp ANTENNA_1644 (.A(net79));
 sg13g2_antennanp ANTENNA_1645 (.A(net79));
 sg13g2_antennanp ANTENNA_1646 (.A(net79));
 sg13g2_antennanp ANTENNA_1647 (.A(net79));
 sg13g2_antennanp ANTENNA_1648 (.A(net79));
 sg13g2_antennanp ANTENNA_1649 (.A(net80));
 sg13g2_antennanp ANTENNA_1650 (.A(net80));
 sg13g2_antennanp ANTENNA_1651 (.A(net80));
 sg13g2_antennanp ANTENNA_1652 (.A(net80));
 sg13g2_antennanp ANTENNA_1653 (.A(net80));
 sg13g2_antennanp ANTENNA_1654 (.A(net80));
 sg13g2_antennanp ANTENNA_1655 (.A(net80));
 sg13g2_antennanp ANTENNA_1656 (.A(net80));
 sg13g2_antennanp ANTENNA_1657 (.A(net80));
 sg13g2_antennanp ANTENNA_1658 (.A(net80));
 sg13g2_antennanp ANTENNA_1659 (.A(net80));
 sg13g2_antennanp ANTENNA_1660 (.A(net80));
 sg13g2_antennanp ANTENNA_1661 (.A(net80));
 sg13g2_antennanp ANTENNA_1662 (.A(net80));
 sg13g2_antennanp ANTENNA_1663 (.A(net82));
 sg13g2_antennanp ANTENNA_1664 (.A(net82));
 sg13g2_antennanp ANTENNA_1665 (.A(net82));
 sg13g2_antennanp ANTENNA_1666 (.A(net82));
 sg13g2_antennanp ANTENNA_1667 (.A(net82));
 sg13g2_antennanp ANTENNA_1668 (.A(net82));
 sg13g2_antennanp ANTENNA_1669 (.A(net82));
 sg13g2_antennanp ANTENNA_1670 (.A(net82));
 sg13g2_antennanp ANTENNA_1671 (.A(net107));
 sg13g2_antennanp ANTENNA_1672 (.A(net107));
 sg13g2_antennanp ANTENNA_1673 (.A(net107));
 sg13g2_antennanp ANTENNA_1674 (.A(net107));
 sg13g2_antennanp ANTENNA_1675 (.A(net107));
 sg13g2_antennanp ANTENNA_1676 (.A(net107));
 sg13g2_antennanp ANTENNA_1677 (.A(net107));
 sg13g2_antennanp ANTENNA_1678 (.A(net107));
 sg13g2_antennanp ANTENNA_1679 (.A(net107));
 sg13g2_antennanp ANTENNA_1680 (.A(net107));
 sg13g2_antennanp ANTENNA_1681 (.A(net107));
 sg13g2_antennanp ANTENNA_1682 (.A(net107));
 sg13g2_antennanp ANTENNA_1683 (.A(net107));
 sg13g2_antennanp ANTENNA_1684 (.A(net107));
 sg13g2_antennanp ANTENNA_1685 (.A(net107));
 sg13g2_antennanp ANTENNA_1686 (.A(net107));
 sg13g2_antennanp ANTENNA_1687 (.A(net107));
 sg13g2_antennanp ANTENNA_1688 (.A(net107));
 sg13g2_antennanp ANTENNA_1689 (.A(net107));
 sg13g2_antennanp ANTENNA_1690 (.A(net107));
 sg13g2_antennanp ANTENNA_1691 (.A(net108));
 sg13g2_antennanp ANTENNA_1692 (.A(net108));
 sg13g2_antennanp ANTENNA_1693 (.A(net108));
 sg13g2_antennanp ANTENNA_1694 (.A(net108));
 sg13g2_antennanp ANTENNA_1695 (.A(net108));
 sg13g2_antennanp ANTENNA_1696 (.A(net108));
 sg13g2_antennanp ANTENNA_1697 (.A(net108));
 sg13g2_antennanp ANTENNA_1698 (.A(net108));
 sg13g2_antennanp ANTENNA_1699 (.A(net108));
 sg13g2_antennanp ANTENNA_1700 (.A(net108));
 sg13g2_antennanp ANTENNA_1701 (.A(net108));
 sg13g2_antennanp ANTENNA_1702 (.A(net108));
 sg13g2_antennanp ANTENNA_1703 (.A(net108));
 sg13g2_antennanp ANTENNA_1704 (.A(net108));
 sg13g2_antennanp ANTENNA_1705 (.A(net108));
 sg13g2_antennanp ANTENNA_1706 (.A(net108));
 sg13g2_antennanp ANTENNA_1707 (.A(net113));
 sg13g2_antennanp ANTENNA_1708 (.A(net113));
 sg13g2_antennanp ANTENNA_1709 (.A(net113));
 sg13g2_antennanp ANTENNA_1710 (.A(net113));
 sg13g2_antennanp ANTENNA_1711 (.A(net113));
 sg13g2_antennanp ANTENNA_1712 (.A(net113));
 sg13g2_antennanp ANTENNA_1713 (.A(net113));
 sg13g2_antennanp ANTENNA_1714 (.A(net113));
 sg13g2_antennanp ANTENNA_1715 (.A(net113));
 sg13g2_antennanp ANTENNA_1716 (.A(net113));
 sg13g2_antennanp ANTENNA_1717 (.A(net113));
 sg13g2_antennanp ANTENNA_1718 (.A(net113));
 sg13g2_antennanp ANTENNA_1719 (.A(net113));
 sg13g2_antennanp ANTENNA_1720 (.A(net113));
 sg13g2_antennanp ANTENNA_1721 (.A(net113));
 sg13g2_antennanp ANTENNA_1722 (.A(net118));
 sg13g2_antennanp ANTENNA_1723 (.A(net118));
 sg13g2_antennanp ANTENNA_1724 (.A(net118));
 sg13g2_antennanp ANTENNA_1725 (.A(net118));
 sg13g2_antennanp ANTENNA_1726 (.A(net118));
 sg13g2_antennanp ANTENNA_1727 (.A(net118));
 sg13g2_antennanp ANTENNA_1728 (.A(net118));
 sg13g2_antennanp ANTENNA_1729 (.A(net118));
 sg13g2_antennanp ANTENNA_1730 (.A(net118));
 sg13g2_antennanp ANTENNA_1731 (.A(net118));
 sg13g2_antennanp ANTENNA_1732 (.A(net118));
 sg13g2_antennanp ANTENNA_1733 (.A(net118));
 sg13g2_antennanp ANTENNA_1734 (.A(net118));
 sg13g2_antennanp ANTENNA_1735 (.A(net118));
 sg13g2_antennanp ANTENNA_1736 (.A(net118));
 sg13g2_antennanp ANTENNA_1737 (.A(net118));
 sg13g2_antennanp ANTENNA_1738 (.A(net118));
 sg13g2_antennanp ANTENNA_1739 (.A(net118));
 sg13g2_antennanp ANTENNA_1740 (.A(net118));
 sg13g2_antennanp ANTENNA_1741 (.A(net118));
 sg13g2_antennanp ANTENNA_1742 (.A(net118));
 sg13g2_antennanp ANTENNA_1743 (.A(net119));
 sg13g2_antennanp ANTENNA_1744 (.A(net119));
 sg13g2_antennanp ANTENNA_1745 (.A(net119));
 sg13g2_antennanp ANTENNA_1746 (.A(net119));
 sg13g2_antennanp ANTENNA_1747 (.A(net119));
 sg13g2_antennanp ANTENNA_1748 (.A(net119));
 sg13g2_antennanp ANTENNA_1749 (.A(net119));
 sg13g2_antennanp ANTENNA_1750 (.A(net119));
 sg13g2_antennanp ANTENNA_1751 (.A(net124));
 sg13g2_antennanp ANTENNA_1752 (.A(net124));
 sg13g2_antennanp ANTENNA_1753 (.A(net124));
 sg13g2_antennanp ANTENNA_1754 (.A(net124));
 sg13g2_antennanp ANTENNA_1755 (.A(net124));
 sg13g2_antennanp ANTENNA_1756 (.A(net124));
 sg13g2_antennanp ANTENNA_1757 (.A(net124));
 sg13g2_antennanp ANTENNA_1758 (.A(net124));
 sg13g2_antennanp ANTENNA_1759 (.A(net127));
 sg13g2_antennanp ANTENNA_1760 (.A(net127));
 sg13g2_antennanp ANTENNA_1761 (.A(net127));
 sg13g2_antennanp ANTENNA_1762 (.A(net127));
 sg13g2_antennanp ANTENNA_1763 (.A(net127));
 sg13g2_antennanp ANTENNA_1764 (.A(net127));
 sg13g2_antennanp ANTENNA_1765 (.A(net127));
 sg13g2_antennanp ANTENNA_1766 (.A(net127));
 sg13g2_antennanp ANTENNA_1767 (.A(net127));
 sg13g2_antennanp ANTENNA_1768 (.A(net127));
 sg13g2_antennanp ANTENNA_1769 (.A(net127));
 sg13g2_antennanp ANTENNA_1770 (.A(net127));
 sg13g2_antennanp ANTENNA_1771 (.A(net127));
 sg13g2_antennanp ANTENNA_1772 (.A(net127));
 sg13g2_antennanp ANTENNA_1773 (.A(net127));
 sg13g2_antennanp ANTENNA_1774 (.A(net368));
 sg13g2_antennanp ANTENNA_1775 (.A(net368));
 sg13g2_antennanp ANTENNA_1776 (.A(net368));
 sg13g2_antennanp ANTENNA_1777 (.A(net368));
 sg13g2_antennanp ANTENNA_1778 (.A(net368));
 sg13g2_antennanp ANTENNA_1779 (.A(net368));
 sg13g2_antennanp ANTENNA_1780 (.A(net368));
 sg13g2_antennanp ANTENNA_1781 (.A(net368));
 sg13g2_antennanp ANTENNA_1782 (.A(net386));
 sg13g2_antennanp ANTENNA_1783 (.A(net386));
 sg13g2_antennanp ANTENNA_1784 (.A(net386));
 sg13g2_antennanp ANTENNA_1785 (.A(net386));
 sg13g2_antennanp ANTENNA_1786 (.A(net386));
 sg13g2_antennanp ANTENNA_1787 (.A(net386));
 sg13g2_antennanp ANTENNA_1788 (.A(net386));
 sg13g2_antennanp ANTENNA_1789 (.A(net386));
 sg13g2_antennanp ANTENNA_1790 (.A(net386));
 sg13g2_antennanp ANTENNA_1791 (.A(net386));
 sg13g2_antennanp ANTENNA_1792 (.A(net386));
 sg13g2_antennanp ANTENNA_1793 (.A(net386));
 sg13g2_antennanp ANTENNA_1794 (.A(net386));
 sg13g2_antennanp ANTENNA_1795 (.A(net386));
 sg13g2_antennanp ANTENNA_1796 (.A(net386));
 sg13g2_antennanp ANTENNA_1797 (.A(net386));
 sg13g2_antennanp ANTENNA_1798 (.A(net386));
 sg13g2_antennanp ANTENNA_1799 (.A(net716));
 sg13g2_antennanp ANTENNA_1800 (.A(net716));
 sg13g2_antennanp ANTENNA_1801 (.A(net716));
 sg13g2_antennanp ANTENNA_1802 (.A(net716));
 sg13g2_antennanp ANTENNA_1803 (.A(net716));
 sg13g2_antennanp ANTENNA_1804 (.A(net716));
 sg13g2_antennanp ANTENNA_1805 (.A(net716));
 sg13g2_antennanp ANTENNA_1806 (.A(net716));
 sg13g2_antennanp ANTENNA_1807 (.A(_00534_));
 sg13g2_antennanp ANTENNA_1808 (.A(_01440_));
 sg13g2_antennanp ANTENNA_1809 (.A(_01440_));
 sg13g2_antennanp ANTENNA_1810 (.A(_01795_));
 sg13g2_antennanp ANTENNA_1811 (.A(_01795_));
 sg13g2_antennanp ANTENNA_1812 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1813 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1814 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1815 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1816 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1817 (.A(_02787_));
 sg13g2_antennanp ANTENNA_1818 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1819 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1820 (.A(_03810_));
 sg13g2_antennanp ANTENNA_1821 (.A(_03821_));
 sg13g2_antennanp ANTENNA_1822 (.A(_03821_));
 sg13g2_antennanp ANTENNA_1823 (.A(_03821_));
 sg13g2_antennanp ANTENNA_1824 (.A(_03821_));
 sg13g2_antennanp ANTENNA_1825 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1826 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1827 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1828 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1829 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1830 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1831 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1832 (.A(_04067_));
 sg13g2_antennanp ANTENNA_1833 (.A(_04077_));
 sg13g2_antennanp ANTENNA_1834 (.A(_04077_));
 sg13g2_antennanp ANTENNA_1835 (.A(_04077_));
 sg13g2_antennanp ANTENNA_1836 (.A(_04077_));
 sg13g2_antennanp ANTENNA_1837 (.A(_04077_));
 sg13g2_antennanp ANTENNA_1838 (.A(_04077_));
 sg13g2_antennanp ANTENNA_1839 (.A(_04242_));
 sg13g2_antennanp ANTENNA_1840 (.A(_04242_));
 sg13g2_antennanp ANTENNA_1841 (.A(_04371_));
 sg13g2_antennanp ANTENNA_1842 (.A(_04378_));
 sg13g2_antennanp ANTENNA_1843 (.A(_04393_));
 sg13g2_antennanp ANTENNA_1844 (.A(_04403_));
 sg13g2_antennanp ANTENNA_1845 (.A(_04411_));
 sg13g2_antennanp ANTENNA_1846 (.A(_04412_));
 sg13g2_antennanp ANTENNA_1847 (.A(_04416_));
 sg13g2_antennanp ANTENNA_1848 (.A(_04419_));
 sg13g2_antennanp ANTENNA_1849 (.A(_04432_));
 sg13g2_antennanp ANTENNA_1850 (.A(_04453_));
 sg13g2_antennanp ANTENNA_1851 (.A(_04481_));
 sg13g2_antennanp ANTENNA_1852 (.A(_04508_));
 sg13g2_antennanp ANTENNA_1853 (.A(_04756_));
 sg13g2_antennanp ANTENNA_1854 (.A(_04773_));
 sg13g2_antennanp ANTENNA_1855 (.A(_04804_));
 sg13g2_antennanp ANTENNA_1856 (.A(_04816_));
 sg13g2_antennanp ANTENNA_1857 (.A(_04828_));
 sg13g2_antennanp ANTENNA_1858 (.A(_04838_));
 sg13g2_antennanp ANTENNA_1859 (.A(_04840_));
 sg13g2_antennanp ANTENNA_1860 (.A(_04842_));
 sg13g2_antennanp ANTENNA_1861 (.A(_04850_));
 sg13g2_antennanp ANTENNA_1862 (.A(_04853_));
 sg13g2_antennanp ANTENNA_1863 (.A(_04860_));
 sg13g2_antennanp ANTENNA_1864 (.A(_04860_));
 sg13g2_antennanp ANTENNA_1865 (.A(_04860_));
 sg13g2_antennanp ANTENNA_1866 (.A(_04914_));
 sg13g2_antennanp ANTENNA_1867 (.A(_04914_));
 sg13g2_antennanp ANTENNA_1868 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1869 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1870 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1871 (.A(_04941_));
 sg13g2_antennanp ANTENNA_1872 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1873 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1874 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1875 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1876 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1877 (.A(_05131_));
 sg13g2_antennanp ANTENNA_1878 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1879 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1880 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1881 (.A(_05416_));
 sg13g2_antennanp ANTENNA_1882 (.A(_05416_));
 sg13g2_antennanp ANTENNA_1883 (.A(_05416_));
 sg13g2_antennanp ANTENNA_1884 (.A(_05757_));
 sg13g2_antennanp ANTENNA_1885 (.A(_05757_));
 sg13g2_antennanp ANTENNA_1886 (.A(_05757_));
 sg13g2_antennanp ANTENNA_1887 (.A(_05757_));
 sg13g2_antennanp ANTENNA_1888 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1889 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1890 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1891 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1892 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1893 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1894 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1895 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1896 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1897 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1898 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1899 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1900 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1901 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1902 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1903 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1904 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1905 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1906 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1907 (.A(_06111_));
 sg13g2_antennanp ANTENNA_1908 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1909 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1910 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1911 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1912 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1913 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1914 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1915 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1916 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1917 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1918 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1919 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1920 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1921 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1922 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1923 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1924 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1925 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1926 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1927 (.A(_06900_));
 sg13g2_antennanp ANTENNA_1928 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1929 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1930 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1931 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1932 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1933 (.A(_07117_));
 sg13g2_antennanp ANTENNA_1934 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1935 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1936 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1937 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1938 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1939 (.A(_08349_));
 sg13g2_antennanp ANTENNA_1940 (.A(_08737_));
 sg13g2_antennanp ANTENNA_1941 (.A(_08737_));
 sg13g2_antennanp ANTENNA_1942 (.A(_08737_));
 sg13g2_antennanp ANTENNA_1943 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1944 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1945 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1946 (.A(_10237_));
 sg13g2_antennanp ANTENNA_1947 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1948 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1949 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1950 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1951 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1952 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1953 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1954 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1955 (.A(_11347_));
 sg13g2_antennanp ANTENNA_1956 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1957 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1958 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1959 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1960 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1961 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1962 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1963 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1964 (.A(_12651_));
 sg13g2_antennanp ANTENNA_1965 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1966 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1967 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1968 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1969 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1970 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1971 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1972 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1973 (.A(_12999_));
 sg13g2_antennanp ANTENNA_1974 (.A(net31));
 sg13g2_antennanp ANTENNA_1975 (.A(net31));
 sg13g2_antennanp ANTENNA_1976 (.A(net31));
 sg13g2_antennanp ANTENNA_1977 (.A(net31));
 sg13g2_antennanp ANTENNA_1978 (.A(net31));
 sg13g2_antennanp ANTENNA_1979 (.A(net31));
 sg13g2_antennanp ANTENNA_1980 (.A(net31));
 sg13g2_antennanp ANTENNA_1981 (.A(net31));
 sg13g2_antennanp ANTENNA_1982 (.A(net31));
 sg13g2_antennanp ANTENNA_1983 (.A(net31));
 sg13g2_antennanp ANTENNA_1984 (.A(net31));
 sg13g2_antennanp ANTENNA_1985 (.A(net31));
 sg13g2_antennanp ANTENNA_1986 (.A(net31));
 sg13g2_antennanp ANTENNA_1987 (.A(net31));
 sg13g2_antennanp ANTENNA_1988 (.A(net31));
 sg13g2_antennanp ANTENNA_1989 (.A(net31));
 sg13g2_antennanp ANTENNA_1990 (.A(net31));
 sg13g2_antennanp ANTENNA_1991 (.A(net31));
 sg13g2_antennanp ANTENNA_1992 (.A(net31));
 sg13g2_antennanp ANTENNA_1993 (.A(net31));
 sg13g2_antennanp ANTENNA_1994 (.A(net31));
 sg13g2_antennanp ANTENNA_1995 (.A(net31));
 sg13g2_antennanp ANTENNA_1996 (.A(net31));
 sg13g2_antennanp ANTENNA_1997 (.A(net31));
 sg13g2_antennanp ANTENNA_1998 (.A(net31));
 sg13g2_antennanp ANTENNA_1999 (.A(net31));
 sg13g2_antennanp ANTENNA_2000 (.A(net43));
 sg13g2_antennanp ANTENNA_2001 (.A(net43));
 sg13g2_antennanp ANTENNA_2002 (.A(net43));
 sg13g2_antennanp ANTENNA_2003 (.A(net43));
 sg13g2_antennanp ANTENNA_2004 (.A(net43));
 sg13g2_antennanp ANTENNA_2005 (.A(net43));
 sg13g2_antennanp ANTENNA_2006 (.A(net43));
 sg13g2_antennanp ANTENNA_2007 (.A(net43));
 sg13g2_antennanp ANTENNA_2008 (.A(net43));
 sg13g2_antennanp ANTENNA_2009 (.A(net43));
 sg13g2_antennanp ANTENNA_2010 (.A(net43));
 sg13g2_antennanp ANTENNA_2011 (.A(net43));
 sg13g2_antennanp ANTENNA_2012 (.A(net43));
 sg13g2_antennanp ANTENNA_2013 (.A(net43));
 sg13g2_antennanp ANTENNA_2014 (.A(net73));
 sg13g2_antennanp ANTENNA_2015 (.A(net73));
 sg13g2_antennanp ANTENNA_2016 (.A(net73));
 sg13g2_antennanp ANTENNA_2017 (.A(net73));
 sg13g2_antennanp ANTENNA_2018 (.A(net73));
 sg13g2_antennanp ANTENNA_2019 (.A(net73));
 sg13g2_antennanp ANTENNA_2020 (.A(net73));
 sg13g2_antennanp ANTENNA_2021 (.A(net73));
 sg13g2_antennanp ANTENNA_2022 (.A(net73));
 sg13g2_antennanp ANTENNA_2023 (.A(net75));
 sg13g2_antennanp ANTENNA_2024 (.A(net75));
 sg13g2_antennanp ANTENNA_2025 (.A(net75));
 sg13g2_antennanp ANTENNA_2026 (.A(net75));
 sg13g2_antennanp ANTENNA_2027 (.A(net75));
 sg13g2_antennanp ANTENNA_2028 (.A(net75));
 sg13g2_antennanp ANTENNA_2029 (.A(net75));
 sg13g2_antennanp ANTENNA_2030 (.A(net75));
 sg13g2_antennanp ANTENNA_2031 (.A(net75));
 sg13g2_antennanp ANTENNA_2032 (.A(net75));
 sg13g2_antennanp ANTENNA_2033 (.A(net75));
 sg13g2_antennanp ANTENNA_2034 (.A(net75));
 sg13g2_antennanp ANTENNA_2035 (.A(net75));
 sg13g2_antennanp ANTENNA_2036 (.A(net75));
 sg13g2_antennanp ANTENNA_2037 (.A(net75));
 sg13g2_antennanp ANTENNA_2038 (.A(net75));
 sg13g2_antennanp ANTENNA_2039 (.A(net75));
 sg13g2_antennanp ANTENNA_2040 (.A(net75));
 sg13g2_antennanp ANTENNA_2041 (.A(net75));
 sg13g2_antennanp ANTENNA_2042 (.A(net75));
 sg13g2_antennanp ANTENNA_2043 (.A(net75));
 sg13g2_antennanp ANTENNA_2044 (.A(net79));
 sg13g2_antennanp ANTENNA_2045 (.A(net79));
 sg13g2_antennanp ANTENNA_2046 (.A(net79));
 sg13g2_antennanp ANTENNA_2047 (.A(net79));
 sg13g2_antennanp ANTENNA_2048 (.A(net79));
 sg13g2_antennanp ANTENNA_2049 (.A(net79));
 sg13g2_antennanp ANTENNA_2050 (.A(net79));
 sg13g2_antennanp ANTENNA_2051 (.A(net79));
 sg13g2_antennanp ANTENNA_2052 (.A(net79));
 sg13g2_antennanp ANTENNA_2053 (.A(net79));
 sg13g2_antennanp ANTENNA_2054 (.A(net79));
 sg13g2_antennanp ANTENNA_2055 (.A(net79));
 sg13g2_antennanp ANTENNA_2056 (.A(net79));
 sg13g2_antennanp ANTENNA_2057 (.A(net79));
 sg13g2_antennanp ANTENNA_2058 (.A(net79));
 sg13g2_antennanp ANTENNA_2059 (.A(net79));
 sg13g2_antennanp ANTENNA_2060 (.A(net79));
 sg13g2_antennanp ANTENNA_2061 (.A(net79));
 sg13g2_antennanp ANTENNA_2062 (.A(net79));
 sg13g2_antennanp ANTENNA_2063 (.A(net79));
 sg13g2_antennanp ANTENNA_2064 (.A(net79));
 sg13g2_antennanp ANTENNA_2065 (.A(net79));
 sg13g2_antennanp ANTENNA_2066 (.A(net79));
 sg13g2_antennanp ANTENNA_2067 (.A(net79));
 sg13g2_antennanp ANTENNA_2068 (.A(net79));
 sg13g2_antennanp ANTENNA_2069 (.A(net79));
 sg13g2_antennanp ANTENNA_2070 (.A(net79));
 sg13g2_antennanp ANTENNA_2071 (.A(net79));
 sg13g2_antennanp ANTENNA_2072 (.A(net79));
 sg13g2_antennanp ANTENNA_2073 (.A(net79));
 sg13g2_antennanp ANTENNA_2074 (.A(net79));
 sg13g2_antennanp ANTENNA_2075 (.A(net79));
 sg13g2_antennanp ANTENNA_2076 (.A(net79));
 sg13g2_antennanp ANTENNA_2077 (.A(net79));
 sg13g2_antennanp ANTENNA_2078 (.A(net79));
 sg13g2_antennanp ANTENNA_2079 (.A(net79));
 sg13g2_antennanp ANTENNA_2080 (.A(net80));
 sg13g2_antennanp ANTENNA_2081 (.A(net80));
 sg13g2_antennanp ANTENNA_2082 (.A(net80));
 sg13g2_antennanp ANTENNA_2083 (.A(net80));
 sg13g2_antennanp ANTENNA_2084 (.A(net80));
 sg13g2_antennanp ANTENNA_2085 (.A(net80));
 sg13g2_antennanp ANTENNA_2086 (.A(net80));
 sg13g2_antennanp ANTENNA_2087 (.A(net80));
 sg13g2_antennanp ANTENNA_2088 (.A(net82));
 sg13g2_antennanp ANTENNA_2089 (.A(net82));
 sg13g2_antennanp ANTENNA_2090 (.A(net82));
 sg13g2_antennanp ANTENNA_2091 (.A(net82));
 sg13g2_antennanp ANTENNA_2092 (.A(net82));
 sg13g2_antennanp ANTENNA_2093 (.A(net82));
 sg13g2_antennanp ANTENNA_2094 (.A(net82));
 sg13g2_antennanp ANTENNA_2095 (.A(net82));
 sg13g2_antennanp ANTENNA_2096 (.A(net82));
 sg13g2_antennanp ANTENNA_2097 (.A(net82));
 sg13g2_antennanp ANTENNA_2098 (.A(net82));
 sg13g2_antennanp ANTENNA_2099 (.A(net82));
 sg13g2_antennanp ANTENNA_2100 (.A(net82));
 sg13g2_antennanp ANTENNA_2101 (.A(net82));
 sg13g2_antennanp ANTENNA_2102 (.A(net82));
 sg13g2_antennanp ANTENNA_2103 (.A(net82));
 sg13g2_antennanp ANTENNA_2104 (.A(net82));
 sg13g2_antennanp ANTENNA_2105 (.A(net103));
 sg13g2_antennanp ANTENNA_2106 (.A(net103));
 sg13g2_antennanp ANTENNA_2107 (.A(net103));
 sg13g2_antennanp ANTENNA_2108 (.A(net103));
 sg13g2_antennanp ANTENNA_2109 (.A(net103));
 sg13g2_antennanp ANTENNA_2110 (.A(net103));
 sg13g2_antennanp ANTENNA_2111 (.A(net103));
 sg13g2_antennanp ANTENNA_2112 (.A(net103));
 sg13g2_antennanp ANTENNA_2113 (.A(net108));
 sg13g2_antennanp ANTENNA_2114 (.A(net108));
 sg13g2_antennanp ANTENNA_2115 (.A(net108));
 sg13g2_antennanp ANTENNA_2116 (.A(net108));
 sg13g2_antennanp ANTENNA_2117 (.A(net108));
 sg13g2_antennanp ANTENNA_2118 (.A(net108));
 sg13g2_antennanp ANTENNA_2119 (.A(net108));
 sg13g2_antennanp ANTENNA_2120 (.A(net108));
 sg13g2_antennanp ANTENNA_2121 (.A(net108));
 sg13g2_antennanp ANTENNA_2122 (.A(net108));
 sg13g2_antennanp ANTENNA_2123 (.A(net108));
 sg13g2_antennanp ANTENNA_2124 (.A(net108));
 sg13g2_antennanp ANTENNA_2125 (.A(net108));
 sg13g2_antennanp ANTENNA_2126 (.A(net108));
 sg13g2_antennanp ANTENNA_2127 (.A(net108));
 sg13g2_antennanp ANTENNA_2128 (.A(net108));
 sg13g2_antennanp ANTENNA_2129 (.A(net113));
 sg13g2_antennanp ANTENNA_2130 (.A(net113));
 sg13g2_antennanp ANTENNA_2131 (.A(net113));
 sg13g2_antennanp ANTENNA_2132 (.A(net113));
 sg13g2_antennanp ANTENNA_2133 (.A(net113));
 sg13g2_antennanp ANTENNA_2134 (.A(net113));
 sg13g2_antennanp ANTENNA_2135 (.A(net113));
 sg13g2_antennanp ANTENNA_2136 (.A(net113));
 sg13g2_antennanp ANTENNA_2137 (.A(net113));
 sg13g2_antennanp ANTENNA_2138 (.A(net113));
 sg13g2_antennanp ANTENNA_2139 (.A(net113));
 sg13g2_antennanp ANTENNA_2140 (.A(net113));
 sg13g2_antennanp ANTENNA_2141 (.A(net113));
 sg13g2_antennanp ANTENNA_2142 (.A(net113));
 sg13g2_antennanp ANTENNA_2143 (.A(net113));
 sg13g2_antennanp ANTENNA_2144 (.A(net118));
 sg13g2_antennanp ANTENNA_2145 (.A(net118));
 sg13g2_antennanp ANTENNA_2146 (.A(net118));
 sg13g2_antennanp ANTENNA_2147 (.A(net118));
 sg13g2_antennanp ANTENNA_2148 (.A(net118));
 sg13g2_antennanp ANTENNA_2149 (.A(net118));
 sg13g2_antennanp ANTENNA_2150 (.A(net118));
 sg13g2_antennanp ANTENNA_2151 (.A(net118));
 sg13g2_antennanp ANTENNA_2152 (.A(net118));
 sg13g2_antennanp ANTENNA_2153 (.A(net118));
 sg13g2_antennanp ANTENNA_2154 (.A(net118));
 sg13g2_antennanp ANTENNA_2155 (.A(net118));
 sg13g2_antennanp ANTENNA_2156 (.A(net118));
 sg13g2_antennanp ANTENNA_2157 (.A(net118));
 sg13g2_antennanp ANTENNA_2158 (.A(net118));
 sg13g2_antennanp ANTENNA_2159 (.A(net118));
 sg13g2_antennanp ANTENNA_2160 (.A(net118));
 sg13g2_antennanp ANTENNA_2161 (.A(net118));
 sg13g2_antennanp ANTENNA_2162 (.A(net118));
 sg13g2_antennanp ANTENNA_2163 (.A(net118));
 sg13g2_antennanp ANTENNA_2164 (.A(net118));
 sg13g2_antennanp ANTENNA_2165 (.A(net124));
 sg13g2_antennanp ANTENNA_2166 (.A(net124));
 sg13g2_antennanp ANTENNA_2167 (.A(net124));
 sg13g2_antennanp ANTENNA_2168 (.A(net124));
 sg13g2_antennanp ANTENNA_2169 (.A(net124));
 sg13g2_antennanp ANTENNA_2170 (.A(net124));
 sg13g2_antennanp ANTENNA_2171 (.A(net124));
 sg13g2_antennanp ANTENNA_2172 (.A(net124));
 sg13g2_antennanp ANTENNA_2173 (.A(net124));
 sg13g2_antennanp ANTENNA_2174 (.A(net124));
 sg13g2_antennanp ANTENNA_2175 (.A(net124));
 sg13g2_antennanp ANTENNA_2176 (.A(net124));
 sg13g2_antennanp ANTENNA_2177 (.A(net124));
 sg13g2_antennanp ANTENNA_2178 (.A(net127));
 sg13g2_antennanp ANTENNA_2179 (.A(net127));
 sg13g2_antennanp ANTENNA_2180 (.A(net127));
 sg13g2_antennanp ANTENNA_2181 (.A(net127));
 sg13g2_antennanp ANTENNA_2182 (.A(net127));
 sg13g2_antennanp ANTENNA_2183 (.A(net127));
 sg13g2_antennanp ANTENNA_2184 (.A(net127));
 sg13g2_antennanp ANTENNA_2185 (.A(net127));
 sg13g2_antennanp ANTENNA_2186 (.A(net127));
 sg13g2_antennanp ANTENNA_2187 (.A(net127));
 sg13g2_antennanp ANTENNA_2188 (.A(net127));
 sg13g2_antennanp ANTENNA_2189 (.A(net127));
 sg13g2_antennanp ANTENNA_2190 (.A(net127));
 sg13g2_antennanp ANTENNA_2191 (.A(net166));
 sg13g2_antennanp ANTENNA_2192 (.A(net166));
 sg13g2_antennanp ANTENNA_2193 (.A(net166));
 sg13g2_antennanp ANTENNA_2194 (.A(net166));
 sg13g2_antennanp ANTENNA_2195 (.A(net166));
 sg13g2_antennanp ANTENNA_2196 (.A(net166));
 sg13g2_antennanp ANTENNA_2197 (.A(net166));
 sg13g2_antennanp ANTENNA_2198 (.A(net166));
 sg13g2_antennanp ANTENNA_2199 (.A(net368));
 sg13g2_antennanp ANTENNA_2200 (.A(net368));
 sg13g2_antennanp ANTENNA_2201 (.A(net368));
 sg13g2_antennanp ANTENNA_2202 (.A(net368));
 sg13g2_antennanp ANTENNA_2203 (.A(net368));
 sg13g2_antennanp ANTENNA_2204 (.A(net368));
 sg13g2_antennanp ANTENNA_2205 (.A(net368));
 sg13g2_antennanp ANTENNA_2206 (.A(net368));
 sg13g2_antennanp ANTENNA_2207 (.A(net368));
 sg13g2_antennanp ANTENNA_2208 (.A(net368));
 sg13g2_antennanp ANTENNA_2209 (.A(net368));
 sg13g2_antennanp ANTENNA_2210 (.A(net368));
 sg13g2_antennanp ANTENNA_2211 (.A(net368));
 sg13g2_antennanp ANTENNA_2212 (.A(net368));
 sg13g2_antennanp ANTENNA_2213 (.A(net368));
 sg13g2_antennanp ANTENNA_2214 (.A(net368));
 sg13g2_antennanp ANTENNA_2215 (.A(net386));
 sg13g2_antennanp ANTENNA_2216 (.A(net386));
 sg13g2_antennanp ANTENNA_2217 (.A(net386));
 sg13g2_antennanp ANTENNA_2218 (.A(net386));
 sg13g2_antennanp ANTENNA_2219 (.A(net386));
 sg13g2_antennanp ANTENNA_2220 (.A(net386));
 sg13g2_antennanp ANTENNA_2221 (.A(net386));
 sg13g2_antennanp ANTENNA_2222 (.A(net386));
 sg13g2_antennanp ANTENNA_2223 (.A(net386));
 sg13g2_antennanp ANTENNA_2224 (.A(net386));
 sg13g2_antennanp ANTENNA_2225 (.A(net386));
 sg13g2_antennanp ANTENNA_2226 (.A(net386));
 sg13g2_antennanp ANTENNA_2227 (.A(net386));
 sg13g2_antennanp ANTENNA_2228 (.A(net386));
 sg13g2_antennanp ANTENNA_2229 (.A(net386));
 sg13g2_antennanp ANTENNA_2230 (.A(net386));
 sg13g2_antennanp ANTENNA_2231 (.A(net386));
 sg13g2_antennanp ANTENNA_2232 (.A(net1002));
 sg13g2_antennanp ANTENNA_2233 (.A(net1002));
 sg13g2_antennanp ANTENNA_2234 (.A(net1002));
 sg13g2_antennanp ANTENNA_2235 (.A(net1002));
 sg13g2_antennanp ANTENNA_2236 (.A(net1002));
 sg13g2_antennanp ANTENNA_2237 (.A(net1002));
 sg13g2_antennanp ANTENNA_2238 (.A(net1002));
 sg13g2_antennanp ANTENNA_2239 (.A(net1002));
 sg13g2_antennanp ANTENNA_2240 (.A(net1002));
 sg13g2_antennanp ANTENNA_2241 (.A(net1002));
 sg13g2_antennanp ANTENNA_2242 (.A(net1002));
 sg13g2_antennanp ANTENNA_2243 (.A(net1002));
 sg13g2_antennanp ANTENNA_2244 (.A(net1002));
 sg13g2_antennanp ANTENNA_2245 (.A(net1002));
 sg13g2_antennanp ANTENNA_2246 (.A(_00534_));
 sg13g2_antennanp ANTENNA_2247 (.A(_01440_));
 sg13g2_antennanp ANTENNA_2248 (.A(_01440_));
 sg13g2_antennanp ANTENNA_2249 (.A(_01795_));
 sg13g2_antennanp ANTENNA_2250 (.A(_01795_));
 sg13g2_antennanp ANTENNA_2251 (.A(_02787_));
 sg13g2_antennanp ANTENNA_2252 (.A(_02787_));
 sg13g2_antennanp ANTENNA_2253 (.A(_02787_));
 sg13g2_antennanp ANTENNA_2254 (.A(_02787_));
 sg13g2_antennanp ANTENNA_2255 (.A(_02787_));
 sg13g2_antennanp ANTENNA_2256 (.A(_02787_));
 sg13g2_antennanp ANTENNA_2257 (.A(_03810_));
 sg13g2_antennanp ANTENNA_2258 (.A(_03810_));
 sg13g2_antennanp ANTENNA_2259 (.A(_03810_));
 sg13g2_antennanp ANTENNA_2260 (.A(_03821_));
 sg13g2_antennanp ANTENNA_2261 (.A(_03821_));
 sg13g2_antennanp ANTENNA_2262 (.A(_03821_));
 sg13g2_antennanp ANTENNA_2263 (.A(_03821_));
 sg13g2_antennanp ANTENNA_2264 (.A(_04067_));
 sg13g2_antennanp ANTENNA_2265 (.A(_04067_));
 sg13g2_antennanp ANTENNA_2266 (.A(_04067_));
 sg13g2_antennanp ANTENNA_2267 (.A(_04067_));
 sg13g2_antennanp ANTENNA_2268 (.A(_04067_));
 sg13g2_antennanp ANTENNA_2269 (.A(_04067_));
 sg13g2_antennanp ANTENNA_2270 (.A(_04067_));
 sg13g2_antennanp ANTENNA_2271 (.A(_04067_));
 sg13g2_antennanp ANTENNA_2272 (.A(_04067_));
 sg13g2_antennanp ANTENNA_2273 (.A(_04077_));
 sg13g2_antennanp ANTENNA_2274 (.A(_04077_));
 sg13g2_antennanp ANTENNA_2275 (.A(_04077_));
 sg13g2_antennanp ANTENNA_2276 (.A(_04077_));
 sg13g2_antennanp ANTENNA_2277 (.A(_04077_));
 sg13g2_antennanp ANTENNA_2278 (.A(_04077_));
 sg13g2_antennanp ANTENNA_2279 (.A(_04242_));
 sg13g2_antennanp ANTENNA_2280 (.A(_04242_));
 sg13g2_antennanp ANTENNA_2281 (.A(_04371_));
 sg13g2_antennanp ANTENNA_2282 (.A(_04378_));
 sg13g2_antennanp ANTENNA_2283 (.A(_04393_));
 sg13g2_antennanp ANTENNA_2284 (.A(_04403_));
 sg13g2_antennanp ANTENNA_2285 (.A(_04411_));
 sg13g2_antennanp ANTENNA_2286 (.A(_04412_));
 sg13g2_antennanp ANTENNA_2287 (.A(_04416_));
 sg13g2_antennanp ANTENNA_2288 (.A(_04419_));
 sg13g2_antennanp ANTENNA_2289 (.A(_04432_));
 sg13g2_antennanp ANTENNA_2290 (.A(_04453_));
 sg13g2_antennanp ANTENNA_2291 (.A(_04481_));
 sg13g2_antennanp ANTENNA_2292 (.A(_04508_));
 sg13g2_antennanp ANTENNA_2293 (.A(_04508_));
 sg13g2_antennanp ANTENNA_2294 (.A(_04756_));
 sg13g2_antennanp ANTENNA_2295 (.A(_04773_));
 sg13g2_antennanp ANTENNA_2296 (.A(_04804_));
 sg13g2_antennanp ANTENNA_2297 (.A(_04816_));
 sg13g2_antennanp ANTENNA_2298 (.A(_04828_));
 sg13g2_antennanp ANTENNA_2299 (.A(_04838_));
 sg13g2_antennanp ANTENNA_2300 (.A(_04840_));
 sg13g2_antennanp ANTENNA_2301 (.A(_04842_));
 sg13g2_antennanp ANTENNA_2302 (.A(_04850_));
 sg13g2_antennanp ANTENNA_2303 (.A(_04853_));
 sg13g2_antennanp ANTENNA_2304 (.A(_04860_));
 sg13g2_antennanp ANTENNA_2305 (.A(_04860_));
 sg13g2_antennanp ANTENNA_2306 (.A(_04860_));
 sg13g2_antennanp ANTENNA_2307 (.A(_04914_));
 sg13g2_antennanp ANTENNA_2308 (.A(_04914_));
 sg13g2_antennanp ANTENNA_2309 (.A(_04941_));
 sg13g2_antennanp ANTENNA_2310 (.A(_04941_));
 sg13g2_antennanp ANTENNA_2311 (.A(_04941_));
 sg13g2_antennanp ANTENNA_2312 (.A(_04941_));
 sg13g2_antennanp ANTENNA_2313 (.A(_05131_));
 sg13g2_antennanp ANTENNA_2314 (.A(_05131_));
 sg13g2_antennanp ANTENNA_2315 (.A(_05131_));
 sg13g2_antennanp ANTENNA_2316 (.A(_05131_));
 sg13g2_antennanp ANTENNA_2317 (.A(_05131_));
 sg13g2_antennanp ANTENNA_2318 (.A(_05131_));
 sg13g2_antennanp ANTENNA_2319 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2320 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2321 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2322 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2323 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2324 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2325 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2326 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2327 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2328 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2329 (.A(_05416_));
 sg13g2_antennanp ANTENNA_2330 (.A(_05416_));
 sg13g2_antennanp ANTENNA_2331 (.A(_05416_));
 sg13g2_antennanp ANTENNA_2332 (.A(_05416_));
 sg13g2_antennanp ANTENNA_2333 (.A(_05416_));
 sg13g2_antennanp ANTENNA_2334 (.A(_05416_));
 sg13g2_antennanp ANTENNA_2335 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2336 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2337 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2338 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2339 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2340 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2341 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2342 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2343 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2344 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2345 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2346 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2347 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2348 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2349 (.A(_06111_));
 sg13g2_antennanp ANTENNA_2350 (.A(_06111_));
 sg13g2_antennanp ANTENNA_2351 (.A(_06111_));
 sg13g2_antennanp ANTENNA_2352 (.A(_06111_));
 sg13g2_antennanp ANTENNA_2353 (.A(_06111_));
 sg13g2_antennanp ANTENNA_2354 (.A(_06111_));
 sg13g2_antennanp ANTENNA_2355 (.A(_06111_));
 sg13g2_antennanp ANTENNA_2356 (.A(_06111_));
 sg13g2_antennanp ANTENNA_2357 (.A(_06111_));
 sg13g2_antennanp ANTENNA_2358 (.A(_06285_));
 sg13g2_antennanp ANTENNA_2359 (.A(_06285_));
 sg13g2_antennanp ANTENNA_2360 (.A(_06285_));
 sg13g2_antennanp ANTENNA_2361 (.A(_06285_));
 sg13g2_antennanp ANTENNA_2362 (.A(_06285_));
 sg13g2_antennanp ANTENNA_2363 (.A(_06285_));
 sg13g2_antennanp ANTENNA_2364 (.A(_06667_));
 sg13g2_antennanp ANTENNA_2365 (.A(_06667_));
 sg13g2_antennanp ANTENNA_2366 (.A(_06667_));
 sg13g2_antennanp ANTENNA_2367 (.A(_06667_));
 sg13g2_antennanp ANTENNA_2368 (.A(_06900_));
 sg13g2_antennanp ANTENNA_2369 (.A(_06900_));
 sg13g2_antennanp ANTENNA_2370 (.A(_06900_));
 sg13g2_antennanp ANTENNA_2371 (.A(_06900_));
 sg13g2_antennanp ANTENNA_2372 (.A(_07117_));
 sg13g2_antennanp ANTENNA_2373 (.A(_07117_));
 sg13g2_antennanp ANTENNA_2374 (.A(_07117_));
 sg13g2_antennanp ANTENNA_2375 (.A(_08349_));
 sg13g2_antennanp ANTENNA_2376 (.A(_08349_));
 sg13g2_antennanp ANTENNA_2377 (.A(_08349_));
 sg13g2_antennanp ANTENNA_2378 (.A(_08349_));
 sg13g2_antennanp ANTENNA_2379 (.A(_08349_));
 sg13g2_antennanp ANTENNA_2380 (.A(_08349_));
 sg13g2_antennanp ANTENNA_2381 (.A(_08737_));
 sg13g2_antennanp ANTENNA_2382 (.A(_08737_));
 sg13g2_antennanp ANTENNA_2383 (.A(_08737_));
 sg13g2_antennanp ANTENNA_2384 (.A(_10237_));
 sg13g2_antennanp ANTENNA_2385 (.A(_10237_));
 sg13g2_antennanp ANTENNA_2386 (.A(_10237_));
 sg13g2_antennanp ANTENNA_2387 (.A(_10237_));
 sg13g2_antennanp ANTENNA_2388 (.A(_10237_));
 sg13g2_antennanp ANTENNA_2389 (.A(_10237_));
 sg13g2_antennanp ANTENNA_2390 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2391 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2392 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2393 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2394 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2395 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2396 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2397 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2398 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2399 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2400 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2401 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2402 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2403 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2404 (.A(_11347_));
 sg13g2_antennanp ANTENNA_2405 (.A(_12651_));
 sg13g2_antennanp ANTENNA_2406 (.A(_12651_));
 sg13g2_antennanp ANTENNA_2407 (.A(_12651_));
 sg13g2_antennanp ANTENNA_2408 (.A(_12651_));
 sg13g2_antennanp ANTENNA_2409 (.A(_12651_));
 sg13g2_antennanp ANTENNA_2410 (.A(_12651_));
 sg13g2_antennanp ANTENNA_2411 (.A(_12651_));
 sg13g2_antennanp ANTENNA_2412 (.A(_12651_));
 sg13g2_antennanp ANTENNA_2413 (.A(_12651_));
 sg13g2_antennanp ANTENNA_2414 (.A(_12999_));
 sg13g2_antennanp ANTENNA_2415 (.A(_12999_));
 sg13g2_antennanp ANTENNA_2416 (.A(_12999_));
 sg13g2_antennanp ANTENNA_2417 (.A(_12999_));
 sg13g2_antennanp ANTENNA_2418 (.A(_12999_));
 sg13g2_antennanp ANTENNA_2419 (.A(_12999_));
 sg13g2_antennanp ANTENNA_2420 (.A(net31));
 sg13g2_antennanp ANTENNA_2421 (.A(net31));
 sg13g2_antennanp ANTENNA_2422 (.A(net31));
 sg13g2_antennanp ANTENNA_2423 (.A(net31));
 sg13g2_antennanp ANTENNA_2424 (.A(net31));
 sg13g2_antennanp ANTENNA_2425 (.A(net31));
 sg13g2_antennanp ANTENNA_2426 (.A(net31));
 sg13g2_antennanp ANTENNA_2427 (.A(net31));
 sg13g2_antennanp ANTENNA_2428 (.A(net31));
 sg13g2_antennanp ANTENNA_2429 (.A(net31));
 sg13g2_antennanp ANTENNA_2430 (.A(net31));
 sg13g2_antennanp ANTENNA_2431 (.A(net31));
 sg13g2_antennanp ANTENNA_2432 (.A(net31));
 sg13g2_antennanp ANTENNA_2433 (.A(net31));
 sg13g2_antennanp ANTENNA_2434 (.A(net31));
 sg13g2_antennanp ANTENNA_2435 (.A(net31));
 sg13g2_antennanp ANTENNA_2436 (.A(net31));
 sg13g2_antennanp ANTENNA_2437 (.A(net31));
 sg13g2_antennanp ANTENNA_2438 (.A(net31));
 sg13g2_antennanp ANTENNA_2439 (.A(net31));
 sg13g2_antennanp ANTENNA_2440 (.A(net31));
 sg13g2_antennanp ANTENNA_2441 (.A(net31));
 sg13g2_antennanp ANTENNA_2442 (.A(net31));
 sg13g2_antennanp ANTENNA_2443 (.A(net31));
 sg13g2_antennanp ANTENNA_2444 (.A(net31));
 sg13g2_antennanp ANTENNA_2445 (.A(net31));
 sg13g2_antennanp ANTENNA_2446 (.A(net43));
 sg13g2_antennanp ANTENNA_2447 (.A(net43));
 sg13g2_antennanp ANTENNA_2448 (.A(net43));
 sg13g2_antennanp ANTENNA_2449 (.A(net43));
 sg13g2_antennanp ANTENNA_2450 (.A(net43));
 sg13g2_antennanp ANTENNA_2451 (.A(net43));
 sg13g2_antennanp ANTENNA_2452 (.A(net43));
 sg13g2_antennanp ANTENNA_2453 (.A(net43));
 sg13g2_antennanp ANTENNA_2454 (.A(net43));
 sg13g2_antennanp ANTENNA_2455 (.A(net73));
 sg13g2_antennanp ANTENNA_2456 (.A(net73));
 sg13g2_antennanp ANTENNA_2457 (.A(net73));
 sg13g2_antennanp ANTENNA_2458 (.A(net73));
 sg13g2_antennanp ANTENNA_2459 (.A(net73));
 sg13g2_antennanp ANTENNA_2460 (.A(net73));
 sg13g2_antennanp ANTENNA_2461 (.A(net73));
 sg13g2_antennanp ANTENNA_2462 (.A(net73));
 sg13g2_antennanp ANTENNA_2463 (.A(net73));
 sg13g2_antennanp ANTENNA_2464 (.A(net75));
 sg13g2_antennanp ANTENNA_2465 (.A(net75));
 sg13g2_antennanp ANTENNA_2466 (.A(net75));
 sg13g2_antennanp ANTENNA_2467 (.A(net75));
 sg13g2_antennanp ANTENNA_2468 (.A(net75));
 sg13g2_antennanp ANTENNA_2469 (.A(net75));
 sg13g2_antennanp ANTENNA_2470 (.A(net75));
 sg13g2_antennanp ANTENNA_2471 (.A(net75));
 sg13g2_antennanp ANTENNA_2472 (.A(net75));
 sg13g2_antennanp ANTENNA_2473 (.A(net75));
 sg13g2_antennanp ANTENNA_2474 (.A(net75));
 sg13g2_antennanp ANTENNA_2475 (.A(net75));
 sg13g2_antennanp ANTENNA_2476 (.A(net75));
 sg13g2_antennanp ANTENNA_2477 (.A(net75));
 sg13g2_antennanp ANTENNA_2478 (.A(net75));
 sg13g2_antennanp ANTENNA_2479 (.A(net75));
 sg13g2_antennanp ANTENNA_2480 (.A(net75));
 sg13g2_antennanp ANTENNA_2481 (.A(net75));
 sg13g2_antennanp ANTENNA_2482 (.A(net75));
 sg13g2_antennanp ANTENNA_2483 (.A(net75));
 sg13g2_antennanp ANTENNA_2484 (.A(net75));
 sg13g2_antennanp ANTENNA_2485 (.A(net79));
 sg13g2_antennanp ANTENNA_2486 (.A(net79));
 sg13g2_antennanp ANTENNA_2487 (.A(net79));
 sg13g2_antennanp ANTENNA_2488 (.A(net79));
 sg13g2_antennanp ANTENNA_2489 (.A(net79));
 sg13g2_antennanp ANTENNA_2490 (.A(net79));
 sg13g2_antennanp ANTENNA_2491 (.A(net79));
 sg13g2_antennanp ANTENNA_2492 (.A(net79));
 sg13g2_antennanp ANTENNA_2493 (.A(net82));
 sg13g2_antennanp ANTENNA_2494 (.A(net82));
 sg13g2_antennanp ANTENNA_2495 (.A(net82));
 sg13g2_antennanp ANTENNA_2496 (.A(net82));
 sg13g2_antennanp ANTENNA_2497 (.A(net82));
 sg13g2_antennanp ANTENNA_2498 (.A(net82));
 sg13g2_antennanp ANTENNA_2499 (.A(net82));
 sg13g2_antennanp ANTENNA_2500 (.A(net82));
 sg13g2_antennanp ANTENNA_2501 (.A(net82));
 sg13g2_antennanp ANTENNA_2502 (.A(net82));
 sg13g2_antennanp ANTENNA_2503 (.A(net82));
 sg13g2_antennanp ANTENNA_2504 (.A(net82));
 sg13g2_antennanp ANTENNA_2505 (.A(net82));
 sg13g2_antennanp ANTENNA_2506 (.A(net103));
 sg13g2_antennanp ANTENNA_2507 (.A(net103));
 sg13g2_antennanp ANTENNA_2508 (.A(net103));
 sg13g2_antennanp ANTENNA_2509 (.A(net103));
 sg13g2_antennanp ANTENNA_2510 (.A(net103));
 sg13g2_antennanp ANTENNA_2511 (.A(net103));
 sg13g2_antennanp ANTENNA_2512 (.A(net103));
 sg13g2_antennanp ANTENNA_2513 (.A(net103));
 sg13g2_antennanp ANTENNA_2514 (.A(net107));
 sg13g2_antennanp ANTENNA_2515 (.A(net107));
 sg13g2_antennanp ANTENNA_2516 (.A(net107));
 sg13g2_antennanp ANTENNA_2517 (.A(net107));
 sg13g2_antennanp ANTENNA_2518 (.A(net107));
 sg13g2_antennanp ANTENNA_2519 (.A(net107));
 sg13g2_antennanp ANTENNA_2520 (.A(net107));
 sg13g2_antennanp ANTENNA_2521 (.A(net107));
 sg13g2_antennanp ANTENNA_2522 (.A(net107));
 sg13g2_antennanp ANTENNA_2523 (.A(net107));
 sg13g2_antennanp ANTENNA_2524 (.A(net107));
 sg13g2_antennanp ANTENNA_2525 (.A(net107));
 sg13g2_antennanp ANTENNA_2526 (.A(net107));
 sg13g2_antennanp ANTENNA_2527 (.A(net107));
 sg13g2_antennanp ANTENNA_2528 (.A(net107));
 sg13g2_antennanp ANTENNA_2529 (.A(net108));
 sg13g2_antennanp ANTENNA_2530 (.A(net108));
 sg13g2_antennanp ANTENNA_2531 (.A(net108));
 sg13g2_antennanp ANTENNA_2532 (.A(net108));
 sg13g2_antennanp ANTENNA_2533 (.A(net108));
 sg13g2_antennanp ANTENNA_2534 (.A(net108));
 sg13g2_antennanp ANTENNA_2535 (.A(net108));
 sg13g2_antennanp ANTENNA_2536 (.A(net108));
 sg13g2_antennanp ANTENNA_2537 (.A(net108));
 sg13g2_antennanp ANTENNA_2538 (.A(net108));
 sg13g2_antennanp ANTENNA_2539 (.A(net108));
 sg13g2_antennanp ANTENNA_2540 (.A(net108));
 sg13g2_antennanp ANTENNA_2541 (.A(net108));
 sg13g2_antennanp ANTENNA_2542 (.A(net108));
 sg13g2_antennanp ANTENNA_2543 (.A(net108));
 sg13g2_antennanp ANTENNA_2544 (.A(net108));
 sg13g2_antennanp ANTENNA_2545 (.A(net108));
 sg13g2_antennanp ANTENNA_2546 (.A(net108));
 sg13g2_antennanp ANTENNA_2547 (.A(net108));
 sg13g2_antennanp ANTENNA_2548 (.A(net108));
 sg13g2_antennanp ANTENNA_2549 (.A(net108));
 sg13g2_antennanp ANTENNA_2550 (.A(net108));
 sg13g2_antennanp ANTENNA_2551 (.A(net108));
 sg13g2_antennanp ANTENNA_2552 (.A(net108));
 sg13g2_antennanp ANTENNA_2553 (.A(net108));
 sg13g2_antennanp ANTENNA_2554 (.A(net108));
 sg13g2_antennanp ANTENNA_2555 (.A(net108));
 sg13g2_antennanp ANTENNA_2556 (.A(net108));
 sg13g2_antennanp ANTENNA_2557 (.A(net108));
 sg13g2_antennanp ANTENNA_2558 (.A(net108));
 sg13g2_antennanp ANTENNA_2559 (.A(net108));
 sg13g2_antennanp ANTENNA_2560 (.A(net108));
 sg13g2_antennanp ANTENNA_2561 (.A(net108));
 sg13g2_antennanp ANTENNA_2562 (.A(net108));
 sg13g2_antennanp ANTENNA_2563 (.A(net108));
 sg13g2_antennanp ANTENNA_2564 (.A(net108));
 sg13g2_antennanp ANTENNA_2565 (.A(net113));
 sg13g2_antennanp ANTENNA_2566 (.A(net113));
 sg13g2_antennanp ANTENNA_2567 (.A(net113));
 sg13g2_antennanp ANTENNA_2568 (.A(net113));
 sg13g2_antennanp ANTENNA_2569 (.A(net113));
 sg13g2_antennanp ANTENNA_2570 (.A(net113));
 sg13g2_antennanp ANTENNA_2571 (.A(net113));
 sg13g2_antennanp ANTENNA_2572 (.A(net113));
 sg13g2_antennanp ANTENNA_2573 (.A(net113));
 sg13g2_antennanp ANTENNA_2574 (.A(net113));
 sg13g2_antennanp ANTENNA_2575 (.A(net113));
 sg13g2_antennanp ANTENNA_2576 (.A(net113));
 sg13g2_antennanp ANTENNA_2577 (.A(net113));
 sg13g2_antennanp ANTENNA_2578 (.A(net113));
 sg13g2_antennanp ANTENNA_2579 (.A(net113));
 sg13g2_antennanp ANTENNA_2580 (.A(net118));
 sg13g2_antennanp ANTENNA_2581 (.A(net118));
 sg13g2_antennanp ANTENNA_2582 (.A(net118));
 sg13g2_antennanp ANTENNA_2583 (.A(net118));
 sg13g2_antennanp ANTENNA_2584 (.A(net118));
 sg13g2_antennanp ANTENNA_2585 (.A(net118));
 sg13g2_antennanp ANTENNA_2586 (.A(net118));
 sg13g2_antennanp ANTENNA_2587 (.A(net118));
 sg13g2_antennanp ANTENNA_2588 (.A(net124));
 sg13g2_antennanp ANTENNA_2589 (.A(net124));
 sg13g2_antennanp ANTENNA_2590 (.A(net124));
 sg13g2_antennanp ANTENNA_2591 (.A(net124));
 sg13g2_antennanp ANTENNA_2592 (.A(net124));
 sg13g2_antennanp ANTENNA_2593 (.A(net124));
 sg13g2_antennanp ANTENNA_2594 (.A(net124));
 sg13g2_antennanp ANTENNA_2595 (.A(net124));
 sg13g2_antennanp ANTENNA_2596 (.A(net124));
 sg13g2_antennanp ANTENNA_2597 (.A(net124));
 sg13g2_antennanp ANTENNA_2598 (.A(net124));
 sg13g2_antennanp ANTENNA_2599 (.A(net124));
 sg13g2_antennanp ANTENNA_2600 (.A(net124));
 sg13g2_antennanp ANTENNA_2601 (.A(net125));
 sg13g2_antennanp ANTENNA_2602 (.A(net125));
 sg13g2_antennanp ANTENNA_2603 (.A(net125));
 sg13g2_antennanp ANTENNA_2604 (.A(net125));
 sg13g2_antennanp ANTENNA_2605 (.A(net125));
 sg13g2_antennanp ANTENNA_2606 (.A(net125));
 sg13g2_antennanp ANTENNA_2607 (.A(net125));
 sg13g2_antennanp ANTENNA_2608 (.A(net125));
 sg13g2_antennanp ANTENNA_2609 (.A(net127));
 sg13g2_antennanp ANTENNA_2610 (.A(net127));
 sg13g2_antennanp ANTENNA_2611 (.A(net127));
 sg13g2_antennanp ANTENNA_2612 (.A(net127));
 sg13g2_antennanp ANTENNA_2613 (.A(net127));
 sg13g2_antennanp ANTENNA_2614 (.A(net127));
 sg13g2_antennanp ANTENNA_2615 (.A(net127));
 sg13g2_antennanp ANTENNA_2616 (.A(net127));
 sg13g2_antennanp ANTENNA_2617 (.A(net127));
 sg13g2_antennanp ANTENNA_2618 (.A(net127));
 sg13g2_antennanp ANTENNA_2619 (.A(net127));
 sg13g2_antennanp ANTENNA_2620 (.A(net127));
 sg13g2_antennanp ANTENNA_2621 (.A(net127));
 sg13g2_antennanp ANTENNA_2622 (.A(net127));
 sg13g2_antennanp ANTENNA_2623 (.A(net127));
 sg13g2_antennanp ANTENNA_2624 (.A(net127));
 sg13g2_antennanp ANTENNA_2625 (.A(net127));
 sg13g2_antennanp ANTENNA_2626 (.A(net127));
 sg13g2_antennanp ANTENNA_2627 (.A(net127));
 sg13g2_antennanp ANTENNA_2628 (.A(net127));
 sg13g2_antennanp ANTENNA_2629 (.A(net127));
 sg13g2_antennanp ANTENNA_2630 (.A(net368));
 sg13g2_antennanp ANTENNA_2631 (.A(net368));
 sg13g2_antennanp ANTENNA_2632 (.A(net368));
 sg13g2_antennanp ANTENNA_2633 (.A(net368));
 sg13g2_antennanp ANTENNA_2634 (.A(net368));
 sg13g2_antennanp ANTENNA_2635 (.A(net368));
 sg13g2_antennanp ANTENNA_2636 (.A(net368));
 sg13g2_antennanp ANTENNA_2637 (.A(net368));
 sg13g2_antennanp ANTENNA_2638 (.A(net368));
 sg13g2_antennanp ANTENNA_2639 (.A(net368));
 sg13g2_antennanp ANTENNA_2640 (.A(net368));
 sg13g2_antennanp ANTENNA_2641 (.A(net368));
 sg13g2_antennanp ANTENNA_2642 (.A(net368));
 sg13g2_antennanp ANTENNA_2643 (.A(net368));
 sg13g2_antennanp ANTENNA_2644 (.A(net368));
 sg13g2_antennanp ANTENNA_2645 (.A(net368));
 sg13g2_antennanp ANTENNA_2646 (.A(net368));
 sg13g2_antennanp ANTENNA_2647 (.A(net368));
 sg13g2_antennanp ANTENNA_2648 (.A(net368));
 sg13g2_antennanp ANTENNA_2649 (.A(net368));
 sg13g2_antennanp ANTENNA_2650 (.A(net368));
 sg13g2_antennanp ANTENNA_2651 (.A(net368));
 sg13g2_antennanp ANTENNA_2652 (.A(net368));
 sg13g2_antennanp ANTENNA_2653 (.A(net368));
 sg13g2_antennanp ANTENNA_2654 (.A(net386));
 sg13g2_antennanp ANTENNA_2655 (.A(net386));
 sg13g2_antennanp ANTENNA_2656 (.A(net386));
 sg13g2_antennanp ANTENNA_2657 (.A(net386));
 sg13g2_antennanp ANTENNA_2658 (.A(net386));
 sg13g2_antennanp ANTENNA_2659 (.A(net386));
 sg13g2_antennanp ANTENNA_2660 (.A(net386));
 sg13g2_antennanp ANTENNA_2661 (.A(net386));
 sg13g2_antennanp ANTENNA_2662 (.A(net386));
 sg13g2_antennanp ANTENNA_2663 (.A(net386));
 sg13g2_antennanp ANTENNA_2664 (.A(net386));
 sg13g2_antennanp ANTENNA_2665 (.A(net386));
 sg13g2_antennanp ANTENNA_2666 (.A(net386));
 sg13g2_antennanp ANTENNA_2667 (.A(net386));
 sg13g2_antennanp ANTENNA_2668 (.A(net386));
 sg13g2_antennanp ANTENNA_2669 (.A(net386));
 sg13g2_antennanp ANTENNA_2670 (.A(net386));
 sg13g2_antennanp ANTENNA_2671 (.A(net1002));
 sg13g2_antennanp ANTENNA_2672 (.A(net1002));
 sg13g2_antennanp ANTENNA_2673 (.A(net1002));
 sg13g2_antennanp ANTENNA_2674 (.A(net1002));
 sg13g2_antennanp ANTENNA_2675 (.A(net1002));
 sg13g2_antennanp ANTENNA_2676 (.A(net1002));
 sg13g2_antennanp ANTENNA_2677 (.A(net1002));
 sg13g2_antennanp ANTENNA_2678 (.A(net1002));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_fill_1 FILLER_0_266 ();
 sg13g2_decap_4 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_4 FILLER_0_300 ();
 sg13g2_fill_2 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_fill_1 FILLER_0_371 ();
 sg13g2_fill_2 FILLER_0_377 ();
 sg13g2_fill_1 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_4 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_decap_8 FILLER_0_449 ();
 sg13g2_fill_2 FILLER_0_456 ();
 sg13g2_decap_8 FILLER_0_466 ();
 sg13g2_fill_1 FILLER_0_497 ();
 sg13g2_fill_1 FILLER_0_506 ();
 sg13g2_decap_8 FILLER_0_537 ();
 sg13g2_decap_8 FILLER_0_544 ();
 sg13g2_decap_8 FILLER_0_551 ();
 sg13g2_decap_8 FILLER_0_558 ();
 sg13g2_decap_8 FILLER_0_565 ();
 sg13g2_decap_8 FILLER_0_572 ();
 sg13g2_decap_4 FILLER_0_579 ();
 sg13g2_fill_2 FILLER_0_583 ();
 sg13g2_decap_8 FILLER_0_601 ();
 sg13g2_decap_8 FILLER_0_608 ();
 sg13g2_decap_8 FILLER_0_615 ();
 sg13g2_decap_8 FILLER_0_622 ();
 sg13g2_decap_8 FILLER_0_629 ();
 sg13g2_decap_8 FILLER_0_636 ();
 sg13g2_decap_8 FILLER_0_643 ();
 sg13g2_fill_2 FILLER_0_650 ();
 sg13g2_fill_1 FILLER_0_652 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_671 ();
 sg13g2_decap_4 FILLER_0_678 ();
 sg13g2_fill_2 FILLER_0_682 ();
 sg13g2_decap_8 FILLER_0_688 ();
 sg13g2_decap_4 FILLER_0_695 ();
 sg13g2_decap_8 FILLER_0_704 ();
 sg13g2_decap_8 FILLER_0_711 ();
 sg13g2_decap_8 FILLER_0_718 ();
 sg13g2_fill_2 FILLER_0_725 ();
 sg13g2_fill_1 FILLER_0_727 ();
 sg13g2_fill_2 FILLER_0_732 ();
 sg13g2_decap_8 FILLER_0_739 ();
 sg13g2_decap_8 FILLER_0_746 ();
 sg13g2_decap_8 FILLER_0_753 ();
 sg13g2_fill_1 FILLER_0_760 ();
 sg13g2_decap_4 FILLER_0_775 ();
 sg13g2_fill_1 FILLER_0_779 ();
 sg13g2_fill_2 FILLER_0_795 ();
 sg13g2_fill_1 FILLER_0_797 ();
 sg13g2_fill_1 FILLER_0_802 ();
 sg13g2_fill_2 FILLER_0_808 ();
 sg13g2_fill_1 FILLER_0_810 ();
 sg13g2_fill_2 FILLER_0_823 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_fill_2 FILLER_0_843 ();
 sg13g2_fill_1 FILLER_0_845 ();
 sg13g2_decap_4 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_880 ();
 sg13g2_fill_2 FILLER_0_887 ();
 sg13g2_fill_1 FILLER_0_889 ();
 sg13g2_decap_4 FILLER_0_894 ();
 sg13g2_fill_2 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_4 FILLER_0_929 ();
 sg13g2_decap_4 FILLER_0_937 ();
 sg13g2_fill_1 FILLER_0_941 ();
 sg13g2_decap_4 FILLER_0_946 ();
 sg13g2_fill_1 FILLER_0_950 ();
 sg13g2_decap_8 FILLER_0_981 ();
 sg13g2_decap_8 FILLER_0_988 ();
 sg13g2_decap_4 FILLER_0_995 ();
 sg13g2_decap_8 FILLER_0_1003 ();
 sg13g2_decap_8 FILLER_0_1023 ();
 sg13g2_decap_8 FILLER_0_1030 ();
 sg13g2_decap_8 FILLER_0_1037 ();
 sg13g2_decap_4 FILLER_0_1049 ();
 sg13g2_decap_8 FILLER_0_1079 ();
 sg13g2_decap_8 FILLER_0_1086 ();
 sg13g2_decap_8 FILLER_0_1093 ();
 sg13g2_decap_8 FILLER_0_1100 ();
 sg13g2_decap_8 FILLER_0_1107 ();
 sg13g2_fill_2 FILLER_0_1114 ();
 sg13g2_fill_1 FILLER_0_1125 ();
 sg13g2_decap_8 FILLER_0_1130 ();
 sg13g2_decap_8 FILLER_0_1150 ();
 sg13g2_decap_8 FILLER_0_1157 ();
 sg13g2_decap_8 FILLER_0_1164 ();
 sg13g2_decap_8 FILLER_0_1171 ();
 sg13g2_decap_8 FILLER_0_1178 ();
 sg13g2_fill_1 FILLER_0_1185 ();
 sg13g2_decap_8 FILLER_0_1212 ();
 sg13g2_decap_8 FILLER_0_1219 ();
 sg13g2_decap_8 FILLER_0_1226 ();
 sg13g2_decap_8 FILLER_0_1233 ();
 sg13g2_decap_8 FILLER_0_1240 ();
 sg13g2_decap_4 FILLER_0_1247 ();
 sg13g2_decap_8 FILLER_0_1255 ();
 sg13g2_decap_8 FILLER_0_1262 ();
 sg13g2_decap_8 FILLER_0_1269 ();
 sg13g2_decap_8 FILLER_0_1276 ();
 sg13g2_decap_8 FILLER_0_1283 ();
 sg13g2_decap_8 FILLER_0_1290 ();
 sg13g2_decap_8 FILLER_0_1297 ();
 sg13g2_decap_8 FILLER_0_1304 ();
 sg13g2_decap_8 FILLER_0_1311 ();
 sg13g2_decap_8 FILLER_0_1318 ();
 sg13g2_decap_8 FILLER_0_1325 ();
 sg13g2_decap_8 FILLER_0_1332 ();
 sg13g2_decap_8 FILLER_0_1339 ();
 sg13g2_decap_8 FILLER_0_1346 ();
 sg13g2_decap_8 FILLER_0_1353 ();
 sg13g2_decap_8 FILLER_0_1360 ();
 sg13g2_decap_8 FILLER_0_1367 ();
 sg13g2_decap_8 FILLER_0_1374 ();
 sg13g2_decap_8 FILLER_0_1381 ();
 sg13g2_decap_8 FILLER_0_1388 ();
 sg13g2_decap_8 FILLER_0_1395 ();
 sg13g2_decap_8 FILLER_0_1402 ();
 sg13g2_decap_8 FILLER_0_1409 ();
 sg13g2_decap_8 FILLER_0_1416 ();
 sg13g2_decap_8 FILLER_0_1423 ();
 sg13g2_decap_8 FILLER_0_1430 ();
 sg13g2_decap_8 FILLER_0_1437 ();
 sg13g2_decap_8 FILLER_0_1444 ();
 sg13g2_decap_8 FILLER_0_1451 ();
 sg13g2_decap_8 FILLER_0_1458 ();
 sg13g2_decap_8 FILLER_0_1465 ();
 sg13g2_decap_8 FILLER_0_1472 ();
 sg13g2_decap_8 FILLER_0_1479 ();
 sg13g2_decap_8 FILLER_0_1486 ();
 sg13g2_decap_8 FILLER_0_1493 ();
 sg13g2_decap_8 FILLER_0_1500 ();
 sg13g2_decap_8 FILLER_0_1507 ();
 sg13g2_decap_8 FILLER_0_1514 ();
 sg13g2_decap_8 FILLER_0_1521 ();
 sg13g2_decap_8 FILLER_0_1528 ();
 sg13g2_decap_8 FILLER_0_1535 ();
 sg13g2_decap_8 FILLER_0_1542 ();
 sg13g2_decap_8 FILLER_0_1549 ();
 sg13g2_decap_8 FILLER_0_1556 ();
 sg13g2_decap_8 FILLER_0_1563 ();
 sg13g2_decap_8 FILLER_0_1570 ();
 sg13g2_decap_8 FILLER_0_1577 ();
 sg13g2_decap_8 FILLER_0_1584 ();
 sg13g2_decap_8 FILLER_0_1591 ();
 sg13g2_decap_8 FILLER_0_1598 ();
 sg13g2_decap_8 FILLER_0_1605 ();
 sg13g2_decap_8 FILLER_0_1612 ();
 sg13g2_decap_8 FILLER_0_1619 ();
 sg13g2_decap_8 FILLER_0_1626 ();
 sg13g2_decap_8 FILLER_0_1633 ();
 sg13g2_decap_8 FILLER_0_1640 ();
 sg13g2_decap_8 FILLER_0_1647 ();
 sg13g2_decap_8 FILLER_0_1654 ();
 sg13g2_decap_8 FILLER_0_1661 ();
 sg13g2_decap_8 FILLER_0_1668 ();
 sg13g2_decap_8 FILLER_0_1675 ();
 sg13g2_decap_8 FILLER_0_1682 ();
 sg13g2_decap_8 FILLER_0_1689 ();
 sg13g2_decap_8 FILLER_0_1696 ();
 sg13g2_decap_8 FILLER_0_1703 ();
 sg13g2_decap_8 FILLER_0_1710 ();
 sg13g2_decap_8 FILLER_0_1717 ();
 sg13g2_decap_8 FILLER_0_1724 ();
 sg13g2_decap_8 FILLER_0_1731 ();
 sg13g2_decap_8 FILLER_0_1738 ();
 sg13g2_decap_8 FILLER_0_1745 ();
 sg13g2_decap_8 FILLER_0_1752 ();
 sg13g2_decap_8 FILLER_0_1759 ();
 sg13g2_decap_8 FILLER_0_1766 ();
 sg13g2_fill_1 FILLER_0_1773 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_4 FILLER_1_333 ();
 sg13g2_fill_1 FILLER_1_337 ();
 sg13g2_decap_4 FILLER_1_351 ();
 sg13g2_fill_1 FILLER_1_355 ();
 sg13g2_fill_1 FILLER_1_361 ();
 sg13g2_fill_1 FILLER_1_382 ();
 sg13g2_decap_4 FILLER_1_387 ();
 sg13g2_fill_1 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_4 FILLER_1_404 ();
 sg13g2_fill_2 FILLER_1_408 ();
 sg13g2_decap_4 FILLER_1_421 ();
 sg13g2_fill_1 FILLER_1_425 ();
 sg13g2_decap_8 FILLER_1_431 ();
 sg13g2_decap_8 FILLER_1_438 ();
 sg13g2_fill_2 FILLER_1_492 ();
 sg13g2_fill_1 FILLER_1_494 ();
 sg13g2_decap_4 FILLER_1_502 ();
 sg13g2_fill_1 FILLER_1_506 ();
 sg13g2_decap_4 FILLER_1_510 ();
 sg13g2_decap_8 FILLER_1_522 ();
 sg13g2_decap_4 FILLER_1_537 ();
 sg13g2_fill_1 FILLER_1_541 ();
 sg13g2_decap_8 FILLER_1_550 ();
 sg13g2_fill_2 FILLER_1_557 ();
 sg13g2_decap_4 FILLER_1_569 ();
 sg13g2_fill_2 FILLER_1_577 ();
 sg13g2_fill_1 FILLER_1_579 ();
 sg13g2_fill_2 FILLER_1_613 ();
 sg13g2_fill_1 FILLER_1_615 ();
 sg13g2_fill_1 FILLER_1_621 ();
 sg13g2_fill_2 FILLER_1_626 ();
 sg13g2_fill_2 FILLER_1_632 ();
 sg13g2_fill_1 FILLER_1_634 ();
 sg13g2_fill_1 FILLER_1_643 ();
 sg13g2_decap_4 FILLER_1_675 ();
 sg13g2_fill_2 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_4 FILLER_1_707 ();
 sg13g2_fill_2 FILLER_1_714 ();
 sg13g2_fill_1 FILLER_1_716 ();
 sg13g2_fill_1 FILLER_1_721 ();
 sg13g2_fill_1 FILLER_1_734 ();
 sg13g2_fill_1 FILLER_1_739 ();
 sg13g2_fill_1 FILLER_1_744 ();
 sg13g2_decap_4 FILLER_1_775 ();
 sg13g2_decap_4 FILLER_1_794 ();
 sg13g2_fill_2 FILLER_1_798 ();
 sg13g2_fill_1 FILLER_1_821 ();
 sg13g2_fill_2 FILLER_1_827 ();
 sg13g2_decap_8 FILLER_1_839 ();
 sg13g2_decap_8 FILLER_1_846 ();
 sg13g2_decap_8 FILLER_1_853 ();
 sg13g2_fill_1 FILLER_1_864 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_fill_2 FILLER_1_889 ();
 sg13g2_fill_2 FILLER_1_900 ();
 sg13g2_fill_1 FILLER_1_917 ();
 sg13g2_fill_1 FILLER_1_929 ();
 sg13g2_fill_1 FILLER_1_935 ();
 sg13g2_fill_2 FILLER_1_949 ();
 sg13g2_fill_1 FILLER_1_951 ();
 sg13g2_decap_4 FILLER_1_956 ();
 sg13g2_fill_2 FILLER_1_973 ();
 sg13g2_fill_1 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_986 ();
 sg13g2_decap_4 FILLER_1_993 ();
 sg13g2_fill_2 FILLER_1_1025 ();
 sg13g2_fill_2 FILLER_1_1050 ();
 sg13g2_decap_4 FILLER_1_1064 ();
 sg13g2_fill_2 FILLER_1_1068 ();
 sg13g2_decap_4 FILLER_1_1074 ();
 sg13g2_fill_1 FILLER_1_1082 ();
 sg13g2_fill_2 FILLER_1_1145 ();
 sg13g2_fill_1 FILLER_1_1147 ();
 sg13g2_fill_2 FILLER_1_1153 ();
 sg13g2_fill_1 FILLER_1_1155 ();
 sg13g2_decap_8 FILLER_1_1161 ();
 sg13g2_decap_8 FILLER_1_1176 ();
 sg13g2_fill_1 FILLER_1_1183 ();
 sg13g2_decap_4 FILLER_1_1188 ();
 sg13g2_fill_2 FILLER_1_1192 ();
 sg13g2_fill_2 FILLER_1_1198 ();
 sg13g2_fill_1 FILLER_1_1200 ();
 sg13g2_decap_4 FILLER_1_1205 ();
 sg13g2_fill_2 FILLER_1_1217 ();
 sg13g2_fill_1 FILLER_1_1219 ();
 sg13g2_decap_8 FILLER_1_1224 ();
 sg13g2_decap_8 FILLER_1_1231 ();
 sg13g2_decap_8 FILLER_1_1238 ();
 sg13g2_fill_1 FILLER_1_1245 ();
 sg13g2_decap_8 FILLER_1_1264 ();
 sg13g2_decap_8 FILLER_1_1271 ();
 sg13g2_decap_8 FILLER_1_1278 ();
 sg13g2_decap_4 FILLER_1_1285 ();
 sg13g2_fill_2 FILLER_1_1289 ();
 sg13g2_decap_8 FILLER_1_1317 ();
 sg13g2_decap_8 FILLER_1_1324 ();
 sg13g2_decap_8 FILLER_1_1331 ();
 sg13g2_decap_8 FILLER_1_1338 ();
 sg13g2_decap_8 FILLER_1_1345 ();
 sg13g2_decap_8 FILLER_1_1352 ();
 sg13g2_decap_8 FILLER_1_1359 ();
 sg13g2_decap_8 FILLER_1_1366 ();
 sg13g2_decap_8 FILLER_1_1373 ();
 sg13g2_decap_8 FILLER_1_1380 ();
 sg13g2_decap_8 FILLER_1_1387 ();
 sg13g2_decap_8 FILLER_1_1394 ();
 sg13g2_decap_8 FILLER_1_1401 ();
 sg13g2_decap_8 FILLER_1_1408 ();
 sg13g2_decap_8 FILLER_1_1415 ();
 sg13g2_decap_8 FILLER_1_1422 ();
 sg13g2_decap_8 FILLER_1_1429 ();
 sg13g2_decap_8 FILLER_1_1436 ();
 sg13g2_decap_8 FILLER_1_1443 ();
 sg13g2_decap_8 FILLER_1_1450 ();
 sg13g2_decap_8 FILLER_1_1457 ();
 sg13g2_decap_8 FILLER_1_1464 ();
 sg13g2_decap_8 FILLER_1_1471 ();
 sg13g2_decap_8 FILLER_1_1478 ();
 sg13g2_decap_8 FILLER_1_1485 ();
 sg13g2_decap_8 FILLER_1_1492 ();
 sg13g2_decap_8 FILLER_1_1499 ();
 sg13g2_decap_8 FILLER_1_1506 ();
 sg13g2_decap_8 FILLER_1_1513 ();
 sg13g2_decap_8 FILLER_1_1520 ();
 sg13g2_decap_8 FILLER_1_1527 ();
 sg13g2_decap_8 FILLER_1_1534 ();
 sg13g2_decap_8 FILLER_1_1541 ();
 sg13g2_decap_8 FILLER_1_1548 ();
 sg13g2_decap_8 FILLER_1_1555 ();
 sg13g2_decap_8 FILLER_1_1562 ();
 sg13g2_decap_8 FILLER_1_1569 ();
 sg13g2_decap_8 FILLER_1_1576 ();
 sg13g2_decap_8 FILLER_1_1583 ();
 sg13g2_decap_8 FILLER_1_1590 ();
 sg13g2_decap_8 FILLER_1_1597 ();
 sg13g2_decap_8 FILLER_1_1604 ();
 sg13g2_decap_8 FILLER_1_1611 ();
 sg13g2_decap_8 FILLER_1_1618 ();
 sg13g2_decap_8 FILLER_1_1625 ();
 sg13g2_decap_8 FILLER_1_1632 ();
 sg13g2_decap_8 FILLER_1_1639 ();
 sg13g2_decap_8 FILLER_1_1646 ();
 sg13g2_decap_8 FILLER_1_1653 ();
 sg13g2_decap_8 FILLER_1_1660 ();
 sg13g2_decap_8 FILLER_1_1667 ();
 sg13g2_decap_8 FILLER_1_1674 ();
 sg13g2_decap_8 FILLER_1_1681 ();
 sg13g2_decap_8 FILLER_1_1688 ();
 sg13g2_decap_8 FILLER_1_1695 ();
 sg13g2_decap_8 FILLER_1_1702 ();
 sg13g2_decap_8 FILLER_1_1709 ();
 sg13g2_decap_8 FILLER_1_1716 ();
 sg13g2_decap_8 FILLER_1_1723 ();
 sg13g2_decap_8 FILLER_1_1730 ();
 sg13g2_decap_8 FILLER_1_1737 ();
 sg13g2_decap_8 FILLER_1_1744 ();
 sg13g2_decap_8 FILLER_1_1751 ();
 sg13g2_decap_8 FILLER_1_1758 ();
 sg13g2_decap_8 FILLER_1_1765 ();
 sg13g2_fill_2 FILLER_1_1772 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_4 FILLER_2_196 ();
 sg13g2_fill_2 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_4 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_226 ();
 sg13g2_fill_1 FILLER_2_233 ();
 sg13g2_decap_4 FILLER_2_243 ();
 sg13g2_fill_1 FILLER_2_247 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_fill_1 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_4 FILLER_2_293 ();
 sg13g2_fill_2 FILLER_2_297 ();
 sg13g2_decap_8 FILLER_2_303 ();
 sg13g2_fill_2 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_fill_2 FILLER_2_333 ();
 sg13g2_decap_4 FILLER_2_339 ();
 sg13g2_fill_2 FILLER_2_343 ();
 sg13g2_fill_2 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_4 FILLER_2_368 ();
 sg13g2_fill_1 FILLER_2_372 ();
 sg13g2_fill_2 FILLER_2_378 ();
 sg13g2_decap_4 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_fill_2 FILLER_2_424 ();
 sg13g2_fill_2 FILLER_2_430 ();
 sg13g2_fill_1 FILLER_2_432 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_4 FILLER_2_445 ();
 sg13g2_fill_1 FILLER_2_449 ();
 sg13g2_fill_1 FILLER_2_454 ();
 sg13g2_fill_2 FILLER_2_460 ();
 sg13g2_decap_4 FILLER_2_488 ();
 sg13g2_fill_1 FILLER_2_492 ();
 sg13g2_decap_8 FILLER_2_508 ();
 sg13g2_fill_2 FILLER_2_515 ();
 sg13g2_decap_4 FILLER_2_526 ();
 sg13g2_fill_2 FILLER_2_530 ();
 sg13g2_decap_4 FILLER_2_537 ();
 sg13g2_fill_1 FILLER_2_541 ();
 sg13g2_fill_2 FILLER_2_547 ();
 sg13g2_fill_1 FILLER_2_549 ();
 sg13g2_decap_8 FILLER_2_559 ();
 sg13g2_fill_1 FILLER_2_566 ();
 sg13g2_fill_2 FILLER_2_572 ();
 sg13g2_fill_2 FILLER_2_594 ();
 sg13g2_fill_2 FILLER_2_604 ();
 sg13g2_fill_1 FILLER_2_606 ();
 sg13g2_fill_2 FILLER_2_626 ();
 sg13g2_fill_2 FILLER_2_639 ();
 sg13g2_fill_1 FILLER_2_641 ();
 sg13g2_fill_1 FILLER_2_647 ();
 sg13g2_fill_1 FILLER_2_652 ();
 sg13g2_decap_4 FILLER_2_662 ();
 sg13g2_fill_2 FILLER_2_666 ();
 sg13g2_decap_4 FILLER_2_672 ();
 sg13g2_fill_2 FILLER_2_680 ();
 sg13g2_fill_1 FILLER_2_686 ();
 sg13g2_fill_1 FILLER_2_691 ();
 sg13g2_fill_1 FILLER_2_696 ();
 sg13g2_fill_1 FILLER_2_702 ();
 sg13g2_fill_2 FILLER_2_708 ();
 sg13g2_fill_2 FILLER_2_715 ();
 sg13g2_fill_2 FILLER_2_723 ();
 sg13g2_decap_8 FILLER_2_730 ();
 sg13g2_decap_8 FILLER_2_737 ();
 sg13g2_decap_8 FILLER_2_744 ();
 sg13g2_decap_4 FILLER_2_751 ();
 sg13g2_fill_1 FILLER_2_755 ();
 sg13g2_decap_4 FILLER_2_760 ();
 sg13g2_fill_2 FILLER_2_764 ();
 sg13g2_fill_1 FILLER_2_781 ();
 sg13g2_fill_2 FILLER_2_787 ();
 sg13g2_fill_2 FILLER_2_794 ();
 sg13g2_fill_1 FILLER_2_839 ();
 sg13g2_decap_8 FILLER_2_852 ();
 sg13g2_fill_1 FILLER_2_859 ();
 sg13g2_fill_2 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_2_883 ();
 sg13g2_decap_8 FILLER_2_894 ();
 sg13g2_fill_2 FILLER_2_901 ();
 sg13g2_fill_1 FILLER_2_903 ();
 sg13g2_fill_1 FILLER_2_934 ();
 sg13g2_fill_1 FILLER_2_939 ();
 sg13g2_fill_1 FILLER_2_946 ();
 sg13g2_fill_1 FILLER_2_952 ();
 sg13g2_decap_4 FILLER_2_980 ();
 sg13g2_fill_1 FILLER_2_984 ();
 sg13g2_decap_4 FILLER_2_989 ();
 sg13g2_fill_2 FILLER_2_993 ();
 sg13g2_decap_4 FILLER_2_999 ();
 sg13g2_fill_1 FILLER_2_1008 ();
 sg13g2_fill_1 FILLER_2_1018 ();
 sg13g2_fill_1 FILLER_2_1024 ();
 sg13g2_fill_1 FILLER_2_1034 ();
 sg13g2_decap_8 FILLER_2_1052 ();
 sg13g2_decap_8 FILLER_2_1059 ();
 sg13g2_decap_8 FILLER_2_1066 ();
 sg13g2_fill_2 FILLER_2_1073 ();
 sg13g2_fill_1 FILLER_2_1075 ();
 sg13g2_fill_1 FILLER_2_1081 ();
 sg13g2_decap_8 FILLER_2_1095 ();
 sg13g2_decap_8 FILLER_2_1102 ();
 sg13g2_fill_1 FILLER_2_1121 ();
 sg13g2_fill_2 FILLER_2_1125 ();
 sg13g2_fill_1 FILLER_2_1127 ();
 sg13g2_fill_2 FILLER_2_1139 ();
 sg13g2_fill_1 FILLER_2_1141 ();
 sg13g2_decap_8 FILLER_2_1150 ();
 sg13g2_fill_2 FILLER_2_1157 ();
 sg13g2_fill_1 FILLER_2_1159 ();
 sg13g2_decap_4 FILLER_2_1167 ();
 sg13g2_decap_4 FILLER_2_1176 ();
 sg13g2_fill_1 FILLER_2_1184 ();
 sg13g2_fill_2 FILLER_2_1189 ();
 sg13g2_fill_1 FILLER_2_1200 ();
 sg13g2_fill_1 FILLER_2_1219 ();
 sg13g2_decap_4 FILLER_2_1256 ();
 sg13g2_fill_1 FILLER_2_1260 ();
 sg13g2_decap_8 FILLER_2_1265 ();
 sg13g2_decap_8 FILLER_2_1272 ();
 sg13g2_decap_8 FILLER_2_1279 ();
 sg13g2_decap_8 FILLER_2_1286 ();
 sg13g2_fill_1 FILLER_2_1293 ();
 sg13g2_fill_2 FILLER_2_1298 ();
 sg13g2_decap_8 FILLER_2_1304 ();
 sg13g2_fill_2 FILLER_2_1311 ();
 sg13g2_fill_1 FILLER_2_1313 ();
 sg13g2_decap_8 FILLER_2_1318 ();
 sg13g2_decap_8 FILLER_2_1325 ();
 sg13g2_decap_8 FILLER_2_1332 ();
 sg13g2_decap_8 FILLER_2_1339 ();
 sg13g2_decap_8 FILLER_2_1346 ();
 sg13g2_decap_8 FILLER_2_1353 ();
 sg13g2_decap_8 FILLER_2_1360 ();
 sg13g2_decap_8 FILLER_2_1367 ();
 sg13g2_decap_8 FILLER_2_1374 ();
 sg13g2_decap_8 FILLER_2_1381 ();
 sg13g2_decap_8 FILLER_2_1388 ();
 sg13g2_decap_8 FILLER_2_1395 ();
 sg13g2_decap_8 FILLER_2_1402 ();
 sg13g2_decap_8 FILLER_2_1409 ();
 sg13g2_decap_8 FILLER_2_1416 ();
 sg13g2_decap_8 FILLER_2_1423 ();
 sg13g2_decap_8 FILLER_2_1430 ();
 sg13g2_decap_8 FILLER_2_1437 ();
 sg13g2_decap_8 FILLER_2_1444 ();
 sg13g2_decap_8 FILLER_2_1451 ();
 sg13g2_decap_8 FILLER_2_1458 ();
 sg13g2_decap_8 FILLER_2_1465 ();
 sg13g2_decap_8 FILLER_2_1472 ();
 sg13g2_decap_8 FILLER_2_1479 ();
 sg13g2_decap_8 FILLER_2_1486 ();
 sg13g2_decap_8 FILLER_2_1493 ();
 sg13g2_decap_8 FILLER_2_1500 ();
 sg13g2_decap_8 FILLER_2_1507 ();
 sg13g2_decap_8 FILLER_2_1514 ();
 sg13g2_decap_8 FILLER_2_1521 ();
 sg13g2_decap_8 FILLER_2_1528 ();
 sg13g2_decap_8 FILLER_2_1535 ();
 sg13g2_decap_8 FILLER_2_1542 ();
 sg13g2_decap_8 FILLER_2_1549 ();
 sg13g2_decap_8 FILLER_2_1556 ();
 sg13g2_decap_8 FILLER_2_1563 ();
 sg13g2_decap_8 FILLER_2_1570 ();
 sg13g2_decap_8 FILLER_2_1577 ();
 sg13g2_decap_8 FILLER_2_1584 ();
 sg13g2_decap_8 FILLER_2_1591 ();
 sg13g2_decap_8 FILLER_2_1598 ();
 sg13g2_decap_8 FILLER_2_1605 ();
 sg13g2_decap_8 FILLER_2_1612 ();
 sg13g2_decap_8 FILLER_2_1619 ();
 sg13g2_decap_8 FILLER_2_1626 ();
 sg13g2_decap_8 FILLER_2_1633 ();
 sg13g2_decap_8 FILLER_2_1640 ();
 sg13g2_decap_8 FILLER_2_1647 ();
 sg13g2_decap_8 FILLER_2_1654 ();
 sg13g2_decap_8 FILLER_2_1661 ();
 sg13g2_decap_8 FILLER_2_1668 ();
 sg13g2_decap_8 FILLER_2_1675 ();
 sg13g2_decap_8 FILLER_2_1682 ();
 sg13g2_decap_8 FILLER_2_1689 ();
 sg13g2_decap_8 FILLER_2_1696 ();
 sg13g2_decap_8 FILLER_2_1703 ();
 sg13g2_decap_8 FILLER_2_1710 ();
 sg13g2_decap_8 FILLER_2_1717 ();
 sg13g2_decap_8 FILLER_2_1724 ();
 sg13g2_decap_8 FILLER_2_1731 ();
 sg13g2_decap_8 FILLER_2_1738 ();
 sg13g2_decap_8 FILLER_2_1745 ();
 sg13g2_decap_8 FILLER_2_1752 ();
 sg13g2_decap_8 FILLER_2_1759 ();
 sg13g2_decap_8 FILLER_2_1766 ();
 sg13g2_fill_1 FILLER_2_1773 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_4 FILLER_3_161 ();
 sg13g2_fill_1 FILLER_3_165 ();
 sg13g2_decap_4 FILLER_3_175 ();
 sg13g2_fill_1 FILLER_3_179 ();
 sg13g2_decap_4 FILLER_3_184 ();
 sg13g2_fill_1 FILLER_3_197 ();
 sg13g2_fill_1 FILLER_3_202 ();
 sg13g2_fill_2 FILLER_3_208 ();
 sg13g2_fill_2 FILLER_3_223 ();
 sg13g2_fill_1 FILLER_3_239 ();
 sg13g2_fill_1 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_fill_1 FILLER_3_299 ();
 sg13g2_fill_2 FILLER_3_308 ();
 sg13g2_fill_2 FILLER_3_317 ();
 sg13g2_fill_1 FILLER_3_319 ();
 sg13g2_decap_4 FILLER_3_328 ();
 sg13g2_fill_2 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_fill_1 FILLER_3_371 ();
 sg13g2_fill_1 FILLER_3_377 ();
 sg13g2_decap_4 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_404 ();
 sg13g2_decap_4 FILLER_3_411 ();
 sg13g2_fill_2 FILLER_3_415 ();
 sg13g2_decap_8 FILLER_3_422 ();
 sg13g2_decap_8 FILLER_3_429 ();
 sg13g2_fill_2 FILLER_3_436 ();
 sg13g2_fill_2 FILLER_3_450 ();
 sg13g2_fill_2 FILLER_3_466 ();
 sg13g2_fill_1 FILLER_3_477 ();
 sg13g2_fill_1 FILLER_3_483 ();
 sg13g2_fill_1 FILLER_3_493 ();
 sg13g2_fill_2 FILLER_3_499 ();
 sg13g2_decap_8 FILLER_3_510 ();
 sg13g2_decap_8 FILLER_3_517 ();
 sg13g2_decap_8 FILLER_3_524 ();
 sg13g2_decap_4 FILLER_3_531 ();
 sg13g2_fill_1 FILLER_3_535 ();
 sg13g2_decap_8 FILLER_3_545 ();
 sg13g2_fill_2 FILLER_3_557 ();
 sg13g2_fill_1 FILLER_3_580 ();
 sg13g2_fill_1 FILLER_3_594 ();
 sg13g2_decap_8 FILLER_3_624 ();
 sg13g2_fill_2 FILLER_3_631 ();
 sg13g2_fill_1 FILLER_3_633 ();
 sg13g2_fill_2 FILLER_3_639 ();
 sg13g2_fill_1 FILLER_3_641 ();
 sg13g2_fill_2 FILLER_3_646 ();
 sg13g2_fill_2 FILLER_3_690 ();
 sg13g2_fill_1 FILLER_3_692 ();
 sg13g2_fill_2 FILLER_3_698 ();
 sg13g2_decap_4 FILLER_3_705 ();
 sg13g2_decap_4 FILLER_3_716 ();
 sg13g2_fill_2 FILLER_3_729 ();
 sg13g2_decap_8 FILLER_3_739 ();
 sg13g2_decap_4 FILLER_3_746 ();
 sg13g2_decap_8 FILLER_3_759 ();
 sg13g2_decap_4 FILLER_3_766 ();
 sg13g2_decap_4 FILLER_3_790 ();
 sg13g2_fill_2 FILLER_3_794 ();
 sg13g2_fill_2 FILLER_3_806 ();
 sg13g2_fill_1 FILLER_3_808 ();
 sg13g2_fill_1 FILLER_3_814 ();
 sg13g2_fill_1 FILLER_3_846 ();
 sg13g2_fill_1 FILLER_3_855 ();
 sg13g2_fill_2 FILLER_3_869 ();
 sg13g2_decap_8 FILLER_3_876 ();
 sg13g2_decap_4 FILLER_3_883 ();
 sg13g2_fill_1 FILLER_3_887 ();
 sg13g2_decap_8 FILLER_3_896 ();
 sg13g2_fill_1 FILLER_3_912 ();
 sg13g2_fill_2 FILLER_3_918 ();
 sg13g2_fill_2 FILLER_3_925 ();
 sg13g2_decap_4 FILLER_3_932 ();
 sg13g2_fill_1 FILLER_3_940 ();
 sg13g2_fill_1 FILLER_3_947 ();
 sg13g2_fill_2 FILLER_3_952 ();
 sg13g2_fill_1 FILLER_3_954 ();
 sg13g2_fill_1 FILLER_3_967 ();
 sg13g2_decap_8 FILLER_3_973 ();
 sg13g2_fill_2 FILLER_3_980 ();
 sg13g2_fill_1 FILLER_3_982 ();
 sg13g2_decap_8 FILLER_3_988 ();
 sg13g2_fill_2 FILLER_3_995 ();
 sg13g2_fill_1 FILLER_3_997 ();
 sg13g2_fill_1 FILLER_3_1006 ();
 sg13g2_decap_8 FILLER_3_1041 ();
 sg13g2_fill_2 FILLER_3_1048 ();
 sg13g2_fill_1 FILLER_3_1050 ();
 sg13g2_decap_8 FILLER_3_1070 ();
 sg13g2_decap_4 FILLER_3_1077 ();
 sg13g2_fill_2 FILLER_3_1081 ();
 sg13g2_fill_1 FILLER_3_1097 ();
 sg13g2_decap_8 FILLER_3_1129 ();
 sg13g2_fill_1 FILLER_3_1136 ();
 sg13g2_fill_2 FILLER_3_1142 ();
 sg13g2_fill_1 FILLER_3_1150 ();
 sg13g2_decap_8 FILLER_3_1163 ();
 sg13g2_decap_8 FILLER_3_1170 ();
 sg13g2_fill_2 FILLER_3_1177 ();
 sg13g2_fill_2 FILLER_3_1198 ();
 sg13g2_fill_1 FILLER_3_1205 ();
 sg13g2_fill_2 FILLER_3_1221 ();
 sg13g2_decap_4 FILLER_3_1228 ();
 sg13g2_fill_1 FILLER_3_1252 ();
 sg13g2_decap_8 FILLER_3_1274 ();
 sg13g2_decap_8 FILLER_3_1281 ();
 sg13g2_fill_2 FILLER_3_1288 ();
 sg13g2_decap_8 FILLER_3_1298 ();
 sg13g2_decap_8 FILLER_3_1305 ();
 sg13g2_fill_2 FILLER_3_1312 ();
 sg13g2_decap_8 FILLER_3_1323 ();
 sg13g2_decap_4 FILLER_3_1330 ();
 sg13g2_decap_8 FILLER_3_1338 ();
 sg13g2_fill_1 FILLER_3_1345 ();
 sg13g2_fill_1 FILLER_3_1355 ();
 sg13g2_decap_8 FILLER_3_1360 ();
 sg13g2_decap_8 FILLER_3_1367 ();
 sg13g2_decap_8 FILLER_3_1374 ();
 sg13g2_decap_8 FILLER_3_1381 ();
 sg13g2_decap_8 FILLER_3_1388 ();
 sg13g2_decap_8 FILLER_3_1395 ();
 sg13g2_decap_8 FILLER_3_1402 ();
 sg13g2_decap_8 FILLER_3_1409 ();
 sg13g2_decap_8 FILLER_3_1416 ();
 sg13g2_decap_8 FILLER_3_1423 ();
 sg13g2_decap_8 FILLER_3_1430 ();
 sg13g2_decap_8 FILLER_3_1437 ();
 sg13g2_decap_8 FILLER_3_1444 ();
 sg13g2_decap_8 FILLER_3_1451 ();
 sg13g2_decap_8 FILLER_3_1458 ();
 sg13g2_decap_8 FILLER_3_1465 ();
 sg13g2_decap_8 FILLER_3_1472 ();
 sg13g2_decap_8 FILLER_3_1479 ();
 sg13g2_decap_8 FILLER_3_1486 ();
 sg13g2_decap_8 FILLER_3_1493 ();
 sg13g2_decap_8 FILLER_3_1500 ();
 sg13g2_decap_8 FILLER_3_1507 ();
 sg13g2_decap_8 FILLER_3_1514 ();
 sg13g2_decap_8 FILLER_3_1521 ();
 sg13g2_decap_8 FILLER_3_1528 ();
 sg13g2_decap_8 FILLER_3_1535 ();
 sg13g2_decap_8 FILLER_3_1542 ();
 sg13g2_decap_8 FILLER_3_1549 ();
 sg13g2_decap_8 FILLER_3_1556 ();
 sg13g2_decap_8 FILLER_3_1563 ();
 sg13g2_decap_8 FILLER_3_1570 ();
 sg13g2_decap_8 FILLER_3_1577 ();
 sg13g2_decap_8 FILLER_3_1584 ();
 sg13g2_decap_8 FILLER_3_1591 ();
 sg13g2_decap_8 FILLER_3_1598 ();
 sg13g2_decap_8 FILLER_3_1605 ();
 sg13g2_decap_8 FILLER_3_1612 ();
 sg13g2_decap_8 FILLER_3_1619 ();
 sg13g2_decap_8 FILLER_3_1626 ();
 sg13g2_decap_8 FILLER_3_1633 ();
 sg13g2_decap_8 FILLER_3_1640 ();
 sg13g2_decap_8 FILLER_3_1647 ();
 sg13g2_decap_8 FILLER_3_1654 ();
 sg13g2_decap_8 FILLER_3_1661 ();
 sg13g2_decap_8 FILLER_3_1668 ();
 sg13g2_decap_8 FILLER_3_1675 ();
 sg13g2_decap_8 FILLER_3_1682 ();
 sg13g2_decap_8 FILLER_3_1689 ();
 sg13g2_decap_8 FILLER_3_1696 ();
 sg13g2_decap_8 FILLER_3_1703 ();
 sg13g2_decap_8 FILLER_3_1710 ();
 sg13g2_decap_8 FILLER_3_1717 ();
 sg13g2_decap_8 FILLER_3_1724 ();
 sg13g2_decap_8 FILLER_3_1731 ();
 sg13g2_decap_8 FILLER_3_1738 ();
 sg13g2_decap_8 FILLER_3_1745 ();
 sg13g2_decap_8 FILLER_3_1752 ();
 sg13g2_decap_8 FILLER_3_1759 ();
 sg13g2_decap_8 FILLER_3_1766 ();
 sg13g2_fill_1 FILLER_3_1773 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_fill_1 FILLER_4_173 ();
 sg13g2_decap_4 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_202 ();
 sg13g2_fill_2 FILLER_4_227 ();
 sg13g2_decap_4 FILLER_4_244 ();
 sg13g2_fill_1 FILLER_4_252 ();
 sg13g2_fill_1 FILLER_4_269 ();
 sg13g2_fill_1 FILLER_4_274 ();
 sg13g2_fill_1 FILLER_4_301 ();
 sg13g2_fill_1 FILLER_4_306 ();
 sg13g2_fill_2 FILLER_4_312 ();
 sg13g2_fill_1 FILLER_4_314 ();
 sg13g2_decap_4 FILLER_4_324 ();
 sg13g2_fill_2 FILLER_4_328 ();
 sg13g2_decap_4 FILLER_4_343 ();
 sg13g2_fill_1 FILLER_4_355 ();
 sg13g2_decap_4 FILLER_4_366 ();
 sg13g2_fill_2 FILLER_4_390 ();
 sg13g2_fill_1 FILLER_4_392 ();
 sg13g2_fill_2 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_422 ();
 sg13g2_fill_2 FILLER_4_435 ();
 sg13g2_fill_1 FILLER_4_441 ();
 sg13g2_fill_1 FILLER_4_452 ();
 sg13g2_decap_8 FILLER_4_471 ();
 sg13g2_fill_1 FILLER_4_487 ();
 sg13g2_fill_2 FILLER_4_503 ();
 sg13g2_fill_2 FILLER_4_514 ();
 sg13g2_decap_8 FILLER_4_521 ();
 sg13g2_decap_8 FILLER_4_528 ();
 sg13g2_decap_8 FILLER_4_535 ();
 sg13g2_decap_8 FILLER_4_542 ();
 sg13g2_decap_8 FILLER_4_549 ();
 sg13g2_fill_2 FILLER_4_556 ();
 sg13g2_fill_1 FILLER_4_558 ();
 sg13g2_decap_8 FILLER_4_564 ();
 sg13g2_fill_2 FILLER_4_571 ();
 sg13g2_fill_1 FILLER_4_595 ();
 sg13g2_fill_1 FILLER_4_599 ();
 sg13g2_fill_2 FILLER_4_605 ();
 sg13g2_fill_2 FILLER_4_611 ();
 sg13g2_fill_1 FILLER_4_613 ();
 sg13g2_fill_2 FILLER_4_619 ();
 sg13g2_fill_2 FILLER_4_626 ();
 sg13g2_fill_1 FILLER_4_628 ();
 sg13g2_decap_8 FILLER_4_634 ();
 sg13g2_fill_1 FILLER_4_641 ();
 sg13g2_fill_1 FILLER_4_647 ();
 sg13g2_fill_1 FILLER_4_656 ();
 sg13g2_fill_2 FILLER_4_669 ();
 sg13g2_fill_2 FILLER_4_686 ();
 sg13g2_fill_1 FILLER_4_688 ();
 sg13g2_fill_1 FILLER_4_694 ();
 sg13g2_fill_2 FILLER_4_700 ();
 sg13g2_fill_1 FILLER_4_706 ();
 sg13g2_fill_2 FILLER_4_715 ();
 sg13g2_fill_2 FILLER_4_722 ();
 sg13g2_fill_2 FILLER_4_729 ();
 sg13g2_decap_8 FILLER_4_736 ();
 sg13g2_fill_1 FILLER_4_743 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_4 FILLER_4_756 ();
 sg13g2_fill_2 FILLER_4_760 ();
 sg13g2_fill_1 FILLER_4_771 ();
 sg13g2_fill_2 FILLER_4_803 ();
 sg13g2_fill_2 FILLER_4_836 ();
 sg13g2_fill_1 FILLER_4_838 ();
 sg13g2_fill_2 FILLER_4_852 ();
 sg13g2_decap_8 FILLER_4_859 ();
 sg13g2_decap_8 FILLER_4_866 ();
 sg13g2_fill_1 FILLER_4_873 ();
 sg13g2_decap_4 FILLER_4_878 ();
 sg13g2_fill_1 FILLER_4_882 ();
 sg13g2_decap_8 FILLER_4_888 ();
 sg13g2_decap_4 FILLER_4_899 ();
 sg13g2_fill_1 FILLER_4_903 ();
 sg13g2_decap_4 FILLER_4_942 ();
 sg13g2_fill_2 FILLER_4_946 ();
 sg13g2_fill_2 FILLER_4_957 ();
 sg13g2_fill_1 FILLER_4_959 ();
 sg13g2_fill_1 FILLER_4_964 ();
 sg13g2_decap_4 FILLER_4_984 ();
 sg13g2_fill_1 FILLER_4_992 ();
 sg13g2_fill_2 FILLER_4_1041 ();
 sg13g2_fill_2 FILLER_4_1048 ();
 sg13g2_fill_2 FILLER_4_1055 ();
 sg13g2_fill_1 FILLER_4_1057 ();
 sg13g2_decap_4 FILLER_4_1062 ();
 sg13g2_fill_1 FILLER_4_1066 ();
 sg13g2_decap_4 FILLER_4_1071 ();
 sg13g2_fill_1 FILLER_4_1083 ();
 sg13g2_fill_1 FILLER_4_1098 ();
 sg13g2_fill_2 FILLER_4_1108 ();
 sg13g2_fill_1 FILLER_4_1119 ();
 sg13g2_fill_2 FILLER_4_1139 ();
 sg13g2_fill_2 FILLER_4_1155 ();
 sg13g2_fill_1 FILLER_4_1157 ();
 sg13g2_fill_1 FILLER_4_1168 ();
 sg13g2_decap_4 FILLER_4_1174 ();
 sg13g2_fill_1 FILLER_4_1178 ();
 sg13g2_decap_4 FILLER_4_1184 ();
 sg13g2_fill_2 FILLER_4_1197 ();
 sg13g2_fill_1 FILLER_4_1199 ();
 sg13g2_fill_1 FILLER_4_1213 ();
 sg13g2_fill_2 FILLER_4_1224 ();
 sg13g2_fill_1 FILLER_4_1226 ();
 sg13g2_fill_1 FILLER_4_1235 ();
 sg13g2_fill_2 FILLER_4_1241 ();
 sg13g2_fill_1 FILLER_4_1248 ();
 sg13g2_fill_1 FILLER_4_1254 ();
 sg13g2_fill_2 FILLER_4_1260 ();
 sg13g2_fill_1 FILLER_4_1262 ();
 sg13g2_fill_1 FILLER_4_1278 ();
 sg13g2_fill_2 FILLER_4_1287 ();
 sg13g2_decap_4 FILLER_4_1298 ();
 sg13g2_fill_2 FILLER_4_1302 ();
 sg13g2_decap_4 FILLER_4_1309 ();
 sg13g2_fill_2 FILLER_4_1313 ();
 sg13g2_fill_2 FILLER_4_1323 ();
 sg13g2_fill_1 FILLER_4_1325 ();
 sg13g2_fill_1 FILLER_4_1340 ();
 sg13g2_fill_2 FILLER_4_1365 ();
 sg13g2_fill_2 FILLER_4_1372 ();
 sg13g2_fill_1 FILLER_4_1374 ();
 sg13g2_fill_1 FILLER_4_1380 ();
 sg13g2_decap_8 FILLER_4_1385 ();
 sg13g2_decap_8 FILLER_4_1392 ();
 sg13g2_decap_8 FILLER_4_1399 ();
 sg13g2_decap_8 FILLER_4_1406 ();
 sg13g2_decap_8 FILLER_4_1413 ();
 sg13g2_decap_8 FILLER_4_1420 ();
 sg13g2_decap_8 FILLER_4_1427 ();
 sg13g2_decap_8 FILLER_4_1434 ();
 sg13g2_decap_8 FILLER_4_1441 ();
 sg13g2_decap_8 FILLER_4_1448 ();
 sg13g2_decap_8 FILLER_4_1455 ();
 sg13g2_decap_8 FILLER_4_1462 ();
 sg13g2_decap_8 FILLER_4_1469 ();
 sg13g2_decap_8 FILLER_4_1476 ();
 sg13g2_decap_8 FILLER_4_1483 ();
 sg13g2_decap_8 FILLER_4_1490 ();
 sg13g2_decap_8 FILLER_4_1497 ();
 sg13g2_decap_8 FILLER_4_1504 ();
 sg13g2_decap_8 FILLER_4_1511 ();
 sg13g2_decap_8 FILLER_4_1518 ();
 sg13g2_decap_8 FILLER_4_1525 ();
 sg13g2_decap_8 FILLER_4_1532 ();
 sg13g2_decap_8 FILLER_4_1539 ();
 sg13g2_decap_8 FILLER_4_1546 ();
 sg13g2_decap_8 FILLER_4_1553 ();
 sg13g2_decap_8 FILLER_4_1560 ();
 sg13g2_decap_8 FILLER_4_1567 ();
 sg13g2_decap_8 FILLER_4_1574 ();
 sg13g2_decap_8 FILLER_4_1581 ();
 sg13g2_decap_8 FILLER_4_1588 ();
 sg13g2_decap_8 FILLER_4_1595 ();
 sg13g2_decap_8 FILLER_4_1602 ();
 sg13g2_decap_8 FILLER_4_1609 ();
 sg13g2_decap_8 FILLER_4_1616 ();
 sg13g2_decap_8 FILLER_4_1623 ();
 sg13g2_decap_8 FILLER_4_1630 ();
 sg13g2_decap_8 FILLER_4_1637 ();
 sg13g2_decap_8 FILLER_4_1644 ();
 sg13g2_decap_8 FILLER_4_1651 ();
 sg13g2_decap_8 FILLER_4_1658 ();
 sg13g2_decap_8 FILLER_4_1665 ();
 sg13g2_decap_8 FILLER_4_1672 ();
 sg13g2_decap_8 FILLER_4_1679 ();
 sg13g2_decap_8 FILLER_4_1686 ();
 sg13g2_decap_8 FILLER_4_1693 ();
 sg13g2_decap_8 FILLER_4_1700 ();
 sg13g2_decap_8 FILLER_4_1707 ();
 sg13g2_decap_8 FILLER_4_1714 ();
 sg13g2_decap_8 FILLER_4_1721 ();
 sg13g2_decap_8 FILLER_4_1728 ();
 sg13g2_decap_8 FILLER_4_1735 ();
 sg13g2_decap_8 FILLER_4_1742 ();
 sg13g2_decap_8 FILLER_4_1749 ();
 sg13g2_decap_8 FILLER_4_1756 ();
 sg13g2_decap_8 FILLER_4_1763 ();
 sg13g2_decap_4 FILLER_4_1770 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_fill_2 FILLER_5_108 ();
 sg13g2_fill_2 FILLER_5_113 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_decap_4 FILLER_5_124 ();
 sg13g2_fill_1 FILLER_5_128 ();
 sg13g2_decap_4 FILLER_5_134 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_fill_1 FILLER_5_150 ();
 sg13g2_decap_4 FILLER_5_167 ();
 sg13g2_fill_2 FILLER_5_171 ();
 sg13g2_fill_2 FILLER_5_178 ();
 sg13g2_fill_1 FILLER_5_180 ();
 sg13g2_fill_2 FILLER_5_189 ();
 sg13g2_fill_1 FILLER_5_204 ();
 sg13g2_decap_8 FILLER_5_213 ();
 sg13g2_fill_2 FILLER_5_220 ();
 sg13g2_decap_4 FILLER_5_232 ();
 sg13g2_fill_2 FILLER_5_241 ();
 sg13g2_fill_2 FILLER_5_248 ();
 sg13g2_decap_4 FILLER_5_269 ();
 sg13g2_fill_2 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_fill_2 FILLER_5_341 ();
 sg13g2_fill_1 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_fill_2 FILLER_5_363 ();
 sg13g2_fill_1 FILLER_5_365 ();
 sg13g2_fill_1 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_decap_8 FILLER_5_407 ();
 sg13g2_fill_2 FILLER_5_414 ();
 sg13g2_fill_1 FILLER_5_416 ();
 sg13g2_fill_2 FILLER_5_436 ();
 sg13g2_fill_1 FILLER_5_438 ();
 sg13g2_fill_1 FILLER_5_444 ();
 sg13g2_fill_1 FILLER_5_450 ();
 sg13g2_fill_1 FILLER_5_460 ();
 sg13g2_fill_1 FILLER_5_470 ();
 sg13g2_fill_2 FILLER_5_474 ();
 sg13g2_decap_8 FILLER_5_485 ();
 sg13g2_decap_8 FILLER_5_492 ();
 sg13g2_fill_2 FILLER_5_499 ();
 sg13g2_fill_2 FILLER_5_521 ();
 sg13g2_fill_1 FILLER_5_590 ();
 sg13g2_fill_2 FILLER_5_621 ();
 sg13g2_fill_1 FILLER_5_623 ();
 sg13g2_decap_4 FILLER_5_641 ();
 sg13g2_fill_1 FILLER_5_645 ();
 sg13g2_decap_4 FILLER_5_651 ();
 sg13g2_fill_2 FILLER_5_674 ();
 sg13g2_fill_1 FILLER_5_676 ();
 sg13g2_fill_2 FILLER_5_689 ();
 sg13g2_fill_2 FILLER_5_696 ();
 sg13g2_fill_2 FILLER_5_703 ();
 sg13g2_fill_2 FILLER_5_710 ();
 sg13g2_fill_1 FILLER_5_712 ();
 sg13g2_fill_2 FILLER_5_718 ();
 sg13g2_fill_1 FILLER_5_720 ();
 sg13g2_fill_2 FILLER_5_726 ();
 sg13g2_decap_8 FILLER_5_733 ();
 sg13g2_fill_2 FILLER_5_740 ();
 sg13g2_fill_1 FILLER_5_751 ();
 sg13g2_decap_4 FILLER_5_778 ();
 sg13g2_fill_1 FILLER_5_782 ();
 sg13g2_decap_4 FILLER_5_788 ();
 sg13g2_fill_2 FILLER_5_792 ();
 sg13g2_fill_2 FILLER_5_803 ();
 sg13g2_fill_2 FILLER_5_814 ();
 sg13g2_fill_1 FILLER_5_816 ();
 sg13g2_fill_2 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_843 ();
 sg13g2_decap_8 FILLER_5_850 ();
 sg13g2_decap_8 FILLER_5_857 ();
 sg13g2_decap_4 FILLER_5_864 ();
 sg13g2_fill_1 FILLER_5_868 ();
 sg13g2_decap_4 FILLER_5_877 ();
 sg13g2_fill_2 FILLER_5_881 ();
 sg13g2_fill_1 FILLER_5_901 ();
 sg13g2_decap_8 FILLER_5_928 ();
 sg13g2_fill_1 FILLER_5_939 ();
 sg13g2_fill_2 FILLER_5_943 ();
 sg13g2_fill_1 FILLER_5_949 ();
 sg13g2_decap_8 FILLER_5_958 ();
 sg13g2_fill_2 FILLER_5_965 ();
 sg13g2_fill_1 FILLER_5_967 ();
 sg13g2_decap_4 FILLER_5_977 ();
 sg13g2_fill_2 FILLER_5_981 ();
 sg13g2_fill_1 FILLER_5_993 ();
 sg13g2_fill_2 FILLER_5_1000 ();
 sg13g2_fill_1 FILLER_5_1002 ();
 sg13g2_fill_2 FILLER_5_1011 ();
 sg13g2_fill_1 FILLER_5_1013 ();
 sg13g2_fill_2 FILLER_5_1022 ();
 sg13g2_fill_2 FILLER_5_1029 ();
 sg13g2_decap_8 FILLER_5_1044 ();
 sg13g2_decap_8 FILLER_5_1051 ();
 sg13g2_decap_8 FILLER_5_1058 ();
 sg13g2_decap_8 FILLER_5_1065 ();
 sg13g2_fill_2 FILLER_5_1072 ();
 sg13g2_fill_2 FILLER_5_1081 ();
 sg13g2_fill_1 FILLER_5_1083 ();
 sg13g2_decap_4 FILLER_5_1089 ();
 sg13g2_fill_1 FILLER_5_1093 ();
 sg13g2_fill_1 FILLER_5_1106 ();
 sg13g2_fill_2 FILLER_5_1122 ();
 sg13g2_decap_4 FILLER_5_1132 ();
 sg13g2_fill_1 FILLER_5_1136 ();
 sg13g2_fill_1 FILLER_5_1142 ();
 sg13g2_fill_1 FILLER_5_1150 ();
 sg13g2_fill_2 FILLER_5_1165 ();
 sg13g2_decap_8 FILLER_5_1172 ();
 sg13g2_decap_8 FILLER_5_1179 ();
 sg13g2_decap_8 FILLER_5_1186 ();
 sg13g2_decap_4 FILLER_5_1193 ();
 sg13g2_fill_1 FILLER_5_1202 ();
 sg13g2_decap_8 FILLER_5_1226 ();
 sg13g2_fill_2 FILLER_5_1233 ();
 sg13g2_fill_2 FILLER_5_1247 ();
 sg13g2_fill_1 FILLER_5_1249 ();
 sg13g2_fill_1 FILLER_5_1259 ();
 sg13g2_decap_8 FILLER_5_1265 ();
 sg13g2_decap_8 FILLER_5_1272 ();
 sg13g2_decap_4 FILLER_5_1279 ();
 sg13g2_fill_1 FILLER_5_1283 ();
 sg13g2_fill_1 FILLER_5_1308 ();
 sg13g2_fill_1 FILLER_5_1313 ();
 sg13g2_fill_1 FILLER_5_1318 ();
 sg13g2_fill_2 FILLER_5_1324 ();
 sg13g2_fill_1 FILLER_5_1339 ();
 sg13g2_fill_1 FILLER_5_1344 ();
 sg13g2_fill_1 FILLER_5_1350 ();
 sg13g2_fill_2 FILLER_5_1356 ();
 sg13g2_fill_2 FILLER_5_1397 ();
 sg13g2_fill_2 FILLER_5_1404 ();
 sg13g2_fill_1 FILLER_5_1406 ();
 sg13g2_fill_2 FILLER_5_1420 ();
 sg13g2_decap_8 FILLER_5_1426 ();
 sg13g2_decap_8 FILLER_5_1433 ();
 sg13g2_decap_8 FILLER_5_1440 ();
 sg13g2_decap_8 FILLER_5_1447 ();
 sg13g2_decap_8 FILLER_5_1454 ();
 sg13g2_decap_8 FILLER_5_1461 ();
 sg13g2_decap_8 FILLER_5_1468 ();
 sg13g2_decap_8 FILLER_5_1475 ();
 sg13g2_decap_8 FILLER_5_1482 ();
 sg13g2_fill_2 FILLER_5_1489 ();
 sg13g2_fill_1 FILLER_5_1491 ();
 sg13g2_decap_8 FILLER_5_1496 ();
 sg13g2_decap_8 FILLER_5_1503 ();
 sg13g2_decap_8 FILLER_5_1510 ();
 sg13g2_decap_8 FILLER_5_1517 ();
 sg13g2_decap_8 FILLER_5_1524 ();
 sg13g2_decap_8 FILLER_5_1531 ();
 sg13g2_decap_8 FILLER_5_1538 ();
 sg13g2_decap_8 FILLER_5_1545 ();
 sg13g2_decap_8 FILLER_5_1552 ();
 sg13g2_decap_8 FILLER_5_1559 ();
 sg13g2_decap_8 FILLER_5_1566 ();
 sg13g2_decap_8 FILLER_5_1573 ();
 sg13g2_decap_8 FILLER_5_1580 ();
 sg13g2_decap_8 FILLER_5_1587 ();
 sg13g2_decap_8 FILLER_5_1594 ();
 sg13g2_decap_8 FILLER_5_1601 ();
 sg13g2_decap_8 FILLER_5_1608 ();
 sg13g2_decap_8 FILLER_5_1615 ();
 sg13g2_decap_8 FILLER_5_1622 ();
 sg13g2_decap_8 FILLER_5_1629 ();
 sg13g2_decap_8 FILLER_5_1636 ();
 sg13g2_decap_8 FILLER_5_1643 ();
 sg13g2_decap_8 FILLER_5_1650 ();
 sg13g2_decap_8 FILLER_5_1657 ();
 sg13g2_decap_8 FILLER_5_1664 ();
 sg13g2_decap_8 FILLER_5_1671 ();
 sg13g2_decap_8 FILLER_5_1678 ();
 sg13g2_decap_8 FILLER_5_1685 ();
 sg13g2_decap_8 FILLER_5_1692 ();
 sg13g2_decap_8 FILLER_5_1699 ();
 sg13g2_decap_8 FILLER_5_1706 ();
 sg13g2_decap_8 FILLER_5_1713 ();
 sg13g2_decap_8 FILLER_5_1720 ();
 sg13g2_decap_8 FILLER_5_1727 ();
 sg13g2_decap_8 FILLER_5_1734 ();
 sg13g2_decap_8 FILLER_5_1741 ();
 sg13g2_decap_8 FILLER_5_1748 ();
 sg13g2_decap_8 FILLER_5_1755 ();
 sg13g2_decap_8 FILLER_5_1762 ();
 sg13g2_decap_4 FILLER_5_1769 ();
 sg13g2_fill_1 FILLER_5_1773 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_91 ();
 sg13g2_fill_1 FILLER_6_109 ();
 sg13g2_fill_1 FILLER_6_139 ();
 sg13g2_fill_1 FILLER_6_154 ();
 sg13g2_fill_1 FILLER_6_164 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_4 FILLER_6_186 ();
 sg13g2_fill_2 FILLER_6_190 ();
 sg13g2_decap_4 FILLER_6_196 ();
 sg13g2_fill_1 FILLER_6_200 ();
 sg13g2_decap_4 FILLER_6_210 ();
 sg13g2_fill_2 FILLER_6_219 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_fill_2 FILLER_6_264 ();
 sg13g2_decap_8 FILLER_6_274 ();
 sg13g2_decap_4 FILLER_6_281 ();
 sg13g2_fill_2 FILLER_6_311 ();
 sg13g2_fill_1 FILLER_6_313 ();
 sg13g2_fill_2 FILLER_6_328 ();
 sg13g2_fill_1 FILLER_6_330 ();
 sg13g2_fill_1 FILLER_6_349 ();
 sg13g2_decap_4 FILLER_6_362 ();
 sg13g2_fill_1 FILLER_6_366 ();
 sg13g2_fill_2 FILLER_6_372 ();
 sg13g2_fill_2 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_6_408 ();
 sg13g2_fill_1 FILLER_6_415 ();
 sg13g2_decap_4 FILLER_6_420 ();
 sg13g2_fill_1 FILLER_6_424 ();
 sg13g2_fill_1 FILLER_6_433 ();
 sg13g2_fill_2 FILLER_6_463 ();
 sg13g2_decap_4 FILLER_6_473 ();
 sg13g2_fill_2 FILLER_6_482 ();
 sg13g2_decap_8 FILLER_6_492 ();
 sg13g2_decap_8 FILLER_6_499 ();
 sg13g2_decap_8 FILLER_6_506 ();
 sg13g2_decap_4 FILLER_6_518 ();
 sg13g2_fill_1 FILLER_6_548 ();
 sg13g2_fill_1 FILLER_6_564 ();
 sg13g2_fill_2 FILLER_6_577 ();
 sg13g2_fill_2 FILLER_6_604 ();
 sg13g2_fill_1 FILLER_6_629 ();
 sg13g2_decap_8 FILLER_6_635 ();
 sg13g2_fill_2 FILLER_6_642 ();
 sg13g2_fill_1 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_649 ();
 sg13g2_decap_8 FILLER_6_660 ();
 sg13g2_fill_1 FILLER_6_667 ();
 sg13g2_fill_1 FILLER_6_673 ();
 sg13g2_fill_2 FILLER_6_679 ();
 sg13g2_fill_1 FILLER_6_681 ();
 sg13g2_fill_1 FILLER_6_708 ();
 sg13g2_fill_1 FILLER_6_713 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_fill_2 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_fill_1 FILLER_6_767 ();
 sg13g2_decap_4 FILLER_6_780 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_fill_1 FILLER_6_795 ();
 sg13g2_fill_1 FILLER_6_807 ();
 sg13g2_fill_2 FILLER_6_812 ();
 sg13g2_fill_2 FILLER_6_819 ();
 sg13g2_fill_1 FILLER_6_834 ();
 sg13g2_fill_1 FILLER_6_839 ();
 sg13g2_decap_8 FILLER_6_845 ();
 sg13g2_decap_4 FILLER_6_852 ();
 sg13g2_fill_1 FILLER_6_856 ();
 sg13g2_decap_8 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_869 ();
 sg13g2_decap_8 FILLER_6_876 ();
 sg13g2_fill_2 FILLER_6_883 ();
 sg13g2_fill_1 FILLER_6_890 ();
 sg13g2_decap_4 FILLER_6_899 ();
 sg13g2_decap_4 FILLER_6_908 ();
 sg13g2_fill_2 FILLER_6_916 ();
 sg13g2_fill_1 FILLER_6_918 ();
 sg13g2_fill_2 FILLER_6_937 ();
 sg13g2_decap_8 FILLER_6_951 ();
 sg13g2_decap_8 FILLER_6_958 ();
 sg13g2_decap_8 FILLER_6_965 ();
 sg13g2_decap_8 FILLER_6_972 ();
 sg13g2_fill_2 FILLER_6_1000 ();
 sg13g2_fill_1 FILLER_6_1002 ();
 sg13g2_fill_2 FILLER_6_1008 ();
 sg13g2_fill_1 FILLER_6_1015 ();
 sg13g2_fill_2 FILLER_6_1020 ();
 sg13g2_fill_1 FILLER_6_1030 ();
 sg13g2_fill_2 FILLER_6_1036 ();
 sg13g2_fill_2 FILLER_6_1043 ();
 sg13g2_decap_8 FILLER_6_1050 ();
 sg13g2_decap_4 FILLER_6_1057 ();
 sg13g2_decap_8 FILLER_6_1068 ();
 sg13g2_fill_1 FILLER_6_1075 ();
 sg13g2_fill_1 FILLER_6_1086 ();
 sg13g2_fill_2 FILLER_6_1116 ();
 sg13g2_fill_1 FILLER_6_1118 ();
 sg13g2_decap_8 FILLER_6_1122 ();
 sg13g2_decap_4 FILLER_6_1173 ();
 sg13g2_fill_1 FILLER_6_1191 ();
 sg13g2_fill_2 FILLER_6_1201 ();
 sg13g2_decap_4 FILLER_6_1216 ();
 sg13g2_fill_1 FILLER_6_1268 ();
 sg13g2_fill_1 FILLER_6_1274 ();
 sg13g2_fill_1 FILLER_6_1284 ();
 sg13g2_fill_2 FILLER_6_1290 ();
 sg13g2_fill_1 FILLER_6_1292 ();
 sg13g2_decap_8 FILLER_6_1298 ();
 sg13g2_decap_4 FILLER_6_1305 ();
 sg13g2_fill_1 FILLER_6_1309 ();
 sg13g2_fill_2 FILLER_6_1315 ();
 sg13g2_fill_1 FILLER_6_1317 ();
 sg13g2_fill_1 FILLER_6_1326 ();
 sg13g2_fill_1 FILLER_6_1340 ();
 sg13g2_fill_1 FILLER_6_1345 ();
 sg13g2_decap_4 FILLER_6_1356 ();
 sg13g2_decap_8 FILLER_6_1369 ();
 sg13g2_fill_2 FILLER_6_1376 ();
 sg13g2_fill_2 FILLER_6_1396 ();
 sg13g2_decap_4 FILLER_6_1403 ();
 sg13g2_fill_2 FILLER_6_1407 ();
 sg13g2_decap_4 FILLER_6_1414 ();
 sg13g2_fill_2 FILLER_6_1418 ();
 sg13g2_fill_1 FILLER_6_1428 ();
 sg13g2_decap_8 FILLER_6_1434 ();
 sg13g2_fill_1 FILLER_6_1441 ();
 sg13g2_fill_1 FILLER_6_1452 ();
 sg13g2_decap_8 FILLER_6_1460 ();
 sg13g2_decap_8 FILLER_6_1467 ();
 sg13g2_fill_2 FILLER_6_1474 ();
 sg13g2_fill_1 FILLER_6_1476 ();
 sg13g2_fill_2 FILLER_6_1482 ();
 sg13g2_decap_8 FILLER_6_1510 ();
 sg13g2_decap_8 FILLER_6_1517 ();
 sg13g2_decap_8 FILLER_6_1524 ();
 sg13g2_decap_8 FILLER_6_1531 ();
 sg13g2_decap_8 FILLER_6_1538 ();
 sg13g2_decap_8 FILLER_6_1545 ();
 sg13g2_decap_8 FILLER_6_1552 ();
 sg13g2_decap_8 FILLER_6_1559 ();
 sg13g2_decap_8 FILLER_6_1566 ();
 sg13g2_decap_8 FILLER_6_1573 ();
 sg13g2_decap_8 FILLER_6_1580 ();
 sg13g2_decap_8 FILLER_6_1587 ();
 sg13g2_decap_8 FILLER_6_1594 ();
 sg13g2_decap_8 FILLER_6_1601 ();
 sg13g2_decap_8 FILLER_6_1608 ();
 sg13g2_decap_8 FILLER_6_1615 ();
 sg13g2_decap_8 FILLER_6_1622 ();
 sg13g2_decap_8 FILLER_6_1629 ();
 sg13g2_decap_8 FILLER_6_1636 ();
 sg13g2_decap_8 FILLER_6_1643 ();
 sg13g2_decap_8 FILLER_6_1650 ();
 sg13g2_decap_8 FILLER_6_1657 ();
 sg13g2_decap_8 FILLER_6_1664 ();
 sg13g2_decap_8 FILLER_6_1671 ();
 sg13g2_decap_8 FILLER_6_1678 ();
 sg13g2_decap_8 FILLER_6_1685 ();
 sg13g2_decap_8 FILLER_6_1692 ();
 sg13g2_decap_8 FILLER_6_1699 ();
 sg13g2_decap_8 FILLER_6_1706 ();
 sg13g2_decap_8 FILLER_6_1713 ();
 sg13g2_decap_8 FILLER_6_1720 ();
 sg13g2_decap_8 FILLER_6_1727 ();
 sg13g2_decap_8 FILLER_6_1734 ();
 sg13g2_decap_8 FILLER_6_1741 ();
 sg13g2_decap_8 FILLER_6_1748 ();
 sg13g2_decap_8 FILLER_6_1755 ();
 sg13g2_decap_8 FILLER_6_1762 ();
 sg13g2_decap_4 FILLER_6_1769 ();
 sg13g2_fill_1 FILLER_6_1773 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_fill_1 FILLER_7_74 ();
 sg13g2_fill_2 FILLER_7_79 ();
 sg13g2_fill_1 FILLER_7_89 ();
 sg13g2_fill_2 FILLER_7_94 ();
 sg13g2_fill_1 FILLER_7_122 ();
 sg13g2_fill_1 FILLER_7_147 ();
 sg13g2_fill_2 FILLER_7_156 ();
 sg13g2_fill_2 FILLER_7_163 ();
 sg13g2_fill_1 FILLER_7_170 ();
 sg13g2_decap_8 FILLER_7_179 ();
 sg13g2_fill_2 FILLER_7_186 ();
 sg13g2_fill_2 FILLER_7_200 ();
 sg13g2_fill_1 FILLER_7_207 ();
 sg13g2_decap_4 FILLER_7_243 ();
 sg13g2_fill_2 FILLER_7_247 ();
 sg13g2_fill_1 FILLER_7_253 ();
 sg13g2_fill_1 FILLER_7_271 ();
 sg13g2_decap_4 FILLER_7_277 ();
 sg13g2_fill_1 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_303 ();
 sg13g2_decap_4 FILLER_7_310 ();
 sg13g2_fill_2 FILLER_7_314 ();
 sg13g2_fill_1 FILLER_7_329 ();
 sg13g2_fill_2 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_fill_1 FILLER_7_372 ();
 sg13g2_decap_4 FILLER_7_378 ();
 sg13g2_fill_1 FILLER_7_382 ();
 sg13g2_fill_2 FILLER_7_388 ();
 sg13g2_fill_1 FILLER_7_390 ();
 sg13g2_fill_1 FILLER_7_395 ();
 sg13g2_fill_2 FILLER_7_410 ();
 sg13g2_fill_1 FILLER_7_412 ();
 sg13g2_fill_1 FILLER_7_442 ();
 sg13g2_fill_1 FILLER_7_452 ();
 sg13g2_fill_1 FILLER_7_473 ();
 sg13g2_fill_2 FILLER_7_478 ();
 sg13g2_fill_2 FILLER_7_484 ();
 sg13g2_fill_1 FILLER_7_486 ();
 sg13g2_decap_8 FILLER_7_495 ();
 sg13g2_decap_4 FILLER_7_502 ();
 sg13g2_fill_2 FILLER_7_506 ();
 sg13g2_fill_2 FILLER_7_516 ();
 sg13g2_fill_1 FILLER_7_518 ();
 sg13g2_decap_4 FILLER_7_523 ();
 sg13g2_fill_2 FILLER_7_527 ();
 sg13g2_fill_2 FILLER_7_545 ();
 sg13g2_fill_2 FILLER_7_558 ();
 sg13g2_fill_2 FILLER_7_582 ();
 sg13g2_fill_2 FILLER_7_589 ();
 sg13g2_fill_1 FILLER_7_617 ();
 sg13g2_fill_2 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_635 ();
 sg13g2_decap_4 FILLER_7_642 ();
 sg13g2_decap_8 FILLER_7_649 ();
 sg13g2_fill_2 FILLER_7_656 ();
 sg13g2_fill_1 FILLER_7_675 ();
 sg13g2_decap_4 FILLER_7_686 ();
 sg13g2_fill_2 FILLER_7_704 ();
 sg13g2_decap_8 FILLER_7_713 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_4 FILLER_7_749 ();
 sg13g2_fill_2 FILLER_7_757 ();
 sg13g2_fill_1 FILLER_7_763 ();
 sg13g2_fill_1 FILLER_7_769 ();
 sg13g2_fill_1 FILLER_7_775 ();
 sg13g2_fill_2 FILLER_7_784 ();
 sg13g2_fill_1 FILLER_7_789 ();
 sg13g2_fill_2 FILLER_7_817 ();
 sg13g2_fill_1 FILLER_7_834 ();
 sg13g2_decap_8 FILLER_7_844 ();
 sg13g2_decap_8 FILLER_7_851 ();
 sg13g2_decap_8 FILLER_7_858 ();
 sg13g2_decap_8 FILLER_7_865 ();
 sg13g2_decap_8 FILLER_7_872 ();
 sg13g2_decap_4 FILLER_7_879 ();
 sg13g2_fill_1 FILLER_7_883 ();
 sg13g2_decap_8 FILLER_7_908 ();
 sg13g2_decap_8 FILLER_7_915 ();
 sg13g2_decap_8 FILLER_7_922 ();
 sg13g2_decap_8 FILLER_7_929 ();
 sg13g2_fill_2 FILLER_7_936 ();
 sg13g2_fill_1 FILLER_7_938 ();
 sg13g2_fill_2 FILLER_7_945 ();
 sg13g2_decap_8 FILLER_7_966 ();
 sg13g2_decap_8 FILLER_7_973 ();
 sg13g2_decap_4 FILLER_7_984 ();
 sg13g2_decap_4 FILLER_7_993 ();
 sg13g2_fill_2 FILLER_7_1002 ();
 sg13g2_decap_4 FILLER_7_1008 ();
 sg13g2_decap_8 FILLER_7_1017 ();
 sg13g2_fill_2 FILLER_7_1028 ();
 sg13g2_fill_1 FILLER_7_1030 ();
 sg13g2_decap_8 FILLER_7_1036 ();
 sg13g2_decap_4 FILLER_7_1043 ();
 sg13g2_decap_4 FILLER_7_1081 ();
 sg13g2_fill_2 FILLER_7_1119 ();
 sg13g2_fill_1 FILLER_7_1121 ();
 sg13g2_decap_4 FILLER_7_1127 ();
 sg13g2_fill_1 FILLER_7_1131 ();
 sg13g2_fill_1 FILLER_7_1146 ();
 sg13g2_decap_8 FILLER_7_1152 ();
 sg13g2_decap_8 FILLER_7_1159 ();
 sg13g2_decap_8 FILLER_7_1166 ();
 sg13g2_decap_8 FILLER_7_1173 ();
 sg13g2_decap_4 FILLER_7_1183 ();
 sg13g2_fill_2 FILLER_7_1187 ();
 sg13g2_fill_1 FILLER_7_1218 ();
 sg13g2_fill_2 FILLER_7_1227 ();
 sg13g2_decap_8 FILLER_7_1234 ();
 sg13g2_fill_2 FILLER_7_1241 ();
 sg13g2_fill_1 FILLER_7_1243 ();
 sg13g2_fill_2 FILLER_7_1248 ();
 sg13g2_fill_1 FILLER_7_1250 ();
 sg13g2_decap_8 FILLER_7_1256 ();
 sg13g2_fill_1 FILLER_7_1263 ();
 sg13g2_fill_2 FILLER_7_1274 ();
 sg13g2_decap_8 FILLER_7_1281 ();
 sg13g2_fill_2 FILLER_7_1288 ();
 sg13g2_decap_4 FILLER_7_1294 ();
 sg13g2_fill_1 FILLER_7_1303 ();
 sg13g2_fill_2 FILLER_7_1314 ();
 sg13g2_fill_2 FILLER_7_1320 ();
 sg13g2_fill_2 FILLER_7_1337 ();
 sg13g2_decap_8 FILLER_7_1345 ();
 sg13g2_decap_8 FILLER_7_1352 ();
 sg13g2_fill_1 FILLER_7_1359 ();
 sg13g2_fill_1 FILLER_7_1374 ();
 sg13g2_decap_8 FILLER_7_1379 ();
 sg13g2_fill_2 FILLER_7_1386 ();
 sg13g2_fill_1 FILLER_7_1388 ();
 sg13g2_decap_8 FILLER_7_1404 ();
 sg13g2_decap_8 FILLER_7_1411 ();
 sg13g2_decap_8 FILLER_7_1418 ();
 sg13g2_decap_8 FILLER_7_1425 ();
 sg13g2_decap_4 FILLER_7_1432 ();
 sg13g2_fill_1 FILLER_7_1458 ();
 sg13g2_fill_2 FILLER_7_1472 ();
 sg13g2_fill_1 FILLER_7_1474 ();
 sg13g2_decap_4 FILLER_7_1485 ();
 sg13g2_decap_8 FILLER_7_1499 ();
 sg13g2_decap_4 FILLER_7_1506 ();
 sg13g2_decap_8 FILLER_7_1514 ();
 sg13g2_decap_8 FILLER_7_1521 ();
 sg13g2_decap_8 FILLER_7_1540 ();
 sg13g2_decap_8 FILLER_7_1547 ();
 sg13g2_fill_1 FILLER_7_1554 ();
 sg13g2_decap_8 FILLER_7_1559 ();
 sg13g2_decap_8 FILLER_7_1566 ();
 sg13g2_decap_8 FILLER_7_1573 ();
 sg13g2_fill_1 FILLER_7_1580 ();
 sg13g2_decap_8 FILLER_7_1585 ();
 sg13g2_decap_8 FILLER_7_1592 ();
 sg13g2_decap_8 FILLER_7_1599 ();
 sg13g2_decap_8 FILLER_7_1606 ();
 sg13g2_decap_8 FILLER_7_1613 ();
 sg13g2_decap_8 FILLER_7_1620 ();
 sg13g2_decap_8 FILLER_7_1627 ();
 sg13g2_decap_8 FILLER_7_1634 ();
 sg13g2_decap_8 FILLER_7_1641 ();
 sg13g2_decap_8 FILLER_7_1648 ();
 sg13g2_decap_8 FILLER_7_1655 ();
 sg13g2_decap_8 FILLER_7_1662 ();
 sg13g2_decap_8 FILLER_7_1669 ();
 sg13g2_decap_8 FILLER_7_1676 ();
 sg13g2_decap_8 FILLER_7_1683 ();
 sg13g2_decap_8 FILLER_7_1690 ();
 sg13g2_decap_8 FILLER_7_1697 ();
 sg13g2_decap_8 FILLER_7_1704 ();
 sg13g2_decap_8 FILLER_7_1711 ();
 sg13g2_decap_8 FILLER_7_1718 ();
 sg13g2_decap_8 FILLER_7_1725 ();
 sg13g2_decap_8 FILLER_7_1732 ();
 sg13g2_decap_8 FILLER_7_1739 ();
 sg13g2_decap_8 FILLER_7_1746 ();
 sg13g2_decap_8 FILLER_7_1753 ();
 sg13g2_decap_8 FILLER_7_1760 ();
 sg13g2_decap_8 FILLER_7_1767 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_fill_1 FILLER_8_70 ();
 sg13g2_fill_2 FILLER_8_75 ();
 sg13g2_fill_1 FILLER_8_123 ();
 sg13g2_fill_2 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_136 ();
 sg13g2_fill_2 FILLER_8_142 ();
 sg13g2_fill_2 FILLER_8_149 ();
 sg13g2_fill_2 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_162 ();
 sg13g2_fill_1 FILLER_8_164 ();
 sg13g2_decap_4 FILLER_8_169 ();
 sg13g2_fill_1 FILLER_8_173 ();
 sg13g2_fill_1 FILLER_8_179 ();
 sg13g2_fill_1 FILLER_8_213 ();
 sg13g2_decap_4 FILLER_8_232 ();
 sg13g2_fill_1 FILLER_8_236 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_fill_2 FILLER_8_256 ();
 sg13g2_fill_1 FILLER_8_258 ();
 sg13g2_decap_4 FILLER_8_264 ();
 sg13g2_fill_2 FILLER_8_278 ();
 sg13g2_fill_1 FILLER_8_297 ();
 sg13g2_fill_1 FILLER_8_305 ();
 sg13g2_fill_1 FILLER_8_315 ();
 sg13g2_fill_2 FILLER_8_353 ();
 sg13g2_fill_2 FILLER_8_363 ();
 sg13g2_fill_2 FILLER_8_382 ();
 sg13g2_fill_2 FILLER_8_388 ();
 sg13g2_decap_4 FILLER_8_411 ();
 sg13g2_fill_1 FILLER_8_445 ();
 sg13g2_fill_1 FILLER_8_459 ();
 sg13g2_fill_2 FILLER_8_472 ();
 sg13g2_fill_1 FILLER_8_474 ();
 sg13g2_decap_4 FILLER_8_483 ();
 sg13g2_fill_2 FILLER_8_487 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_508 ();
 sg13g2_decap_8 FILLER_8_515 ();
 sg13g2_decap_8 FILLER_8_522 ();
 sg13g2_decap_8 FILLER_8_529 ();
 sg13g2_fill_1 FILLER_8_536 ();
 sg13g2_fill_1 FILLER_8_603 ();
 sg13g2_fill_2 FILLER_8_617 ();
 sg13g2_fill_1 FILLER_8_640 ();
 sg13g2_fill_1 FILLER_8_645 ();
 sg13g2_fill_2 FILLER_8_657 ();
 sg13g2_decap_8 FILLER_8_678 ();
 sg13g2_decap_8 FILLER_8_685 ();
 sg13g2_decap_4 FILLER_8_692 ();
 sg13g2_decap_8 FILLER_8_731 ();
 sg13g2_decap_4 FILLER_8_738 ();
 sg13g2_fill_1 FILLER_8_742 ();
 sg13g2_fill_2 FILLER_8_759 ();
 sg13g2_fill_1 FILLER_8_778 ();
 sg13g2_fill_1 FILLER_8_810 ();
 sg13g2_fill_1 FILLER_8_819 ();
 sg13g2_fill_2 FILLER_8_826 ();
 sg13g2_fill_2 FILLER_8_832 ();
 sg13g2_decap_4 FILLER_8_844 ();
 sg13g2_fill_2 FILLER_8_848 ();
 sg13g2_fill_2 FILLER_8_854 ();
 sg13g2_fill_2 FILLER_8_871 ();
 sg13g2_fill_1 FILLER_8_873 ();
 sg13g2_decap_4 FILLER_8_887 ();
 sg13g2_fill_1 FILLER_8_903 ();
 sg13g2_fill_2 FILLER_8_926 ();
 sg13g2_fill_2 FILLER_8_945 ();
 sg13g2_fill_1 FILLER_8_947 ();
 sg13g2_decap_4 FILLER_8_954 ();
 sg13g2_fill_1 FILLER_8_958 ();
 sg13g2_decap_4 FILLER_8_968 ();
 sg13g2_fill_1 FILLER_8_972 ();
 sg13g2_decap_4 FILLER_8_978 ();
 sg13g2_fill_2 FILLER_8_982 ();
 sg13g2_decap_8 FILLER_8_988 ();
 sg13g2_fill_1 FILLER_8_1005 ();
 sg13g2_fill_1 FILLER_8_1012 ();
 sg13g2_decap_8 FILLER_8_1018 ();
 sg13g2_fill_2 FILLER_8_1025 ();
 sg13g2_decap_8 FILLER_8_1048 ();
 sg13g2_decap_4 FILLER_8_1055 ();
 sg13g2_decap_4 FILLER_8_1091 ();
 sg13g2_fill_2 FILLER_8_1095 ();
 sg13g2_decap_8 FILLER_8_1109 ();
 sg13g2_fill_1 FILLER_8_1116 ();
 sg13g2_fill_2 FILLER_8_1141 ();
 sg13g2_fill_1 FILLER_8_1143 ();
 sg13g2_decap_4 FILLER_8_1155 ();
 sg13g2_fill_2 FILLER_8_1159 ();
 sg13g2_decap_8 FILLER_8_1165 ();
 sg13g2_decap_8 FILLER_8_1172 ();
 sg13g2_decap_4 FILLER_8_1179 ();
 sg13g2_fill_1 FILLER_8_1183 ();
 sg13g2_fill_1 FILLER_8_1196 ();
 sg13g2_decap_4 FILLER_8_1202 ();
 sg13g2_fill_1 FILLER_8_1206 ();
 sg13g2_decap_8 FILLER_8_1216 ();
 sg13g2_decap_8 FILLER_8_1223 ();
 sg13g2_decap_8 FILLER_8_1230 ();
 sg13g2_fill_2 FILLER_8_1237 ();
 sg13g2_fill_1 FILLER_8_1239 ();
 sg13g2_fill_1 FILLER_8_1250 ();
 sg13g2_fill_2 FILLER_8_1256 ();
 sg13g2_fill_2 FILLER_8_1262 ();
 sg13g2_fill_2 FILLER_8_1269 ();
 sg13g2_fill_2 FILLER_8_1297 ();
 sg13g2_decap_4 FILLER_8_1304 ();
 sg13g2_decap_4 FILLER_8_1334 ();
 sg13g2_fill_1 FILLER_8_1347 ();
 sg13g2_fill_2 FILLER_8_1365 ();
 sg13g2_fill_2 FILLER_8_1384 ();
 sg13g2_fill_1 FILLER_8_1386 ();
 sg13g2_fill_2 FILLER_8_1397 ();
 sg13g2_fill_1 FILLER_8_1399 ();
 sg13g2_decap_8 FILLER_8_1426 ();
 sg13g2_fill_1 FILLER_8_1433 ();
 sg13g2_decap_4 FILLER_8_1484 ();
 sg13g2_fill_2 FILLER_8_1505 ();
 sg13g2_fill_1 FILLER_8_1513 ();
 sg13g2_decap_4 FILLER_8_1552 ();
 sg13g2_fill_2 FILLER_8_1556 ();
 sg13g2_decap_8 FILLER_8_1563 ();
 sg13g2_decap_8 FILLER_8_1570 ();
 sg13g2_decap_8 FILLER_8_1577 ();
 sg13g2_decap_8 FILLER_8_1584 ();
 sg13g2_decap_8 FILLER_8_1591 ();
 sg13g2_decap_8 FILLER_8_1598 ();
 sg13g2_decap_8 FILLER_8_1605 ();
 sg13g2_decap_8 FILLER_8_1612 ();
 sg13g2_decap_8 FILLER_8_1619 ();
 sg13g2_decap_8 FILLER_8_1626 ();
 sg13g2_decap_8 FILLER_8_1633 ();
 sg13g2_decap_8 FILLER_8_1640 ();
 sg13g2_decap_8 FILLER_8_1647 ();
 sg13g2_fill_2 FILLER_8_1654 ();
 sg13g2_decap_8 FILLER_8_1664 ();
 sg13g2_decap_8 FILLER_8_1671 ();
 sg13g2_decap_8 FILLER_8_1678 ();
 sg13g2_decap_8 FILLER_8_1685 ();
 sg13g2_decap_8 FILLER_8_1692 ();
 sg13g2_decap_8 FILLER_8_1699 ();
 sg13g2_decap_8 FILLER_8_1706 ();
 sg13g2_decap_8 FILLER_8_1713 ();
 sg13g2_decap_8 FILLER_8_1720 ();
 sg13g2_decap_8 FILLER_8_1727 ();
 sg13g2_decap_8 FILLER_8_1734 ();
 sg13g2_decap_8 FILLER_8_1741 ();
 sg13g2_decap_8 FILLER_8_1748 ();
 sg13g2_decap_8 FILLER_8_1755 ();
 sg13g2_decap_8 FILLER_8_1762 ();
 sg13g2_decap_4 FILLER_8_1769 ();
 sg13g2_fill_1 FILLER_8_1773 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_fill_2 FILLER_9_53 ();
 sg13g2_fill_1 FILLER_9_58 ();
 sg13g2_fill_2 FILLER_9_63 ();
 sg13g2_fill_1 FILLER_9_70 ();
 sg13g2_fill_1 FILLER_9_76 ();
 sg13g2_fill_1 FILLER_9_85 ();
 sg13g2_fill_2 FILLER_9_117 ();
 sg13g2_fill_2 FILLER_9_129 ();
 sg13g2_fill_1 FILLER_9_137 ();
 sg13g2_fill_2 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_150 ();
 sg13g2_fill_2 FILLER_9_199 ();
 sg13g2_fill_2 FILLER_9_206 ();
 sg13g2_fill_1 FILLER_9_212 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_fill_1 FILLER_9_286 ();
 sg13g2_fill_1 FILLER_9_295 ();
 sg13g2_fill_2 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_376 ();
 sg13g2_fill_2 FILLER_9_391 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_fill_1 FILLER_9_409 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_4 FILLER_9_461 ();
 sg13g2_fill_2 FILLER_9_465 ();
 sg13g2_decap_8 FILLER_9_487 ();
 sg13g2_fill_1 FILLER_9_494 ();
 sg13g2_decap_8 FILLER_9_521 ();
 sg13g2_fill_2 FILLER_9_528 ();
 sg13g2_fill_1 FILLER_9_567 ();
 sg13g2_fill_2 FILLER_9_588 ();
 sg13g2_fill_1 FILLER_9_594 ();
 sg13g2_fill_2 FILLER_9_620 ();
 sg13g2_fill_1 FILLER_9_628 ();
 sg13g2_fill_1 FILLER_9_667 ();
 sg13g2_fill_1 FILLER_9_673 ();
 sg13g2_decap_4 FILLER_9_695 ();
 sg13g2_fill_2 FILLER_9_699 ();
 sg13g2_decap_8 FILLER_9_706 ();
 sg13g2_fill_2 FILLER_9_721 ();
 sg13g2_fill_1 FILLER_9_740 ();
 sg13g2_fill_2 FILLER_9_749 ();
 sg13g2_fill_2 FILLER_9_784 ();
 sg13g2_fill_1 FILLER_9_786 ();
 sg13g2_fill_2 FILLER_9_795 ();
 sg13g2_fill_1 FILLER_9_815 ();
 sg13g2_decap_8 FILLER_9_823 ();
 sg13g2_fill_1 FILLER_9_830 ();
 sg13g2_decap_4 FILLER_9_865 ();
 sg13g2_fill_1 FILLER_9_883 ();
 sg13g2_decap_4 FILLER_9_909 ();
 sg13g2_fill_1 FILLER_9_913 ();
 sg13g2_fill_2 FILLER_9_927 ();
 sg13g2_decap_8 FILLER_9_933 ();
 sg13g2_fill_2 FILLER_9_948 ();
 sg13g2_fill_1 FILLER_9_950 ();
 sg13g2_fill_2 FILLER_9_977 ();
 sg13g2_fill_1 FILLER_9_979 ();
 sg13g2_decap_4 FILLER_9_1004 ();
 sg13g2_fill_2 FILLER_9_1013 ();
 sg13g2_decap_8 FILLER_9_1027 ();
 sg13g2_fill_2 FILLER_9_1034 ();
 sg13g2_fill_1 FILLER_9_1036 ();
 sg13g2_fill_2 FILLER_9_1062 ();
 sg13g2_decap_4 FILLER_9_1088 ();
 sg13g2_fill_2 FILLER_9_1092 ();
 sg13g2_decap_4 FILLER_9_1115 ();
 sg13g2_fill_1 FILLER_9_1124 ();
 sg13g2_decap_8 FILLER_9_1145 ();
 sg13g2_decap_8 FILLER_9_1152 ();
 sg13g2_decap_8 FILLER_9_1159 ();
 sg13g2_fill_1 FILLER_9_1166 ();
 sg13g2_fill_1 FILLER_9_1172 ();
 sg13g2_fill_1 FILLER_9_1189 ();
 sg13g2_fill_1 FILLER_9_1195 ();
 sg13g2_fill_1 FILLER_9_1242 ();
 sg13g2_fill_2 FILLER_9_1262 ();
 sg13g2_decap_8 FILLER_9_1290 ();
 sg13g2_decap_4 FILLER_9_1297 ();
 sg13g2_fill_2 FILLER_9_1301 ();
 sg13g2_decap_8 FILLER_9_1311 ();
 sg13g2_fill_2 FILLER_9_1318 ();
 sg13g2_fill_1 FILLER_9_1320 ();
 sg13g2_fill_2 FILLER_9_1333 ();
 sg13g2_fill_1 FILLER_9_1335 ();
 sg13g2_fill_1 FILLER_9_1340 ();
 sg13g2_fill_2 FILLER_9_1372 ();
 sg13g2_fill_1 FILLER_9_1374 ();
 sg13g2_decap_4 FILLER_9_1379 ();
 sg13g2_fill_2 FILLER_9_1383 ();
 sg13g2_fill_1 FILLER_9_1392 ();
 sg13g2_decap_8 FILLER_9_1425 ();
 sg13g2_fill_1 FILLER_9_1456 ();
 sg13g2_decap_4 FILLER_9_1462 ();
 sg13g2_fill_2 FILLER_9_1466 ();
 sg13g2_fill_2 FILLER_9_1475 ();
 sg13g2_fill_1 FILLER_9_1494 ();
 sg13g2_fill_1 FILLER_9_1505 ();
 sg13g2_decap_4 FILLER_9_1536 ();
 sg13g2_fill_2 FILLER_9_1559 ();
 sg13g2_fill_1 FILLER_9_1561 ();
 sg13g2_decap_8 FILLER_9_1570 ();
 sg13g2_decap_8 FILLER_9_1577 ();
 sg13g2_decap_8 FILLER_9_1584 ();
 sg13g2_decap_8 FILLER_9_1596 ();
 sg13g2_decap_4 FILLER_9_1603 ();
 sg13g2_fill_1 FILLER_9_1607 ();
 sg13g2_decap_8 FILLER_9_1613 ();
 sg13g2_decap_8 FILLER_9_1620 ();
 sg13g2_decap_8 FILLER_9_1627 ();
 sg13g2_decap_4 FILLER_9_1634 ();
 sg13g2_decap_8 FILLER_9_1643 ();
 sg13g2_decap_8 FILLER_9_1650 ();
 sg13g2_decap_4 FILLER_9_1657 ();
 sg13g2_decap_8 FILLER_9_1665 ();
 sg13g2_decap_8 FILLER_9_1672 ();
 sg13g2_decap_8 FILLER_9_1679 ();
 sg13g2_decap_8 FILLER_9_1686 ();
 sg13g2_decap_8 FILLER_9_1693 ();
 sg13g2_decap_8 FILLER_9_1700 ();
 sg13g2_decap_8 FILLER_9_1707 ();
 sg13g2_decap_8 FILLER_9_1714 ();
 sg13g2_decap_8 FILLER_9_1721 ();
 sg13g2_decap_8 FILLER_9_1728 ();
 sg13g2_decap_8 FILLER_9_1735 ();
 sg13g2_decap_8 FILLER_9_1742 ();
 sg13g2_decap_8 FILLER_9_1749 ();
 sg13g2_decap_8 FILLER_9_1756 ();
 sg13g2_decap_8 FILLER_9_1763 ();
 sg13g2_decap_4 FILLER_9_1770 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_fill_1 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_31 ();
 sg13g2_decap_8 FILLER_10_38 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_fill_1 FILLER_10_71 ();
 sg13g2_fill_1 FILLER_10_89 ();
 sg13g2_fill_2 FILLER_10_104 ();
 sg13g2_decap_4 FILLER_10_173 ();
 sg13g2_fill_1 FILLER_10_177 ();
 sg13g2_fill_2 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_202 ();
 sg13g2_fill_2 FILLER_10_220 ();
 sg13g2_fill_1 FILLER_10_222 ();
 sg13g2_fill_1 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_247 ();
 sg13g2_decap_8 FILLER_10_251 ();
 sg13g2_fill_2 FILLER_10_258 ();
 sg13g2_fill_2 FILLER_10_285 ();
 sg13g2_decap_4 FILLER_10_295 ();
 sg13g2_decap_4 FILLER_10_311 ();
 sg13g2_fill_1 FILLER_10_315 ();
 sg13g2_fill_2 FILLER_10_349 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_388 ();
 sg13g2_decap_4 FILLER_10_410 ();
 sg13g2_fill_2 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_449 ();
 sg13g2_fill_2 FILLER_10_456 ();
 sg13g2_fill_1 FILLER_10_458 ();
 sg13g2_fill_2 FILLER_10_476 ();
 sg13g2_fill_1 FILLER_10_478 ();
 sg13g2_decap_4 FILLER_10_486 ();
 sg13g2_fill_1 FILLER_10_490 ();
 sg13g2_fill_2 FILLER_10_496 ();
 sg13g2_decap_8 FILLER_10_502 ();
 sg13g2_decap_8 FILLER_10_509 ();
 sg13g2_decap_8 FILLER_10_516 ();
 sg13g2_fill_2 FILLER_10_523 ();
 sg13g2_fill_1 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_533 ();
 sg13g2_fill_1 FILLER_10_553 ();
 sg13g2_fill_1 FILLER_10_567 ();
 sg13g2_fill_1 FILLER_10_593 ();
 sg13g2_fill_1 FILLER_10_631 ();
 sg13g2_decap_8 FILLER_10_636 ();
 sg13g2_fill_1 FILLER_10_643 ();
 sg13g2_fill_2 FILLER_10_663 ();
 sg13g2_fill_1 FILLER_10_681 ();
 sg13g2_fill_1 FILLER_10_690 ();
 sg13g2_fill_1 FILLER_10_699 ();
 sg13g2_decap_4 FILLER_10_708 ();
 sg13g2_decap_8 FILLER_10_733 ();
 sg13g2_fill_2 FILLER_10_740 ();
 sg13g2_decap_4 FILLER_10_763 ();
 sg13g2_decap_4 FILLER_10_776 ();
 sg13g2_fill_1 FILLER_10_780 ();
 sg13g2_fill_2 FILLER_10_799 ();
 sg13g2_fill_1 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_825 ();
 sg13g2_decap_8 FILLER_10_832 ();
 sg13g2_decap_4 FILLER_10_839 ();
 sg13g2_fill_1 FILLER_10_843 ();
 sg13g2_decap_8 FILLER_10_853 ();
 sg13g2_decap_4 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_10_897 ();
 sg13g2_fill_1 FILLER_10_904 ();
 sg13g2_decap_4 FILLER_10_916 ();
 sg13g2_fill_1 FILLER_10_920 ();
 sg13g2_fill_2 FILLER_10_926 ();
 sg13g2_fill_1 FILLER_10_928 ();
 sg13g2_fill_2 FILLER_10_933 ();
 sg13g2_decap_4 FILLER_10_940 ();
 sg13g2_fill_1 FILLER_10_944 ();
 sg13g2_decap_4 FILLER_10_953 ();
 sg13g2_fill_1 FILLER_10_957 ();
 sg13g2_fill_2 FILLER_10_968 ();
 sg13g2_fill_1 FILLER_10_1004 ();
 sg13g2_decap_4 FILLER_10_1015 ();
 sg13g2_fill_2 FILLER_10_1019 ();
 sg13g2_decap_4 FILLER_10_1029 ();
 sg13g2_fill_2 FILLER_10_1049 ();
 sg13g2_fill_1 FILLER_10_1051 ();
 sg13g2_fill_1 FILLER_10_1057 ();
 sg13g2_decap_8 FILLER_10_1062 ();
 sg13g2_fill_1 FILLER_10_1069 ();
 sg13g2_fill_2 FILLER_10_1079 ();
 sg13g2_decap_8 FILLER_10_1085 ();
 sg13g2_decap_8 FILLER_10_1092 ();
 sg13g2_fill_2 FILLER_10_1099 ();
 sg13g2_fill_1 FILLER_10_1101 ();
 sg13g2_decap_8 FILLER_10_1118 ();
 sg13g2_decap_8 FILLER_10_1138 ();
 sg13g2_decap_8 FILLER_10_1145 ();
 sg13g2_fill_2 FILLER_10_1152 ();
 sg13g2_fill_1 FILLER_10_1165 ();
 sg13g2_decap_8 FILLER_10_1182 ();
 sg13g2_decap_4 FILLER_10_1220 ();
 sg13g2_fill_1 FILLER_10_1224 ();
 sg13g2_decap_8 FILLER_10_1233 ();
 sg13g2_decap_8 FILLER_10_1240 ();
 sg13g2_decap_8 FILLER_10_1247 ();
 sg13g2_fill_2 FILLER_10_1254 ();
 sg13g2_decap_4 FILLER_10_1265 ();
 sg13g2_fill_1 FILLER_10_1269 ();
 sg13g2_decap_8 FILLER_10_1274 ();
 sg13g2_decap_8 FILLER_10_1281 ();
 sg13g2_fill_1 FILLER_10_1288 ();
 sg13g2_fill_2 FILLER_10_1297 ();
 sg13g2_fill_1 FILLER_10_1329 ();
 sg13g2_decap_8 FILLER_10_1335 ();
 sg13g2_decap_4 FILLER_10_1342 ();
 sg13g2_fill_2 FILLER_10_1346 ();
 sg13g2_fill_2 FILLER_10_1352 ();
 sg13g2_decap_8 FILLER_10_1361 ();
 sg13g2_decap_4 FILLER_10_1376 ();
 sg13g2_fill_1 FILLER_10_1380 ();
 sg13g2_decap_4 FILLER_10_1384 ();
 sg13g2_fill_1 FILLER_10_1410 ();
 sg13g2_decap_8 FILLER_10_1432 ();
 sg13g2_fill_1 FILLER_10_1444 ();
 sg13g2_fill_1 FILLER_10_1470 ();
 sg13g2_fill_1 FILLER_10_1479 ();
 sg13g2_fill_1 FILLER_10_1515 ();
 sg13g2_fill_2 FILLER_10_1551 ();
 sg13g2_fill_1 FILLER_10_1566 ();
 sg13g2_decap_8 FILLER_10_1593 ();
 sg13g2_decap_4 FILLER_10_1600 ();
 sg13g2_fill_2 FILLER_10_1604 ();
 sg13g2_decap_8 FILLER_10_1614 ();
 sg13g2_decap_8 FILLER_10_1621 ();
 sg13g2_decap_4 FILLER_10_1628 ();
 sg13g2_decap_8 FILLER_10_1636 ();
 sg13g2_decap_8 FILLER_10_1643 ();
 sg13g2_decap_8 FILLER_10_1650 ();
 sg13g2_decap_4 FILLER_10_1657 ();
 sg13g2_fill_1 FILLER_10_1661 ();
 sg13g2_decap_8 FILLER_10_1667 ();
 sg13g2_decap_8 FILLER_10_1674 ();
 sg13g2_decap_8 FILLER_10_1681 ();
 sg13g2_decap_8 FILLER_10_1688 ();
 sg13g2_decap_8 FILLER_10_1695 ();
 sg13g2_decap_8 FILLER_10_1702 ();
 sg13g2_decap_8 FILLER_10_1709 ();
 sg13g2_decap_4 FILLER_10_1716 ();
 sg13g2_fill_1 FILLER_10_1720 ();
 sg13g2_decap_8 FILLER_10_1725 ();
 sg13g2_decap_8 FILLER_10_1732 ();
 sg13g2_decap_8 FILLER_10_1739 ();
 sg13g2_decap_8 FILLER_10_1746 ();
 sg13g2_decap_8 FILLER_10_1753 ();
 sg13g2_decap_8 FILLER_10_1760 ();
 sg13g2_decap_8 FILLER_10_1767 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_fill_2 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_44 ();
 sg13g2_fill_2 FILLER_11_50 ();
 sg13g2_decap_4 FILLER_11_57 ();
 sg13g2_fill_2 FILLER_11_61 ();
 sg13g2_fill_1 FILLER_11_67 ();
 sg13g2_fill_2 FILLER_11_72 ();
 sg13g2_fill_1 FILLER_11_114 ();
 sg13g2_fill_2 FILLER_11_177 ();
 sg13g2_fill_2 FILLER_11_192 ();
 sg13g2_decap_8 FILLER_11_198 ();
 sg13g2_decap_8 FILLER_11_205 ();
 sg13g2_decap_8 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_219 ();
 sg13g2_decap_8 FILLER_11_230 ();
 sg13g2_decap_4 FILLER_11_237 ();
 sg13g2_fill_1 FILLER_11_241 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_decap_4 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_276 ();
 sg13g2_fill_2 FILLER_11_293 ();
 sg13g2_fill_1 FILLER_11_295 ();
 sg13g2_fill_1 FILLER_11_299 ();
 sg13g2_fill_1 FILLER_11_358 ();
 sg13g2_fill_2 FILLER_11_380 ();
 sg13g2_fill_2 FILLER_11_385 ();
 sg13g2_fill_1 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_fill_2 FILLER_11_417 ();
 sg13g2_fill_1 FILLER_11_419 ();
 sg13g2_fill_1 FILLER_11_425 ();
 sg13g2_fill_2 FILLER_11_456 ();
 sg13g2_fill_1 FILLER_11_476 ();
 sg13g2_fill_2 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_510 ();
 sg13g2_decap_4 FILLER_11_517 ();
 sg13g2_decap_4 FILLER_11_547 ();
 sg13g2_fill_1 FILLER_11_554 ();
 sg13g2_fill_2 FILLER_11_571 ();
 sg13g2_fill_2 FILLER_11_577 ();
 sg13g2_fill_1 FILLER_11_599 ();
 sg13g2_fill_2 FILLER_11_608 ();
 sg13g2_fill_1 FILLER_11_651 ();
 sg13g2_fill_2 FILLER_11_655 ();
 sg13g2_fill_1 FILLER_11_668 ();
 sg13g2_fill_1 FILLER_11_673 ();
 sg13g2_decap_4 FILLER_11_687 ();
 sg13g2_decap_8 FILLER_11_695 ();
 sg13g2_fill_1 FILLER_11_719 ();
 sg13g2_fill_1 FILLER_11_731 ();
 sg13g2_decap_4 FILLER_11_758 ();
 sg13g2_fill_1 FILLER_11_766 ();
 sg13g2_fill_2 FILLER_11_778 ();
 sg13g2_fill_1 FILLER_11_780 ();
 sg13g2_fill_1 FILLER_11_803 ();
 sg13g2_fill_1 FILLER_11_812 ();
 sg13g2_fill_1 FILLER_11_818 ();
 sg13g2_fill_2 FILLER_11_823 ();
 sg13g2_fill_2 FILLER_11_833 ();
 sg13g2_decap_4 FILLER_11_840 ();
 sg13g2_fill_2 FILLER_11_844 ();
 sg13g2_decap_4 FILLER_11_850 ();
 sg13g2_fill_1 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_872 ();
 sg13g2_fill_1 FILLER_11_881 ();
 sg13g2_fill_1 FILLER_11_932 ();
 sg13g2_decap_4 FILLER_11_955 ();
 sg13g2_fill_2 FILLER_11_959 ();
 sg13g2_decap_8 FILLER_11_969 ();
 sg13g2_fill_1 FILLER_11_976 ();
 sg13g2_decap_4 FILLER_11_987 ();
 sg13g2_fill_1 FILLER_11_991 ();
 sg13g2_decap_8 FILLER_11_1014 ();
 sg13g2_fill_2 FILLER_11_1036 ();
 sg13g2_decap_4 FILLER_11_1043 ();
 sg13g2_fill_2 FILLER_11_1096 ();
 sg13g2_fill_1 FILLER_11_1098 ();
 sg13g2_fill_2 FILLER_11_1104 ();
 sg13g2_fill_1 FILLER_11_1106 ();
 sg13g2_fill_1 FILLER_11_1117 ();
 sg13g2_fill_1 FILLER_11_1124 ();
 sg13g2_decap_4 FILLER_11_1141 ();
 sg13g2_fill_1 FILLER_11_1145 ();
 sg13g2_decap_8 FILLER_11_1154 ();
 sg13g2_decap_4 FILLER_11_1161 ();
 sg13g2_fill_1 FILLER_11_1165 ();
 sg13g2_decap_8 FILLER_11_1195 ();
 sg13g2_fill_1 FILLER_11_1202 ();
 sg13g2_decap_4 FILLER_11_1219 ();
 sg13g2_fill_1 FILLER_11_1223 ();
 sg13g2_fill_1 FILLER_11_1237 ();
 sg13g2_decap_4 FILLER_11_1246 ();
 sg13g2_decap_8 FILLER_11_1271 ();
 sg13g2_decap_8 FILLER_11_1278 ();
 sg13g2_fill_1 FILLER_11_1285 ();
 sg13g2_fill_2 FILLER_11_1289 ();
 sg13g2_decap_8 FILLER_11_1328 ();
 sg13g2_decap_4 FILLER_11_1335 ();
 sg13g2_fill_2 FILLER_11_1339 ();
 sg13g2_fill_2 FILLER_11_1357 ();
 sg13g2_decap_8 FILLER_11_1367 ();
 sg13g2_fill_1 FILLER_11_1374 ();
 sg13g2_decap_4 FILLER_11_1379 ();
 sg13g2_fill_1 FILLER_11_1414 ();
 sg13g2_fill_1 FILLER_11_1420 ();
 sg13g2_decap_8 FILLER_11_1438 ();
 sg13g2_decap_8 FILLER_11_1445 ();
 sg13g2_fill_2 FILLER_11_1469 ();
 sg13g2_fill_1 FILLER_11_1483 ();
 sg13g2_fill_2 FILLER_11_1517 ();
 sg13g2_fill_1 FILLER_11_1524 ();
 sg13g2_fill_2 FILLER_11_1534 ();
 sg13g2_fill_1 FILLER_11_1558 ();
 sg13g2_fill_1 FILLER_11_1570 ();
 sg13g2_decap_8 FILLER_11_1580 ();
 sg13g2_fill_1 FILLER_11_1587 ();
 sg13g2_decap_8 FILLER_11_1592 ();
 sg13g2_decap_8 FILLER_11_1599 ();
 sg13g2_decap_4 FILLER_11_1606 ();
 sg13g2_fill_1 FILLER_11_1610 ();
 sg13g2_decap_8 FILLER_11_1615 ();
 sg13g2_decap_8 FILLER_11_1622 ();
 sg13g2_decap_8 FILLER_11_1629 ();
 sg13g2_decap_8 FILLER_11_1636 ();
 sg13g2_fill_2 FILLER_11_1643 ();
 sg13g2_fill_1 FILLER_11_1645 ();
 sg13g2_decap_4 FILLER_11_1651 ();
 sg13g2_fill_1 FILLER_11_1655 ();
 sg13g2_fill_1 FILLER_11_1661 ();
 sg13g2_decap_8 FILLER_11_1666 ();
 sg13g2_decap_8 FILLER_11_1673 ();
 sg13g2_decap_8 FILLER_11_1680 ();
 sg13g2_decap_8 FILLER_11_1687 ();
 sg13g2_decap_8 FILLER_11_1694 ();
 sg13g2_decap_8 FILLER_11_1701 ();
 sg13g2_decap_8 FILLER_11_1708 ();
 sg13g2_decap_8 FILLER_11_1715 ();
 sg13g2_decap_8 FILLER_11_1722 ();
 sg13g2_decap_8 FILLER_11_1729 ();
 sg13g2_decap_8 FILLER_11_1736 ();
 sg13g2_decap_8 FILLER_11_1743 ();
 sg13g2_decap_8 FILLER_11_1750 ();
 sg13g2_decap_8 FILLER_11_1757 ();
 sg13g2_decap_8 FILLER_11_1764 ();
 sg13g2_fill_2 FILLER_11_1771 ();
 sg13g2_fill_1 FILLER_11_1773 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_25 ();
 sg13g2_decap_4 FILLER_12_57 ();
 sg13g2_fill_1 FILLER_12_61 ();
 sg13g2_fill_1 FILLER_12_67 ();
 sg13g2_fill_1 FILLER_12_76 ();
 sg13g2_fill_1 FILLER_12_89 ();
 sg13g2_fill_1 FILLER_12_119 ();
 sg13g2_fill_1 FILLER_12_134 ();
 sg13g2_fill_1 FILLER_12_150 ();
 sg13g2_fill_2 FILLER_12_181 ();
 sg13g2_decap_4 FILLER_12_220 ();
 sg13g2_fill_2 FILLER_12_224 ();
 sg13g2_fill_1 FILLER_12_231 ();
 sg13g2_fill_2 FILLER_12_252 ();
 sg13g2_fill_2 FILLER_12_259 ();
 sg13g2_fill_2 FILLER_12_265 ();
 sg13g2_fill_1 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_fill_2 FILLER_12_323 ();
 sg13g2_fill_1 FILLER_12_325 ();
 sg13g2_fill_2 FILLER_12_336 ();
 sg13g2_fill_1 FILLER_12_349 ();
 sg13g2_fill_2 FILLER_12_373 ();
 sg13g2_fill_2 FILLER_12_388 ();
 sg13g2_fill_1 FILLER_12_393 ();
 sg13g2_fill_2 FILLER_12_413 ();
 sg13g2_fill_2 FILLER_12_419 ();
 sg13g2_decap_8 FILLER_12_431 ();
 sg13g2_decap_8 FILLER_12_438 ();
 sg13g2_fill_1 FILLER_12_445 ();
 sg13g2_decap_8 FILLER_12_477 ();
 sg13g2_fill_2 FILLER_12_484 ();
 sg13g2_decap_8 FILLER_12_500 ();
 sg13g2_fill_1 FILLER_12_507 ();
 sg13g2_decap_4 FILLER_12_516 ();
 sg13g2_fill_2 FILLER_12_520 ();
 sg13g2_decap_8 FILLER_12_538 ();
 sg13g2_decap_8 FILLER_12_545 ();
 sg13g2_decap_8 FILLER_12_556 ();
 sg13g2_fill_2 FILLER_12_570 ();
 sg13g2_decap_4 FILLER_12_597 ();
 sg13g2_fill_1 FILLER_12_612 ();
 sg13g2_decap_4 FILLER_12_657 ();
 sg13g2_fill_1 FILLER_12_661 ();
 sg13g2_decap_4 FILLER_12_666 ();
 sg13g2_decap_4 FILLER_12_697 ();
 sg13g2_fill_1 FILLER_12_701 ();
 sg13g2_decap_4 FILLER_12_710 ();
 sg13g2_decap_4 FILLER_12_719 ();
 sg13g2_fill_1 FILLER_12_723 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_fill_1 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_740 ();
 sg13g2_decap_8 FILLER_12_747 ();
 sg13g2_decap_4 FILLER_12_754 ();
 sg13g2_fill_1 FILLER_12_758 ();
 sg13g2_fill_1 FILLER_12_764 ();
 sg13g2_fill_2 FILLER_12_770 ();
 sg13g2_fill_2 FILLER_12_808 ();
 sg13g2_fill_1 FILLER_12_816 ();
 sg13g2_fill_1 FILLER_12_827 ();
 sg13g2_fill_2 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_842 ();
 sg13g2_fill_2 FILLER_12_849 ();
 sg13g2_fill_1 FILLER_12_851 ();
 sg13g2_decap_4 FILLER_12_860 ();
 sg13g2_fill_1 FILLER_12_868 ();
 sg13g2_decap_4 FILLER_12_874 ();
 sg13g2_fill_2 FILLER_12_887 ();
 sg13g2_fill_1 FILLER_12_894 ();
 sg13g2_fill_2 FILLER_12_899 ();
 sg13g2_fill_2 FILLER_12_934 ();
 sg13g2_decap_8 FILLER_12_947 ();
 sg13g2_fill_1 FILLER_12_954 ();
 sg13g2_decap_8 FILLER_12_960 ();
 sg13g2_decap_8 FILLER_12_967 ();
 sg13g2_fill_2 FILLER_12_974 ();
 sg13g2_decap_4 FILLER_12_987 ();
 sg13g2_fill_1 FILLER_12_991 ();
 sg13g2_fill_2 FILLER_12_1000 ();
 sg13g2_decap_8 FILLER_12_1007 ();
 sg13g2_decap_8 FILLER_12_1014 ();
 sg13g2_fill_2 FILLER_12_1021 ();
 sg13g2_fill_1 FILLER_12_1023 ();
 sg13g2_decap_8 FILLER_12_1037 ();
 sg13g2_decap_4 FILLER_12_1044 ();
 sg13g2_fill_2 FILLER_12_1048 ();
 sg13g2_decap_8 FILLER_12_1065 ();
 sg13g2_decap_8 FILLER_12_1072 ();
 sg13g2_fill_2 FILLER_12_1079 ();
 sg13g2_fill_2 FILLER_12_1125 ();
 sg13g2_fill_1 FILLER_12_1141 ();
 sg13g2_decap_8 FILLER_12_1151 ();
 sg13g2_decap_4 FILLER_12_1158 ();
 sg13g2_fill_1 FILLER_12_1162 ();
 sg13g2_decap_4 FILLER_12_1167 ();
 sg13g2_fill_2 FILLER_12_1176 ();
 sg13g2_fill_2 FILLER_12_1183 ();
 sg13g2_decap_8 FILLER_12_1219 ();
 sg13g2_decap_4 FILLER_12_1226 ();
 sg13g2_fill_2 FILLER_12_1230 ();
 sg13g2_fill_1 FILLER_12_1237 ();
 sg13g2_fill_2 FILLER_12_1257 ();
 sg13g2_decap_8 FILLER_12_1263 ();
 sg13g2_decap_4 FILLER_12_1278 ();
 sg13g2_fill_2 FILLER_12_1287 ();
 sg13g2_fill_1 FILLER_12_1289 ();
 sg13g2_decap_8 FILLER_12_1295 ();
 sg13g2_fill_1 FILLER_12_1302 ();
 sg13g2_fill_2 FILLER_12_1339 ();
 sg13g2_fill_1 FILLER_12_1351 ();
 sg13g2_decap_8 FILLER_12_1372 ();
 sg13g2_decap_4 FILLER_12_1379 ();
 sg13g2_fill_2 FILLER_12_1383 ();
 sg13g2_decap_4 FILLER_12_1389 ();
 sg13g2_fill_2 FILLER_12_1396 ();
 sg13g2_fill_1 FILLER_12_1398 ();
 sg13g2_fill_1 FILLER_12_1408 ();
 sg13g2_fill_1 FILLER_12_1423 ();
 sg13g2_fill_2 FILLER_12_1430 ();
 sg13g2_fill_1 FILLER_12_1432 ();
 sg13g2_decap_8 FILLER_12_1438 ();
 sg13g2_fill_1 FILLER_12_1465 ();
 sg13g2_fill_2 FILLER_12_1498 ();
 sg13g2_fill_1 FILLER_12_1534 ();
 sg13g2_fill_1 FILLER_12_1549 ();
 sg13g2_fill_2 FILLER_12_1556 ();
 sg13g2_fill_1 FILLER_12_1566 ();
 sg13g2_fill_2 FILLER_12_1577 ();
 sg13g2_decap_8 FILLER_12_1584 ();
 sg13g2_fill_1 FILLER_12_1591 ();
 sg13g2_decap_4 FILLER_12_1609 ();
 sg13g2_fill_2 FILLER_12_1622 ();
 sg13g2_fill_2 FILLER_12_1634 ();
 sg13g2_fill_1 FILLER_12_1636 ();
 sg13g2_fill_1 FILLER_12_1644 ();
 sg13g2_fill_2 FILLER_12_1650 ();
 sg13g2_fill_2 FILLER_12_1662 ();
 sg13g2_decap_8 FILLER_12_1668 ();
 sg13g2_decap_8 FILLER_12_1675 ();
 sg13g2_decap_8 FILLER_12_1682 ();
 sg13g2_decap_8 FILLER_12_1689 ();
 sg13g2_decap_8 FILLER_12_1696 ();
 sg13g2_decap_8 FILLER_12_1703 ();
 sg13g2_decap_8 FILLER_12_1710 ();
 sg13g2_decap_8 FILLER_12_1717 ();
 sg13g2_decap_8 FILLER_12_1724 ();
 sg13g2_decap_8 FILLER_12_1731 ();
 sg13g2_decap_8 FILLER_12_1738 ();
 sg13g2_decap_8 FILLER_12_1745 ();
 sg13g2_decap_8 FILLER_12_1752 ();
 sg13g2_decap_8 FILLER_12_1759 ();
 sg13g2_decap_8 FILLER_12_1766 ();
 sg13g2_fill_1 FILLER_12_1773 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_37 ();
 sg13g2_decap_8 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_51 ();
 sg13g2_fill_2 FILLER_13_56 ();
 sg13g2_fill_2 FILLER_13_66 ();
 sg13g2_fill_2 FILLER_13_95 ();
 sg13g2_fill_2 FILLER_13_118 ();
 sg13g2_fill_1 FILLER_13_128 ();
 sg13g2_fill_2 FILLER_13_179 ();
 sg13g2_fill_1 FILLER_13_191 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_fill_2 FILLER_13_271 ();
 sg13g2_fill_2 FILLER_13_333 ();
 sg13g2_fill_1 FILLER_13_335 ();
 sg13g2_fill_1 FILLER_13_341 ();
 sg13g2_fill_2 FILLER_13_346 ();
 sg13g2_fill_1 FILLER_13_348 ();
 sg13g2_fill_1 FILLER_13_353 ();
 sg13g2_fill_1 FILLER_13_359 ();
 sg13g2_fill_1 FILLER_13_375 ();
 sg13g2_fill_2 FILLER_13_380 ();
 sg13g2_fill_2 FILLER_13_390 ();
 sg13g2_fill_1 FILLER_13_398 ();
 sg13g2_fill_2 FILLER_13_404 ();
 sg13g2_decap_8 FILLER_13_436 ();
 sg13g2_decap_8 FILLER_13_443 ();
 sg13g2_decap_4 FILLER_13_450 ();
 sg13g2_fill_2 FILLER_13_462 ();
 sg13g2_fill_1 FILLER_13_464 ();
 sg13g2_decap_8 FILLER_13_479 ();
 sg13g2_decap_4 FILLER_13_486 ();
 sg13g2_fill_2 FILLER_13_490 ();
 sg13g2_decap_4 FILLER_13_495 ();
 sg13g2_fill_1 FILLER_13_499 ();
 sg13g2_fill_2 FILLER_13_503 ();
 sg13g2_fill_1 FILLER_13_505 ();
 sg13g2_decap_4 FILLER_13_511 ();
 sg13g2_fill_1 FILLER_13_515 ();
 sg13g2_decap_4 FILLER_13_529 ();
 sg13g2_fill_2 FILLER_13_533 ();
 sg13g2_decap_8 FILLER_13_543 ();
 sg13g2_fill_2 FILLER_13_550 ();
 sg13g2_decap_4 FILLER_13_599 ();
 sg13g2_fill_2 FILLER_13_611 ();
 sg13g2_fill_1 FILLER_13_636 ();
 sg13g2_fill_1 FILLER_13_641 ();
 sg13g2_decap_4 FILLER_13_650 ();
 sg13g2_fill_2 FILLER_13_654 ();
 sg13g2_fill_1 FILLER_13_668 ();
 sg13g2_fill_2 FILLER_13_682 ();
 sg13g2_fill_2 FILLER_13_700 ();
 sg13g2_fill_1 FILLER_13_712 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_fill_1 FILLER_13_735 ();
 sg13g2_decap_4 FILLER_13_740 ();
 sg13g2_fill_1 FILLER_13_791 ();
 sg13g2_fill_2 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_4 FILLER_13_844 ();
 sg13g2_fill_1 FILLER_13_881 ();
 sg13g2_fill_2 FILLER_13_890 ();
 sg13g2_fill_1 FILLER_13_892 ();
 sg13g2_fill_1 FILLER_13_912 ();
 sg13g2_fill_1 FILLER_13_921 ();
 sg13g2_fill_2 FILLER_13_938 ();
 sg13g2_decap_4 FILLER_13_970 ();
 sg13g2_fill_2 FILLER_13_974 ();
 sg13g2_decap_8 FILLER_13_989 ();
 sg13g2_decap_4 FILLER_13_1000 ();
 sg13g2_fill_2 FILLER_13_1004 ();
 sg13g2_fill_2 FILLER_13_1032 ();
 sg13g2_fill_2 FILLER_13_1063 ();
 sg13g2_fill_1 FILLER_13_1065 ();
 sg13g2_decap_8 FILLER_13_1074 ();
 sg13g2_fill_1 FILLER_13_1088 ();
 sg13g2_decap_4 FILLER_13_1097 ();
 sg13g2_fill_1 FILLER_13_1124 ();
 sg13g2_decap_8 FILLER_13_1151 ();
 sg13g2_decap_4 FILLER_13_1158 ();
 sg13g2_fill_2 FILLER_13_1162 ();
 sg13g2_fill_2 FILLER_13_1168 ();
 sg13g2_fill_1 FILLER_13_1170 ();
 sg13g2_fill_2 FILLER_13_1179 ();
 sg13g2_fill_1 FILLER_13_1181 ();
 sg13g2_fill_2 FILLER_13_1186 ();
 sg13g2_fill_1 FILLER_13_1188 ();
 sg13g2_fill_2 FILLER_13_1212 ();
 sg13g2_fill_2 FILLER_13_1218 ();
 sg13g2_fill_1 FILLER_13_1220 ();
 sg13g2_fill_2 FILLER_13_1226 ();
 sg13g2_fill_1 FILLER_13_1228 ();
 sg13g2_decap_8 FILLER_13_1265 ();
 sg13g2_decap_4 FILLER_13_1272 ();
 sg13g2_fill_1 FILLER_13_1276 ();
 sg13g2_fill_1 FILLER_13_1321 ();
 sg13g2_fill_1 FILLER_13_1387 ();
 sg13g2_decap_4 FILLER_13_1392 ();
 sg13g2_fill_2 FILLER_13_1396 ();
 sg13g2_decap_8 FILLER_13_1403 ();
 sg13g2_fill_1 FILLER_13_1410 ();
 sg13g2_decap_4 FILLER_13_1421 ();
 sg13g2_fill_2 FILLER_13_1425 ();
 sg13g2_fill_2 FILLER_13_1440 ();
 sg13g2_decap_8 FILLER_13_1447 ();
 sg13g2_decap_8 FILLER_13_1454 ();
 sg13g2_fill_1 FILLER_13_1482 ();
 sg13g2_fill_1 FILLER_13_1495 ();
 sg13g2_fill_2 FILLER_13_1508 ();
 sg13g2_decap_8 FILLER_13_1585 ();
 sg13g2_fill_1 FILLER_13_1597 ();
 sg13g2_fill_2 FILLER_13_1603 ();
 sg13g2_fill_1 FILLER_13_1605 ();
 sg13g2_fill_1 FILLER_13_1614 ();
 sg13g2_fill_2 FILLER_13_1640 ();
 sg13g2_decap_4 FILLER_13_1656 ();
 sg13g2_decap_8 FILLER_13_1663 ();
 sg13g2_decap_4 FILLER_13_1670 ();
 sg13g2_decap_8 FILLER_13_1678 ();
 sg13g2_decap_4 FILLER_13_1685 ();
 sg13g2_fill_1 FILLER_13_1689 ();
 sg13g2_decap_8 FILLER_13_1694 ();
 sg13g2_decap_8 FILLER_13_1701 ();
 sg13g2_decap_8 FILLER_13_1708 ();
 sg13g2_decap_8 FILLER_13_1715 ();
 sg13g2_decap_8 FILLER_13_1722 ();
 sg13g2_decap_8 FILLER_13_1729 ();
 sg13g2_decap_8 FILLER_13_1736 ();
 sg13g2_decap_8 FILLER_13_1743 ();
 sg13g2_decap_8 FILLER_13_1750 ();
 sg13g2_decap_8 FILLER_13_1757 ();
 sg13g2_decap_8 FILLER_13_1764 ();
 sg13g2_fill_2 FILLER_13_1771 ();
 sg13g2_fill_1 FILLER_13_1773 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_22 ();
 sg13g2_fill_2 FILLER_14_55 ();
 sg13g2_decap_4 FILLER_14_61 ();
 sg13g2_fill_1 FILLER_14_65 ();
 sg13g2_fill_1 FILLER_14_90 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_fill_1 FILLER_14_165 ();
 sg13g2_fill_2 FILLER_14_180 ();
 sg13g2_fill_2 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_fill_1 FILLER_14_247 ();
 sg13g2_fill_2 FILLER_14_260 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_fill_1 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_fill_2 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_decap_4 FILLER_14_318 ();
 sg13g2_decap_4 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_360 ();
 sg13g2_fill_1 FILLER_14_366 ();
 sg13g2_fill_2 FILLER_14_398 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_decap_8 FILLER_14_418 ();
 sg13g2_decap_8 FILLER_14_425 ();
 sg13g2_decap_8 FILLER_14_432 ();
 sg13g2_fill_1 FILLER_14_439 ();
 sg13g2_decap_4 FILLER_14_445 ();
 sg13g2_fill_2 FILLER_14_449 ();
 sg13g2_fill_1 FILLER_14_459 ();
 sg13g2_decap_4 FILLER_14_474 ();
 sg13g2_fill_1 FILLER_14_478 ();
 sg13g2_decap_4 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_529 ();
 sg13g2_decap_8 FILLER_14_536 ();
 sg13g2_decap_4 FILLER_14_543 ();
 sg13g2_fill_1 FILLER_14_547 ();
 sg13g2_fill_2 FILLER_14_589 ();
 sg13g2_decap_4 FILLER_14_599 ();
 sg13g2_fill_2 FILLER_14_667 ();
 sg13g2_fill_2 FILLER_14_673 ();
 sg13g2_fill_1 FILLER_14_675 ();
 sg13g2_fill_2 FILLER_14_682 ();
 sg13g2_fill_1 FILLER_14_684 ();
 sg13g2_fill_2 FILLER_14_693 ();
 sg13g2_fill_1 FILLER_14_695 ();
 sg13g2_fill_1 FILLER_14_714 ();
 sg13g2_fill_2 FILLER_14_759 ();
 sg13g2_fill_1 FILLER_14_761 ();
 sg13g2_fill_1 FILLER_14_766 ();
 sg13g2_fill_2 FILLER_14_780 ();
 sg13g2_fill_2 FILLER_14_787 ();
 sg13g2_decap_4 FILLER_14_850 ();
 sg13g2_fill_1 FILLER_14_854 ();
 sg13g2_fill_2 FILLER_14_859 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_fill_2 FILLER_14_887 ();
 sg13g2_fill_1 FILLER_14_889 ();
 sg13g2_decap_8 FILLER_14_894 ();
 sg13g2_fill_2 FILLER_14_901 ();
 sg13g2_fill_1 FILLER_14_903 ();
 sg13g2_fill_2 FILLER_14_926 ();
 sg13g2_fill_1 FILLER_14_928 ();
 sg13g2_fill_2 FILLER_14_946 ();
 sg13g2_fill_1 FILLER_14_967 ();
 sg13g2_fill_2 FILLER_14_975 ();
 sg13g2_decap_4 FILLER_14_982 ();
 sg13g2_decap_4 FILLER_14_990 ();
 sg13g2_fill_1 FILLER_14_994 ();
 sg13g2_fill_2 FILLER_14_1000 ();
 sg13g2_decap_4 FILLER_14_1015 ();
 sg13g2_fill_1 FILLER_14_1019 ();
 sg13g2_decap_8 FILLER_14_1043 ();
 sg13g2_decap_8 FILLER_14_1050 ();
 sg13g2_fill_2 FILLER_14_1057 ();
 sg13g2_fill_1 FILLER_14_1059 ();
 sg13g2_fill_2 FILLER_14_1065 ();
 sg13g2_fill_1 FILLER_14_1073 ();
 sg13g2_fill_1 FILLER_14_1078 ();
 sg13g2_decap_4 FILLER_14_1105 ();
 sg13g2_decap_4 FILLER_14_1115 ();
 sg13g2_fill_2 FILLER_14_1124 ();
 sg13g2_fill_1 FILLER_14_1126 ();
 sg13g2_fill_1 FILLER_14_1136 ();
 sg13g2_decap_8 FILLER_14_1142 ();
 sg13g2_fill_2 FILLER_14_1149 ();
 sg13g2_fill_1 FILLER_14_1151 ();
 sg13g2_fill_2 FILLER_14_1182 ();
 sg13g2_fill_1 FILLER_14_1184 ();
 sg13g2_fill_2 FILLER_14_1207 ();
 sg13g2_decap_8 FILLER_14_1235 ();
 sg13g2_decap_8 FILLER_14_1242 ();
 sg13g2_fill_1 FILLER_14_1254 ();
 sg13g2_fill_2 FILLER_14_1269 ();
 sg13g2_fill_1 FILLER_14_1271 ();
 sg13g2_decap_8 FILLER_14_1343 ();
 sg13g2_fill_2 FILLER_14_1350 ();
 sg13g2_fill_2 FILLER_14_1355 ();
 sg13g2_fill_2 FILLER_14_1364 ();
 sg13g2_fill_2 FILLER_14_1383 ();
 sg13g2_fill_1 FILLER_14_1385 ();
 sg13g2_fill_1 FILLER_14_1391 ();
 sg13g2_fill_1 FILLER_14_1397 ();
 sg13g2_decap_4 FILLER_14_1402 ();
 sg13g2_fill_2 FILLER_14_1406 ();
 sg13g2_decap_4 FILLER_14_1413 ();
 sg13g2_fill_1 FILLER_14_1417 ();
 sg13g2_decap_8 FILLER_14_1422 ();
 sg13g2_fill_2 FILLER_14_1429 ();
 sg13g2_decap_8 FILLER_14_1448 ();
 sg13g2_fill_1 FILLER_14_1455 ();
 sg13g2_fill_2 FILLER_14_1516 ();
 sg13g2_fill_2 FILLER_14_1566 ();
 sg13g2_fill_2 FILLER_14_1584 ();
 sg13g2_fill_1 FILLER_14_1586 ();
 sg13g2_decap_4 FILLER_14_1618 ();
 sg13g2_fill_1 FILLER_14_1622 ();
 sg13g2_fill_1 FILLER_14_1634 ();
 sg13g2_fill_1 FILLER_14_1686 ();
 sg13g2_decap_8 FILLER_14_1692 ();
 sg13g2_decap_8 FILLER_14_1699 ();
 sg13g2_decap_8 FILLER_14_1706 ();
 sg13g2_decap_8 FILLER_14_1713 ();
 sg13g2_decap_8 FILLER_14_1720 ();
 sg13g2_decap_8 FILLER_14_1727 ();
 sg13g2_decap_8 FILLER_14_1734 ();
 sg13g2_decap_8 FILLER_14_1741 ();
 sg13g2_decap_8 FILLER_14_1748 ();
 sg13g2_decap_8 FILLER_14_1755 ();
 sg13g2_decap_8 FILLER_14_1762 ();
 sg13g2_decap_4 FILLER_14_1769 ();
 sg13g2_fill_1 FILLER_14_1773 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_4 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_fill_2 FILLER_15_60 ();
 sg13g2_fill_1 FILLER_15_89 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_fill_2 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_154 ();
 sg13g2_fill_1 FILLER_15_165 ();
 sg13g2_fill_1 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_2 FILLER_15_209 ();
 sg13g2_fill_2 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_271 ();
 sg13g2_decap_4 FILLER_15_293 ();
 sg13g2_fill_2 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_320 ();
 sg13g2_fill_2 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_361 ();
 sg13g2_fill_1 FILLER_15_385 ();
 sg13g2_fill_1 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_414 ();
 sg13g2_fill_1 FILLER_15_421 ();
 sg13g2_decap_4 FILLER_15_479 ();
 sg13g2_fill_2 FILLER_15_483 ();
 sg13g2_decap_4 FILLER_15_489 ();
 sg13g2_fill_1 FILLER_15_507 ();
 sg13g2_decap_4 FILLER_15_512 ();
 sg13g2_fill_2 FILLER_15_516 ();
 sg13g2_fill_2 FILLER_15_521 ();
 sg13g2_fill_1 FILLER_15_523 ();
 sg13g2_fill_1 FILLER_15_537 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_fill_2 FILLER_15_550 ();
 sg13g2_fill_1 FILLER_15_552 ();
 sg13g2_fill_2 FILLER_15_573 ();
 sg13g2_fill_1 FILLER_15_575 ();
 sg13g2_fill_2 FILLER_15_580 ();
 sg13g2_fill_1 FILLER_15_582 ();
 sg13g2_fill_2 FILLER_15_597 ();
 sg13g2_fill_2 FILLER_15_635 ();
 sg13g2_fill_1 FILLER_15_660 ();
 sg13g2_decap_8 FILLER_15_666 ();
 sg13g2_fill_2 FILLER_15_673 ();
 sg13g2_fill_1 FILLER_15_683 ();
 sg13g2_decap_4 FILLER_15_689 ();
 sg13g2_decap_8 FILLER_15_706 ();
 sg13g2_fill_2 FILLER_15_713 ();
 sg13g2_decap_8 FILLER_15_723 ();
 sg13g2_fill_2 FILLER_15_730 ();
 sg13g2_fill_1 FILLER_15_732 ();
 sg13g2_decap_8 FILLER_15_737 ();
 sg13g2_fill_2 FILLER_15_744 ();
 sg13g2_fill_2 FILLER_15_771 ();
 sg13g2_fill_1 FILLER_15_801 ();
 sg13g2_fill_2 FILLER_15_819 ();
 sg13g2_fill_1 FILLER_15_821 ();
 sg13g2_fill_2 FILLER_15_831 ();
 sg13g2_decap_8 FILLER_15_837 ();
 sg13g2_decap_8 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_851 ();
 sg13g2_fill_2 FILLER_15_858 ();
 sg13g2_decap_8 FILLER_15_865 ();
 sg13g2_decap_8 FILLER_15_872 ();
 sg13g2_fill_2 FILLER_15_879 ();
 sg13g2_fill_1 FILLER_15_881 ();
 sg13g2_decap_8 FILLER_15_890 ();
 sg13g2_fill_1 FILLER_15_897 ();
 sg13g2_decap_4 FILLER_15_902 ();
 sg13g2_fill_1 FILLER_15_906 ();
 sg13g2_fill_1 FILLER_15_929 ();
 sg13g2_decap_4 FILLER_15_934 ();
 sg13g2_decap_8 FILLER_15_944 ();
 sg13g2_fill_2 FILLER_15_951 ();
 sg13g2_fill_1 FILLER_15_953 ();
 sg13g2_decap_8 FILLER_15_998 ();
 sg13g2_fill_1 FILLER_15_1005 ();
 sg13g2_decap_4 FILLER_15_1011 ();
 sg13g2_fill_1 FILLER_15_1015 ();
 sg13g2_fill_2 FILLER_15_1027 ();
 sg13g2_fill_1 FILLER_15_1029 ();
 sg13g2_fill_1 FILLER_15_1048 ();
 sg13g2_fill_2 FILLER_15_1065 ();
 sg13g2_fill_2 FILLER_15_1075 ();
 sg13g2_fill_1 FILLER_15_1077 ();
 sg13g2_fill_1 FILLER_15_1101 ();
 sg13g2_fill_2 FILLER_15_1110 ();
 sg13g2_fill_1 FILLER_15_1112 ();
 sg13g2_fill_2 FILLER_15_1121 ();
 sg13g2_decap_8 FILLER_15_1158 ();
 sg13g2_decap_4 FILLER_15_1181 ();
 sg13g2_fill_1 FILLER_15_1185 ();
 sg13g2_decap_8 FILLER_15_1190 ();
 sg13g2_decap_4 FILLER_15_1197 ();
 sg13g2_fill_1 FILLER_15_1201 ();
 sg13g2_decap_8 FILLER_15_1215 ();
 sg13g2_fill_2 FILLER_15_1227 ();
 sg13g2_fill_1 FILLER_15_1229 ();
 sg13g2_fill_1 FILLER_15_1241 ();
 sg13g2_fill_1 FILLER_15_1253 ();
 sg13g2_fill_2 FILLER_15_1259 ();
 sg13g2_fill_1 FILLER_15_1270 ();
 sg13g2_fill_1 FILLER_15_1275 ();
 sg13g2_fill_2 FILLER_15_1280 ();
 sg13g2_decap_4 FILLER_15_1291 ();
 sg13g2_fill_1 FILLER_15_1295 ();
 sg13g2_decap_4 FILLER_15_1300 ();
 sg13g2_fill_1 FILLER_15_1309 ();
 sg13g2_decap_4 FILLER_15_1328 ();
 sg13g2_decap_8 FILLER_15_1335 ();
 sg13g2_fill_2 FILLER_15_1354 ();
 sg13g2_fill_1 FILLER_15_1356 ();
 sg13g2_fill_1 FILLER_15_1399 ();
 sg13g2_decap_8 FILLER_15_1405 ();
 sg13g2_decap_8 FILLER_15_1416 ();
 sg13g2_decap_4 FILLER_15_1423 ();
 sg13g2_fill_2 FILLER_15_1427 ();
 sg13g2_fill_2 FILLER_15_1437 ();
 sg13g2_fill_2 FILLER_15_1443 ();
 sg13g2_fill_2 FILLER_15_1454 ();
 sg13g2_fill_1 FILLER_15_1456 ();
 sg13g2_fill_2 FILLER_15_1472 ();
 sg13g2_fill_1 FILLER_15_1474 ();
 sg13g2_fill_1 FILLER_15_1479 ();
 sg13g2_fill_1 FILLER_15_1499 ();
 sg13g2_fill_1 FILLER_15_1536 ();
 sg13g2_fill_1 FILLER_15_1545 ();
 sg13g2_fill_1 FILLER_15_1553 ();
 sg13g2_fill_1 FILLER_15_1570 ();
 sg13g2_fill_2 FILLER_15_1587 ();
 sg13g2_fill_2 FILLER_15_1613 ();
 sg13g2_decap_4 FILLER_15_1625 ();
 sg13g2_fill_1 FILLER_15_1629 ();
 sg13g2_fill_2 FILLER_15_1644 ();
 sg13g2_fill_2 FILLER_15_1650 ();
 sg13g2_fill_1 FILLER_15_1652 ();
 sg13g2_decap_4 FILLER_15_1658 ();
 sg13g2_fill_1 FILLER_15_1662 ();
 sg13g2_fill_2 FILLER_15_1677 ();
 sg13g2_fill_1 FILLER_15_1679 ();
 sg13g2_fill_1 FILLER_15_1697 ();
 sg13g2_decap_4 FILLER_15_1703 ();
 sg13g2_decap_8 FILLER_15_1716 ();
 sg13g2_decap_8 FILLER_15_1723 ();
 sg13g2_decap_8 FILLER_15_1730 ();
 sg13g2_decap_8 FILLER_15_1737 ();
 sg13g2_decap_8 FILLER_15_1744 ();
 sg13g2_decap_8 FILLER_15_1751 ();
 sg13g2_decap_8 FILLER_15_1758 ();
 sg13g2_decap_8 FILLER_15_1765 ();
 sg13g2_fill_2 FILLER_15_1772 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_fill_2 FILLER_16_18 ();
 sg13g2_decap_8 FILLER_16_24 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_64 ();
 sg13g2_fill_1 FILLER_16_66 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_fill_1 FILLER_16_85 ();
 sg13g2_fill_1 FILLER_16_106 ();
 sg13g2_fill_1 FILLER_16_118 ();
 sg13g2_fill_2 FILLER_16_190 ();
 sg13g2_fill_1 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_decap_4 FILLER_16_263 ();
 sg13g2_fill_1 FILLER_16_267 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_292 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_decap_4 FILLER_16_329 ();
 sg13g2_fill_1 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_fill_2 FILLER_16_366 ();
 sg13g2_decap_4 FILLER_16_424 ();
 sg13g2_fill_1 FILLER_16_428 ();
 sg13g2_decap_4 FILLER_16_445 ();
 sg13g2_fill_1 FILLER_16_465 ();
 sg13g2_fill_1 FILLER_16_475 ();
 sg13g2_fill_1 FILLER_16_484 ();
 sg13g2_fill_1 FILLER_16_490 ();
 sg13g2_fill_1 FILLER_16_499 ();
 sg13g2_fill_2 FILLER_16_505 ();
 sg13g2_fill_1 FILLER_16_507 ();
 sg13g2_fill_2 FILLER_16_512 ();
 sg13g2_fill_2 FILLER_16_533 ();
 sg13g2_fill_1 FILLER_16_568 ();
 sg13g2_decap_8 FILLER_16_575 ();
 sg13g2_fill_2 FILLER_16_598 ();
 sg13g2_fill_1 FILLER_16_600 ();
 sg13g2_fill_2 FILLER_16_614 ();
 sg13g2_fill_2 FILLER_16_638 ();
 sg13g2_decap_8 FILLER_16_670 ();
 sg13g2_fill_2 FILLER_16_698 ();
 sg13g2_decap_4 FILLER_16_708 ();
 sg13g2_decap_8 FILLER_16_720 ();
 sg13g2_fill_2 FILLER_16_727 ();
 sg13g2_fill_1 FILLER_16_729 ();
 sg13g2_decap_8 FILLER_16_740 ();
 sg13g2_decap_8 FILLER_16_747 ();
 sg13g2_fill_1 FILLER_16_754 ();
 sg13g2_decap_4 FILLER_16_759 ();
 sg13g2_fill_1 FILLER_16_763 ();
 sg13g2_fill_1 FILLER_16_785 ();
 sg13g2_fill_2 FILLER_16_798 ();
 sg13g2_fill_1 FILLER_16_808 ();
 sg13g2_fill_2 FILLER_16_822 ();
 sg13g2_fill_1 FILLER_16_824 ();
 sg13g2_fill_1 FILLER_16_830 ();
 sg13g2_decap_8 FILLER_16_839 ();
 sg13g2_fill_2 FILLER_16_846 ();
 sg13g2_decap_8 FILLER_16_864 ();
 sg13g2_decap_4 FILLER_16_871 ();
 sg13g2_decap_8 FILLER_16_883 ();
 sg13g2_decap_8 FILLER_16_890 ();
 sg13g2_decap_4 FILLER_16_897 ();
 sg13g2_fill_2 FILLER_16_906 ();
 sg13g2_decap_8 FILLER_16_921 ();
 sg13g2_fill_2 FILLER_16_947 ();
 sg13g2_fill_1 FILLER_16_949 ();
 sg13g2_decap_8 FILLER_16_958 ();
 sg13g2_decap_8 FILLER_16_965 ();
 sg13g2_decap_8 FILLER_16_972 ();
 sg13g2_decap_8 FILLER_16_979 ();
 sg13g2_fill_1 FILLER_16_986 ();
 sg13g2_decap_8 FILLER_16_1022 ();
 sg13g2_fill_2 FILLER_16_1029 ();
 sg13g2_fill_1 FILLER_16_1031 ();
 sg13g2_decap_8 FILLER_16_1038 ();
 sg13g2_decap_8 FILLER_16_1045 ();
 sg13g2_fill_2 FILLER_16_1066 ();
 sg13g2_fill_1 FILLER_16_1068 ();
 sg13g2_fill_2 FILLER_16_1088 ();
 sg13g2_fill_1 FILLER_16_1090 ();
 sg13g2_decap_4 FILLER_16_1105 ();
 sg13g2_fill_1 FILLER_16_1109 ();
 sg13g2_fill_1 FILLER_16_1115 ();
 sg13g2_decap_4 FILLER_16_1136 ();
 sg13g2_fill_1 FILLER_16_1140 ();
 sg13g2_fill_1 FILLER_16_1153 ();
 sg13g2_decap_4 FILLER_16_1185 ();
 sg13g2_decap_4 FILLER_16_1193 ();
 sg13g2_fill_1 FILLER_16_1197 ();
 sg13g2_decap_4 FILLER_16_1203 ();
 sg13g2_fill_1 FILLER_16_1207 ();
 sg13g2_decap_8 FILLER_16_1212 ();
 sg13g2_decap_8 FILLER_16_1219 ();
 sg13g2_fill_1 FILLER_16_1226 ();
 sg13g2_fill_1 FILLER_16_1248 ();
 sg13g2_fill_2 FILLER_16_1253 ();
 sg13g2_fill_1 FILLER_16_1259 ();
 sg13g2_decap_4 FILLER_16_1296 ();
 sg13g2_decap_4 FILLER_16_1307 ();
 sg13g2_fill_2 FILLER_16_1320 ();
 sg13g2_fill_1 FILLER_16_1322 ();
 sg13g2_fill_1 FILLER_16_1327 ();
 sg13g2_fill_1 FILLER_16_1349 ();
 sg13g2_decap_8 FILLER_16_1364 ();
 sg13g2_fill_2 FILLER_16_1371 ();
 sg13g2_fill_1 FILLER_16_1373 ();
 sg13g2_decap_8 FILLER_16_1378 ();
 sg13g2_fill_2 FILLER_16_1385 ();
 sg13g2_fill_2 FILLER_16_1419 ();
 sg13g2_fill_1 FILLER_16_1425 ();
 sg13g2_fill_1 FILLER_16_1468 ();
 sg13g2_fill_2 FILLER_16_1474 ();
 sg13g2_fill_1 FILLER_16_1482 ();
 sg13g2_fill_1 FILLER_16_1488 ();
 sg13g2_fill_2 FILLER_16_1494 ();
 sg13g2_fill_1 FILLER_16_1500 ();
 sg13g2_fill_2 FILLER_16_1510 ();
 sg13g2_fill_1 FILLER_16_1532 ();
 sg13g2_fill_2 FILLER_16_1542 ();
 sg13g2_decap_4 FILLER_16_1584 ();
 sg13g2_decap_8 FILLER_16_1594 ();
 sg13g2_decap_4 FILLER_16_1601 ();
 sg13g2_fill_1 FILLER_16_1609 ();
 sg13g2_fill_2 FILLER_16_1615 ();
 sg13g2_fill_1 FILLER_16_1617 ();
 sg13g2_decap_8 FILLER_16_1627 ();
 sg13g2_fill_1 FILLER_16_1634 ();
 sg13g2_decap_4 FILLER_16_1647 ();
 sg13g2_decap_4 FILLER_16_1668 ();
 sg13g2_fill_2 FILLER_16_1672 ();
 sg13g2_fill_1 FILLER_16_1678 ();
 sg13g2_fill_2 FILLER_16_1692 ();
 sg13g2_fill_1 FILLER_16_1701 ();
 sg13g2_decap_8 FILLER_16_1707 ();
 sg13g2_decap_8 FILLER_16_1714 ();
 sg13g2_decap_8 FILLER_16_1721 ();
 sg13g2_decap_8 FILLER_16_1728 ();
 sg13g2_decap_8 FILLER_16_1735 ();
 sg13g2_decap_8 FILLER_16_1742 ();
 sg13g2_decap_8 FILLER_16_1749 ();
 sg13g2_decap_8 FILLER_16_1756 ();
 sg13g2_decap_8 FILLER_16_1763 ();
 sg13g2_decap_4 FILLER_16_1770 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_decap_4 FILLER_17_86 ();
 sg13g2_fill_2 FILLER_17_93 ();
 sg13g2_fill_1 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_139 ();
 sg13g2_fill_2 FILLER_17_146 ();
 sg13g2_fill_2 FILLER_17_165 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_197 ();
 sg13g2_decap_4 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_261 ();
 sg13g2_decap_4 FILLER_17_270 ();
 sg13g2_fill_2 FILLER_17_274 ();
 sg13g2_fill_2 FILLER_17_287 ();
 sg13g2_fill_1 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_fill_1 FILLER_17_387 ();
 sg13g2_fill_1 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_decap_4 FILLER_17_441 ();
 sg13g2_fill_2 FILLER_17_445 ();
 sg13g2_decap_8 FILLER_17_470 ();
 sg13g2_fill_1 FILLER_17_498 ();
 sg13g2_decap_4 FILLER_17_504 ();
 sg13g2_fill_2 FILLER_17_536 ();
 sg13g2_decap_4 FILLER_17_547 ();
 sg13g2_fill_1 FILLER_17_556 ();
 sg13g2_fill_2 FILLER_17_570 ();
 sg13g2_decap_8 FILLER_17_576 ();
 sg13g2_fill_1 FILLER_17_583 ();
 sg13g2_decap_4 FILLER_17_604 ();
 sg13g2_fill_1 FILLER_17_608 ();
 sg13g2_fill_1 FILLER_17_617 ();
 sg13g2_fill_1 FILLER_17_628 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_fill_1 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_670 ();
 sg13g2_fill_1 FILLER_17_677 ();
 sg13g2_fill_2 FILLER_17_681 ();
 sg13g2_fill_1 FILLER_17_683 ();
 sg13g2_decap_8 FILLER_17_698 ();
 sg13g2_decap_4 FILLER_17_716 ();
 sg13g2_fill_1 FILLER_17_720 ();
 sg13g2_decap_8 FILLER_17_729 ();
 sg13g2_fill_1 FILLER_17_736 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_4 FILLER_17_749 ();
 sg13g2_fill_2 FILLER_17_753 ();
 sg13g2_fill_2 FILLER_17_759 ();
 sg13g2_fill_1 FILLER_17_761 ();
 sg13g2_fill_1 FILLER_17_767 ();
 sg13g2_fill_1 FILLER_17_781 ();
 sg13g2_fill_2 FILLER_17_787 ();
 sg13g2_fill_1 FILLER_17_797 ();
 sg13g2_fill_1 FILLER_17_804 ();
 sg13g2_fill_2 FILLER_17_810 ();
 sg13g2_fill_1 FILLER_17_818 ();
 sg13g2_fill_2 FILLER_17_827 ();
 sg13g2_decap_4 FILLER_17_843 ();
 sg13g2_decap_4 FILLER_17_866 ();
 sg13g2_fill_2 FILLER_17_870 ();
 sg13g2_decap_8 FILLER_17_880 ();
 sg13g2_decap_8 FILLER_17_887 ();
 sg13g2_decap_8 FILLER_17_894 ();
 sg13g2_fill_2 FILLER_17_905 ();
 sg13g2_fill_2 FILLER_17_912 ();
 sg13g2_fill_1 FILLER_17_914 ();
 sg13g2_fill_2 FILLER_17_940 ();
 sg13g2_fill_1 FILLER_17_942 ();
 sg13g2_decap_8 FILLER_17_948 ();
 sg13g2_fill_2 FILLER_17_955 ();
 sg13g2_fill_2 FILLER_17_962 ();
 sg13g2_fill_1 FILLER_17_968 ();
 sg13g2_fill_1 FILLER_17_987 ();
 sg13g2_fill_1 FILLER_17_992 ();
 sg13g2_fill_1 FILLER_17_999 ();
 sg13g2_fill_2 FILLER_17_1010 ();
 sg13g2_fill_1 FILLER_17_1012 ();
 sg13g2_fill_1 FILLER_17_1022 ();
 sg13g2_fill_1 FILLER_17_1027 ();
 sg13g2_decap_8 FILLER_17_1032 ();
 sg13g2_decap_8 FILLER_17_1039 ();
 sg13g2_fill_2 FILLER_17_1046 ();
 sg13g2_fill_1 FILLER_17_1048 ();
 sg13g2_decap_8 FILLER_17_1106 ();
 sg13g2_decap_8 FILLER_17_1113 ();
 sg13g2_fill_1 FILLER_17_1120 ();
 sg13g2_fill_2 FILLER_17_1129 ();
 sg13g2_fill_1 FILLER_17_1131 ();
 sg13g2_fill_1 FILLER_17_1140 ();
 sg13g2_fill_1 FILLER_17_1146 ();
 sg13g2_fill_1 FILLER_17_1160 ();
 sg13g2_fill_2 FILLER_17_1192 ();
 sg13g2_fill_1 FILLER_17_1194 ();
 sg13g2_decap_8 FILLER_17_1207 ();
 sg13g2_decap_8 FILLER_17_1214 ();
 sg13g2_decap_8 FILLER_17_1221 ();
 sg13g2_fill_2 FILLER_17_1228 ();
 sg13g2_fill_2 FILLER_17_1261 ();
 sg13g2_decap_4 FILLER_17_1272 ();
 sg13g2_fill_2 FILLER_17_1276 ();
 sg13g2_decap_4 FILLER_17_1286 ();
 sg13g2_decap_8 FILLER_17_1318 ();
 sg13g2_fill_2 FILLER_17_1325 ();
 sg13g2_fill_1 FILLER_17_1327 ();
 sg13g2_decap_8 FILLER_17_1336 ();
 sg13g2_decap_4 FILLER_17_1381 ();
 sg13g2_fill_1 FILLER_17_1385 ();
 sg13g2_fill_2 FILLER_17_1391 ();
 sg13g2_decap_8 FILLER_17_1397 ();
 sg13g2_fill_1 FILLER_17_1404 ();
 sg13g2_fill_1 FILLER_17_1421 ();
 sg13g2_fill_2 FILLER_17_1447 ();
 sg13g2_decap_4 FILLER_17_1465 ();
 sg13g2_fill_2 FILLER_17_1474 ();
 sg13g2_fill_2 FILLER_17_1499 ();
 sg13g2_fill_1 FILLER_17_1516 ();
 sg13g2_fill_1 FILLER_17_1520 ();
 sg13g2_fill_2 FILLER_17_1563 ();
 sg13g2_decap_8 FILLER_17_1575 ();
 sg13g2_fill_1 FILLER_17_1582 ();
 sg13g2_fill_1 FILLER_17_1591 ();
 sg13g2_fill_1 FILLER_17_1596 ();
 sg13g2_decap_8 FILLER_17_1610 ();
 sg13g2_decap_8 FILLER_17_1617 ();
 sg13g2_fill_2 FILLER_17_1624 ();
 sg13g2_fill_1 FILLER_17_1651 ();
 sg13g2_fill_1 FILLER_17_1667 ();
 sg13g2_fill_1 FILLER_17_1673 ();
 sg13g2_decap_4 FILLER_17_1689 ();
 sg13g2_fill_2 FILLER_17_1698 ();
 sg13g2_decap_8 FILLER_17_1710 ();
 sg13g2_decap_8 FILLER_17_1717 ();
 sg13g2_decap_8 FILLER_17_1724 ();
 sg13g2_decap_8 FILLER_17_1731 ();
 sg13g2_decap_8 FILLER_17_1738 ();
 sg13g2_decap_8 FILLER_17_1745 ();
 sg13g2_decap_8 FILLER_17_1752 ();
 sg13g2_decap_8 FILLER_17_1759 ();
 sg13g2_decap_8 FILLER_17_1766 ();
 sg13g2_fill_1 FILLER_17_1773 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_27 ();
 sg13g2_fill_2 FILLER_18_41 ();
 sg13g2_fill_1 FILLER_18_54 ();
 sg13g2_fill_1 FILLER_18_69 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_4 FILLER_18_91 ();
 sg13g2_fill_2 FILLER_18_95 ();
 sg13g2_fill_1 FILLER_18_111 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_2 FILLER_18_212 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_decap_4 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_272 ();
 sg13g2_fill_2 FILLER_18_278 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_fill_2 FILLER_18_302 ();
 sg13g2_decap_4 FILLER_18_312 ();
 sg13g2_fill_2 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_322 ();
 sg13g2_decap_4 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_340 ();
 sg13g2_decap_4 FILLER_18_346 ();
 sg13g2_fill_1 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_367 ();
 sg13g2_fill_1 FILLER_18_369 ();
 sg13g2_fill_1 FILLER_18_386 ();
 sg13g2_fill_2 FILLER_18_397 ();
 sg13g2_fill_2 FILLER_18_414 ();
 sg13g2_fill_1 FILLER_18_416 ();
 sg13g2_fill_2 FILLER_18_421 ();
 sg13g2_decap_8 FILLER_18_431 ();
 sg13g2_decap_8 FILLER_18_438 ();
 sg13g2_decap_8 FILLER_18_445 ();
 sg13g2_decap_8 FILLER_18_452 ();
 sg13g2_decap_4 FILLER_18_459 ();
 sg13g2_fill_2 FILLER_18_463 ();
 sg13g2_decap_8 FILLER_18_468 ();
 sg13g2_fill_2 FILLER_18_475 ();
 sg13g2_fill_1 FILLER_18_477 ();
 sg13g2_decap_8 FILLER_18_486 ();
 sg13g2_decap_8 FILLER_18_493 ();
 sg13g2_decap_4 FILLER_18_500 ();
 sg13g2_fill_2 FILLER_18_512 ();
 sg13g2_fill_2 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_545 ();
 sg13g2_decap_4 FILLER_18_552 ();
 sg13g2_fill_1 FILLER_18_556 ();
 sg13g2_decap_8 FILLER_18_566 ();
 sg13g2_decap_8 FILLER_18_573 ();
 sg13g2_decap_4 FILLER_18_580 ();
 sg13g2_decap_4 FILLER_18_588 ();
 sg13g2_decap_4 FILLER_18_603 ();
 sg13g2_decap_8 FILLER_18_610 ();
 sg13g2_fill_2 FILLER_18_642 ();
 sg13g2_decap_8 FILLER_18_648 ();
 sg13g2_decap_8 FILLER_18_660 ();
 sg13g2_decap_8 FILLER_18_667 ();
 sg13g2_fill_2 FILLER_18_674 ();
 sg13g2_fill_1 FILLER_18_676 ();
 sg13g2_decap_4 FILLER_18_688 ();
 sg13g2_fill_2 FILLER_18_700 ();
 sg13g2_decap_4 FILLER_18_709 ();
 sg13g2_fill_2 FILLER_18_713 ();
 sg13g2_decap_8 FILLER_18_732 ();
 sg13g2_decap_8 FILLER_18_739 ();
 sg13g2_decap_4 FILLER_18_746 ();
 sg13g2_fill_1 FILLER_18_757 ();
 sg13g2_fill_2 FILLER_18_785 ();
 sg13g2_fill_1 FILLER_18_787 ();
 sg13g2_fill_1 FILLER_18_795 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_4 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_decap_4 FILLER_18_861 ();
 sg13g2_fill_2 FILLER_18_865 ();
 sg13g2_decap_4 FILLER_18_895 ();
 sg13g2_decap_8 FILLER_18_915 ();
 sg13g2_decap_8 FILLER_18_922 ();
 sg13g2_fill_1 FILLER_18_929 ();
 sg13g2_decap_8 FILLER_18_950 ();
 sg13g2_fill_1 FILLER_18_961 ();
 sg13g2_decap_4 FILLER_18_967 ();
 sg13g2_fill_1 FILLER_18_971 ();
 sg13g2_fill_1 FILLER_18_985 ();
 sg13g2_fill_1 FILLER_18_991 ();
 sg13g2_fill_1 FILLER_18_1008 ();
 sg13g2_decap_8 FILLER_18_1029 ();
 sg13g2_decap_8 FILLER_18_1036 ();
 sg13g2_decap_8 FILLER_18_1043 ();
 sg13g2_decap_4 FILLER_18_1050 ();
 sg13g2_fill_2 FILLER_18_1065 ();
 sg13g2_fill_1 FILLER_18_1081 ();
 sg13g2_decap_8 FILLER_18_1087 ();
 sg13g2_decap_8 FILLER_18_1094 ();
 sg13g2_fill_2 FILLER_18_1101 ();
 sg13g2_fill_1 FILLER_18_1103 ();
 sg13g2_fill_1 FILLER_18_1125 ();
 sg13g2_fill_1 FILLER_18_1130 ();
 sg13g2_fill_1 FILLER_18_1135 ();
 sg13g2_decap_8 FILLER_18_1140 ();
 sg13g2_decap_4 FILLER_18_1147 ();
 sg13g2_fill_1 FILLER_18_1151 ();
 sg13g2_fill_1 FILLER_18_1208 ();
 sg13g2_decap_8 FILLER_18_1214 ();
 sg13g2_decap_4 FILLER_18_1221 ();
 sg13g2_fill_2 FILLER_18_1229 ();
 sg13g2_fill_2 FILLER_18_1239 ();
 sg13g2_decap_4 FILLER_18_1249 ();
 sg13g2_fill_2 FILLER_18_1253 ();
 sg13g2_fill_2 FILLER_18_1273 ();
 sg13g2_decap_4 FILLER_18_1283 ();
 sg13g2_fill_1 FILLER_18_1294 ();
 sg13g2_decap_8 FILLER_18_1327 ();
 sg13g2_decap_4 FILLER_18_1334 ();
 sg13g2_fill_1 FILLER_18_1338 ();
 sg13g2_decap_8 FILLER_18_1372 ();
 sg13g2_decap_4 FILLER_18_1379 ();
 sg13g2_fill_2 FILLER_18_1383 ();
 sg13g2_decap_8 FILLER_18_1389 ();
 sg13g2_decap_8 FILLER_18_1396 ();
 sg13g2_decap_4 FILLER_18_1403 ();
 sg13g2_fill_1 FILLER_18_1407 ();
 sg13g2_decap_4 FILLER_18_1416 ();
 sg13g2_fill_1 FILLER_18_1420 ();
 sg13g2_fill_2 FILLER_18_1429 ();
 sg13g2_fill_1 FILLER_18_1437 ();
 sg13g2_decap_4 FILLER_18_1469 ();
 sg13g2_fill_2 FILLER_18_1473 ();
 sg13g2_decap_4 FILLER_18_1480 ();
 sg13g2_fill_1 FILLER_18_1520 ();
 sg13g2_fill_2 FILLER_18_1536 ();
 sg13g2_decap_8 FILLER_18_1567 ();
 sg13g2_fill_1 FILLER_18_1582 ();
 sg13g2_decap_8 FILLER_18_1608 ();
 sg13g2_decap_8 FILLER_18_1615 ();
 sg13g2_fill_1 FILLER_18_1635 ();
 sg13g2_fill_2 FILLER_18_1640 ();
 sg13g2_fill_1 FILLER_18_1642 ();
 sg13g2_decap_8 FILLER_18_1648 ();
 sg13g2_decap_4 FILLER_18_1655 ();
 sg13g2_fill_1 FILLER_18_1659 ();
 sg13g2_fill_1 FILLER_18_1665 ();
 sg13g2_fill_2 FILLER_18_1671 ();
 sg13g2_fill_1 FILLER_18_1678 ();
 sg13g2_fill_1 FILLER_18_1699 ();
 sg13g2_fill_1 FILLER_18_1704 ();
 sg13g2_decap_8 FILLER_18_1724 ();
 sg13g2_decap_8 FILLER_18_1731 ();
 sg13g2_decap_8 FILLER_18_1738 ();
 sg13g2_decap_8 FILLER_18_1745 ();
 sg13g2_decap_8 FILLER_18_1752 ();
 sg13g2_decap_8 FILLER_18_1759 ();
 sg13g2_decap_8 FILLER_18_1766 ();
 sg13g2_fill_1 FILLER_18_1773 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_11 ();
 sg13g2_fill_2 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_24 ();
 sg13g2_decap_4 FILLER_19_31 ();
 sg13g2_decap_4 FILLER_19_73 ();
 sg13g2_decap_4 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_89 ();
 sg13g2_decap_4 FILLER_19_94 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_124 ();
 sg13g2_fill_2 FILLER_19_183 ();
 sg13g2_fill_1 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_215 ();
 sg13g2_decap_4 FILLER_19_222 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_fill_2 FILLER_19_235 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_361 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_decap_4 FILLER_19_392 ();
 sg13g2_fill_2 FILLER_19_409 ();
 sg13g2_fill_1 FILLER_19_419 ();
 sg13g2_fill_1 FILLER_19_428 ();
 sg13g2_fill_1 FILLER_19_437 ();
 sg13g2_fill_2 FILLER_19_459 ();
 sg13g2_decap_4 FILLER_19_465 ();
 sg13g2_fill_1 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_474 ();
 sg13g2_decap_8 FILLER_19_481 ();
 sg13g2_decap_8 FILLER_19_488 ();
 sg13g2_fill_1 FILLER_19_495 ();
 sg13g2_fill_1 FILLER_19_501 ();
 sg13g2_fill_2 FILLER_19_523 ();
 sg13g2_decap_4 FILLER_19_559 ();
 sg13g2_fill_2 FILLER_19_563 ();
 sg13g2_decap_8 FILLER_19_573 ();
 sg13g2_fill_1 FILLER_19_580 ();
 sg13g2_decap_8 FILLER_19_612 ();
 sg13g2_decap_8 FILLER_19_619 ();
 sg13g2_fill_2 FILLER_19_626 ();
 sg13g2_fill_2 FILLER_19_636 ();
 sg13g2_fill_1 FILLER_19_638 ();
 sg13g2_decap_8 FILLER_19_704 ();
 sg13g2_fill_2 FILLER_19_711 ();
 sg13g2_decap_8 FILLER_19_718 ();
 sg13g2_decap_4 FILLER_19_725 ();
 sg13g2_fill_2 FILLER_19_729 ();
 sg13g2_decap_4 FILLER_19_735 ();
 sg13g2_fill_2 FILLER_19_765 ();
 sg13g2_fill_1 FILLER_19_775 ();
 sg13g2_fill_2 FILLER_19_794 ();
 sg13g2_decap_8 FILLER_19_817 ();
 sg13g2_decap_4 FILLER_19_824 ();
 sg13g2_fill_1 FILLER_19_828 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_fill_2 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_870 ();
 sg13g2_decap_8 FILLER_19_877 ();
 sg13g2_fill_1 FILLER_19_884 ();
 sg13g2_decap_8 FILLER_19_919 ();
 sg13g2_decap_8 FILLER_19_926 ();
 sg13g2_fill_1 FILLER_19_933 ();
 sg13g2_decap_8 FILLER_19_950 ();
 sg13g2_decap_8 FILLER_19_957 ();
 sg13g2_decap_8 FILLER_19_964 ();
 sg13g2_decap_8 FILLER_19_971 ();
 sg13g2_decap_4 FILLER_19_978 ();
 sg13g2_fill_1 FILLER_19_982 ();
 sg13g2_fill_2 FILLER_19_988 ();
 sg13g2_fill_2 FILLER_19_997 ();
 sg13g2_fill_2 FILLER_19_1004 ();
 sg13g2_fill_1 FILLER_19_1006 ();
 sg13g2_decap_4 FILLER_19_1012 ();
 sg13g2_fill_2 FILLER_19_1016 ();
 sg13g2_decap_4 FILLER_19_1024 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_19_1045 ();
 sg13g2_fill_2 FILLER_19_1052 ();
 sg13g2_fill_2 FILLER_19_1068 ();
 sg13g2_fill_1 FILLER_19_1070 ();
 sg13g2_fill_1 FILLER_19_1075 ();
 sg13g2_fill_2 FILLER_19_1081 ();
 sg13g2_fill_2 FILLER_19_1091 ();
 sg13g2_fill_2 FILLER_19_1102 ();
 sg13g2_fill_1 FILLER_19_1104 ();
 sg13g2_fill_2 FILLER_19_1115 ();
 sg13g2_fill_1 FILLER_19_1117 ();
 sg13g2_fill_2 FILLER_19_1123 ();
 sg13g2_fill_1 FILLER_19_1125 ();
 sg13g2_decap_8 FILLER_19_1136 ();
 sg13g2_decap_8 FILLER_19_1143 ();
 sg13g2_fill_1 FILLER_19_1150 ();
 sg13g2_fill_1 FILLER_19_1160 ();
 sg13g2_fill_2 FILLER_19_1171 ();
 sg13g2_decap_4 FILLER_19_1181 ();
 sg13g2_decap_8 FILLER_19_1189 ();
 sg13g2_fill_2 FILLER_19_1229 ();
 sg13g2_decap_8 FILLER_19_1237 ();
 sg13g2_decap_8 FILLER_19_1244 ();
 sg13g2_fill_2 FILLER_19_1259 ();
 sg13g2_fill_1 FILLER_19_1261 ();
 sg13g2_decap_4 FILLER_19_1270 ();
 sg13g2_fill_2 FILLER_19_1274 ();
 sg13g2_decap_8 FILLER_19_1281 ();
 sg13g2_decap_4 FILLER_19_1323 ();
 sg13g2_fill_1 FILLER_19_1327 ();
 sg13g2_decap_8 FILLER_19_1337 ();
 sg13g2_decap_4 FILLER_19_1344 ();
 sg13g2_fill_1 FILLER_19_1348 ();
 sg13g2_decap_4 FILLER_19_1353 ();
 sg13g2_fill_1 FILLER_19_1357 ();
 sg13g2_fill_1 FILLER_19_1363 ();
 sg13g2_decap_4 FILLER_19_1385 ();
 sg13g2_decap_8 FILLER_19_1397 ();
 sg13g2_decap_8 FILLER_19_1404 ();
 sg13g2_fill_2 FILLER_19_1411 ();
 sg13g2_fill_1 FILLER_19_1413 ();
 sg13g2_fill_1 FILLER_19_1424 ();
 sg13g2_fill_1 FILLER_19_1430 ();
 sg13g2_fill_1 FILLER_19_1441 ();
 sg13g2_fill_1 FILLER_19_1446 ();
 sg13g2_fill_1 FILLER_19_1453 ();
 sg13g2_fill_2 FILLER_19_1463 ();
 sg13g2_fill_1 FILLER_19_1465 ();
 sg13g2_decap_8 FILLER_19_1471 ();
 sg13g2_fill_2 FILLER_19_1478 ();
 sg13g2_fill_1 FILLER_19_1480 ();
 sg13g2_fill_2 FILLER_19_1493 ();
 sg13g2_fill_1 FILLER_19_1563 ();
 sg13g2_fill_2 FILLER_19_1572 ();
 sg13g2_fill_1 FILLER_19_1574 ();
 sg13g2_decap_4 FILLER_19_1583 ();
 sg13g2_fill_1 FILLER_19_1587 ();
 sg13g2_fill_1 FILLER_19_1622 ();
 sg13g2_decap_4 FILLER_19_1631 ();
 sg13g2_fill_1 FILLER_19_1635 ();
 sg13g2_decap_8 FILLER_19_1641 ();
 sg13g2_fill_2 FILLER_19_1648 ();
 sg13g2_fill_2 FILLER_19_1668 ();
 sg13g2_fill_2 FILLER_19_1680 ();
 sg13g2_fill_1 FILLER_19_1682 ();
 sg13g2_decap_4 FILLER_19_1688 ();
 sg13g2_fill_2 FILLER_19_1692 ();
 sg13g2_fill_2 FILLER_19_1699 ();
 sg13g2_fill_1 FILLER_19_1701 ();
 sg13g2_decap_4 FILLER_19_1707 ();
 sg13g2_fill_2 FILLER_19_1711 ();
 sg13g2_fill_1 FILLER_19_1718 ();
 sg13g2_decap_4 FILLER_19_1723 ();
 sg13g2_decap_4 FILLER_19_1732 ();
 sg13g2_decap_8 FILLER_19_1745 ();
 sg13g2_decap_8 FILLER_19_1752 ();
 sg13g2_decap_8 FILLER_19_1759 ();
 sg13g2_decap_8 FILLER_19_1766 ();
 sg13g2_fill_1 FILLER_19_1773 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_30 ();
 sg13g2_fill_1 FILLER_20_32 ();
 sg13g2_fill_1 FILLER_20_61 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_87 ();
 sg13g2_decap_8 FILLER_20_94 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_1 FILLER_20_121 ();
 sg13g2_decap_4 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_135 ();
 sg13g2_fill_1 FILLER_20_140 ();
 sg13g2_decap_4 FILLER_20_149 ();
 sg13g2_fill_1 FILLER_20_153 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_decap_4 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_220 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_decap_4 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_342 ();
 sg13g2_fill_1 FILLER_20_349 ();
 sg13g2_fill_2 FILLER_20_358 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_fill_2 FILLER_20_398 ();
 sg13g2_fill_1 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_404 ();
 sg13g2_decap_8 FILLER_20_419 ();
 sg13g2_decap_8 FILLER_20_426 ();
 sg13g2_decap_8 FILLER_20_433 ();
 sg13g2_decap_8 FILLER_20_440 ();
 sg13g2_fill_1 FILLER_20_447 ();
 sg13g2_fill_2 FILLER_20_470 ();
 sg13g2_fill_1 FILLER_20_472 ();
 sg13g2_decap_8 FILLER_20_492 ();
 sg13g2_fill_2 FILLER_20_499 ();
 sg13g2_decap_4 FILLER_20_510 ();
 sg13g2_fill_2 FILLER_20_535 ();
 sg13g2_decap_4 FILLER_20_545 ();
 sg13g2_fill_1 FILLER_20_549 ();
 sg13g2_decap_8 FILLER_20_559 ();
 sg13g2_decap_8 FILLER_20_566 ();
 sg13g2_fill_1 FILLER_20_573 ();
 sg13g2_decap_4 FILLER_20_608 ();
 sg13g2_decap_8 FILLER_20_622 ();
 sg13g2_fill_2 FILLER_20_629 ();
 sg13g2_decap_8 FILLER_20_635 ();
 sg13g2_fill_1 FILLER_20_642 ();
 sg13g2_fill_1 FILLER_20_647 ();
 sg13g2_decap_4 FILLER_20_652 ();
 sg13g2_fill_1 FILLER_20_656 ();
 sg13g2_fill_2 FILLER_20_661 ();
 sg13g2_fill_1 FILLER_20_663 ();
 sg13g2_decap_8 FILLER_20_668 ();
 sg13g2_decap_4 FILLER_20_675 ();
 sg13g2_fill_2 FILLER_20_719 ();
 sg13g2_decap_4 FILLER_20_726 ();
 sg13g2_fill_1 FILLER_20_735 ();
 sg13g2_fill_1 FILLER_20_753 ();
 sg13g2_fill_2 FILLER_20_770 ();
 sg13g2_fill_1 FILLER_20_782 ();
 sg13g2_fill_1 FILLER_20_788 ();
 sg13g2_fill_2 FILLER_20_794 ();
 sg13g2_fill_1 FILLER_20_796 ();
 sg13g2_fill_1 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_820 ();
 sg13g2_fill_1 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_836 ();
 sg13g2_decap_8 FILLER_20_843 ();
 sg13g2_decap_8 FILLER_20_850 ();
 sg13g2_decap_8 FILLER_20_857 ();
 sg13g2_decap_8 FILLER_20_864 ();
 sg13g2_decap_8 FILLER_20_871 ();
 sg13g2_decap_4 FILLER_20_878 ();
 sg13g2_fill_1 FILLER_20_882 ();
 sg13g2_fill_2 FILLER_20_887 ();
 sg13g2_decap_8 FILLER_20_894 ();
 sg13g2_fill_2 FILLER_20_901 ();
 sg13g2_fill_2 FILLER_20_908 ();
 sg13g2_fill_1 FILLER_20_910 ();
 sg13g2_decap_8 FILLER_20_919 ();
 sg13g2_decap_8 FILLER_20_926 ();
 sg13g2_decap_8 FILLER_20_933 ();
 sg13g2_fill_2 FILLER_20_940 ();
 sg13g2_fill_1 FILLER_20_942 ();
 sg13g2_decap_4 FILLER_20_951 ();
 sg13g2_fill_2 FILLER_20_955 ();
 sg13g2_decap_8 FILLER_20_971 ();
 sg13g2_fill_2 FILLER_20_978 ();
 sg13g2_fill_1 FILLER_20_980 ();
 sg13g2_decap_4 FILLER_20_994 ();
 sg13g2_fill_1 FILLER_20_1003 ();
 sg13g2_fill_2 FILLER_20_1030 ();
 sg13g2_decap_4 FILLER_20_1036 ();
 sg13g2_fill_1 FILLER_20_1040 ();
 sg13g2_fill_1 FILLER_20_1059 ();
 sg13g2_fill_1 FILLER_20_1070 ();
 sg13g2_fill_1 FILLER_20_1076 ();
 sg13g2_fill_1 FILLER_20_1087 ();
 sg13g2_decap_4 FILLER_20_1098 ();
 sg13g2_fill_1 FILLER_20_1102 ();
 sg13g2_decap_8 FILLER_20_1180 ();
 sg13g2_fill_2 FILLER_20_1187 ();
 sg13g2_decap_8 FILLER_20_1198 ();
 sg13g2_decap_4 FILLER_20_1205 ();
 sg13g2_fill_2 FILLER_20_1209 ();
 sg13g2_decap_4 FILLER_20_1225 ();
 sg13g2_fill_1 FILLER_20_1229 ();
 sg13g2_decap_8 FILLER_20_1234 ();
 sg13g2_decap_8 FILLER_20_1241 ();
 sg13g2_decap_8 FILLER_20_1248 ();
 sg13g2_decap_8 FILLER_20_1255 ();
 sg13g2_decap_4 FILLER_20_1262 ();
 sg13g2_fill_1 FILLER_20_1271 ();
 sg13g2_fill_2 FILLER_20_1287 ();
 sg13g2_fill_1 FILLER_20_1289 ();
 sg13g2_fill_2 FILLER_20_1308 ();
 sg13g2_fill_1 FILLER_20_1310 ();
 sg13g2_fill_2 FILLER_20_1337 ();
 sg13g2_fill_1 FILLER_20_1339 ();
 sg13g2_decap_4 FILLER_20_1392 ();
 sg13g2_decap_8 FILLER_20_1409 ();
 sg13g2_fill_2 FILLER_20_1416 ();
 sg13g2_fill_2 FILLER_20_1430 ();
 sg13g2_fill_1 FILLER_20_1432 ();
 sg13g2_decap_8 FILLER_20_1464 ();
 sg13g2_fill_1 FILLER_20_1481 ();
 sg13g2_fill_1 FILLER_20_1491 ();
 sg13g2_fill_2 FILLER_20_1500 ();
 sg13g2_decap_4 FILLER_20_1516 ();
 sg13g2_fill_1 FILLER_20_1520 ();
 sg13g2_decap_4 FILLER_20_1529 ();
 sg13g2_fill_1 FILLER_20_1533 ();
 sg13g2_fill_1 FILLER_20_1539 ();
 sg13g2_fill_2 FILLER_20_1549 ();
 sg13g2_fill_1 FILLER_20_1566 ();
 sg13g2_fill_1 FILLER_20_1572 ();
 sg13g2_fill_2 FILLER_20_1581 ();
 sg13g2_decap_8 FILLER_20_1596 ();
 sg13g2_decap_8 FILLER_20_1603 ();
 sg13g2_decap_8 FILLER_20_1613 ();
 sg13g2_decap_8 FILLER_20_1620 ();
 sg13g2_fill_2 FILLER_20_1627 ();
 sg13g2_fill_2 FILLER_20_1637 ();
 sg13g2_decap_8 FILLER_20_1647 ();
 sg13g2_fill_2 FILLER_20_1654 ();
 sg13g2_fill_1 FILLER_20_1656 ();
 sg13g2_decap_8 FILLER_20_1716 ();
 sg13g2_decap_8 FILLER_20_1723 ();
 sg13g2_decap_8 FILLER_20_1734 ();
 sg13g2_decap_4 FILLER_20_1741 ();
 sg13g2_decap_8 FILLER_20_1748 ();
 sg13g2_decap_8 FILLER_20_1755 ();
 sg13g2_decap_8 FILLER_20_1762 ();
 sg13g2_decap_4 FILLER_20_1769 ();
 sg13g2_fill_1 FILLER_20_1773 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_20 ();
 sg13g2_fill_1 FILLER_21_22 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_fill_1 FILLER_21_50 ();
 sg13g2_decap_4 FILLER_21_68 ();
 sg13g2_decap_4 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_136 ();
 sg13g2_decap_4 FILLER_21_155 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_184 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_216 ();
 sg13g2_fill_2 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_244 ();
 sg13g2_decap_4 FILLER_21_249 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_275 ();
 sg13g2_fill_2 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_282 ();
 sg13g2_decap_8 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_4 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_fill_2 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_fill_2 FILLER_21_396 ();
 sg13g2_fill_1 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_415 ();
 sg13g2_fill_2 FILLER_21_445 ();
 sg13g2_fill_2 FILLER_21_465 ();
 sg13g2_fill_1 FILLER_21_472 ();
 sg13g2_decap_4 FILLER_21_487 ();
 sg13g2_fill_2 FILLER_21_533 ();
 sg13g2_fill_2 FILLER_21_548 ();
 sg13g2_decap_8 FILLER_21_554 ();
 sg13g2_decap_8 FILLER_21_561 ();
 sg13g2_fill_2 FILLER_21_568 ();
 sg13g2_fill_1 FILLER_21_570 ();
 sg13g2_fill_1 FILLER_21_575 ();
 sg13g2_decap_4 FILLER_21_581 ();
 sg13g2_fill_2 FILLER_21_585 ();
 sg13g2_fill_2 FILLER_21_598 ();
 sg13g2_fill_1 FILLER_21_600 ();
 sg13g2_decap_4 FILLER_21_616 ();
 sg13g2_fill_1 FILLER_21_625 ();
 sg13g2_fill_1 FILLER_21_631 ();
 sg13g2_fill_1 FILLER_21_637 ();
 sg13g2_fill_1 FILLER_21_651 ();
 sg13g2_fill_2 FILLER_21_657 ();
 sg13g2_decap_8 FILLER_21_664 ();
 sg13g2_fill_2 FILLER_21_671 ();
 sg13g2_fill_1 FILLER_21_673 ();
 sg13g2_fill_1 FILLER_21_693 ();
 sg13g2_fill_1 FILLER_21_713 ();
 sg13g2_fill_1 FILLER_21_725 ();
 sg13g2_fill_1 FILLER_21_731 ();
 sg13g2_fill_1 FILLER_21_754 ();
 sg13g2_fill_2 FILLER_21_775 ();
 sg13g2_fill_1 FILLER_21_782 ();
 sg13g2_decap_8 FILLER_21_820 ();
 sg13g2_decap_4 FILLER_21_827 ();
 sg13g2_fill_1 FILLER_21_831 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_4 FILLER_21_847 ();
 sg13g2_fill_1 FILLER_21_851 ();
 sg13g2_fill_2 FILLER_21_882 ();
 sg13g2_fill_1 FILLER_21_884 ();
 sg13g2_decap_4 FILLER_21_890 ();
 sg13g2_decap_8 FILLER_21_902 ();
 sg13g2_fill_2 FILLER_21_925 ();
 sg13g2_decap_4 FILLER_21_932 ();
 sg13g2_fill_2 FILLER_21_936 ();
 sg13g2_decap_8 FILLER_21_946 ();
 sg13g2_fill_1 FILLER_21_953 ();
 sg13g2_decap_8 FILLER_21_965 ();
 sg13g2_fill_1 FILLER_21_972 ();
 sg13g2_fill_2 FILLER_21_999 ();
 sg13g2_decap_4 FILLER_21_1006 ();
 sg13g2_fill_1 FILLER_21_1010 ();
 sg13g2_decap_4 FILLER_21_1015 ();
 sg13g2_decap_4 FILLER_21_1023 ();
 sg13g2_fill_1 FILLER_21_1027 ();
 sg13g2_fill_1 FILLER_21_1033 ();
 sg13g2_fill_2 FILLER_21_1046 ();
 sg13g2_decap_8 FILLER_21_1051 ();
 sg13g2_decap_8 FILLER_21_1058 ();
 sg13g2_decap_8 FILLER_21_1065 ();
 sg13g2_fill_2 FILLER_21_1072 ();
 sg13g2_fill_1 FILLER_21_1074 ();
 sg13g2_decap_8 FILLER_21_1089 ();
 sg13g2_fill_2 FILLER_21_1096 ();
 sg13g2_decap_8 FILLER_21_1120 ();
 sg13g2_decap_8 FILLER_21_1127 ();
 sg13g2_decap_4 FILLER_21_1138 ();
 sg13g2_fill_1 FILLER_21_1142 ();
 sg13g2_decap_4 FILLER_21_1156 ();
 sg13g2_fill_1 FILLER_21_1160 ();
 sg13g2_fill_1 FILLER_21_1177 ();
 sg13g2_decap_8 FILLER_21_1182 ();
 sg13g2_decap_8 FILLER_21_1189 ();
 sg13g2_fill_2 FILLER_21_1196 ();
 sg13g2_fill_1 FILLER_21_1198 ();
 sg13g2_decap_8 FILLER_21_1207 ();
 sg13g2_decap_8 FILLER_21_1214 ();
 sg13g2_fill_2 FILLER_21_1221 ();
 sg13g2_fill_1 FILLER_21_1223 ();
 sg13g2_fill_2 FILLER_21_1239 ();
 sg13g2_decap_8 FILLER_21_1245 ();
 sg13g2_decap_8 FILLER_21_1260 ();
 sg13g2_decap_8 FILLER_21_1267 ();
 sg13g2_decap_8 FILLER_21_1274 ();
 sg13g2_fill_1 FILLER_21_1281 ();
 sg13g2_fill_1 FILLER_21_1319 ();
 sg13g2_fill_1 FILLER_21_1324 ();
 sg13g2_fill_2 FILLER_21_1330 ();
 sg13g2_decap_4 FILLER_21_1336 ();
 sg13g2_fill_2 FILLER_21_1346 ();
 sg13g2_fill_2 FILLER_21_1360 ();
 sg13g2_fill_2 FILLER_21_1374 ();
 sg13g2_fill_1 FILLER_21_1376 ();
 sg13g2_fill_1 FILLER_21_1385 ();
 sg13g2_decap_8 FILLER_21_1408 ();
 sg13g2_decap_8 FILLER_21_1415 ();
 sg13g2_decap_8 FILLER_21_1426 ();
 sg13g2_decap_4 FILLER_21_1433 ();
 sg13g2_fill_2 FILLER_21_1437 ();
 sg13g2_decap_8 FILLER_21_1447 ();
 sg13g2_decap_8 FILLER_21_1454 ();
 sg13g2_fill_2 FILLER_21_1466 ();
 sg13g2_fill_2 FILLER_21_1473 ();
 sg13g2_fill_1 FILLER_21_1475 ();
 sg13g2_fill_1 FILLER_21_1481 ();
 sg13g2_fill_1 FILLER_21_1508 ();
 sg13g2_decap_4 FILLER_21_1536 ();
 sg13g2_fill_2 FILLER_21_1540 ();
 sg13g2_fill_1 FILLER_21_1553 ();
 sg13g2_decap_4 FILLER_21_1600 ();
 sg13g2_decap_8 FILLER_21_1626 ();
 sg13g2_decap_4 FILLER_21_1638 ();
 sg13g2_fill_2 FILLER_21_1642 ();
 sg13g2_decap_4 FILLER_21_1652 ();
 sg13g2_decap_8 FILLER_21_1664 ();
 sg13g2_decap_4 FILLER_21_1671 ();
 sg13g2_fill_1 FILLER_21_1675 ();
 sg13g2_fill_1 FILLER_21_1681 ();
 sg13g2_fill_1 FILLER_21_1693 ();
 sg13g2_decap_8 FILLER_21_1729 ();
 sg13g2_decap_8 FILLER_21_1736 ();
 sg13g2_decap_8 FILLER_21_1743 ();
 sg13g2_decap_8 FILLER_21_1750 ();
 sg13g2_decap_8 FILLER_21_1757 ();
 sg13g2_decap_8 FILLER_21_1764 ();
 sg13g2_fill_2 FILLER_21_1771 ();
 sg13g2_fill_1 FILLER_21_1773 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_9 ();
 sg13g2_fill_2 FILLER_22_24 ();
 sg13g2_fill_1 FILLER_22_30 ();
 sg13g2_fill_2 FILLER_22_46 ();
 sg13g2_decap_4 FILLER_22_59 ();
 sg13g2_fill_1 FILLER_22_63 ();
 sg13g2_fill_2 FILLER_22_69 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_fill_2 FILLER_22_136 ();
 sg13g2_fill_1 FILLER_22_138 ();
 sg13g2_decap_4 FILLER_22_144 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_1 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_4 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_230 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_4 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_265 ();
 sg13g2_decap_8 FILLER_22_276 ();
 sg13g2_decap_4 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_287 ();
 sg13g2_fill_2 FILLER_22_309 ();
 sg13g2_fill_1 FILLER_22_311 ();
 sg13g2_fill_2 FILLER_22_336 ();
 sg13g2_fill_1 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_370 ();
 sg13g2_fill_2 FILLER_22_379 ();
 sg13g2_decap_4 FILLER_22_389 ();
 sg13g2_fill_2 FILLER_22_401 ();
 sg13g2_decap_4 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_22_416 ();
 sg13g2_fill_1 FILLER_22_432 ();
 sg13g2_fill_1 FILLER_22_438 ();
 sg13g2_fill_1 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_453 ();
 sg13g2_fill_2 FILLER_22_460 ();
 sg13g2_decap_4 FILLER_22_471 ();
 sg13g2_decap_4 FILLER_22_480 ();
 sg13g2_fill_2 FILLER_22_484 ();
 sg13g2_fill_2 FILLER_22_507 ();
 sg13g2_fill_2 FILLER_22_514 ();
 sg13g2_decap_8 FILLER_22_521 ();
 sg13g2_decap_4 FILLER_22_528 ();
 sg13g2_fill_2 FILLER_22_536 ();
 sg13g2_fill_1 FILLER_22_542 ();
 sg13g2_decap_8 FILLER_22_559 ();
 sg13g2_decap_4 FILLER_22_566 ();
 sg13g2_fill_1 FILLER_22_590 ();
 sg13g2_decap_8 FILLER_22_596 ();
 sg13g2_fill_1 FILLER_22_603 ();
 sg13g2_fill_2 FILLER_22_611 ();
 sg13g2_fill_1 FILLER_22_613 ();
 sg13g2_fill_2 FILLER_22_645 ();
 sg13g2_fill_1 FILLER_22_647 ();
 sg13g2_decap_8 FILLER_22_656 ();
 sg13g2_decap_4 FILLER_22_663 ();
 sg13g2_fill_2 FILLER_22_667 ();
 sg13g2_decap_8 FILLER_22_673 ();
 sg13g2_fill_1 FILLER_22_704 ();
 sg13g2_fill_1 FILLER_22_734 ();
 sg13g2_fill_1 FILLER_22_746 ();
 sg13g2_fill_2 FILLER_22_752 ();
 sg13g2_fill_1 FILLER_22_754 ();
 sg13g2_fill_1 FILLER_22_770 ();
 sg13g2_decap_4 FILLER_22_787 ();
 sg13g2_fill_1 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_4 FILLER_22_816 ();
 sg13g2_fill_2 FILLER_22_820 ();
 sg13g2_fill_2 FILLER_22_836 ();
 sg13g2_decap_8 FILLER_22_846 ();
 sg13g2_decap_8 FILLER_22_853 ();
 sg13g2_fill_2 FILLER_22_860 ();
 sg13g2_decap_4 FILLER_22_866 ();
 sg13g2_fill_1 FILLER_22_870 ();
 sg13g2_decap_8 FILLER_22_886 ();
 sg13g2_fill_1 FILLER_22_893 ();
 sg13g2_decap_4 FILLER_22_897 ();
 sg13g2_fill_1 FILLER_22_909 ();
 sg13g2_decap_4 FILLER_22_939 ();
 sg13g2_fill_2 FILLER_22_943 ();
 sg13g2_fill_2 FILLER_22_975 ();
 sg13g2_fill_1 FILLER_22_977 ();
 sg13g2_fill_1 FILLER_22_991 ();
 sg13g2_fill_1 FILLER_22_996 ();
 sg13g2_decap_8 FILLER_22_1006 ();
 sg13g2_decap_8 FILLER_22_1013 ();
 sg13g2_fill_1 FILLER_22_1024 ();
 sg13g2_decap_4 FILLER_22_1040 ();
 sg13g2_decap_4 FILLER_22_1049 ();
 sg13g2_fill_1 FILLER_22_1061 ();
 sg13g2_fill_2 FILLER_22_1077 ();
 sg13g2_fill_1 FILLER_22_1079 ();
 sg13g2_decap_4 FILLER_22_1088 ();
 sg13g2_fill_1 FILLER_22_1092 ();
 sg13g2_decap_4 FILLER_22_1112 ();
 sg13g2_decap_8 FILLER_22_1119 ();
 sg13g2_fill_2 FILLER_22_1126 ();
 sg13g2_fill_1 FILLER_22_1128 ();
 sg13g2_decap_4 FILLER_22_1133 ();
 sg13g2_fill_2 FILLER_22_1137 ();
 sg13g2_decap_8 FILLER_22_1144 ();
 sg13g2_decap_4 FILLER_22_1151 ();
 sg13g2_fill_2 FILLER_22_1155 ();
 sg13g2_decap_4 FILLER_22_1160 ();
 sg13g2_decap_8 FILLER_22_1209 ();
 sg13g2_fill_2 FILLER_22_1216 ();
 sg13g2_fill_1 FILLER_22_1218 ();
 sg13g2_decap_4 FILLER_22_1232 ();
 sg13g2_fill_1 FILLER_22_1240 ();
 sg13g2_fill_2 FILLER_22_1247 ();
 sg13g2_decap_8 FILLER_22_1259 ();
 sg13g2_fill_1 FILLER_22_1266 ();
 sg13g2_fill_2 FILLER_22_1289 ();
 sg13g2_fill_2 FILLER_22_1302 ();
 sg13g2_fill_1 FILLER_22_1304 ();
 sg13g2_decap_8 FILLER_22_1318 ();
 sg13g2_decap_4 FILLER_22_1325 ();
 sg13g2_fill_2 FILLER_22_1329 ();
 sg13g2_fill_1 FILLER_22_1377 ();
 sg13g2_fill_2 FILLER_22_1390 ();
 sg13g2_fill_1 FILLER_22_1392 ();
 sg13g2_decap_8 FILLER_22_1398 ();
 sg13g2_fill_1 FILLER_22_1405 ();
 sg13g2_decap_8 FILLER_22_1428 ();
 sg13g2_fill_2 FILLER_22_1435 ();
 sg13g2_fill_1 FILLER_22_1437 ();
 sg13g2_decap_8 FILLER_22_1442 ();
 sg13g2_decap_8 FILLER_22_1449 ();
 sg13g2_decap_8 FILLER_22_1456 ();
 sg13g2_fill_1 FILLER_22_1463 ();
 sg13g2_fill_2 FILLER_22_1477 ();
 sg13g2_fill_1 FILLER_22_1479 ();
 sg13g2_fill_2 FILLER_22_1485 ();
 sg13g2_fill_1 FILLER_22_1487 ();
 sg13g2_fill_2 FILLER_22_1508 ();
 sg13g2_decap_8 FILLER_22_1514 ();
 sg13g2_decap_4 FILLER_22_1521 ();
 sg13g2_fill_2 FILLER_22_1525 ();
 sg13g2_decap_8 FILLER_22_1531 ();
 sg13g2_decap_4 FILLER_22_1538 ();
 sg13g2_fill_1 FILLER_22_1547 ();
 sg13g2_fill_2 FILLER_22_1556 ();
 sg13g2_fill_1 FILLER_22_1558 ();
 sg13g2_fill_1 FILLER_22_1572 ();
 sg13g2_fill_1 FILLER_22_1582 ();
 sg13g2_decap_4 FILLER_22_1586 ();
 sg13g2_fill_2 FILLER_22_1595 ();
 sg13g2_fill_1 FILLER_22_1601 ();
 sg13g2_fill_1 FILLER_22_1607 ();
 sg13g2_decap_8 FILLER_22_1615 ();
 sg13g2_fill_1 FILLER_22_1622 ();
 sg13g2_decap_4 FILLER_22_1627 ();
 sg13g2_fill_1 FILLER_22_1631 ();
 sg13g2_decap_8 FILLER_22_1640 ();
 sg13g2_decap_4 FILLER_22_1647 ();
 sg13g2_fill_1 FILLER_22_1651 ();
 sg13g2_fill_2 FILLER_22_1656 ();
 sg13g2_fill_2 FILLER_22_1666 ();
 sg13g2_fill_2 FILLER_22_1673 ();
 sg13g2_fill_1 FILLER_22_1675 ();
 sg13g2_fill_1 FILLER_22_1743 ();
 sg13g2_decap_8 FILLER_22_1748 ();
 sg13g2_decap_8 FILLER_22_1755 ();
 sg13g2_decap_8 FILLER_22_1762 ();
 sg13g2_decap_4 FILLER_22_1769 ();
 sg13g2_fill_1 FILLER_22_1773 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_32 ();
 sg13g2_fill_1 FILLER_23_46 ();
 sg13g2_decap_4 FILLER_23_74 ();
 sg13g2_fill_1 FILLER_23_78 ();
 sg13g2_fill_1 FILLER_23_89 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_fill_2 FILLER_23_120 ();
 sg13g2_fill_1 FILLER_23_137 ();
 sg13g2_decap_4 FILLER_23_142 ();
 sg13g2_fill_2 FILLER_23_151 ();
 sg13g2_fill_1 FILLER_23_158 ();
 sg13g2_fill_2 FILLER_23_164 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_177 ();
 sg13g2_decap_4 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_188 ();
 sg13g2_decap_4 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_205 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_decap_4 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_decap_8 FILLER_23_265 ();
 sg13g2_decap_8 FILLER_23_272 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_4 FILLER_23_291 ();
 sg13g2_fill_2 FILLER_23_299 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_4 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_fill_1 FILLER_23_392 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_2 FILLER_23_418 ();
 sg13g2_decap_4 FILLER_23_444 ();
 sg13g2_fill_2 FILLER_23_453 ();
 sg13g2_fill_2 FILLER_23_463 ();
 sg13g2_decap_8 FILLER_23_481 ();
 sg13g2_decap_4 FILLER_23_493 ();
 sg13g2_fill_1 FILLER_23_497 ();
 sg13g2_fill_2 FILLER_23_502 ();
 sg13g2_decap_8 FILLER_23_515 ();
 sg13g2_decap_4 FILLER_23_522 ();
 sg13g2_fill_2 FILLER_23_541 ();
 sg13g2_fill_1 FILLER_23_563 ();
 sg13g2_decap_4 FILLER_23_568 ();
 sg13g2_decap_8 FILLER_23_594 ();
 sg13g2_fill_2 FILLER_23_601 ();
 sg13g2_fill_1 FILLER_23_603 ();
 sg13g2_fill_1 FILLER_23_608 ();
 sg13g2_fill_1 FILLER_23_615 ();
 sg13g2_fill_1 FILLER_23_624 ();
 sg13g2_fill_2 FILLER_23_631 ();
 sg13g2_fill_1 FILLER_23_641 ();
 sg13g2_fill_1 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_657 ();
 sg13g2_decap_8 FILLER_23_664 ();
 sg13g2_decap_4 FILLER_23_671 ();
 sg13g2_fill_1 FILLER_23_675 ();
 sg13g2_fill_1 FILLER_23_680 ();
 sg13g2_fill_1 FILLER_23_701 ();
 sg13g2_fill_2 FILLER_23_720 ();
 sg13g2_fill_2 FILLER_23_735 ();
 sg13g2_fill_1 FILLER_23_799 ();
 sg13g2_fill_1 FILLER_23_803 ();
 sg13g2_fill_2 FILLER_23_809 ();
 sg13g2_fill_1 FILLER_23_811 ();
 sg13g2_fill_2 FILLER_23_824 ();
 sg13g2_fill_1 FILLER_23_826 ();
 sg13g2_decap_4 FILLER_23_839 ();
 sg13g2_fill_2 FILLER_23_843 ();
 sg13g2_decap_4 FILLER_23_884 ();
 sg13g2_decap_8 FILLER_23_903 ();
 sg13g2_decap_8 FILLER_23_929 ();
 sg13g2_fill_2 FILLER_23_936 ();
 sg13g2_fill_1 FILLER_23_938 ();
 sg13g2_fill_2 FILLER_23_943 ();
 sg13g2_fill_1 FILLER_23_945 ();
 sg13g2_decap_8 FILLER_23_962 ();
 sg13g2_decap_4 FILLER_23_969 ();
 sg13g2_fill_2 FILLER_23_981 ();
 sg13g2_decap_4 FILLER_23_1004 ();
 sg13g2_fill_1 FILLER_23_1008 ();
 sg13g2_decap_4 FILLER_23_1035 ();
 sg13g2_fill_1 FILLER_23_1039 ();
 sg13g2_decap_4 FILLER_23_1053 ();
 sg13g2_fill_1 FILLER_23_1061 ();
 sg13g2_decap_4 FILLER_23_1070 ();
 sg13g2_fill_2 FILLER_23_1089 ();
 sg13g2_fill_1 FILLER_23_1091 ();
 sg13g2_decap_8 FILLER_23_1097 ();
 sg13g2_fill_2 FILLER_23_1104 ();
 sg13g2_decap_8 FILLER_23_1111 ();
 sg13g2_decap_8 FILLER_23_1118 ();
 sg13g2_fill_2 FILLER_23_1125 ();
 sg13g2_fill_1 FILLER_23_1127 ();
 sg13g2_decap_4 FILLER_23_1133 ();
 sg13g2_fill_1 FILLER_23_1137 ();
 sg13g2_decap_8 FILLER_23_1185 ();
 sg13g2_fill_1 FILLER_23_1192 ();
 sg13g2_decap_8 FILLER_23_1214 ();
 sg13g2_fill_2 FILLER_23_1221 ();
 sg13g2_fill_1 FILLER_23_1223 ();
 sg13g2_decap_8 FILLER_23_1232 ();
 sg13g2_fill_1 FILLER_23_1244 ();
 sg13g2_fill_1 FILLER_23_1254 ();
 sg13g2_decap_8 FILLER_23_1287 ();
 sg13g2_fill_2 FILLER_23_1294 ();
 sg13g2_decap_8 FILLER_23_1312 ();
 sg13g2_decap_8 FILLER_23_1319 ();
 sg13g2_fill_1 FILLER_23_1372 ();
 sg13g2_decap_8 FILLER_23_1388 ();
 sg13g2_decap_8 FILLER_23_1395 ();
 sg13g2_decap_4 FILLER_23_1402 ();
 sg13g2_fill_2 FILLER_23_1406 ();
 sg13g2_fill_1 FILLER_23_1441 ();
 sg13g2_decap_8 FILLER_23_1450 ();
 sg13g2_fill_1 FILLER_23_1457 ();
 sg13g2_decap_4 FILLER_23_1466 ();
 sg13g2_decap_8 FILLER_23_1474 ();
 sg13g2_fill_1 FILLER_23_1481 ();
 sg13g2_fill_2 FILLER_23_1495 ();
 sg13g2_fill_1 FILLER_23_1497 ();
 sg13g2_decap_4 FILLER_23_1529 ();
 sg13g2_fill_1 FILLER_23_1533 ();
 sg13g2_fill_2 FILLER_23_1537 ();
 sg13g2_fill_1 FILLER_23_1539 ();
 sg13g2_fill_2 FILLER_23_1544 ();
 sg13g2_fill_1 FILLER_23_1546 ();
 sg13g2_fill_1 FILLER_23_1556 ();
 sg13g2_fill_1 FILLER_23_1568 ();
 sg13g2_decap_4 FILLER_23_1587 ();
 sg13g2_fill_2 FILLER_23_1591 ();
 sg13g2_decap_4 FILLER_23_1597 ();
 sg13g2_fill_2 FILLER_23_1601 ();
 sg13g2_fill_1 FILLER_23_1626 ();
 sg13g2_fill_1 FILLER_23_1640 ();
 sg13g2_decap_8 FILLER_23_1646 ();
 sg13g2_decap_8 FILLER_23_1653 ();
 sg13g2_fill_2 FILLER_23_1660 ();
 sg13g2_fill_1 FILLER_23_1662 ();
 sg13g2_fill_2 FILLER_23_1682 ();
 sg13g2_fill_2 FILLER_23_1703 ();
 sg13g2_decap_8 FILLER_23_1760 ();
 sg13g2_decap_8 FILLER_23_1767 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_32 ();
 sg13g2_fill_1 FILLER_24_36 ();
 sg13g2_decap_8 FILLER_24_47 ();
 sg13g2_fill_1 FILLER_24_54 ();
 sg13g2_decap_4 FILLER_24_76 ();
 sg13g2_fill_1 FILLER_24_80 ();
 sg13g2_fill_2 FILLER_24_86 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_fill_2 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_110 ();
 sg13g2_fill_1 FILLER_24_121 ();
 sg13g2_fill_1 FILLER_24_135 ();
 sg13g2_decap_4 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_fill_2 FILLER_24_166 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_decap_8 FILLER_24_211 ();
 sg13g2_fill_1 FILLER_24_218 ();
 sg13g2_decap_4 FILLER_24_223 ();
 sg13g2_fill_2 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_326 ();
 sg13g2_fill_1 FILLER_24_331 ();
 sg13g2_decap_4 FILLER_24_337 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_decap_4 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_351 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_2 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_4 FILLER_24_402 ();
 sg13g2_fill_1 FILLER_24_416 ();
 sg13g2_fill_1 FILLER_24_422 ();
 sg13g2_fill_1 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_433 ();
 sg13g2_decap_8 FILLER_24_449 ();
 sg13g2_decap_8 FILLER_24_456 ();
 sg13g2_fill_2 FILLER_24_463 ();
 sg13g2_fill_1 FILLER_24_465 ();
 sg13g2_fill_2 FILLER_24_488 ();
 sg13g2_fill_1 FILLER_24_490 ();
 sg13g2_decap_4 FILLER_24_499 ();
 sg13g2_decap_8 FILLER_24_519 ();
 sg13g2_fill_2 FILLER_24_526 ();
 sg13g2_fill_2 FILLER_24_548 ();
 sg13g2_fill_1 FILLER_24_550 ();
 sg13g2_decap_8 FILLER_24_559 ();
 sg13g2_decap_8 FILLER_24_566 ();
 sg13g2_decap_4 FILLER_24_573 ();
 sg13g2_fill_1 FILLER_24_577 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_605 ();
 sg13g2_decap_8 FILLER_24_619 ();
 sg13g2_decap_4 FILLER_24_626 ();
 sg13g2_fill_1 FILLER_24_630 ();
 sg13g2_fill_2 FILLER_24_647 ();
 sg13g2_decap_4 FILLER_24_654 ();
 sg13g2_decap_8 FILLER_24_666 ();
 sg13g2_fill_2 FILLER_24_673 ();
 sg13g2_fill_1 FILLER_24_675 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_4 FILLER_24_708 ();
 sg13g2_fill_1 FILLER_24_712 ();
 sg13g2_fill_2 FILLER_24_727 ();
 sg13g2_fill_1 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_741 ();
 sg13g2_decap_8 FILLER_24_748 ();
 sg13g2_decap_8 FILLER_24_755 ();
 sg13g2_fill_1 FILLER_24_762 ();
 sg13g2_decap_4 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_fill_2 FILLER_24_791 ();
 sg13g2_fill_2 FILLER_24_797 ();
 sg13g2_fill_1 FILLER_24_828 ();
 sg13g2_fill_1 FILLER_24_837 ();
 sg13g2_decap_8 FILLER_24_851 ();
 sg13g2_decap_8 FILLER_24_858 ();
 sg13g2_decap_4 FILLER_24_865 ();
 sg13g2_fill_2 FILLER_24_869 ();
 sg13g2_fill_2 FILLER_24_892 ();
 sg13g2_fill_1 FILLER_24_894 ();
 sg13g2_decap_8 FILLER_24_904 ();
 sg13g2_decap_4 FILLER_24_911 ();
 sg13g2_fill_2 FILLER_24_915 ();
 sg13g2_decap_4 FILLER_24_923 ();
 sg13g2_decap_4 FILLER_24_931 ();
 sg13g2_fill_2 FILLER_24_935 ();
 sg13g2_fill_1 FILLER_24_949 ();
 sg13g2_fill_2 FILLER_24_955 ();
 sg13g2_fill_1 FILLER_24_957 ();
 sg13g2_decap_8 FILLER_24_962 ();
 sg13g2_decap_4 FILLER_24_969 ();
 sg13g2_fill_2 FILLER_24_973 ();
 sg13g2_fill_2 FILLER_24_983 ();
 sg13g2_decap_8 FILLER_24_988 ();
 sg13g2_fill_2 FILLER_24_995 ();
 sg13g2_fill_1 FILLER_24_1001 ();
 sg13g2_fill_1 FILLER_24_1038 ();
 sg13g2_decap_4 FILLER_24_1043 ();
 sg13g2_fill_2 FILLER_24_1047 ();
 sg13g2_fill_1 FILLER_24_1054 ();
 sg13g2_fill_2 FILLER_24_1060 ();
 sg13g2_fill_1 FILLER_24_1067 ();
 sg13g2_decap_8 FILLER_24_1092 ();
 sg13g2_fill_1 FILLER_24_1117 ();
 sg13g2_decap_8 FILLER_24_1126 ();
 sg13g2_decap_8 FILLER_24_1133 ();
 sg13g2_fill_2 FILLER_24_1140 ();
 sg13g2_decap_4 FILLER_24_1150 ();
 sg13g2_fill_2 FILLER_24_1184 ();
 sg13g2_decap_4 FILLER_24_1191 ();
 sg13g2_fill_2 FILLER_24_1195 ();
 sg13g2_fill_2 FILLER_24_1206 ();
 sg13g2_fill_2 FILLER_24_1213 ();
 sg13g2_fill_1 FILLER_24_1215 ();
 sg13g2_decap_4 FILLER_24_1220 ();
 sg13g2_decap_8 FILLER_24_1250 ();
 sg13g2_fill_2 FILLER_24_1262 ();
 sg13g2_decap_4 FILLER_24_1286 ();
 sg13g2_fill_2 FILLER_24_1290 ();
 sg13g2_fill_1 FILLER_24_1318 ();
 sg13g2_fill_2 FILLER_24_1323 ();
 sg13g2_fill_1 FILLER_24_1345 ();
 sg13g2_fill_1 FILLER_24_1371 ();
 sg13g2_fill_1 FILLER_24_1382 ();
 sg13g2_fill_1 FILLER_24_1393 ();
 sg13g2_fill_1 FILLER_24_1399 ();
 sg13g2_fill_2 FILLER_24_1404 ();
 sg13g2_decap_4 FILLER_24_1411 ();
 sg13g2_fill_2 FILLER_24_1415 ();
 sg13g2_decap_8 FILLER_24_1439 ();
 sg13g2_decap_4 FILLER_24_1446 ();
 sg13g2_decap_8 FILLER_24_1459 ();
 sg13g2_fill_1 FILLER_24_1470 ();
 sg13g2_decap_8 FILLER_24_1476 ();
 sg13g2_fill_1 FILLER_24_1483 ();
 sg13g2_fill_1 FILLER_24_1499 ();
 sg13g2_fill_2 FILLER_24_1566 ();
 sg13g2_fill_1 FILLER_24_1568 ();
 sg13g2_fill_2 FILLER_24_1573 ();
 sg13g2_fill_1 FILLER_24_1575 ();
 sg13g2_fill_2 FILLER_24_1587 ();
 sg13g2_fill_1 FILLER_24_1593 ();
 sg13g2_fill_2 FILLER_24_1630 ();
 sg13g2_fill_1 FILLER_24_1632 ();
 sg13g2_decap_8 FILLER_24_1642 ();
 sg13g2_decap_4 FILLER_24_1649 ();
 sg13g2_fill_1 FILLER_24_1683 ();
 sg13g2_decap_8 FILLER_24_1694 ();
 sg13g2_fill_2 FILLER_24_1701 ();
 sg13g2_fill_1 FILLER_24_1703 ();
 sg13g2_fill_2 FILLER_24_1712 ();
 sg13g2_fill_1 FILLER_24_1738 ();
 sg13g2_fill_2 FILLER_24_1743 ();
 sg13g2_fill_1 FILLER_24_1750 ();
 sg13g2_fill_1 FILLER_24_1755 ();
 sg13g2_fill_2 FILLER_24_1761 ();
 sg13g2_decap_4 FILLER_24_1768 ();
 sg13g2_fill_2 FILLER_24_1772 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_fill_2 FILLER_25_18 ();
 sg13g2_fill_1 FILLER_25_20 ();
 sg13g2_decap_8 FILLER_25_29 ();
 sg13g2_decap_8 FILLER_25_36 ();
 sg13g2_decap_8 FILLER_25_43 ();
 sg13g2_fill_2 FILLER_25_50 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_61 ();
 sg13g2_decap_8 FILLER_25_76 ();
 sg13g2_decap_8 FILLER_25_100 ();
 sg13g2_decap_4 FILLER_25_107 ();
 sg13g2_fill_2 FILLER_25_111 ();
 sg13g2_fill_2 FILLER_25_117 ();
 sg13g2_decap_4 FILLER_25_122 ();
 sg13g2_fill_2 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_decap_8 FILLER_25_176 ();
 sg13g2_decap_4 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_fill_2 FILLER_25_206 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_decap_8 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_decap_4 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_285 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_decap_8 FILLER_25_298 ();
 sg13g2_fill_1 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_321 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_decap_4 FILLER_25_337 ();
 sg13g2_fill_2 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_fill_1 FILLER_25_399 ();
 sg13g2_decap_4 FILLER_25_439 ();
 sg13g2_fill_1 FILLER_25_443 ();
 sg13g2_decap_4 FILLER_25_448 ();
 sg13g2_fill_1 FILLER_25_481 ();
 sg13g2_fill_2 FILLER_25_486 ();
 sg13g2_fill_1 FILLER_25_488 ();
 sg13g2_fill_2 FILLER_25_493 ();
 sg13g2_fill_1 FILLER_25_495 ();
 sg13g2_decap_8 FILLER_25_501 ();
 sg13g2_fill_2 FILLER_25_515 ();
 sg13g2_fill_1 FILLER_25_517 ();
 sg13g2_decap_8 FILLER_25_565 ();
 sg13g2_decap_8 FILLER_25_572 ();
 sg13g2_decap_8 FILLER_25_579 ();
 sg13g2_decap_4 FILLER_25_586 ();
 sg13g2_fill_2 FILLER_25_608 ();
 sg13g2_fill_1 FILLER_25_610 ();
 sg13g2_fill_2 FILLER_25_619 ();
 sg13g2_fill_1 FILLER_25_621 ();
 sg13g2_fill_2 FILLER_25_627 ();
 sg13g2_decap_4 FILLER_25_634 ();
 sg13g2_fill_1 FILLER_25_645 ();
 sg13g2_fill_2 FILLER_25_680 ();
 sg13g2_decap_4 FILLER_25_727 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_4 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_764 ();
 sg13g2_decap_8 FILLER_25_771 ();
 sg13g2_fill_2 FILLER_25_778 ();
 sg13g2_fill_1 FILLER_25_780 ();
 sg13g2_fill_2 FILLER_25_795 ();
 sg13g2_decap_4 FILLER_25_807 ();
 sg13g2_fill_1 FILLER_25_811 ();
 sg13g2_fill_1 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_830 ();
 sg13g2_fill_2 FILLER_25_837 ();
 sg13g2_fill_1 FILLER_25_839 ();
 sg13g2_decap_8 FILLER_25_850 ();
 sg13g2_decap_8 FILLER_25_857 ();
 sg13g2_decap_4 FILLER_25_864 ();
 sg13g2_fill_2 FILLER_25_877 ();
 sg13g2_fill_1 FILLER_25_888 ();
 sg13g2_fill_2 FILLER_25_907 ();
 sg13g2_decap_4 FILLER_25_914 ();
 sg13g2_fill_2 FILLER_25_918 ();
 sg13g2_decap_4 FILLER_25_954 ();
 sg13g2_fill_1 FILLER_25_958 ();
 sg13g2_decap_4 FILLER_25_967 ();
 sg13g2_fill_2 FILLER_25_971 ();
 sg13g2_fill_1 FILLER_25_994 ();
 sg13g2_fill_2 FILLER_25_1003 ();
 sg13g2_decap_8 FILLER_25_1015 ();
 sg13g2_decap_8 FILLER_25_1022 ();
 sg13g2_decap_4 FILLER_25_1029 ();
 sg13g2_fill_2 FILLER_25_1033 ();
 sg13g2_fill_2 FILLER_25_1039 ();
 sg13g2_fill_1 FILLER_25_1041 ();
 sg13g2_decap_8 FILLER_25_1050 ();
 sg13g2_fill_1 FILLER_25_1072 ();
 sg13g2_decap_8 FILLER_25_1078 ();
 sg13g2_fill_1 FILLER_25_1085 ();
 sg13g2_decap_8 FILLER_25_1095 ();
 sg13g2_decap_8 FILLER_25_1102 ();
 sg13g2_fill_1 FILLER_25_1109 ();
 sg13g2_fill_2 FILLER_25_1120 ();
 sg13g2_fill_1 FILLER_25_1122 ();
 sg13g2_decap_4 FILLER_25_1128 ();
 sg13g2_fill_2 FILLER_25_1136 ();
 sg13g2_decap_4 FILLER_25_1154 ();
 sg13g2_decap_8 FILLER_25_1163 ();
 sg13g2_decap_8 FILLER_25_1170 ();
 sg13g2_decap_8 FILLER_25_1177 ();
 sg13g2_decap_4 FILLER_25_1184 ();
 sg13g2_fill_2 FILLER_25_1188 ();
 sg13g2_decap_4 FILLER_25_1206 ();
 sg13g2_fill_2 FILLER_25_1210 ();
 sg13g2_decap_4 FILLER_25_1221 ();
 sg13g2_fill_1 FILLER_25_1225 ();
 sg13g2_fill_1 FILLER_25_1231 ();
 sg13g2_fill_2 FILLER_25_1250 ();
 sg13g2_fill_1 FILLER_25_1263 ();
 sg13g2_fill_2 FILLER_25_1280 ();
 sg13g2_decap_4 FILLER_25_1287 ();
 sg13g2_fill_1 FILLER_25_1299 ();
 sg13g2_decap_4 FILLER_25_1309 ();
 sg13g2_fill_2 FILLER_25_1332 ();
 sg13g2_fill_1 FILLER_25_1339 ();
 sg13g2_fill_1 FILLER_25_1372 ();
 sg13g2_decap_4 FILLER_25_1389 ();
 sg13g2_decap_8 FILLER_25_1417 ();
 sg13g2_decap_4 FILLER_25_1424 ();
 sg13g2_decap_4 FILLER_25_1436 ();
 sg13g2_fill_2 FILLER_25_1440 ();
 sg13g2_decap_8 FILLER_25_1459 ();
 sg13g2_decap_4 FILLER_25_1466 ();
 sg13g2_fill_2 FILLER_25_1481 ();
 sg13g2_decap_4 FILLER_25_1493 ();
 sg13g2_decap_4 FILLER_25_1505 ();
 sg13g2_decap_8 FILLER_25_1523 ();
 sg13g2_fill_1 FILLER_25_1530 ();
 sg13g2_fill_1 FILLER_25_1557 ();
 sg13g2_decap_8 FILLER_25_1567 ();
 sg13g2_decap_8 FILLER_25_1574 ();
 sg13g2_decap_8 FILLER_25_1581 ();
 sg13g2_decap_4 FILLER_25_1588 ();
 sg13g2_fill_1 FILLER_25_1592 ();
 sg13g2_fill_1 FILLER_25_1598 ();
 sg13g2_fill_2 FILLER_25_1617 ();
 sg13g2_fill_1 FILLER_25_1624 ();
 sg13g2_decap_4 FILLER_25_1643 ();
 sg13g2_fill_1 FILLER_25_1680 ();
 sg13g2_decap_4 FILLER_25_1700 ();
 sg13g2_decap_4 FILLER_25_1709 ();
 sg13g2_fill_2 FILLER_25_1713 ();
 sg13g2_fill_1 FILLER_25_1730 ();
 sg13g2_fill_1 FILLER_25_1740 ();
 sg13g2_fill_2 FILLER_25_1760 ();
 sg13g2_decap_4 FILLER_25_1768 ();
 sg13g2_fill_2 FILLER_25_1772 ();
 sg13g2_fill_2 FILLER_26_31 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_decap_4 FILLER_26_55 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_72 ();
 sg13g2_decap_4 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_127 ();
 sg13g2_fill_2 FILLER_26_157 ();
 sg13g2_fill_2 FILLER_26_163 ();
 sg13g2_decap_8 FILLER_26_173 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_fill_2 FILLER_26_243 ();
 sg13g2_fill_1 FILLER_26_245 ();
 sg13g2_decap_4 FILLER_26_262 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_288 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_decap_4 FILLER_26_302 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_fill_2 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_341 ();
 sg13g2_fill_2 FILLER_26_355 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_fill_1 FILLER_26_397 ();
 sg13g2_fill_1 FILLER_26_423 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_26_440 ();
 sg13g2_decap_4 FILLER_26_498 ();
 sg13g2_fill_1 FILLER_26_507 ();
 sg13g2_fill_1 FILLER_26_520 ();
 sg13g2_fill_1 FILLER_26_530 ();
 sg13g2_fill_2 FILLER_26_546 ();
 sg13g2_fill_1 FILLER_26_554 ();
 sg13g2_fill_2 FILLER_26_565 ();
 sg13g2_fill_1 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_573 ();
 sg13g2_decap_8 FILLER_26_580 ();
 sg13g2_decap_8 FILLER_26_587 ();
 sg13g2_fill_2 FILLER_26_594 ();
 sg13g2_fill_1 FILLER_26_601 ();
 sg13g2_fill_1 FILLER_26_607 ();
 sg13g2_fill_1 FILLER_26_613 ();
 sg13g2_fill_1 FILLER_26_622 ();
 sg13g2_fill_2 FILLER_26_629 ();
 sg13g2_fill_2 FILLER_26_639 ();
 sg13g2_decap_8 FILLER_26_656 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_fill_2 FILLER_26_670 ();
 sg13g2_fill_1 FILLER_26_672 ();
 sg13g2_fill_2 FILLER_26_677 ();
 sg13g2_fill_2 FILLER_26_684 ();
 sg13g2_fill_2 FILLER_26_691 ();
 sg13g2_fill_1 FILLER_26_703 ();
 sg13g2_decap_8 FILLER_26_720 ();
 sg13g2_decap_8 FILLER_26_727 ();
 sg13g2_decap_4 FILLER_26_734 ();
 sg13g2_fill_1 FILLER_26_738 ();
 sg13g2_decap_4 FILLER_26_747 ();
 sg13g2_fill_1 FILLER_26_751 ();
 sg13g2_fill_2 FILLER_26_761 ();
 sg13g2_fill_1 FILLER_26_767 ();
 sg13g2_decap_4 FILLER_26_788 ();
 sg13g2_decap_4 FILLER_26_796 ();
 sg13g2_fill_1 FILLER_26_809 ();
 sg13g2_decap_4 FILLER_26_837 ();
 sg13g2_fill_1 FILLER_26_841 ();
 sg13g2_decap_4 FILLER_26_851 ();
 sg13g2_fill_2 FILLER_26_855 ();
 sg13g2_decap_8 FILLER_26_877 ();
 sg13g2_decap_4 FILLER_26_884 ();
 sg13g2_fill_1 FILLER_26_888 ();
 sg13g2_fill_2 FILLER_26_895 ();
 sg13g2_decap_4 FILLER_26_906 ();
 sg13g2_fill_2 FILLER_26_919 ();
 sg13g2_decap_8 FILLER_26_939 ();
 sg13g2_decap_8 FILLER_26_946 ();
 sg13g2_decap_8 FILLER_26_953 ();
 sg13g2_decap_4 FILLER_26_960 ();
 sg13g2_fill_2 FILLER_26_964 ();
 sg13g2_decap_8 FILLER_26_974 ();
 sg13g2_decap_4 FILLER_26_986 ();
 sg13g2_fill_1 FILLER_26_999 ();
 sg13g2_fill_1 FILLER_26_1004 ();
 sg13g2_decap_8 FILLER_26_1016 ();
 sg13g2_fill_2 FILLER_26_1035 ();
 sg13g2_decap_4 FILLER_26_1046 ();
 sg13g2_fill_1 FILLER_26_1050 ();
 sg13g2_decap_8 FILLER_26_1056 ();
 sg13g2_fill_2 FILLER_26_1063 ();
 sg13g2_fill_2 FILLER_26_1077 ();
 sg13g2_decap_4 FILLER_26_1083 ();
 sg13g2_decap_4 FILLER_26_1100 ();
 sg13g2_fill_1 FILLER_26_1129 ();
 sg13g2_fill_2 FILLER_26_1153 ();
 sg13g2_decap_8 FILLER_26_1166 ();
 sg13g2_decap_4 FILLER_26_1181 ();
 sg13g2_fill_2 FILLER_26_1185 ();
 sg13g2_decap_8 FILLER_26_1191 ();
 sg13g2_decap_8 FILLER_26_1198 ();
 sg13g2_decap_8 FILLER_26_1218 ();
 sg13g2_decap_4 FILLER_26_1225 ();
 sg13g2_decap_4 FILLER_26_1233 ();
 sg13g2_fill_2 FILLER_26_1241 ();
 sg13g2_fill_1 FILLER_26_1243 ();
 sg13g2_decap_4 FILLER_26_1260 ();
 sg13g2_fill_2 FILLER_26_1264 ();
 sg13g2_fill_2 FILLER_26_1271 ();
 sg13g2_fill_1 FILLER_26_1273 ();
 sg13g2_decap_4 FILLER_26_1286 ();
 sg13g2_decap_4 FILLER_26_1298 ();
 sg13g2_fill_2 FILLER_26_1313 ();
 sg13g2_fill_1 FILLER_26_1344 ();
 sg13g2_fill_2 FILLER_26_1365 ();
 sg13g2_fill_2 FILLER_26_1397 ();
 sg13g2_fill_1 FILLER_26_1399 ();
 sg13g2_fill_2 FILLER_26_1406 ();
 sg13g2_decap_4 FILLER_26_1416 ();
 sg13g2_fill_2 FILLER_26_1420 ();
 sg13g2_decap_4 FILLER_26_1427 ();
 sg13g2_fill_1 FILLER_26_1431 ();
 sg13g2_decap_4 FILLER_26_1437 ();
 sg13g2_fill_2 FILLER_26_1441 ();
 sg13g2_decap_8 FILLER_26_1447 ();
 sg13g2_decap_4 FILLER_26_1454 ();
 sg13g2_fill_2 FILLER_26_1458 ();
 sg13g2_decap_4 FILLER_26_1491 ();
 sg13g2_fill_2 FILLER_26_1495 ();
 sg13g2_fill_1 FILLER_26_1501 ();
 sg13g2_decap_8 FILLER_26_1519 ();
 sg13g2_fill_2 FILLER_26_1531 ();
 sg13g2_fill_2 FILLER_26_1556 ();
 sg13g2_fill_1 FILLER_26_1558 ();
 sg13g2_fill_2 FILLER_26_1576 ();
 sg13g2_decap_4 FILLER_26_1586 ();
 sg13g2_fill_1 FILLER_26_1590 ();
 sg13g2_fill_1 FILLER_26_1606 ();
 sg13g2_fill_1 FILLER_26_1617 ();
 sg13g2_fill_2 FILLER_26_1630 ();
 sg13g2_fill_2 FILLER_26_1636 ();
 sg13g2_fill_1 FILLER_26_1641 ();
 sg13g2_fill_1 FILLER_26_1655 ();
 sg13g2_decap_8 FILLER_26_1664 ();
 sg13g2_decap_4 FILLER_26_1680 ();
 sg13g2_fill_2 FILLER_26_1684 ();
 sg13g2_decap_8 FILLER_26_1690 ();
 sg13g2_decap_8 FILLER_26_1697 ();
 sg13g2_decap_8 FILLER_26_1704 ();
 sg13g2_decap_4 FILLER_26_1711 ();
 sg13g2_fill_1 FILLER_26_1715 ();
 sg13g2_fill_2 FILLER_26_1725 ();
 sg13g2_fill_1 FILLER_26_1727 ();
 sg13g2_decap_8 FILLER_26_1733 ();
 sg13g2_fill_2 FILLER_26_1740 ();
 sg13g2_fill_1 FILLER_26_1742 ();
 sg13g2_fill_2 FILLER_26_1751 ();
 sg13g2_decap_4 FILLER_26_1758 ();
 sg13g2_decap_4 FILLER_26_1769 ();
 sg13g2_fill_1 FILLER_26_1773 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_9 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_fill_2 FILLER_27_40 ();
 sg13g2_fill_1 FILLER_27_47 ();
 sg13g2_fill_1 FILLER_27_53 ();
 sg13g2_fill_2 FILLER_27_62 ();
 sg13g2_fill_1 FILLER_27_64 ();
 sg13g2_fill_1 FILLER_27_69 ();
 sg13g2_fill_2 FILLER_27_75 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_103 ();
 sg13g2_fill_2 FILLER_27_113 ();
 sg13g2_fill_1 FILLER_27_115 ();
 sg13g2_fill_1 FILLER_27_139 ();
 sg13g2_fill_2 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_157 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_176 ();
 sg13g2_decap_4 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_fill_1 FILLER_27_218 ();
 sg13g2_fill_2 FILLER_27_227 ();
 sg13g2_decap_8 FILLER_27_241 ();
 sg13g2_decap_4 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_252 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_decap_8 FILLER_27_281 ();
 sg13g2_fill_2 FILLER_27_305 ();
 sg13g2_fill_1 FILLER_27_307 ();
 sg13g2_decap_4 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_fill_2 FILLER_27_378 ();
 sg13g2_fill_1 FILLER_27_433 ();
 sg13g2_fill_2 FILLER_27_438 ();
 sg13g2_decap_8 FILLER_27_445 ();
 sg13g2_fill_1 FILLER_27_452 ();
 sg13g2_fill_2 FILLER_27_457 ();
 sg13g2_fill_1 FILLER_27_459 ();
 sg13g2_fill_1 FILLER_27_473 ();
 sg13g2_decap_8 FILLER_27_478 ();
 sg13g2_decap_4 FILLER_27_485 ();
 sg13g2_fill_2 FILLER_27_489 ();
 sg13g2_fill_1 FILLER_27_500 ();
 sg13g2_fill_1 FILLER_27_532 ();
 sg13g2_fill_2 FILLER_27_544 ();
 sg13g2_fill_1 FILLER_27_551 ();
 sg13g2_fill_1 FILLER_27_561 ();
 sg13g2_fill_1 FILLER_27_566 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_fill_1 FILLER_27_595 ();
 sg13g2_fill_2 FILLER_27_604 ();
 sg13g2_fill_1 FILLER_27_606 ();
 sg13g2_decap_8 FILLER_27_611 ();
 sg13g2_fill_1 FILLER_27_618 ();
 sg13g2_decap_4 FILLER_27_622 ();
 sg13g2_fill_2 FILLER_27_626 ();
 sg13g2_fill_1 FILLER_27_647 ();
 sg13g2_decap_8 FILLER_27_659 ();
 sg13g2_fill_2 FILLER_27_666 ();
 sg13g2_fill_1 FILLER_27_668 ();
 sg13g2_decap_8 FILLER_27_697 ();
 sg13g2_fill_2 FILLER_27_704 ();
 sg13g2_fill_1 FILLER_27_706 ();
 sg13g2_decap_8 FILLER_27_724 ();
 sg13g2_decap_4 FILLER_27_731 ();
 sg13g2_fill_1 FILLER_27_788 ();
 sg13g2_fill_1 FILLER_27_822 ();
 sg13g2_decap_4 FILLER_27_832 ();
 sg13g2_fill_2 FILLER_27_836 ();
 sg13g2_fill_1 FILLER_27_848 ();
 sg13g2_fill_1 FILLER_27_858 ();
 sg13g2_fill_1 FILLER_27_863 ();
 sg13g2_decap_4 FILLER_27_885 ();
 sg13g2_decap_4 FILLER_27_906 ();
 sg13g2_fill_1 FILLER_27_910 ();
 sg13g2_fill_1 FILLER_27_930 ();
 sg13g2_fill_1 FILLER_27_937 ();
 sg13g2_fill_1 FILLER_27_944 ();
 sg13g2_decap_8 FILLER_27_953 ();
 sg13g2_fill_1 FILLER_27_960 ();
 sg13g2_decap_8 FILLER_27_969 ();
 sg13g2_fill_2 FILLER_27_976 ();
 sg13g2_fill_2 FILLER_27_982 ();
 sg13g2_fill_2 FILLER_27_988 ();
 sg13g2_fill_2 FILLER_27_995 ();
 sg13g2_decap_4 FILLER_27_1006 ();
 sg13g2_fill_1 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_fill_1 FILLER_27_1024 ();
 sg13g2_fill_1 FILLER_27_1034 ();
 sg13g2_decap_4 FILLER_27_1040 ();
 sg13g2_fill_1 FILLER_27_1044 ();
 sg13g2_fill_2 FILLER_27_1049 ();
 sg13g2_decap_8 FILLER_27_1055 ();
 sg13g2_fill_1 FILLER_27_1062 ();
 sg13g2_fill_1 FILLER_27_1071 ();
 sg13g2_decap_4 FILLER_27_1077 ();
 sg13g2_decap_4 FILLER_27_1090 ();
 sg13g2_decap_8 FILLER_27_1102 ();
 sg13g2_decap_8 FILLER_27_1109 ();
 sg13g2_fill_2 FILLER_27_1116 ();
 sg13g2_decap_8 FILLER_27_1122 ();
 sg13g2_decap_8 FILLER_27_1129 ();
 sg13g2_fill_1 FILLER_27_1136 ();
 sg13g2_decap_4 FILLER_27_1158 ();
 sg13g2_fill_1 FILLER_27_1162 ();
 sg13g2_decap_4 FILLER_27_1171 ();
 sg13g2_decap_8 FILLER_27_1184 ();
 sg13g2_decap_4 FILLER_27_1191 ();
 sg13g2_decap_8 FILLER_27_1220 ();
 sg13g2_fill_1 FILLER_27_1227 ();
 sg13g2_decap_4 FILLER_27_1232 ();
 sg13g2_decap_4 FILLER_27_1248 ();
 sg13g2_decap_4 FILLER_27_1263 ();
 sg13g2_fill_2 FILLER_27_1267 ();
 sg13g2_decap_8 FILLER_27_1282 ();
 sg13g2_decap_8 FILLER_27_1289 ();
 sg13g2_fill_1 FILLER_27_1296 ();
 sg13g2_fill_2 FILLER_27_1310 ();
 sg13g2_fill_1 FILLER_27_1315 ();
 sg13g2_fill_2 FILLER_27_1323 ();
 sg13g2_fill_2 FILLER_27_1380 ();
 sg13g2_decap_4 FILLER_27_1432 ();
 sg13g2_fill_1 FILLER_27_1471 ();
 sg13g2_fill_1 FILLER_27_1484 ();
 sg13g2_fill_1 FILLER_27_1493 ();
 sg13g2_fill_2 FILLER_27_1499 ();
 sg13g2_fill_1 FILLER_27_1501 ();
 sg13g2_fill_1 FILLER_27_1507 ();
 sg13g2_fill_1 FILLER_27_1511 ();
 sg13g2_decap_4 FILLER_27_1515 ();
 sg13g2_fill_1 FILLER_27_1519 ();
 sg13g2_fill_1 FILLER_27_1525 ();
 sg13g2_fill_2 FILLER_27_1530 ();
 sg13g2_fill_1 FILLER_27_1532 ();
 sg13g2_fill_2 FILLER_27_1559 ();
 sg13g2_decap_4 FILLER_27_1565 ();
 sg13g2_decap_8 FILLER_27_1573 ();
 sg13g2_decap_8 FILLER_27_1580 ();
 sg13g2_decap_4 FILLER_27_1587 ();
 sg13g2_decap_4 FILLER_27_1601 ();
 sg13g2_fill_2 FILLER_27_1610 ();
 sg13g2_fill_2 FILLER_27_1620 ();
 sg13g2_fill_2 FILLER_27_1627 ();
 sg13g2_decap_4 FILLER_27_1634 ();
 sg13g2_fill_1 FILLER_27_1638 ();
 sg13g2_decap_8 FILLER_27_1643 ();
 sg13g2_fill_1 FILLER_27_1655 ();
 sg13g2_fill_1 FILLER_27_1664 ();
 sg13g2_fill_1 FILLER_27_1673 ();
 sg13g2_decap_8 FILLER_27_1678 ();
 sg13g2_decap_4 FILLER_27_1685 ();
 sg13g2_decap_8 FILLER_27_1701 ();
 sg13g2_fill_2 FILLER_27_1708 ();
 sg13g2_fill_2 FILLER_27_1738 ();
 sg13g2_decap_4 FILLER_27_1753 ();
 sg13g2_fill_1 FILLER_27_1762 ();
 sg13g2_decap_4 FILLER_27_1768 ();
 sg13g2_fill_2 FILLER_27_1772 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_26 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_58 ();
 sg13g2_fill_1 FILLER_28_64 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_95 ();
 sg13g2_fill_1 FILLER_28_97 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_118 ();
 sg13g2_decap_4 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_165 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_decap_4 FILLER_28_183 ();
 sg13g2_fill_2 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_4 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_252 ();
 sg13g2_fill_1 FILLER_28_254 ();
 sg13g2_decap_4 FILLER_28_263 ();
 sg13g2_fill_2 FILLER_28_292 ();
 sg13g2_fill_2 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_318 ();
 sg13g2_fill_1 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_348 ();
 sg13g2_decap_4 FILLER_28_408 ();
 sg13g2_fill_1 FILLER_28_412 ();
 sg13g2_fill_2 FILLER_28_431 ();
 sg13g2_fill_1 FILLER_28_437 ();
 sg13g2_fill_2 FILLER_28_457 ();
 sg13g2_fill_1 FILLER_28_459 ();
 sg13g2_fill_2 FILLER_28_463 ();
 sg13g2_fill_2 FILLER_28_521 ();
 sg13g2_fill_1 FILLER_28_523 ();
 sg13g2_fill_2 FILLER_28_527 ();
 sg13g2_fill_1 FILLER_28_529 ();
 sg13g2_fill_1 FILLER_28_549 ();
 sg13g2_fill_2 FILLER_28_555 ();
 sg13g2_decap_8 FILLER_28_562 ();
 sg13g2_decap_8 FILLER_28_569 ();
 sg13g2_decap_8 FILLER_28_576 ();
 sg13g2_fill_1 FILLER_28_583 ();
 sg13g2_fill_1 FILLER_28_592 ();
 sg13g2_fill_2 FILLER_28_617 ();
 sg13g2_fill_1 FILLER_28_619 ();
 sg13g2_decap_8 FILLER_28_661 ();
 sg13g2_decap_8 FILLER_28_668 ();
 sg13g2_decap_4 FILLER_28_675 ();
 sg13g2_fill_1 FILLER_28_679 ();
 sg13g2_decap_4 FILLER_28_684 ();
 sg13g2_fill_2 FILLER_28_688 ();
 sg13g2_decap_8 FILLER_28_699 ();
 sg13g2_fill_1 FILLER_28_718 ();
 sg13g2_fill_2 FILLER_28_724 ();
 sg13g2_fill_1 FILLER_28_726 ();
 sg13g2_fill_2 FILLER_28_740 ();
 sg13g2_fill_1 FILLER_28_742 ();
 sg13g2_fill_1 FILLER_28_784 ();
 sg13g2_fill_1 FILLER_28_792 ();
 sg13g2_fill_1 FILLER_28_798 ();
 sg13g2_fill_1 FILLER_28_810 ();
 sg13g2_fill_2 FILLER_28_822 ();
 sg13g2_fill_1 FILLER_28_824 ();
 sg13g2_decap_8 FILLER_28_834 ();
 sg13g2_decap_8 FILLER_28_841 ();
 sg13g2_decap_8 FILLER_28_848 ();
 sg13g2_decap_4 FILLER_28_855 ();
 sg13g2_fill_1 FILLER_28_872 ();
 sg13g2_fill_1 FILLER_28_881 ();
 sg13g2_fill_1 FILLER_28_885 ();
 sg13g2_decap_4 FILLER_28_910 ();
 sg13g2_fill_2 FILLER_28_914 ();
 sg13g2_decap_8 FILLER_28_932 ();
 sg13g2_decap_4 FILLER_28_939 ();
 sg13g2_fill_2 FILLER_28_943 ();
 sg13g2_fill_2 FILLER_28_953 ();
 sg13g2_fill_1 FILLER_28_955 ();
 sg13g2_decap_8 FILLER_28_998 ();
 sg13g2_decap_4 FILLER_28_1005 ();
 sg13g2_fill_1 FILLER_28_1009 ();
 sg13g2_decap_8 FILLER_28_1018 ();
 sg13g2_decap_8 FILLER_28_1033 ();
 sg13g2_decap_8 FILLER_28_1040 ();
 sg13g2_fill_1 FILLER_28_1047 ();
 sg13g2_decap_4 FILLER_28_1064 ();
 sg13g2_fill_1 FILLER_28_1093 ();
 sg13g2_fill_2 FILLER_28_1129 ();
 sg13g2_fill_1 FILLER_28_1131 ();
 sg13g2_fill_1 FILLER_28_1157 ();
 sg13g2_decap_4 FILLER_28_1171 ();
 sg13g2_fill_2 FILLER_28_1188 ();
 sg13g2_fill_1 FILLER_28_1190 ();
 sg13g2_decap_8 FILLER_28_1201 ();
 sg13g2_decap_8 FILLER_28_1208 ();
 sg13g2_decap_8 FILLER_28_1215 ();
 sg13g2_decap_4 FILLER_28_1230 ();
 sg13g2_fill_2 FILLER_28_1234 ();
 sg13g2_fill_2 FILLER_28_1244 ();
 sg13g2_fill_1 FILLER_28_1256 ();
 sg13g2_decap_8 FILLER_28_1260 ();
 sg13g2_decap_8 FILLER_28_1267 ();
 sg13g2_fill_2 FILLER_28_1274 ();
 sg13g2_fill_2 FILLER_28_1280 ();
 sg13g2_fill_1 FILLER_28_1303 ();
 sg13g2_fill_2 FILLER_28_1312 ();
 sg13g2_fill_1 FILLER_28_1385 ();
 sg13g2_decap_8 FILLER_28_1432 ();
 sg13g2_decap_8 FILLER_28_1439 ();
 sg13g2_decap_8 FILLER_28_1446 ();
 sg13g2_fill_1 FILLER_28_1457 ();
 sg13g2_fill_2 FILLER_28_1463 ();
 sg13g2_fill_1 FILLER_28_1468 ();
 sg13g2_fill_2 FILLER_28_1477 ();
 sg13g2_fill_2 FILLER_28_1493 ();
 sg13g2_fill_2 FILLER_28_1500 ();
 sg13g2_decap_8 FILLER_28_1510 ();
 sg13g2_fill_1 FILLER_28_1517 ();
 sg13g2_fill_1 FILLER_28_1524 ();
 sg13g2_fill_2 FILLER_28_1532 ();
 sg13g2_fill_1 FILLER_28_1545 ();
 sg13g2_decap_4 FILLER_28_1570 ();
 sg13g2_fill_1 FILLER_28_1574 ();
 sg13g2_decap_4 FILLER_28_1585 ();
 sg13g2_fill_1 FILLER_28_1589 ();
 sg13g2_fill_2 FILLER_28_1595 ();
 sg13g2_decap_8 FILLER_28_1610 ();
 sg13g2_decap_8 FILLER_28_1617 ();
 sg13g2_fill_2 FILLER_28_1624 ();
 sg13g2_fill_1 FILLER_28_1630 ();
 sg13g2_decap_8 FILLER_28_1636 ();
 sg13g2_fill_2 FILLER_28_1643 ();
 sg13g2_fill_1 FILLER_28_1645 ();
 sg13g2_fill_2 FILLER_28_1654 ();
 sg13g2_fill_1 FILLER_28_1656 ();
 sg13g2_decap_4 FILLER_28_1665 ();
 sg13g2_decap_4 FILLER_28_1674 ();
 sg13g2_fill_1 FILLER_28_1678 ();
 sg13g2_decap_4 FILLER_28_1709 ();
 sg13g2_fill_2 FILLER_28_1713 ();
 sg13g2_fill_1 FILLER_28_1718 ();
 sg13g2_fill_1 FILLER_28_1724 ();
 sg13g2_fill_1 FILLER_28_1736 ();
 sg13g2_fill_1 FILLER_28_1742 ();
 sg13g2_fill_1 FILLER_28_1748 ();
 sg13g2_fill_1 FILLER_28_1754 ();
 sg13g2_decap_8 FILLER_28_1765 ();
 sg13g2_fill_2 FILLER_28_1772 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_19 ();
 sg13g2_decap_8 FILLER_29_34 ();
 sg13g2_decap_8 FILLER_29_41 ();
 sg13g2_fill_2 FILLER_29_52 ();
 sg13g2_decap_4 FILLER_29_64 ();
 sg13g2_decap_8 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_decap_8 FILLER_29_101 ();
 sg13g2_fill_2 FILLER_29_108 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_decap_4 FILLER_29_117 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_207 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_240 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_fill_2 FILLER_29_260 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_2 FILLER_29_281 ();
 sg13g2_fill_1 FILLER_29_288 ();
 sg13g2_fill_2 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_311 ();
 sg13g2_decap_4 FILLER_29_318 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_fill_2 FILLER_29_344 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_fill_2 FILLER_29_356 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_decap_4 FILLER_29_364 ();
 sg13g2_fill_1 FILLER_29_368 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_1 FILLER_29_402 ();
 sg13g2_fill_2 FILLER_29_412 ();
 sg13g2_fill_1 FILLER_29_420 ();
 sg13g2_decap_4 FILLER_29_433 ();
 sg13g2_fill_1 FILLER_29_437 ();
 sg13g2_decap_4 FILLER_29_447 ();
 sg13g2_fill_1 FILLER_29_451 ();
 sg13g2_decap_8 FILLER_29_481 ();
 sg13g2_decap_8 FILLER_29_488 ();
 sg13g2_decap_8 FILLER_29_499 ();
 sg13g2_fill_2 FILLER_29_506 ();
 sg13g2_fill_1 FILLER_29_517 ();
 sg13g2_fill_2 FILLER_29_535 ();
 sg13g2_decap_4 FILLER_29_561 ();
 sg13g2_fill_2 FILLER_29_565 ();
 sg13g2_decap_8 FILLER_29_571 ();
 sg13g2_decap_8 FILLER_29_578 ();
 sg13g2_decap_8 FILLER_29_585 ();
 sg13g2_fill_1 FILLER_29_596 ();
 sg13g2_decap_8 FILLER_29_601 ();
 sg13g2_decap_4 FILLER_29_608 ();
 sg13g2_decap_4 FILLER_29_673 ();
 sg13g2_fill_2 FILLER_29_718 ();
 sg13g2_fill_1 FILLER_29_720 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_4 FILLER_29_749 ();
 sg13g2_fill_1 FILLER_29_753 ();
 sg13g2_decap_8 FILLER_29_759 ();
 sg13g2_decap_4 FILLER_29_766 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_decap_4 FILLER_29_788 ();
 sg13g2_fill_1 FILLER_29_797 ();
 sg13g2_fill_1 FILLER_29_804 ();
 sg13g2_fill_2 FILLER_29_810 ();
 sg13g2_fill_1 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_817 ();
 sg13g2_decap_8 FILLER_29_829 ();
 sg13g2_fill_2 FILLER_29_836 ();
 sg13g2_fill_1 FILLER_29_838 ();
 sg13g2_fill_1 FILLER_29_886 ();
 sg13g2_decap_8 FILLER_29_895 ();
 sg13g2_decap_4 FILLER_29_902 ();
 sg13g2_fill_1 FILLER_29_906 ();
 sg13g2_decap_4 FILLER_29_917 ();
 sg13g2_fill_1 FILLER_29_921 ();
 sg13g2_decap_8 FILLER_29_932 ();
 sg13g2_decap_8 FILLER_29_939 ();
 sg13g2_decap_8 FILLER_29_946 ();
 sg13g2_fill_1 FILLER_29_953 ();
 sg13g2_decap_8 FILLER_29_958 ();
 sg13g2_decap_4 FILLER_29_991 ();
 sg13g2_fill_2 FILLER_29_1010 ();
 sg13g2_fill_1 FILLER_29_1017 ();
 sg13g2_decap_8 FILLER_29_1054 ();
 sg13g2_fill_2 FILLER_29_1061 ();
 sg13g2_fill_1 FILLER_29_1063 ();
 sg13g2_decap_8 FILLER_29_1085 ();
 sg13g2_decap_4 FILLER_29_1092 ();
 sg13g2_fill_1 FILLER_29_1096 ();
 sg13g2_fill_2 FILLER_29_1105 ();
 sg13g2_decap_8 FILLER_29_1115 ();
 sg13g2_decap_4 FILLER_29_1122 ();
 sg13g2_fill_1 FILLER_29_1139 ();
 sg13g2_fill_1 FILLER_29_1150 ();
 sg13g2_decap_4 FILLER_29_1164 ();
 sg13g2_fill_2 FILLER_29_1181 ();
 sg13g2_fill_1 FILLER_29_1183 ();
 sg13g2_decap_8 FILLER_29_1215 ();
 sg13g2_decap_4 FILLER_29_1222 ();
 sg13g2_fill_2 FILLER_29_1226 ();
 sg13g2_decap_4 FILLER_29_1236 ();
 sg13g2_fill_2 FILLER_29_1264 ();
 sg13g2_fill_1 FILLER_29_1266 ();
 sg13g2_decap_8 FILLER_29_1287 ();
 sg13g2_decap_8 FILLER_29_1298 ();
 sg13g2_fill_2 FILLER_29_1305 ();
 sg13g2_fill_2 FILLER_29_1323 ();
 sg13g2_fill_1 FILLER_29_1360 ();
 sg13g2_decap_8 FILLER_29_1369 ();
 sg13g2_fill_2 FILLER_29_1376 ();
 sg13g2_fill_1 FILLER_29_1378 ();
 sg13g2_fill_2 FILLER_29_1417 ();
 sg13g2_fill_2 FILLER_29_1439 ();
 sg13g2_fill_2 FILLER_29_1445 ();
 sg13g2_fill_1 FILLER_29_1453 ();
 sg13g2_fill_1 FILLER_29_1473 ();
 sg13g2_decap_4 FILLER_29_1491 ();
 sg13g2_fill_2 FILLER_29_1495 ();
 sg13g2_fill_2 FILLER_29_1517 ();
 sg13g2_fill_1 FILLER_29_1519 ();
 sg13g2_fill_1 FILLER_29_1533 ();
 sg13g2_fill_2 FILLER_29_1592 ();
 sg13g2_fill_1 FILLER_29_1594 ();
 sg13g2_decap_4 FILLER_29_1608 ();
 sg13g2_fill_2 FILLER_29_1612 ();
 sg13g2_fill_1 FILLER_29_1620 ();
 sg13g2_fill_1 FILLER_29_1626 ();
 sg13g2_decap_8 FILLER_29_1639 ();
 sg13g2_decap_4 FILLER_29_1646 ();
 sg13g2_fill_2 FILLER_29_1650 ();
 sg13g2_decap_8 FILLER_29_1657 ();
 sg13g2_decap_8 FILLER_29_1664 ();
 sg13g2_decap_8 FILLER_29_1678 ();
 sg13g2_decap_4 FILLER_29_1685 ();
 sg13g2_fill_1 FILLER_29_1718 ();
 sg13g2_fill_1 FILLER_29_1724 ();
 sg13g2_fill_1 FILLER_29_1730 ();
 sg13g2_fill_1 FILLER_29_1736 ();
 sg13g2_fill_1 FILLER_29_1741 ();
 sg13g2_fill_1 FILLER_29_1747 ();
 sg13g2_fill_1 FILLER_29_1756 ();
 sg13g2_decap_8 FILLER_29_1764 ();
 sg13g2_fill_2 FILLER_29_1771 ();
 sg13g2_fill_1 FILLER_29_1773 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_24 ();
 sg13g2_fill_1 FILLER_30_39 ();
 sg13g2_fill_1 FILLER_30_48 ();
 sg13g2_decap_8 FILLER_30_75 ();
 sg13g2_decap_8 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_89 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_114 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_129 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_4 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_decap_4 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_fill_2 FILLER_30_255 ();
 sg13g2_fill_1 FILLER_30_257 ();
 sg13g2_decap_4 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_299 ();
 sg13g2_decap_8 FILLER_30_310 ();
 sg13g2_decap_8 FILLER_30_317 ();
 sg13g2_decap_4 FILLER_30_324 ();
 sg13g2_decap_4 FILLER_30_332 ();
 sg13g2_fill_1 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_fill_1 FILLER_30_349 ();
 sg13g2_fill_2 FILLER_30_366 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_30_423 ();
 sg13g2_decap_4 FILLER_30_439 ();
 sg13g2_fill_2 FILLER_30_443 ();
 sg13g2_fill_1 FILLER_30_449 ();
 sg13g2_fill_2 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_4 FILLER_30_490 ();
 sg13g2_fill_2 FILLER_30_494 ();
 sg13g2_decap_4 FILLER_30_502 ();
 sg13g2_fill_2 FILLER_30_506 ();
 sg13g2_decap_4 FILLER_30_517 ();
 sg13g2_fill_1 FILLER_30_521 ();
 sg13g2_decap_8 FILLER_30_530 ();
 sg13g2_decap_4 FILLER_30_537 ();
 sg13g2_fill_2 FILLER_30_548 ();
 sg13g2_fill_1 FILLER_30_560 ();
 sg13g2_decap_4 FILLER_30_569 ();
 sg13g2_decap_4 FILLER_30_581 ();
 sg13g2_decap_4 FILLER_30_590 ();
 sg13g2_fill_2 FILLER_30_599 ();
 sg13g2_decap_4 FILLER_30_611 ();
 sg13g2_fill_1 FILLER_30_615 ();
 sg13g2_fill_2 FILLER_30_647 ();
 sg13g2_fill_1 FILLER_30_649 ();
 sg13g2_decap_4 FILLER_30_654 ();
 sg13g2_decap_4 FILLER_30_662 ();
 sg13g2_fill_1 FILLER_30_666 ();
 sg13g2_fill_2 FILLER_30_693 ();
 sg13g2_decap_4 FILLER_30_703 ();
 sg13g2_fill_1 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_717 ();
 sg13g2_decap_8 FILLER_30_737 ();
 sg13g2_decap_8 FILLER_30_744 ();
 sg13g2_decap_8 FILLER_30_751 ();
 sg13g2_decap_4 FILLER_30_758 ();
 sg13g2_fill_2 FILLER_30_762 ();
 sg13g2_decap_8 FILLER_30_778 ();
 sg13g2_fill_1 FILLER_30_799 ();
 sg13g2_fill_1 FILLER_30_805 ();
 sg13g2_fill_1 FILLER_30_814 ();
 sg13g2_fill_1 FILLER_30_819 ();
 sg13g2_fill_2 FILLER_30_824 ();
 sg13g2_decap_4 FILLER_30_831 ();
 sg13g2_decap_4 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_848 ();
 sg13g2_decap_8 FILLER_30_855 ();
 sg13g2_decap_4 FILLER_30_862 ();
 sg13g2_fill_2 FILLER_30_877 ();
 sg13g2_fill_1 FILLER_30_890 ();
 sg13g2_decap_4 FILLER_30_907 ();
 sg13g2_fill_2 FILLER_30_916 ();
 sg13g2_fill_2 FILLER_30_923 ();
 sg13g2_fill_1 FILLER_30_925 ();
 sg13g2_decap_4 FILLER_30_934 ();
 sg13g2_fill_1 FILLER_30_942 ();
 sg13g2_decap_8 FILLER_30_959 ();
 sg13g2_decap_8 FILLER_30_966 ();
 sg13g2_decap_8 FILLER_30_973 ();
 sg13g2_decap_4 FILLER_30_980 ();
 sg13g2_fill_1 FILLER_30_984 ();
 sg13g2_fill_2 FILLER_30_989 ();
 sg13g2_fill_1 FILLER_30_991 ();
 sg13g2_decap_8 FILLER_30_996 ();
 sg13g2_decap_8 FILLER_30_1013 ();
 sg13g2_decap_4 FILLER_30_1020 ();
 sg13g2_fill_2 FILLER_30_1024 ();
 sg13g2_decap_4 FILLER_30_1030 ();
 sg13g2_fill_1 FILLER_30_1034 ();
 sg13g2_fill_2 FILLER_30_1039 ();
 sg13g2_fill_1 FILLER_30_1041 ();
 sg13g2_decap_4 FILLER_30_1046 ();
 sg13g2_fill_1 FILLER_30_1054 ();
 sg13g2_decap_4 FILLER_30_1059 ();
 sg13g2_decap_8 FILLER_30_1074 ();
 sg13g2_decap_8 FILLER_30_1081 ();
 sg13g2_decap_4 FILLER_30_1098 ();
 sg13g2_fill_1 FILLER_30_1102 ();
 sg13g2_decap_4 FILLER_30_1108 ();
 sg13g2_fill_2 FILLER_30_1112 ();
 sg13g2_fill_1 FILLER_30_1140 ();
 sg13g2_fill_1 FILLER_30_1146 ();
 sg13g2_decap_8 FILLER_30_1156 ();
 sg13g2_decap_4 FILLER_30_1163 ();
 sg13g2_fill_2 FILLER_30_1172 ();
 sg13g2_fill_1 FILLER_30_1174 ();
 sg13g2_fill_1 FILLER_30_1183 ();
 sg13g2_decap_4 FILLER_30_1192 ();
 sg13g2_decap_8 FILLER_30_1200 ();
 sg13g2_decap_8 FILLER_30_1207 ();
 sg13g2_decap_8 FILLER_30_1214 ();
 sg13g2_fill_1 FILLER_30_1221 ();
 sg13g2_fill_1 FILLER_30_1234 ();
 sg13g2_fill_2 FILLER_30_1257 ();
 sg13g2_decap_8 FILLER_30_1264 ();
 sg13g2_fill_2 FILLER_30_1271 ();
 sg13g2_decap_8 FILLER_30_1277 ();
 sg13g2_fill_2 FILLER_30_1284 ();
 sg13g2_fill_2 FILLER_30_1306 ();
 sg13g2_fill_1 FILLER_30_1308 ();
 sg13g2_fill_1 FILLER_30_1317 ();
 sg13g2_fill_1 FILLER_30_1337 ();
 sg13g2_fill_1 FILLER_30_1342 ();
 sg13g2_fill_2 FILLER_30_1361 ();
 sg13g2_decap_8 FILLER_30_1374 ();
 sg13g2_decap_8 FILLER_30_1381 ();
 sg13g2_fill_1 FILLER_30_1388 ();
 sg13g2_decap_4 FILLER_30_1405 ();
 sg13g2_fill_1 FILLER_30_1409 ();
 sg13g2_decap_4 FILLER_30_1415 ();
 sg13g2_decap_4 FILLER_30_1433 ();
 sg13g2_fill_2 FILLER_30_1437 ();
 sg13g2_fill_2 FILLER_30_1444 ();
 sg13g2_fill_1 FILLER_30_1446 ();
 sg13g2_fill_2 FILLER_30_1455 ();
 sg13g2_fill_1 FILLER_30_1457 ();
 sg13g2_fill_1 FILLER_30_1474 ();
 sg13g2_decap_8 FILLER_30_1479 ();
 sg13g2_decap_8 FILLER_30_1486 ();
 sg13g2_decap_4 FILLER_30_1498 ();
 sg13g2_fill_1 FILLER_30_1518 ();
 sg13g2_fill_1 FILLER_30_1532 ();
 sg13g2_fill_1 FILLER_30_1537 ();
 sg13g2_decap_4 FILLER_30_1543 ();
 sg13g2_decap_8 FILLER_30_1553 ();
 sg13g2_decap_4 FILLER_30_1560 ();
 sg13g2_fill_2 FILLER_30_1564 ();
 sg13g2_decap_8 FILLER_30_1574 ();
 sg13g2_decap_4 FILLER_30_1581 ();
 sg13g2_fill_2 FILLER_30_1585 ();
 sg13g2_fill_2 FILLER_30_1615 ();
 sg13g2_fill_1 FILLER_30_1617 ();
 sg13g2_fill_2 FILLER_30_1642 ();
 sg13g2_fill_1 FILLER_30_1652 ();
 sg13g2_fill_1 FILLER_30_1708 ();
 sg13g2_decap_8 FILLER_30_1728 ();
 sg13g2_fill_1 FILLER_30_1735 ();
 sg13g2_fill_2 FILLER_30_1739 ();
 sg13g2_fill_1 FILLER_30_1741 ();
 sg13g2_fill_1 FILLER_30_1747 ();
 sg13g2_decap_8 FILLER_30_1760 ();
 sg13g2_decap_8 FILLER_30_1767 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_30 ();
 sg13g2_decap_4 FILLER_31_37 ();
 sg13g2_fill_2 FILLER_31_44 ();
 sg13g2_decap_4 FILLER_31_54 ();
 sg13g2_decap_8 FILLER_31_62 ();
 sg13g2_decap_4 FILLER_31_69 ();
 sg13g2_decap_4 FILLER_31_83 ();
 sg13g2_fill_2 FILLER_31_87 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_125 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_decap_4 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_decap_4 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_decap_8 FILLER_31_255 ();
 sg13g2_fill_2 FILLER_31_267 ();
 sg13g2_decap_4 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_335 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_354 ();
 sg13g2_fill_1 FILLER_31_383 ();
 sg13g2_fill_2 FILLER_31_397 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_fill_1 FILLER_31_414 ();
 sg13g2_fill_2 FILLER_31_435 ();
 sg13g2_fill_1 FILLER_31_463 ();
 sg13g2_decap_8 FILLER_31_471 ();
 sg13g2_fill_2 FILLER_31_478 ();
 sg13g2_fill_2 FILLER_31_485 ();
 sg13g2_fill_2 FILLER_31_493 ();
 sg13g2_fill_1 FILLER_31_495 ();
 sg13g2_fill_1 FILLER_31_516 ();
 sg13g2_fill_1 FILLER_31_544 ();
 sg13g2_fill_1 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_568 ();
 sg13g2_decap_4 FILLER_31_575 ();
 sg13g2_fill_1 FILLER_31_579 ();
 sg13g2_fill_1 FILLER_31_585 ();
 sg13g2_decap_4 FILLER_31_606 ();
 sg13g2_fill_1 FILLER_31_610 ();
 sg13g2_fill_1 FILLER_31_687 ();
 sg13g2_fill_1 FILLER_31_693 ();
 sg13g2_fill_1 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_720 ();
 sg13g2_decap_8 FILLER_31_731 ();
 sg13g2_decap_4 FILLER_31_738 ();
 sg13g2_fill_2 FILLER_31_742 ();
 sg13g2_fill_1 FILLER_31_771 ();
 sg13g2_fill_2 FILLER_31_784 ();
 sg13g2_fill_1 FILLER_31_786 ();
 sg13g2_fill_1 FILLER_31_790 ();
 sg13g2_decap_4 FILLER_31_808 ();
 sg13g2_fill_1 FILLER_31_827 ();
 sg13g2_fill_1 FILLER_31_832 ();
 sg13g2_fill_1 FILLER_31_838 ();
 sg13g2_fill_1 FILLER_31_843 ();
 sg13g2_fill_2 FILLER_31_849 ();
 sg13g2_fill_1 FILLER_31_851 ();
 sg13g2_decap_8 FILLER_31_857 ();
 sg13g2_decap_4 FILLER_31_864 ();
 sg13g2_fill_1 FILLER_31_868 ();
 sg13g2_decap_8 FILLER_31_875 ();
 sg13g2_decap_4 FILLER_31_882 ();
 sg13g2_fill_2 FILLER_31_891 ();
 sg13g2_fill_1 FILLER_31_893 ();
 sg13g2_decap_4 FILLER_31_902 ();
 sg13g2_fill_1 FILLER_31_906 ();
 sg13g2_decap_4 FILLER_31_919 ();
 sg13g2_decap_4 FILLER_31_927 ();
 sg13g2_decap_8 FILLER_31_935 ();
 sg13g2_decap_4 FILLER_31_942 ();
 sg13g2_fill_1 FILLER_31_950 ();
 sg13g2_decap_4 FILLER_31_967 ();
 sg13g2_fill_1 FILLER_31_987 ();
 sg13g2_decap_4 FILLER_31_999 ();
 sg13g2_fill_1 FILLER_31_1029 ();
 sg13g2_decap_8 FILLER_31_1034 ();
 sg13g2_fill_2 FILLER_31_1041 ();
 sg13g2_fill_1 FILLER_31_1047 ();
 sg13g2_fill_1 FILLER_31_1057 ();
 sg13g2_decap_8 FILLER_31_1068 ();
 sg13g2_fill_1 FILLER_31_1075 ();
 sg13g2_fill_2 FILLER_31_1103 ();
 sg13g2_fill_1 FILLER_31_1105 ();
 sg13g2_decap_8 FILLER_31_1111 ();
 sg13g2_decap_8 FILLER_31_1118 ();
 sg13g2_fill_2 FILLER_31_1125 ();
 sg13g2_decap_8 FILLER_31_1131 ();
 sg13g2_fill_2 FILLER_31_1156 ();
 sg13g2_fill_1 FILLER_31_1158 ();
 sg13g2_decap_8 FILLER_31_1207 ();
 sg13g2_decap_4 FILLER_31_1214 ();
 sg13g2_fill_1 FILLER_31_1239 ();
 sg13g2_fill_1 FILLER_31_1245 ();
 sg13g2_fill_1 FILLER_31_1252 ();
 sg13g2_decap_4 FILLER_31_1266 ();
 sg13g2_fill_1 FILLER_31_1270 ();
 sg13g2_decap_8 FILLER_31_1276 ();
 sg13g2_decap_4 FILLER_31_1283 ();
 sg13g2_fill_1 FILLER_31_1287 ();
 sg13g2_fill_1 FILLER_31_1296 ();
 sg13g2_decap_4 FILLER_31_1325 ();
 sg13g2_fill_1 FILLER_31_1329 ();
 sg13g2_fill_1 FILLER_31_1342 ();
 sg13g2_fill_1 FILLER_31_1362 ();
 sg13g2_fill_1 FILLER_31_1371 ();
 sg13g2_decap_4 FILLER_31_1377 ();
 sg13g2_fill_1 FILLER_31_1381 ();
 sg13g2_decap_8 FILLER_31_1387 ();
 sg13g2_decap_4 FILLER_31_1394 ();
 sg13g2_fill_2 FILLER_31_1406 ();
 sg13g2_fill_1 FILLER_31_1408 ();
 sg13g2_decap_8 FILLER_31_1420 ();
 sg13g2_fill_1 FILLER_31_1427 ();
 sg13g2_fill_2 FILLER_31_1442 ();
 sg13g2_decap_4 FILLER_31_1449 ();
 sg13g2_fill_2 FILLER_31_1453 ();
 sg13g2_fill_2 FILLER_31_1470 ();
 sg13g2_decap_8 FILLER_31_1477 ();
 sg13g2_decap_8 FILLER_31_1484 ();
 sg13g2_fill_1 FILLER_31_1491 ();
 sg13g2_decap_8 FILLER_31_1516 ();
 sg13g2_fill_2 FILLER_31_1523 ();
 sg13g2_decap_8 FILLER_31_1530 ();
 sg13g2_fill_1 FILLER_31_1537 ();
 sg13g2_decap_8 FILLER_31_1548 ();
 sg13g2_decap_8 FILLER_31_1555 ();
 sg13g2_fill_2 FILLER_31_1562 ();
 sg13g2_decap_8 FILLER_31_1572 ();
 sg13g2_decap_8 FILLER_31_1579 ();
 sg13g2_fill_2 FILLER_31_1586 ();
 sg13g2_fill_2 FILLER_31_1598 ();
 sg13g2_decap_8 FILLER_31_1613 ();
 sg13g2_decap_4 FILLER_31_1620 ();
 sg13g2_fill_2 FILLER_31_1628 ();
 sg13g2_fill_2 FILLER_31_1648 ();
 sg13g2_fill_2 FILLER_31_1655 ();
 sg13g2_fill_1 FILLER_31_1675 ();
 sg13g2_fill_2 FILLER_31_1689 ();
 sg13g2_fill_1 FILLER_31_1691 ();
 sg13g2_fill_1 FILLER_31_1726 ();
 sg13g2_fill_1 FILLER_31_1761 ();
 sg13g2_decap_8 FILLER_31_1767 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_27 ();
 sg13g2_decap_4 FILLER_32_59 ();
 sg13g2_decap_4 FILLER_32_71 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_decap_4 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_96 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_122 ();
 sg13g2_fill_1 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_decap_4 FILLER_32_162 ();
 sg13g2_decap_8 FILLER_32_184 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_fill_2 FILLER_32_202 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_decap_8 FILLER_32_236 ();
 sg13g2_fill_2 FILLER_32_243 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_1 FILLER_32_283 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_331 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_382 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_394 ();
 sg13g2_decap_4 FILLER_32_398 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_1 FILLER_32_409 ();
 sg13g2_fill_2 FILLER_32_414 ();
 sg13g2_fill_1 FILLER_32_420 ();
 sg13g2_decap_4 FILLER_32_427 ();
 sg13g2_fill_2 FILLER_32_448 ();
 sg13g2_fill_1 FILLER_32_450 ();
 sg13g2_fill_2 FILLER_32_456 ();
 sg13g2_fill_1 FILLER_32_461 ();
 sg13g2_decap_8 FILLER_32_470 ();
 sg13g2_fill_1 FILLER_32_484 ();
 sg13g2_fill_1 FILLER_32_498 ();
 sg13g2_fill_2 FILLER_32_517 ();
 sg13g2_fill_1 FILLER_32_519 ();
 sg13g2_fill_1 FILLER_32_529 ();
 sg13g2_fill_2 FILLER_32_538 ();
 sg13g2_fill_1 FILLER_32_540 ();
 sg13g2_fill_2 FILLER_32_567 ();
 sg13g2_fill_1 FILLER_32_578 ();
 sg13g2_fill_2 FILLER_32_583 ();
 sg13g2_fill_1 FILLER_32_585 ();
 sg13g2_decap_4 FILLER_32_616 ();
 sg13g2_fill_2 FILLER_32_620 ();
 sg13g2_fill_2 FILLER_32_634 ();
 sg13g2_decap_4 FILLER_32_645 ();
 sg13g2_decap_8 FILLER_32_653 ();
 sg13g2_decap_4 FILLER_32_660 ();
 sg13g2_fill_1 FILLER_32_664 ();
 sg13g2_fill_2 FILLER_32_669 ();
 sg13g2_fill_2 FILLER_32_676 ();
 sg13g2_fill_1 FILLER_32_682 ();
 sg13g2_fill_1 FILLER_32_711 ();
 sg13g2_fill_1 FILLER_32_717 ();
 sg13g2_fill_2 FILLER_32_723 ();
 sg13g2_fill_1 FILLER_32_725 ();
 sg13g2_fill_2 FILLER_32_732 ();
 sg13g2_decap_4 FILLER_32_742 ();
 sg13g2_fill_1 FILLER_32_746 ();
 sg13g2_decap_4 FILLER_32_755 ();
 sg13g2_fill_1 FILLER_32_759 ();
 sg13g2_fill_1 FILLER_32_765 ();
 sg13g2_fill_1 FILLER_32_774 ();
 sg13g2_fill_1 FILLER_32_780 ();
 sg13g2_decap_4 FILLER_32_794 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_fill_2 FILLER_32_822 ();
 sg13g2_fill_2 FILLER_32_829 ();
 sg13g2_fill_2 FILLER_32_848 ();
 sg13g2_fill_1 FILLER_32_850 ();
 sg13g2_decap_8 FILLER_32_857 ();
 sg13g2_fill_2 FILLER_32_864 ();
 sg13g2_fill_1 FILLER_32_871 ();
 sg13g2_fill_2 FILLER_32_896 ();
 sg13g2_fill_1 FILLER_32_902 ();
 sg13g2_fill_2 FILLER_32_932 ();
 sg13g2_fill_2 FILLER_32_938 ();
 sg13g2_fill_1 FILLER_32_940 ();
 sg13g2_decap_8 FILLER_32_951 ();
 sg13g2_fill_2 FILLER_32_967 ();
 sg13g2_fill_1 FILLER_32_969 ();
 sg13g2_fill_2 FILLER_32_989 ();
 sg13g2_fill_2 FILLER_32_1005 ();
 sg13g2_decap_8 FILLER_32_1011 ();
 sg13g2_decap_4 FILLER_32_1018 ();
 sg13g2_fill_1 FILLER_32_1022 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_fill_2 FILLER_32_1047 ();
 sg13g2_fill_2 FILLER_32_1053 ();
 sg13g2_fill_1 FILLER_32_1055 ();
 sg13g2_fill_1 FILLER_32_1061 ();
 sg13g2_fill_1 FILLER_32_1067 ();
 sg13g2_fill_1 FILLER_32_1076 ();
 sg13g2_fill_1 FILLER_32_1082 ();
 sg13g2_decap_4 FILLER_32_1093 ();
 sg13g2_fill_1 FILLER_32_1115 ();
 sg13g2_decap_8 FILLER_32_1120 ();
 sg13g2_decap_8 FILLER_32_1127 ();
 sg13g2_decap_8 FILLER_32_1134 ();
 sg13g2_fill_1 FILLER_32_1154 ();
 sg13g2_fill_2 FILLER_32_1160 ();
 sg13g2_fill_1 FILLER_32_1162 ();
 sg13g2_fill_2 FILLER_32_1172 ();
 sg13g2_fill_1 FILLER_32_1195 ();
 sg13g2_fill_1 FILLER_32_1204 ();
 sg13g2_fill_1 FILLER_32_1215 ();
 sg13g2_fill_2 FILLER_32_1220 ();
 sg13g2_fill_1 FILLER_32_1222 ();
 sg13g2_fill_2 FILLER_32_1227 ();
 sg13g2_fill_1 FILLER_32_1229 ();
 sg13g2_decap_4 FILLER_32_1240 ();
 sg13g2_fill_2 FILLER_32_1265 ();
 sg13g2_decap_8 FILLER_32_1275 ();
 sg13g2_decap_8 FILLER_32_1282 ();
 sg13g2_decap_4 FILLER_32_1289 ();
 sg13g2_fill_2 FILLER_32_1293 ();
 sg13g2_fill_2 FILLER_32_1299 ();
 sg13g2_fill_2 FILLER_32_1305 ();
 sg13g2_fill_1 FILLER_32_1307 ();
 sg13g2_fill_1 FILLER_32_1313 ();
 sg13g2_fill_1 FILLER_32_1317 ();
 sg13g2_fill_1 FILLER_32_1340 ();
 sg13g2_fill_1 FILLER_32_1359 ();
 sg13g2_fill_1 FILLER_32_1365 ();
 sg13g2_fill_2 FILLER_32_1378 ();
 sg13g2_fill_1 FILLER_32_1380 ();
 sg13g2_fill_2 FILLER_32_1390 ();
 sg13g2_fill_1 FILLER_32_1392 ();
 sg13g2_fill_1 FILLER_32_1401 ();
 sg13g2_decap_8 FILLER_32_1418 ();
 sg13g2_decap_4 FILLER_32_1425 ();
 sg13g2_fill_2 FILLER_32_1429 ();
 sg13g2_decap_8 FILLER_32_1439 ();
 sg13g2_decap_8 FILLER_32_1446 ();
 sg13g2_fill_2 FILLER_32_1473 ();
 sg13g2_fill_1 FILLER_32_1475 ();
 sg13g2_decap_8 FILLER_32_1495 ();
 sg13g2_fill_1 FILLER_32_1502 ();
 sg13g2_decap_4 FILLER_32_1511 ();
 sg13g2_fill_1 FILLER_32_1515 ();
 sg13g2_decap_4 FILLER_32_1521 ();
 sg13g2_fill_1 FILLER_32_1525 ();
 sg13g2_fill_1 FILLER_32_1530 ();
 sg13g2_decap_4 FILLER_32_1547 ();
 sg13g2_decap_8 FILLER_32_1564 ();
 sg13g2_decap_8 FILLER_32_1576 ();
 sg13g2_fill_1 FILLER_32_1583 ();
 sg13g2_fill_2 FILLER_32_1606 ();
 sg13g2_decap_4 FILLER_32_1613 ();
 sg13g2_fill_1 FILLER_32_1617 ();
 sg13g2_decap_8 FILLER_32_1622 ();
 sg13g2_fill_2 FILLER_32_1629 ();
 sg13g2_fill_1 FILLER_32_1631 ();
 sg13g2_fill_2 FILLER_32_1637 ();
 sg13g2_fill_2 FILLER_32_1661 ();
 sg13g2_fill_1 FILLER_32_1668 ();
 sg13g2_fill_1 FILLER_32_1684 ();
 sg13g2_fill_2 FILLER_32_1690 ();
 sg13g2_fill_2 FILLER_32_1695 ();
 sg13g2_decap_4 FILLER_32_1711 ();
 sg13g2_fill_1 FILLER_32_1715 ();
 sg13g2_decap_4 FILLER_32_1724 ();
 sg13g2_fill_1 FILLER_32_1728 ();
 sg13g2_decap_4 FILLER_32_1755 ();
 sg13g2_decap_8 FILLER_32_1763 ();
 sg13g2_decap_4 FILLER_32_1770 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_46 ();
 sg13g2_decap_8 FILLER_33_62 ();
 sg13g2_fill_1 FILLER_33_69 ();
 sg13g2_decap_4 FILLER_33_74 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_fill_2 FILLER_33_109 ();
 sg13g2_fill_1 FILLER_33_122 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_decap_4 FILLER_33_167 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_200 ();
 sg13g2_fill_1 FILLER_33_202 ();
 sg13g2_decap_8 FILLER_33_209 ();
 sg13g2_decap_8 FILLER_33_216 ();
 sg13g2_decap_4 FILLER_33_223 ();
 sg13g2_fill_2 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_decap_4 FILLER_33_253 ();
 sg13g2_decap_4 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_274 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_4 FILLER_33_415 ();
 sg13g2_fill_1 FILLER_33_419 ();
 sg13g2_decap_4 FILLER_33_431 ();
 sg13g2_fill_2 FILLER_33_459 ();
 sg13g2_fill_2 FILLER_33_465 ();
 sg13g2_decap_4 FILLER_33_472 ();
 sg13g2_fill_1 FILLER_33_476 ();
 sg13g2_decap_4 FILLER_33_481 ();
 sg13g2_fill_2 FILLER_33_485 ();
 sg13g2_fill_2 FILLER_33_497 ();
 sg13g2_decap_4 FILLER_33_532 ();
 sg13g2_fill_1 FILLER_33_536 ();
 sg13g2_fill_2 FILLER_33_550 ();
 sg13g2_fill_1 FILLER_33_552 ();
 sg13g2_fill_2 FILLER_33_566 ();
 sg13g2_fill_1 FILLER_33_568 ();
 sg13g2_decap_4 FILLER_33_577 ();
 sg13g2_decap_4 FILLER_33_589 ();
 sg13g2_fill_2 FILLER_33_598 ();
 sg13g2_fill_1 FILLER_33_600 ();
 sg13g2_fill_2 FILLER_33_609 ();
 sg13g2_fill_1 FILLER_33_611 ();
 sg13g2_fill_2 FILLER_33_620 ();
 sg13g2_fill_1 FILLER_33_622 ();
 sg13g2_fill_1 FILLER_33_639 ();
 sg13g2_decap_4 FILLER_33_644 ();
 sg13g2_fill_1 FILLER_33_648 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_fill_1 FILLER_33_665 ();
 sg13g2_fill_1 FILLER_33_675 ();
 sg13g2_fill_2 FILLER_33_684 ();
 sg13g2_fill_1 FILLER_33_694 ();
 sg13g2_fill_2 FILLER_33_700 ();
 sg13g2_fill_1 FILLER_33_702 ();
 sg13g2_fill_2 FILLER_33_708 ();
 sg13g2_fill_1 FILLER_33_710 ();
 sg13g2_fill_2 FILLER_33_751 ();
 sg13g2_fill_2 FILLER_33_761 ();
 sg13g2_decap_4 FILLER_33_788 ();
 sg13g2_fill_1 FILLER_33_811 ();
 sg13g2_fill_1 FILLER_33_817 ();
 sg13g2_decap_4 FILLER_33_829 ();
 sg13g2_fill_2 FILLER_33_837 ();
 sg13g2_fill_1 FILLER_33_839 ();
 sg13g2_fill_2 FILLER_33_845 ();
 sg13g2_fill_2 FILLER_33_852 ();
 sg13g2_fill_1 FILLER_33_854 ();
 sg13g2_fill_2 FILLER_33_859 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_33_881 ();
 sg13g2_decap_8 FILLER_33_892 ();
 sg13g2_fill_2 FILLER_33_899 ();
 sg13g2_fill_1 FILLER_33_901 ();
 sg13g2_fill_2 FILLER_33_910 ();
 sg13g2_fill_1 FILLER_33_912 ();
 sg13g2_fill_1 FILLER_33_923 ();
 sg13g2_fill_1 FILLER_33_934 ();
 sg13g2_decap_8 FILLER_33_943 ();
 sg13g2_decap_4 FILLER_33_950 ();
 sg13g2_fill_1 FILLER_33_978 ();
 sg13g2_fill_1 FILLER_33_984 ();
 sg13g2_fill_2 FILLER_33_988 ();
 sg13g2_decap_8 FILLER_33_1058 ();
 sg13g2_decap_8 FILLER_33_1065 ();
 sg13g2_decap_8 FILLER_33_1077 ();
 sg13g2_decap_8 FILLER_33_1084 ();
 sg13g2_fill_2 FILLER_33_1091 ();
 sg13g2_fill_2 FILLER_33_1096 ();
 sg13g2_fill_1 FILLER_33_1098 ();
 sg13g2_decap_8 FILLER_33_1124 ();
 sg13g2_decap_4 FILLER_33_1131 ();
 sg13g2_fill_1 FILLER_33_1159 ();
 sg13g2_decap_4 FILLER_33_1169 ();
 sg13g2_fill_1 FILLER_33_1173 ();
 sg13g2_decap_8 FILLER_33_1178 ();
 sg13g2_decap_4 FILLER_33_1185 ();
 sg13g2_fill_2 FILLER_33_1207 ();
 sg13g2_fill_1 FILLER_33_1209 ();
 sg13g2_decap_4 FILLER_33_1217 ();
 sg13g2_fill_1 FILLER_33_1221 ();
 sg13g2_decap_4 FILLER_33_1233 ();
 sg13g2_fill_2 FILLER_33_1237 ();
 sg13g2_fill_1 FILLER_33_1247 ();
 sg13g2_fill_1 FILLER_33_1253 ();
 sg13g2_decap_4 FILLER_33_1275 ();
 sg13g2_fill_2 FILLER_33_1279 ();
 sg13g2_decap_4 FILLER_33_1295 ();
 sg13g2_fill_2 FILLER_33_1304 ();
 sg13g2_fill_1 FILLER_33_1306 ();
 sg13g2_decap_4 FILLER_33_1312 ();
 sg13g2_fill_1 FILLER_33_1321 ();
 sg13g2_decap_4 FILLER_33_1327 ();
 sg13g2_fill_1 FILLER_33_1344 ();
 sg13g2_fill_1 FILLER_33_1356 ();
 sg13g2_fill_1 FILLER_33_1367 ();
 sg13g2_fill_1 FILLER_33_1377 ();
 sg13g2_fill_2 FILLER_33_1400 ();
 sg13g2_decap_4 FILLER_33_1434 ();
 sg13g2_fill_1 FILLER_33_1471 ();
 sg13g2_decap_4 FILLER_33_1478 ();
 sg13g2_decap_4 FILLER_33_1489 ();
 sg13g2_fill_2 FILLER_33_1493 ();
 sg13g2_decap_4 FILLER_33_1503 ();
 sg13g2_fill_2 FILLER_33_1512 ();
 sg13g2_fill_1 FILLER_33_1514 ();
 sg13g2_decap_8 FILLER_33_1519 ();
 sg13g2_fill_2 FILLER_33_1526 ();
 sg13g2_fill_1 FILLER_33_1544 ();
 sg13g2_fill_2 FILLER_33_1559 ();
 sg13g2_fill_1 FILLER_33_1561 ();
 sg13g2_decap_8 FILLER_33_1575 ();
 sg13g2_decap_8 FILLER_33_1590 ();
 sg13g2_decap_8 FILLER_33_1597 ();
 sg13g2_fill_2 FILLER_33_1604 ();
 sg13g2_decap_4 FILLER_33_1622 ();
 sg13g2_fill_2 FILLER_33_1626 ();
 sg13g2_fill_2 FILLER_33_1632 ();
 sg13g2_fill_1 FILLER_33_1651 ();
 sg13g2_fill_1 FILLER_33_1667 ();
 sg13g2_fill_1 FILLER_33_1676 ();
 sg13g2_decap_8 FILLER_33_1698 ();
 sg13g2_decap_8 FILLER_33_1705 ();
 sg13g2_decap_4 FILLER_33_1712 ();
 sg13g2_fill_2 FILLER_33_1721 ();
 sg13g2_decap_8 FILLER_33_1758 ();
 sg13g2_decap_8 FILLER_33_1765 ();
 sg13g2_fill_2 FILLER_33_1772 ();
 sg13g2_fill_2 FILLER_34_30 ();
 sg13g2_fill_2 FILLER_34_53 ();
 sg13g2_decap_4 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_69 ();
 sg13g2_fill_1 FILLER_34_85 ();
 sg13g2_fill_1 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_152 ();
 sg13g2_decap_8 FILLER_34_180 ();
 sg13g2_decap_8 FILLER_34_187 ();
 sg13g2_fill_1 FILLER_34_199 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_fill_2 FILLER_34_219 ();
 sg13g2_decap_8 FILLER_34_226 ();
 sg13g2_decap_8 FILLER_34_233 ();
 sg13g2_decap_8 FILLER_34_240 ();
 sg13g2_decap_8 FILLER_34_247 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_decap_8 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_303 ();
 sg13g2_decap_8 FILLER_34_310 ();
 sg13g2_decap_4 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_404 ();
 sg13g2_decap_8 FILLER_34_411 ();
 sg13g2_fill_2 FILLER_34_418 ();
 sg13g2_fill_1 FILLER_34_420 ();
 sg13g2_fill_2 FILLER_34_431 ();
 sg13g2_decap_4 FILLER_34_451 ();
 sg13g2_decap_8 FILLER_34_465 ();
 sg13g2_decap_8 FILLER_34_472 ();
 sg13g2_decap_8 FILLER_34_479 ();
 sg13g2_decap_4 FILLER_34_486 ();
 sg13g2_fill_2 FILLER_34_499 ();
 sg13g2_fill_1 FILLER_34_501 ();
 sg13g2_decap_8 FILLER_34_513 ();
 sg13g2_decap_8 FILLER_34_520 ();
 sg13g2_fill_2 FILLER_34_527 ();
 sg13g2_fill_1 FILLER_34_529 ();
 sg13g2_fill_2 FILLER_34_535 ();
 sg13g2_fill_1 FILLER_34_537 ();
 sg13g2_decap_4 FILLER_34_546 ();
 sg13g2_fill_2 FILLER_34_550 ();
 sg13g2_decap_4 FILLER_34_557 ();
 sg13g2_decap_8 FILLER_34_569 ();
 sg13g2_fill_1 FILLER_34_576 ();
 sg13g2_fill_2 FILLER_34_585 ();
 sg13g2_fill_1 FILLER_34_587 ();
 sg13g2_fill_2 FILLER_34_593 ();
 sg13g2_fill_1 FILLER_34_595 ();
 sg13g2_fill_1 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_618 ();
 sg13g2_fill_2 FILLER_34_625 ();
 sg13g2_decap_8 FILLER_34_636 ();
 sg13g2_fill_2 FILLER_34_643 ();
 sg13g2_decap_4 FILLER_34_658 ();
 sg13g2_fill_2 FILLER_34_662 ();
 sg13g2_fill_1 FILLER_34_668 ();
 sg13g2_fill_2 FILLER_34_697 ();
 sg13g2_fill_2 FILLER_34_705 ();
 sg13g2_fill_1 FILLER_34_707 ();
 sg13g2_fill_2 FILLER_34_731 ();
 sg13g2_fill_2 FILLER_34_741 ();
 sg13g2_fill_2 FILLER_34_752 ();
 sg13g2_fill_1 FILLER_34_766 ();
 sg13g2_fill_2 FILLER_34_780 ();
 sg13g2_fill_1 FILLER_34_790 ();
 sg13g2_fill_2 FILLER_34_804 ();
 sg13g2_fill_1 FILLER_34_806 ();
 sg13g2_fill_2 FILLER_34_826 ();
 sg13g2_fill_1 FILLER_34_828 ();
 sg13g2_decap_4 FILLER_34_834 ();
 sg13g2_decap_8 FILLER_34_842 ();
 sg13g2_fill_2 FILLER_34_849 ();
 sg13g2_fill_1 FILLER_34_851 ();
 sg13g2_decap_4 FILLER_34_880 ();
 sg13g2_decap_8 FILLER_34_889 ();
 sg13g2_fill_2 FILLER_34_912 ();
 sg13g2_fill_1 FILLER_34_921 ();
 sg13g2_fill_2 FILLER_34_927 ();
 sg13g2_fill_1 FILLER_34_935 ();
 sg13g2_fill_2 FILLER_34_941 ();
 sg13g2_decap_8 FILLER_34_948 ();
 sg13g2_fill_2 FILLER_34_955 ();
 sg13g2_fill_1 FILLER_34_957 ();
 sg13g2_fill_1 FILLER_34_975 ();
 sg13g2_fill_1 FILLER_34_984 ();
 sg13g2_fill_1 FILLER_34_990 ();
 sg13g2_fill_2 FILLER_34_1007 ();
 sg13g2_fill_1 FILLER_34_1014 ();
 sg13g2_fill_1 FILLER_34_1020 ();
 sg13g2_decap_8 FILLER_34_1026 ();
 sg13g2_decap_8 FILLER_34_1033 ();
 sg13g2_decap_8 FILLER_34_1040 ();
 sg13g2_decap_8 FILLER_34_1047 ();
 sg13g2_decap_4 FILLER_34_1107 ();
 sg13g2_decap_8 FILLER_34_1116 ();
 sg13g2_decap_4 FILLER_34_1123 ();
 sg13g2_fill_2 FILLER_34_1127 ();
 sg13g2_fill_1 FILLER_34_1164 ();
 sg13g2_fill_2 FILLER_34_1169 ();
 sg13g2_decap_4 FILLER_34_1176 ();
 sg13g2_fill_1 FILLER_34_1180 ();
 sg13g2_fill_2 FILLER_34_1186 ();
 sg13g2_fill_1 FILLER_34_1188 ();
 sg13g2_decap_4 FILLER_34_1194 ();
 sg13g2_fill_1 FILLER_34_1198 ();
 sg13g2_fill_1 FILLER_34_1204 ();
 sg13g2_decap_4 FILLER_34_1210 ();
 sg13g2_fill_1 FILLER_34_1227 ();
 sg13g2_fill_1 FILLER_34_1233 ();
 sg13g2_fill_1 FILLER_34_1238 ();
 sg13g2_fill_1 FILLER_34_1253 ();
 sg13g2_decap_8 FILLER_34_1264 ();
 sg13g2_fill_1 FILLER_34_1271 ();
 sg13g2_decap_8 FILLER_34_1277 ();
 sg13g2_fill_2 FILLER_34_1284 ();
 sg13g2_fill_1 FILLER_34_1296 ();
 sg13g2_fill_1 FILLER_34_1301 ();
 sg13g2_fill_1 FILLER_34_1327 ();
 sg13g2_fill_1 FILLER_34_1338 ();
 sg13g2_decap_8 FILLER_34_1371 ();
 sg13g2_fill_2 FILLER_34_1378 ();
 sg13g2_fill_1 FILLER_34_1393 ();
 sg13g2_fill_2 FILLER_34_1398 ();
 sg13g2_decap_8 FILLER_34_1423 ();
 sg13g2_decap_4 FILLER_34_1430 ();
 sg13g2_decap_8 FILLER_34_1439 ();
 sg13g2_decap_8 FILLER_34_1446 ();
 sg13g2_decap_4 FILLER_34_1453 ();
 sg13g2_fill_1 FILLER_34_1457 ();
 sg13g2_decap_4 FILLER_34_1468 ();
 sg13g2_fill_1 FILLER_34_1477 ();
 sg13g2_fill_2 FILLER_34_1490 ();
 sg13g2_decap_4 FILLER_34_1519 ();
 sg13g2_decap_8 FILLER_34_1527 ();
 sg13g2_fill_2 FILLER_34_1534 ();
 sg13g2_decap_4 FILLER_34_1541 ();
 sg13g2_fill_1 FILLER_34_1545 ();
 sg13g2_decap_8 FILLER_34_1554 ();
 sg13g2_decap_4 FILLER_34_1574 ();
 sg13g2_fill_1 FILLER_34_1625 ();
 sg13g2_decap_8 FILLER_34_1630 ();
 sg13g2_fill_2 FILLER_34_1649 ();
 sg13g2_fill_2 FILLER_34_1694 ();
 sg13g2_decap_8 FILLER_34_1708 ();
 sg13g2_decap_4 FILLER_34_1715 ();
 sg13g2_fill_2 FILLER_34_1719 ();
 sg13g2_fill_1 FILLER_34_1735 ();
 sg13g2_decap_8 FILLER_34_1748 ();
 sg13g2_decap_8 FILLER_34_1755 ();
 sg13g2_decap_8 FILLER_34_1762 ();
 sg13g2_decap_4 FILLER_34_1769 ();
 sg13g2_fill_1 FILLER_34_1773 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_decap_4 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_18 ();
 sg13g2_fill_2 FILLER_35_24 ();
 sg13g2_decap_4 FILLER_35_30 ();
 sg13g2_fill_1 FILLER_35_34 ();
 sg13g2_fill_2 FILLER_35_48 ();
 sg13g2_fill_2 FILLER_35_55 ();
 sg13g2_fill_1 FILLER_35_57 ();
 sg13g2_decap_4 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_67 ();
 sg13g2_fill_2 FILLER_35_82 ();
 sg13g2_fill_1 FILLER_35_110 ();
 sg13g2_fill_2 FILLER_35_141 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_decap_4 FILLER_35_179 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_decap_8 FILLER_35_201 ();
 sg13g2_fill_1 FILLER_35_225 ();
 sg13g2_fill_2 FILLER_35_236 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_258 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_decap_4 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_306 ();
 sg13g2_decap_8 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_320 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_fill_2 FILLER_35_383 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_4 FILLER_35_441 ();
 sg13g2_fill_2 FILLER_35_457 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_fill_2 FILLER_35_483 ();
 sg13g2_fill_1 FILLER_35_485 ();
 sg13g2_fill_2 FILLER_35_500 ();
 sg13g2_decap_8 FILLER_35_509 ();
 sg13g2_fill_2 FILLER_35_516 ();
 sg13g2_decap_4 FILLER_35_527 ();
 sg13g2_fill_2 FILLER_35_531 ();
 sg13g2_decap_8 FILLER_35_559 ();
 sg13g2_decap_8 FILLER_35_566 ();
 sg13g2_decap_4 FILLER_35_573 ();
 sg13g2_decap_8 FILLER_35_585 ();
 sg13g2_decap_4 FILLER_35_592 ();
 sg13g2_fill_1 FILLER_35_611 ();
 sg13g2_decap_4 FILLER_35_624 ();
 sg13g2_fill_2 FILLER_35_628 ();
 sg13g2_decap_8 FILLER_35_641 ();
 sg13g2_decap_4 FILLER_35_648 ();
 sg13g2_fill_2 FILLER_35_660 ();
 sg13g2_fill_1 FILLER_35_670 ();
 sg13g2_fill_1 FILLER_35_679 ();
 sg13g2_fill_2 FILLER_35_703 ();
 sg13g2_decap_8 FILLER_35_710 ();
 sg13g2_fill_1 FILLER_35_717 ();
 sg13g2_fill_1 FILLER_35_721 ();
 sg13g2_decap_4 FILLER_35_730 ();
 sg13g2_fill_1 FILLER_35_734 ();
 sg13g2_decap_4 FILLER_35_740 ();
 sg13g2_fill_2 FILLER_35_744 ();
 sg13g2_fill_2 FILLER_35_758 ();
 sg13g2_decap_4 FILLER_35_797 ();
 sg13g2_fill_1 FILLER_35_801 ();
 sg13g2_fill_1 FILLER_35_818 ();
 sg13g2_fill_1 FILLER_35_830 ();
 sg13g2_fill_1 FILLER_35_845 ();
 sg13g2_fill_2 FILLER_35_850 ();
 sg13g2_fill_1 FILLER_35_862 ();
 sg13g2_fill_1 FILLER_35_874 ();
 sg13g2_fill_2 FILLER_35_887 ();
 sg13g2_fill_2 FILLER_35_909 ();
 sg13g2_fill_1 FILLER_35_911 ();
 sg13g2_fill_2 FILLER_35_924 ();
 sg13g2_fill_1 FILLER_35_926 ();
 sg13g2_decap_8 FILLER_35_950 ();
 sg13g2_fill_1 FILLER_35_962 ();
 sg13g2_fill_1 FILLER_35_970 ();
 sg13g2_fill_2 FILLER_35_979 ();
 sg13g2_fill_2 FILLER_35_1030 ();
 sg13g2_fill_1 FILLER_35_1032 ();
 sg13g2_fill_2 FILLER_35_1044 ();
 sg13g2_decap_4 FILLER_35_1051 ();
 sg13g2_fill_1 FILLER_35_1055 ();
 sg13g2_decap_4 FILLER_35_1061 ();
 sg13g2_fill_2 FILLER_35_1081 ();
 sg13g2_fill_1 FILLER_35_1096 ();
 sg13g2_fill_1 FILLER_35_1111 ();
 sg13g2_fill_2 FILLER_35_1129 ();
 sg13g2_fill_2 FILLER_35_1134 ();
 sg13g2_fill_2 FILLER_35_1140 ();
 sg13g2_fill_1 FILLER_35_1158 ();
 sg13g2_fill_1 FILLER_35_1162 ();
 sg13g2_fill_1 FILLER_35_1168 ();
 sg13g2_decap_8 FILLER_35_1173 ();
 sg13g2_decap_4 FILLER_35_1195 ();
 sg13g2_fill_2 FILLER_35_1199 ();
 sg13g2_decap_8 FILLER_35_1209 ();
 sg13g2_decap_4 FILLER_35_1216 ();
 sg13g2_fill_1 FILLER_35_1220 ();
 sg13g2_decap_4 FILLER_35_1225 ();
 sg13g2_decap_4 FILLER_35_1241 ();
 sg13g2_fill_1 FILLER_35_1277 ();
 sg13g2_decap_4 FILLER_35_1299 ();
 sg13g2_fill_1 FILLER_35_1307 ();
 sg13g2_fill_1 FILLER_35_1312 ();
 sg13g2_fill_2 FILLER_35_1317 ();
 sg13g2_fill_2 FILLER_35_1324 ();
 sg13g2_fill_1 FILLER_35_1332 ();
 sg13g2_fill_2 FILLER_35_1351 ();
 sg13g2_decap_8 FILLER_35_1367 ();
 sg13g2_fill_2 FILLER_35_1374 ();
 sg13g2_fill_2 FILLER_35_1389 ();
 sg13g2_fill_1 FILLER_35_1399 ();
 sg13g2_fill_1 FILLER_35_1406 ();
 sg13g2_fill_1 FILLER_35_1417 ();
 sg13g2_decap_8 FILLER_35_1422 ();
 sg13g2_fill_1 FILLER_35_1429 ();
 sg13g2_decap_8 FILLER_35_1435 ();
 sg13g2_fill_1 FILLER_35_1442 ();
 sg13g2_fill_2 FILLER_35_1451 ();
 sg13g2_fill_2 FILLER_35_1458 ();
 sg13g2_fill_1 FILLER_35_1460 ();
 sg13g2_fill_2 FILLER_35_1469 ();
 sg13g2_fill_1 FILLER_35_1476 ();
 sg13g2_decap_4 FILLER_35_1483 ();
 sg13g2_fill_1 FILLER_35_1503 ();
 sg13g2_fill_1 FILLER_35_1511 ();
 sg13g2_fill_2 FILLER_35_1517 ();
 sg13g2_fill_1 FILLER_35_1554 ();
 sg13g2_decap_4 FILLER_35_1563 ();
 sg13g2_fill_2 FILLER_35_1567 ();
 sg13g2_decap_4 FILLER_35_1573 ();
 sg13g2_decap_8 FILLER_35_1582 ();
 sg13g2_decap_8 FILLER_35_1589 ();
 sg13g2_decap_8 FILLER_35_1596 ();
 sg13g2_fill_1 FILLER_35_1603 ();
 sg13g2_fill_1 FILLER_35_1612 ();
 sg13g2_decap_4 FILLER_35_1621 ();
 sg13g2_decap_8 FILLER_35_1637 ();
 sg13g2_fill_1 FILLER_35_1644 ();
 sg13g2_fill_1 FILLER_35_1657 ();
 sg13g2_fill_1 FILLER_35_1665 ();
 sg13g2_fill_1 FILLER_35_1709 ();
 sg13g2_decap_8 FILLER_35_1715 ();
 sg13g2_fill_2 FILLER_35_1722 ();
 sg13g2_fill_1 FILLER_35_1728 ();
 sg13g2_decap_8 FILLER_35_1764 ();
 sg13g2_fill_2 FILLER_35_1771 ();
 sg13g2_fill_1 FILLER_35_1773 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_12 ();
 sg13g2_decap_8 FILLER_36_26 ();
 sg13g2_decap_4 FILLER_36_37 ();
 sg13g2_fill_2 FILLER_36_60 ();
 sg13g2_fill_1 FILLER_36_67 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_decap_8 FILLER_36_94 ();
 sg13g2_fill_1 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_130 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_decap_4 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_204 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_fill_2 FILLER_36_221 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_fill_2 FILLER_36_241 ();
 sg13g2_decap_4 FILLER_36_248 ();
 sg13g2_fill_1 FILLER_36_252 ();
 sg13g2_decap_4 FILLER_36_258 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_decap_8 FILLER_36_268 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_282 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_fill_1 FILLER_36_349 ();
 sg13g2_fill_1 FILLER_36_379 ();
 sg13g2_fill_2 FILLER_36_387 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_407 ();
 sg13g2_fill_2 FILLER_36_411 ();
 sg13g2_fill_1 FILLER_36_421 ();
 sg13g2_fill_2 FILLER_36_448 ();
 sg13g2_decap_4 FILLER_36_458 ();
 sg13g2_fill_1 FILLER_36_462 ();
 sg13g2_fill_2 FILLER_36_500 ();
 sg13g2_fill_2 FILLER_36_536 ();
 sg13g2_fill_1 FILLER_36_538 ();
 sg13g2_decap_8 FILLER_36_547 ();
 sg13g2_fill_2 FILLER_36_554 ();
 sg13g2_decap_4 FILLER_36_577 ();
 sg13g2_fill_1 FILLER_36_581 ();
 sg13g2_fill_2 FILLER_36_624 ();
 sg13g2_fill_1 FILLER_36_636 ();
 sg13g2_decap_8 FILLER_36_641 ();
 sg13g2_decap_4 FILLER_36_662 ();
 sg13g2_fill_1 FILLER_36_670 ();
 sg13g2_fill_1 FILLER_36_679 ();
 sg13g2_fill_2 FILLER_36_690 ();
 sg13g2_fill_1 FILLER_36_692 ();
 sg13g2_decap_4 FILLER_36_714 ();
 sg13g2_fill_2 FILLER_36_718 ();
 sg13g2_fill_2 FILLER_36_728 ();
 sg13g2_fill_1 FILLER_36_730 ();
 sg13g2_decap_8 FILLER_36_735 ();
 sg13g2_decap_4 FILLER_36_746 ();
 sg13g2_fill_2 FILLER_36_766 ();
 sg13g2_fill_2 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_796 ();
 sg13g2_decap_4 FILLER_36_803 ();
 sg13g2_decap_8 FILLER_36_811 ();
 sg13g2_fill_1 FILLER_36_818 ();
 sg13g2_decap_8 FILLER_36_836 ();
 sg13g2_decap_8 FILLER_36_843 ();
 sg13g2_fill_1 FILLER_36_875 ();
 sg13g2_fill_1 FILLER_36_885 ();
 sg13g2_decap_4 FILLER_36_892 ();
 sg13g2_fill_2 FILLER_36_896 ();
 sg13g2_fill_2 FILLER_36_903 ();
 sg13g2_fill_1 FILLER_36_905 ();
 sg13g2_fill_1 FILLER_36_914 ();
 sg13g2_fill_1 FILLER_36_923 ();
 sg13g2_fill_1 FILLER_36_931 ();
 sg13g2_fill_2 FILLER_36_936 ();
 sg13g2_fill_1 FILLER_36_938 ();
 sg13g2_decap_8 FILLER_36_943 ();
 sg13g2_decap_4 FILLER_36_950 ();
 sg13g2_decap_4 FILLER_36_966 ();
 sg13g2_fill_2 FILLER_36_986 ();
 sg13g2_decap_4 FILLER_36_1000 ();
 sg13g2_fill_1 FILLER_36_1004 ();
 sg13g2_decap_4 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1025 ();
 sg13g2_decap_8 FILLER_36_1032 ();
 sg13g2_decap_8 FILLER_36_1039 ();
 sg13g2_fill_1 FILLER_36_1046 ();
 sg13g2_fill_1 FILLER_36_1063 ();
 sg13g2_fill_1 FILLER_36_1074 ();
 sg13g2_fill_1 FILLER_36_1095 ();
 sg13g2_fill_1 FILLER_36_1101 ();
 sg13g2_fill_1 FILLER_36_1107 ();
 sg13g2_fill_1 FILLER_36_1113 ();
 sg13g2_decap_4 FILLER_36_1133 ();
 sg13g2_fill_1 FILLER_36_1137 ();
 sg13g2_fill_1 FILLER_36_1164 ();
 sg13g2_decap_4 FILLER_36_1168 ();
 sg13g2_fill_2 FILLER_36_1185 ();
 sg13g2_fill_2 FILLER_36_1197 ();
 sg13g2_fill_2 FILLER_36_1208 ();
 sg13g2_fill_1 FILLER_36_1210 ();
 sg13g2_decap_4 FILLER_36_1243 ();
 sg13g2_fill_2 FILLER_36_1247 ();
 sg13g2_decap_8 FILLER_36_1258 ();
 sg13g2_decap_8 FILLER_36_1265 ();
 sg13g2_fill_1 FILLER_36_1272 ();
 sg13g2_decap_4 FILLER_36_1304 ();
 sg13g2_fill_2 FILLER_36_1320 ();
 sg13g2_fill_1 FILLER_36_1326 ();
 sg13g2_decap_4 FILLER_36_1337 ();
 sg13g2_fill_2 FILLER_36_1354 ();
 sg13g2_decap_4 FILLER_36_1360 ();
 sg13g2_fill_1 FILLER_36_1364 ();
 sg13g2_fill_1 FILLER_36_1369 ();
 sg13g2_decap_8 FILLER_36_1383 ();
 sg13g2_fill_1 FILLER_36_1390 ();
 sg13g2_decap_8 FILLER_36_1396 ();
 sg13g2_fill_1 FILLER_36_1403 ();
 sg13g2_decap_8 FILLER_36_1408 ();
 sg13g2_fill_1 FILLER_36_1415 ();
 sg13g2_fill_1 FILLER_36_1419 ();
 sg13g2_decap_8 FILLER_36_1425 ();
 sg13g2_fill_1 FILLER_36_1432 ();
 sg13g2_fill_1 FILLER_36_1437 ();
 sg13g2_fill_2 FILLER_36_1454 ();
 sg13g2_fill_1 FILLER_36_1456 ();
 sg13g2_decap_4 FILLER_36_1490 ();
 sg13g2_fill_2 FILLER_36_1494 ();
 sg13g2_decap_8 FILLER_36_1517 ();
 sg13g2_fill_2 FILLER_36_1524 ();
 sg13g2_decap_4 FILLER_36_1530 ();
 sg13g2_fill_1 FILLER_36_1550 ();
 sg13g2_fill_1 FILLER_36_1560 ();
 sg13g2_fill_1 FILLER_36_1569 ();
 sg13g2_fill_1 FILLER_36_1602 ();
 sg13g2_decap_4 FILLER_36_1607 ();
 sg13g2_fill_2 FILLER_36_1611 ();
 sg13g2_fill_2 FILLER_36_1627 ();
 sg13g2_fill_1 FILLER_36_1629 ();
 sg13g2_fill_1 FILLER_36_1634 ();
 sg13g2_fill_1 FILLER_36_1650 ();
 sg13g2_fill_1 FILLER_36_1656 ();
 sg13g2_fill_1 FILLER_36_1660 ();
 sg13g2_decap_8 FILLER_36_1716 ();
 sg13g2_decap_4 FILLER_36_1727 ();
 sg13g2_fill_1 FILLER_36_1731 ();
 sg13g2_decap_4 FILLER_36_1737 ();
 sg13g2_decap_4 FILLER_36_1759 ();
 sg13g2_fill_2 FILLER_36_1763 ();
 sg13g2_decap_4 FILLER_36_1769 ();
 sg13g2_fill_1 FILLER_36_1773 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_18 ();
 sg13g2_decap_8 FILLER_37_44 ();
 sg13g2_decap_4 FILLER_37_51 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_decap_4 FILLER_37_72 ();
 sg13g2_fill_2 FILLER_37_76 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_111 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_125 ();
 sg13g2_fill_1 FILLER_37_131 ();
 sg13g2_decap_8 FILLER_37_142 ();
 sg13g2_decap_8 FILLER_37_149 ();
 sg13g2_decap_4 FILLER_37_156 ();
 sg13g2_fill_2 FILLER_37_160 ();
 sg13g2_decap_8 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_180 ();
 sg13g2_fill_2 FILLER_37_187 ();
 sg13g2_decap_4 FILLER_37_222 ();
 sg13g2_fill_1 FILLER_37_233 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_275 ();
 sg13g2_fill_1 FILLER_37_282 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_321 ();
 sg13g2_fill_2 FILLER_37_334 ();
 sg13g2_fill_2 FILLER_37_383 ();
 sg13g2_fill_1 FILLER_37_385 ();
 sg13g2_fill_2 FILLER_37_404 ();
 sg13g2_decap_8 FILLER_37_411 ();
 sg13g2_fill_1 FILLER_37_418 ();
 sg13g2_decap_4 FILLER_37_440 ();
 sg13g2_fill_2 FILLER_37_444 ();
 sg13g2_decap_4 FILLER_37_450 ();
 sg13g2_decap_8 FILLER_37_458 ();
 sg13g2_decap_8 FILLER_37_465 ();
 sg13g2_decap_4 FILLER_37_476 ();
 sg13g2_fill_2 FILLER_37_480 ();
 sg13g2_fill_1 FILLER_37_495 ();
 sg13g2_decap_4 FILLER_37_511 ();
 sg13g2_fill_1 FILLER_37_515 ();
 sg13g2_fill_1 FILLER_37_524 ();
 sg13g2_decap_4 FILLER_37_533 ();
 sg13g2_fill_1 FILLER_37_537 ();
 sg13g2_fill_2 FILLER_37_559 ();
 sg13g2_decap_4 FILLER_37_574 ();
 sg13g2_fill_1 FILLER_37_578 ();
 sg13g2_decap_8 FILLER_37_584 ();
 sg13g2_decap_8 FILLER_37_591 ();
 sg13g2_fill_2 FILLER_37_639 ();
 sg13g2_fill_1 FILLER_37_641 ();
 sg13g2_fill_1 FILLER_37_647 ();
 sg13g2_decap_4 FILLER_37_653 ();
 sg13g2_fill_1 FILLER_37_660 ();
 sg13g2_fill_1 FILLER_37_670 ();
 sg13g2_decap_4 FILLER_37_675 ();
 sg13g2_fill_2 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_4 FILLER_37_714 ();
 sg13g2_fill_2 FILLER_37_718 ();
 sg13g2_decap_4 FILLER_37_728 ();
 sg13g2_decap_4 FILLER_37_762 ();
 sg13g2_decap_8 FILLER_37_804 ();
 sg13g2_decap_8 FILLER_37_815 ();
 sg13g2_fill_1 FILLER_37_822 ();
 sg13g2_decap_4 FILLER_37_831 ();
 sg13g2_fill_1 FILLER_37_835 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_4 FILLER_37_847 ();
 sg13g2_decap_4 FILLER_37_855 ();
 sg13g2_fill_1 FILLER_37_867 ();
 sg13g2_fill_2 FILLER_37_880 ();
 sg13g2_fill_2 FILLER_37_904 ();
 sg13g2_fill_1 FILLER_37_906 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_decap_4 FILLER_37_924 ();
 sg13g2_fill_2 FILLER_37_928 ();
 sg13g2_decap_4 FILLER_37_936 ();
 sg13g2_fill_2 FILLER_37_940 ();
 sg13g2_decap_8 FILLER_37_947 ();
 sg13g2_decap_4 FILLER_37_954 ();
 sg13g2_fill_2 FILLER_37_958 ();
 sg13g2_decap_4 FILLER_37_968 ();
 sg13g2_fill_1 FILLER_37_972 ();
 sg13g2_fill_2 FILLER_37_988 ();
 sg13g2_fill_1 FILLER_37_1003 ();
 sg13g2_decap_8 FILLER_37_1008 ();
 sg13g2_fill_2 FILLER_37_1015 ();
 sg13g2_fill_1 FILLER_37_1024 ();
 sg13g2_decap_4 FILLER_37_1030 ();
 sg13g2_fill_2 FILLER_37_1047 ();
 sg13g2_fill_1 FILLER_37_1074 ();
 sg13g2_decap_4 FILLER_37_1091 ();
 sg13g2_fill_1 FILLER_37_1103 ();
 sg13g2_fill_1 FILLER_37_1109 ();
 sg13g2_fill_1 FILLER_37_1115 ();
 sg13g2_fill_2 FILLER_37_1125 ();
 sg13g2_fill_1 FILLER_37_1127 ();
 sg13g2_decap_8 FILLER_37_1137 ();
 sg13g2_decap_8 FILLER_37_1144 ();
 sg13g2_fill_2 FILLER_37_1151 ();
 sg13g2_fill_1 FILLER_37_1153 ();
 sg13g2_decap_4 FILLER_37_1159 ();
 sg13g2_fill_2 FILLER_37_1163 ();
 sg13g2_fill_1 FILLER_37_1189 ();
 sg13g2_decap_8 FILLER_37_1210 ();
 sg13g2_decap_8 FILLER_37_1222 ();
 sg13g2_decap_8 FILLER_37_1229 ();
 sg13g2_decap_8 FILLER_37_1236 ();
 sg13g2_decap_8 FILLER_37_1243 ();
 sg13g2_fill_1 FILLER_37_1250 ();
 sg13g2_fill_2 FILLER_37_1258 ();
 sg13g2_decap_8 FILLER_37_1280 ();
 sg13g2_decap_8 FILLER_37_1361 ();
 sg13g2_fill_1 FILLER_37_1368 ();
 sg13g2_decap_4 FILLER_37_1378 ();
 sg13g2_fill_2 FILLER_37_1382 ();
 sg13g2_decap_8 FILLER_37_1388 ();
 sg13g2_fill_1 FILLER_37_1395 ();
 sg13g2_fill_1 FILLER_37_1401 ();
 sg13g2_decap_4 FILLER_37_1412 ();
 sg13g2_fill_1 FILLER_37_1416 ();
 sg13g2_decap_8 FILLER_37_1422 ();
 sg13g2_fill_1 FILLER_37_1429 ();
 sg13g2_decap_8 FILLER_37_1439 ();
 sg13g2_decap_8 FILLER_37_1450 ();
 sg13g2_fill_1 FILLER_37_1457 ();
 sg13g2_fill_2 FILLER_37_1471 ();
 sg13g2_decap_8 FILLER_37_1481 ();
 sg13g2_decap_8 FILLER_37_1488 ();
 sg13g2_fill_2 FILLER_37_1499 ();
 sg13g2_fill_2 FILLER_37_1506 ();
 sg13g2_decap_8 FILLER_37_1513 ();
 sg13g2_fill_2 FILLER_37_1520 ();
 sg13g2_decap_8 FILLER_37_1526 ();
 sg13g2_decap_4 FILLER_37_1533 ();
 sg13g2_decap_4 FILLER_37_1550 ();
 sg13g2_fill_1 FILLER_37_1554 ();
 sg13g2_fill_1 FILLER_37_1571 ();
 sg13g2_fill_2 FILLER_37_1586 ();
 sg13g2_decap_8 FILLER_37_1601 ();
 sg13g2_fill_2 FILLER_37_1608 ();
 sg13g2_fill_1 FILLER_37_1610 ();
 sg13g2_fill_1 FILLER_37_1625 ();
 sg13g2_fill_2 FILLER_37_1637 ();
 sg13g2_fill_1 FILLER_37_1639 ();
 sg13g2_fill_1 FILLER_37_1653 ();
 sg13g2_fill_2 FILLER_37_1668 ();
 sg13g2_fill_1 FILLER_37_1675 ();
 sg13g2_decap_8 FILLER_37_1684 ();
 sg13g2_decap_8 FILLER_37_1691 ();
 sg13g2_fill_1 FILLER_37_1698 ();
 sg13g2_decap_8 FILLER_37_1715 ();
 sg13g2_decap_4 FILLER_37_1722 ();
 sg13g2_decap_4 FILLER_37_1731 ();
 sg13g2_fill_2 FILLER_37_1735 ();
 sg13g2_decap_8 FILLER_37_1767 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_11 ();
 sg13g2_decap_4 FILLER_38_17 ();
 sg13g2_fill_1 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_32 ();
 sg13g2_fill_2 FILLER_38_36 ();
 sg13g2_fill_2 FILLER_38_51 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_decap_8 FILLER_38_78 ();
 sg13g2_fill_1 FILLER_38_85 ();
 sg13g2_decap_4 FILLER_38_95 ();
 sg13g2_fill_2 FILLER_38_104 ();
 sg13g2_fill_2 FILLER_38_120 ();
 sg13g2_fill_1 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_138 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_decap_4 FILLER_38_205 ();
 sg13g2_fill_1 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_decap_8 FILLER_38_484 ();
 sg13g2_decap_4 FILLER_38_491 ();
 sg13g2_decap_4 FILLER_38_516 ();
 sg13g2_fill_1 FILLER_38_520 ();
 sg13g2_fill_2 FILLER_38_542 ();
 sg13g2_decap_8 FILLER_38_599 ();
 sg13g2_decap_8 FILLER_38_606 ();
 sg13g2_decap_8 FILLER_38_613 ();
 sg13g2_decap_4 FILLER_38_620 ();
 sg13g2_decap_8 FILLER_38_653 ();
 sg13g2_fill_2 FILLER_38_660 ();
 sg13g2_fill_1 FILLER_38_692 ();
 sg13g2_decap_8 FILLER_38_698 ();
 sg13g2_fill_1 FILLER_38_710 ();
 sg13g2_fill_2 FILLER_38_715 ();
 sg13g2_decap_8 FILLER_38_727 ();
 sg13g2_fill_2 FILLER_38_734 ();
 sg13g2_fill_1 FILLER_38_736 ();
 sg13g2_decap_4 FILLER_38_745 ();
 sg13g2_fill_1 FILLER_38_749 ();
 sg13g2_fill_1 FILLER_38_771 ();
 sg13g2_fill_2 FILLER_38_786 ();
 sg13g2_fill_1 FILLER_38_792 ();
 sg13g2_fill_1 FILLER_38_811 ();
 sg13g2_decap_8 FILLER_38_817 ();
 sg13g2_decap_8 FILLER_38_824 ();
 sg13g2_decap_8 FILLER_38_831 ();
 sg13g2_decap_4 FILLER_38_838 ();
 sg13g2_decap_4 FILLER_38_846 ();
 sg13g2_fill_1 FILLER_38_850 ();
 sg13g2_fill_1 FILLER_38_862 ();
 sg13g2_fill_2 FILLER_38_896 ();
 sg13g2_decap_8 FILLER_38_919 ();
 sg13g2_fill_2 FILLER_38_926 ();
 sg13g2_decap_8 FILLER_38_932 ();
 sg13g2_fill_2 FILLER_38_939 ();
 sg13g2_fill_1 FILLER_38_941 ();
 sg13g2_fill_2 FILLER_38_947 ();
 sg13g2_decap_8 FILLER_38_974 ();
 sg13g2_fill_1 FILLER_38_981 ();
 sg13g2_decap_4 FILLER_38_991 ();
 sg13g2_decap_8 FILLER_38_1048 ();
 sg13g2_decap_8 FILLER_38_1055 ();
 sg13g2_fill_2 FILLER_38_1062 ();
 sg13g2_fill_1 FILLER_38_1064 ();
 sg13g2_fill_1 FILLER_38_1079 ();
 sg13g2_decap_4 FILLER_38_1083 ();
 sg13g2_fill_2 FILLER_38_1087 ();
 sg13g2_fill_2 FILLER_38_1094 ();
 sg13g2_decap_8 FILLER_38_1108 ();
 sg13g2_decap_8 FILLER_38_1115 ();
 sg13g2_fill_2 FILLER_38_1122 ();
 sg13g2_decap_4 FILLER_38_1133 ();
 sg13g2_fill_1 FILLER_38_1137 ();
 sg13g2_decap_4 FILLER_38_1147 ();
 sg13g2_fill_1 FILLER_38_1151 ();
 sg13g2_fill_2 FILLER_38_1156 ();
 sg13g2_fill_1 FILLER_38_1158 ();
 sg13g2_fill_2 FILLER_38_1162 ();
 sg13g2_fill_2 FILLER_38_1175 ();
 sg13g2_fill_2 FILLER_38_1182 ();
 sg13g2_decap_8 FILLER_38_1192 ();
 sg13g2_decap_4 FILLER_38_1199 ();
 sg13g2_fill_2 FILLER_38_1203 ();
 sg13g2_fill_2 FILLER_38_1233 ();
 sg13g2_fill_2 FILLER_38_1263 ();
 sg13g2_fill_2 FILLER_38_1291 ();
 sg13g2_fill_1 FILLER_38_1293 ();
 sg13g2_fill_1 FILLER_38_1303 ();
 sg13g2_decap_8 FILLER_38_1338 ();
 sg13g2_decap_4 FILLER_38_1345 ();
 sg13g2_decap_4 FILLER_38_1353 ();
 sg13g2_fill_1 FILLER_38_1357 ();
 sg13g2_decap_4 FILLER_38_1367 ();
 sg13g2_fill_2 FILLER_38_1371 ();
 sg13g2_decap_8 FILLER_38_1451 ();
 sg13g2_fill_2 FILLER_38_1458 ();
 sg13g2_fill_1 FILLER_38_1460 ();
 sg13g2_fill_2 FILLER_38_1469 ();
 sg13g2_decap_4 FILLER_38_1484 ();
 sg13g2_fill_1 FILLER_38_1488 ();
 sg13g2_decap_8 FILLER_38_1493 ();
 sg13g2_fill_2 FILLER_38_1500 ();
 sg13g2_decap_4 FILLER_38_1515 ();
 sg13g2_fill_1 FILLER_38_1527 ();
 sg13g2_fill_2 FILLER_38_1533 ();
 sg13g2_decap_8 FILLER_38_1547 ();
 sg13g2_decap_4 FILLER_38_1554 ();
 sg13g2_fill_1 FILLER_38_1558 ();
 sg13g2_decap_8 FILLER_38_1577 ();
 sg13g2_decap_4 FILLER_38_1584 ();
 sg13g2_fill_2 FILLER_38_1595 ();
 sg13g2_fill_1 FILLER_38_1597 ();
 sg13g2_decap_8 FILLER_38_1603 ();
 sg13g2_fill_2 FILLER_38_1610 ();
 sg13g2_fill_2 FILLER_38_1621 ();
 sg13g2_decap_8 FILLER_38_1638 ();
 sg13g2_fill_1 FILLER_38_1645 ();
 sg13g2_decap_4 FILLER_38_1669 ();
 sg13g2_fill_2 FILLER_38_1690 ();
 sg13g2_decap_8 FILLER_38_1718 ();
 sg13g2_fill_1 FILLER_38_1756 ();
 sg13g2_fill_1 FILLER_38_1762 ();
 sg13g2_decap_4 FILLER_38_1768 ();
 sg13g2_fill_2 FILLER_38_1772 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_11 ();
 sg13g2_fill_2 FILLER_39_21 ();
 sg13g2_fill_1 FILLER_39_32 ();
 sg13g2_fill_1 FILLER_39_37 ();
 sg13g2_decap_4 FILLER_39_46 ();
 sg13g2_fill_2 FILLER_39_50 ();
 sg13g2_decap_8 FILLER_39_60 ();
 sg13g2_decap_4 FILLER_39_67 ();
 sg13g2_decap_4 FILLER_39_97 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_decap_8 FILLER_39_116 ();
 sg13g2_fill_1 FILLER_39_123 ();
 sg13g2_decap_8 FILLER_39_164 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_fill_2 FILLER_39_182 ();
 sg13g2_decap_4 FILLER_39_201 ();
 sg13g2_fill_1 FILLER_39_205 ();
 sg13g2_decap_8 FILLER_39_222 ();
 sg13g2_fill_2 FILLER_39_229 ();
 sg13g2_fill_1 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_250 ();
 sg13g2_decap_4 FILLER_39_257 ();
 sg13g2_fill_1 FILLER_39_261 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_fill_2 FILLER_39_284 ();
 sg13g2_fill_1 FILLER_39_286 ();
 sg13g2_decap_8 FILLER_39_296 ();
 sg13g2_fill_1 FILLER_39_303 ();
 sg13g2_decap_4 FILLER_39_312 ();
 sg13g2_fill_1 FILLER_39_316 ();
 sg13g2_fill_2 FILLER_39_321 ();
 sg13g2_fill_1 FILLER_39_335 ();
 sg13g2_fill_2 FILLER_39_362 ();
 sg13g2_fill_1 FILLER_39_388 ();
 sg13g2_fill_2 FILLER_39_396 ();
 sg13g2_fill_1 FILLER_39_407 ();
 sg13g2_decap_4 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_459 ();
 sg13g2_decap_8 FILLER_39_466 ();
 sg13g2_decap_8 FILLER_39_473 ();
 sg13g2_decap_8 FILLER_39_480 ();
 sg13g2_fill_2 FILLER_39_492 ();
 sg13g2_fill_1 FILLER_39_494 ();
 sg13g2_decap_8 FILLER_39_516 ();
 sg13g2_decap_4 FILLER_39_523 ();
 sg13g2_fill_2 FILLER_39_527 ();
 sg13g2_fill_2 FILLER_39_547 ();
 sg13g2_fill_1 FILLER_39_594 ();
 sg13g2_decap_4 FILLER_39_616 ();
 sg13g2_fill_1 FILLER_39_620 ();
 sg13g2_fill_1 FILLER_39_625 ();
 sg13g2_decap_8 FILLER_39_661 ();
 sg13g2_decap_8 FILLER_39_668 ();
 sg13g2_decap_4 FILLER_39_675 ();
 sg13g2_fill_1 FILLER_39_683 ();
 sg13g2_decap_4 FILLER_39_734 ();
 sg13g2_decap_4 FILLER_39_741 ();
 sg13g2_fill_2 FILLER_39_787 ();
 sg13g2_fill_1 FILLER_39_794 ();
 sg13g2_fill_2 FILLER_39_840 ();
 sg13g2_fill_2 FILLER_39_866 ();
 sg13g2_fill_1 FILLER_39_876 ();
 sg13g2_fill_2 FILLER_39_888 ();
 sg13g2_decap_8 FILLER_39_899 ();
 sg13g2_fill_2 FILLER_39_906 ();
 sg13g2_decap_8 FILLER_39_912 ();
 sg13g2_fill_2 FILLER_39_919 ();
 sg13g2_fill_2 FILLER_39_952 ();
 sg13g2_decap_8 FILLER_39_958 ();
 sg13g2_fill_2 FILLER_39_965 ();
 sg13g2_decap_8 FILLER_39_972 ();
 sg13g2_decap_4 FILLER_39_979 ();
 sg13g2_fill_2 FILLER_39_983 ();
 sg13g2_fill_1 FILLER_39_990 ();
 sg13g2_fill_1 FILLER_39_1004 ();
 sg13g2_fill_2 FILLER_39_1018 ();
 sg13g2_fill_2 FILLER_39_1024 ();
 sg13g2_fill_1 FILLER_39_1026 ();
 sg13g2_fill_2 FILLER_39_1058 ();
 sg13g2_decap_4 FILLER_39_1064 ();
 sg13g2_fill_2 FILLER_39_1068 ();
 sg13g2_fill_1 FILLER_39_1074 ();
 sg13g2_decap_4 FILLER_39_1080 ();
 sg13g2_decap_4 FILLER_39_1088 ();
 sg13g2_fill_2 FILLER_39_1092 ();
 sg13g2_decap_8 FILLER_39_1133 ();
 sg13g2_fill_1 FILLER_39_1143 ();
 sg13g2_decap_8 FILLER_39_1175 ();
 sg13g2_decap_4 FILLER_39_1182 ();
 sg13g2_decap_8 FILLER_39_1201 ();
 sg13g2_decap_8 FILLER_39_1208 ();
 sg13g2_decap_8 FILLER_39_1215 ();
 sg13g2_decap_4 FILLER_39_1222 ();
 sg13g2_fill_1 FILLER_39_1226 ();
 sg13g2_decap_8 FILLER_39_1271 ();
 sg13g2_fill_2 FILLER_39_1278 ();
 sg13g2_fill_2 FILLER_39_1293 ();
 sg13g2_fill_1 FILLER_39_1299 ();
 sg13g2_fill_1 FILLER_39_1306 ();
 sg13g2_fill_2 FILLER_39_1314 ();
 sg13g2_fill_1 FILLER_39_1316 ();
 sg13g2_decap_8 FILLER_39_1321 ();
 sg13g2_decap_8 FILLER_39_1328 ();
 sg13g2_decap_8 FILLER_39_1335 ();
 sg13g2_fill_1 FILLER_39_1355 ();
 sg13g2_decap_8 FILLER_39_1390 ();
 sg13g2_decap_4 FILLER_39_1397 ();
 sg13g2_fill_1 FILLER_39_1401 ();
 sg13g2_fill_2 FILLER_39_1415 ();
 sg13g2_fill_1 FILLER_39_1417 ();
 sg13g2_decap_8 FILLER_39_1427 ();
 sg13g2_fill_1 FILLER_39_1434 ();
 sg13g2_decap_8 FILLER_39_1444 ();
 sg13g2_decap_4 FILLER_39_1451 ();
 sg13g2_fill_2 FILLER_39_1460 ();
 sg13g2_decap_8 FILLER_39_1486 ();
 sg13g2_decap_8 FILLER_39_1493 ();
 sg13g2_fill_2 FILLER_39_1522 ();
 sg13g2_decap_8 FILLER_39_1528 ();
 sg13g2_fill_2 FILLER_39_1535 ();
 sg13g2_decap_8 FILLER_39_1545 ();
 sg13g2_fill_1 FILLER_39_1552 ();
 sg13g2_fill_2 FILLER_39_1569 ();
 sg13g2_decap_8 FILLER_39_1586 ();
 sg13g2_decap_8 FILLER_39_1593 ();
 sg13g2_fill_1 FILLER_39_1600 ();
 sg13g2_decap_8 FILLER_39_1605 ();
 sg13g2_decap_8 FILLER_39_1612 ();
 sg13g2_decap_8 FILLER_39_1634 ();
 sg13g2_decap_8 FILLER_39_1641 ();
 sg13g2_fill_2 FILLER_39_1648 ();
 sg13g2_fill_2 FILLER_39_1667 ();
 sg13g2_fill_1 FILLER_39_1669 ();
 sg13g2_decap_8 FILLER_39_1674 ();
 sg13g2_fill_1 FILLER_39_1691 ();
 sg13g2_decap_8 FILLER_39_1697 ();
 sg13g2_decap_4 FILLER_39_1704 ();
 sg13g2_fill_1 FILLER_39_1708 ();
 sg13g2_decap_8 FILLER_39_1714 ();
 sg13g2_decap_8 FILLER_39_1726 ();
 sg13g2_fill_2 FILLER_39_1747 ();
 sg13g2_fill_1 FILLER_39_1749 ();
 sg13g2_fill_1 FILLER_39_1760 ();
 sg13g2_decap_8 FILLER_39_1766 ();
 sg13g2_fill_1 FILLER_39_1773 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_12 ();
 sg13g2_decap_4 FILLER_40_21 ();
 sg13g2_fill_1 FILLER_40_25 ();
 sg13g2_fill_1 FILLER_40_40 ();
 sg13g2_decap_8 FILLER_40_57 ();
 sg13g2_fill_2 FILLER_40_64 ();
 sg13g2_decap_4 FILLER_40_71 ();
 sg13g2_fill_2 FILLER_40_75 ();
 sg13g2_decap_4 FILLER_40_93 ();
 sg13g2_fill_2 FILLER_40_97 ();
 sg13g2_decap_8 FILLER_40_107 ();
 sg13g2_decap_8 FILLER_40_114 ();
 sg13g2_decap_8 FILLER_40_121 ();
 sg13g2_fill_2 FILLER_40_128 ();
 sg13g2_decap_8 FILLER_40_138 ();
 sg13g2_fill_2 FILLER_40_145 ();
 sg13g2_fill_1 FILLER_40_147 ();
 sg13g2_fill_1 FILLER_40_161 ();
 sg13g2_fill_2 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_188 ();
 sg13g2_fill_2 FILLER_40_195 ();
 sg13g2_fill_1 FILLER_40_197 ();
 sg13g2_fill_2 FILLER_40_209 ();
 sg13g2_fill_1 FILLER_40_211 ();
 sg13g2_fill_2 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_227 ();
 sg13g2_fill_1 FILLER_40_234 ();
 sg13g2_fill_2 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_291 ();
 sg13g2_decap_8 FILLER_40_298 ();
 sg13g2_decap_8 FILLER_40_305 ();
 sg13g2_fill_2 FILLER_40_312 ();
 sg13g2_fill_1 FILLER_40_314 ();
 sg13g2_fill_1 FILLER_40_336 ();
 sg13g2_fill_1 FILLER_40_345 ();
 sg13g2_fill_2 FILLER_40_349 ();
 sg13g2_fill_1 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_4 FILLER_40_490 ();
 sg13g2_fill_1 FILLER_40_494 ();
 sg13g2_decap_8 FILLER_40_498 ();
 sg13g2_fill_1 FILLER_40_531 ();
 sg13g2_fill_1 FILLER_40_546 ();
 sg13g2_fill_2 FILLER_40_571 ();
 sg13g2_decap_4 FILLER_40_612 ();
 sg13g2_fill_2 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_676 ();
 sg13g2_fill_2 FILLER_40_683 ();
 sg13g2_fill_1 FILLER_40_685 ();
 sg13g2_fill_2 FILLER_40_691 ();
 sg13g2_fill_2 FILLER_40_697 ();
 sg13g2_fill_1 FILLER_40_699 ();
 sg13g2_decap_4 FILLER_40_704 ();
 sg13g2_decap_4 FILLER_40_726 ();
 sg13g2_fill_1 FILLER_40_734 ();
 sg13g2_fill_2 FILLER_40_774 ();
 sg13g2_decap_4 FILLER_40_806 ();
 sg13g2_fill_2 FILLER_40_810 ();
 sg13g2_fill_1 FILLER_40_821 ();
 sg13g2_decap_8 FILLER_40_831 ();
 sg13g2_decap_8 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_873 ();
 sg13g2_decap_4 FILLER_40_924 ();
 sg13g2_decap_8 FILLER_40_953 ();
 sg13g2_decap_8 FILLER_40_960 ();
 sg13g2_fill_2 FILLER_40_967 ();
 sg13g2_fill_1 FILLER_40_969 ();
 sg13g2_decap_8 FILLER_40_978 ();
 sg13g2_fill_1 FILLER_40_1016 ();
 sg13g2_decap_8 FILLER_40_1040 ();
 sg13g2_decap_4 FILLER_40_1047 ();
 sg13g2_fill_1 FILLER_40_1051 ();
 sg13g2_decap_4 FILLER_40_1067 ();
 sg13g2_fill_1 FILLER_40_1071 ();
 sg13g2_decap_4 FILLER_40_1127 ();
 sg13g2_fill_1 FILLER_40_1131 ();
 sg13g2_fill_1 FILLER_40_1143 ();
 sg13g2_fill_2 FILLER_40_1170 ();
 sg13g2_fill_1 FILLER_40_1197 ();
 sg13g2_decap_4 FILLER_40_1202 ();
 sg13g2_fill_2 FILLER_40_1206 ();
 sg13g2_decap_8 FILLER_40_1213 ();
 sg13g2_fill_2 FILLER_40_1220 ();
 sg13g2_fill_1 FILLER_40_1235 ();
 sg13g2_decap_8 FILLER_40_1248 ();
 sg13g2_decap_4 FILLER_40_1255 ();
 sg13g2_decap_8 FILLER_40_1264 ();
 sg13g2_fill_1 FILLER_40_1271 ();
 sg13g2_decap_4 FILLER_40_1302 ();
 sg13g2_fill_1 FILLER_40_1306 ();
 sg13g2_fill_2 FILLER_40_1317 ();
 sg13g2_fill_2 FILLER_40_1325 ();
 sg13g2_fill_1 FILLER_40_1332 ();
 sg13g2_decap_4 FILLER_40_1338 ();
 sg13g2_fill_1 FILLER_40_1358 ();
 sg13g2_decap_4 FILLER_40_1368 ();
 sg13g2_fill_1 FILLER_40_1372 ();
 sg13g2_fill_1 FILLER_40_1408 ();
 sg13g2_decap_4 FILLER_40_1431 ();
 sg13g2_fill_2 FILLER_40_1435 ();
 sg13g2_fill_1 FILLER_40_1466 ();
 sg13g2_fill_2 FILLER_40_1472 ();
 sg13g2_fill_1 FILLER_40_1474 ();
 sg13g2_decap_4 FILLER_40_1495 ();
 sg13g2_fill_1 FILLER_40_1508 ();
 sg13g2_fill_1 FILLER_40_1514 ();
 sg13g2_fill_1 FILLER_40_1555 ();
 sg13g2_decap_4 FILLER_40_1564 ();
 sg13g2_fill_1 FILLER_40_1568 ();
 sg13g2_decap_8 FILLER_40_1582 ();
 sg13g2_decap_8 FILLER_40_1589 ();
 sg13g2_decap_8 FILLER_40_1596 ();
 sg13g2_decap_8 FILLER_40_1603 ();
 sg13g2_decap_8 FILLER_40_1610 ();
 sg13g2_decap_8 FILLER_40_1617 ();
 sg13g2_decap_8 FILLER_40_1624 ();
 sg13g2_decap_4 FILLER_40_1631 ();
 sg13g2_fill_1 FILLER_40_1635 ();
 sg13g2_decap_4 FILLER_40_1648 ();
 sg13g2_fill_1 FILLER_40_1652 ();
 sg13g2_decap_8 FILLER_40_1666 ();
 sg13g2_fill_2 FILLER_40_1673 ();
 sg13g2_fill_1 FILLER_40_1675 ();
 sg13g2_fill_2 FILLER_40_1692 ();
 sg13g2_decap_8 FILLER_40_1703 ();
 sg13g2_fill_2 FILLER_40_1710 ();
 sg13g2_fill_1 FILLER_40_1712 ();
 sg13g2_fill_1 FILLER_40_1736 ();
 sg13g2_fill_2 FILLER_40_1757 ();
 sg13g2_decap_8 FILLER_40_1764 ();
 sg13g2_fill_2 FILLER_40_1771 ();
 sg13g2_fill_1 FILLER_40_1773 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_39 ();
 sg13g2_decap_8 FILLER_41_76 ();
 sg13g2_decap_8 FILLER_41_83 ();
 sg13g2_decap_8 FILLER_41_99 ();
 sg13g2_decap_4 FILLER_41_106 ();
 sg13g2_fill_1 FILLER_41_121 ();
 sg13g2_decap_8 FILLER_41_130 ();
 sg13g2_decap_4 FILLER_41_137 ();
 sg13g2_fill_1 FILLER_41_141 ();
 sg13g2_fill_1 FILLER_41_175 ();
 sg13g2_fill_1 FILLER_41_202 ();
 sg13g2_decap_4 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_223 ();
 sg13g2_fill_1 FILLER_41_241 ();
 sg13g2_decap_4 FILLER_41_248 ();
 sg13g2_fill_1 FILLER_41_252 ();
 sg13g2_fill_2 FILLER_41_264 ();
 sg13g2_fill_1 FILLER_41_266 ();
 sg13g2_fill_1 FILLER_41_309 ();
 sg13g2_fill_2 FILLER_41_318 ();
 sg13g2_fill_1 FILLER_41_324 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_fill_2 FILLER_41_420 ();
 sg13g2_fill_2 FILLER_41_442 ();
 sg13g2_fill_2 FILLER_41_449 ();
 sg13g2_fill_1 FILLER_41_451 ();
 sg13g2_decap_4 FILLER_41_457 ();
 sg13g2_fill_2 FILLER_41_461 ();
 sg13g2_decap_8 FILLER_41_505 ();
 sg13g2_decap_8 FILLER_41_512 ();
 sg13g2_decap_4 FILLER_41_519 ();
 sg13g2_fill_2 FILLER_41_523 ();
 sg13g2_fill_2 FILLER_41_533 ();
 sg13g2_fill_1 FILLER_41_543 ();
 sg13g2_fill_2 FILLER_41_558 ();
 sg13g2_fill_2 FILLER_41_579 ();
 sg13g2_fill_1 FILLER_41_646 ();
 sg13g2_fill_1 FILLER_41_663 ();
 sg13g2_decap_4 FILLER_41_676 ();
 sg13g2_fill_1 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_691 ();
 sg13g2_decap_4 FILLER_41_700 ();
 sg13g2_fill_1 FILLER_41_704 ();
 sg13g2_decap_8 FILLER_41_710 ();
 sg13g2_decap_8 FILLER_41_717 ();
 sg13g2_decap_8 FILLER_41_724 ();
 sg13g2_decap_8 FILLER_41_731 ();
 sg13g2_decap_4 FILLER_41_738 ();
 sg13g2_fill_2 FILLER_41_742 ();
 sg13g2_fill_1 FILLER_41_762 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_4 FILLER_41_798 ();
 sg13g2_decap_4 FILLER_41_807 ();
 sg13g2_decap_4 FILLER_41_815 ();
 sg13g2_fill_1 FILLER_41_819 ();
 sg13g2_fill_1 FILLER_41_838 ();
 sg13g2_fill_1 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_849 ();
 sg13g2_decap_4 FILLER_41_856 ();
 sg13g2_fill_1 FILLER_41_860 ();
 sg13g2_decap_4 FILLER_41_866 ();
 sg13g2_decap_8 FILLER_41_874 ();
 sg13g2_decap_4 FILLER_41_881 ();
 sg13g2_fill_2 FILLER_41_885 ();
 sg13g2_decap_4 FILLER_41_891 ();
 sg13g2_fill_2 FILLER_41_895 ();
 sg13g2_fill_2 FILLER_41_901 ();
 sg13g2_fill_1 FILLER_41_903 ();
 sg13g2_fill_2 FILLER_41_916 ();
 sg13g2_fill_1 FILLER_41_918 ();
 sg13g2_decap_4 FILLER_41_929 ();
 sg13g2_fill_1 FILLER_41_933 ();
 sg13g2_decap_8 FILLER_41_943 ();
 sg13g2_decap_4 FILLER_41_950 ();
 sg13g2_fill_1 FILLER_41_954 ();
 sg13g2_decap_4 FILLER_41_967 ();
 sg13g2_decap_4 FILLER_41_979 ();
 sg13g2_fill_2 FILLER_41_996 ();
 sg13g2_fill_1 FILLER_41_998 ();
 sg13g2_decap_4 FILLER_41_1003 ();
 sg13g2_fill_2 FILLER_41_1011 ();
 sg13g2_fill_1 FILLER_41_1013 ();
 sg13g2_decap_4 FILLER_41_1026 ();
 sg13g2_fill_2 FILLER_41_1030 ();
 sg13g2_decap_8 FILLER_41_1036 ();
 sg13g2_decap_4 FILLER_41_1043 ();
 sg13g2_fill_2 FILLER_41_1047 ();
 sg13g2_fill_1 FILLER_41_1069 ();
 sg13g2_fill_1 FILLER_41_1078 ();
 sg13g2_fill_2 FILLER_41_1083 ();
 sg13g2_fill_1 FILLER_41_1085 ();
 sg13g2_fill_2 FILLER_41_1095 ();
 sg13g2_fill_1 FILLER_41_1097 ();
 sg13g2_fill_1 FILLER_41_1105 ();
 sg13g2_decap_8 FILLER_41_1109 ();
 sg13g2_decap_8 FILLER_41_1116 ();
 sg13g2_decap_4 FILLER_41_1123 ();
 sg13g2_fill_1 FILLER_41_1127 ();
 sg13g2_decap_4 FILLER_41_1132 ();
 sg13g2_fill_1 FILLER_41_1136 ();
 sg13g2_fill_1 FILLER_41_1150 ();
 sg13g2_fill_1 FILLER_41_1155 ();
 sg13g2_fill_2 FILLER_41_1218 ();
 sg13g2_fill_1 FILLER_41_1220 ();
 sg13g2_decap_8 FILLER_41_1236 ();
 sg13g2_decap_8 FILLER_41_1243 ();
 sg13g2_fill_1 FILLER_41_1250 ();
 sg13g2_fill_2 FILLER_41_1256 ();
 sg13g2_fill_1 FILLER_41_1258 ();
 sg13g2_fill_2 FILLER_41_1266 ();
 sg13g2_fill_1 FILLER_41_1268 ();
 sg13g2_decap_8 FILLER_41_1277 ();
 sg13g2_decap_8 FILLER_41_1284 ();
 sg13g2_decap_8 FILLER_41_1291 ();
 sg13g2_decap_8 FILLER_41_1298 ();
 sg13g2_decap_8 FILLER_41_1305 ();
 sg13g2_decap_8 FILLER_41_1312 ();
 sg13g2_decap_8 FILLER_41_1319 ();
 sg13g2_decap_8 FILLER_41_1326 ();
 sg13g2_decap_8 FILLER_41_1333 ();
 sg13g2_decap_8 FILLER_41_1344 ();
 sg13g2_decap_8 FILLER_41_1351 ();
 sg13g2_fill_1 FILLER_41_1358 ();
 sg13g2_decap_4 FILLER_41_1364 ();
 sg13g2_fill_1 FILLER_41_1368 ();
 sg13g2_decap_8 FILLER_41_1374 ();
 sg13g2_fill_2 FILLER_41_1381 ();
 sg13g2_fill_1 FILLER_41_1383 ();
 sg13g2_decap_8 FILLER_41_1429 ();
 sg13g2_decap_8 FILLER_41_1436 ();
 sg13g2_decap_4 FILLER_41_1443 ();
 sg13g2_fill_2 FILLER_41_1447 ();
 sg13g2_fill_1 FILLER_41_1458 ();
 sg13g2_fill_1 FILLER_41_1463 ();
 sg13g2_fill_2 FILLER_41_1474 ();
 sg13g2_fill_2 FILLER_41_1481 ();
 sg13g2_fill_2 FILLER_41_1491 ();
 sg13g2_decap_4 FILLER_41_1497 ();
 sg13g2_fill_2 FILLER_41_1501 ();
 sg13g2_decap_8 FILLER_41_1514 ();
 sg13g2_fill_1 FILLER_41_1521 ();
 sg13g2_fill_1 FILLER_41_1532 ();
 sg13g2_fill_1 FILLER_41_1538 ();
 sg13g2_fill_1 FILLER_41_1544 ();
 sg13g2_fill_2 FILLER_41_1553 ();
 sg13g2_decap_8 FILLER_41_1583 ();
 sg13g2_decap_8 FILLER_41_1590 ();
 sg13g2_decap_4 FILLER_41_1597 ();
 sg13g2_decap_8 FILLER_41_1648 ();
 sg13g2_decap_8 FILLER_41_1655 ();
 sg13g2_fill_2 FILLER_41_1662 ();
 sg13g2_decap_8 FILLER_41_1672 ();
 sg13g2_fill_2 FILLER_41_1679 ();
 sg13g2_fill_1 FILLER_41_1681 ();
 sg13g2_decap_4 FILLER_41_1698 ();
 sg13g2_fill_1 FILLER_41_1707 ();
 sg13g2_fill_2 FILLER_41_1725 ();
 sg13g2_fill_1 FILLER_41_1732 ();
 sg13g2_decap_8 FILLER_41_1764 ();
 sg13g2_fill_2 FILLER_41_1771 ();
 sg13g2_fill_1 FILLER_41_1773 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_14 ();
 sg13g2_fill_1 FILLER_42_16 ();
 sg13g2_decap_4 FILLER_42_21 ();
 sg13g2_fill_1 FILLER_42_25 ();
 sg13g2_fill_2 FILLER_42_36 ();
 sg13g2_fill_1 FILLER_42_38 ();
 sg13g2_fill_1 FILLER_42_43 ();
 sg13g2_fill_2 FILLER_42_49 ();
 sg13g2_fill_1 FILLER_42_51 ();
 sg13g2_fill_1 FILLER_42_57 ();
 sg13g2_decap_8 FILLER_42_65 ();
 sg13g2_fill_2 FILLER_42_72 ();
 sg13g2_decap_4 FILLER_42_79 ();
 sg13g2_fill_2 FILLER_42_83 ();
 sg13g2_fill_2 FILLER_42_90 ();
 sg13g2_fill_1 FILLER_42_92 ();
 sg13g2_fill_2 FILLER_42_102 ();
 sg13g2_fill_1 FILLER_42_104 ();
 sg13g2_decap_8 FILLER_42_131 ();
 sg13g2_fill_2 FILLER_42_138 ();
 sg13g2_fill_1 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_149 ();
 sg13g2_decap_4 FILLER_42_156 ();
 sg13g2_fill_2 FILLER_42_160 ();
 sg13g2_decap_8 FILLER_42_172 ();
 sg13g2_decap_4 FILLER_42_179 ();
 sg13g2_decap_8 FILLER_42_190 ();
 sg13g2_decap_8 FILLER_42_197 ();
 sg13g2_decap_8 FILLER_42_204 ();
 sg13g2_decap_8 FILLER_42_211 ();
 sg13g2_fill_2 FILLER_42_218 ();
 sg13g2_decap_8 FILLER_42_228 ();
 sg13g2_decap_4 FILLER_42_243 ();
 sg13g2_fill_1 FILLER_42_247 ();
 sg13g2_fill_1 FILLER_42_275 ();
 sg13g2_decap_8 FILLER_42_288 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_decap_4 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_313 ();
 sg13g2_decap_4 FILLER_42_320 ();
 sg13g2_fill_1 FILLER_42_341 ();
 sg13g2_fill_2 FILLER_42_355 ();
 sg13g2_fill_1 FILLER_42_364 ();
 sg13g2_fill_2 FILLER_42_369 ();
 sg13g2_fill_1 FILLER_42_383 ();
 sg13g2_decap_8 FILLER_42_418 ();
 sg13g2_decap_8 FILLER_42_425 ();
 sg13g2_decap_8 FILLER_42_432 ();
 sg13g2_decap_8 FILLER_42_439 ();
 sg13g2_decap_8 FILLER_42_446 ();
 sg13g2_decap_8 FILLER_42_453 ();
 sg13g2_decap_8 FILLER_42_460 ();
 sg13g2_decap_8 FILLER_42_467 ();
 sg13g2_decap_4 FILLER_42_474 ();
 sg13g2_fill_1 FILLER_42_478 ();
 sg13g2_decap_8 FILLER_42_484 ();
 sg13g2_decap_4 FILLER_42_491 ();
 sg13g2_fill_2 FILLER_42_505 ();
 sg13g2_fill_2 FILLER_42_579 ();
 sg13g2_fill_1 FILLER_42_625 ();
 sg13g2_fill_1 FILLER_42_636 ();
 sg13g2_fill_1 FILLER_42_650 ();
 sg13g2_decap_8 FILLER_42_682 ();
 sg13g2_fill_2 FILLER_42_689 ();
 sg13g2_fill_1 FILLER_42_691 ();
 sg13g2_decap_8 FILLER_42_720 ();
 sg13g2_decap_4 FILLER_42_727 ();
 sg13g2_fill_1 FILLER_42_735 ();
 sg13g2_fill_2 FILLER_42_744 ();
 sg13g2_fill_1 FILLER_42_751 ();
 sg13g2_fill_2 FILLER_42_786 ();
 sg13g2_fill_2 FILLER_42_796 ();
 sg13g2_fill_1 FILLER_42_798 ();
 sg13g2_fill_2 FILLER_42_812 ();
 sg13g2_fill_1 FILLER_42_814 ();
 sg13g2_fill_1 FILLER_42_819 ();
 sg13g2_fill_1 FILLER_42_826 ();
 sg13g2_fill_2 FILLER_42_837 ();
 sg13g2_decap_8 FILLER_42_857 ();
 sg13g2_decap_4 FILLER_42_864 ();
 sg13g2_fill_1 FILLER_42_868 ();
 sg13g2_decap_8 FILLER_42_884 ();
 sg13g2_fill_2 FILLER_42_891 ();
 sg13g2_fill_1 FILLER_42_893 ();
 sg13g2_decap_4 FILLER_42_925 ();
 sg13g2_decap_4 FILLER_42_933 ();
 sg13g2_decap_4 FILLER_42_942 ();
 sg13g2_fill_1 FILLER_42_946 ();
 sg13g2_decap_8 FILLER_42_983 ();
 sg13g2_fill_2 FILLER_42_990 ();
 sg13g2_decap_8 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_42_1035 ();
 sg13g2_decap_8 FILLER_42_1042 ();
 sg13g2_fill_2 FILLER_42_1049 ();
 sg13g2_fill_1 FILLER_42_1051 ();
 sg13g2_fill_1 FILLER_42_1055 ();
 sg13g2_decap_4 FILLER_42_1060 ();
 sg13g2_decap_8 FILLER_42_1209 ();
 sg13g2_decap_4 FILLER_42_1216 ();
 sg13g2_fill_1 FILLER_42_1220 ();
 sg13g2_decap_4 FILLER_42_1246 ();
 sg13g2_fill_1 FILLER_42_1275 ();
 sg13g2_decap_8 FILLER_42_1280 ();
 sg13g2_fill_2 FILLER_42_1287 ();
 sg13g2_decap_8 FILLER_42_1319 ();
 sg13g2_decap_4 FILLER_42_1326 ();
 sg13g2_fill_2 FILLER_42_1330 ();
 sg13g2_decap_4 FILLER_42_1363 ();
 sg13g2_fill_2 FILLER_42_1367 ();
 sg13g2_decap_8 FILLER_42_1374 ();
 sg13g2_decap_4 FILLER_42_1381 ();
 sg13g2_fill_2 FILLER_42_1385 ();
 sg13g2_fill_2 FILLER_42_1412 ();
 sg13g2_fill_1 FILLER_42_1414 ();
 sg13g2_fill_1 FILLER_42_1419 ();
 sg13g2_fill_2 FILLER_42_1428 ();
 sg13g2_fill_2 FILLER_42_1435 ();
 sg13g2_fill_1 FILLER_42_1437 ();
 sg13g2_fill_1 FILLER_42_1451 ();
 sg13g2_fill_2 FILLER_42_1457 ();
 sg13g2_fill_1 FILLER_42_1459 ();
 sg13g2_decap_8 FILLER_42_1479 ();
 sg13g2_decap_8 FILLER_42_1486 ();
 sg13g2_decap_8 FILLER_42_1493 ();
 sg13g2_decap_8 FILLER_42_1500 ();
 sg13g2_fill_2 FILLER_42_1516 ();
 sg13g2_fill_1 FILLER_42_1518 ();
 sg13g2_fill_2 FILLER_42_1533 ();
 sg13g2_fill_1 FILLER_42_1535 ();
 sg13g2_decap_8 FILLER_42_1549 ();
 sg13g2_fill_2 FILLER_42_1572 ();
 sg13g2_decap_4 FILLER_42_1605 ();
 sg13g2_decap_8 FILLER_42_1614 ();
 sg13g2_decap_4 FILLER_42_1621 ();
 sg13g2_fill_1 FILLER_42_1660 ();
 sg13g2_fill_1 FILLER_42_1670 ();
 sg13g2_fill_1 FILLER_42_1678 ();
 sg13g2_fill_1 FILLER_42_1687 ();
 sg13g2_decap_4 FILLER_42_1694 ();
 sg13g2_fill_1 FILLER_42_1698 ();
 sg13g2_fill_2 FILLER_42_1703 ();
 sg13g2_fill_2 FILLER_42_1711 ();
 sg13g2_fill_2 FILLER_42_1726 ();
 sg13g2_fill_2 FILLER_42_1742 ();
 sg13g2_decap_8 FILLER_42_1756 ();
 sg13g2_decap_8 FILLER_42_1763 ();
 sg13g2_decap_4 FILLER_42_1770 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_11 ();
 sg13g2_fill_2 FILLER_43_15 ();
 sg13g2_fill_2 FILLER_43_45 ();
 sg13g2_decap_4 FILLER_43_65 ();
 sg13g2_fill_2 FILLER_43_78 ();
 sg13g2_decap_8 FILLER_43_87 ();
 sg13g2_fill_1 FILLER_43_94 ();
 sg13g2_decap_4 FILLER_43_103 ();
 sg13g2_fill_1 FILLER_43_107 ();
 sg13g2_fill_1 FILLER_43_128 ();
 sg13g2_decap_4 FILLER_43_137 ();
 sg13g2_fill_2 FILLER_43_149 ();
 sg13g2_fill_1 FILLER_43_151 ();
 sg13g2_fill_2 FILLER_43_156 ();
 sg13g2_fill_2 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_165 ();
 sg13g2_fill_2 FILLER_43_176 ();
 sg13g2_fill_1 FILLER_43_178 ();
 sg13g2_fill_2 FILLER_43_201 ();
 sg13g2_fill_1 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_233 ();
 sg13g2_decap_8 FILLER_43_240 ();
 sg13g2_decap_4 FILLER_43_247 ();
 sg13g2_decap_4 FILLER_43_291 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_4 FILLER_43_308 ();
 sg13g2_fill_2 FILLER_43_312 ();
 sg13g2_fill_1 FILLER_43_342 ();
 sg13g2_decap_8 FILLER_43_388 ();
 sg13g2_fill_2 FILLER_43_395 ();
 sg13g2_fill_1 FILLER_43_397 ();
 sg13g2_decap_8 FILLER_43_405 ();
 sg13g2_fill_2 FILLER_43_412 ();
 sg13g2_fill_2 FILLER_43_418 ();
 sg13g2_decap_4 FILLER_43_424 ();
 sg13g2_fill_1 FILLER_43_428 ();
 sg13g2_decap_8 FILLER_43_465 ();
 sg13g2_decap_8 FILLER_43_472 ();
 sg13g2_decap_4 FILLER_43_479 ();
 sg13g2_fill_1 FILLER_43_483 ();
 sg13g2_decap_4 FILLER_43_489 ();
 sg13g2_fill_1 FILLER_43_493 ();
 sg13g2_fill_2 FILLER_43_498 ();
 sg13g2_fill_1 FILLER_43_500 ();
 sg13g2_decap_8 FILLER_43_548 ();
 sg13g2_decap_4 FILLER_43_569 ();
 sg13g2_fill_2 FILLER_43_573 ();
 sg13g2_fill_1 FILLER_43_584 ();
 sg13g2_fill_2 FILLER_43_601 ();
 sg13g2_fill_2 FILLER_43_669 ();
 sg13g2_fill_1 FILLER_43_701 ();
 sg13g2_fill_2 FILLER_43_706 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_8 FILLER_43_725 ();
 sg13g2_decap_4 FILLER_43_732 ();
 sg13g2_fill_2 FILLER_43_823 ();
 sg13g2_fill_2 FILLER_43_869 ();
 sg13g2_decap_8 FILLER_43_885 ();
 sg13g2_decap_4 FILLER_43_892 ();
 sg13g2_fill_1 FILLER_43_896 ();
 sg13g2_decap_8 FILLER_43_905 ();
 sg13g2_decap_8 FILLER_43_922 ();
 sg13g2_fill_2 FILLER_43_929 ();
 sg13g2_fill_1 FILLER_43_931 ();
 sg13g2_decap_4 FILLER_43_936 ();
 sg13g2_fill_2 FILLER_43_940 ();
 sg13g2_decap_4 FILLER_43_972 ();
 sg13g2_decap_8 FILLER_43_1033 ();
 sg13g2_decap_8 FILLER_43_1040 ();
 sg13g2_decap_4 FILLER_43_1047 ();
 sg13g2_fill_2 FILLER_43_1051 ();
 sg13g2_decap_4 FILLER_43_1057 ();
 sg13g2_fill_2 FILLER_43_1061 ();
 sg13g2_fill_2 FILLER_43_1075 ();
 sg13g2_fill_2 FILLER_43_1086 ();
 sg13g2_fill_1 FILLER_43_1088 ();
 sg13g2_decap_8 FILLER_43_1102 ();
 sg13g2_fill_1 FILLER_43_1109 ();
 sg13g2_decap_4 FILLER_43_1115 ();
 sg13g2_fill_1 FILLER_43_1119 ();
 sg13g2_decap_8 FILLER_43_1123 ();
 sg13g2_fill_2 FILLER_43_1130 ();
 sg13g2_fill_1 FILLER_43_1132 ();
 sg13g2_fill_2 FILLER_43_1180 ();
 sg13g2_fill_1 FILLER_43_1182 ();
 sg13g2_decap_8 FILLER_43_1204 ();
 sg13g2_fill_1 FILLER_43_1211 ();
 sg13g2_decap_8 FILLER_43_1240 ();
 sg13g2_decap_4 FILLER_43_1247 ();
 sg13g2_fill_2 FILLER_43_1251 ();
 sg13g2_fill_1 FILLER_43_1258 ();
 sg13g2_fill_1 FILLER_43_1268 ();
 sg13g2_decap_8 FILLER_43_1295 ();
 sg13g2_decap_8 FILLER_43_1302 ();
 sg13g2_decap_4 FILLER_43_1309 ();
 sg13g2_decap_8 FILLER_43_1318 ();
 sg13g2_decap_4 FILLER_43_1325 ();
 sg13g2_fill_1 FILLER_43_1329 ();
 sg13g2_decap_4 FILLER_43_1351 ();
 sg13g2_fill_2 FILLER_43_1359 ();
 sg13g2_decap_8 FILLER_43_1387 ();
 sg13g2_decap_4 FILLER_43_1394 ();
 sg13g2_fill_1 FILLER_43_1398 ();
 sg13g2_decap_8 FILLER_43_1403 ();
 sg13g2_decap_8 FILLER_43_1410 ();
 sg13g2_decap_8 FILLER_43_1417 ();
 sg13g2_fill_2 FILLER_43_1424 ();
 sg13g2_fill_2 FILLER_43_1438 ();
 sg13g2_fill_1 FILLER_43_1449 ();
 sg13g2_fill_2 FILLER_43_1454 ();
 sg13g2_fill_1 FILLER_43_1460 ();
 sg13g2_fill_2 FILLER_43_1487 ();
 sg13g2_decap_8 FILLER_43_1493 ();
 sg13g2_decap_4 FILLER_43_1500 ();
 sg13g2_fill_1 FILLER_43_1504 ();
 sg13g2_decap_4 FILLER_43_1526 ();
 sg13g2_fill_2 FILLER_43_1530 ();
 sg13g2_decap_8 FILLER_43_1550 ();
 sg13g2_fill_1 FILLER_43_1557 ();
 sg13g2_decap_4 FILLER_43_1570 ();
 sg13g2_fill_2 FILLER_43_1582 ();
 sg13g2_decap_4 FILLER_43_1591 ();
 sg13g2_fill_2 FILLER_43_1595 ();
 sg13g2_fill_2 FILLER_43_1601 ();
 sg13g2_fill_1 FILLER_43_1603 ();
 sg13g2_decap_8 FILLER_43_1609 ();
 sg13g2_fill_1 FILLER_43_1616 ();
 sg13g2_decap_4 FILLER_43_1621 ();
 sg13g2_decap_8 FILLER_43_1640 ();
 sg13g2_fill_2 FILLER_43_1647 ();
 sg13g2_fill_1 FILLER_43_1657 ();
 sg13g2_fill_1 FILLER_43_1666 ();
 sg13g2_fill_1 FILLER_43_1689 ();
 sg13g2_fill_2 FILLER_43_1700 ();
 sg13g2_fill_2 FILLER_43_1720 ();
 sg13g2_fill_2 FILLER_43_1733 ();
 sg13g2_fill_2 FILLER_43_1739 ();
 sg13g2_fill_1 FILLER_43_1753 ();
 sg13g2_decap_8 FILLER_43_1758 ();
 sg13g2_decap_8 FILLER_43_1765 ();
 sg13g2_fill_2 FILLER_43_1772 ();
 sg13g2_decap_8 FILLER_44_30 ();
 sg13g2_fill_1 FILLER_44_37 ();
 sg13g2_fill_1 FILLER_44_43 ();
 sg13g2_fill_1 FILLER_44_54 ();
 sg13g2_fill_2 FILLER_44_69 ();
 sg13g2_fill_1 FILLER_44_71 ();
 sg13g2_decap_8 FILLER_44_83 ();
 sg13g2_decap_4 FILLER_44_95 ();
 sg13g2_fill_1 FILLER_44_107 ();
 sg13g2_fill_2 FILLER_44_116 ();
 sg13g2_fill_2 FILLER_44_132 ();
 sg13g2_fill_1 FILLER_44_134 ();
 sg13g2_fill_1 FILLER_44_158 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_fill_2 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_192 ();
 sg13g2_fill_2 FILLER_44_199 ();
 sg13g2_fill_2 FILLER_44_232 ();
 sg13g2_decap_4 FILLER_44_255 ();
 sg13g2_fill_1 FILLER_44_259 ();
 sg13g2_decap_4 FILLER_44_268 ();
 sg13g2_fill_1 FILLER_44_272 ();
 sg13g2_decap_8 FILLER_44_278 ();
 sg13g2_decap_8 FILLER_44_285 ();
 sg13g2_decap_4 FILLER_44_292 ();
 sg13g2_fill_2 FILLER_44_300 ();
 sg13g2_fill_2 FILLER_44_310 ();
 sg13g2_fill_1 FILLER_44_312 ();
 sg13g2_fill_1 FILLER_44_348 ();
 sg13g2_fill_1 FILLER_44_355 ();
 sg13g2_fill_1 FILLER_44_394 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_fill_1 FILLER_44_458 ();
 sg13g2_fill_2 FILLER_44_520 ();
 sg13g2_decap_4 FILLER_44_544 ();
 sg13g2_fill_1 FILLER_44_548 ();
 sg13g2_fill_1 FILLER_44_554 ();
 sg13g2_decap_8 FILLER_44_572 ();
 sg13g2_fill_1 FILLER_44_579 ();
 sg13g2_fill_1 FILLER_44_593 ();
 sg13g2_fill_2 FILLER_44_599 ();
 sg13g2_fill_1 FILLER_44_610 ();
 sg13g2_fill_2 FILLER_44_632 ();
 sg13g2_fill_2 FILLER_44_640 ();
 sg13g2_fill_2 FILLER_44_664 ();
 sg13g2_decap_8 FILLER_44_701 ();
 sg13g2_decap_4 FILLER_44_708 ();
 sg13g2_fill_2 FILLER_44_712 ();
 sg13g2_fill_2 FILLER_44_740 ();
 sg13g2_fill_1 FILLER_44_742 ();
 sg13g2_fill_2 FILLER_44_760 ();
 sg13g2_fill_2 FILLER_44_765 ();
 sg13g2_fill_2 FILLER_44_781 ();
 sg13g2_fill_1 FILLER_44_822 ();
 sg13g2_fill_2 FILLER_44_828 ();
 sg13g2_fill_2 FILLER_44_842 ();
 sg13g2_decap_4 FILLER_44_852 ();
 sg13g2_fill_2 FILLER_44_856 ();
 sg13g2_fill_2 FILLER_44_874 ();
 sg13g2_decap_4 FILLER_44_881 ();
 sg13g2_decap_4 FILLER_44_898 ();
 sg13g2_fill_2 FILLER_44_902 ();
 sg13g2_decap_4 FILLER_44_926 ();
 sg13g2_decap_8 FILLER_44_977 ();
 sg13g2_decap_8 FILLER_44_988 ();
 sg13g2_fill_2 FILLER_44_995 ();
 sg13g2_decap_4 FILLER_44_1002 ();
 sg13g2_fill_1 FILLER_44_1006 ();
 sg13g2_decap_8 FILLER_44_1031 ();
 sg13g2_decap_8 FILLER_44_1038 ();
 sg13g2_fill_1 FILLER_44_1045 ();
 sg13g2_decap_4 FILLER_44_1059 ();
 sg13g2_fill_1 FILLER_44_1068 ();
 sg13g2_decap_4 FILLER_44_1141 ();
 sg13g2_fill_1 FILLER_44_1169 ();
 sg13g2_decap_8 FILLER_44_1234 ();
 sg13g2_decap_4 FILLER_44_1241 ();
 sg13g2_fill_1 FILLER_44_1245 ();
 sg13g2_fill_1 FILLER_44_1258 ();
 sg13g2_fill_1 FILLER_44_1269 ();
 sg13g2_fill_2 FILLER_44_1281 ();
 sg13g2_decap_8 FILLER_44_1299 ();
 sg13g2_decap_8 FILLER_44_1306 ();
 sg13g2_decap_8 FILLER_44_1313 ();
 sg13g2_decap_8 FILLER_44_1320 ();
 sg13g2_decap_8 FILLER_44_1327 ();
 sg13g2_decap_4 FILLER_44_1343 ();
 sg13g2_decap_4 FILLER_44_1356 ();
 sg13g2_decap_8 FILLER_44_1402 ();
 sg13g2_decap_8 FILLER_44_1409 ();
 sg13g2_decap_4 FILLER_44_1416 ();
 sg13g2_fill_1 FILLER_44_1420 ();
 sg13g2_decap_8 FILLER_44_1456 ();
 sg13g2_decap_4 FILLER_44_1463 ();
 sg13g2_fill_1 FILLER_44_1467 ();
 sg13g2_fill_2 FILLER_44_1476 ();
 sg13g2_fill_2 FILLER_44_1482 ();
 sg13g2_fill_1 FILLER_44_1484 ();
 sg13g2_fill_2 FILLER_44_1506 ();
 sg13g2_fill_1 FILLER_44_1508 ();
 sg13g2_fill_2 FILLER_44_1517 ();
 sg13g2_decap_8 FILLER_44_1523 ();
 sg13g2_decap_4 FILLER_44_1530 ();
 sg13g2_fill_1 FILLER_44_1534 ();
 sg13g2_fill_2 FILLER_44_1552 ();
 sg13g2_fill_1 FILLER_44_1554 ();
 sg13g2_fill_1 FILLER_44_1567 ();
 sg13g2_decap_8 FILLER_44_1572 ();
 sg13g2_decap_8 FILLER_44_1579 ();
 sg13g2_fill_1 FILLER_44_1586 ();
 sg13g2_fill_1 FILLER_44_1592 ();
 sg13g2_decap_8 FILLER_44_1615 ();
 sg13g2_decap_4 FILLER_44_1622 ();
 sg13g2_fill_1 FILLER_44_1646 ();
 sg13g2_fill_2 FILLER_44_1656 ();
 sg13g2_decap_8 FILLER_44_1668 ();
 sg13g2_decap_8 FILLER_44_1675 ();
 sg13g2_decap_8 FILLER_44_1682 ();
 sg13g2_fill_2 FILLER_44_1689 ();
 sg13g2_fill_1 FILLER_44_1691 ();
 sg13g2_fill_1 FILLER_44_1710 ();
 sg13g2_fill_2 FILLER_44_1719 ();
 sg13g2_fill_1 FILLER_44_1743 ();
 sg13g2_fill_1 FILLER_44_1755 ();
 sg13g2_decap_8 FILLER_44_1763 ();
 sg13g2_decap_4 FILLER_44_1770 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_11 ();
 sg13g2_decap_8 FILLER_45_18 ();
 sg13g2_decap_4 FILLER_45_25 ();
 sg13g2_fill_1 FILLER_45_62 ();
 sg13g2_fill_1 FILLER_45_94 ();
 sg13g2_fill_2 FILLER_45_116 ();
 sg13g2_decap_8 FILLER_45_130 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_fill_2 FILLER_45_175 ();
 sg13g2_fill_1 FILLER_45_177 ();
 sg13g2_decap_8 FILLER_45_190 ();
 sg13g2_decap_8 FILLER_45_197 ();
 sg13g2_fill_2 FILLER_45_204 ();
 sg13g2_decap_8 FILLER_45_214 ();
 sg13g2_decap_4 FILLER_45_221 ();
 sg13g2_fill_2 FILLER_45_230 ();
 sg13g2_fill_1 FILLER_45_232 ();
 sg13g2_decap_8 FILLER_45_237 ();
 sg13g2_decap_8 FILLER_45_244 ();
 sg13g2_fill_2 FILLER_45_251 ();
 sg13g2_fill_1 FILLER_45_274 ();
 sg13g2_fill_2 FILLER_45_280 ();
 sg13g2_fill_1 FILLER_45_282 ();
 sg13g2_decap_4 FILLER_45_289 ();
 sg13g2_decap_4 FILLER_45_297 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_fill_1 FILLER_45_307 ();
 sg13g2_fill_1 FILLER_45_316 ();
 sg13g2_fill_1 FILLER_45_322 ();
 sg13g2_fill_1 FILLER_45_328 ();
 sg13g2_fill_1 FILLER_45_359 ();
 sg13g2_fill_2 FILLER_45_390 ();
 sg13g2_decap_4 FILLER_45_396 ();
 sg13g2_decap_8 FILLER_45_451 ();
 sg13g2_decap_8 FILLER_45_458 ();
 sg13g2_decap_4 FILLER_45_465 ();
 sg13g2_fill_1 FILLER_45_469 ();
 sg13g2_decap_4 FILLER_45_516 ();
 sg13g2_decap_8 FILLER_45_538 ();
 sg13g2_decap_8 FILLER_45_545 ();
 sg13g2_fill_2 FILLER_45_556 ();
 sg13g2_decap_4 FILLER_45_567 ();
 sg13g2_fill_1 FILLER_45_571 ();
 sg13g2_fill_1 FILLER_45_577 ();
 sg13g2_fill_2 FILLER_45_582 ();
 sg13g2_fill_1 FILLER_45_589 ();
 sg13g2_fill_2 FILLER_45_604 ();
 sg13g2_fill_2 FILLER_45_617 ();
 sg13g2_fill_2 FILLER_45_665 ();
 sg13g2_decap_4 FILLER_45_703 ();
 sg13g2_fill_1 FILLER_45_707 ();
 sg13g2_fill_1 FILLER_45_721 ();
 sg13g2_decap_8 FILLER_45_727 ();
 sg13g2_fill_1 FILLER_45_734 ();
 sg13g2_fill_1 FILLER_45_739 ();
 sg13g2_fill_1 FILLER_45_745 ();
 sg13g2_fill_2 FILLER_45_760 ();
 sg13g2_fill_2 FILLER_45_773 ();
 sg13g2_fill_1 FILLER_45_775 ();
 sg13g2_fill_1 FILLER_45_781 ();
 sg13g2_fill_1 FILLER_45_791 ();
 sg13g2_decap_4 FILLER_45_796 ();
 sg13g2_fill_2 FILLER_45_800 ();
 sg13g2_fill_2 FILLER_45_822 ();
 sg13g2_decap_8 FILLER_45_846 ();
 sg13g2_decap_4 FILLER_45_913 ();
 sg13g2_fill_1 FILLER_45_917 ();
 sg13g2_decap_8 FILLER_45_939 ();
 sg13g2_decap_8 FILLER_45_946 ();
 sg13g2_decap_4 FILLER_45_953 ();
 sg13g2_fill_1 FILLER_45_957 ();
 sg13g2_decap_8 FILLER_45_979 ();
 sg13g2_decap_8 FILLER_45_986 ();
 sg13g2_decap_4 FILLER_45_993 ();
 sg13g2_fill_1 FILLER_45_997 ();
 sg13g2_decap_8 FILLER_45_1035 ();
 sg13g2_decap_8 FILLER_45_1042 ();
 sg13g2_decap_8 FILLER_45_1049 ();
 sg13g2_decap_4 FILLER_45_1056 ();
 sg13g2_fill_2 FILLER_45_1060 ();
 sg13g2_decap_4 FILLER_45_1067 ();
 sg13g2_decap_8 FILLER_45_1075 ();
 sg13g2_decap_8 FILLER_45_1082 ();
 sg13g2_fill_1 FILLER_45_1089 ();
 sg13g2_fill_1 FILLER_45_1094 ();
 sg13g2_fill_2 FILLER_45_1099 ();
 sg13g2_decap_4 FILLER_45_1136 ();
 sg13g2_fill_2 FILLER_45_1140 ();
 sg13g2_decap_8 FILLER_45_1154 ();
 sg13g2_fill_1 FILLER_45_1161 ();
 sg13g2_decap_4 FILLER_45_1219 ();
 sg13g2_fill_1 FILLER_45_1258 ();
 sg13g2_decap_4 FILLER_45_1328 ();
 sg13g2_fill_2 FILLER_45_1332 ();
 sg13g2_decap_4 FILLER_45_1339 ();
 sg13g2_fill_1 FILLER_45_1362 ();
 sg13g2_decap_8 FILLER_45_1408 ();
 sg13g2_fill_2 FILLER_45_1420 ();
 sg13g2_fill_1 FILLER_45_1422 ();
 sg13g2_fill_2 FILLER_45_1439 ();
 sg13g2_fill_2 FILLER_45_1446 ();
 sg13g2_fill_2 FILLER_45_1464 ();
 sg13g2_fill_2 FILLER_45_1472 ();
 sg13g2_fill_2 FILLER_45_1482 ();
 sg13g2_fill_2 FILLER_45_1488 ();
 sg13g2_fill_1 FILLER_45_1490 ();
 sg13g2_fill_2 FILLER_45_1499 ();
 sg13g2_fill_1 FILLER_45_1501 ();
 sg13g2_decap_8 FILLER_45_1523 ();
 sg13g2_fill_2 FILLER_45_1530 ();
 sg13g2_fill_1 FILLER_45_1532 ();
 sg13g2_fill_2 FILLER_45_1543 ();
 sg13g2_decap_4 FILLER_45_1574 ();
 sg13g2_decap_4 FILLER_45_1604 ();
 sg13g2_decap_8 FILLER_45_1613 ();
 sg13g2_fill_1 FILLER_45_1642 ();
 sg13g2_decap_4 FILLER_45_1656 ();
 sg13g2_fill_2 FILLER_45_1660 ();
 sg13g2_decap_4 FILLER_45_1666 ();
 sg13g2_fill_1 FILLER_45_1670 ();
 sg13g2_decap_8 FILLER_45_1676 ();
 sg13g2_decap_8 FILLER_45_1683 ();
 sg13g2_fill_2 FILLER_45_1694 ();
 sg13g2_fill_1 FILLER_45_1696 ();
 sg13g2_fill_2 FILLER_45_1722 ();
 sg13g2_fill_1 FILLER_45_1734 ();
 sg13g2_fill_1 FILLER_45_1751 ();
 sg13g2_fill_1 FILLER_45_1757 ();
 sg13g2_decap_8 FILLER_45_1763 ();
 sg13g2_decap_4 FILLER_45_1770 ();
 sg13g2_decap_8 FILLER_46_26 ();
 sg13g2_decap_8 FILLER_46_37 ();
 sg13g2_fill_2 FILLER_46_44 ();
 sg13g2_fill_1 FILLER_46_46 ();
 sg13g2_fill_2 FILLER_46_60 ();
 sg13g2_fill_2 FILLER_46_65 ();
 sg13g2_fill_1 FILLER_46_67 ();
 sg13g2_fill_1 FILLER_46_72 ();
 sg13g2_fill_2 FILLER_46_86 ();
 sg13g2_fill_1 FILLER_46_88 ();
 sg13g2_decap_8 FILLER_46_132 ();
 sg13g2_decap_8 FILLER_46_176 ();
 sg13g2_decap_8 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_190 ();
 sg13g2_decap_8 FILLER_46_195 ();
 sg13g2_decap_4 FILLER_46_206 ();
 sg13g2_decap_8 FILLER_46_223 ();
 sg13g2_fill_1 FILLER_46_234 ();
 sg13g2_fill_2 FILLER_46_239 ();
 sg13g2_fill_1 FILLER_46_241 ();
 sg13g2_fill_2 FILLER_46_258 ();
 sg13g2_fill_2 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_283 ();
 sg13g2_decap_4 FILLER_46_301 ();
 sg13g2_fill_1 FILLER_46_305 ();
 sg13g2_decap_8 FILLER_46_314 ();
 sg13g2_decap_4 FILLER_46_321 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_fill_2 FILLER_46_344 ();
 sg13g2_fill_1 FILLER_46_354 ();
 sg13g2_fill_1 FILLER_46_363 ();
 sg13g2_decap_4 FILLER_46_401 ();
 sg13g2_fill_2 FILLER_46_417 ();
 sg13g2_decap_8 FILLER_46_454 ();
 sg13g2_decap_4 FILLER_46_461 ();
 sg13g2_fill_1 FILLER_46_465 ();
 sg13g2_decap_8 FILLER_46_487 ();
 sg13g2_fill_1 FILLER_46_494 ();
 sg13g2_decap_8 FILLER_46_516 ();
 sg13g2_decap_8 FILLER_46_523 ();
 sg13g2_decap_4 FILLER_46_530 ();
 sg13g2_decap_4 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_583 ();
 sg13g2_fill_2 FILLER_46_590 ();
 sg13g2_fill_2 FILLER_46_606 ();
 sg13g2_fill_1 FILLER_46_629 ();
 sg13g2_fill_1 FILLER_46_648 ();
 sg13g2_fill_1 FILLER_46_653 ();
 sg13g2_fill_1 FILLER_46_660 ();
 sg13g2_fill_2 FILLER_46_680 ();
 sg13g2_decap_4 FILLER_46_690 ();
 sg13g2_fill_1 FILLER_46_694 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_4 FILLER_46_714 ();
 sg13g2_fill_2 FILLER_46_718 ();
 sg13g2_fill_2 FILLER_46_728 ();
 sg13g2_fill_1 FILLER_46_730 ();
 sg13g2_fill_2 FILLER_46_757 ();
 sg13g2_decap_8 FILLER_46_802 ();
 sg13g2_fill_1 FILLER_46_817 ();
 sg13g2_fill_1 FILLER_46_830 ();
 sg13g2_decap_4 FILLER_46_838 ();
 sg13g2_fill_1 FILLER_46_842 ();
 sg13g2_decap_4 FILLER_46_848 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_fill_1 FILLER_46_862 ();
 sg13g2_fill_2 FILLER_46_871 ();
 sg13g2_fill_1 FILLER_46_877 ();
 sg13g2_decap_8 FILLER_46_900 ();
 sg13g2_decap_4 FILLER_46_937 ();
 sg13g2_decap_8 FILLER_46_973 ();
 sg13g2_fill_1 FILLER_46_980 ();
 sg13g2_decap_8 FILLER_46_999 ();
 sg13g2_fill_2 FILLER_46_1006 ();
 sg13g2_decap_8 FILLER_46_1012 ();
 sg13g2_fill_2 FILLER_46_1019 ();
 sg13g2_fill_1 FILLER_46_1021 ();
 sg13g2_fill_2 FILLER_46_1026 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_decap_4 FILLER_46_1046 ();
 sg13g2_fill_2 FILLER_46_1050 ();
 sg13g2_decap_4 FILLER_46_1055 ();
 sg13g2_fill_1 FILLER_46_1059 ();
 sg13g2_decap_4 FILLER_46_1075 ();
 sg13g2_fill_1 FILLER_46_1079 ();
 sg13g2_decap_8 FILLER_46_1096 ();
 sg13g2_decap_4 FILLER_46_1103 ();
 sg13g2_fill_1 FILLER_46_1107 ();
 sg13g2_decap_4 FILLER_46_1113 ();
 sg13g2_decap_8 FILLER_46_1121 ();
 sg13g2_decap_8 FILLER_46_1133 ();
 sg13g2_decap_4 FILLER_46_1140 ();
 sg13g2_fill_1 FILLER_46_1144 ();
 sg13g2_decap_8 FILLER_46_1148 ();
 sg13g2_decap_8 FILLER_46_1155 ();
 sg13g2_fill_1 FILLER_46_1197 ();
 sg13g2_fill_1 FILLER_46_1258 ();
 sg13g2_fill_2 FILLER_46_1276 ();
 sg13g2_fill_1 FILLER_46_1288 ();
 sg13g2_fill_2 FILLER_46_1301 ();
 sg13g2_fill_1 FILLER_46_1303 ();
 sg13g2_decap_4 FILLER_46_1343 ();
 sg13g2_fill_2 FILLER_46_1347 ();
 sg13g2_fill_1 FILLER_46_1365 ();
 sg13g2_decap_8 FILLER_46_1401 ();
 sg13g2_decap_8 FILLER_46_1408 ();
 sg13g2_fill_2 FILLER_46_1415 ();
 sg13g2_fill_1 FILLER_46_1417 ();
 sg13g2_fill_1 FILLER_46_1433 ();
 sg13g2_decap_4 FILLER_46_1445 ();
 sg13g2_fill_1 FILLER_46_1449 ();
 sg13g2_decap_8 FILLER_46_1455 ();
 sg13g2_decap_8 FILLER_46_1462 ();
 sg13g2_fill_2 FILLER_46_1469 ();
 sg13g2_fill_1 FILLER_46_1471 ();
 sg13g2_fill_2 FILLER_46_1486 ();
 sg13g2_decap_8 FILLER_46_1496 ();
 sg13g2_decap_8 FILLER_46_1503 ();
 sg13g2_decap_8 FILLER_46_1510 ();
 sg13g2_decap_4 FILLER_46_1522 ();
 sg13g2_fill_2 FILLER_46_1526 ();
 sg13g2_fill_2 FILLER_46_1534 ();
 sg13g2_fill_1 FILLER_46_1544 ();
 sg13g2_fill_1 FILLER_46_1561 ();
 sg13g2_fill_1 FILLER_46_1566 ();
 sg13g2_fill_1 FILLER_46_1577 ();
 sg13g2_fill_1 FILLER_46_1591 ();
 sg13g2_fill_2 FILLER_46_1596 ();
 sg13g2_fill_1 FILLER_46_1598 ();
 sg13g2_decap_8 FILLER_46_1609 ();
 sg13g2_decap_4 FILLER_46_1616 ();
 sg13g2_decap_8 FILLER_46_1632 ();
 sg13g2_decap_8 FILLER_46_1639 ();
 sg13g2_decap_8 FILLER_46_1646 ();
 sg13g2_fill_2 FILLER_46_1687 ();
 sg13g2_fill_1 FILLER_46_1689 ();
 sg13g2_fill_2 FILLER_46_1695 ();
 sg13g2_decap_4 FILLER_46_1701 ();
 sg13g2_fill_2 FILLER_46_1713 ();
 sg13g2_fill_1 FILLER_46_1736 ();
 sg13g2_fill_1 FILLER_46_1741 ();
 sg13g2_fill_1 FILLER_46_1757 ();
 sg13g2_fill_1 FILLER_46_1763 ();
 sg13g2_decap_4 FILLER_46_1768 ();
 sg13g2_fill_2 FILLER_46_1772 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_11 ();
 sg13g2_fill_2 FILLER_47_18 ();
 sg13g2_fill_1 FILLER_47_20 ();
 sg13g2_decap_4 FILLER_47_26 ();
 sg13g2_fill_2 FILLER_47_30 ();
 sg13g2_fill_2 FILLER_47_37 ();
 sg13g2_decap_4 FILLER_47_44 ();
 sg13g2_fill_1 FILLER_47_48 ();
 sg13g2_fill_2 FILLER_47_54 ();
 sg13g2_decap_4 FILLER_47_65 ();
 sg13g2_fill_1 FILLER_47_69 ();
 sg13g2_decap_4 FILLER_47_75 ();
 sg13g2_decap_8 FILLER_47_92 ();
 sg13g2_decap_4 FILLER_47_99 ();
 sg13g2_fill_2 FILLER_47_103 ();
 sg13g2_fill_2 FILLER_47_108 ();
 sg13g2_fill_1 FILLER_47_110 ();
 sg13g2_fill_2 FILLER_47_117 ();
 sg13g2_decap_4 FILLER_47_127 ();
 sg13g2_fill_2 FILLER_47_131 ();
 sg13g2_decap_4 FILLER_47_142 ();
 sg13g2_fill_1 FILLER_47_146 ();
 sg13g2_decap_8 FILLER_47_155 ();
 sg13g2_fill_1 FILLER_47_162 ();
 sg13g2_decap_8 FILLER_47_176 ();
 sg13g2_fill_1 FILLER_47_183 ();
 sg13g2_fill_1 FILLER_47_193 ();
 sg13g2_fill_2 FILLER_47_204 ();
 sg13g2_fill_1 FILLER_47_210 ();
 sg13g2_fill_2 FILLER_47_226 ();
 sg13g2_fill_1 FILLER_47_228 ();
 sg13g2_fill_2 FILLER_47_233 ();
 sg13g2_fill_1 FILLER_47_235 ();
 sg13g2_fill_2 FILLER_47_247 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_decap_4 FILLER_47_258 ();
 sg13g2_fill_2 FILLER_47_262 ();
 sg13g2_fill_2 FILLER_47_274 ();
 sg13g2_decap_4 FILLER_47_280 ();
 sg13g2_fill_1 FILLER_47_289 ();
 sg13g2_decap_4 FILLER_47_299 ();
 sg13g2_fill_1 FILLER_47_303 ();
 sg13g2_fill_1 FILLER_47_308 ();
 sg13g2_fill_2 FILLER_47_377 ();
 sg13g2_fill_2 FILLER_47_389 ();
 sg13g2_fill_1 FILLER_47_421 ();
 sg13g2_fill_2 FILLER_47_443 ();
 sg13g2_fill_1 FILLER_47_445 ();
 sg13g2_fill_1 FILLER_47_480 ();
 sg13g2_decap_8 FILLER_47_486 ();
 sg13g2_decap_8 FILLER_47_493 ();
 sg13g2_decap_8 FILLER_47_500 ();
 sg13g2_decap_8 FILLER_47_507 ();
 sg13g2_decap_4 FILLER_47_514 ();
 sg13g2_decap_8 FILLER_47_544 ();
 sg13g2_decap_4 FILLER_47_551 ();
 sg13g2_fill_2 FILLER_47_555 ();
 sg13g2_fill_1 FILLER_47_591 ();
 sg13g2_decap_4 FILLER_47_596 ();
 sg13g2_fill_1 FILLER_47_616 ();
 sg13g2_fill_2 FILLER_47_629 ();
 sg13g2_fill_1 FILLER_47_645 ();
 sg13g2_fill_1 FILLER_47_654 ();
 sg13g2_decap_4 FILLER_47_690 ();
 sg13g2_fill_1 FILLER_47_694 ();
 sg13g2_decap_8 FILLER_47_711 ();
 sg13g2_fill_2 FILLER_47_718 ();
 sg13g2_fill_1 FILLER_47_729 ();
 sg13g2_decap_4 FILLER_47_741 ();
 sg13g2_fill_1 FILLER_47_745 ();
 sg13g2_fill_2 FILLER_47_766 ();
 sg13g2_fill_2 FILLER_47_786 ();
 sg13g2_fill_1 FILLER_47_788 ();
 sg13g2_fill_2 FILLER_47_818 ();
 sg13g2_fill_1 FILLER_47_820 ();
 sg13g2_fill_2 FILLER_47_825 ();
 sg13g2_fill_1 FILLER_47_827 ();
 sg13g2_fill_1 FILLER_47_868 ();
 sg13g2_decap_4 FILLER_47_872 ();
 sg13g2_fill_2 FILLER_47_876 ();
 sg13g2_fill_2 FILLER_47_881 ();
 sg13g2_fill_1 FILLER_47_883 ();
 sg13g2_fill_1 FILLER_47_900 ();
 sg13g2_decap_8 FILLER_47_919 ();
 sg13g2_decap_8 FILLER_47_926 ();
 sg13g2_decap_8 FILLER_47_933 ();
 sg13g2_decap_8 FILLER_47_940 ();
 sg13g2_fill_2 FILLER_47_988 ();
 sg13g2_decap_4 FILLER_47_995 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_fill_2 FILLER_47_1022 ();
 sg13g2_fill_1 FILLER_47_1024 ();
 sg13g2_fill_2 FILLER_47_1029 ();
 sg13g2_fill_2 FILLER_47_1039 ();
 sg13g2_fill_1 FILLER_47_1055 ();
 sg13g2_fill_1 FILLER_47_1069 ();
 sg13g2_decap_4 FILLER_47_1087 ();
 sg13g2_decap_8 FILLER_47_1120 ();
 sg13g2_decap_8 FILLER_47_1127 ();
 sg13g2_decap_8 FILLER_47_1134 ();
 sg13g2_fill_2 FILLER_47_1141 ();
 sg13g2_fill_1 FILLER_47_1143 ();
 sg13g2_fill_2 FILLER_47_1162 ();
 sg13g2_fill_1 FILLER_47_1164 ();
 sg13g2_decap_4 FILLER_47_1173 ();
 sg13g2_fill_1 FILLER_47_1177 ();
 sg13g2_fill_2 FILLER_47_1183 ();
 sg13g2_fill_1 FILLER_47_1200 ();
 sg13g2_fill_1 FILLER_47_1209 ();
 sg13g2_fill_2 FILLER_47_1224 ();
 sg13g2_fill_2 FILLER_47_1235 ();
 sg13g2_fill_1 FILLER_47_1237 ();
 sg13g2_fill_2 FILLER_47_1251 ();
 sg13g2_fill_1 FILLER_47_1270 ();
 sg13g2_fill_1 FILLER_47_1301 ();
 sg13g2_decap_4 FILLER_47_1307 ();
 sg13g2_fill_1 FILLER_47_1330 ();
 sg13g2_fill_2 FILLER_47_1340 ();
 sg13g2_fill_1 FILLER_47_1342 ();
 sg13g2_decap_4 FILLER_47_1351 ();
 sg13g2_fill_1 FILLER_47_1355 ();
 sg13g2_fill_1 FILLER_47_1374 ();
 sg13g2_fill_2 FILLER_47_1385 ();
 sg13g2_fill_1 FILLER_47_1387 ();
 sg13g2_fill_1 FILLER_47_1414 ();
 sg13g2_fill_1 FILLER_47_1420 ();
 sg13g2_fill_2 FILLER_47_1425 ();
 sg13g2_fill_2 FILLER_47_1432 ();
 sg13g2_decap_8 FILLER_47_1455 ();
 sg13g2_decap_8 FILLER_47_1462 ();
 sg13g2_decap_4 FILLER_47_1469 ();
 sg13g2_decap_8 FILLER_47_1487 ();
 sg13g2_decap_8 FILLER_47_1494 ();
 sg13g2_decap_4 FILLER_47_1501 ();
 sg13g2_fill_2 FILLER_47_1505 ();
 sg13g2_decap_8 FILLER_47_1525 ();
 sg13g2_decap_4 FILLER_47_1532 ();
 sg13g2_fill_2 FILLER_47_1541 ();
 sg13g2_decap_8 FILLER_47_1571 ();
 sg13g2_fill_1 FILLER_47_1578 ();
 sg13g2_decap_4 FILLER_47_1605 ();
 sg13g2_decap_8 FILLER_47_1613 ();
 sg13g2_fill_1 FILLER_47_1620 ();
 sg13g2_decap_4 FILLER_47_1629 ();
 sg13g2_fill_2 FILLER_47_1633 ();
 sg13g2_decap_8 FILLER_47_1656 ();
 sg13g2_decap_8 FILLER_47_1663 ();
 sg13g2_fill_2 FILLER_47_1670 ();
 sg13g2_fill_2 FILLER_47_1680 ();
 sg13g2_fill_2 FILLER_47_1690 ();
 sg13g2_fill_2 FILLER_47_1697 ();
 sg13g2_fill_1 FILLER_47_1699 ();
 sg13g2_decap_4 FILLER_47_1710 ();
 sg13g2_fill_1 FILLER_47_1719 ();
 sg13g2_fill_2 FILLER_47_1729 ();
 sg13g2_decap_4 FILLER_47_1743 ();
 sg13g2_decap_8 FILLER_47_1757 ();
 sg13g2_decap_8 FILLER_47_1764 ();
 sg13g2_fill_2 FILLER_47_1771 ();
 sg13g2_fill_1 FILLER_47_1773 ();
 sg13g2_fill_2 FILLER_48_55 ();
 sg13g2_fill_2 FILLER_48_88 ();
 sg13g2_fill_2 FILLER_48_117 ();
 sg13g2_fill_2 FILLER_48_125 ();
 sg13g2_fill_2 FILLER_48_143 ();
 sg13g2_decap_4 FILLER_48_185 ();
 sg13g2_fill_1 FILLER_48_189 ();
 sg13g2_fill_2 FILLER_48_198 ();
 sg13g2_fill_1 FILLER_48_205 ();
 sg13g2_fill_2 FILLER_48_212 ();
 sg13g2_fill_1 FILLER_48_214 ();
 sg13g2_decap_8 FILLER_48_221 ();
 sg13g2_fill_2 FILLER_48_228 ();
 sg13g2_fill_1 FILLER_48_230 ();
 sg13g2_decap_4 FILLER_48_244 ();
 sg13g2_fill_1 FILLER_48_248 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_fill_2 FILLER_48_282 ();
 sg13g2_fill_1 FILLER_48_284 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_fill_2 FILLER_48_298 ();
 sg13g2_decap_4 FILLER_48_305 ();
 sg13g2_fill_1 FILLER_48_309 ();
 sg13g2_fill_2 FILLER_48_320 ();
 sg13g2_decap_4 FILLER_48_329 ();
 sg13g2_fill_1 FILLER_48_333 ();
 sg13g2_fill_1 FILLER_48_339 ();
 sg13g2_fill_1 FILLER_48_363 ();
 sg13g2_fill_1 FILLER_48_374 ();
 sg13g2_fill_1 FILLER_48_391 ();
 sg13g2_fill_1 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_405 ();
 sg13g2_fill_1 FILLER_48_407 ();
 sg13g2_fill_1 FILLER_48_416 ();
 sg13g2_decap_4 FILLER_48_431 ();
 sg13g2_fill_2 FILLER_48_435 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_4 FILLER_48_448 ();
 sg13g2_fill_1 FILLER_48_452 ();
 sg13g2_decap_8 FILLER_48_474 ();
 sg13g2_fill_1 FILLER_48_481 ();
 sg13g2_fill_2 FILLER_48_487 ();
 sg13g2_fill_1 FILLER_48_489 ();
 sg13g2_decap_8 FILLER_48_515 ();
 sg13g2_fill_2 FILLER_48_522 ();
 sg13g2_fill_1 FILLER_48_524 ();
 sg13g2_fill_2 FILLER_48_529 ();
 sg13g2_fill_1 FILLER_48_538 ();
 sg13g2_fill_2 FILLER_48_569 ();
 sg13g2_fill_1 FILLER_48_571 ();
 sg13g2_fill_1 FILLER_48_576 ();
 sg13g2_fill_2 FILLER_48_587 ();
 sg13g2_fill_1 FILLER_48_589 ();
 sg13g2_fill_1 FILLER_48_609 ();
 sg13g2_fill_2 FILLER_48_646 ();
 sg13g2_fill_1 FILLER_48_678 ();
 sg13g2_fill_2 FILLER_48_687 ();
 sg13g2_fill_2 FILLER_48_694 ();
 sg13g2_fill_1 FILLER_48_709 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_fill_1 FILLER_48_721 ();
 sg13g2_decap_4 FILLER_48_738 ();
 sg13g2_fill_2 FILLER_48_742 ();
 sg13g2_fill_1 FILLER_48_761 ();
 sg13g2_decap_8 FILLER_48_767 ();
 sg13g2_decap_8 FILLER_48_774 ();
 sg13g2_fill_2 FILLER_48_785 ();
 sg13g2_fill_1 FILLER_48_787 ();
 sg13g2_fill_1 FILLER_48_793 ();
 sg13g2_decap_8 FILLER_48_799 ();
 sg13g2_decap_8 FILLER_48_806 ();
 sg13g2_fill_1 FILLER_48_813 ();
 sg13g2_fill_2 FILLER_48_826 ();
 sg13g2_fill_1 FILLER_48_831 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_4 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_fill_1 FILLER_48_895 ();
 sg13g2_decap_8 FILLER_48_900 ();
 sg13g2_fill_1 FILLER_48_907 ();
 sg13g2_decap_8 FILLER_48_921 ();
 sg13g2_decap_4 FILLER_48_938 ();
 sg13g2_fill_2 FILLER_48_949 ();
 sg13g2_fill_1 FILLER_48_951 ();
 sg13g2_fill_1 FILLER_48_955 ();
 sg13g2_fill_2 FILLER_48_967 ();
 sg13g2_decap_4 FILLER_48_974 ();
 sg13g2_decap_8 FILLER_48_982 ();
 sg13g2_fill_2 FILLER_48_1012 ();
 sg13g2_fill_1 FILLER_48_1014 ();
 sg13g2_decap_4 FILLER_48_1020 ();
 sg13g2_fill_2 FILLER_48_1032 ();
 sg13g2_fill_1 FILLER_48_1058 ();
 sg13g2_decap_4 FILLER_48_1069 ();
 sg13g2_fill_2 FILLER_48_1080 ();
 sg13g2_fill_1 FILLER_48_1082 ();
 sg13g2_decap_4 FILLER_48_1089 ();
 sg13g2_decap_4 FILLER_48_1099 ();
 sg13g2_fill_2 FILLER_48_1103 ();
 sg13g2_decap_4 FILLER_48_1112 ();
 sg13g2_fill_2 FILLER_48_1132 ();
 sg13g2_decap_8 FILLER_48_1138 ();
 sg13g2_fill_2 FILLER_48_1145 ();
 sg13g2_fill_1 FILLER_48_1147 ();
 sg13g2_fill_1 FILLER_48_1152 ();
 sg13g2_decap_4 FILLER_48_1159 ();
 sg13g2_fill_2 FILLER_48_1167 ();
 sg13g2_fill_1 FILLER_48_1183 ();
 sg13g2_fill_2 FILLER_48_1188 ();
 sg13g2_fill_2 FILLER_48_1194 ();
 sg13g2_decap_8 FILLER_48_1217 ();
 sg13g2_decap_4 FILLER_48_1224 ();
 sg13g2_fill_2 FILLER_48_1228 ();
 sg13g2_fill_2 FILLER_48_1261 ();
 sg13g2_decap_8 FILLER_48_1276 ();
 sg13g2_decap_4 FILLER_48_1283 ();
 sg13g2_fill_2 FILLER_48_1287 ();
 sg13g2_fill_2 FILLER_48_1297 ();
 sg13g2_fill_1 FILLER_48_1307 ();
 sg13g2_fill_2 FILLER_48_1319 ();
 sg13g2_fill_1 FILLER_48_1329 ();
 sg13g2_fill_1 FILLER_48_1369 ();
 sg13g2_decap_8 FILLER_48_1380 ();
 sg13g2_decap_8 FILLER_48_1387 ();
 sg13g2_decap_8 FILLER_48_1394 ();
 sg13g2_decap_4 FILLER_48_1401 ();
 sg13g2_fill_2 FILLER_48_1405 ();
 sg13g2_decap_8 FILLER_48_1412 ();
 sg13g2_fill_2 FILLER_48_1419 ();
 sg13g2_fill_1 FILLER_48_1421 ();
 sg13g2_fill_1 FILLER_48_1452 ();
 sg13g2_decap_8 FILLER_48_1461 ();
 sg13g2_decap_4 FILLER_48_1468 ();
 sg13g2_decap_8 FILLER_48_1486 ();
 sg13g2_decap_4 FILLER_48_1493 ();
 sg13g2_decap_4 FILLER_48_1505 ();
 sg13g2_fill_2 FILLER_48_1523 ();
 sg13g2_decap_4 FILLER_48_1529 ();
 sg13g2_fill_2 FILLER_48_1541 ();
 sg13g2_fill_1 FILLER_48_1543 ();
 sg13g2_fill_1 FILLER_48_1556 ();
 sg13g2_fill_2 FILLER_48_1573 ();
 sg13g2_fill_2 FILLER_48_1583 ();
 sg13g2_decap_4 FILLER_48_1589 ();
 sg13g2_fill_1 FILLER_48_1593 ();
 sg13g2_decap_8 FILLER_48_1599 ();
 sg13g2_decap_4 FILLER_48_1606 ();
 sg13g2_fill_2 FILLER_48_1610 ();
 sg13g2_fill_1 FILLER_48_1625 ();
 sg13g2_decap_4 FILLER_48_1638 ();
 sg13g2_fill_1 FILLER_48_1642 ();
 sg13g2_decap_4 FILLER_48_1651 ();
 sg13g2_fill_1 FILLER_48_1655 ();
 sg13g2_decap_8 FILLER_48_1664 ();
 sg13g2_decap_4 FILLER_48_1671 ();
 sg13g2_decap_8 FILLER_48_1691 ();
 sg13g2_fill_1 FILLER_48_1698 ();
 sg13g2_fill_2 FILLER_48_1704 ();
 sg13g2_decap_8 FILLER_48_1733 ();
 sg13g2_fill_2 FILLER_48_1740 ();
 sg13g2_fill_1 FILLER_48_1742 ();
 sg13g2_decap_8 FILLER_48_1751 ();
 sg13g2_decap_8 FILLER_48_1758 ();
 sg13g2_decap_8 FILLER_48_1765 ();
 sg13g2_fill_2 FILLER_48_1772 ();
 sg13g2_decap_8 FILLER_49_3 ();
 sg13g2_decap_8 FILLER_49_10 ();
 sg13g2_decap_4 FILLER_49_17 ();
 sg13g2_decap_4 FILLER_49_71 ();
 sg13g2_fill_1 FILLER_49_79 ();
 sg13g2_fill_1 FILLER_49_87 ();
 sg13g2_fill_2 FILLER_49_118 ();
 sg13g2_fill_1 FILLER_49_134 ();
 sg13g2_fill_1 FILLER_49_169 ();
 sg13g2_decap_8 FILLER_49_197 ();
 sg13g2_decap_4 FILLER_49_204 ();
 sg13g2_fill_1 FILLER_49_208 ();
 sg13g2_decap_4 FILLER_49_224 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_fill_1 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_257 ();
 sg13g2_decap_8 FILLER_49_264 ();
 sg13g2_fill_1 FILLER_49_271 ();
 sg13g2_fill_1 FILLER_49_281 ();
 sg13g2_fill_2 FILLER_49_309 ();
 sg13g2_decap_8 FILLER_49_316 ();
 sg13g2_decap_8 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_330 ();
 sg13g2_fill_1 FILLER_49_332 ();
 sg13g2_fill_1 FILLER_49_342 ();
 sg13g2_decap_8 FILLER_49_349 ();
 sg13g2_decap_8 FILLER_49_356 ();
 sg13g2_decap_4 FILLER_49_363 ();
 sg13g2_fill_1 FILLER_49_367 ();
 sg13g2_fill_2 FILLER_49_380 ();
 sg13g2_fill_2 FILLER_49_390 ();
 sg13g2_decap_4 FILLER_49_431 ();
 sg13g2_decap_4 FILLER_49_440 ();
 sg13g2_fill_1 FILLER_49_453 ();
 sg13g2_decap_8 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_480 ();
 sg13g2_decap_4 FILLER_49_495 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_fill_1 FILLER_49_511 ();
 sg13g2_fill_2 FILLER_49_522 ();
 sg13g2_fill_2 FILLER_49_529 ();
 sg13g2_fill_1 FILLER_49_547 ();
 sg13g2_fill_1 FILLER_49_562 ();
 sg13g2_fill_2 FILLER_49_584 ();
 sg13g2_fill_1 FILLER_49_586 ();
 sg13g2_decap_4 FILLER_49_595 ();
 sg13g2_fill_1 FILLER_49_599 ();
 sg13g2_fill_1 FILLER_49_605 ();
 sg13g2_fill_1 FILLER_49_615 ();
 sg13g2_fill_1 FILLER_49_631 ();
 sg13g2_fill_2 FILLER_49_639 ();
 sg13g2_fill_1 FILLER_49_645 ();
 sg13g2_fill_2 FILLER_49_653 ();
 sg13g2_fill_1 FILLER_49_659 ();
 sg13g2_fill_1 FILLER_49_663 ();
 sg13g2_fill_1 FILLER_49_682 ();
 sg13g2_fill_1 FILLER_49_688 ();
 sg13g2_fill_1 FILLER_49_695 ();
 sg13g2_fill_1 FILLER_49_702 ();
 sg13g2_fill_1 FILLER_49_708 ();
 sg13g2_decap_8 FILLER_49_718 ();
 sg13g2_decap_8 FILLER_49_725 ();
 sg13g2_fill_1 FILLER_49_732 ();
 sg13g2_fill_2 FILLER_49_737 ();
 sg13g2_fill_2 FILLER_49_745 ();
 sg13g2_decap_4 FILLER_49_765 ();
 sg13g2_fill_1 FILLER_49_774 ();
 sg13g2_fill_1 FILLER_49_780 ();
 sg13g2_fill_2 FILLER_49_785 ();
 sg13g2_fill_1 FILLER_49_799 ();
 sg13g2_fill_2 FILLER_49_805 ();
 sg13g2_fill_1 FILLER_49_819 ();
 sg13g2_fill_2 FILLER_49_825 ();
 sg13g2_fill_2 FILLER_49_831 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_fill_1 FILLER_49_866 ();
 sg13g2_decap_4 FILLER_49_871 ();
 sg13g2_fill_1 FILLER_49_880 ();
 sg13g2_decap_4 FILLER_49_886 ();
 sg13g2_fill_2 FILLER_49_902 ();
 sg13g2_decap_4 FILLER_49_915 ();
 sg13g2_fill_1 FILLER_49_919 ();
 sg13g2_decap_8 FILLER_49_928 ();
 sg13g2_fill_2 FILLER_49_935 ();
 sg13g2_fill_1 FILLER_49_937 ();
 sg13g2_fill_2 FILLER_49_942 ();
 sg13g2_fill_2 FILLER_49_949 ();
 sg13g2_fill_1 FILLER_49_951 ();
 sg13g2_fill_2 FILLER_49_958 ();
 sg13g2_fill_2 FILLER_49_965 ();
 sg13g2_fill_2 FILLER_49_991 ();
 sg13g2_fill_2 FILLER_49_998 ();
 sg13g2_decap_4 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1017 ();
 sg13g2_fill_2 FILLER_49_1033 ();
 sg13g2_fill_2 FILLER_49_1064 ();
 sg13g2_fill_2 FILLER_49_1071 ();
 sg13g2_fill_2 FILLER_49_1079 ();
 sg13g2_fill_1 FILLER_49_1081 ();
 sg13g2_decap_8 FILLER_49_1086 ();
 sg13g2_decap_8 FILLER_49_1093 ();
 sg13g2_decap_4 FILLER_49_1100 ();
 sg13g2_fill_1 FILLER_49_1104 ();
 sg13g2_fill_2 FILLER_49_1150 ();
 sg13g2_fill_2 FILLER_49_1175 ();
 sg13g2_fill_1 FILLER_49_1177 ();
 sg13g2_decap_4 FILLER_49_1208 ();
 sg13g2_fill_1 FILLER_49_1212 ();
 sg13g2_fill_1 FILLER_49_1221 ();
 sg13g2_fill_1 FILLER_49_1230 ();
 sg13g2_fill_2 FILLER_49_1252 ();
 sg13g2_decap_4 FILLER_49_1278 ();
 sg13g2_fill_2 FILLER_49_1290 ();
 sg13g2_decap_8 FILLER_49_1317 ();
 sg13g2_fill_2 FILLER_49_1324 ();
 sg13g2_fill_1 FILLER_49_1326 ();
 sg13g2_fill_2 FILLER_49_1342 ();
 sg13g2_decap_8 FILLER_49_1349 ();
 sg13g2_fill_2 FILLER_49_1395 ();
 sg13g2_decap_4 FILLER_49_1402 ();
 sg13g2_fill_2 FILLER_49_1406 ();
 sg13g2_fill_2 FILLER_49_1412 ();
 sg13g2_decap_8 FILLER_49_1422 ();
 sg13g2_fill_2 FILLER_49_1434 ();
 sg13g2_decap_8 FILLER_49_1462 ();
 sg13g2_fill_2 FILLER_49_1469 ();
 sg13g2_decap_4 FILLER_49_1486 ();
 sg13g2_fill_1 FILLER_49_1519 ();
 sg13g2_fill_2 FILLER_49_1548 ();
 sg13g2_fill_1 FILLER_49_1550 ();
 sg13g2_decap_8 FILLER_49_1556 ();
 sg13g2_decap_8 FILLER_49_1563 ();
 sg13g2_fill_2 FILLER_49_1570 ();
 sg13g2_fill_1 FILLER_49_1572 ();
 sg13g2_decap_8 FILLER_49_1591 ();
 sg13g2_fill_2 FILLER_49_1598 ();
 sg13g2_decap_4 FILLER_49_1604 ();
 sg13g2_fill_1 FILLER_49_1608 ();
 sg13g2_fill_2 FILLER_49_1612 ();
 sg13g2_fill_2 FILLER_49_1629 ();
 sg13g2_fill_1 FILLER_49_1631 ();
 sg13g2_decap_8 FILLER_49_1635 ();
 sg13g2_decap_8 FILLER_49_1642 ();
 sg13g2_fill_2 FILLER_49_1649 ();
 sg13g2_fill_1 FILLER_49_1651 ();
 sg13g2_fill_1 FILLER_49_1665 ();
 sg13g2_fill_2 FILLER_49_1720 ();
 sg13g2_fill_2 FILLER_49_1744 ();
 sg13g2_decap_8 FILLER_49_1751 ();
 sg13g2_decap_8 FILLER_49_1758 ();
 sg13g2_decap_8 FILLER_49_1765 ();
 sg13g2_fill_2 FILLER_49_1772 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_31 ();
 sg13g2_fill_1 FILLER_50_33 ();
 sg13g2_fill_1 FILLER_50_38 ();
 sg13g2_fill_1 FILLER_50_47 ();
 sg13g2_fill_1 FILLER_50_66 ();
 sg13g2_fill_1 FILLER_50_81 ();
 sg13g2_fill_1 FILLER_50_95 ();
 sg13g2_fill_1 FILLER_50_143 ();
 sg13g2_fill_1 FILLER_50_169 ();
 sg13g2_fill_2 FILLER_50_188 ();
 sg13g2_fill_2 FILLER_50_214 ();
 sg13g2_fill_1 FILLER_50_232 ();
 sg13g2_fill_2 FILLER_50_237 ();
 sg13g2_fill_2 FILLER_50_247 ();
 sg13g2_fill_1 FILLER_50_254 ();
 sg13g2_decap_8 FILLER_50_265 ();
 sg13g2_decap_4 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_276 ();
 sg13g2_decap_8 FILLER_50_286 ();
 sg13g2_decap_8 FILLER_50_293 ();
 sg13g2_decap_4 FILLER_50_300 ();
 sg13g2_fill_2 FILLER_50_309 ();
 sg13g2_fill_2 FILLER_50_327 ();
 sg13g2_fill_1 FILLER_50_329 ();
 sg13g2_fill_2 FILLER_50_340 ();
 sg13g2_decap_4 FILLER_50_346 ();
 sg13g2_fill_2 FILLER_50_350 ();
 sg13g2_decap_8 FILLER_50_393 ();
 sg13g2_decap_8 FILLER_50_404 ();
 sg13g2_fill_2 FILLER_50_411 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_fill_1 FILLER_50_441 ();
 sg13g2_decap_8 FILLER_50_446 ();
 sg13g2_fill_2 FILLER_50_453 ();
 sg13g2_fill_1 FILLER_50_455 ();
 sg13g2_fill_1 FILLER_50_464 ();
 sg13g2_decap_8 FILLER_50_473 ();
 sg13g2_decap_4 FILLER_50_480 ();
 sg13g2_decap_4 FILLER_50_499 ();
 sg13g2_fill_2 FILLER_50_527 ();
 sg13g2_fill_2 FILLER_50_538 ();
 sg13g2_fill_1 FILLER_50_567 ();
 sg13g2_fill_2 FILLER_50_589 ();
 sg13g2_fill_1 FILLER_50_591 ();
 sg13g2_fill_2 FILLER_50_605 ();
 sg13g2_fill_1 FILLER_50_607 ();
 sg13g2_fill_1 FILLER_50_629 ();
 sg13g2_fill_2 FILLER_50_641 ();
 sg13g2_fill_1 FILLER_50_661 ();
 sg13g2_fill_1 FILLER_50_679 ();
 sg13g2_fill_2 FILLER_50_694 ();
 sg13g2_fill_1 FILLER_50_705 ();
 sg13g2_fill_2 FILLER_50_711 ();
 sg13g2_decap_8 FILLER_50_717 ();
 sg13g2_decap_8 FILLER_50_724 ();
 sg13g2_decap_8 FILLER_50_755 ();
 sg13g2_fill_1 FILLER_50_767 ();
 sg13g2_decap_8 FILLER_50_772 ();
 sg13g2_fill_2 FILLER_50_779 ();
 sg13g2_fill_1 FILLER_50_797 ();
 sg13g2_fill_1 FILLER_50_803 ();
 sg13g2_fill_1 FILLER_50_812 ();
 sg13g2_fill_1 FILLER_50_830 ();
 sg13g2_fill_1 FILLER_50_839 ();
 sg13g2_fill_1 FILLER_50_862 ();
 sg13g2_fill_1 FILLER_50_871 ();
 sg13g2_decap_4 FILLER_50_884 ();
 sg13g2_fill_2 FILLER_50_893 ();
 sg13g2_fill_1 FILLER_50_899 ();
 sg13g2_fill_2 FILLER_50_904 ();
 sg13g2_fill_2 FILLER_50_917 ();
 sg13g2_decap_8 FILLER_50_928 ();
 sg13g2_decap_8 FILLER_50_935 ();
 sg13g2_fill_1 FILLER_50_942 ();
 sg13g2_decap_8 FILLER_50_952 ();
 sg13g2_decap_8 FILLER_50_963 ();
 sg13g2_fill_2 FILLER_50_970 ();
 sg13g2_fill_1 FILLER_50_972 ();
 sg13g2_fill_2 FILLER_50_978 ();
 sg13g2_fill_1 FILLER_50_980 ();
 sg13g2_decap_4 FILLER_50_999 ();
 sg13g2_fill_2 FILLER_50_1003 ();
 sg13g2_decap_8 FILLER_50_1009 ();
 sg13g2_decap_8 FILLER_50_1016 ();
 sg13g2_decap_8 FILLER_50_1023 ();
 sg13g2_fill_2 FILLER_50_1030 ();
 sg13g2_fill_1 FILLER_50_1032 ();
 sg13g2_fill_1 FILLER_50_1048 ();
 sg13g2_decap_8 FILLER_50_1054 ();
 sg13g2_fill_2 FILLER_50_1061 ();
 sg13g2_decap_8 FILLER_50_1079 ();
 sg13g2_fill_2 FILLER_50_1086 ();
 sg13g2_fill_1 FILLER_50_1088 ();
 sg13g2_fill_2 FILLER_50_1094 ();
 sg13g2_decap_8 FILLER_50_1100 ();
 sg13g2_fill_1 FILLER_50_1117 ();
 sg13g2_fill_2 FILLER_50_1130 ();
 sg13g2_fill_2 FILLER_50_1175 ();
 sg13g2_decap_4 FILLER_50_1187 ();
 sg13g2_fill_1 FILLER_50_1191 ();
 sg13g2_fill_1 FILLER_50_1197 ();
 sg13g2_fill_2 FILLER_50_1202 ();
 sg13g2_decap_8 FILLER_50_1212 ();
 sg13g2_decap_4 FILLER_50_1234 ();
 sg13g2_fill_1 FILLER_50_1238 ();
 sg13g2_fill_1 FILLER_50_1265 ();
 sg13g2_fill_2 FILLER_50_1272 ();
 sg13g2_fill_2 FILLER_50_1282 ();
 sg13g2_fill_2 FILLER_50_1295 ();
 sg13g2_decap_4 FILLER_50_1327 ();
 sg13g2_fill_2 FILLER_50_1331 ();
 sg13g2_decap_8 FILLER_50_1355 ();
 sg13g2_decap_4 FILLER_50_1371 ();
 sg13g2_fill_2 FILLER_50_1388 ();
 sg13g2_decap_4 FILLER_50_1399 ();
 sg13g2_fill_2 FILLER_50_1409 ();
 sg13g2_fill_1 FILLER_50_1415 ();
 sg13g2_fill_2 FILLER_50_1427 ();
 sg13g2_fill_1 FILLER_50_1429 ();
 sg13g2_fill_2 FILLER_50_1434 ();
 sg13g2_decap_8 FILLER_50_1452 ();
 sg13g2_decap_8 FILLER_50_1459 ();
 sg13g2_decap_8 FILLER_50_1466 ();
 sg13g2_decap_4 FILLER_50_1473 ();
 sg13g2_fill_1 FILLER_50_1481 ();
 sg13g2_decap_8 FILLER_50_1487 ();
 sg13g2_fill_2 FILLER_50_1494 ();
 sg13g2_fill_1 FILLER_50_1496 ();
 sg13g2_fill_1 FILLER_50_1505 ();
 sg13g2_decap_8 FILLER_50_1515 ();
 sg13g2_fill_2 FILLER_50_1522 ();
 sg13g2_fill_2 FILLER_50_1537 ();
 sg13g2_fill_1 FILLER_50_1539 ();
 sg13g2_decap_8 FILLER_50_1564 ();
 sg13g2_fill_1 FILLER_50_1581 ();
 sg13g2_fill_1 FILLER_50_1591 ();
 sg13g2_fill_1 FILLER_50_1635 ();
 sg13g2_decap_4 FILLER_50_1645 ();
 sg13g2_decap_4 FILLER_50_1665 ();
 sg13g2_decap_8 FILLER_50_1676 ();
 sg13g2_fill_1 FILLER_50_1683 ();
 sg13g2_decap_4 FILLER_50_1698 ();
 sg13g2_fill_2 FILLER_50_1707 ();
 sg13g2_fill_2 FILLER_50_1714 ();
 sg13g2_fill_1 FILLER_50_1734 ();
 sg13g2_fill_2 FILLER_50_1752 ();
 sg13g2_fill_1 FILLER_50_1754 ();
 sg13g2_decap_8 FILLER_50_1760 ();
 sg13g2_decap_8 FILLER_50_1767 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_11 ();
 sg13g2_decap_8 FILLER_51_18 ();
 sg13g2_fill_1 FILLER_51_25 ();
 sg13g2_decap_8 FILLER_51_33 ();
 sg13g2_decap_4 FILLER_51_48 ();
 sg13g2_fill_1 FILLER_51_52 ();
 sg13g2_fill_1 FILLER_51_57 ();
 sg13g2_fill_1 FILLER_51_70 ();
 sg13g2_fill_2 FILLER_51_89 ();
 sg13g2_fill_1 FILLER_51_97 ();
 sg13g2_fill_2 FILLER_51_102 ();
 sg13g2_fill_1 FILLER_51_146 ();
 sg13g2_fill_2 FILLER_51_160 ();
 sg13g2_decap_8 FILLER_51_213 ();
 sg13g2_fill_2 FILLER_51_220 ();
 sg13g2_decap_8 FILLER_51_238 ();
 sg13g2_decap_4 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_261 ();
 sg13g2_decap_8 FILLER_51_268 ();
 sg13g2_decap_8 FILLER_51_275 ();
 sg13g2_decap_8 FILLER_51_282 ();
 sg13g2_decap_4 FILLER_51_296 ();
 sg13g2_fill_1 FILLER_51_300 ();
 sg13g2_fill_1 FILLER_51_306 ();
 sg13g2_decap_8 FILLER_51_311 ();
 sg13g2_decap_4 FILLER_51_318 ();
 sg13g2_fill_1 FILLER_51_322 ();
 sg13g2_decap_8 FILLER_51_345 ();
 sg13g2_decap_4 FILLER_51_352 ();
 sg13g2_fill_2 FILLER_51_385 ();
 sg13g2_fill_1 FILLER_51_387 ();
 sg13g2_fill_2 FILLER_51_396 ();
 sg13g2_fill_1 FILLER_51_398 ();
 sg13g2_fill_1 FILLER_51_418 ();
 sg13g2_fill_2 FILLER_51_436 ();
 sg13g2_decap_4 FILLER_51_460 ();
 sg13g2_decap_8 FILLER_51_471 ();
 sg13g2_decap_4 FILLER_51_478 ();
 sg13g2_fill_2 FILLER_51_482 ();
 sg13g2_fill_2 FILLER_51_492 ();
 sg13g2_fill_1 FILLER_51_494 ();
 sg13g2_decap_4 FILLER_51_499 ();
 sg13g2_decap_8 FILLER_51_535 ();
 sg13g2_fill_1 FILLER_51_547 ();
 sg13g2_decap_8 FILLER_51_572 ();
 sg13g2_fill_2 FILLER_51_579 ();
 sg13g2_decap_8 FILLER_51_598 ();
 sg13g2_fill_2 FILLER_51_605 ();
 sg13g2_fill_1 FILLER_51_607 ();
 sg13g2_fill_1 FILLER_51_625 ();
 sg13g2_fill_1 FILLER_51_632 ();
 sg13g2_fill_1 FILLER_51_638 ();
 sg13g2_fill_2 FILLER_51_652 ();
 sg13g2_fill_1 FILLER_51_676 ();
 sg13g2_fill_1 FILLER_51_685 ();
 sg13g2_fill_1 FILLER_51_698 ();
 sg13g2_decap_4 FILLER_51_714 ();
 sg13g2_fill_1 FILLER_51_718 ();
 sg13g2_decap_8 FILLER_51_723 ();
 sg13g2_decap_8 FILLER_51_730 ();
 sg13g2_decap_8 FILLER_51_737 ();
 sg13g2_decap_8 FILLER_51_744 ();
 sg13g2_decap_4 FILLER_51_751 ();
 sg13g2_decap_4 FILLER_51_780 ();
 sg13g2_fill_2 FILLER_51_784 ();
 sg13g2_fill_1 FILLER_51_794 ();
 sg13g2_fill_2 FILLER_51_801 ();
 sg13g2_decap_4 FILLER_51_808 ();
 sg13g2_fill_2 FILLER_51_812 ();
 sg13g2_fill_2 FILLER_51_820 ();
 sg13g2_fill_2 FILLER_51_825 ();
 sg13g2_fill_2 FILLER_51_841 ();
 sg13g2_fill_2 FILLER_51_847 ();
 sg13g2_decap_4 FILLER_51_862 ();
 sg13g2_fill_1 FILLER_51_871 ();
 sg13g2_decap_4 FILLER_51_889 ();
 sg13g2_fill_1 FILLER_51_898 ();
 sg13g2_fill_1 FILLER_51_905 ();
 sg13g2_fill_1 FILLER_51_911 ();
 sg13g2_fill_1 FILLER_51_923 ();
 sg13g2_decap_4 FILLER_51_929 ();
 sg13g2_fill_2 FILLER_51_933 ();
 sg13g2_decap_4 FILLER_51_939 ();
 sg13g2_fill_1 FILLER_51_943 ();
 sg13g2_fill_1 FILLER_51_984 ();
 sg13g2_fill_1 FILLER_51_989 ();
 sg13g2_decap_8 FILLER_51_1006 ();
 sg13g2_fill_2 FILLER_51_1013 ();
 sg13g2_fill_1 FILLER_51_1015 ();
 sg13g2_fill_1 FILLER_51_1032 ();
 sg13g2_fill_1 FILLER_51_1042 ();
 sg13g2_fill_2 FILLER_51_1048 ();
 sg13g2_fill_1 FILLER_51_1055 ();
 sg13g2_fill_2 FILLER_51_1062 ();
 sg13g2_fill_2 FILLER_51_1069 ();
 sg13g2_fill_2 FILLER_51_1075 ();
 sg13g2_fill_1 FILLER_51_1077 ();
 sg13g2_fill_1 FILLER_51_1086 ();
 sg13g2_fill_1 FILLER_51_1095 ();
 sg13g2_fill_2 FILLER_51_1100 ();
 sg13g2_fill_2 FILLER_51_1110 ();
 sg13g2_fill_1 FILLER_51_1112 ();
 sg13g2_fill_2 FILLER_51_1127 ();
 sg13g2_fill_2 FILLER_51_1134 ();
 sg13g2_fill_1 FILLER_51_1136 ();
 sg13g2_fill_2 FILLER_51_1162 ();
 sg13g2_fill_1 FILLER_51_1164 ();
 sg13g2_fill_1 FILLER_51_1170 ();
 sg13g2_fill_2 FILLER_51_1181 ();
 sg13g2_fill_2 FILLER_51_1187 ();
 sg13g2_fill_2 FILLER_51_1194 ();
 sg13g2_fill_1 FILLER_51_1196 ();
 sg13g2_decap_8 FILLER_51_1210 ();
 sg13g2_decap_8 FILLER_51_1217 ();
 sg13g2_decap_8 FILLER_51_1224 ();
 sg13g2_fill_2 FILLER_51_1231 ();
 sg13g2_fill_1 FILLER_51_1233 ();
 sg13g2_fill_1 FILLER_51_1257 ();
 sg13g2_fill_1 FILLER_51_1277 ();
 sg13g2_fill_2 FILLER_51_1305 ();
 sg13g2_fill_1 FILLER_51_1322 ();
 sg13g2_fill_1 FILLER_51_1326 ();
 sg13g2_decap_8 FILLER_51_1339 ();
 sg13g2_decap_4 FILLER_51_1346 ();
 sg13g2_fill_2 FILLER_51_1362 ();
 sg13g2_fill_1 FILLER_51_1364 ();
 sg13g2_decap_8 FILLER_51_1373 ();
 sg13g2_fill_1 FILLER_51_1380 ();
 sg13g2_fill_1 FILLER_51_1384 ();
 sg13g2_fill_2 FILLER_51_1390 ();
 sg13g2_fill_2 FILLER_51_1399 ();
 sg13g2_decap_8 FILLER_51_1415 ();
 sg13g2_decap_8 FILLER_51_1422 ();
 sg13g2_fill_2 FILLER_51_1429 ();
 sg13g2_decap_8 FILLER_51_1436 ();
 sg13g2_fill_1 FILLER_51_1443 ();
 sg13g2_decap_8 FILLER_51_1457 ();
 sg13g2_decap_8 FILLER_51_1464 ();
 sg13g2_fill_1 FILLER_51_1471 ();
 sg13g2_fill_2 FILLER_51_1514 ();
 sg13g2_fill_1 FILLER_51_1529 ();
 sg13g2_fill_2 FILLER_51_1535 ();
 sg13g2_fill_2 FILLER_51_1545 ();
 sg13g2_decap_4 FILLER_51_1560 ();
 sg13g2_fill_1 FILLER_51_1564 ();
 sg13g2_fill_2 FILLER_51_1575 ();
 sg13g2_fill_1 FILLER_51_1599 ();
 sg13g2_fill_1 FILLER_51_1617 ();
 sg13g2_fill_2 FILLER_51_1652 ();
 sg13g2_decap_8 FILLER_51_1664 ();
 sg13g2_decap_4 FILLER_51_1671 ();
 sg13g2_fill_2 FILLER_51_1675 ();
 sg13g2_fill_2 FILLER_51_1681 ();
 sg13g2_fill_1 FILLER_51_1683 ();
 sg13g2_fill_1 FILLER_51_1695 ();
 sg13g2_decap_4 FILLER_51_1701 ();
 sg13g2_fill_2 FILLER_51_1709 ();
 sg13g2_fill_1 FILLER_51_1711 ();
 sg13g2_decap_4 FILLER_51_1721 ();
 sg13g2_fill_2 FILLER_51_1725 ();
 sg13g2_decap_4 FILLER_51_1732 ();
 sg13g2_fill_1 FILLER_51_1746 ();
 sg13g2_decap_8 FILLER_51_1767 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_14 ();
 sg13g2_fill_1 FILLER_52_32 ();
 sg13g2_decap_4 FILLER_52_37 ();
 sg13g2_fill_2 FILLER_52_46 ();
 sg13g2_fill_1 FILLER_52_48 ();
 sg13g2_fill_1 FILLER_52_54 ();
 sg13g2_fill_2 FILLER_52_69 ();
 sg13g2_fill_1 FILLER_52_71 ();
 sg13g2_fill_1 FILLER_52_89 ();
 sg13g2_fill_1 FILLER_52_145 ();
 sg13g2_fill_1 FILLER_52_154 ();
 sg13g2_fill_1 FILLER_52_169 ();
 sg13g2_fill_2 FILLER_52_173 ();
 sg13g2_decap_8 FILLER_52_191 ();
 sg13g2_decap_8 FILLER_52_198 ();
 sg13g2_decap_8 FILLER_52_205 ();
 sg13g2_decap_8 FILLER_52_212 ();
 sg13g2_decap_4 FILLER_52_219 ();
 sg13g2_decap_4 FILLER_52_239 ();
 sg13g2_fill_1 FILLER_52_243 ();
 sg13g2_fill_1 FILLER_52_252 ();
 sg13g2_fill_2 FILLER_52_257 ();
 sg13g2_fill_1 FILLER_52_277 ();
 sg13g2_fill_2 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_296 ();
 sg13g2_decap_8 FILLER_52_309 ();
 sg13g2_fill_2 FILLER_52_316 ();
 sg13g2_fill_1 FILLER_52_343 ();
 sg13g2_decap_8 FILLER_52_352 ();
 sg13g2_decap_8 FILLER_52_359 ();
 sg13g2_decap_8 FILLER_52_366 ();
 sg13g2_fill_2 FILLER_52_373 ();
 sg13g2_fill_1 FILLER_52_375 ();
 sg13g2_fill_1 FILLER_52_392 ();
 sg13g2_fill_1 FILLER_52_396 ();
 sg13g2_fill_2 FILLER_52_444 ();
 sg13g2_fill_2 FILLER_52_473 ();
 sg13g2_fill_1 FILLER_52_475 ();
 sg13g2_decap_8 FILLER_52_481 ();
 sg13g2_fill_1 FILLER_52_488 ();
 sg13g2_fill_2 FILLER_52_504 ();
 sg13g2_fill_1 FILLER_52_506 ();
 sg13g2_decap_8 FILLER_52_525 ();
 sg13g2_fill_2 FILLER_52_532 ();
 sg13g2_fill_2 FILLER_52_550 ();
 sg13g2_fill_1 FILLER_52_552 ();
 sg13g2_decap_4 FILLER_52_568 ();
 sg13g2_fill_1 FILLER_52_572 ();
 sg13g2_decap_4 FILLER_52_577 ();
 sg13g2_fill_2 FILLER_52_589 ();
 sg13g2_fill_1 FILLER_52_591 ();
 sg13g2_decap_8 FILLER_52_605 ();
 sg13g2_decap_8 FILLER_52_612 ();
 sg13g2_fill_2 FILLER_52_619 ();
 sg13g2_fill_1 FILLER_52_621 ();
 sg13g2_fill_2 FILLER_52_627 ();
 sg13g2_fill_1 FILLER_52_629 ();
 sg13g2_fill_1 FILLER_52_639 ();
 sg13g2_fill_2 FILLER_52_651 ();
 sg13g2_fill_2 FILLER_52_658 ();
 sg13g2_fill_1 FILLER_52_669 ();
 sg13g2_fill_1 FILLER_52_680 ();
 sg13g2_decap_4 FILLER_52_693 ();
 sg13g2_fill_1 FILLER_52_697 ();
 sg13g2_decap_8 FILLER_52_722 ();
 sg13g2_fill_2 FILLER_52_729 ();
 sg13g2_decap_4 FILLER_52_744 ();
 sg13g2_fill_2 FILLER_52_763 ();
 sg13g2_fill_1 FILLER_52_765 ();
 sg13g2_fill_1 FILLER_52_771 ();
 sg13g2_decap_8 FILLER_52_803 ();
 sg13g2_decap_4 FILLER_52_810 ();
 sg13g2_fill_2 FILLER_52_814 ();
 sg13g2_fill_1 FILLER_52_832 ();
 sg13g2_fill_2 FILLER_52_847 ();
 sg13g2_fill_1 FILLER_52_858 ();
 sg13g2_fill_2 FILLER_52_863 ();
 sg13g2_decap_4 FILLER_52_873 ();
 sg13g2_fill_1 FILLER_52_904 ();
 sg13g2_decap_8 FILLER_52_909 ();
 sg13g2_decap_8 FILLER_52_916 ();
 sg13g2_decap_8 FILLER_52_923 ();
 sg13g2_decap_8 FILLER_52_930 ();
 sg13g2_fill_1 FILLER_52_937 ();
 sg13g2_fill_2 FILLER_52_967 ();
 sg13g2_fill_1 FILLER_52_969 ();
 sg13g2_decap_8 FILLER_52_975 ();
 sg13g2_decap_8 FILLER_52_982 ();
 sg13g2_fill_1 FILLER_52_989 ();
 sg13g2_decap_4 FILLER_52_994 ();
 sg13g2_decap_8 FILLER_52_1012 ();
 sg13g2_fill_2 FILLER_52_1019 ();
 sg13g2_decap_4 FILLER_52_1031 ();
 sg13g2_fill_1 FILLER_52_1035 ();
 sg13g2_fill_2 FILLER_52_1050 ();
 sg13g2_decap_4 FILLER_52_1059 ();
 sg13g2_decap_4 FILLER_52_1071 ();
 sg13g2_decap_4 FILLER_52_1083 ();
 sg13g2_decap_8 FILLER_52_1115 ();
 sg13g2_fill_2 FILLER_52_1122 ();
 sg13g2_decap_8 FILLER_52_1127 ();
 sg13g2_decap_8 FILLER_52_1134 ();
 sg13g2_decap_8 FILLER_52_1141 ();
 sg13g2_decap_4 FILLER_52_1148 ();
 sg13g2_fill_1 FILLER_52_1152 ();
 sg13g2_decap_4 FILLER_52_1161 ();
 sg13g2_fill_1 FILLER_52_1174 ();
 sg13g2_fill_1 FILLER_52_1180 ();
 sg13g2_fill_1 FILLER_52_1185 ();
 sg13g2_fill_1 FILLER_52_1196 ();
 sg13g2_fill_1 FILLER_52_1201 ();
 sg13g2_decap_4 FILLER_52_1210 ();
 sg13g2_fill_2 FILLER_52_1214 ();
 sg13g2_decap_8 FILLER_52_1224 ();
 sg13g2_fill_2 FILLER_52_1231 ();
 sg13g2_fill_1 FILLER_52_1263 ();
 sg13g2_fill_1 FILLER_52_1273 ();
 sg13g2_fill_1 FILLER_52_1304 ();
 sg13g2_fill_2 FILLER_52_1342 ();
 sg13g2_decap_8 FILLER_52_1352 ();
 sg13g2_decap_4 FILLER_52_1359 ();
 sg13g2_fill_1 FILLER_52_1363 ();
 sg13g2_fill_1 FILLER_52_1386 ();
 sg13g2_decap_8 FILLER_52_1392 ();
 sg13g2_decap_8 FILLER_52_1399 ();
 sg13g2_fill_2 FILLER_52_1417 ();
 sg13g2_fill_1 FILLER_52_1419 ();
 sg13g2_fill_2 FILLER_52_1425 ();
 sg13g2_fill_2 FILLER_52_1439 ();
 sg13g2_decap_8 FILLER_52_1458 ();
 sg13g2_decap_4 FILLER_52_1465 ();
 sg13g2_fill_1 FILLER_52_1469 ();
 sg13g2_fill_1 FILLER_52_1493 ();
 sg13g2_fill_1 FILLER_52_1504 ();
 sg13g2_fill_1 FILLER_52_1510 ();
 sg13g2_fill_2 FILLER_52_1530 ();
 sg13g2_fill_1 FILLER_52_1578 ();
 sg13g2_fill_1 FILLER_52_1586 ();
 sg13g2_fill_1 FILLER_52_1612 ();
 sg13g2_fill_1 FILLER_52_1627 ();
 sg13g2_fill_2 FILLER_52_1642 ();
 sg13g2_fill_1 FILLER_52_1644 ();
 sg13g2_fill_1 FILLER_52_1648 ();
 sg13g2_decap_4 FILLER_52_1654 ();
 sg13g2_fill_1 FILLER_52_1658 ();
 sg13g2_fill_1 FILLER_52_1673 ();
 sg13g2_fill_2 FILLER_52_1684 ();
 sg13g2_fill_1 FILLER_52_1686 ();
 sg13g2_fill_1 FILLER_52_1691 ();
 sg13g2_fill_2 FILLER_52_1716 ();
 sg13g2_fill_1 FILLER_52_1718 ();
 sg13g2_decap_8 FILLER_52_1725 ();
 sg13g2_fill_2 FILLER_52_1732 ();
 sg13g2_fill_1 FILLER_52_1734 ();
 sg13g2_fill_2 FILLER_52_1740 ();
 sg13g2_decap_4 FILLER_52_1762 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_18 ();
 sg13g2_fill_1 FILLER_53_30 ();
 sg13g2_fill_2 FILLER_53_36 ();
 sg13g2_fill_1 FILLER_53_46 ();
 sg13g2_fill_2 FILLER_53_55 ();
 sg13g2_decap_4 FILLER_53_80 ();
 sg13g2_fill_1 FILLER_53_93 ();
 sg13g2_fill_1 FILLER_53_158 ();
 sg13g2_fill_1 FILLER_53_169 ();
 sg13g2_fill_2 FILLER_53_176 ();
 sg13g2_decap_8 FILLER_53_197 ();
 sg13g2_decap_8 FILLER_53_204 ();
 sg13g2_decap_8 FILLER_53_211 ();
 sg13g2_decap_8 FILLER_53_218 ();
 sg13g2_decap_8 FILLER_53_225 ();
 sg13g2_decap_8 FILLER_53_232 ();
 sg13g2_fill_1 FILLER_53_243 ();
 sg13g2_decap_4 FILLER_53_277 ();
 sg13g2_decap_8 FILLER_53_290 ();
 sg13g2_decap_8 FILLER_53_297 ();
 sg13g2_decap_8 FILLER_53_304 ();
 sg13g2_fill_2 FILLER_53_311 ();
 sg13g2_fill_1 FILLER_53_313 ();
 sg13g2_fill_2 FILLER_53_328 ();
 sg13g2_fill_1 FILLER_53_330 ();
 sg13g2_fill_2 FILLER_53_350 ();
 sg13g2_fill_2 FILLER_53_369 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_fill_2 FILLER_53_438 ();
 sg13g2_fill_1 FILLER_53_440 ();
 sg13g2_fill_1 FILLER_53_451 ();
 sg13g2_decap_4 FILLER_53_456 ();
 sg13g2_fill_2 FILLER_53_474 ();
 sg13g2_decap_4 FILLER_53_481 ();
 sg13g2_fill_1 FILLER_53_485 ();
 sg13g2_decap_4 FILLER_53_527 ();
 sg13g2_fill_1 FILLER_53_531 ();
 sg13g2_decap_8 FILLER_53_537 ();
 sg13g2_decap_8 FILLER_53_544 ();
 sg13g2_decap_8 FILLER_53_551 ();
 sg13g2_fill_2 FILLER_53_558 ();
 sg13g2_fill_2 FILLER_53_578 ();
 sg13g2_fill_2 FILLER_53_592 ();
 sg13g2_fill_1 FILLER_53_607 ();
 sg13g2_fill_2 FILLER_53_616 ();
 sg13g2_fill_1 FILLER_53_618 ();
 sg13g2_decap_8 FILLER_53_623 ();
 sg13g2_decap_8 FILLER_53_630 ();
 sg13g2_fill_1 FILLER_53_637 ();
 sg13g2_fill_2 FILLER_53_644 ();
 sg13g2_fill_1 FILLER_53_651 ();
 sg13g2_fill_2 FILLER_53_674 ();
 sg13g2_fill_1 FILLER_53_676 ();
 sg13g2_fill_2 FILLER_53_683 ();
 sg13g2_decap_8 FILLER_53_690 ();
 sg13g2_decap_4 FILLER_53_697 ();
 sg13g2_decap_4 FILLER_53_708 ();
 sg13g2_decap_4 FILLER_53_721 ();
 sg13g2_fill_1 FILLER_53_725 ();
 sg13g2_fill_1 FILLER_53_731 ();
 sg13g2_decap_4 FILLER_53_740 ();
 sg13g2_fill_2 FILLER_53_757 ();
 sg13g2_decap_4 FILLER_53_764 ();
 sg13g2_fill_2 FILLER_53_768 ();
 sg13g2_decap_8 FILLER_53_800 ();
 sg13g2_decap_8 FILLER_53_807 ();
 sg13g2_decap_8 FILLER_53_814 ();
 sg13g2_fill_2 FILLER_53_821 ();
 sg13g2_fill_1 FILLER_53_823 ();
 sg13g2_fill_2 FILLER_53_833 ();
 sg13g2_fill_1 FILLER_53_835 ();
 sg13g2_fill_2 FILLER_53_862 ();
 sg13g2_fill_1 FILLER_53_864 ();
 sg13g2_fill_1 FILLER_53_884 ();
 sg13g2_decap_4 FILLER_53_889 ();
 sg13g2_fill_2 FILLER_53_903 ();
 sg13g2_decap_4 FILLER_53_931 ();
 sg13g2_decap_8 FILLER_53_938 ();
 sg13g2_decap_8 FILLER_53_945 ();
 sg13g2_fill_1 FILLER_53_952 ();
 sg13g2_fill_1 FILLER_53_965 ();
 sg13g2_decap_8 FILLER_53_976 ();
 sg13g2_decap_4 FILLER_53_983 ();
 sg13g2_fill_2 FILLER_53_987 ();
 sg13g2_fill_1 FILLER_53_1002 ();
 sg13g2_fill_2 FILLER_53_1036 ();
 sg13g2_fill_1 FILLER_53_1038 ();
 sg13g2_fill_2 FILLER_53_1049 ();
 sg13g2_decap_8 FILLER_53_1082 ();
 sg13g2_fill_2 FILLER_53_1097 ();
 sg13g2_fill_1 FILLER_53_1099 ();
 sg13g2_fill_1 FILLER_53_1104 ();
 sg13g2_fill_1 FILLER_53_1110 ();
 sg13g2_decap_4 FILLER_53_1116 ();
 sg13g2_fill_1 FILLER_53_1120 ();
 sg13g2_decap_4 FILLER_53_1151 ();
 sg13g2_fill_1 FILLER_53_1155 ();
 sg13g2_decap_8 FILLER_53_1160 ();
 sg13g2_fill_2 FILLER_53_1188 ();
 sg13g2_fill_1 FILLER_53_1190 ();
 sg13g2_decap_8 FILLER_53_1199 ();
 sg13g2_fill_2 FILLER_53_1206 ();
 sg13g2_decap_8 FILLER_53_1221 ();
 sg13g2_fill_2 FILLER_53_1228 ();
 sg13g2_fill_2 FILLER_53_1253 ();
 sg13g2_fill_1 FILLER_53_1255 ();
 sg13g2_fill_1 FILLER_53_1306 ();
 sg13g2_decap_4 FILLER_53_1312 ();
 sg13g2_fill_1 FILLER_53_1316 ();
 sg13g2_fill_2 FILLER_53_1346 ();
 sg13g2_fill_1 FILLER_53_1353 ();
 sg13g2_fill_2 FILLER_53_1394 ();
 sg13g2_decap_4 FILLER_53_1426 ();
 sg13g2_fill_1 FILLER_53_1430 ();
 sg13g2_fill_1 FILLER_53_1439 ();
 sg13g2_fill_2 FILLER_53_1463 ();
 sg13g2_fill_1 FILLER_53_1465 ();
 sg13g2_decap_8 FILLER_53_1473 ();
 sg13g2_decap_8 FILLER_53_1480 ();
 sg13g2_fill_2 FILLER_53_1487 ();
 sg13g2_fill_1 FILLER_53_1489 ();
 sg13g2_decap_8 FILLER_53_1515 ();
 sg13g2_fill_1 FILLER_53_1522 ();
 sg13g2_fill_2 FILLER_53_1531 ();
 sg13g2_fill_1 FILLER_53_1533 ();
 sg13g2_decap_8 FILLER_53_1539 ();
 sg13g2_fill_2 FILLER_53_1546 ();
 sg13g2_fill_1 FILLER_53_1548 ();
 sg13g2_fill_2 FILLER_53_1562 ();
 sg13g2_fill_1 FILLER_53_1612 ();
 sg13g2_fill_1 FILLER_53_1621 ();
 sg13g2_fill_2 FILLER_53_1643 ();
 sg13g2_fill_1 FILLER_53_1664 ();
 sg13g2_decap_8 FILLER_53_1681 ();
 sg13g2_decap_4 FILLER_53_1694 ();
 sg13g2_fill_1 FILLER_53_1698 ();
 sg13g2_fill_2 FILLER_53_1716 ();
 sg13g2_fill_2 FILLER_53_1723 ();
 sg13g2_fill_1 FILLER_53_1725 ();
 sg13g2_fill_2 FILLER_53_1732 ();
 sg13g2_fill_1 FILLER_53_1734 ();
 sg13g2_fill_2 FILLER_53_1740 ();
 sg13g2_fill_1 FILLER_53_1750 ();
 sg13g2_decap_4 FILLER_53_1760 ();
 sg13g2_decap_4 FILLER_53_1769 ();
 sg13g2_fill_1 FILLER_53_1773 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_4 FILLER_54_14 ();
 sg13g2_fill_2 FILLER_54_18 ();
 sg13g2_fill_1 FILLER_54_36 ();
 sg13g2_fill_1 FILLER_54_42 ();
 sg13g2_fill_2 FILLER_54_136 ();
 sg13g2_fill_1 FILLER_54_138 ();
 sg13g2_decap_8 FILLER_54_144 ();
 sg13g2_decap_8 FILLER_54_151 ();
 sg13g2_fill_1 FILLER_54_158 ();
 sg13g2_fill_1 FILLER_54_206 ();
 sg13g2_decap_4 FILLER_54_220 ();
 sg13g2_decap_8 FILLER_54_228 ();
 sg13g2_fill_2 FILLER_54_235 ();
 sg13g2_fill_2 FILLER_54_245 ();
 sg13g2_fill_1 FILLER_54_252 ();
 sg13g2_decap_8 FILLER_54_257 ();
 sg13g2_fill_2 FILLER_54_264 ();
 sg13g2_decap_4 FILLER_54_279 ();
 sg13g2_fill_1 FILLER_54_297 ();
 sg13g2_fill_1 FILLER_54_303 ();
 sg13g2_fill_1 FILLER_54_309 ();
 sg13g2_fill_1 FILLER_54_315 ();
 sg13g2_fill_1 FILLER_54_325 ();
 sg13g2_fill_2 FILLER_54_350 ();
 sg13g2_fill_1 FILLER_54_352 ();
 sg13g2_fill_2 FILLER_54_374 ();
 sg13g2_fill_2 FILLER_54_383 ();
 sg13g2_fill_1 FILLER_54_393 ();
 sg13g2_fill_2 FILLER_54_405 ();
 sg13g2_fill_2 FILLER_54_415 ();
 sg13g2_fill_1 FILLER_54_433 ();
 sg13g2_decap_8 FILLER_54_478 ();
 sg13g2_decap_4 FILLER_54_493 ();
 sg13g2_decap_4 FILLER_54_505 ();
 sg13g2_fill_1 FILLER_54_509 ();
 sg13g2_fill_1 FILLER_54_541 ();
 sg13g2_decap_4 FILLER_54_545 ();
 sg13g2_decap_4 FILLER_54_553 ();
 sg13g2_fill_1 FILLER_54_585 ();
 sg13g2_decap_8 FILLER_54_599 ();
 sg13g2_fill_2 FILLER_54_606 ();
 sg13g2_decap_8 FILLER_54_617 ();
 sg13g2_decap_4 FILLER_54_624 ();
 sg13g2_fill_2 FILLER_54_628 ();
 sg13g2_fill_2 FILLER_54_644 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_1 FILLER_54_692 ();
 sg13g2_decap_8 FILLER_54_699 ();
 sg13g2_decap_4 FILLER_54_724 ();
 sg13g2_fill_1 FILLER_54_728 ();
 sg13g2_decap_8 FILLER_54_741 ();
 sg13g2_decap_4 FILLER_54_748 ();
 sg13g2_fill_2 FILLER_54_752 ();
 sg13g2_decap_4 FILLER_54_758 ();
 sg13g2_fill_2 FILLER_54_762 ();
 sg13g2_fill_1 FILLER_54_772 ();
 sg13g2_fill_2 FILLER_54_786 ();
 sg13g2_fill_1 FILLER_54_788 ();
 sg13g2_decap_8 FILLER_54_802 ();
 sg13g2_fill_2 FILLER_54_809 ();
 sg13g2_fill_1 FILLER_54_811 ();
 sg13g2_decap_4 FILLER_54_820 ();
 sg13g2_fill_1 FILLER_54_824 ();
 sg13g2_decap_8 FILLER_54_854 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_decap_8 FILLER_54_866 ();
 sg13g2_fill_1 FILLER_54_873 ();
 sg13g2_decap_8 FILLER_54_882 ();
 sg13g2_decap_4 FILLER_54_909 ();
 sg13g2_decap_4 FILLER_54_932 ();
 sg13g2_decap_4 FILLER_54_940 ();
 sg13g2_fill_1 FILLER_54_944 ();
 sg13g2_fill_1 FILLER_54_974 ();
 sg13g2_decap_4 FILLER_54_1030 ();
 sg13g2_fill_1 FILLER_54_1034 ();
 sg13g2_decap_8 FILLER_54_1043 ();
 sg13g2_fill_1 FILLER_54_1066 ();
 sg13g2_decap_4 FILLER_54_1076 ();
 sg13g2_decap_4 FILLER_54_1097 ();
 sg13g2_fill_2 FILLER_54_1101 ();
 sg13g2_decap_4 FILLER_54_1124 ();
 sg13g2_fill_2 FILLER_54_1132 ();
 sg13g2_fill_1 FILLER_54_1134 ();
 sg13g2_fill_1 FILLER_54_1138 ();
 sg13g2_fill_2 FILLER_54_1151 ();
 sg13g2_fill_1 FILLER_54_1153 ();
 sg13g2_fill_2 FILLER_54_1159 ();
 sg13g2_fill_1 FILLER_54_1161 ();
 sg13g2_decap_4 FILLER_54_1170 ();
 sg13g2_fill_2 FILLER_54_1174 ();
 sg13g2_decap_8 FILLER_54_1187 ();
 sg13g2_fill_1 FILLER_54_1194 ();
 sg13g2_fill_2 FILLER_54_1203 ();
 sg13g2_decap_8 FILLER_54_1230 ();
 sg13g2_decap_4 FILLER_54_1237 ();
 sg13g2_fill_2 FILLER_54_1241 ();
 sg13g2_decap_4 FILLER_54_1262 ();
 sg13g2_fill_1 FILLER_54_1266 ();
 sg13g2_fill_1 FILLER_54_1271 ();
 sg13g2_decap_8 FILLER_54_1284 ();
 sg13g2_fill_1 FILLER_54_1301 ();
 sg13g2_decap_4 FILLER_54_1306 ();
 sg13g2_fill_1 FILLER_54_1310 ();
 sg13g2_fill_2 FILLER_54_1334 ();
 sg13g2_fill_2 FILLER_54_1348 ();
 sg13g2_fill_2 FILLER_54_1371 ();
 sg13g2_fill_1 FILLER_54_1373 ();
 sg13g2_decap_8 FILLER_54_1380 ();
 sg13g2_decap_8 FILLER_54_1391 ();
 sg13g2_decap_4 FILLER_54_1398 ();
 sg13g2_fill_2 FILLER_54_1402 ();
 sg13g2_decap_4 FILLER_54_1419 ();
 sg13g2_decap_8 FILLER_54_1434 ();
 sg13g2_decap_8 FILLER_54_1441 ();
 sg13g2_decap_8 FILLER_54_1448 ();
 sg13g2_fill_1 FILLER_54_1455 ();
 sg13g2_fill_1 FILLER_54_1469 ();
 sg13g2_decap_4 FILLER_54_1480 ();
 sg13g2_fill_2 FILLER_54_1489 ();
 sg13g2_decap_4 FILLER_54_1510 ();
 sg13g2_decap_4 FILLER_54_1527 ();
 sg13g2_fill_2 FILLER_54_1531 ();
 sg13g2_decap_4 FILLER_54_1541 ();
 sg13g2_fill_1 FILLER_54_1545 ();
 sg13g2_fill_2 FILLER_54_1551 ();
 sg13g2_decap_4 FILLER_54_1571 ();
 sg13g2_fill_2 FILLER_54_1575 ();
 sg13g2_decap_8 FILLER_54_1584 ();
 sg13g2_fill_1 FILLER_54_1591 ();
 sg13g2_fill_2 FILLER_54_1597 ();
 sg13g2_fill_2 FILLER_54_1607 ();
 sg13g2_fill_1 FILLER_54_1628 ();
 sg13g2_fill_1 FILLER_54_1639 ();
 sg13g2_fill_2 FILLER_54_1643 ();
 sg13g2_fill_1 FILLER_54_1661 ();
 sg13g2_decap_8 FILLER_54_1687 ();
 sg13g2_decap_8 FILLER_54_1710 ();
 sg13g2_fill_2 FILLER_54_1717 ();
 sg13g2_fill_1 FILLER_54_1719 ();
 sg13g2_fill_1 FILLER_54_1730 ();
 sg13g2_fill_1 FILLER_54_1752 ();
 sg13g2_fill_1 FILLER_54_1758 ();
 sg13g2_decap_8 FILLER_54_1767 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_4 FILLER_55_14 ();
 sg13g2_fill_2 FILLER_55_18 ();
 sg13g2_fill_1 FILLER_55_30 ();
 sg13g2_fill_1 FILLER_55_64 ();
 sg13g2_fill_1 FILLER_55_122 ();
 sg13g2_fill_2 FILLER_55_139 ();
 sg13g2_fill_1 FILLER_55_141 ();
 sg13g2_fill_2 FILLER_55_160 ();
 sg13g2_decap_8 FILLER_55_167 ();
 sg13g2_decap_8 FILLER_55_174 ();
 sg13g2_decap_8 FILLER_55_181 ();
 sg13g2_fill_1 FILLER_55_188 ();
 sg13g2_fill_2 FILLER_55_197 ();
 sg13g2_decap_4 FILLER_55_205 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_fill_1 FILLER_55_233 ();
 sg13g2_fill_1 FILLER_55_242 ();
 sg13g2_decap_8 FILLER_55_256 ();
 sg13g2_decap_4 FILLER_55_263 ();
 sg13g2_fill_1 FILLER_55_267 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_4 FILLER_55_287 ();
 sg13g2_decap_4 FILLER_55_300 ();
 sg13g2_fill_2 FILLER_55_308 ();
 sg13g2_fill_1 FILLER_55_310 ();
 sg13g2_fill_2 FILLER_55_317 ();
 sg13g2_fill_1 FILLER_55_319 ();
 sg13g2_decap_4 FILLER_55_332 ();
 sg13g2_fill_2 FILLER_55_336 ();
 sg13g2_fill_1 FILLER_55_350 ();
 sg13g2_fill_1 FILLER_55_364 ();
 sg13g2_fill_1 FILLER_55_370 ();
 sg13g2_fill_1 FILLER_55_378 ();
 sg13g2_fill_2 FILLER_55_394 ();
 sg13g2_decap_8 FILLER_55_431 ();
 sg13g2_fill_1 FILLER_55_438 ();
 sg13g2_decap_4 FILLER_55_444 ();
 sg13g2_decap_8 FILLER_55_453 ();
 sg13g2_fill_2 FILLER_55_472 ();
 sg13g2_decap_4 FILLER_55_479 ();
 sg13g2_decap_8 FILLER_55_504 ();
 sg13g2_decap_4 FILLER_55_511 ();
 sg13g2_fill_1 FILLER_55_523 ();
 sg13g2_fill_2 FILLER_55_527 ();
 sg13g2_fill_1 FILLER_55_529 ();
 sg13g2_decap_8 FILLER_55_574 ();
 sg13g2_decap_4 FILLER_55_581 ();
 sg13g2_decap_8 FILLER_55_597 ();
 sg13g2_decap_8 FILLER_55_604 ();
 sg13g2_decap_8 FILLER_55_611 ();
 sg13g2_decap_8 FILLER_55_618 ();
 sg13g2_decap_4 FILLER_55_625 ();
 sg13g2_decap_4 FILLER_55_639 ();
 sg13g2_fill_1 FILLER_55_643 ();
 sg13g2_fill_2 FILLER_55_652 ();
 sg13g2_fill_1 FILLER_55_671 ();
 sg13g2_fill_1 FILLER_55_677 ();
 sg13g2_fill_1 FILLER_55_686 ();
 sg13g2_fill_1 FILLER_55_701 ();
 sg13g2_decap_8 FILLER_55_723 ();
 sg13g2_decap_8 FILLER_55_730 ();
 sg13g2_decap_8 FILLER_55_737 ();
 sg13g2_decap_8 FILLER_55_744 ();
 sg13g2_decap_4 FILLER_55_751 ();
 sg13g2_fill_1 FILLER_55_755 ();
 sg13g2_fill_2 FILLER_55_786 ();
 sg13g2_fill_1 FILLER_55_788 ();
 sg13g2_decap_4 FILLER_55_803 ();
 sg13g2_fill_1 FILLER_55_820 ();
 sg13g2_decap_4 FILLER_55_827 ();
 sg13g2_fill_2 FILLER_55_841 ();
 sg13g2_fill_1 FILLER_55_843 ();
 sg13g2_fill_2 FILLER_55_857 ();
 sg13g2_fill_2 FILLER_55_863 ();
 sg13g2_fill_2 FILLER_55_869 ();
 sg13g2_decap_4 FILLER_55_883 ();
 sg13g2_fill_2 FILLER_55_887 ();
 sg13g2_decap_8 FILLER_55_904 ();
 sg13g2_decap_4 FILLER_55_911 ();
 sg13g2_fill_1 FILLER_55_915 ();
 sg13g2_fill_2 FILLER_55_932 ();
 sg13g2_fill_1 FILLER_55_934 ();
 sg13g2_fill_2 FILLER_55_946 ();
 sg13g2_decap_4 FILLER_55_964 ();
 sg13g2_decap_8 FILLER_55_973 ();
 sg13g2_decap_4 FILLER_55_980 ();
 sg13g2_fill_2 FILLER_55_984 ();
 sg13g2_fill_1 FILLER_55_991 ();
 sg13g2_fill_1 FILLER_55_997 ();
 sg13g2_fill_2 FILLER_55_1027 ();
 sg13g2_fill_1 FILLER_55_1029 ();
 sg13g2_fill_1 FILLER_55_1054 ();
 sg13g2_fill_2 FILLER_55_1058 ();
 sg13g2_fill_1 FILLER_55_1060 ();
 sg13g2_fill_2 FILLER_55_1069 ();
 sg13g2_fill_1 FILLER_55_1110 ();
 sg13g2_fill_1 FILLER_55_1119 ();
 sg13g2_decap_8 FILLER_55_1124 ();
 sg13g2_decap_4 FILLER_55_1131 ();
 sg13g2_fill_1 FILLER_55_1135 ();
 sg13g2_fill_1 FILLER_55_1148 ();
 sg13g2_fill_2 FILLER_55_1154 ();
 sg13g2_fill_1 FILLER_55_1164 ();
 sg13g2_decap_4 FILLER_55_1184 ();
 sg13g2_fill_1 FILLER_55_1188 ();
 sg13g2_fill_2 FILLER_55_1202 ();
 sg13g2_fill_1 FILLER_55_1204 ();
 sg13g2_decap_4 FILLER_55_1213 ();
 sg13g2_decap_4 FILLER_55_1221 ();
 sg13g2_fill_2 FILLER_55_1225 ();
 sg13g2_fill_1 FILLER_55_1235 ();
 sg13g2_decap_4 FILLER_55_1278 ();
 sg13g2_fill_2 FILLER_55_1282 ();
 sg13g2_fill_1 FILLER_55_1310 ();
 sg13g2_fill_1 FILLER_55_1317 ();
 sg13g2_fill_1 FILLER_55_1329 ();
 sg13g2_fill_2 FILLER_55_1338 ();
 sg13g2_fill_2 FILLER_55_1358 ();
 sg13g2_fill_1 FILLER_55_1360 ();
 sg13g2_fill_2 FILLER_55_1384 ();
 sg13g2_fill_1 FILLER_55_1386 ();
 sg13g2_decap_8 FILLER_55_1429 ();
 sg13g2_decap_8 FILLER_55_1436 ();
 sg13g2_decap_8 FILLER_55_1443 ();
 sg13g2_fill_2 FILLER_55_1450 ();
 sg13g2_fill_1 FILLER_55_1452 ();
 sg13g2_fill_2 FILLER_55_1483 ();
 sg13g2_fill_1 FILLER_55_1485 ();
 sg13g2_fill_2 FILLER_55_1504 ();
 sg13g2_fill_2 FILLER_55_1532 ();
 sg13g2_fill_1 FILLER_55_1534 ();
 sg13g2_decap_8 FILLER_55_1539 ();
 sg13g2_fill_2 FILLER_55_1546 ();
 sg13g2_fill_1 FILLER_55_1548 ();
 sg13g2_fill_2 FILLER_55_1554 ();
 sg13g2_fill_1 FILLER_55_1556 ();
 sg13g2_decap_8 FILLER_55_1579 ();
 sg13g2_fill_2 FILLER_55_1586 ();
 sg13g2_decap_8 FILLER_55_1592 ();
 sg13g2_decap_8 FILLER_55_1608 ();
 sg13g2_fill_1 FILLER_55_1615 ();
 sg13g2_fill_2 FILLER_55_1634 ();
 sg13g2_fill_2 FILLER_55_1648 ();
 sg13g2_fill_1 FILLER_55_1670 ();
 sg13g2_fill_2 FILLER_55_1692 ();
 sg13g2_fill_1 FILLER_55_1747 ();
 sg13g2_decap_4 FILLER_55_1752 ();
 sg13g2_fill_2 FILLER_55_1761 ();
 sg13g2_decap_4 FILLER_55_1768 ();
 sg13g2_fill_2 FILLER_55_1772 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_16 ();
 sg13g2_fill_1 FILLER_56_28 ();
 sg13g2_fill_1 FILLER_56_45 ();
 sg13g2_fill_2 FILLER_56_51 ();
 sg13g2_fill_1 FILLER_56_72 ();
 sg13g2_fill_1 FILLER_56_89 ();
 sg13g2_fill_2 FILLER_56_94 ();
 sg13g2_fill_2 FILLER_56_125 ();
 sg13g2_fill_1 FILLER_56_131 ();
 sg13g2_fill_2 FILLER_56_151 ();
 sg13g2_decap_8 FILLER_56_163 ();
 sg13g2_decap_8 FILLER_56_170 ();
 sg13g2_decap_4 FILLER_56_177 ();
 sg13g2_decap_8 FILLER_56_189 ();
 sg13g2_fill_2 FILLER_56_204 ();
 sg13g2_fill_1 FILLER_56_206 ();
 sg13g2_fill_2 FILLER_56_235 ();
 sg13g2_fill_1 FILLER_56_237 ();
 sg13g2_decap_8 FILLER_56_266 ();
 sg13g2_fill_2 FILLER_56_273 ();
 sg13g2_fill_2 FILLER_56_285 ();
 sg13g2_fill_1 FILLER_56_317 ();
 sg13g2_fill_2 FILLER_56_333 ();
 sg13g2_fill_1 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_340 ();
 sg13g2_decap_8 FILLER_56_345 ();
 sg13g2_decap_8 FILLER_56_352 ();
 sg13g2_fill_2 FILLER_56_363 ();
 sg13g2_fill_1 FILLER_56_370 ();
 sg13g2_fill_1 FILLER_56_389 ();
 sg13g2_fill_1 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_436 ();
 sg13g2_decap_8 FILLER_56_455 ();
 sg13g2_decap_8 FILLER_56_462 ();
 sg13g2_fill_2 FILLER_56_469 ();
 sg13g2_decap_8 FILLER_56_501 ();
 sg13g2_decap_4 FILLER_56_508 ();
 sg13g2_fill_1 FILLER_56_515 ();
 sg13g2_decap_8 FILLER_56_531 ();
 sg13g2_decap_8 FILLER_56_538 ();
 sg13g2_decap_4 FILLER_56_545 ();
 sg13g2_fill_2 FILLER_56_549 ();
 sg13g2_decap_4 FILLER_56_580 ();
 sg13g2_decap_4 FILLER_56_592 ();
 sg13g2_decap_8 FILLER_56_610 ();
 sg13g2_fill_2 FILLER_56_617 ();
 sg13g2_fill_2 FILLER_56_634 ();
 sg13g2_fill_1 FILLER_56_636 ();
 sg13g2_fill_1 FILLER_56_645 ();
 sg13g2_fill_1 FILLER_56_654 ();
 sg13g2_fill_2 FILLER_56_663 ();
 sg13g2_fill_1 FILLER_56_701 ();
 sg13g2_fill_2 FILLER_56_712 ();
 sg13g2_decap_8 FILLER_56_734 ();
 sg13g2_fill_2 FILLER_56_741 ();
 sg13g2_fill_1 FILLER_56_743 ();
 sg13g2_fill_1 FILLER_56_774 ();
 sg13g2_fill_1 FILLER_56_780 ();
 sg13g2_fill_2 FILLER_56_807 ();
 sg13g2_decap_4 FILLER_56_814 ();
 sg13g2_fill_2 FILLER_56_818 ();
 sg13g2_decap_8 FILLER_56_824 ();
 sg13g2_fill_2 FILLER_56_847 ();
 sg13g2_fill_1 FILLER_56_886 ();
 sg13g2_decap_4 FILLER_56_891 ();
 sg13g2_fill_2 FILLER_56_895 ();
 sg13g2_decap_4 FILLER_56_911 ();
 sg13g2_decap_4 FILLER_56_921 ();
 sg13g2_fill_2 FILLER_56_925 ();
 sg13g2_fill_2 FILLER_56_948 ();
 sg13g2_fill_1 FILLER_56_950 ();
 sg13g2_fill_1 FILLER_56_959 ();
 sg13g2_decap_8 FILLER_56_973 ();
 sg13g2_decap_8 FILLER_56_980 ();
 sg13g2_fill_1 FILLER_56_987 ();
 sg13g2_fill_2 FILLER_56_996 ();
 sg13g2_fill_1 FILLER_56_1051 ();
 sg13g2_decap_8 FILLER_56_1073 ();
 sg13g2_fill_2 FILLER_56_1080 ();
 sg13g2_fill_1 FILLER_56_1096 ();
 sg13g2_fill_1 FILLER_56_1101 ();
 sg13g2_fill_1 FILLER_56_1105 ();
 sg13g2_fill_1 FILLER_56_1116 ();
 sg13g2_fill_1 FILLER_56_1121 ();
 sg13g2_fill_1 FILLER_56_1127 ();
 sg13g2_fill_2 FILLER_56_1132 ();
 sg13g2_decap_4 FILLER_56_1141 ();
 sg13g2_fill_2 FILLER_56_1148 ();
 sg13g2_fill_1 FILLER_56_1182 ();
 sg13g2_fill_1 FILLER_56_1187 ();
 sg13g2_decap_8 FILLER_56_1196 ();
 sg13g2_fill_2 FILLER_56_1203 ();
 sg13g2_decap_4 FILLER_56_1214 ();
 sg13g2_fill_2 FILLER_56_1218 ();
 sg13g2_fill_2 FILLER_56_1224 ();
 sg13g2_fill_1 FILLER_56_1226 ();
 sg13g2_fill_2 FILLER_56_1232 ();
 sg13g2_fill_1 FILLER_56_1234 ();
 sg13g2_fill_2 FILLER_56_1240 ();
 sg13g2_decap_4 FILLER_56_1265 ();
 sg13g2_fill_1 FILLER_56_1269 ();
 sg13g2_fill_1 FILLER_56_1288 ();
 sg13g2_fill_1 FILLER_56_1309 ();
 sg13g2_fill_2 FILLER_56_1316 ();
 sg13g2_fill_2 FILLER_56_1335 ();
 sg13g2_fill_2 FILLER_56_1370 ();
 sg13g2_fill_2 FILLER_56_1377 ();
 sg13g2_fill_1 FILLER_56_1379 ();
 sg13g2_fill_1 FILLER_56_1424 ();
 sg13g2_fill_1 FILLER_56_1430 ();
 sg13g2_fill_2 FILLER_56_1436 ();
 sg13g2_fill_1 FILLER_56_1443 ();
 sg13g2_fill_2 FILLER_56_1462 ();
 sg13g2_fill_2 FILLER_56_1470 ();
 sg13g2_fill_1 FILLER_56_1481 ();
 sg13g2_fill_2 FILLER_56_1490 ();
 sg13g2_fill_2 FILLER_56_1498 ();
 sg13g2_fill_2 FILLER_56_1514 ();
 sg13g2_fill_2 FILLER_56_1520 ();
 sg13g2_fill_1 FILLER_56_1522 ();
 sg13g2_fill_1 FILLER_56_1528 ();
 sg13g2_decap_8 FILLER_56_1550 ();
 sg13g2_fill_2 FILLER_56_1557 ();
 sg13g2_decap_4 FILLER_56_1576 ();
 sg13g2_decap_4 FILLER_56_1614 ();
 sg13g2_decap_4 FILLER_56_1623 ();
 sg13g2_fill_1 FILLER_56_1627 ();
 sg13g2_fill_1 FILLER_56_1635 ();
 sg13g2_fill_2 FILLER_56_1649 ();
 sg13g2_fill_2 FILLER_56_1671 ();
 sg13g2_fill_1 FILLER_56_1702 ();
 sg13g2_fill_1 FILLER_56_1708 ();
 sg13g2_fill_2 FILLER_56_1714 ();
 sg13g2_fill_2 FILLER_56_1724 ();
 sg13g2_decap_8 FILLER_56_1733 ();
 sg13g2_decap_8 FILLER_56_1740 ();
 sg13g2_decap_8 FILLER_56_1747 ();
 sg13g2_decap_8 FILLER_56_1754 ();
 sg13g2_decap_8 FILLER_56_1761 ();
 sg13g2_decap_4 FILLER_56_1768 ();
 sg13g2_fill_2 FILLER_56_1772 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_4 ();
 sg13g2_fill_1 FILLER_57_21 ();
 sg13g2_fill_2 FILLER_57_27 ();
 sg13g2_fill_1 FILLER_57_39 ();
 sg13g2_fill_2 FILLER_57_49 ();
 sg13g2_fill_1 FILLER_57_51 ();
 sg13g2_decap_4 FILLER_57_57 ();
 sg13g2_fill_2 FILLER_57_61 ();
 sg13g2_fill_2 FILLER_57_78 ();
 sg13g2_decap_8 FILLER_57_107 ();
 sg13g2_decap_4 FILLER_57_114 ();
 sg13g2_fill_2 FILLER_57_118 ();
 sg13g2_fill_2 FILLER_57_125 ();
 sg13g2_fill_2 FILLER_57_132 ();
 sg13g2_fill_1 FILLER_57_146 ();
 sg13g2_decap_8 FILLER_57_152 ();
 sg13g2_decap_8 FILLER_57_159 ();
 sg13g2_decap_8 FILLER_57_166 ();
 sg13g2_fill_2 FILLER_57_173 ();
 sg13g2_fill_2 FILLER_57_193 ();
 sg13g2_fill_1 FILLER_57_195 ();
 sg13g2_fill_2 FILLER_57_204 ();
 sg13g2_fill_1 FILLER_57_206 ();
 sg13g2_fill_1 FILLER_57_220 ();
 sg13g2_decap_8 FILLER_57_260 ();
 sg13g2_decap_8 FILLER_57_267 ();
 sg13g2_decap_4 FILLER_57_274 ();
 sg13g2_fill_1 FILLER_57_278 ();
 sg13g2_decap_4 FILLER_57_301 ();
 sg13g2_fill_1 FILLER_57_305 ();
 sg13g2_decap_8 FILLER_57_310 ();
 sg13g2_decap_4 FILLER_57_317 ();
 sg13g2_fill_1 FILLER_57_321 ();
 sg13g2_fill_1 FILLER_57_340 ();
 sg13g2_decap_4 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_fill_1 FILLER_57_389 ();
 sg13g2_fill_2 FILLER_57_400 ();
 sg13g2_fill_1 FILLER_57_452 ();
 sg13g2_decap_8 FILLER_57_457 ();
 sg13g2_decap_4 FILLER_57_464 ();
 sg13g2_fill_2 FILLER_57_468 ();
 sg13g2_decap_4 FILLER_57_478 ();
 sg13g2_fill_1 FILLER_57_482 ();
 sg13g2_fill_2 FILLER_57_488 ();
 sg13g2_fill_1 FILLER_57_490 ();
 sg13g2_decap_8 FILLER_57_495 ();
 sg13g2_fill_2 FILLER_57_506 ();
 sg13g2_fill_2 FILLER_57_526 ();
 sg13g2_decap_4 FILLER_57_545 ();
 sg13g2_fill_2 FILLER_57_557 ();
 sg13g2_fill_1 FILLER_57_566 ();
 sg13g2_fill_1 FILLER_57_572 ();
 sg13g2_fill_2 FILLER_57_591 ();
 sg13g2_fill_1 FILLER_57_593 ();
 sg13g2_fill_1 FILLER_57_598 ();
 sg13g2_decap_8 FILLER_57_607 ();
 sg13g2_fill_2 FILLER_57_614 ();
 sg13g2_fill_1 FILLER_57_616 ();
 sg13g2_fill_1 FILLER_57_624 ();
 sg13g2_fill_1 FILLER_57_638 ();
 sg13g2_decap_4 FILLER_57_643 ();
 sg13g2_fill_2 FILLER_57_661 ();
 sg13g2_decap_8 FILLER_57_694 ();
 sg13g2_fill_1 FILLER_57_701 ();
 sg13g2_decap_4 FILLER_57_711 ();
 sg13g2_decap_8 FILLER_57_719 ();
 sg13g2_fill_1 FILLER_57_726 ();
 sg13g2_decap_4 FILLER_57_743 ();
 sg13g2_fill_1 FILLER_57_747 ();
 sg13g2_decap_8 FILLER_57_752 ();
 sg13g2_fill_2 FILLER_57_759 ();
 sg13g2_decap_8 FILLER_57_771 ();
 sg13g2_decap_4 FILLER_57_825 ();
 sg13g2_fill_2 FILLER_57_829 ();
 sg13g2_decap_8 FILLER_57_843 ();
 sg13g2_decap_8 FILLER_57_850 ();
 sg13g2_decap_4 FILLER_57_857 ();
 sg13g2_fill_2 FILLER_57_883 ();
 sg13g2_decap_8 FILLER_57_890 ();
 sg13g2_decap_8 FILLER_57_903 ();
 sg13g2_decap_8 FILLER_57_910 ();
 sg13g2_fill_1 FILLER_57_922 ();
 sg13g2_fill_1 FILLER_57_927 ();
 sg13g2_fill_2 FILLER_57_936 ();
 sg13g2_fill_1 FILLER_57_938 ();
 sg13g2_fill_1 FILLER_57_944 ();
 sg13g2_decap_8 FILLER_57_950 ();
 sg13g2_fill_1 FILLER_57_957 ();
 sg13g2_decap_8 FILLER_57_966 ();
 sg13g2_decap_4 FILLER_57_973 ();
 sg13g2_fill_1 FILLER_57_977 ();
 sg13g2_fill_2 FILLER_57_982 ();
 sg13g2_fill_1 FILLER_57_984 ();
 sg13g2_decap_8 FILLER_57_990 ();
 sg13g2_fill_1 FILLER_57_997 ();
 sg13g2_decap_8 FILLER_57_1003 ();
 sg13g2_decap_8 FILLER_57_1010 ();
 sg13g2_fill_1 FILLER_57_1023 ();
 sg13g2_fill_1 FILLER_57_1051 ();
 sg13g2_fill_2 FILLER_57_1087 ();
 sg13g2_fill_1 FILLER_57_1089 ();
 sg13g2_fill_2 FILLER_57_1100 ();
 sg13g2_fill_2 FILLER_57_1127 ();
 sg13g2_decap_4 FILLER_57_1140 ();
 sg13g2_fill_1 FILLER_57_1144 ();
 sg13g2_decap_8 FILLER_57_1149 ();
 sg13g2_fill_2 FILLER_57_1156 ();
 sg13g2_fill_1 FILLER_57_1158 ();
 sg13g2_decap_4 FILLER_57_1164 ();
 sg13g2_fill_1 FILLER_57_1172 ();
 sg13g2_decap_4 FILLER_57_1201 ();
 sg13g2_fill_2 FILLER_57_1219 ();
 sg13g2_fill_1 FILLER_57_1221 ();
 sg13g2_decap_8 FILLER_57_1226 ();
 sg13g2_fill_2 FILLER_57_1249 ();
 sg13g2_fill_2 FILLER_57_1255 ();
 sg13g2_fill_2 FILLER_57_1265 ();
 sg13g2_fill_1 FILLER_57_1267 ();
 sg13g2_fill_2 FILLER_57_1273 ();
 sg13g2_fill_1 FILLER_57_1286 ();
 sg13g2_fill_2 FILLER_57_1301 ();
 sg13g2_fill_2 FILLER_57_1306 ();
 sg13g2_fill_1 FILLER_57_1330 ();
 sg13g2_decap_4 FILLER_57_1373 ();
 sg13g2_fill_1 FILLER_57_1388 ();
 sg13g2_fill_1 FILLER_57_1398 ();
 sg13g2_decap_4 FILLER_57_1406 ();
 sg13g2_fill_2 FILLER_57_1436 ();
 sg13g2_fill_2 FILLER_57_1442 ();
 sg13g2_fill_1 FILLER_57_1444 ();
 sg13g2_decap_8 FILLER_57_1450 ();
 sg13g2_decap_4 FILLER_57_1457 ();
 sg13g2_fill_2 FILLER_57_1466 ();
 sg13g2_decap_4 FILLER_57_1516 ();
 sg13g2_fill_1 FILLER_57_1520 ();
 sg13g2_fill_2 FILLER_57_1526 ();
 sg13g2_decap_4 FILLER_57_1554 ();
 sg13g2_fill_2 FILLER_57_1558 ();
 sg13g2_decap_8 FILLER_57_1578 ();
 sg13g2_decap_8 FILLER_57_1585 ();
 sg13g2_decap_8 FILLER_57_1592 ();
 sg13g2_decap_4 FILLER_57_1599 ();
 sg13g2_fill_2 FILLER_57_1603 ();
 sg13g2_decap_8 FILLER_57_1609 ();
 sg13g2_decap_4 FILLER_57_1628 ();
 sg13g2_fill_1 FILLER_57_1632 ();
 sg13g2_decap_4 FILLER_57_1641 ();
 sg13g2_fill_1 FILLER_57_1645 ();
 sg13g2_fill_1 FILLER_57_1667 ();
 sg13g2_fill_1 FILLER_57_1672 ();
 sg13g2_fill_1 FILLER_57_1678 ();
 sg13g2_fill_2 FILLER_57_1692 ();
 sg13g2_fill_1 FILLER_57_1709 ();
 sg13g2_decap_8 FILLER_57_1720 ();
 sg13g2_fill_1 FILLER_57_1727 ();
 sg13g2_decap_8 FILLER_57_1737 ();
 sg13g2_decap_8 FILLER_57_1744 ();
 sg13g2_decap_8 FILLER_57_1751 ();
 sg13g2_decap_8 FILLER_57_1758 ();
 sg13g2_decap_8 FILLER_57_1765 ();
 sg13g2_fill_2 FILLER_57_1772 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_9 ();
 sg13g2_decap_8 FILLER_58_27 ();
 sg13g2_fill_1 FILLER_58_38 ();
 sg13g2_decap_4 FILLER_58_54 ();
 sg13g2_fill_1 FILLER_58_58 ();
 sg13g2_decap_4 FILLER_58_64 ();
 sg13g2_decap_8 FILLER_58_80 ();
 sg13g2_decap_4 FILLER_58_91 ();
 sg13g2_fill_2 FILLER_58_95 ();
 sg13g2_decap_8 FILLER_58_102 ();
 sg13g2_decap_4 FILLER_58_109 ();
 sg13g2_fill_1 FILLER_58_113 ();
 sg13g2_decap_8 FILLER_58_124 ();
 sg13g2_fill_1 FILLER_58_131 ();
 sg13g2_fill_1 FILLER_58_139 ();
 sg13g2_decap_4 FILLER_58_159 ();
 sg13g2_fill_1 FILLER_58_163 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_fill_1 FILLER_58_175 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_decap_4 FILLER_58_194 ();
 sg13g2_fill_2 FILLER_58_198 ();
 sg13g2_fill_1 FILLER_58_226 ();
 sg13g2_fill_1 FILLER_58_232 ();
 sg13g2_fill_2 FILLER_58_241 ();
 sg13g2_fill_2 FILLER_58_251 ();
 sg13g2_fill_1 FILLER_58_261 ();
 sg13g2_fill_2 FILLER_58_267 ();
 sg13g2_fill_2 FILLER_58_276 ();
 sg13g2_fill_2 FILLER_58_283 ();
 sg13g2_fill_1 FILLER_58_285 ();
 sg13g2_decap_8 FILLER_58_290 ();
 sg13g2_fill_2 FILLER_58_297 ();
 sg13g2_fill_2 FILLER_58_303 ();
 sg13g2_decap_8 FILLER_58_309 ();
 sg13g2_decap_4 FILLER_58_316 ();
 sg13g2_fill_2 FILLER_58_320 ();
 sg13g2_decap_4 FILLER_58_327 ();
 sg13g2_decap_8 FILLER_58_345 ();
 sg13g2_fill_2 FILLER_58_352 ();
 sg13g2_fill_2 FILLER_58_399 ();
 sg13g2_decap_8 FILLER_58_416 ();
 sg13g2_fill_1 FILLER_58_423 ();
 sg13g2_fill_1 FILLER_58_436 ();
 sg13g2_fill_1 FILLER_58_446 ();
 sg13g2_fill_2 FILLER_58_457 ();
 sg13g2_decap_4 FILLER_58_471 ();
 sg13g2_fill_2 FILLER_58_475 ();
 sg13g2_fill_2 FILLER_58_485 ();
 sg13g2_decap_4 FILLER_58_492 ();
 sg13g2_fill_2 FILLER_58_496 ();
 sg13g2_fill_1 FILLER_58_503 ();
 sg13g2_fill_2 FILLER_58_523 ();
 sg13g2_fill_1 FILLER_58_567 ();
 sg13g2_decap_8 FILLER_58_590 ();
 sg13g2_fill_2 FILLER_58_597 ();
 sg13g2_fill_1 FILLER_58_599 ();
 sg13g2_fill_2 FILLER_58_606 ();
 sg13g2_fill_1 FILLER_58_608 ();
 sg13g2_decap_8 FILLER_58_612 ();
 sg13g2_decap_8 FILLER_58_619 ();
 sg13g2_fill_1 FILLER_58_626 ();
 sg13g2_decap_8 FILLER_58_637 ();
 sg13g2_decap_4 FILLER_58_644 ();
 sg13g2_fill_1 FILLER_58_648 ();
 sg13g2_decap_4 FILLER_58_677 ();
 sg13g2_decap_4 FILLER_58_736 ();
 sg13g2_fill_2 FILLER_58_740 ();
 sg13g2_fill_2 FILLER_58_751 ();
 sg13g2_decap_8 FILLER_58_758 ();
 sg13g2_decap_8 FILLER_58_765 ();
 sg13g2_fill_2 FILLER_58_772 ();
 sg13g2_decap_8 FILLER_58_778 ();
 sg13g2_decap_8 FILLER_58_785 ();
 sg13g2_decap_4 FILLER_58_792 ();
 sg13g2_fill_1 FILLER_58_796 ();
 sg13g2_fill_2 FILLER_58_801 ();
 sg13g2_fill_1 FILLER_58_803 ();
 sg13g2_decap_8 FILLER_58_809 ();
 sg13g2_decap_8 FILLER_58_816 ();
 sg13g2_decap_4 FILLER_58_823 ();
 sg13g2_decap_8 FILLER_58_831 ();
 sg13g2_decap_8 FILLER_58_843 ();
 sg13g2_decap_8 FILLER_58_850 ();
 sg13g2_fill_2 FILLER_58_857 ();
 sg13g2_fill_1 FILLER_58_905 ();
 sg13g2_fill_2 FILLER_58_909 ();
 sg13g2_fill_1 FILLER_58_911 ();
 sg13g2_fill_1 FILLER_58_920 ();
 sg13g2_decap_8 FILLER_58_924 ();
 sg13g2_decap_4 FILLER_58_931 ();
 sg13g2_decap_8 FILLER_58_988 ();
 sg13g2_decap_8 FILLER_58_1003 ();
 sg13g2_fill_2 FILLER_58_1010 ();
 sg13g2_fill_1 FILLER_58_1012 ();
 sg13g2_fill_2 FILLER_58_1034 ();
 sg13g2_fill_2 FILLER_58_1041 ();
 sg13g2_fill_1 FILLER_58_1051 ();
 sg13g2_fill_1 FILLER_58_1066 ();
 sg13g2_fill_1 FILLER_58_1096 ();
 sg13g2_decap_8 FILLER_58_1110 ();
 sg13g2_decap_8 FILLER_58_1117 ();
 sg13g2_fill_2 FILLER_58_1129 ();
 sg13g2_fill_1 FILLER_58_1131 ();
 sg13g2_fill_2 FILLER_58_1143 ();
 sg13g2_fill_1 FILLER_58_1202 ();
 sg13g2_fill_2 FILLER_58_1241 ();
 sg13g2_fill_1 FILLER_58_1243 ();
 sg13g2_decap_8 FILLER_58_1249 ();
 sg13g2_fill_1 FILLER_58_1256 ();
 sg13g2_fill_1 FILLER_58_1262 ();
 sg13g2_fill_2 FILLER_58_1268 ();
 sg13g2_decap_8 FILLER_58_1289 ();
 sg13g2_fill_1 FILLER_58_1309 ();
 sg13g2_fill_1 FILLER_58_1332 ();
 sg13g2_fill_2 FILLER_58_1350 ();
 sg13g2_fill_1 FILLER_58_1364 ();
 sg13g2_fill_1 FILLER_58_1370 ();
 sg13g2_decap_4 FILLER_58_1394 ();
 sg13g2_fill_2 FILLER_58_1398 ();
 sg13g2_decap_8 FILLER_58_1404 ();
 sg13g2_decap_4 FILLER_58_1411 ();
 sg13g2_fill_2 FILLER_58_1425 ();
 sg13g2_fill_1 FILLER_58_1435 ();
 sg13g2_fill_2 FILLER_58_1466 ();
 sg13g2_fill_1 FILLER_58_1492 ();
 sg13g2_fill_1 FILLER_58_1507 ();
 sg13g2_fill_2 FILLER_58_1512 ();
 sg13g2_fill_1 FILLER_58_1528 ();
 sg13g2_fill_1 FILLER_58_1533 ();
 sg13g2_decap_4 FILLER_58_1542 ();
 sg13g2_fill_2 FILLER_58_1546 ();
 sg13g2_fill_1 FILLER_58_1556 ();
 sg13g2_decap_8 FILLER_58_1560 ();
 sg13g2_decap_4 FILLER_58_1573 ();
 sg13g2_decap_8 FILLER_58_1589 ();
 sg13g2_fill_1 FILLER_58_1596 ();
 sg13g2_decap_8 FILLER_58_1601 ();
 sg13g2_decap_4 FILLER_58_1608 ();
 sg13g2_fill_1 FILLER_58_1633 ();
 sg13g2_decap_8 FILLER_58_1642 ();
 sg13g2_decap_8 FILLER_58_1649 ();
 sg13g2_decap_4 FILLER_58_1656 ();
 sg13g2_fill_2 FILLER_58_1678 ();
 sg13g2_fill_1 FILLER_58_1680 ();
 sg13g2_fill_1 FILLER_58_1693 ();
 sg13g2_decap_8 FILLER_58_1707 ();
 sg13g2_fill_2 FILLER_58_1718 ();
 sg13g2_fill_1 FILLER_58_1720 ();
 sg13g2_decap_8 FILLER_58_1743 ();
 sg13g2_decap_8 FILLER_58_1750 ();
 sg13g2_decap_8 FILLER_58_1757 ();
 sg13g2_decap_8 FILLER_58_1764 ();
 sg13g2_fill_2 FILLER_58_1771 ();
 sg13g2_fill_1 FILLER_58_1773 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_38 ();
 sg13g2_decap_8 FILLER_59_45 ();
 sg13g2_decap_4 FILLER_59_52 ();
 sg13g2_fill_2 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_67 ();
 sg13g2_decap_8 FILLER_59_74 ();
 sg13g2_decap_8 FILLER_59_81 ();
 sg13g2_fill_2 FILLER_59_88 ();
 sg13g2_fill_1 FILLER_59_90 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_fill_1 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_124 ();
 sg13g2_decap_8 FILLER_59_131 ();
 sg13g2_fill_2 FILLER_59_138 ();
 sg13g2_fill_1 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_170 ();
 sg13g2_decap_4 FILLER_59_200 ();
 sg13g2_decap_8 FILLER_59_212 ();
 sg13g2_decap_4 FILLER_59_219 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_decap_4 FILLER_59_275 ();
 sg13g2_decap_4 FILLER_59_305 ();
 sg13g2_fill_2 FILLER_59_309 ();
 sg13g2_fill_1 FILLER_59_319 ();
 sg13g2_decap_8 FILLER_59_325 ();
 sg13g2_decap_4 FILLER_59_332 ();
 sg13g2_fill_2 FILLER_59_348 ();
 sg13g2_fill_1 FILLER_59_375 ();
 sg13g2_fill_2 FILLER_59_391 ();
 sg13g2_fill_1 FILLER_59_396 ();
 sg13g2_decap_4 FILLER_59_424 ();
 sg13g2_fill_2 FILLER_59_428 ();
 sg13g2_fill_1 FILLER_59_442 ();
 sg13g2_decap_8 FILLER_59_447 ();
 sg13g2_decap_8 FILLER_59_459 ();
 sg13g2_decap_8 FILLER_59_466 ();
 sg13g2_fill_2 FILLER_59_473 ();
 sg13g2_decap_8 FILLER_59_491 ();
 sg13g2_decap_4 FILLER_59_498 ();
 sg13g2_fill_2 FILLER_59_502 ();
 sg13g2_fill_1 FILLER_59_508 ();
 sg13g2_decap_8 FILLER_59_520 ();
 sg13g2_decap_8 FILLER_59_536 ();
 sg13g2_decap_8 FILLER_59_543 ();
 sg13g2_decap_8 FILLER_59_550 ();
 sg13g2_decap_8 FILLER_59_557 ();
 sg13g2_fill_2 FILLER_59_564 ();
 sg13g2_fill_2 FILLER_59_574 ();
 sg13g2_fill_1 FILLER_59_576 ();
 sg13g2_fill_2 FILLER_59_585 ();
 sg13g2_fill_2 FILLER_59_609 ();
 sg13g2_fill_2 FILLER_59_619 ();
 sg13g2_decap_4 FILLER_59_629 ();
 sg13g2_fill_1 FILLER_59_633 ();
 sg13g2_decap_8 FILLER_59_642 ();
 sg13g2_fill_1 FILLER_59_649 ();
 sg13g2_fill_2 FILLER_59_654 ();
 sg13g2_decap_8 FILLER_59_672 ();
 sg13g2_fill_2 FILLER_59_679 ();
 sg13g2_fill_1 FILLER_59_681 ();
 sg13g2_decap_8 FILLER_59_690 ();
 sg13g2_decap_8 FILLER_59_697 ();
 sg13g2_fill_1 FILLER_59_704 ();
 sg13g2_fill_2 FILLER_59_713 ();
 sg13g2_fill_1 FILLER_59_756 ();
 sg13g2_fill_2 FILLER_59_771 ();
 sg13g2_fill_1 FILLER_59_773 ();
 sg13g2_decap_4 FILLER_59_779 ();
 sg13g2_fill_1 FILLER_59_783 ();
 sg13g2_decap_4 FILLER_59_792 ();
 sg13g2_fill_2 FILLER_59_796 ();
 sg13g2_decap_8 FILLER_59_803 ();
 sg13g2_decap_8 FILLER_59_810 ();
 sg13g2_decap_8 FILLER_59_817 ();
 sg13g2_decap_8 FILLER_59_845 ();
 sg13g2_decap_8 FILLER_59_852 ();
 sg13g2_decap_4 FILLER_59_859 ();
 sg13g2_fill_1 FILLER_59_863 ();
 sg13g2_fill_2 FILLER_59_894 ();
 sg13g2_fill_1 FILLER_59_896 ();
 sg13g2_fill_2 FILLER_59_913 ();
 sg13g2_decap_4 FILLER_59_931 ();
 sg13g2_decap_4 FILLER_59_960 ();
 sg13g2_decap_4 FILLER_59_988 ();
 sg13g2_decap_4 FILLER_59_996 ();
 sg13g2_decap_4 FILLER_59_1009 ();
 sg13g2_fill_1 FILLER_59_1013 ();
 sg13g2_decap_4 FILLER_59_1019 ();
 sg13g2_fill_1 FILLER_59_1023 ();
 sg13g2_decap_8 FILLER_59_1032 ();
 sg13g2_fill_2 FILLER_59_1039 ();
 sg13g2_fill_1 FILLER_59_1041 ();
 sg13g2_fill_2 FILLER_59_1050 ();
 sg13g2_fill_2 FILLER_59_1081 ();
 sg13g2_fill_1 FILLER_59_1083 ();
 sg13g2_fill_2 FILLER_59_1093 ();
 sg13g2_decap_4 FILLER_59_1103 ();
 sg13g2_fill_2 FILLER_59_1107 ();
 sg13g2_decap_8 FILLER_59_1117 ();
 sg13g2_fill_2 FILLER_59_1124 ();
 sg13g2_fill_2 FILLER_59_1145 ();
 sg13g2_decap_8 FILLER_59_1161 ();
 sg13g2_fill_1 FILLER_59_1207 ();
 sg13g2_fill_2 FILLER_59_1212 ();
 sg13g2_fill_1 FILLER_59_1218 ();
 sg13g2_decap_8 FILLER_59_1240 ();
 sg13g2_fill_2 FILLER_59_1247 ();
 sg13g2_fill_1 FILLER_59_1249 ();
 sg13g2_fill_1 FILLER_59_1258 ();
 sg13g2_fill_1 FILLER_59_1264 ();
 sg13g2_decap_4 FILLER_59_1280 ();
 sg13g2_fill_1 FILLER_59_1284 ();
 sg13g2_decap_8 FILLER_59_1292 ();
 sg13g2_fill_2 FILLER_59_1299 ();
 sg13g2_fill_2 FILLER_59_1320 ();
 sg13g2_fill_1 FILLER_59_1353 ();
 sg13g2_fill_2 FILLER_59_1359 ();
 sg13g2_fill_2 FILLER_59_1369 ();
 sg13g2_fill_1 FILLER_59_1371 ();
 sg13g2_fill_2 FILLER_59_1380 ();
 sg13g2_decap_8 FILLER_59_1390 ();
 sg13g2_decap_8 FILLER_59_1402 ();
 sg13g2_fill_1 FILLER_59_1409 ();
 sg13g2_fill_1 FILLER_59_1418 ();
 sg13g2_fill_2 FILLER_59_1435 ();
 sg13g2_fill_1 FILLER_59_1443 ();
 sg13g2_decap_8 FILLER_59_1448 ();
 sg13g2_fill_2 FILLER_59_1455 ();
 sg13g2_decap_4 FILLER_59_1462 ();
 sg13g2_fill_1 FILLER_59_1466 ();
 sg13g2_fill_1 FILLER_59_1512 ();
 sg13g2_decap_8 FILLER_59_1534 ();
 sg13g2_fill_2 FILLER_59_1541 ();
 sg13g2_fill_1 FILLER_59_1543 ();
 sg13g2_decap_8 FILLER_59_1549 ();
 sg13g2_fill_1 FILLER_59_1556 ();
 sg13g2_decap_8 FILLER_59_1562 ();
 sg13g2_fill_2 FILLER_59_1569 ();
 sg13g2_decap_4 FILLER_59_1576 ();
 sg13g2_fill_1 FILLER_59_1580 ();
 sg13g2_decap_8 FILLER_59_1595 ();
 sg13g2_fill_2 FILLER_59_1602 ();
 sg13g2_fill_1 FILLER_59_1604 ();
 sg13g2_fill_2 FILLER_59_1615 ();
 sg13g2_fill_1 FILLER_59_1617 ();
 sg13g2_fill_2 FILLER_59_1623 ();
 sg13g2_fill_1 FILLER_59_1630 ();
 sg13g2_fill_2 FILLER_59_1635 ();
 sg13g2_decap_8 FILLER_59_1642 ();
 sg13g2_fill_2 FILLER_59_1658 ();
 sg13g2_fill_1 FILLER_59_1697 ();
 sg13g2_fill_2 FILLER_59_1708 ();
 sg13g2_fill_2 FILLER_59_1714 ();
 sg13g2_fill_2 FILLER_59_1723 ();
 sg13g2_decap_8 FILLER_59_1729 ();
 sg13g2_decap_8 FILLER_59_1736 ();
 sg13g2_decap_8 FILLER_59_1743 ();
 sg13g2_decap_8 FILLER_59_1750 ();
 sg13g2_decap_8 FILLER_59_1757 ();
 sg13g2_decap_8 FILLER_59_1764 ();
 sg13g2_fill_2 FILLER_59_1771 ();
 sg13g2_fill_1 FILLER_59_1773 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_9 ();
 sg13g2_fill_2 FILLER_60_20 ();
 sg13g2_fill_1 FILLER_60_27 ();
 sg13g2_fill_2 FILLER_60_36 ();
 sg13g2_fill_1 FILLER_60_38 ();
 sg13g2_fill_1 FILLER_60_47 ();
 sg13g2_fill_2 FILLER_60_56 ();
 sg13g2_fill_2 FILLER_60_68 ();
 sg13g2_decap_8 FILLER_60_74 ();
 sg13g2_fill_1 FILLER_60_81 ();
 sg13g2_fill_2 FILLER_60_90 ();
 sg13g2_fill_1 FILLER_60_92 ();
 sg13g2_fill_1 FILLER_60_101 ();
 sg13g2_fill_1 FILLER_60_110 ();
 sg13g2_fill_2 FILLER_60_115 ();
 sg13g2_fill_1 FILLER_60_122 ();
 sg13g2_decap_8 FILLER_60_128 ();
 sg13g2_fill_1 FILLER_60_135 ();
 sg13g2_fill_1 FILLER_60_156 ();
 sg13g2_fill_1 FILLER_60_163 ();
 sg13g2_fill_2 FILLER_60_173 ();
 sg13g2_fill_1 FILLER_60_175 ();
 sg13g2_fill_2 FILLER_60_191 ();
 sg13g2_fill_1 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_199 ();
 sg13g2_fill_2 FILLER_60_219 ();
 sg13g2_fill_1 FILLER_60_221 ();
 sg13g2_decap_8 FILLER_60_235 ();
 sg13g2_fill_2 FILLER_60_242 ();
 sg13g2_decap_8 FILLER_60_256 ();
 sg13g2_decap_8 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_decap_4 FILLER_60_287 ();
 sg13g2_fill_1 FILLER_60_291 ();
 sg13g2_decap_4 FILLER_60_300 ();
 sg13g2_decap_4 FILLER_60_321 ();
 sg13g2_fill_2 FILLER_60_325 ();
 sg13g2_decap_8 FILLER_60_331 ();
 sg13g2_fill_1 FILLER_60_351 ();
 sg13g2_fill_2 FILLER_60_383 ();
 sg13g2_fill_2 FILLER_60_401 ();
 sg13g2_fill_2 FILLER_60_445 ();
 sg13g2_fill_1 FILLER_60_447 ();
 sg13g2_decap_8 FILLER_60_465 ();
 sg13g2_fill_2 FILLER_60_472 ();
 sg13g2_fill_2 FILLER_60_482 ();
 sg13g2_fill_1 FILLER_60_484 ();
 sg13g2_fill_2 FILLER_60_498 ();
 sg13g2_fill_1 FILLER_60_508 ();
 sg13g2_decap_8 FILLER_60_515 ();
 sg13g2_decap_4 FILLER_60_522 ();
 sg13g2_fill_1 FILLER_60_526 ();
 sg13g2_fill_2 FILLER_60_532 ();
 sg13g2_decap_8 FILLER_60_541 ();
 sg13g2_decap_4 FILLER_60_548 ();
 sg13g2_decap_8 FILLER_60_564 ();
 sg13g2_decap_8 FILLER_60_571 ();
 sg13g2_decap_8 FILLER_60_578 ();
 sg13g2_decap_4 FILLER_60_585 ();
 sg13g2_fill_2 FILLER_60_589 ();
 sg13g2_decap_4 FILLER_60_596 ();
 sg13g2_fill_2 FILLER_60_600 ();
 sg13g2_fill_2 FILLER_60_606 ();
 sg13g2_decap_4 FILLER_60_617 ();
 sg13g2_decap_4 FILLER_60_631 ();
 sg13g2_fill_2 FILLER_60_635 ();
 sg13g2_fill_1 FILLER_60_642 ();
 sg13g2_fill_2 FILLER_60_648 ();
 sg13g2_fill_2 FILLER_60_670 ();
 sg13g2_fill_1 FILLER_60_672 ();
 sg13g2_decap_4 FILLER_60_700 ();
 sg13g2_decap_8 FILLER_60_708 ();
 sg13g2_fill_2 FILLER_60_715 ();
 sg13g2_fill_1 FILLER_60_717 ();
 sg13g2_fill_1 FILLER_60_735 ();
 sg13g2_decap_4 FILLER_60_741 ();
 sg13g2_fill_2 FILLER_60_760 ();
 sg13g2_fill_1 FILLER_60_762 ();
 sg13g2_decap_8 FILLER_60_775 ();
 sg13g2_decap_8 FILLER_60_782 ();
 sg13g2_fill_1 FILLER_60_789 ();
 sg13g2_fill_2 FILLER_60_803 ();
 sg13g2_fill_1 FILLER_60_805 ();
 sg13g2_fill_1 FILLER_60_812 ();
 sg13g2_fill_2 FILLER_60_821 ();
 sg13g2_fill_1 FILLER_60_823 ();
 sg13g2_fill_2 FILLER_60_840 ();
 sg13g2_fill_1 FILLER_60_848 ();
 sg13g2_decap_4 FILLER_60_869 ();
 sg13g2_fill_2 FILLER_60_878 ();
 sg13g2_decap_8 FILLER_60_905 ();
 sg13g2_decap_4 FILLER_60_912 ();
 sg13g2_fill_2 FILLER_60_916 ();
 sg13g2_decap_8 FILLER_60_927 ();
 sg13g2_fill_2 FILLER_60_934 ();
 sg13g2_decap_8 FILLER_60_951 ();
 sg13g2_decap_8 FILLER_60_958 ();
 sg13g2_decap_8 FILLER_60_965 ();
 sg13g2_fill_2 FILLER_60_972 ();
 sg13g2_fill_1 FILLER_60_974 ();
 sg13g2_fill_1 FILLER_60_983 ();
 sg13g2_fill_1 FILLER_60_988 ();
 sg13g2_fill_1 FILLER_60_993 ();
 sg13g2_fill_1 FILLER_60_1006 ();
 sg13g2_fill_2 FILLER_60_1017 ();
 sg13g2_decap_4 FILLER_60_1024 ();
 sg13g2_fill_2 FILLER_60_1028 ();
 sg13g2_decap_8 FILLER_60_1034 ();
 sg13g2_decap_4 FILLER_60_1041 ();
 sg13g2_fill_2 FILLER_60_1050 ();
 sg13g2_decap_8 FILLER_60_1066 ();
 sg13g2_decap_4 FILLER_60_1081 ();
 sg13g2_decap_4 FILLER_60_1090 ();
 sg13g2_fill_1 FILLER_60_1117 ();
 sg13g2_decap_4 FILLER_60_1122 ();
 sg13g2_fill_1 FILLER_60_1126 ();
 sg13g2_fill_2 FILLER_60_1131 ();
 sg13g2_fill_2 FILLER_60_1152 ();
 sg13g2_decap_4 FILLER_60_1171 ();
 sg13g2_fill_1 FILLER_60_1175 ();
 sg13g2_fill_2 FILLER_60_1203 ();
 sg13g2_fill_1 FILLER_60_1205 ();
 sg13g2_decap_8 FILLER_60_1232 ();
 sg13g2_decap_8 FILLER_60_1251 ();
 sg13g2_decap_4 FILLER_60_1258 ();
 sg13g2_fill_2 FILLER_60_1262 ();
 sg13g2_decap_4 FILLER_60_1268 ();
 sg13g2_fill_1 FILLER_60_1272 ();
 sg13g2_fill_2 FILLER_60_1283 ();
 sg13g2_fill_2 FILLER_60_1290 ();
 sg13g2_fill_2 FILLER_60_1300 ();
 sg13g2_fill_2 FILLER_60_1309 ();
 sg13g2_decap_4 FILLER_60_1324 ();
 sg13g2_fill_2 FILLER_60_1328 ();
 sg13g2_fill_1 FILLER_60_1364 ();
 sg13g2_decap_4 FILLER_60_1375 ();
 sg13g2_fill_1 FILLER_60_1384 ();
 sg13g2_fill_2 FILLER_60_1413 ();
 sg13g2_fill_1 FILLER_60_1415 ();
 sg13g2_fill_2 FILLER_60_1437 ();
 sg13g2_fill_2 FILLER_60_1452 ();
 sg13g2_fill_1 FILLER_60_1454 ();
 sg13g2_decap_4 FILLER_60_1460 ();
 sg13g2_fill_1 FILLER_60_1464 ();
 sg13g2_fill_2 FILLER_60_1470 ();
 sg13g2_fill_1 FILLER_60_1476 ();
 sg13g2_fill_1 FILLER_60_1481 ();
 sg13g2_fill_1 FILLER_60_1490 ();
 sg13g2_fill_2 FILLER_60_1521 ();
 sg13g2_fill_2 FILLER_60_1553 ();
 sg13g2_fill_1 FILLER_60_1555 ();
 sg13g2_fill_2 FILLER_60_1576 ();
 sg13g2_fill_2 FILLER_60_1595 ();
 sg13g2_fill_2 FILLER_60_1605 ();
 sg13g2_fill_1 FILLER_60_1629 ();
 sg13g2_fill_1 FILLER_60_1635 ();
 sg13g2_decap_8 FILLER_60_1640 ();
 sg13g2_decap_8 FILLER_60_1647 ();
 sg13g2_decap_8 FILLER_60_1654 ();
 sg13g2_decap_8 FILLER_60_1661 ();
 sg13g2_decap_8 FILLER_60_1668 ();
 sg13g2_decap_4 FILLER_60_1675 ();
 sg13g2_decap_4 FILLER_60_1688 ();
 sg13g2_fill_2 FILLER_60_1692 ();
 sg13g2_decap_4 FILLER_60_1697 ();
 sg13g2_fill_2 FILLER_60_1701 ();
 sg13g2_fill_1 FILLER_60_1708 ();
 sg13g2_decap_8 FILLER_60_1713 ();
 sg13g2_decap_8 FILLER_60_1720 ();
 sg13g2_decap_8 FILLER_60_1727 ();
 sg13g2_decap_8 FILLER_60_1734 ();
 sg13g2_decap_8 FILLER_60_1741 ();
 sg13g2_decap_8 FILLER_60_1748 ();
 sg13g2_decap_8 FILLER_60_1755 ();
 sg13g2_decap_8 FILLER_60_1762 ();
 sg13g2_decap_4 FILLER_60_1769 ();
 sg13g2_fill_1 FILLER_60_1773 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_11 ();
 sg13g2_decap_8 FILLER_61_18 ();
 sg13g2_decap_8 FILLER_61_25 ();
 sg13g2_fill_1 FILLER_61_32 ();
 sg13g2_fill_2 FILLER_61_41 ();
 sg13g2_fill_1 FILLER_61_54 ();
 sg13g2_fill_2 FILLER_61_59 ();
 sg13g2_decap_8 FILLER_61_66 ();
 sg13g2_fill_2 FILLER_61_91 ();
 sg13g2_decap_4 FILLER_61_107 ();
 sg13g2_fill_1 FILLER_61_111 ();
 sg13g2_fill_2 FILLER_61_117 ();
 sg13g2_fill_2 FILLER_61_124 ();
 sg13g2_decap_4 FILLER_61_131 ();
 sg13g2_fill_1 FILLER_61_139 ();
 sg13g2_fill_1 FILLER_61_145 ();
 sg13g2_fill_1 FILLER_61_151 ();
 sg13g2_fill_1 FILLER_61_157 ();
 sg13g2_fill_1 FILLER_61_163 ();
 sg13g2_fill_2 FILLER_61_179 ();
 sg13g2_decap_4 FILLER_61_185 ();
 sg13g2_decap_4 FILLER_61_194 ();
 sg13g2_decap_4 FILLER_61_202 ();
 sg13g2_decap_4 FILLER_61_219 ();
 sg13g2_fill_1 FILLER_61_223 ();
 sg13g2_fill_1 FILLER_61_232 ();
 sg13g2_decap_8 FILLER_61_240 ();
 sg13g2_decap_8 FILLER_61_281 ();
 sg13g2_fill_1 FILLER_61_292 ();
 sg13g2_fill_1 FILLER_61_303 ();
 sg13g2_fill_2 FILLER_61_319 ();
 sg13g2_decap_8 FILLER_61_325 ();
 sg13g2_decap_8 FILLER_61_332 ();
 sg13g2_fill_2 FILLER_61_339 ();
 sg13g2_fill_1 FILLER_61_379 ();
 sg13g2_fill_2 FILLER_61_391 ();
 sg13g2_fill_2 FILLER_61_409 ();
 sg13g2_fill_2 FILLER_61_420 ();
 sg13g2_decap_8 FILLER_61_426 ();
 sg13g2_fill_2 FILLER_61_433 ();
 sg13g2_fill_2 FILLER_61_449 ();
 sg13g2_decap_8 FILLER_61_474 ();
 sg13g2_fill_2 FILLER_61_481 ();
 sg13g2_decap_8 FILLER_61_493 ();
 sg13g2_decap_8 FILLER_61_500 ();
 sg13g2_fill_1 FILLER_61_526 ();
 sg13g2_fill_1 FILLER_61_535 ();
 sg13g2_fill_1 FILLER_61_541 ();
 sg13g2_fill_1 FILLER_61_550 ();
 sg13g2_fill_2 FILLER_61_556 ();
 sg13g2_fill_2 FILLER_61_566 ();
 sg13g2_fill_2 FILLER_61_576 ();
 sg13g2_fill_1 FILLER_61_578 ();
 sg13g2_decap_4 FILLER_61_583 ();
 sg13g2_fill_2 FILLER_61_587 ();
 sg13g2_decap_8 FILLER_61_593 ();
 sg13g2_fill_2 FILLER_61_600 ();
 sg13g2_fill_1 FILLER_61_602 ();
 sg13g2_fill_1 FILLER_61_607 ();
 sg13g2_decap_8 FILLER_61_616 ();
 sg13g2_fill_2 FILLER_61_627 ();
 sg13g2_fill_1 FILLER_61_629 ();
 sg13g2_fill_1 FILLER_61_639 ();
 sg13g2_fill_1 FILLER_61_645 ();
 sg13g2_fill_1 FILLER_61_650 ();
 sg13g2_fill_1 FILLER_61_656 ();
 sg13g2_decap_4 FILLER_61_679 ();
 sg13g2_decap_4 FILLER_61_700 ();
 sg13g2_fill_1 FILLER_61_704 ();
 sg13g2_decap_8 FILLER_61_708 ();
 sg13g2_decap_8 FILLER_61_715 ();
 sg13g2_decap_4 FILLER_61_736 ();
 sg13g2_fill_2 FILLER_61_740 ();
 sg13g2_fill_1 FILLER_61_754 ();
 sg13g2_fill_2 FILLER_61_761 ();
 sg13g2_fill_1 FILLER_61_763 ();
 sg13g2_decap_8 FILLER_61_782 ();
 sg13g2_decap_8 FILLER_61_789 ();
 sg13g2_decap_8 FILLER_61_800 ();
 sg13g2_fill_2 FILLER_61_814 ();
 sg13g2_fill_1 FILLER_61_816 ();
 sg13g2_fill_1 FILLER_61_838 ();
 sg13g2_decap_8 FILLER_61_844 ();
 sg13g2_decap_4 FILLER_61_851 ();
 sg13g2_fill_1 FILLER_61_855 ();
 sg13g2_fill_1 FILLER_61_866 ();
 sg13g2_fill_1 FILLER_61_875 ();
 sg13g2_fill_1 FILLER_61_897 ();
 sg13g2_decap_4 FILLER_61_919 ();
 sg13g2_fill_2 FILLER_61_927 ();
 sg13g2_fill_1 FILLER_61_929 ();
 sg13g2_decap_8 FILLER_61_938 ();
 sg13g2_fill_1 FILLER_61_945 ();
 sg13g2_decap_4 FILLER_61_961 ();
 sg13g2_fill_2 FILLER_61_1006 ();
 sg13g2_decap_4 FILLER_61_1025 ();
 sg13g2_decap_8 FILLER_61_1052 ();
 sg13g2_decap_8 FILLER_61_1059 ();
 sg13g2_fill_2 FILLER_61_1066 ();
 sg13g2_fill_2 FILLER_61_1089 ();
 sg13g2_fill_1 FILLER_61_1104 ();
 sg13g2_fill_1 FILLER_61_1110 ();
 sg13g2_fill_1 FILLER_61_1117 ();
 sg13g2_fill_2 FILLER_61_1123 ();
 sg13g2_decap_4 FILLER_61_1135 ();
 sg13g2_fill_2 FILLER_61_1139 ();
 sg13g2_fill_2 FILLER_61_1162 ();
 sg13g2_fill_1 FILLER_61_1168 ();
 sg13g2_fill_1 FILLER_61_1181 ();
 sg13g2_fill_2 FILLER_61_1217 ();
 sg13g2_decap_8 FILLER_61_1228 ();
 sg13g2_decap_8 FILLER_61_1235 ();
 sg13g2_fill_2 FILLER_61_1242 ();
 sg13g2_decap_8 FILLER_61_1249 ();
 sg13g2_decap_8 FILLER_61_1256 ();
 sg13g2_decap_8 FILLER_61_1263 ();
 sg13g2_fill_1 FILLER_61_1270 ();
 sg13g2_decap_4 FILLER_61_1276 ();
 sg13g2_fill_1 FILLER_61_1280 ();
 sg13g2_fill_2 FILLER_61_1294 ();
 sg13g2_fill_1 FILLER_61_1312 ();
 sg13g2_fill_1 FILLER_61_1323 ();
 sg13g2_fill_1 FILLER_61_1329 ();
 sg13g2_decap_4 FILLER_61_1335 ();
 sg13g2_fill_2 FILLER_61_1339 ();
 sg13g2_decap_4 FILLER_61_1345 ();
 sg13g2_fill_1 FILLER_61_1349 ();
 sg13g2_decap_4 FILLER_61_1355 ();
 sg13g2_fill_1 FILLER_61_1359 ();
 sg13g2_fill_1 FILLER_61_1365 ();
 sg13g2_decap_4 FILLER_61_1375 ();
 sg13g2_fill_2 FILLER_61_1384 ();
 sg13g2_fill_1 FILLER_61_1386 ();
 sg13g2_fill_2 FILLER_61_1401 ();
 sg13g2_decap_8 FILLER_61_1407 ();
 sg13g2_decap_4 FILLER_61_1414 ();
 sg13g2_fill_1 FILLER_61_1418 ();
 sg13g2_decap_4 FILLER_61_1422 ();
 sg13g2_fill_1 FILLER_61_1439 ();
 sg13g2_fill_2 FILLER_61_1446 ();
 sg13g2_fill_1 FILLER_61_1448 ();
 sg13g2_decap_8 FILLER_61_1473 ();
 sg13g2_decap_4 FILLER_61_1480 ();
 sg13g2_fill_2 FILLER_61_1518 ();
 sg13g2_fill_2 FILLER_61_1536 ();
 sg13g2_fill_1 FILLER_61_1542 ();
 sg13g2_fill_2 FILLER_61_1548 ();
 sg13g2_fill_1 FILLER_61_1550 ();
 sg13g2_decap_8 FILLER_61_1556 ();
 sg13g2_fill_1 FILLER_61_1563 ();
 sg13g2_fill_1 FILLER_61_1576 ();
 sg13g2_fill_1 FILLER_61_1581 ();
 sg13g2_fill_2 FILLER_61_1596 ();
 sg13g2_fill_1 FILLER_61_1598 ();
 sg13g2_decap_4 FILLER_61_1604 ();
 sg13g2_fill_2 FILLER_61_1623 ();
 sg13g2_decap_8 FILLER_61_1629 ();
 sg13g2_fill_1 FILLER_61_1654 ();
 sg13g2_decap_8 FILLER_61_1660 ();
 sg13g2_decap_4 FILLER_61_1667 ();
 sg13g2_decap_4 FILLER_61_1679 ();
 sg13g2_fill_2 FILLER_61_1683 ();
 sg13g2_decap_8 FILLER_61_1715 ();
 sg13g2_decap_8 FILLER_61_1722 ();
 sg13g2_decap_8 FILLER_61_1729 ();
 sg13g2_decap_8 FILLER_61_1736 ();
 sg13g2_decap_8 FILLER_61_1743 ();
 sg13g2_decap_8 FILLER_61_1750 ();
 sg13g2_decap_8 FILLER_61_1757 ();
 sg13g2_decap_8 FILLER_61_1764 ();
 sg13g2_fill_2 FILLER_61_1771 ();
 sg13g2_fill_1 FILLER_61_1773 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_20 ();
 sg13g2_fill_2 FILLER_62_27 ();
 sg13g2_fill_2 FILLER_62_39 ();
 sg13g2_decap_4 FILLER_62_60 ();
 sg13g2_fill_2 FILLER_62_88 ();
 sg13g2_fill_1 FILLER_62_90 ();
 sg13g2_fill_1 FILLER_62_95 ();
 sg13g2_fill_1 FILLER_62_108 ();
 sg13g2_decap_8 FILLER_62_125 ();
 sg13g2_decap_8 FILLER_62_162 ();
 sg13g2_fill_1 FILLER_62_169 ();
 sg13g2_fill_1 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_201 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_fill_2 FILLER_62_225 ();
 sg13g2_fill_1 FILLER_62_227 ();
 sg13g2_fill_1 FILLER_62_233 ();
 sg13g2_fill_1 FILLER_62_242 ();
 sg13g2_fill_1 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_fill_1 FILLER_62_273 ();
 sg13g2_decap_4 FILLER_62_279 ();
 sg13g2_fill_1 FILLER_62_283 ();
 sg13g2_decap_4 FILLER_62_289 ();
 sg13g2_fill_1 FILLER_62_293 ();
 sg13g2_fill_1 FILLER_62_319 ();
 sg13g2_fill_2 FILLER_62_325 ();
 sg13g2_fill_1 FILLER_62_327 ();
 sg13g2_decap_8 FILLER_62_333 ();
 sg13g2_decap_8 FILLER_62_340 ();
 sg13g2_fill_1 FILLER_62_347 ();
 sg13g2_fill_2 FILLER_62_358 ();
 sg13g2_fill_1 FILLER_62_378 ();
 sg13g2_fill_2 FILLER_62_400 ();
 sg13g2_fill_2 FILLER_62_412 ();
 sg13g2_decap_8 FILLER_62_426 ();
 sg13g2_fill_2 FILLER_62_433 ();
 sg13g2_fill_1 FILLER_62_435 ();
 sg13g2_decap_4 FILLER_62_441 ();
 sg13g2_decap_8 FILLER_62_449 ();
 sg13g2_fill_1 FILLER_62_456 ();
 sg13g2_decap_4 FILLER_62_462 ();
 sg13g2_fill_2 FILLER_62_466 ();
 sg13g2_fill_2 FILLER_62_485 ();
 sg13g2_decap_8 FILLER_62_495 ();
 sg13g2_decap_8 FILLER_62_502 ();
 sg13g2_fill_2 FILLER_62_509 ();
 sg13g2_fill_1 FILLER_62_511 ();
 sg13g2_fill_1 FILLER_62_516 ();
 sg13g2_decap_4 FILLER_62_535 ();
 sg13g2_decap_8 FILLER_62_547 ();
 sg13g2_fill_2 FILLER_62_554 ();
 sg13g2_decap_8 FILLER_62_564 ();
 sg13g2_decap_8 FILLER_62_598 ();
 sg13g2_decap_8 FILLER_62_605 ();
 sg13g2_fill_2 FILLER_62_612 ();
 sg13g2_fill_2 FILLER_62_618 ();
 sg13g2_decap_8 FILLER_62_631 ();
 sg13g2_fill_2 FILLER_62_638 ();
 sg13g2_fill_1 FILLER_62_640 ();
 sg13g2_fill_1 FILLER_62_645 ();
 sg13g2_decap_4 FILLER_62_658 ();
 sg13g2_fill_1 FILLER_62_662 ();
 sg13g2_decap_4 FILLER_62_669 ();
 sg13g2_fill_1 FILLER_62_678 ();
 sg13g2_decap_8 FILLER_62_694 ();
 sg13g2_decap_8 FILLER_62_701 ();
 sg13g2_decap_8 FILLER_62_708 ();
 sg13g2_decap_4 FILLER_62_715 ();
 sg13g2_fill_1 FILLER_62_719 ();
 sg13g2_fill_2 FILLER_62_735 ();
 sg13g2_fill_1 FILLER_62_743 ();
 sg13g2_decap_8 FILLER_62_782 ();
 sg13g2_fill_2 FILLER_62_789 ();
 sg13g2_fill_1 FILLER_62_791 ();
 sg13g2_decap_4 FILLER_62_796 ();
 sg13g2_decap_8 FILLER_62_804 ();
 sg13g2_fill_2 FILLER_62_811 ();
 sg13g2_fill_1 FILLER_62_813 ();
 sg13g2_decap_4 FILLER_62_823 ();
 sg13g2_fill_2 FILLER_62_859 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_4 FILLER_62_875 ();
 sg13g2_fill_1 FILLER_62_884 ();
 sg13g2_fill_1 FILLER_62_889 ();
 sg13g2_fill_2 FILLER_62_902 ();
 sg13g2_fill_1 FILLER_62_904 ();
 sg13g2_decap_8 FILLER_62_926 ();
 sg13g2_fill_1 FILLER_62_933 ();
 sg13g2_decap_4 FILLER_62_939 ();
 sg13g2_decap_8 FILLER_62_947 ();
 sg13g2_decap_8 FILLER_62_954 ();
 sg13g2_decap_4 FILLER_62_961 ();
 sg13g2_fill_1 FILLER_62_965 ();
 sg13g2_decap_8 FILLER_62_976 ();
 sg13g2_fill_2 FILLER_62_983 ();
 sg13g2_fill_1 FILLER_62_985 ();
 sg13g2_decap_4 FILLER_62_1000 ();
 sg13g2_decap_8 FILLER_62_1012 ();
 sg13g2_decap_8 FILLER_62_1019 ();
 sg13g2_decap_8 FILLER_62_1026 ();
 sg13g2_decap_4 FILLER_62_1033 ();
 sg13g2_fill_2 FILLER_62_1037 ();
 sg13g2_fill_2 FILLER_62_1044 ();
 sg13g2_decap_4 FILLER_62_1064 ();
 sg13g2_fill_1 FILLER_62_1078 ();
 sg13g2_decap_8 FILLER_62_1086 ();
 sg13g2_decap_4 FILLER_62_1093 ();
 sg13g2_fill_1 FILLER_62_1102 ();
 sg13g2_decap_8 FILLER_62_1113 ();
 sg13g2_fill_2 FILLER_62_1120 ();
 sg13g2_fill_1 FILLER_62_1122 ();
 sg13g2_decap_8 FILLER_62_1138 ();
 sg13g2_fill_2 FILLER_62_1145 ();
 sg13g2_fill_1 FILLER_62_1147 ();
 sg13g2_decap_8 FILLER_62_1156 ();
 sg13g2_decap_4 FILLER_62_1163 ();
 sg13g2_fill_1 FILLER_62_1167 ();
 sg13g2_fill_2 FILLER_62_1177 ();
 sg13g2_decap_4 FILLER_62_1188 ();
 sg13g2_fill_1 FILLER_62_1192 ();
 sg13g2_fill_2 FILLER_62_1218 ();
 sg13g2_decap_8 FILLER_62_1228 ();
 sg13g2_fill_2 FILLER_62_1235 ();
 sg13g2_decap_8 FILLER_62_1245 ();
 sg13g2_fill_2 FILLER_62_1252 ();
 sg13g2_fill_1 FILLER_62_1258 ();
 sg13g2_decap_4 FILLER_62_1288 ();
 sg13g2_fill_2 FILLER_62_1296 ();
 sg13g2_fill_2 FILLER_62_1303 ();
 sg13g2_fill_1 FILLER_62_1311 ();
 sg13g2_fill_2 FILLER_62_1322 ();
 sg13g2_fill_1 FILLER_62_1324 ();
 sg13g2_decap_8 FILLER_62_1330 ();
 sg13g2_decap_8 FILLER_62_1337 ();
 sg13g2_decap_8 FILLER_62_1344 ();
 sg13g2_fill_2 FILLER_62_1362 ();
 sg13g2_fill_1 FILLER_62_1364 ();
 sg13g2_decap_8 FILLER_62_1410 ();
 sg13g2_fill_2 FILLER_62_1417 ();
 sg13g2_fill_1 FILLER_62_1419 ();
 sg13g2_fill_2 FILLER_62_1442 ();
 sg13g2_fill_1 FILLER_62_1476 ();
 sg13g2_fill_1 FILLER_62_1481 ();
 sg13g2_fill_2 FILLER_62_1494 ();
 sg13g2_fill_1 FILLER_62_1496 ();
 sg13g2_decap_4 FILLER_62_1529 ();
 sg13g2_decap_4 FILLER_62_1538 ();
 sg13g2_decap_8 FILLER_62_1546 ();
 sg13g2_decap_4 FILLER_62_1553 ();
 sg13g2_fill_1 FILLER_62_1571 ();
 sg13g2_fill_2 FILLER_62_1610 ();
 sg13g2_decap_8 FILLER_62_1622 ();
 sg13g2_fill_2 FILLER_62_1629 ();
 sg13g2_fill_1 FILLER_62_1631 ();
 sg13g2_fill_1 FILLER_62_1645 ();
 sg13g2_fill_2 FILLER_62_1662 ();
 sg13g2_fill_2 FILLER_62_1694 ();
 sg13g2_fill_1 FILLER_62_1696 ();
 sg13g2_decap_8 FILLER_62_1701 ();
 sg13g2_decap_8 FILLER_62_1713 ();
 sg13g2_fill_1 FILLER_62_1720 ();
 sg13g2_decap_8 FILLER_62_1724 ();
 sg13g2_decap_8 FILLER_62_1731 ();
 sg13g2_decap_8 FILLER_62_1738 ();
 sg13g2_decap_8 FILLER_62_1745 ();
 sg13g2_decap_8 FILLER_62_1752 ();
 sg13g2_decap_8 FILLER_62_1759 ();
 sg13g2_decap_8 FILLER_62_1766 ();
 sg13g2_fill_1 FILLER_62_1773 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_28 ();
 sg13g2_fill_1 FILLER_63_30 ();
 sg13g2_fill_1 FILLER_63_35 ();
 sg13g2_fill_2 FILLER_63_48 ();
 sg13g2_fill_1 FILLER_63_50 ();
 sg13g2_fill_1 FILLER_63_57 ();
 sg13g2_fill_1 FILLER_63_67 ();
 sg13g2_decap_8 FILLER_63_73 ();
 sg13g2_fill_2 FILLER_63_85 ();
 sg13g2_fill_2 FILLER_63_96 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_decap_8 FILLER_63_123 ();
 sg13g2_decap_8 FILLER_63_130 ();
 sg13g2_fill_2 FILLER_63_137 ();
 sg13g2_decap_4 FILLER_63_143 ();
 sg13g2_fill_1 FILLER_63_151 ();
 sg13g2_fill_2 FILLER_63_164 ();
 sg13g2_fill_2 FILLER_63_190 ();
 sg13g2_decap_8 FILLER_63_200 ();
 sg13g2_decap_8 FILLER_63_207 ();
 sg13g2_fill_1 FILLER_63_225 ();
 sg13g2_fill_2 FILLER_63_236 ();
 sg13g2_decap_4 FILLER_63_249 ();
 sg13g2_decap_4 FILLER_63_258 ();
 sg13g2_fill_1 FILLER_63_262 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_310 ();
 sg13g2_decap_8 FILLER_63_321 ();
 sg13g2_decap_8 FILLER_63_328 ();
 sg13g2_fill_1 FILLER_63_335 ();
 sg13g2_fill_1 FILLER_63_344 ();
 sg13g2_decap_4 FILLER_63_350 ();
 sg13g2_fill_2 FILLER_63_354 ();
 sg13g2_fill_1 FILLER_63_384 ();
 sg13g2_fill_1 FILLER_63_398 ();
 sg13g2_decap_4 FILLER_63_403 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_2 FILLER_63_412 ();
 sg13g2_fill_1 FILLER_63_414 ();
 sg13g2_fill_2 FILLER_63_449 ();
 sg13g2_fill_1 FILLER_63_451 ();
 sg13g2_fill_2 FILLER_63_499 ();
 sg13g2_decap_8 FILLER_63_506 ();
 sg13g2_fill_1 FILLER_63_513 ();
 sg13g2_decap_8 FILLER_63_519 ();
 sg13g2_fill_1 FILLER_63_526 ();
 sg13g2_fill_1 FILLER_63_533 ();
 sg13g2_fill_1 FILLER_63_542 ();
 sg13g2_fill_2 FILLER_63_555 ();
 sg13g2_decap_4 FILLER_63_562 ();
 sg13g2_fill_1 FILLER_63_566 ();
 sg13g2_fill_1 FILLER_63_571 ();
 sg13g2_fill_2 FILLER_63_577 ();
 sg13g2_decap_4 FILLER_63_596 ();
 sg13g2_fill_1 FILLER_63_608 ();
 sg13g2_fill_1 FILLER_63_618 ();
 sg13g2_fill_2 FILLER_63_623 ();
 sg13g2_fill_1 FILLER_63_633 ();
 sg13g2_fill_1 FILLER_63_649 ();
 sg13g2_fill_1 FILLER_63_654 ();
 sg13g2_decap_4 FILLER_63_660 ();
 sg13g2_fill_2 FILLER_63_683 ();
 sg13g2_fill_2 FILLER_63_694 ();
 sg13g2_decap_8 FILLER_63_700 ();
 sg13g2_fill_1 FILLER_63_707 ();
 sg13g2_fill_2 FILLER_63_719 ();
 sg13g2_decap_8 FILLER_63_729 ();
 sg13g2_decap_8 FILLER_63_736 ();
 sg13g2_decap_4 FILLER_63_743 ();
 sg13g2_fill_2 FILLER_63_747 ();
 sg13g2_decap_4 FILLER_63_758 ();
 sg13g2_fill_2 FILLER_63_762 ();
 sg13g2_decap_8 FILLER_63_778 ();
 sg13g2_decap_4 FILLER_63_785 ();
 sg13g2_fill_1 FILLER_63_789 ();
 sg13g2_fill_1 FILLER_63_799 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_fill_2 FILLER_63_812 ();
 sg13g2_decap_4 FILLER_63_828 ();
 sg13g2_decap_8 FILLER_63_865 ();
 sg13g2_decap_8 FILLER_63_877 ();
 sg13g2_fill_2 FILLER_63_889 ();
 sg13g2_fill_2 FILLER_63_902 ();
 sg13g2_fill_1 FILLER_63_904 ();
 sg13g2_decap_8 FILLER_63_926 ();
 sg13g2_decap_8 FILLER_63_933 ();
 sg13g2_decap_4 FILLER_63_940 ();
 sg13g2_fill_2 FILLER_63_944 ();
 sg13g2_decap_8 FILLER_63_950 ();
 sg13g2_fill_2 FILLER_63_957 ();
 sg13g2_fill_2 FILLER_63_967 ();
 sg13g2_fill_1 FILLER_63_969 ();
 sg13g2_fill_1 FILLER_63_975 ();
 sg13g2_decap_8 FILLER_63_1015 ();
 sg13g2_decap_8 FILLER_63_1022 ();
 sg13g2_decap_8 FILLER_63_1029 ();
 sg13g2_fill_2 FILLER_63_1036 ();
 sg13g2_fill_2 FILLER_63_1046 ();
 sg13g2_fill_1 FILLER_63_1077 ();
 sg13g2_fill_2 FILLER_63_1092 ();
 sg13g2_fill_1 FILLER_63_1094 ();
 sg13g2_fill_1 FILLER_63_1104 ();
 sg13g2_fill_2 FILLER_63_1116 ();
 sg13g2_decap_4 FILLER_63_1129 ();
 sg13g2_decap_4 FILLER_63_1154 ();
 sg13g2_fill_1 FILLER_63_1158 ();
 sg13g2_fill_1 FILLER_63_1171 ();
 sg13g2_decap_8 FILLER_63_1197 ();
 sg13g2_fill_2 FILLER_63_1204 ();
 sg13g2_fill_1 FILLER_63_1212 ();
 sg13g2_fill_2 FILLER_63_1240 ();
 sg13g2_fill_1 FILLER_63_1242 ();
 sg13g2_fill_2 FILLER_63_1248 ();
 sg13g2_fill_1 FILLER_63_1250 ();
 sg13g2_fill_1 FILLER_63_1255 ();
 sg13g2_fill_1 FILLER_63_1262 ();
 sg13g2_fill_1 FILLER_63_1268 ();
 sg13g2_fill_2 FILLER_63_1274 ();
 sg13g2_decap_8 FILLER_63_1281 ();
 sg13g2_decap_4 FILLER_63_1288 ();
 sg13g2_fill_1 FILLER_63_1292 ();
 sg13g2_decap_4 FILLER_63_1299 ();
 sg13g2_fill_1 FILLER_63_1308 ();
 sg13g2_fill_1 FILLER_63_1314 ();
 sg13g2_decap_8 FILLER_63_1325 ();
 sg13g2_decap_8 FILLER_63_1339 ();
 sg13g2_decap_8 FILLER_63_1346 ();
 sg13g2_decap_8 FILLER_63_1362 ();
 sg13g2_decap_8 FILLER_63_1369 ();
 sg13g2_decap_4 FILLER_63_1376 ();
 sg13g2_fill_2 FILLER_63_1380 ();
 sg13g2_fill_1 FILLER_63_1408 ();
 sg13g2_fill_1 FILLER_63_1419 ();
 sg13g2_decap_4 FILLER_63_1424 ();
 sg13g2_fill_1 FILLER_63_1458 ();
 sg13g2_decap_4 FILLER_63_1477 ();
 sg13g2_fill_2 FILLER_63_1481 ();
 sg13g2_fill_1 FILLER_63_1512 ();
 sg13g2_fill_1 FILLER_63_1518 ();
 sg13g2_fill_1 FILLER_63_1541 ();
 sg13g2_decap_8 FILLER_63_1550 ();
 sg13g2_decap_8 FILLER_63_1557 ();
 sg13g2_decap_8 FILLER_63_1564 ();
 sg13g2_fill_1 FILLER_63_1571 ();
 sg13g2_fill_2 FILLER_63_1585 ();
 sg13g2_fill_1 FILLER_63_1587 ();
 sg13g2_fill_2 FILLER_63_1601 ();
 sg13g2_fill_1 FILLER_63_1603 ();
 sg13g2_decap_8 FILLER_63_1628 ();
 sg13g2_fill_2 FILLER_63_1681 ();
 sg13g2_fill_2 FILLER_63_1687 ();
 sg13g2_fill_2 FILLER_63_1693 ();
 sg13g2_fill_1 FILLER_63_1695 ();
 sg13g2_fill_2 FILLER_63_1701 ();
 sg13g2_decap_8 FILLER_63_1708 ();
 sg13g2_decap_8 FILLER_63_1715 ();
 sg13g2_decap_8 FILLER_63_1722 ();
 sg13g2_decap_8 FILLER_63_1729 ();
 sg13g2_decap_8 FILLER_63_1736 ();
 sg13g2_decap_8 FILLER_63_1743 ();
 sg13g2_decap_8 FILLER_63_1750 ();
 sg13g2_decap_8 FILLER_63_1757 ();
 sg13g2_decap_8 FILLER_63_1764 ();
 sg13g2_fill_2 FILLER_63_1771 ();
 sg13g2_fill_1 FILLER_63_1773 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_4 FILLER_64_21 ();
 sg13g2_fill_2 FILLER_64_25 ();
 sg13g2_decap_8 FILLER_64_31 ();
 sg13g2_fill_1 FILLER_64_38 ();
 sg13g2_fill_2 FILLER_64_60 ();
 sg13g2_decap_4 FILLER_64_77 ();
 sg13g2_fill_2 FILLER_64_81 ();
 sg13g2_decap_8 FILLER_64_88 ();
 sg13g2_decap_4 FILLER_64_95 ();
 sg13g2_decap_4 FILLER_64_104 ();
 sg13g2_decap_8 FILLER_64_130 ();
 sg13g2_decap_8 FILLER_64_137 ();
 sg13g2_decap_8 FILLER_64_152 ();
 sg13g2_decap_8 FILLER_64_159 ();
 sg13g2_fill_1 FILLER_64_166 ();
 sg13g2_decap_8 FILLER_64_177 ();
 sg13g2_fill_2 FILLER_64_190 ();
 sg13g2_decap_8 FILLER_64_195 ();
 sg13g2_fill_1 FILLER_64_202 ();
 sg13g2_fill_2 FILLER_64_212 ();
 sg13g2_fill_1 FILLER_64_226 ();
 sg13g2_fill_2 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_237 ();
 sg13g2_fill_2 FILLER_64_242 ();
 sg13g2_fill_1 FILLER_64_249 ();
 sg13g2_decap_8 FILLER_64_255 ();
 sg13g2_decap_8 FILLER_64_262 ();
 sg13g2_decap_4 FILLER_64_269 ();
 sg13g2_decap_8 FILLER_64_278 ();
 sg13g2_decap_4 FILLER_64_285 ();
 sg13g2_fill_2 FILLER_64_289 ();
 sg13g2_fill_1 FILLER_64_307 ();
 sg13g2_decap_4 FILLER_64_326 ();
 sg13g2_fill_2 FILLER_64_330 ();
 sg13g2_fill_2 FILLER_64_346 ();
 sg13g2_decap_8 FILLER_64_353 ();
 sg13g2_decap_4 FILLER_64_365 ();
 sg13g2_fill_2 FILLER_64_374 ();
 sg13g2_fill_2 FILLER_64_379 ();
 sg13g2_fill_1 FILLER_64_388 ();
 sg13g2_decap_4 FILLER_64_419 ();
 sg13g2_fill_1 FILLER_64_423 ();
 sg13g2_decap_8 FILLER_64_433 ();
 sg13g2_decap_8 FILLER_64_440 ();
 sg13g2_decap_8 FILLER_64_447 ();
 sg13g2_decap_4 FILLER_64_454 ();
 sg13g2_decap_8 FILLER_64_462 ();
 sg13g2_decap_4 FILLER_64_469 ();
 sg13g2_decap_8 FILLER_64_477 ();
 sg13g2_decap_4 FILLER_64_484 ();
 sg13g2_fill_2 FILLER_64_496 ();
 sg13g2_decap_8 FILLER_64_503 ();
 sg13g2_decap_8 FILLER_64_519 ();
 sg13g2_decap_8 FILLER_64_526 ();
 sg13g2_fill_2 FILLER_64_533 ();
 sg13g2_fill_1 FILLER_64_543 ();
 sg13g2_fill_2 FILLER_64_549 ();
 sg13g2_decap_4 FILLER_64_561 ();
 sg13g2_fill_1 FILLER_64_565 ();
 sg13g2_decap_4 FILLER_64_570 ();
 sg13g2_fill_2 FILLER_64_574 ();
 sg13g2_fill_2 FILLER_64_581 ();
 sg13g2_fill_1 FILLER_64_583 ();
 sg13g2_decap_8 FILLER_64_651 ();
 sg13g2_decap_8 FILLER_64_663 ();
 sg13g2_decap_8 FILLER_64_670 ();
 sg13g2_fill_2 FILLER_64_677 ();
 sg13g2_fill_2 FILLER_64_684 ();
 sg13g2_decap_8 FILLER_64_701 ();
 sg13g2_fill_1 FILLER_64_708 ();
 sg13g2_fill_1 FILLER_64_725 ();
 sg13g2_fill_2 FILLER_64_743 ();
 sg13g2_fill_1 FILLER_64_745 ();
 sg13g2_fill_1 FILLER_64_756 ();
 sg13g2_fill_1 FILLER_64_762 ();
 sg13g2_fill_1 FILLER_64_772 ();
 sg13g2_decap_4 FILLER_64_827 ();
 sg13g2_fill_1 FILLER_64_831 ();
 sg13g2_fill_2 FILLER_64_846 ();
 sg13g2_fill_1 FILLER_64_848 ();
 sg13g2_decap_4 FILLER_64_854 ();
 sg13g2_decap_8 FILLER_64_863 ();
 sg13g2_decap_8 FILLER_64_870 ();
 sg13g2_fill_1 FILLER_64_877 ();
 sg13g2_fill_2 FILLER_64_890 ();
 sg13g2_decap_8 FILLER_64_925 ();
 sg13g2_decap_4 FILLER_64_932 ();
 sg13g2_fill_2 FILLER_64_936 ();
 sg13g2_decap_4 FILLER_64_956 ();
 sg13g2_fill_2 FILLER_64_960 ();
 sg13g2_fill_1 FILLER_64_970 ();
 sg13g2_fill_2 FILLER_64_975 ();
 sg13g2_fill_1 FILLER_64_977 ();
 sg13g2_fill_1 FILLER_64_994 ();
 sg13g2_fill_2 FILLER_64_999 ();
 sg13g2_fill_1 FILLER_64_1001 ();
 sg13g2_fill_2 FILLER_64_1006 ();
 sg13g2_fill_1 FILLER_64_1008 ();
 sg13g2_decap_8 FILLER_64_1017 ();
 sg13g2_decap_8 FILLER_64_1024 ();
 sg13g2_fill_2 FILLER_64_1035 ();
 sg13g2_fill_1 FILLER_64_1037 ();
 sg13g2_fill_2 FILLER_64_1070 ();
 sg13g2_decap_8 FILLER_64_1076 ();
 sg13g2_decap_4 FILLER_64_1083 ();
 sg13g2_fill_1 FILLER_64_1087 ();
 sg13g2_decap_8 FILLER_64_1111 ();
 sg13g2_decap_8 FILLER_64_1118 ();
 sg13g2_decap_4 FILLER_64_1125 ();
 sg13g2_fill_2 FILLER_64_1129 ();
 sg13g2_decap_8 FILLER_64_1134 ();
 sg13g2_decap_8 FILLER_64_1141 ();
 sg13g2_decap_8 FILLER_64_1148 ();
 sg13g2_decap_8 FILLER_64_1155 ();
 sg13g2_fill_2 FILLER_64_1162 ();
 sg13g2_decap_4 FILLER_64_1169 ();
 sg13g2_fill_1 FILLER_64_1173 ();
 sg13g2_fill_1 FILLER_64_1187 ();
 sg13g2_fill_2 FILLER_64_1193 ();
 sg13g2_fill_1 FILLER_64_1200 ();
 sg13g2_decap_8 FILLER_64_1206 ();
 sg13g2_decap_8 FILLER_64_1213 ();
 sg13g2_decap_8 FILLER_64_1220 ();
 sg13g2_decap_8 FILLER_64_1227 ();
 sg13g2_decap_4 FILLER_64_1234 ();
 sg13g2_decap_8 FILLER_64_1247 ();
 sg13g2_fill_2 FILLER_64_1254 ();
 sg13g2_fill_2 FILLER_64_1264 ();
 sg13g2_fill_1 FILLER_64_1266 ();
 sg13g2_decap_8 FILLER_64_1279 ();
 sg13g2_fill_2 FILLER_64_1286 ();
 sg13g2_fill_1 FILLER_64_1288 ();
 sg13g2_fill_1 FILLER_64_1294 ();
 sg13g2_decap_4 FILLER_64_1325 ();
 sg13g2_decap_8 FILLER_64_1339 ();
 sg13g2_decap_8 FILLER_64_1346 ();
 sg13g2_fill_1 FILLER_64_1353 ();
 sg13g2_fill_1 FILLER_64_1374 ();
 sg13g2_fill_2 FILLER_64_1380 ();
 sg13g2_decap_8 FILLER_64_1418 ();
 sg13g2_decap_8 FILLER_64_1439 ();
 sg13g2_fill_1 FILLER_64_1460 ();
 sg13g2_decap_8 FILLER_64_1472 ();
 sg13g2_fill_1 FILLER_64_1479 ();
 sg13g2_fill_2 FILLER_64_1499 ();
 sg13g2_fill_1 FILLER_64_1501 ();
 sg13g2_decap_8 FILLER_64_1507 ();
 sg13g2_decap_4 FILLER_64_1514 ();
 sg13g2_decap_4 FILLER_64_1526 ();
 sg13g2_fill_1 FILLER_64_1530 ();
 sg13g2_decap_4 FILLER_64_1539 ();
 sg13g2_fill_1 FILLER_64_1543 ();
 sg13g2_decap_4 FILLER_64_1552 ();
 sg13g2_decap_8 FILLER_64_1569 ();
 sg13g2_fill_2 FILLER_64_1576 ();
 sg13g2_decap_4 FILLER_64_1582 ();
 sg13g2_fill_1 FILLER_64_1586 ();
 sg13g2_fill_1 FILLER_64_1595 ();
 sg13g2_decap_8 FILLER_64_1613 ();
 sg13g2_fill_2 FILLER_64_1620 ();
 sg13g2_fill_2 FILLER_64_1626 ();
 sg13g2_fill_1 FILLER_64_1642 ();
 sg13g2_fill_2 FILLER_64_1669 ();
 sg13g2_decap_4 FILLER_64_1697 ();
 sg13g2_fill_1 FILLER_64_1701 ();
 sg13g2_decap_8 FILLER_64_1719 ();
 sg13g2_decap_8 FILLER_64_1726 ();
 sg13g2_decap_8 FILLER_64_1733 ();
 sg13g2_decap_8 FILLER_64_1740 ();
 sg13g2_decap_8 FILLER_64_1747 ();
 sg13g2_decap_8 FILLER_64_1754 ();
 sg13g2_decap_8 FILLER_64_1761 ();
 sg13g2_decap_4 FILLER_64_1768 ();
 sg13g2_fill_2 FILLER_64_1772 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_4 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_18 ();
 sg13g2_decap_4 FILLER_65_46 ();
 sg13g2_fill_1 FILLER_65_54 ();
 sg13g2_fill_2 FILLER_65_65 ();
 sg13g2_fill_1 FILLER_65_72 ();
 sg13g2_decap_4 FILLER_65_79 ();
 sg13g2_fill_2 FILLER_65_83 ();
 sg13g2_fill_1 FILLER_65_90 ();
 sg13g2_decap_4 FILLER_65_103 ();
 sg13g2_fill_2 FILLER_65_112 ();
 sg13g2_fill_1 FILLER_65_114 ();
 sg13g2_decap_4 FILLER_65_123 ();
 sg13g2_fill_2 FILLER_65_127 ();
 sg13g2_fill_1 FILLER_65_139 ();
 sg13g2_fill_1 FILLER_65_146 ();
 sg13g2_fill_2 FILLER_65_152 ();
 sg13g2_fill_1 FILLER_65_193 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_fill_1 FILLER_65_247 ();
 sg13g2_fill_2 FILLER_65_252 ();
 sg13g2_fill_1 FILLER_65_254 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_4 FILLER_65_280 ();
 sg13g2_decap_4 FILLER_65_290 ();
 sg13g2_fill_1 FILLER_65_294 ();
 sg13g2_decap_4 FILLER_65_308 ();
 sg13g2_fill_2 FILLER_65_312 ();
 sg13g2_decap_4 FILLER_65_326 ();
 sg13g2_fill_1 FILLER_65_330 ();
 sg13g2_fill_1 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_370 ();
 sg13g2_decap_8 FILLER_65_377 ();
 sg13g2_fill_1 FILLER_65_384 ();
 sg13g2_decap_4 FILLER_65_393 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_fill_2 FILLER_65_449 ();
 sg13g2_fill_2 FILLER_65_456 ();
 sg13g2_fill_1 FILLER_65_458 ();
 sg13g2_fill_1 FILLER_65_464 ();
 sg13g2_fill_2 FILLER_65_470 ();
 sg13g2_fill_1 FILLER_65_472 ();
 sg13g2_fill_1 FILLER_65_480 ();
 sg13g2_fill_2 FILLER_65_511 ();
 sg13g2_fill_2 FILLER_65_520 ();
 sg13g2_fill_1 FILLER_65_550 ();
 sg13g2_fill_2 FILLER_65_560 ();
 sg13g2_fill_1 FILLER_65_562 ();
 sg13g2_fill_1 FILLER_65_567 ();
 sg13g2_fill_2 FILLER_65_573 ();
 sg13g2_fill_1 FILLER_65_575 ();
 sg13g2_fill_2 FILLER_65_598 ();
 sg13g2_fill_2 FILLER_65_625 ();
 sg13g2_decap_8 FILLER_65_641 ();
 sg13g2_fill_1 FILLER_65_680 ();
 sg13g2_decap_8 FILLER_65_694 ();
 sg13g2_decap_8 FILLER_65_701 ();
 sg13g2_decap_4 FILLER_65_708 ();
 sg13g2_decap_4 FILLER_65_718 ();
 sg13g2_fill_2 FILLER_65_725 ();
 sg13g2_fill_2 FILLER_65_745 ();
 sg13g2_fill_1 FILLER_65_747 ();
 sg13g2_fill_2 FILLER_65_768 ();
 sg13g2_fill_1 FILLER_65_795 ();
 sg13g2_fill_2 FILLER_65_801 ();
 sg13g2_decap_8 FILLER_65_808 ();
 sg13g2_fill_2 FILLER_65_815 ();
 sg13g2_decap_4 FILLER_65_821 ();
 sg13g2_fill_2 FILLER_65_829 ();
 sg13g2_fill_1 FILLER_65_831 ();
 sg13g2_fill_2 FILLER_65_840 ();
 sg13g2_fill_2 FILLER_65_846 ();
 sg13g2_fill_1 FILLER_65_848 ();
 sg13g2_fill_1 FILLER_65_864 ();
 sg13g2_fill_1 FILLER_65_870 ();
 sg13g2_fill_1 FILLER_65_886 ();
 sg13g2_fill_2 FILLER_65_899 ();
 sg13g2_fill_1 FILLER_65_901 ();
 sg13g2_fill_2 FILLER_65_907 ();
 sg13g2_fill_1 FILLER_65_914 ();
 sg13g2_fill_1 FILLER_65_935 ();
 sg13g2_fill_2 FILLER_65_942 ();
 sg13g2_fill_1 FILLER_65_944 ();
 sg13g2_fill_2 FILLER_65_974 ();
 sg13g2_fill_1 FILLER_65_976 ();
 sg13g2_fill_1 FILLER_65_986 ();
 sg13g2_decap_8 FILLER_65_1017 ();
 sg13g2_fill_2 FILLER_65_1024 ();
 sg13g2_fill_2 FILLER_65_1031 ();
 sg13g2_decap_4 FILLER_65_1073 ();
 sg13g2_decap_4 FILLER_65_1081 ();
 sg13g2_decap_8 FILLER_65_1102 ();
 sg13g2_decap_8 FILLER_65_1109 ();
 sg13g2_fill_1 FILLER_65_1116 ();
 sg13g2_decap_8 FILLER_65_1159 ();
 sg13g2_fill_1 FILLER_65_1171 ();
 sg13g2_fill_1 FILLER_65_1181 ();
 sg13g2_fill_2 FILLER_65_1223 ();
 sg13g2_fill_1 FILLER_65_1225 ();
 sg13g2_fill_2 FILLER_65_1230 ();
 sg13g2_fill_1 FILLER_65_1232 ();
 sg13g2_decap_4 FILLER_65_1250 ();
 sg13g2_fill_1 FILLER_65_1254 ();
 sg13g2_fill_2 FILLER_65_1263 ();
 sg13g2_fill_1 FILLER_65_1274 ();
 sg13g2_decap_8 FILLER_65_1288 ();
 sg13g2_decap_8 FILLER_65_1295 ();
 sg13g2_fill_1 FILLER_65_1302 ();
 sg13g2_decap_8 FILLER_65_1318 ();
 sg13g2_decap_4 FILLER_65_1325 ();
 sg13g2_fill_1 FILLER_65_1329 ();
 sg13g2_fill_2 FILLER_65_1340 ();
 sg13g2_fill_1 FILLER_65_1342 ();
 sg13g2_decap_8 FILLER_65_1352 ();
 sg13g2_fill_1 FILLER_65_1368 ();
 sg13g2_fill_1 FILLER_65_1374 ();
 sg13g2_fill_1 FILLER_65_1379 ();
 sg13g2_fill_1 FILLER_65_1396 ();
 sg13g2_fill_2 FILLER_65_1419 ();
 sg13g2_decap_8 FILLER_65_1425 ();
 sg13g2_fill_1 FILLER_65_1432 ();
 sg13g2_decap_8 FILLER_65_1441 ();
 sg13g2_decap_8 FILLER_65_1454 ();
 sg13g2_fill_1 FILLER_65_1461 ();
 sg13g2_fill_1 FILLER_65_1470 ();
 sg13g2_decap_4 FILLER_65_1476 ();
 sg13g2_fill_2 FILLER_65_1485 ();
 sg13g2_fill_1 FILLER_65_1495 ();
 sg13g2_decap_8 FILLER_65_1504 ();
 sg13g2_decap_8 FILLER_65_1511 ();
 sg13g2_decap_8 FILLER_65_1518 ();
 sg13g2_fill_1 FILLER_65_1541 ();
 sg13g2_fill_2 FILLER_65_1554 ();
 sg13g2_fill_1 FILLER_65_1556 ();
 sg13g2_decap_8 FILLER_65_1561 ();
 sg13g2_decap_8 FILLER_65_1568 ();
 sg13g2_decap_8 FILLER_65_1575 ();
 sg13g2_fill_1 FILLER_65_1592 ();
 sg13g2_fill_1 FILLER_65_1598 ();
 sg13g2_fill_1 FILLER_65_1605 ();
 sg13g2_fill_1 FILLER_65_1612 ();
 sg13g2_fill_1 FILLER_65_1617 ();
 sg13g2_fill_1 FILLER_65_1623 ();
 sg13g2_fill_1 FILLER_65_1629 ();
 sg13g2_fill_2 FILLER_65_1649 ();
 sg13g2_fill_1 FILLER_65_1689 ();
 sg13g2_decap_4 FILLER_65_1694 ();
 sg13g2_decap_8 FILLER_65_1715 ();
 sg13g2_decap_8 FILLER_65_1722 ();
 sg13g2_decap_8 FILLER_65_1729 ();
 sg13g2_decap_8 FILLER_65_1736 ();
 sg13g2_decap_8 FILLER_65_1743 ();
 sg13g2_decap_8 FILLER_65_1750 ();
 sg13g2_decap_8 FILLER_65_1757 ();
 sg13g2_decap_8 FILLER_65_1764 ();
 sg13g2_fill_2 FILLER_65_1771 ();
 sg13g2_fill_1 FILLER_65_1773 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_35 ();
 sg13g2_fill_2 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_44 ();
 sg13g2_fill_2 FILLER_66_50 ();
 sg13g2_fill_1 FILLER_66_52 ();
 sg13g2_fill_2 FILLER_66_101 ();
 sg13g2_fill_1 FILLER_66_103 ();
 sg13g2_fill_1 FILLER_66_112 ();
 sg13g2_decap_4 FILLER_66_118 ();
 sg13g2_fill_1 FILLER_66_122 ();
 sg13g2_fill_2 FILLER_66_140 ();
 sg13g2_fill_2 FILLER_66_157 ();
 sg13g2_fill_1 FILLER_66_164 ();
 sg13g2_fill_1 FILLER_66_176 ();
 sg13g2_fill_1 FILLER_66_202 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_fill_2 FILLER_66_231 ();
 sg13g2_fill_1 FILLER_66_233 ();
 sg13g2_fill_2 FILLER_66_256 ();
 sg13g2_fill_1 FILLER_66_258 ();
 sg13g2_fill_2 FILLER_66_278 ();
 sg13g2_fill_1 FILLER_66_280 ();
 sg13g2_fill_1 FILLER_66_285 ();
 sg13g2_fill_1 FILLER_66_291 ();
 sg13g2_fill_1 FILLER_66_303 ();
 sg13g2_fill_1 FILLER_66_329 ();
 sg13g2_decap_8 FILLER_66_351 ();
 sg13g2_decap_8 FILLER_66_358 ();
 sg13g2_decap_8 FILLER_66_365 ();
 sg13g2_decap_8 FILLER_66_372 ();
 sg13g2_fill_2 FILLER_66_379 ();
 sg13g2_fill_2 FILLER_66_397 ();
 sg13g2_fill_1 FILLER_66_399 ();
 sg13g2_decap_8 FILLER_66_419 ();
 sg13g2_decap_8 FILLER_66_426 ();
 sg13g2_fill_2 FILLER_66_433 ();
 sg13g2_fill_1 FILLER_66_435 ();
 sg13g2_fill_1 FILLER_66_468 ();
 sg13g2_fill_2 FILLER_66_474 ();
 sg13g2_fill_2 FILLER_66_490 ();
 sg13g2_decap_8 FILLER_66_533 ();
 sg13g2_decap_4 FILLER_66_540 ();
 sg13g2_decap_4 FILLER_66_554 ();
 sg13g2_fill_2 FILLER_66_580 ();
 sg13g2_decap_8 FILLER_66_600 ();
 sg13g2_decap_4 FILLER_66_607 ();
 sg13g2_fill_1 FILLER_66_616 ();
 sg13g2_fill_2 FILLER_66_639 ();
 sg13g2_fill_2 FILLER_66_648 ();
 sg13g2_fill_2 FILLER_66_671 ();
 sg13g2_fill_1 FILLER_66_673 ();
 sg13g2_fill_1 FILLER_66_688 ();
 sg13g2_fill_1 FILLER_66_695 ();
 sg13g2_fill_2 FILLER_66_704 ();
 sg13g2_decap_8 FILLER_66_714 ();
 sg13g2_decap_8 FILLER_66_725 ();
 sg13g2_decap_4 FILLER_66_732 ();
 sg13g2_fill_1 FILLER_66_736 ();
 sg13g2_fill_2 FILLER_66_754 ();
 sg13g2_fill_1 FILLER_66_756 ();
 sg13g2_fill_2 FILLER_66_806 ();
 sg13g2_decap_4 FILLER_66_812 ();
 sg13g2_fill_1 FILLER_66_816 ();
 sg13g2_decap_4 FILLER_66_826 ();
 sg13g2_fill_2 FILLER_66_830 ();
 sg13g2_decap_8 FILLER_66_837 ();
 sg13g2_fill_1 FILLER_66_844 ();
 sg13g2_fill_2 FILLER_66_868 ();
 sg13g2_fill_1 FILLER_66_870 ();
 sg13g2_fill_2 FILLER_66_879 ();
 sg13g2_fill_2 FILLER_66_889 ();
 sg13g2_fill_1 FILLER_66_891 ();
 sg13g2_decap_4 FILLER_66_909 ();
 sg13g2_decap_8 FILLER_66_921 ();
 sg13g2_fill_2 FILLER_66_928 ();
 sg13g2_fill_1 FILLER_66_930 ();
 sg13g2_fill_2 FILLER_66_943 ();
 sg13g2_fill_2 FILLER_66_970 ();
 sg13g2_fill_1 FILLER_66_972 ();
 sg13g2_fill_2 FILLER_66_978 ();
 sg13g2_fill_1 FILLER_66_980 ();
 sg13g2_fill_2 FILLER_66_989 ();
 sg13g2_decap_8 FILLER_66_1000 ();
 sg13g2_fill_2 FILLER_66_1007 ();
 sg13g2_fill_1 FILLER_66_1009 ();
 sg13g2_decap_4 FILLER_66_1023 ();
 sg13g2_fill_2 FILLER_66_1037 ();
 sg13g2_fill_1 FILLER_66_1039 ();
 sg13g2_decap_8 FILLER_66_1048 ();
 sg13g2_decap_4 FILLER_66_1055 ();
 sg13g2_fill_2 FILLER_66_1059 ();
 sg13g2_decap_4 FILLER_66_1065 ();
 sg13g2_fill_2 FILLER_66_1079 ();
 sg13g2_fill_1 FILLER_66_1081 ();
 sg13g2_decap_8 FILLER_66_1096 ();
 sg13g2_decap_8 FILLER_66_1112 ();
 sg13g2_decap_4 FILLER_66_1119 ();
 sg13g2_decap_8 FILLER_66_1126 ();
 sg13g2_fill_1 FILLER_66_1133 ();
 sg13g2_decap_8 FILLER_66_1138 ();
 sg13g2_fill_1 FILLER_66_1145 ();
 sg13g2_fill_1 FILLER_66_1151 ();
 sg13g2_fill_2 FILLER_66_1156 ();
 sg13g2_decap_4 FILLER_66_1189 ();
 sg13g2_fill_2 FILLER_66_1193 ();
 sg13g2_decap_8 FILLER_66_1205 ();
 sg13g2_decap_4 FILLER_66_1212 ();
 sg13g2_decap_4 FILLER_66_1224 ();
 sg13g2_fill_2 FILLER_66_1237 ();
 sg13g2_decap_4 FILLER_66_1244 ();
 sg13g2_fill_1 FILLER_66_1270 ();
 sg13g2_fill_2 FILLER_66_1275 ();
 sg13g2_decap_8 FILLER_66_1287 ();
 sg13g2_decap_8 FILLER_66_1294 ();
 sg13g2_decap_8 FILLER_66_1315 ();
 sg13g2_decap_4 FILLER_66_1322 ();
 sg13g2_fill_2 FILLER_66_1326 ();
 sg13g2_fill_2 FILLER_66_1337 ();
 sg13g2_fill_1 FILLER_66_1339 ();
 sg13g2_decap_8 FILLER_66_1355 ();
 sg13g2_decap_4 FILLER_66_1367 ();
 sg13g2_fill_1 FILLER_66_1371 ();
 sg13g2_fill_1 FILLER_66_1380 ();
 sg13g2_fill_1 FILLER_66_1391 ();
 sg13g2_decap_8 FILLER_66_1401 ();
 sg13g2_decap_8 FILLER_66_1408 ();
 sg13g2_decap_8 FILLER_66_1415 ();
 sg13g2_decap_8 FILLER_66_1422 ();
 sg13g2_fill_2 FILLER_66_1429 ();
 sg13g2_decap_8 FILLER_66_1437 ();
 sg13g2_decap_8 FILLER_66_1444 ();
 sg13g2_decap_4 FILLER_66_1451 ();
 sg13g2_fill_2 FILLER_66_1468 ();
 sg13g2_fill_1 FILLER_66_1470 ();
 sg13g2_decap_4 FILLER_66_1481 ();
 sg13g2_fill_2 FILLER_66_1485 ();
 sg13g2_decap_4 FILLER_66_1492 ();
 sg13g2_fill_2 FILLER_66_1496 ();
 sg13g2_fill_1 FILLER_66_1510 ();
 sg13g2_decap_4 FILLER_66_1519 ();
 sg13g2_fill_1 FILLER_66_1523 ();
 sg13g2_fill_2 FILLER_66_1532 ();
 sg13g2_fill_1 FILLER_66_1534 ();
 sg13g2_fill_2 FILLER_66_1540 ();
 sg13g2_fill_2 FILLER_66_1548 ();
 sg13g2_fill_1 FILLER_66_1575 ();
 sg13g2_fill_2 FILLER_66_1586 ();
 sg13g2_fill_1 FILLER_66_1588 ();
 sg13g2_fill_2 FILLER_66_1598 ();
 sg13g2_fill_2 FILLER_66_1610 ();
 sg13g2_fill_1 FILLER_66_1612 ();
 sg13g2_decap_4 FILLER_66_1620 ();
 sg13g2_fill_1 FILLER_66_1657 ();
 sg13g2_fill_1 FILLER_66_1668 ();
 sg13g2_decap_8 FILLER_66_1690 ();
 sg13g2_decap_8 FILLER_66_1697 ();
 sg13g2_decap_8 FILLER_66_1704 ();
 sg13g2_decap_8 FILLER_66_1711 ();
 sg13g2_decap_8 FILLER_66_1718 ();
 sg13g2_fill_2 FILLER_66_1725 ();
 sg13g2_fill_1 FILLER_66_1727 ();
 sg13g2_decap_8 FILLER_66_1732 ();
 sg13g2_decap_8 FILLER_66_1739 ();
 sg13g2_decap_8 FILLER_66_1746 ();
 sg13g2_decap_8 FILLER_66_1753 ();
 sg13g2_decap_8 FILLER_66_1760 ();
 sg13g2_decap_8 FILLER_66_1767 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_4 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_fill_1 FILLER_67_109 ();
 sg13g2_fill_1 FILLER_67_115 ();
 sg13g2_fill_2 FILLER_67_133 ();
 sg13g2_fill_2 FILLER_67_145 ();
 sg13g2_fill_1 FILLER_67_162 ();
 sg13g2_fill_2 FILLER_67_172 ();
 sg13g2_fill_2 FILLER_67_193 ();
 sg13g2_fill_2 FILLER_67_224 ();
 sg13g2_fill_2 FILLER_67_231 ();
 sg13g2_fill_2 FILLER_67_243 ();
 sg13g2_decap_4 FILLER_67_263 ();
 sg13g2_decap_4 FILLER_67_280 ();
 sg13g2_fill_1 FILLER_67_284 ();
 sg13g2_fill_2 FILLER_67_297 ();
 sg13g2_fill_1 FILLER_67_310 ();
 sg13g2_fill_1 FILLER_67_330 ();
 sg13g2_fill_1 FILLER_67_341 ();
 sg13g2_decap_4 FILLER_67_347 ();
 sg13g2_decap_8 FILLER_67_416 ();
 sg13g2_fill_2 FILLER_67_423 ();
 sg13g2_fill_2 FILLER_67_442 ();
 sg13g2_fill_1 FILLER_67_449 ();
 sg13g2_fill_2 FILLER_67_455 ();
 sg13g2_decap_4 FILLER_67_461 ();
 sg13g2_fill_2 FILLER_67_465 ();
 sg13g2_decap_4 FILLER_67_472 ();
 sg13g2_fill_1 FILLER_67_495 ();
 sg13g2_fill_1 FILLER_67_509 ();
 sg13g2_fill_2 FILLER_67_515 ();
 sg13g2_fill_2 FILLER_67_525 ();
 sg13g2_fill_2 FILLER_67_535 ();
 sg13g2_fill_1 FILLER_67_565 ();
 sg13g2_decap_8 FILLER_67_570 ();
 sg13g2_decap_4 FILLER_67_577 ();
 sg13g2_fill_1 FILLER_67_585 ();
 sg13g2_fill_2 FILLER_67_616 ();
 sg13g2_fill_1 FILLER_67_618 ();
 sg13g2_decap_8 FILLER_67_627 ();
 sg13g2_fill_2 FILLER_67_634 ();
 sg13g2_fill_2 FILLER_67_641 ();
 sg13g2_fill_2 FILLER_67_652 ();
 sg13g2_decap_4 FILLER_67_659 ();
 sg13g2_fill_2 FILLER_67_663 ();
 sg13g2_fill_1 FILLER_67_670 ();
 sg13g2_decap_8 FILLER_67_675 ();
 sg13g2_decap_4 FILLER_67_682 ();
 sg13g2_fill_2 FILLER_67_686 ();
 sg13g2_fill_1 FILLER_67_691 ();
 sg13g2_decap_4 FILLER_67_722 ();
 sg13g2_decap_4 FILLER_67_730 ();
 sg13g2_fill_2 FILLER_67_734 ();
 sg13g2_fill_2 FILLER_67_787 ();
 sg13g2_decap_8 FILLER_67_832 ();
 sg13g2_fill_2 FILLER_67_839 ();
 sg13g2_fill_1 FILLER_67_841 ();
 sg13g2_fill_2 FILLER_67_850 ();
 sg13g2_fill_1 FILLER_67_852 ();
 sg13g2_decap_8 FILLER_67_871 ();
 sg13g2_fill_1 FILLER_67_882 ();
 sg13g2_decap_8 FILLER_67_906 ();
 sg13g2_fill_2 FILLER_67_913 ();
 sg13g2_fill_1 FILLER_67_915 ();
 sg13g2_decap_4 FILLER_67_924 ();
 sg13g2_fill_1 FILLER_67_928 ();
 sg13g2_fill_1 FILLER_67_934 ();
 sg13g2_fill_2 FILLER_67_945 ();
 sg13g2_fill_1 FILLER_67_947 ();
 sg13g2_fill_1 FILLER_67_961 ();
 sg13g2_decap_8 FILLER_67_979 ();
 sg13g2_decap_4 FILLER_67_986 ();
 sg13g2_fill_2 FILLER_67_990 ();
 sg13g2_fill_1 FILLER_67_999 ();
 sg13g2_decap_8 FILLER_67_1005 ();
 sg13g2_decap_8 FILLER_67_1012 ();
 sg13g2_decap_4 FILLER_67_1019 ();
 sg13g2_fill_1 FILLER_67_1027 ();
 sg13g2_decap_8 FILLER_67_1068 ();
 sg13g2_decap_8 FILLER_67_1075 ();
 sg13g2_decap_8 FILLER_67_1082 ();
 sg13g2_fill_2 FILLER_67_1089 ();
 sg13g2_fill_1 FILLER_67_1091 ();
 sg13g2_decap_8 FILLER_67_1101 ();
 sg13g2_decap_8 FILLER_67_1117 ();
 sg13g2_fill_2 FILLER_67_1124 ();
 sg13g2_fill_1 FILLER_67_1126 ();
 sg13g2_fill_2 FILLER_67_1141 ();
 sg13g2_fill_2 FILLER_67_1155 ();
 sg13g2_fill_2 FILLER_67_1165 ();
 sg13g2_fill_1 FILLER_67_1183 ();
 sg13g2_decap_4 FILLER_67_1190 ();
 sg13g2_decap_8 FILLER_67_1202 ();
 sg13g2_decap_8 FILLER_67_1209 ();
 sg13g2_decap_8 FILLER_67_1216 ();
 sg13g2_decap_4 FILLER_67_1223 ();
 sg13g2_fill_1 FILLER_67_1227 ();
 sg13g2_fill_2 FILLER_67_1242 ();
 sg13g2_fill_1 FILLER_67_1257 ();
 sg13g2_decap_8 FILLER_67_1292 ();
 sg13g2_decap_8 FILLER_67_1299 ();
 sg13g2_decap_8 FILLER_67_1306 ();
 sg13g2_fill_2 FILLER_67_1313 ();
 sg13g2_decap_8 FILLER_67_1319 ();
 sg13g2_decap_8 FILLER_67_1326 ();
 sg13g2_fill_1 FILLER_67_1333 ();
 sg13g2_fill_1 FILLER_67_1339 ();
 sg13g2_fill_1 FILLER_67_1348 ();
 sg13g2_fill_1 FILLER_67_1384 ();
 sg13g2_fill_1 FILLER_67_1400 ();
 sg13g2_fill_2 FILLER_67_1415 ();
 sg13g2_fill_1 FILLER_67_1417 ();
 sg13g2_fill_2 FILLER_67_1426 ();
 sg13g2_fill_2 FILLER_67_1447 ();
 sg13g2_fill_1 FILLER_67_1449 ();
 sg13g2_decap_4 FILLER_67_1469 ();
 sg13g2_fill_1 FILLER_67_1473 ();
 sg13g2_decap_8 FILLER_67_1488 ();
 sg13g2_decap_8 FILLER_67_1495 ();
 sg13g2_decap_8 FILLER_67_1502 ();
 sg13g2_decap_8 FILLER_67_1509 ();
 sg13g2_decap_8 FILLER_67_1516 ();
 sg13g2_fill_2 FILLER_67_1523 ();
 sg13g2_decap_4 FILLER_67_1551 ();
 sg13g2_fill_1 FILLER_67_1573 ();
 sg13g2_decap_8 FILLER_67_1579 ();
 sg13g2_decap_4 FILLER_67_1586 ();
 sg13g2_fill_1 FILLER_67_1605 ();
 sg13g2_fill_1 FILLER_67_1625 ();
 sg13g2_fill_2 FILLER_67_1634 ();
 sg13g2_fill_1 FILLER_67_1644 ();
 sg13g2_fill_1 FILLER_67_1656 ();
 sg13g2_fill_1 FILLER_67_1666 ();
 sg13g2_fill_2 FILLER_67_1671 ();
 sg13g2_fill_1 FILLER_67_1673 ();
 sg13g2_decap_8 FILLER_67_1677 ();
 sg13g2_decap_8 FILLER_67_1684 ();
 sg13g2_decap_8 FILLER_67_1695 ();
 sg13g2_decap_8 FILLER_67_1702 ();
 sg13g2_decap_8 FILLER_67_1709 ();
 sg13g2_decap_4 FILLER_67_1716 ();
 sg13g2_fill_1 FILLER_67_1720 ();
 sg13g2_decap_8 FILLER_67_1747 ();
 sg13g2_decap_8 FILLER_67_1754 ();
 sg13g2_decap_8 FILLER_67_1761 ();
 sg13g2_decap_4 FILLER_67_1768 ();
 sg13g2_fill_2 FILLER_67_1772 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_fill_2 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_37 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_fill_2 FILLER_68_63 ();
 sg13g2_fill_1 FILLER_68_65 ();
 sg13g2_decap_4 FILLER_68_70 ();
 sg13g2_fill_2 FILLER_68_74 ();
 sg13g2_decap_8 FILLER_68_80 ();
 sg13g2_fill_1 FILLER_68_87 ();
 sg13g2_fill_1 FILLER_68_108 ();
 sg13g2_fill_1 FILLER_68_117 ();
 sg13g2_fill_1 FILLER_68_152 ();
 sg13g2_fill_2 FILLER_68_157 ();
 sg13g2_fill_1 FILLER_68_165 ();
 sg13g2_fill_1 FILLER_68_173 ();
 sg13g2_fill_2 FILLER_68_178 ();
 sg13g2_fill_2 FILLER_68_188 ();
 sg13g2_fill_2 FILLER_68_201 ();
 sg13g2_decap_8 FILLER_68_246 ();
 sg13g2_decap_8 FILLER_68_253 ();
 sg13g2_decap_4 FILLER_68_260 ();
 sg13g2_fill_1 FILLER_68_264 ();
 sg13g2_decap_8 FILLER_68_278 ();
 sg13g2_fill_1 FILLER_68_285 ();
 sg13g2_fill_1 FILLER_68_299 ();
 sg13g2_fill_2 FILLER_68_315 ();
 sg13g2_fill_1 FILLER_68_343 ();
 sg13g2_fill_1 FILLER_68_374 ();
 sg13g2_fill_2 FILLER_68_387 ();
 sg13g2_decap_8 FILLER_68_408 ();
 sg13g2_decap_4 FILLER_68_415 ();
 sg13g2_fill_1 FILLER_68_419 ();
 sg13g2_decap_8 FILLER_68_429 ();
 sg13g2_decap_8 FILLER_68_436 ();
 sg13g2_fill_1 FILLER_68_446 ();
 sg13g2_decap_4 FILLER_68_467 ();
 sg13g2_fill_1 FILLER_68_471 ();
 sg13g2_decap_4 FILLER_68_479 ();
 sg13g2_fill_1 FILLER_68_510 ();
 sg13g2_decap_8 FILLER_68_522 ();
 sg13g2_fill_1 FILLER_68_547 ();
 sg13g2_fill_1 FILLER_68_559 ();
 sg13g2_fill_1 FILLER_68_590 ();
 sg13g2_decap_4 FILLER_68_599 ();
 sg13g2_fill_1 FILLER_68_603 ();
 sg13g2_fill_1 FILLER_68_616 ();
 sg13g2_fill_2 FILLER_68_648 ();
 sg13g2_fill_2 FILLER_68_658 ();
 sg13g2_fill_2 FILLER_68_673 ();
 sg13g2_fill_1 FILLER_68_683 ();
 sg13g2_fill_1 FILLER_68_693 ();
 sg13g2_fill_1 FILLER_68_699 ();
 sg13g2_decap_4 FILLER_68_704 ();
 sg13g2_fill_1 FILLER_68_708 ();
 sg13g2_fill_1 FILLER_68_729 ();
 sg13g2_fill_2 FILLER_68_737 ();
 sg13g2_fill_2 FILLER_68_817 ();
 sg13g2_fill_1 FILLER_68_819 ();
 sg13g2_fill_2 FILLER_68_828 ();
 sg13g2_decap_4 FILLER_68_839 ();
 sg13g2_decap_8 FILLER_68_847 ();
 sg13g2_decap_8 FILLER_68_854 ();
 sg13g2_decap_4 FILLER_68_861 ();
 sg13g2_decap_4 FILLER_68_877 ();
 sg13g2_fill_2 FILLER_68_881 ();
 sg13g2_decap_8 FILLER_68_905 ();
 sg13g2_decap_8 FILLER_68_912 ();
 sg13g2_fill_2 FILLER_68_919 ();
 sg13g2_decap_4 FILLER_68_938 ();
 sg13g2_fill_2 FILLER_68_942 ();
 sg13g2_decap_8 FILLER_68_962 ();
 sg13g2_decap_8 FILLER_68_977 ();
 sg13g2_fill_2 FILLER_68_984 ();
 sg13g2_decap_4 FILLER_68_1012 ();
 sg13g2_fill_1 FILLER_68_1016 ();
 sg13g2_decap_4 FILLER_68_1029 ();
 sg13g2_decap_8 FILLER_68_1046 ();
 sg13g2_fill_2 FILLER_68_1053 ();
 sg13g2_fill_2 FILLER_68_1060 ();
 sg13g2_fill_1 FILLER_68_1067 ();
 sg13g2_decap_4 FILLER_68_1085 ();
 sg13g2_fill_1 FILLER_68_1089 ();
 sg13g2_decap_4 FILLER_68_1116 ();
 sg13g2_fill_2 FILLER_68_1120 ();
 sg13g2_fill_2 FILLER_68_1135 ();
 sg13g2_fill_1 FILLER_68_1137 ();
 sg13g2_decap_4 FILLER_68_1149 ();
 sg13g2_fill_1 FILLER_68_1157 ();
 sg13g2_fill_2 FILLER_68_1166 ();
 sg13g2_fill_2 FILLER_68_1183 ();
 sg13g2_fill_2 FILLER_68_1206 ();
 sg13g2_fill_1 FILLER_68_1208 ();
 sg13g2_decap_8 FILLER_68_1223 ();
 sg13g2_decap_8 FILLER_68_1230 ();
 sg13g2_fill_2 FILLER_68_1237 ();
 sg13g2_fill_1 FILLER_68_1239 ();
 sg13g2_fill_2 FILLER_68_1260 ();
 sg13g2_fill_1 FILLER_68_1262 ();
 sg13g2_fill_2 FILLER_68_1276 ();
 sg13g2_decap_8 FILLER_68_1286 ();
 sg13g2_decap_8 FILLER_68_1293 ();
 sg13g2_fill_1 FILLER_68_1300 ();
 sg13g2_decap_4 FILLER_68_1311 ();
 sg13g2_fill_2 FILLER_68_1315 ();
 sg13g2_fill_2 FILLER_68_1325 ();
 sg13g2_fill_2 FILLER_68_1344 ();
 sg13g2_decap_4 FILLER_68_1351 ();
 sg13g2_decap_4 FILLER_68_1373 ();
 sg13g2_fill_1 FILLER_68_1377 ();
 sg13g2_fill_2 FILLER_68_1396 ();
 sg13g2_fill_1 FILLER_68_1398 ();
 sg13g2_decap_8 FILLER_68_1403 ();
 sg13g2_fill_2 FILLER_68_1421 ();
 sg13g2_fill_2 FILLER_68_1447 ();
 sg13g2_fill_1 FILLER_68_1449 ();
 sg13g2_decap_8 FILLER_68_1485 ();
 sg13g2_decap_4 FILLER_68_1492 ();
 sg13g2_decap_4 FILLER_68_1512 ();
 sg13g2_fill_1 FILLER_68_1521 ();
 sg13g2_fill_1 FILLER_68_1530 ();
 sg13g2_decap_8 FILLER_68_1536 ();
 sg13g2_decap_8 FILLER_68_1543 ();
 sg13g2_decap_4 FILLER_68_1550 ();
 sg13g2_fill_2 FILLER_68_1564 ();
 sg13g2_fill_2 FILLER_68_1575 ();
 sg13g2_fill_1 FILLER_68_1593 ();
 sg13g2_fill_1 FILLER_68_1603 ();
 sg13g2_fill_1 FILLER_68_1617 ();
 sg13g2_fill_2 FILLER_68_1622 ();
 sg13g2_decap_8 FILLER_68_1628 ();
 sg13g2_decap_8 FILLER_68_1635 ();
 sg13g2_fill_2 FILLER_68_1642 ();
 sg13g2_fill_1 FILLER_68_1644 ();
 sg13g2_fill_2 FILLER_68_1648 ();
 sg13g2_fill_1 FILLER_68_1663 ();
 sg13g2_fill_1 FILLER_68_1722 ();
 sg13g2_decap_4 FILLER_68_1731 ();
 sg13g2_fill_2 FILLER_68_1735 ();
 sg13g2_decap_8 FILLER_68_1741 ();
 sg13g2_decap_8 FILLER_68_1752 ();
 sg13g2_decap_8 FILLER_68_1759 ();
 sg13g2_decap_8 FILLER_68_1766 ();
 sg13g2_fill_1 FILLER_68_1773 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_fill_2 FILLER_69_35 ();
 sg13g2_fill_1 FILLER_69_37 ();
 sg13g2_fill_2 FILLER_69_69 ();
 sg13g2_fill_2 FILLER_69_97 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_4 FILLER_69_119 ();
 sg13g2_fill_1 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_131 ();
 sg13g2_fill_1 FILLER_69_170 ();
 sg13g2_fill_1 FILLER_69_176 ();
 sg13g2_fill_1 FILLER_69_193 ();
 sg13g2_fill_1 FILLER_69_208 ();
 sg13g2_fill_1 FILLER_69_213 ();
 sg13g2_fill_1 FILLER_69_218 ();
 sg13g2_decap_8 FILLER_69_223 ();
 sg13g2_decap_8 FILLER_69_230 ();
 sg13g2_decap_8 FILLER_69_250 ();
 sg13g2_decap_8 FILLER_69_257 ();
 sg13g2_fill_1 FILLER_69_264 ();
 sg13g2_fill_2 FILLER_69_292 ();
 sg13g2_fill_2 FILLER_69_342 ();
 sg13g2_fill_2 FILLER_69_364 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_fill_1 FILLER_69_399 ();
 sg13g2_fill_2 FILLER_69_429 ();
 sg13g2_fill_1 FILLER_69_431 ();
 sg13g2_fill_1 FILLER_69_442 ();
 sg13g2_fill_1 FILLER_69_452 ();
 sg13g2_fill_1 FILLER_69_458 ();
 sg13g2_fill_2 FILLER_69_463 ();
 sg13g2_fill_1 FILLER_69_465 ();
 sg13g2_fill_2 FILLER_69_471 ();
 sg13g2_fill_1 FILLER_69_473 ();
 sg13g2_decap_4 FILLER_69_479 ();
 sg13g2_decap_8 FILLER_69_492 ();
 sg13g2_decap_4 FILLER_69_499 ();
 sg13g2_fill_1 FILLER_69_503 ();
 sg13g2_decap_4 FILLER_69_519 ();
 sg13g2_fill_1 FILLER_69_523 ();
 sg13g2_decap_8 FILLER_69_583 ();
 sg13g2_decap_8 FILLER_69_590 ();
 sg13g2_fill_2 FILLER_69_597 ();
 sg13g2_decap_8 FILLER_69_603 ();
 sg13g2_decap_8 FILLER_69_610 ();
 sg13g2_fill_1 FILLER_69_617 ();
 sg13g2_fill_1 FILLER_69_622 ();
 sg13g2_fill_1 FILLER_69_657 ();
 sg13g2_decap_4 FILLER_69_666 ();
 sg13g2_fill_2 FILLER_69_670 ();
 sg13g2_fill_2 FILLER_69_684 ();
 sg13g2_fill_1 FILLER_69_686 ();
 sg13g2_decap_8 FILLER_69_692 ();
 sg13g2_decap_8 FILLER_69_699 ();
 sg13g2_fill_2 FILLER_69_706 ();
 sg13g2_fill_1 FILLER_69_708 ();
 sg13g2_fill_2 FILLER_69_719 ();
 sg13g2_fill_1 FILLER_69_730 ();
 sg13g2_fill_2 FILLER_69_736 ();
 sg13g2_fill_2 FILLER_69_757 ();
 sg13g2_fill_1 FILLER_69_777 ();
 sg13g2_fill_1 FILLER_69_786 ();
 sg13g2_fill_2 FILLER_69_806 ();
 sg13g2_decap_8 FILLER_69_829 ();
 sg13g2_decap_8 FILLER_69_850 ();
 sg13g2_decap_8 FILLER_69_857 ();
 sg13g2_fill_1 FILLER_69_864 ();
 sg13g2_decap_4 FILLER_69_870 ();
 sg13g2_fill_1 FILLER_69_874 ();
 sg13g2_decap_4 FILLER_69_889 ();
 sg13g2_decap_4 FILLER_69_902 ();
 sg13g2_fill_2 FILLER_69_906 ();
 sg13g2_decap_8 FILLER_69_912 ();
 sg13g2_fill_2 FILLER_69_919 ();
 sg13g2_fill_2 FILLER_69_929 ();
 sg13g2_fill_2 FILLER_69_939 ();
 sg13g2_decap_8 FILLER_69_954 ();
 sg13g2_decap_8 FILLER_69_961 ();
 sg13g2_decap_8 FILLER_69_968 ();
 sg13g2_decap_4 FILLER_69_975 ();
 sg13g2_decap_8 FILLER_69_993 ();
 sg13g2_decap_8 FILLER_69_1000 ();
 sg13g2_fill_2 FILLER_69_1007 ();
 sg13g2_decap_8 FILLER_69_1013 ();
 sg13g2_fill_2 FILLER_69_1020 ();
 sg13g2_fill_1 FILLER_69_1030 ();
 sg13g2_fill_1 FILLER_69_1039 ();
 sg13g2_fill_1 FILLER_69_1044 ();
 sg13g2_fill_1 FILLER_69_1049 ();
 sg13g2_decap_4 FILLER_69_1067 ();
 sg13g2_fill_1 FILLER_69_1071 ();
 sg13g2_decap_8 FILLER_69_1085 ();
 sg13g2_fill_2 FILLER_69_1092 ();
 sg13g2_fill_1 FILLER_69_1094 ();
 sg13g2_fill_1 FILLER_69_1123 ();
 sg13g2_fill_2 FILLER_69_1133 ();
 sg13g2_fill_1 FILLER_69_1135 ();
 sg13g2_fill_2 FILLER_69_1149 ();
 sg13g2_decap_8 FILLER_69_1156 ();
 sg13g2_fill_2 FILLER_69_1163 ();
 sg13g2_fill_1 FILLER_69_1165 ();
 sg13g2_fill_1 FILLER_69_1171 ();
 sg13g2_fill_2 FILLER_69_1178 ();
 sg13g2_fill_2 FILLER_69_1195 ();
 sg13g2_fill_2 FILLER_69_1217 ();
 sg13g2_decap_8 FILLER_69_1223 ();
 sg13g2_decap_8 FILLER_69_1230 ();
 sg13g2_decap_8 FILLER_69_1237 ();
 sg13g2_decap_8 FILLER_69_1244 ();
 sg13g2_decap_4 FILLER_69_1251 ();
 sg13g2_fill_1 FILLER_69_1255 ();
 sg13g2_fill_1 FILLER_69_1260 ();
 sg13g2_fill_1 FILLER_69_1268 ();
 sg13g2_fill_2 FILLER_69_1274 ();
 sg13g2_fill_1 FILLER_69_1280 ();
 sg13g2_fill_1 FILLER_69_1289 ();
 sg13g2_fill_2 FILLER_69_1295 ();
 sg13g2_fill_1 FILLER_69_1297 ();
 sg13g2_fill_1 FILLER_69_1312 ();
 sg13g2_decap_8 FILLER_69_1345 ();
 sg13g2_decap_8 FILLER_69_1356 ();
 sg13g2_decap_8 FILLER_69_1363 ();
 sg13g2_fill_2 FILLER_69_1370 ();
 sg13g2_fill_1 FILLER_69_1386 ();
 sg13g2_fill_2 FILLER_69_1392 ();
 sg13g2_decap_4 FILLER_69_1411 ();
 sg13g2_fill_1 FILLER_69_1415 ();
 sg13g2_fill_2 FILLER_69_1424 ();
 sg13g2_fill_2 FILLER_69_1430 ();
 sg13g2_fill_1 FILLER_69_1432 ();
 sg13g2_fill_1 FILLER_69_1438 ();
 sg13g2_fill_1 FILLER_69_1446 ();
 sg13g2_decap_8 FILLER_69_1463 ();
 sg13g2_fill_2 FILLER_69_1470 ();
 sg13g2_fill_1 FILLER_69_1472 ();
 sg13g2_decap_4 FILLER_69_1486 ();
 sg13g2_decap_8 FILLER_69_1498 ();
 sg13g2_fill_1 FILLER_69_1505 ();
 sg13g2_fill_1 FILLER_69_1514 ();
 sg13g2_decap_4 FILLER_69_1523 ();
 sg13g2_fill_1 FILLER_69_1527 ();
 sg13g2_fill_2 FILLER_69_1554 ();
 sg13g2_fill_2 FILLER_69_1560 ();
 sg13g2_fill_2 FILLER_69_1567 ();
 sg13g2_fill_2 FILLER_69_1582 ();
 sg13g2_fill_1 FILLER_69_1588 ();
 sg13g2_decap_8 FILLER_69_1628 ();
 sg13g2_decap_8 FILLER_69_1635 ();
 sg13g2_fill_2 FILLER_69_1642 ();
 sg13g2_fill_1 FILLER_69_1644 ();
 sg13g2_fill_1 FILLER_69_1657 ();
 sg13g2_decap_8 FILLER_69_1684 ();
 sg13g2_decap_8 FILLER_69_1695 ();
 sg13g2_decap_8 FILLER_69_1702 ();
 sg13g2_fill_2 FILLER_69_1709 ();
 sg13g2_fill_1 FILLER_69_1730 ();
 sg13g2_fill_2 FILLER_69_1739 ();
 sg13g2_fill_2 FILLER_69_1771 ();
 sg13g2_fill_1 FILLER_69_1773 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_4 FILLER_70_39 ();
 sg13g2_fill_1 FILLER_70_43 ();
 sg13g2_decap_8 FILLER_70_48 ();
 sg13g2_decap_8 FILLER_70_55 ();
 sg13g2_fill_1 FILLER_70_62 ();
 sg13g2_decap_4 FILLER_70_67 ();
 sg13g2_fill_2 FILLER_70_71 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_4 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_105 ();
 sg13g2_fill_1 FILLER_70_112 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_fill_2 FILLER_70_125 ();
 sg13g2_fill_2 FILLER_70_137 ();
 sg13g2_fill_1 FILLER_70_139 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_237 ();
 sg13g2_fill_2 FILLER_70_280 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_decap_4 FILLER_70_301 ();
 sg13g2_fill_2 FILLER_70_317 ();
 sg13g2_fill_2 FILLER_70_323 ();
 sg13g2_decap_8 FILLER_70_333 ();
 sg13g2_fill_2 FILLER_70_340 ();
 sg13g2_fill_1 FILLER_70_342 ();
 sg13g2_fill_2 FILLER_70_347 ();
 sg13g2_decap_8 FILLER_70_375 ();
 sg13g2_fill_1 FILLER_70_382 ();
 sg13g2_decap_8 FILLER_70_386 ();
 sg13g2_fill_1 FILLER_70_393 ();
 sg13g2_fill_2 FILLER_70_398 ();
 sg13g2_decap_4 FILLER_70_408 ();
 sg13g2_fill_2 FILLER_70_412 ();
 sg13g2_fill_1 FILLER_70_418 ();
 sg13g2_fill_1 FILLER_70_424 ();
 sg13g2_fill_2 FILLER_70_446 ();
 sg13g2_decap_8 FILLER_70_510 ();
 sg13g2_decap_4 FILLER_70_517 ();
 sg13g2_fill_1 FILLER_70_521 ();
 sg13g2_fill_2 FILLER_70_525 ();
 sg13g2_fill_2 FILLER_70_566 ();
 sg13g2_decap_8 FILLER_70_579 ();
 sg13g2_fill_2 FILLER_70_586 ();
 sg13g2_decap_8 FILLER_70_593 ();
 sg13g2_decap_4 FILLER_70_600 ();
 sg13g2_decap_4 FILLER_70_607 ();
 sg13g2_fill_2 FILLER_70_611 ();
 sg13g2_fill_1 FILLER_70_673 ();
 sg13g2_fill_2 FILLER_70_685 ();
 sg13g2_fill_2 FILLER_70_691 ();
 sg13g2_decap_4 FILLER_70_708 ();
 sg13g2_fill_1 FILLER_70_728 ();
 sg13g2_fill_1 FILLER_70_734 ();
 sg13g2_fill_1 FILLER_70_745 ();
 sg13g2_fill_1 FILLER_70_757 ();
 sg13g2_fill_1 FILLER_70_768 ();
 sg13g2_decap_8 FILLER_70_806 ();
 sg13g2_fill_2 FILLER_70_813 ();
 sg13g2_fill_1 FILLER_70_815 ();
 sg13g2_fill_2 FILLER_70_832 ();
 sg13g2_fill_1 FILLER_70_842 ();
 sg13g2_decap_4 FILLER_70_858 ();
 sg13g2_fill_1 FILLER_70_867 ();
 sg13g2_decap_8 FILLER_70_878 ();
 sg13g2_decap_8 FILLER_70_890 ();
 sg13g2_decap_4 FILLER_70_897 ();
 sg13g2_decap_8 FILLER_70_905 ();
 sg13g2_fill_2 FILLER_70_912 ();
 sg13g2_fill_2 FILLER_70_919 ();
 sg13g2_fill_1 FILLER_70_921 ();
 sg13g2_fill_1 FILLER_70_965 ();
 sg13g2_decap_8 FILLER_70_971 ();
 sg13g2_decap_4 FILLER_70_978 ();
 sg13g2_fill_2 FILLER_70_982 ();
 sg13g2_fill_1 FILLER_70_997 ();
 sg13g2_fill_2 FILLER_70_1003 ();
 sg13g2_fill_1 FILLER_70_1005 ();
 sg13g2_decap_8 FILLER_70_1011 ();
 sg13g2_decap_8 FILLER_70_1018 ();
 sg13g2_decap_4 FILLER_70_1041 ();
 sg13g2_fill_1 FILLER_70_1045 ();
 sg13g2_fill_1 FILLER_70_1051 ();
 sg13g2_fill_2 FILLER_70_1066 ();
 sg13g2_fill_1 FILLER_70_1091 ();
 sg13g2_decap_4 FILLER_70_1108 ();
 sg13g2_fill_2 FILLER_70_1112 ();
 sg13g2_fill_1 FILLER_70_1121 ();
 sg13g2_fill_1 FILLER_70_1127 ();
 sg13g2_decap_8 FILLER_70_1133 ();
 sg13g2_decap_4 FILLER_70_1148 ();
 sg13g2_fill_1 FILLER_70_1152 ();
 sg13g2_fill_1 FILLER_70_1157 ();
 sg13g2_fill_2 FILLER_70_1185 ();
 sg13g2_fill_1 FILLER_70_1220 ();
 sg13g2_decap_4 FILLER_70_1226 ();
 sg13g2_fill_1 FILLER_70_1230 ();
 sg13g2_fill_1 FILLER_70_1235 ();
 sg13g2_decap_4 FILLER_70_1241 ();
 sg13g2_fill_1 FILLER_70_1245 ();
 sg13g2_fill_1 FILLER_70_1297 ();
 sg13g2_decap_8 FILLER_70_1306 ();
 sg13g2_fill_1 FILLER_70_1313 ();
 sg13g2_fill_2 FILLER_70_1319 ();
 sg13g2_fill_1 FILLER_70_1321 ();
 sg13g2_fill_2 FILLER_70_1327 ();
 sg13g2_fill_2 FILLER_70_1337 ();
 sg13g2_decap_8 FILLER_70_1347 ();
 sg13g2_decap_8 FILLER_70_1362 ();
 sg13g2_decap_8 FILLER_70_1369 ();
 sg13g2_decap_8 FILLER_70_1376 ();
 sg13g2_decap_8 FILLER_70_1383 ();
 sg13g2_decap_4 FILLER_70_1390 ();
 sg13g2_decap_4 FILLER_70_1404 ();
 sg13g2_fill_1 FILLER_70_1418 ();
 sg13g2_fill_1 FILLER_70_1426 ();
 sg13g2_fill_1 FILLER_70_1432 ();
 sg13g2_decap_4 FILLER_70_1455 ();
 sg13g2_decap_8 FILLER_70_1463 ();
 sg13g2_fill_2 FILLER_70_1470 ();
 sg13g2_fill_2 FILLER_70_1482 ();
 sg13g2_decap_8 FILLER_70_1488 ();
 sg13g2_decap_8 FILLER_70_1495 ();
 sg13g2_decap_8 FILLER_70_1502 ();
 sg13g2_decap_4 FILLER_70_1509 ();
 sg13g2_fill_1 FILLER_70_1526 ();
 sg13g2_fill_2 FILLER_70_1547 ();
 sg13g2_fill_1 FILLER_70_1578 ();
 sg13g2_fill_2 FILLER_70_1587 ();
 sg13g2_fill_2 FILLER_70_1610 ();
 sg13g2_decap_8 FILLER_70_1620 ();
 sg13g2_decap_4 FILLER_70_1627 ();
 sg13g2_decap_8 FILLER_70_1665 ();
 sg13g2_fill_2 FILLER_70_1672 ();
 sg13g2_fill_2 FILLER_70_1678 ();
 sg13g2_decap_8 FILLER_70_1706 ();
 sg13g2_decap_4 FILLER_70_1721 ();
 sg13g2_fill_1 FILLER_70_1725 ();
 sg13g2_fill_2 FILLER_70_1730 ();
 sg13g2_fill_1 FILLER_70_1736 ();
 sg13g2_decap_8 FILLER_70_1741 ();
 sg13g2_decap_8 FILLER_70_1748 ();
 sg13g2_decap_8 FILLER_70_1755 ();
 sg13g2_decap_8 FILLER_70_1762 ();
 sg13g2_decap_4 FILLER_70_1769 ();
 sg13g2_fill_1 FILLER_70_1773 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_54 ();
 sg13g2_decap_4 FILLER_71_61 ();
 sg13g2_fill_2 FILLER_71_65 ();
 sg13g2_decap_8 FILLER_71_85 ();
 sg13g2_decap_4 FILLER_71_92 ();
 sg13g2_fill_1 FILLER_71_96 ();
 sg13g2_fill_2 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_152 ();
 sg13g2_fill_2 FILLER_71_188 ();
 sg13g2_fill_2 FILLER_71_199 ();
 sg13g2_fill_1 FILLER_71_201 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_224 ();
 sg13g2_fill_2 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_237 ();
 sg13g2_decap_8 FILLER_71_244 ();
 sg13g2_decap_8 FILLER_71_251 ();
 sg13g2_fill_2 FILLER_71_258 ();
 sg13g2_fill_1 FILLER_71_260 ();
 sg13g2_fill_2 FILLER_71_265 ();
 sg13g2_fill_1 FILLER_71_267 ();
 sg13g2_fill_2 FILLER_71_272 ();
 sg13g2_decap_8 FILLER_71_278 ();
 sg13g2_fill_1 FILLER_71_285 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_fill_2 FILLER_71_308 ();
 sg13g2_fill_1 FILLER_71_336 ();
 sg13g2_fill_2 FILLER_71_342 ();
 sg13g2_fill_1 FILLER_71_362 ();
 sg13g2_fill_2 FILLER_71_373 ();
 sg13g2_decap_4 FILLER_71_386 ();
 sg13g2_fill_2 FILLER_71_390 ();
 sg13g2_decap_4 FILLER_71_396 ();
 sg13g2_fill_1 FILLER_71_400 ();
 sg13g2_decap_4 FILLER_71_409 ();
 sg13g2_fill_1 FILLER_71_434 ();
 sg13g2_fill_2 FILLER_71_476 ();
 sg13g2_decap_4 FILLER_71_492 ();
 sg13g2_fill_1 FILLER_71_496 ();
 sg13g2_decap_4 FILLER_71_507 ();
 sg13g2_fill_1 FILLER_71_511 ();
 sg13g2_fill_1 FILLER_71_521 ();
 sg13g2_fill_2 FILLER_71_562 ();
 sg13g2_fill_2 FILLER_71_574 ();
 sg13g2_fill_1 FILLER_71_576 ();
 sg13g2_decap_4 FILLER_71_581 ();
 sg13g2_fill_1 FILLER_71_585 ();
 sg13g2_fill_1 FILLER_71_594 ();
 sg13g2_fill_2 FILLER_71_599 ();
 sg13g2_fill_1 FILLER_71_605 ();
 sg13g2_fill_2 FILLER_71_610 ();
 sg13g2_fill_2 FILLER_71_617 ();
 sg13g2_fill_2 FILLER_71_627 ();
 sg13g2_fill_1 FILLER_71_634 ();
 sg13g2_fill_1 FILLER_71_662 ();
 sg13g2_decap_8 FILLER_71_676 ();
 sg13g2_decap_8 FILLER_71_683 ();
 sg13g2_decap_8 FILLER_71_690 ();
 sg13g2_decap_8 FILLER_71_706 ();
 sg13g2_decap_8 FILLER_71_713 ();
 sg13g2_fill_2 FILLER_71_720 ();
 sg13g2_fill_1 FILLER_71_722 ();
 sg13g2_decap_4 FILLER_71_735 ();
 sg13g2_decap_4 FILLER_71_744 ();
 sg13g2_fill_1 FILLER_71_759 ();
 sg13g2_fill_1 FILLER_71_764 ();
 sg13g2_fill_1 FILLER_71_769 ();
 sg13g2_fill_2 FILLER_71_789 ();
 sg13g2_decap_8 FILLER_71_806 ();
 sg13g2_decap_8 FILLER_71_813 ();
 sg13g2_decap_4 FILLER_71_820 ();
 sg13g2_fill_1 FILLER_71_824 ();
 sg13g2_decap_4 FILLER_71_833 ();
 sg13g2_fill_2 FILLER_71_837 ();
 sg13g2_decap_8 FILLER_71_853 ();
 sg13g2_decap_8 FILLER_71_860 ();
 sg13g2_decap_8 FILLER_71_867 ();
 sg13g2_decap_8 FILLER_71_879 ();
 sg13g2_decap_8 FILLER_71_891 ();
 sg13g2_decap_8 FILLER_71_898 ();
 sg13g2_fill_2 FILLER_71_905 ();
 sg13g2_fill_1 FILLER_71_907 ();
 sg13g2_fill_1 FILLER_71_916 ();
 sg13g2_fill_1 FILLER_71_922 ();
 sg13g2_fill_1 FILLER_71_929 ();
 sg13g2_fill_1 FILLER_71_941 ();
 sg13g2_fill_2 FILLER_71_956 ();
 sg13g2_decap_8 FILLER_71_971 ();
 sg13g2_fill_1 FILLER_71_978 ();
 sg13g2_fill_2 FILLER_71_999 ();
 sg13g2_fill_1 FILLER_71_1001 ();
 sg13g2_decap_8 FILLER_71_1015 ();
 sg13g2_decap_8 FILLER_71_1022 ();
 sg13g2_decap_8 FILLER_71_1029 ();
 sg13g2_decap_4 FILLER_71_1036 ();
 sg13g2_fill_1 FILLER_71_1040 ();
 sg13g2_fill_2 FILLER_71_1049 ();
 sg13g2_fill_1 FILLER_71_1051 ();
 sg13g2_decap_8 FILLER_71_1089 ();
 sg13g2_fill_2 FILLER_71_1096 ();
 sg13g2_fill_1 FILLER_71_1098 ();
 sg13g2_decap_4 FILLER_71_1104 ();
 sg13g2_fill_1 FILLER_71_1108 ();
 sg13g2_decap_4 FILLER_71_1113 ();
 sg13g2_decap_4 FILLER_71_1125 ();
 sg13g2_decap_8 FILLER_71_1133 ();
 sg13g2_fill_2 FILLER_71_1193 ();
 sg13g2_fill_1 FILLER_71_1199 ();
 sg13g2_fill_2 FILLER_71_1220 ();
 sg13g2_decap_8 FILLER_71_1241 ();
 sg13g2_fill_2 FILLER_71_1256 ();
 sg13g2_fill_2 FILLER_71_1262 ();
 sg13g2_fill_1 FILLER_71_1264 ();
 sg13g2_fill_1 FILLER_71_1286 ();
 sg13g2_decap_8 FILLER_71_1296 ();
 sg13g2_decap_4 FILLER_71_1303 ();
 sg13g2_decap_8 FILLER_71_1310 ();
 sg13g2_decap_8 FILLER_71_1317 ();
 sg13g2_decap_8 FILLER_71_1324 ();
 sg13g2_fill_1 FILLER_71_1336 ();
 sg13g2_fill_2 FILLER_71_1345 ();
 sg13g2_fill_1 FILLER_71_1347 ();
 sg13g2_decap_8 FILLER_71_1357 ();
 sg13g2_decap_4 FILLER_71_1364 ();
 sg13g2_decap_4 FILLER_71_1373 ();
 sg13g2_fill_1 FILLER_71_1377 ();
 sg13g2_decap_4 FILLER_71_1383 ();
 sg13g2_fill_2 FILLER_71_1387 ();
 sg13g2_decap_4 FILLER_71_1403 ();
 sg13g2_decap_8 FILLER_71_1418 ();
 sg13g2_fill_1 FILLER_71_1438 ();
 sg13g2_fill_1 FILLER_71_1449 ();
 sg13g2_fill_2 FILLER_71_1473 ();
 sg13g2_decap_8 FILLER_71_1488 ();
 sg13g2_decap_4 FILLER_71_1495 ();
 sg13g2_decap_8 FILLER_71_1534 ();
 sg13g2_decap_4 FILLER_71_1541 ();
 sg13g2_fill_1 FILLER_71_1545 ();
 sg13g2_decap_4 FILLER_71_1591 ();
 sg13g2_fill_1 FILLER_71_1595 ();
 sg13g2_fill_1 FILLER_71_1601 ();
 sg13g2_decap_4 FILLER_71_1607 ();
 sg13g2_decap_8 FILLER_71_1619 ();
 sg13g2_decap_8 FILLER_71_1626 ();
 sg13g2_fill_1 FILLER_71_1633 ();
 sg13g2_decap_4 FILLER_71_1638 ();
 sg13g2_decap_4 FILLER_71_1658 ();
 sg13g2_fill_2 FILLER_71_1691 ();
 sg13g2_decap_8 FILLER_71_1708 ();
 sg13g2_fill_2 FILLER_71_1715 ();
 sg13g2_fill_1 FILLER_71_1717 ();
 sg13g2_decap_8 FILLER_71_1748 ();
 sg13g2_decap_8 FILLER_71_1755 ();
 sg13g2_decap_8 FILLER_71_1762 ();
 sg13g2_decap_4 FILLER_71_1769 ();
 sg13g2_fill_1 FILLER_71_1773 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_fill_1 FILLER_72_42 ();
 sg13g2_decap_4 FILLER_72_69 ();
 sg13g2_fill_2 FILLER_72_73 ();
 sg13g2_fill_1 FILLER_72_79 ();
 sg13g2_fill_1 FILLER_72_84 ();
 sg13g2_fill_2 FILLER_72_90 ();
 sg13g2_decap_4 FILLER_72_102 ();
 sg13g2_decap_4 FILLER_72_118 ();
 sg13g2_fill_1 FILLER_72_122 ();
 sg13g2_decap_4 FILLER_72_134 ();
 sg13g2_fill_2 FILLER_72_138 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_fill_2 FILLER_72_224 ();
 sg13g2_fill_2 FILLER_72_256 ();
 sg13g2_fill_1 FILLER_72_258 ();
 sg13g2_fill_2 FILLER_72_264 ();
 sg13g2_fill_1 FILLER_72_266 ();
 sg13g2_fill_2 FILLER_72_271 ();
 sg13g2_fill_1 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_314 ();
 sg13g2_decap_8 FILLER_72_321 ();
 sg13g2_decap_4 FILLER_72_328 ();
 sg13g2_fill_2 FILLER_72_332 ();
 sg13g2_fill_2 FILLER_72_347 ();
 sg13g2_fill_2 FILLER_72_376 ();
 sg13g2_decap_8 FILLER_72_415 ();
 sg13g2_fill_2 FILLER_72_427 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_fill_1 FILLER_72_438 ();
 sg13g2_decap_8 FILLER_72_443 ();
 sg13g2_decap_8 FILLER_72_450 ();
 sg13g2_decap_8 FILLER_72_457 ();
 sg13g2_fill_1 FILLER_72_464 ();
 sg13g2_fill_1 FILLER_72_469 ();
 sg13g2_decap_8 FILLER_72_478 ();
 sg13g2_decap_4 FILLER_72_485 ();
 sg13g2_fill_2 FILLER_72_489 ();
 sg13g2_fill_2 FILLER_72_500 ();
 sg13g2_fill_2 FILLER_72_505 ();
 sg13g2_fill_2 FILLER_72_512 ();
 sg13g2_fill_1 FILLER_72_543 ();
 sg13g2_decap_8 FILLER_72_565 ();
 sg13g2_decap_4 FILLER_72_572 ();
 sg13g2_decap_4 FILLER_72_607 ();
 sg13g2_fill_2 FILLER_72_615 ();
 sg13g2_fill_1 FILLER_72_617 ();
 sg13g2_fill_1 FILLER_72_656 ();
 sg13g2_fill_1 FILLER_72_670 ();
 sg13g2_decap_8 FILLER_72_676 ();
 sg13g2_decap_4 FILLER_72_683 ();
 sg13g2_fill_2 FILLER_72_687 ();
 sg13g2_fill_1 FILLER_72_712 ();
 sg13g2_decap_4 FILLER_72_721 ();
 sg13g2_decap_8 FILLER_72_733 ();
 sg13g2_decap_8 FILLER_72_740 ();
 sg13g2_decap_4 FILLER_72_747 ();
 sg13g2_fill_1 FILLER_72_751 ();
 sg13g2_fill_2 FILLER_72_765 ();
 sg13g2_fill_1 FILLER_72_786 ();
 sg13g2_fill_2 FILLER_72_800 ();
 sg13g2_decap_8 FILLER_72_807 ();
 sg13g2_fill_1 FILLER_72_826 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_decap_4 FILLER_72_878 ();
 sg13g2_fill_1 FILLER_72_882 ();
 sg13g2_fill_1 FILLER_72_910 ();
 sg13g2_fill_1 FILLER_72_928 ();
 sg13g2_fill_2 FILLER_72_952 ();
 sg13g2_decap_8 FILLER_72_963 ();
 sg13g2_decap_8 FILLER_72_970 ();
 sg13g2_fill_1 FILLER_72_994 ();
 sg13g2_fill_2 FILLER_72_1005 ();
 sg13g2_fill_2 FILLER_72_1022 ();
 sg13g2_fill_2 FILLER_72_1037 ();
 sg13g2_fill_1 FILLER_72_1039 ();
 sg13g2_fill_2 FILLER_72_1045 ();
 sg13g2_fill_1 FILLER_72_1047 ();
 sg13g2_decap_8 FILLER_72_1061 ();
 sg13g2_decap_8 FILLER_72_1068 ();
 sg13g2_decap_4 FILLER_72_1075 ();
 sg13g2_decap_4 FILLER_72_1084 ();
 sg13g2_fill_1 FILLER_72_1102 ();
 sg13g2_decap_8 FILLER_72_1127 ();
 sg13g2_decap_8 FILLER_72_1134 ();
 sg13g2_decap_4 FILLER_72_1156 ();
 sg13g2_fill_2 FILLER_72_1179 ();
 sg13g2_fill_1 FILLER_72_1190 ();
 sg13g2_fill_2 FILLER_72_1227 ();
 sg13g2_fill_1 FILLER_72_1229 ();
 sg13g2_fill_1 FILLER_72_1247 ();
 sg13g2_decap_4 FILLER_72_1252 ();
 sg13g2_fill_1 FILLER_72_1256 ();
 sg13g2_fill_1 FILLER_72_1262 ();
 sg13g2_fill_2 FILLER_72_1272 ();
 sg13g2_fill_1 FILLER_72_1274 ();
 sg13g2_decap_4 FILLER_72_1285 ();
 sg13g2_fill_1 FILLER_72_1289 ();
 sg13g2_fill_1 FILLER_72_1308 ();
 sg13g2_fill_1 FILLER_72_1313 ();
 sg13g2_decap_8 FILLER_72_1319 ();
 sg13g2_decap_8 FILLER_72_1326 ();
 sg13g2_fill_1 FILLER_72_1333 ();
 sg13g2_fill_1 FILLER_72_1337 ();
 sg13g2_decap_8 FILLER_72_1360 ();
 sg13g2_decap_8 FILLER_72_1367 ();
 sg13g2_fill_1 FILLER_72_1379 ();
 sg13g2_fill_2 FILLER_72_1390 ();
 sg13g2_fill_2 FILLER_72_1397 ();
 sg13g2_fill_1 FILLER_72_1418 ();
 sg13g2_fill_2 FILLER_72_1437 ();
 sg13g2_fill_2 FILLER_72_1448 ();
 sg13g2_fill_2 FILLER_72_1470 ();
 sg13g2_fill_1 FILLER_72_1472 ();
 sg13g2_fill_1 FILLER_72_1478 ();
 sg13g2_decap_4 FILLER_72_1494 ();
 sg13g2_fill_1 FILLER_72_1498 ();
 sg13g2_fill_2 FILLER_72_1504 ();
 sg13g2_fill_1 FILLER_72_1506 ();
 sg13g2_decap_8 FILLER_72_1511 ();
 sg13g2_fill_1 FILLER_72_1518 ();
 sg13g2_decap_8 FILLER_72_1527 ();
 sg13g2_decap_8 FILLER_72_1534 ();
 sg13g2_fill_2 FILLER_72_1541 ();
 sg13g2_fill_1 FILLER_72_1543 ();
 sg13g2_fill_1 FILLER_72_1573 ();
 sg13g2_decap_8 FILLER_72_1583 ();
 sg13g2_decap_8 FILLER_72_1590 ();
 sg13g2_fill_2 FILLER_72_1602 ();
 sg13g2_fill_2 FILLER_72_1646 ();
 sg13g2_decap_8 FILLER_72_1653 ();
 sg13g2_fill_1 FILLER_72_1660 ();
 sg13g2_fill_1 FILLER_72_1673 ();
 sg13g2_decap_8 FILLER_72_1704 ();
 sg13g2_decap_8 FILLER_72_1711 ();
 sg13g2_decap_8 FILLER_72_1718 ();
 sg13g2_fill_1 FILLER_72_1725 ();
 sg13g2_decap_8 FILLER_72_1730 ();
 sg13g2_decap_8 FILLER_72_1737 ();
 sg13g2_decap_8 FILLER_72_1744 ();
 sg13g2_decap_8 FILLER_72_1751 ();
 sg13g2_decap_8 FILLER_72_1758 ();
 sg13g2_decap_8 FILLER_72_1765 ();
 sg13g2_fill_2 FILLER_72_1772 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_54 ();
 sg13g2_fill_2 FILLER_73_61 ();
 sg13g2_fill_2 FILLER_73_73 ();
 sg13g2_fill_1 FILLER_73_75 ();
 sg13g2_decap_8 FILLER_73_81 ();
 sg13g2_fill_2 FILLER_73_88 ();
 sg13g2_decap_8 FILLER_73_128 ();
 sg13g2_fill_2 FILLER_73_135 ();
 sg13g2_fill_1 FILLER_73_137 ();
 sg13g2_decap_4 FILLER_73_142 ();
 sg13g2_fill_2 FILLER_73_146 ();
 sg13g2_fill_1 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_190 ();
 sg13g2_fill_1 FILLER_73_201 ();
 sg13g2_decap_8 FILLER_73_209 ();
 sg13g2_decap_8 FILLER_73_228 ();
 sg13g2_fill_2 FILLER_73_235 ();
 sg13g2_fill_1 FILLER_73_256 ();
 sg13g2_fill_1 FILLER_73_262 ();
 sg13g2_fill_2 FILLER_73_267 ();
 sg13g2_fill_1 FILLER_73_305 ();
 sg13g2_fill_2 FILLER_73_326 ();
 sg13g2_fill_1 FILLER_73_328 ();
 sg13g2_decap_4 FILLER_73_333 ();
 sg13g2_fill_1 FILLER_73_342 ();
 sg13g2_fill_1 FILLER_73_369 ();
 sg13g2_decap_4 FILLER_73_385 ();
 sg13g2_fill_1 FILLER_73_389 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_decap_8 FILLER_73_427 ();
 sg13g2_decap_8 FILLER_73_434 ();
 sg13g2_decap_8 FILLER_73_441 ();
 sg13g2_decap_8 FILLER_73_448 ();
 sg13g2_decap_8 FILLER_73_455 ();
 sg13g2_decap_8 FILLER_73_462 ();
 sg13g2_decap_4 FILLER_73_469 ();
 sg13g2_fill_2 FILLER_73_473 ();
 sg13g2_fill_2 FILLER_73_522 ();
 sg13g2_fill_1 FILLER_73_538 ();
 sg13g2_fill_1 FILLER_73_551 ();
 sg13g2_decap_4 FILLER_73_559 ();
 sg13g2_fill_1 FILLER_73_563 ();
 sg13g2_decap_8 FILLER_73_569 ();
 sg13g2_fill_1 FILLER_73_576 ();
 sg13g2_fill_2 FILLER_73_582 ();
 sg13g2_fill_1 FILLER_73_588 ();
 sg13g2_fill_2 FILLER_73_593 ();
 sg13g2_fill_1 FILLER_73_595 ();
 sg13g2_fill_2 FILLER_73_609 ();
 sg13g2_fill_1 FILLER_73_611 ();
 sg13g2_fill_2 FILLER_73_617 ();
 sg13g2_fill_1 FILLER_73_634 ();
 sg13g2_decap_4 FILLER_73_667 ();
 sg13g2_fill_2 FILLER_73_675 ();
 sg13g2_decap_4 FILLER_73_681 ();
 sg13g2_fill_2 FILLER_73_685 ();
 sg13g2_fill_1 FILLER_73_692 ();
 sg13g2_fill_2 FILLER_73_745 ();
 sg13g2_fill_2 FILLER_73_758 ();
 sg13g2_decap_4 FILLER_73_772 ();
 sg13g2_fill_2 FILLER_73_791 ();
 sg13g2_fill_1 FILLER_73_793 ();
 sg13g2_fill_2 FILLER_73_797 ();
 sg13g2_fill_2 FILLER_73_803 ();
 sg13g2_fill_2 FILLER_73_809 ();
 sg13g2_fill_1 FILLER_73_811 ();
 sg13g2_fill_1 FILLER_73_815 ();
 sg13g2_fill_1 FILLER_73_855 ();
 sg13g2_decap_8 FILLER_73_866 ();
 sg13g2_decap_8 FILLER_73_873 ();
 sg13g2_fill_2 FILLER_73_880 ();
 sg13g2_fill_1 FILLER_73_891 ();
 sg13g2_fill_1 FILLER_73_905 ();
 sg13g2_fill_1 FILLER_73_914 ();
 sg13g2_fill_2 FILLER_73_929 ();
 sg13g2_fill_1 FILLER_73_947 ();
 sg13g2_fill_2 FILLER_73_970 ();
 sg13g2_fill_1 FILLER_73_972 ();
 sg13g2_fill_2 FILLER_73_989 ();
 sg13g2_fill_1 FILLER_73_999 ();
 sg13g2_fill_1 FILLER_73_1013 ();
 sg13g2_decap_4 FILLER_73_1026 ();
 sg13g2_fill_1 FILLER_73_1030 ();
 sg13g2_decap_4 FILLER_73_1048 ();
 sg13g2_fill_1 FILLER_73_1057 ();
 sg13g2_fill_2 FILLER_73_1062 ();
 sg13g2_fill_1 FILLER_73_1069 ();
 sg13g2_fill_2 FILLER_73_1076 ();
 sg13g2_fill_1 FILLER_73_1104 ();
 sg13g2_decap_8 FILLER_73_1127 ();
 sg13g2_fill_1 FILLER_73_1134 ();
 sg13g2_fill_2 FILLER_73_1155 ();
 sg13g2_fill_1 FILLER_73_1170 ();
 sg13g2_fill_2 FILLER_73_1177 ();
 sg13g2_fill_1 FILLER_73_1198 ();
 sg13g2_fill_1 FILLER_73_1207 ();
 sg13g2_decap_8 FILLER_73_1223 ();
 sg13g2_decap_8 FILLER_73_1230 ();
 sg13g2_decap_8 FILLER_73_1237 ();
 sg13g2_decap_4 FILLER_73_1244 ();
 sg13g2_fill_1 FILLER_73_1248 ();
 sg13g2_decap_4 FILLER_73_1254 ();
 sg13g2_fill_2 FILLER_73_1258 ();
 sg13g2_fill_1 FILLER_73_1273 ();
 sg13g2_fill_1 FILLER_73_1278 ();
 sg13g2_fill_2 FILLER_73_1331 ();
 sg13g2_fill_1 FILLER_73_1333 ();
 sg13g2_decap_4 FILLER_73_1346 ();
 sg13g2_decap_8 FILLER_73_1366 ();
 sg13g2_decap_4 FILLER_73_1373 ();
 sg13g2_fill_1 FILLER_73_1385 ();
 sg13g2_fill_2 FILLER_73_1408 ();
 sg13g2_fill_1 FILLER_73_1418 ();
 sg13g2_fill_1 FILLER_73_1432 ();
 sg13g2_decap_8 FILLER_73_1505 ();
 sg13g2_fill_2 FILLER_73_1525 ();
 sg13g2_fill_1 FILLER_73_1527 ();
 sg13g2_decap_8 FILLER_73_1532 ();
 sg13g2_fill_2 FILLER_73_1542 ();
 sg13g2_fill_1 FILLER_73_1544 ();
 sg13g2_decap_4 FILLER_73_1552 ();
 sg13g2_fill_2 FILLER_73_1556 ();
 sg13g2_decap_8 FILLER_73_1563 ();
 sg13g2_decap_8 FILLER_73_1570 ();
 sg13g2_fill_2 FILLER_73_1577 ();
 sg13g2_decap_8 FILLER_73_1605 ();
 sg13g2_decap_8 FILLER_73_1612 ();
 sg13g2_decap_8 FILLER_73_1619 ();
 sg13g2_fill_2 FILLER_73_1626 ();
 sg13g2_fill_2 FILLER_73_1632 ();
 sg13g2_fill_2 FILLER_73_1645 ();
 sg13g2_decap_8 FILLER_73_1655 ();
 sg13g2_decap_8 FILLER_73_1662 ();
 sg13g2_fill_1 FILLER_73_1674 ();
 sg13g2_decap_8 FILLER_73_1685 ();
 sg13g2_decap_4 FILLER_73_1692 ();
 sg13g2_fill_2 FILLER_73_1717 ();
 sg13g2_decap_8 FILLER_73_1745 ();
 sg13g2_decap_8 FILLER_73_1752 ();
 sg13g2_decap_8 FILLER_73_1759 ();
 sg13g2_decap_8 FILLER_73_1766 ();
 sg13g2_fill_1 FILLER_73_1773 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_fill_1 FILLER_74_58 ();
 sg13g2_decap_4 FILLER_74_63 ();
 sg13g2_fill_1 FILLER_74_67 ();
 sg13g2_fill_1 FILLER_74_97 ();
 sg13g2_fill_2 FILLER_74_102 ();
 sg13g2_fill_1 FILLER_74_104 ();
 sg13g2_decap_4 FILLER_74_131 ();
 sg13g2_fill_1 FILLER_74_135 ();
 sg13g2_decap_4 FILLER_74_141 ();
 sg13g2_fill_2 FILLER_74_150 ();
 sg13g2_fill_1 FILLER_74_152 ();
 sg13g2_fill_2 FILLER_74_161 ();
 sg13g2_fill_1 FILLER_74_163 ();
 sg13g2_fill_2 FILLER_74_189 ();
 sg13g2_fill_2 FILLER_74_196 ();
 sg13g2_fill_2 FILLER_74_201 ();
 sg13g2_fill_1 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_230 ();
 sg13g2_fill_1 FILLER_74_240 ();
 sg13g2_fill_1 FILLER_74_249 ();
 sg13g2_decap_8 FILLER_74_264 ();
 sg13g2_fill_1 FILLER_74_271 ();
 sg13g2_fill_2 FILLER_74_283 ();
 sg13g2_fill_1 FILLER_74_298 ();
 sg13g2_fill_2 FILLER_74_307 ();
 sg13g2_fill_1 FILLER_74_314 ();
 sg13g2_fill_1 FILLER_74_324 ();
 sg13g2_decap_8 FILLER_74_332 ();
 sg13g2_decap_8 FILLER_74_339 ();
 sg13g2_fill_2 FILLER_74_346 ();
 sg13g2_fill_1 FILLER_74_348 ();
 sg13g2_decap_4 FILLER_74_353 ();
 sg13g2_fill_1 FILLER_74_360 ();
 sg13g2_decap_8 FILLER_74_400 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_fill_1 FILLER_74_409 ();
 sg13g2_decap_4 FILLER_74_417 ();
 sg13g2_fill_2 FILLER_74_421 ();
 sg13g2_fill_1 FILLER_74_426 ();
 sg13g2_decap_8 FILLER_74_432 ();
 sg13g2_fill_2 FILLER_74_439 ();
 sg13g2_decap_8 FILLER_74_451 ();
 sg13g2_decap_4 FILLER_74_458 ();
 sg13g2_decap_8 FILLER_74_474 ();
 sg13g2_decap_4 FILLER_74_481 ();
 sg13g2_fill_1 FILLER_74_489 ();
 sg13g2_decap_8 FILLER_74_494 ();
 sg13g2_fill_2 FILLER_74_501 ();
 sg13g2_fill_1 FILLER_74_503 ();
 sg13g2_decap_4 FILLER_74_515 ();
 sg13g2_decap_8 FILLER_74_523 ();
 sg13g2_decap_8 FILLER_74_530 ();
 sg13g2_decap_8 FILLER_74_537 ();
 sg13g2_decap_8 FILLER_74_544 ();
 sg13g2_fill_2 FILLER_74_551 ();
 sg13g2_fill_1 FILLER_74_553 ();
 sg13g2_fill_2 FILLER_74_562 ();
 sg13g2_fill_1 FILLER_74_564 ();
 sg13g2_decap_8 FILLER_74_570 ();
 sg13g2_fill_1 FILLER_74_577 ();
 sg13g2_fill_1 FILLER_74_597 ();
 sg13g2_fill_1 FILLER_74_607 ();
 sg13g2_fill_1 FILLER_74_618 ();
 sg13g2_decap_8 FILLER_74_661 ();
 sg13g2_decap_8 FILLER_74_668 ();
 sg13g2_decap_8 FILLER_74_675 ();
 sg13g2_fill_2 FILLER_74_682 ();
 sg13g2_fill_1 FILLER_74_684 ();
 sg13g2_fill_2 FILLER_74_701 ();
 sg13g2_decap_4 FILLER_74_708 ();
 sg13g2_fill_1 FILLER_74_712 ();
 sg13g2_fill_1 FILLER_74_729 ();
 sg13g2_fill_1 FILLER_74_735 ();
 sg13g2_fill_1 FILLER_74_741 ();
 sg13g2_fill_1 FILLER_74_750 ();
 sg13g2_fill_1 FILLER_74_759 ();
 sg13g2_fill_2 FILLER_74_766 ();
 sg13g2_fill_2 FILLER_74_773 ();
 sg13g2_fill_1 FILLER_74_786 ();
 sg13g2_fill_2 FILLER_74_796 ();
 sg13g2_fill_1 FILLER_74_802 ();
 sg13g2_fill_1 FILLER_74_813 ();
 sg13g2_fill_2 FILLER_74_820 ();
 sg13g2_fill_2 FILLER_74_827 ();
 sg13g2_fill_2 FILLER_74_850 ();
 sg13g2_fill_1 FILLER_74_852 ();
 sg13g2_decap_8 FILLER_74_868 ();
 sg13g2_decap_8 FILLER_74_875 ();
 sg13g2_fill_1 FILLER_74_882 ();
 sg13g2_decap_4 FILLER_74_888 ();
 sg13g2_fill_2 FILLER_74_892 ();
 sg13g2_decap_8 FILLER_74_903 ();
 sg13g2_fill_2 FILLER_74_926 ();
 sg13g2_fill_2 FILLER_74_932 ();
 sg13g2_fill_1 FILLER_74_956 ();
 sg13g2_fill_1 FILLER_74_962 ();
 sg13g2_fill_1 FILLER_74_967 ();
 sg13g2_fill_1 FILLER_74_983 ();
 sg13g2_fill_1 FILLER_74_1000 ();
 sg13g2_fill_2 FILLER_74_1009 ();
 sg13g2_decap_8 FILLER_74_1019 ();
 sg13g2_decap_8 FILLER_74_1026 ();
 sg13g2_decap_8 FILLER_74_1033 ();
 sg13g2_decap_8 FILLER_74_1040 ();
 sg13g2_fill_2 FILLER_74_1047 ();
 sg13g2_fill_1 FILLER_74_1049 ();
 sg13g2_fill_1 FILLER_74_1063 ();
 sg13g2_decap_8 FILLER_74_1068 ();
 sg13g2_fill_1 FILLER_74_1075 ();
 sg13g2_fill_2 FILLER_74_1081 ();
 sg13g2_decap_8 FILLER_74_1108 ();
 sg13g2_decap_8 FILLER_74_1115 ();
 sg13g2_decap_8 FILLER_74_1122 ();
 sg13g2_fill_2 FILLER_74_1134 ();
 sg13g2_fill_1 FILLER_74_1136 ();
 sg13g2_fill_2 FILLER_74_1142 ();
 sg13g2_fill_1 FILLER_74_1144 ();
 sg13g2_fill_1 FILLER_74_1164 ();
 sg13g2_fill_2 FILLER_74_1191 ();
 sg13g2_decap_4 FILLER_74_1222 ();
 sg13g2_decap_8 FILLER_74_1230 ();
 sg13g2_fill_2 FILLER_74_1237 ();
 sg13g2_fill_1 FILLER_74_1239 ();
 sg13g2_decap_4 FILLER_74_1249 ();
 sg13g2_decap_8 FILLER_74_1257 ();
 sg13g2_fill_2 FILLER_74_1282 ();
 sg13g2_fill_1 FILLER_74_1284 ();
 sg13g2_fill_2 FILLER_74_1289 ();
 sg13g2_fill_1 FILLER_74_1291 ();
 sg13g2_fill_1 FILLER_74_1303 ();
 sg13g2_fill_1 FILLER_74_1323 ();
 sg13g2_fill_1 FILLER_74_1336 ();
 sg13g2_decap_8 FILLER_74_1341 ();
 sg13g2_fill_2 FILLER_74_1348 ();
 sg13g2_decap_8 FILLER_74_1363 ();
 sg13g2_decap_4 FILLER_74_1370 ();
 sg13g2_decap_4 FILLER_74_1382 ();
 sg13g2_decap_4 FILLER_74_1390 ();
 sg13g2_fill_2 FILLER_74_1394 ();
 sg13g2_decap_8 FILLER_74_1407 ();
 sg13g2_decap_4 FILLER_74_1414 ();
 sg13g2_fill_2 FILLER_74_1440 ();
 sg13g2_fill_1 FILLER_74_1447 ();
 sg13g2_fill_2 FILLER_74_1472 ();
 sg13g2_decap_8 FILLER_74_1490 ();
 sg13g2_fill_2 FILLER_74_1497 ();
 sg13g2_decap_8 FILLER_74_1529 ();
 sg13g2_decap_8 FILLER_74_1536 ();
 sg13g2_decap_8 FILLER_74_1543 ();
 sg13g2_decap_8 FILLER_74_1550 ();
 sg13g2_decap_4 FILLER_74_1583 ();
 sg13g2_fill_1 FILLER_74_1587 ();
 sg13g2_decap_4 FILLER_74_1592 ();
 sg13g2_fill_2 FILLER_74_1596 ();
 sg13g2_fill_2 FILLER_74_1641 ();
 sg13g2_fill_1 FILLER_74_1646 ();
 sg13g2_decap_4 FILLER_74_1660 ();
 sg13g2_fill_2 FILLER_74_1664 ();
 sg13g2_fill_2 FILLER_74_1680 ();
 sg13g2_fill_1 FILLER_74_1682 ();
 sg13g2_fill_2 FILLER_74_1709 ();
 sg13g2_decap_4 FILLER_74_1723 ();
 sg13g2_fill_2 FILLER_74_1739 ();
 sg13g2_fill_1 FILLER_74_1741 ();
 sg13g2_decap_4 FILLER_74_1768 ();
 sg13g2_fill_2 FILLER_74_1772 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_4 FILLER_75_70 ();
 sg13g2_fill_2 FILLER_75_74 ();
 sg13g2_decap_4 FILLER_75_80 ();
 sg13g2_fill_2 FILLER_75_84 ();
 sg13g2_fill_2 FILLER_75_89 ();
 sg13g2_decap_8 FILLER_75_103 ();
 sg13g2_decap_8 FILLER_75_110 ();
 sg13g2_fill_1 FILLER_75_117 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_fill_1 FILLER_75_171 ();
 sg13g2_decap_4 FILLER_75_178 ();
 sg13g2_fill_1 FILLER_75_182 ();
 sg13g2_fill_2 FILLER_75_188 ();
 sg13g2_fill_2 FILLER_75_195 ();
 sg13g2_fill_1 FILLER_75_197 ();
 sg13g2_fill_1 FILLER_75_209 ();
 sg13g2_decap_4 FILLER_75_214 ();
 sg13g2_fill_1 FILLER_75_218 ();
 sg13g2_fill_2 FILLER_75_223 ();
 sg13g2_fill_1 FILLER_75_225 ();
 sg13g2_fill_1 FILLER_75_233 ();
 sg13g2_decap_4 FILLER_75_243 ();
 sg13g2_fill_1 FILLER_75_271 ();
 sg13g2_decap_4 FILLER_75_282 ();
 sg13g2_fill_2 FILLER_75_312 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_decap_8 FILLER_75_339 ();
 sg13g2_decap_8 FILLER_75_346 ();
 sg13g2_fill_2 FILLER_75_353 ();
 sg13g2_fill_1 FILLER_75_355 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_decap_8 FILLER_75_367 ();
 sg13g2_fill_2 FILLER_75_374 ();
 sg13g2_decap_8 FILLER_75_380 ();
 sg13g2_decap_8 FILLER_75_387 ();
 sg13g2_fill_2 FILLER_75_394 ();
 sg13g2_decap_4 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_404 ();
 sg13g2_fill_2 FILLER_75_440 ();
 sg13g2_fill_1 FILLER_75_447 ();
 sg13g2_fill_2 FILLER_75_458 ();
 sg13g2_fill_1 FILLER_75_460 ();
 sg13g2_decap_4 FILLER_75_470 ();
 sg13g2_fill_2 FILLER_75_474 ();
 sg13g2_fill_2 FILLER_75_490 ();
 sg13g2_decap_8 FILLER_75_504 ();
 sg13g2_fill_2 FILLER_75_537 ();
 sg13g2_decap_8 FILLER_75_543 ();
 sg13g2_fill_1 FILLER_75_550 ();
 sg13g2_fill_2 FILLER_75_571 ();
 sg13g2_fill_1 FILLER_75_573 ();
 sg13g2_fill_2 FILLER_75_579 ();
 sg13g2_fill_1 FILLER_75_581 ();
 sg13g2_decap_4 FILLER_75_595 ();
 sg13g2_fill_2 FILLER_75_599 ();
 sg13g2_decap_4 FILLER_75_618 ();
 sg13g2_fill_1 FILLER_75_622 ();
 sg13g2_decap_4 FILLER_75_642 ();
 sg13g2_fill_1 FILLER_75_659 ();
 sg13g2_fill_1 FILLER_75_664 ();
 sg13g2_decap_4 FILLER_75_696 ();
 sg13g2_decap_4 FILLER_75_705 ();
 sg13g2_fill_1 FILLER_75_709 ();
 sg13g2_fill_2 FILLER_75_715 ();
 sg13g2_fill_1 FILLER_75_722 ();
 sg13g2_fill_2 FILLER_75_784 ();
 sg13g2_fill_1 FILLER_75_812 ();
 sg13g2_fill_1 FILLER_75_826 ();
 sg13g2_fill_2 FILLER_75_840 ();
 sg13g2_fill_1 FILLER_75_847 ();
 sg13g2_fill_2 FILLER_75_856 ();
 sg13g2_decap_8 FILLER_75_871 ();
 sg13g2_fill_2 FILLER_75_878 ();
 sg13g2_decap_8 FILLER_75_893 ();
 sg13g2_decap_8 FILLER_75_900 ();
 sg13g2_decap_8 FILLER_75_907 ();
 sg13g2_fill_2 FILLER_75_914 ();
 sg13g2_fill_1 FILLER_75_916 ();
 sg13g2_fill_1 FILLER_75_939 ();
 sg13g2_fill_1 FILLER_75_945 ();
 sg13g2_fill_1 FILLER_75_958 ();
 sg13g2_fill_1 FILLER_75_980 ();
 sg13g2_fill_1 FILLER_75_986 ();
 sg13g2_decap_8 FILLER_75_992 ();
 sg13g2_fill_1 FILLER_75_1015 ();
 sg13g2_decap_4 FILLER_75_1019 ();
 sg13g2_decap_4 FILLER_75_1031 ();
 sg13g2_fill_2 FILLER_75_1035 ();
 sg13g2_fill_2 FILLER_75_1043 ();
 sg13g2_decap_4 FILLER_75_1059 ();
 sg13g2_decap_8 FILLER_75_1067 ();
 sg13g2_decap_8 FILLER_75_1094 ();
 sg13g2_decap_8 FILLER_75_1101 ();
 sg13g2_decap_8 FILLER_75_1108 ();
 sg13g2_decap_8 FILLER_75_1115 ();
 sg13g2_decap_8 FILLER_75_1122 ();
 sg13g2_decap_8 FILLER_75_1129 ();
 sg13g2_decap_8 FILLER_75_1136 ();
 sg13g2_decap_4 FILLER_75_1147 ();
 sg13g2_fill_2 FILLER_75_1151 ();
 sg13g2_decap_4 FILLER_75_1224 ();
 sg13g2_fill_1 FILLER_75_1228 ();
 sg13g2_fill_1 FILLER_75_1243 ();
 sg13g2_fill_2 FILLER_75_1248 ();
 sg13g2_fill_2 FILLER_75_1255 ();
 sg13g2_fill_1 FILLER_75_1257 ();
 sg13g2_fill_2 FILLER_75_1262 ();
 sg13g2_decap_8 FILLER_75_1277 ();
 sg13g2_fill_2 FILLER_75_1284 ();
 sg13g2_fill_1 FILLER_75_1286 ();
 sg13g2_fill_2 FILLER_75_1290 ();
 sg13g2_fill_1 FILLER_75_1308 ();
 sg13g2_fill_2 FILLER_75_1352 ();
 sg13g2_fill_1 FILLER_75_1354 ();
 sg13g2_fill_2 FILLER_75_1370 ();
 sg13g2_fill_1 FILLER_75_1372 ();
 sg13g2_decap_8 FILLER_75_1377 ();
 sg13g2_decap_8 FILLER_75_1384 ();
 sg13g2_fill_2 FILLER_75_1411 ();
 sg13g2_fill_1 FILLER_75_1413 ();
 sg13g2_fill_2 FILLER_75_1422 ();
 sg13g2_fill_1 FILLER_75_1424 ();
 sg13g2_fill_2 FILLER_75_1462 ();
 sg13g2_fill_1 FILLER_75_1471 ();
 sg13g2_decap_8 FILLER_75_1479 ();
 sg13g2_decap_4 FILLER_75_1486 ();
 sg13g2_fill_2 FILLER_75_1490 ();
 sg13g2_decap_8 FILLER_75_1496 ();
 sg13g2_decap_8 FILLER_75_1503 ();
 sg13g2_decap_8 FILLER_75_1510 ();
 sg13g2_fill_2 FILLER_75_1517 ();
 sg13g2_fill_1 FILLER_75_1519 ();
 sg13g2_fill_2 FILLER_75_1546 ();
 sg13g2_fill_2 FILLER_75_1556 ();
 sg13g2_fill_1 FILLER_75_1558 ();
 sg13g2_fill_2 FILLER_75_1564 ();
 sg13g2_decap_8 FILLER_75_1570 ();
 sg13g2_fill_2 FILLER_75_1577 ();
 sg13g2_fill_1 FILLER_75_1579 ();
 sg13g2_decap_8 FILLER_75_1584 ();
 sg13g2_decap_8 FILLER_75_1591 ();
 sg13g2_decap_8 FILLER_75_1598 ();
 sg13g2_decap_4 FILLER_75_1605 ();
 sg13g2_fill_1 FILLER_75_1645 ();
 sg13g2_decap_8 FILLER_75_1655 ();
 sg13g2_decap_4 FILLER_75_1662 ();
 sg13g2_fill_1 FILLER_75_1666 ();
 sg13g2_fill_2 FILLER_75_1673 ();
 sg13g2_fill_1 FILLER_75_1675 ();
 sg13g2_fill_2 FILLER_75_1688 ();
 sg13g2_fill_1 FILLER_75_1690 ();
 sg13g2_decap_8 FILLER_75_1695 ();
 sg13g2_fill_2 FILLER_75_1702 ();
 sg13g2_fill_1 FILLER_75_1712 ();
 sg13g2_decap_8 FILLER_75_1718 ();
 sg13g2_decap_8 FILLER_75_1725 ();
 sg13g2_decap_8 FILLER_75_1732 ();
 sg13g2_decap_8 FILLER_75_1739 ();
 sg13g2_fill_2 FILLER_75_1746 ();
 sg13g2_fill_1 FILLER_75_1752 ();
 sg13g2_fill_2 FILLER_75_1757 ();
 sg13g2_fill_1 FILLER_75_1759 ();
 sg13g2_decap_8 FILLER_75_1764 ();
 sg13g2_fill_2 FILLER_75_1771 ();
 sg13g2_fill_1 FILLER_75_1773 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_4 FILLER_76_21 ();
 sg13g2_fill_2 FILLER_76_25 ();
 sg13g2_fill_1 FILLER_76_93 ();
 sg13g2_fill_1 FILLER_76_99 ();
 sg13g2_fill_1 FILLER_76_103 ();
 sg13g2_decap_4 FILLER_76_139 ();
 sg13g2_fill_1 FILLER_76_143 ();
 sg13g2_fill_1 FILLER_76_149 ();
 sg13g2_fill_1 FILLER_76_154 ();
 sg13g2_fill_1 FILLER_76_163 ();
 sg13g2_fill_2 FILLER_76_176 ();
 sg13g2_fill_1 FILLER_76_178 ();
 sg13g2_decap_4 FILLER_76_195 ();
 sg13g2_fill_2 FILLER_76_199 ();
 sg13g2_fill_1 FILLER_76_223 ();
 sg13g2_decap_8 FILLER_76_242 ();
 sg13g2_decap_8 FILLER_76_249 ();
 sg13g2_fill_2 FILLER_76_256 ();
 sg13g2_fill_1 FILLER_76_273 ();
 sg13g2_fill_1 FILLER_76_278 ();
 sg13g2_fill_1 FILLER_76_284 ();
 sg13g2_fill_1 FILLER_76_289 ();
 sg13g2_decap_4 FILLER_76_343 ();
 sg13g2_fill_2 FILLER_76_347 ();
 sg13g2_decap_4 FILLER_76_376 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_4 FILLER_76_392 ();
 sg13g2_fill_1 FILLER_76_401 ();
 sg13g2_fill_1 FILLER_76_412 ();
 sg13g2_fill_1 FILLER_76_418 ();
 sg13g2_fill_1 FILLER_76_427 ();
 sg13g2_fill_2 FILLER_76_443 ();
 sg13g2_fill_1 FILLER_76_471 ();
 sg13g2_fill_1 FILLER_76_477 ();
 sg13g2_fill_2 FILLER_76_483 ();
 sg13g2_fill_2 FILLER_76_496 ();
 sg13g2_fill_1 FILLER_76_498 ();
 sg13g2_decap_8 FILLER_76_507 ();
 sg13g2_fill_2 FILLER_76_514 ();
 sg13g2_decap_4 FILLER_76_520 ();
 sg13g2_fill_1 FILLER_76_524 ();
 sg13g2_fill_1 FILLER_76_530 ();
 sg13g2_decap_4 FILLER_76_544 ();
 sg13g2_fill_2 FILLER_76_552 ();
 sg13g2_fill_2 FILLER_76_558 ();
 sg13g2_fill_2 FILLER_76_567 ();
 sg13g2_fill_2 FILLER_76_576 ();
 sg13g2_fill_1 FILLER_76_578 ();
 sg13g2_fill_1 FILLER_76_588 ();
 sg13g2_decap_8 FILLER_76_616 ();
 sg13g2_decap_8 FILLER_76_623 ();
 sg13g2_decap_4 FILLER_76_630 ();
 sg13g2_decap_4 FILLER_76_637 ();
 sg13g2_fill_1 FILLER_76_641 ();
 sg13g2_fill_2 FILLER_76_652 ();
 sg13g2_fill_1 FILLER_76_672 ();
 sg13g2_decap_4 FILLER_76_689 ();
 sg13g2_fill_1 FILLER_76_693 ();
 sg13g2_fill_1 FILLER_76_713 ();
 sg13g2_fill_1 FILLER_76_722 ();
 sg13g2_fill_1 FILLER_76_734 ();
 sg13g2_fill_2 FILLER_76_745 ();
 sg13g2_fill_1 FILLER_76_762 ();
 sg13g2_fill_2 FILLER_76_769 ();
 sg13g2_decap_8 FILLER_76_802 ();
 sg13g2_fill_1 FILLER_76_814 ();
 sg13g2_fill_2 FILLER_76_835 ();
 sg13g2_fill_1 FILLER_76_843 ();
 sg13g2_fill_2 FILLER_76_864 ();
 sg13g2_fill_1 FILLER_76_866 ();
 sg13g2_fill_2 FILLER_76_872 ();
 sg13g2_fill_1 FILLER_76_874 ();
 sg13g2_decap_8 FILLER_76_888 ();
 sg13g2_fill_2 FILLER_76_895 ();
 sg13g2_fill_1 FILLER_76_897 ();
 sg13g2_fill_1 FILLER_76_919 ();
 sg13g2_fill_1 FILLER_76_929 ();
 sg13g2_fill_2 FILLER_76_935 ();
 sg13g2_decap_4 FILLER_76_978 ();
 sg13g2_fill_2 FILLER_76_995 ();
 sg13g2_decap_4 FILLER_76_1002 ();
 sg13g2_fill_2 FILLER_76_1011 ();
 sg13g2_decap_4 FILLER_76_1021 ();
 sg13g2_fill_1 FILLER_76_1030 ();
 sg13g2_decap_8 FILLER_76_1058 ();
 sg13g2_decap_8 FILLER_76_1065 ();
 sg13g2_decap_4 FILLER_76_1072 ();
 sg13g2_fill_1 FILLER_76_1076 ();
 sg13g2_fill_1 FILLER_76_1086 ();
 sg13g2_decap_4 FILLER_76_1103 ();
 sg13g2_fill_2 FILLER_76_1111 ();
 sg13g2_fill_1 FILLER_76_1113 ();
 sg13g2_decap_4 FILLER_76_1122 ();
 sg13g2_fill_1 FILLER_76_1126 ();
 sg13g2_decap_4 FILLER_76_1131 ();
 sg13g2_fill_1 FILLER_76_1135 ();
 sg13g2_decap_8 FILLER_76_1141 ();
 sg13g2_fill_1 FILLER_76_1148 ();
 sg13g2_fill_1 FILLER_76_1189 ();
 sg13g2_fill_1 FILLER_76_1206 ();
 sg13g2_fill_2 FILLER_76_1227 ();
 sg13g2_fill_1 FILLER_76_1229 ();
 sg13g2_fill_1 FILLER_76_1302 ();
 sg13g2_fill_1 FILLER_76_1322 ();
 sg13g2_fill_2 FILLER_76_1348 ();
 sg13g2_fill_1 FILLER_76_1350 ();
 sg13g2_decap_4 FILLER_76_1372 ();
 sg13g2_fill_2 FILLER_76_1381 ();
 sg13g2_fill_1 FILLER_76_1383 ();
 sg13g2_decap_8 FILLER_76_1389 ();
 sg13g2_decap_8 FILLER_76_1401 ();
 sg13g2_decap_8 FILLER_76_1408 ();
 sg13g2_fill_2 FILLER_76_1453 ();
 sg13g2_decap_8 FILLER_76_1460 ();
 sg13g2_decap_8 FILLER_76_1467 ();
 sg13g2_decap_8 FILLER_76_1474 ();
 sg13g2_decap_4 FILLER_76_1481 ();
 sg13g2_fill_2 FILLER_76_1511 ();
 sg13g2_fill_1 FILLER_76_1518 ();
 sg13g2_fill_2 FILLER_76_1544 ();
 sg13g2_fill_1 FILLER_76_1546 ();
 sg13g2_decap_8 FILLER_76_1558 ();
 sg13g2_decap_8 FILLER_76_1599 ();
 sg13g2_decap_8 FILLER_76_1606 ();
 sg13g2_decap_8 FILLER_76_1617 ();
 sg13g2_fill_2 FILLER_76_1624 ();
 sg13g2_fill_1 FILLER_76_1626 ();
 sg13g2_fill_2 FILLER_76_1631 ();
 sg13g2_decap_8 FILLER_76_1650 ();
 sg13g2_decap_8 FILLER_76_1660 ();
 sg13g2_decap_4 FILLER_76_1667 ();
 sg13g2_fill_2 FILLER_76_1677 ();
 sg13g2_decap_4 FILLER_76_1713 ();
 sg13g2_decap_4 FILLER_76_1721 ();
 sg13g2_fill_2 FILLER_76_1725 ();
 sg13g2_fill_2 FILLER_76_1739 ();
 sg13g2_fill_2 FILLER_76_1771 ();
 sg13g2_fill_1 FILLER_76_1773 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_11 ();
 sg13g2_decap_8 FILLER_77_18 ();
 sg13g2_decap_8 FILLER_77_25 ();
 sg13g2_decap_8 FILLER_77_40 ();
 sg13g2_fill_2 FILLER_77_47 ();
 sg13g2_decap_4 FILLER_77_65 ();
 sg13g2_decap_8 FILLER_77_73 ();
 sg13g2_decap_4 FILLER_77_80 ();
 sg13g2_fill_1 FILLER_77_84 ();
 sg13g2_fill_2 FILLER_77_89 ();
 sg13g2_decap_4 FILLER_77_97 ();
 sg13g2_fill_1 FILLER_77_101 ();
 sg13g2_fill_1 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_118 ();
 sg13g2_decap_4 FILLER_77_125 ();
 sg13g2_fill_2 FILLER_77_129 ();
 sg13g2_fill_1 FILLER_77_135 ();
 sg13g2_decap_8 FILLER_77_145 ();
 sg13g2_decap_8 FILLER_77_152 ();
 sg13g2_fill_2 FILLER_77_159 ();
 sg13g2_fill_1 FILLER_77_161 ();
 sg13g2_fill_1 FILLER_77_166 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_fill_1 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_fill_2 FILLER_77_203 ();
 sg13g2_fill_1 FILLER_77_205 ();
 sg13g2_fill_2 FILLER_77_215 ();
 sg13g2_fill_1 FILLER_77_243 ();
 sg13g2_fill_1 FILLER_77_275 ();
 sg13g2_fill_2 FILLER_77_280 ();
 sg13g2_fill_1 FILLER_77_282 ();
 sg13g2_fill_2 FILLER_77_288 ();
 sg13g2_fill_2 FILLER_77_299 ();
 sg13g2_fill_1 FILLER_77_333 ();
 sg13g2_decap_8 FILLER_77_338 ();
 sg13g2_decap_4 FILLER_77_345 ();
 sg13g2_fill_2 FILLER_77_349 ();
 sg13g2_decap_8 FILLER_77_356 ();
 sg13g2_decap_4 FILLER_77_363 ();
 sg13g2_fill_1 FILLER_77_367 ();
 sg13g2_fill_2 FILLER_77_373 ();
 sg13g2_fill_1 FILLER_77_375 ();
 sg13g2_fill_2 FILLER_77_395 ();
 sg13g2_fill_1 FILLER_77_401 ();
 sg13g2_fill_1 FILLER_77_421 ();
 sg13g2_fill_1 FILLER_77_428 ();
 sg13g2_fill_1 FILLER_77_434 ();
 sg13g2_fill_2 FILLER_77_458 ();
 sg13g2_fill_1 FILLER_77_460 ();
 sg13g2_decap_8 FILLER_77_464 ();
 sg13g2_fill_1 FILLER_77_481 ();
 sg13g2_fill_1 FILLER_77_486 ();
 sg13g2_decap_8 FILLER_77_506 ();
 sg13g2_fill_2 FILLER_77_513 ();
 sg13g2_fill_1 FILLER_77_515 ();
 sg13g2_fill_1 FILLER_77_532 ();
 sg13g2_fill_1 FILLER_77_542 ();
 sg13g2_fill_2 FILLER_77_548 ();
 sg13g2_fill_2 FILLER_77_580 ();
 sg13g2_fill_2 FILLER_77_586 ();
 sg13g2_fill_1 FILLER_77_588 ();
 sg13g2_fill_2 FILLER_77_592 ();
 sg13g2_fill_1 FILLER_77_594 ();
 sg13g2_decap_8 FILLER_77_638 ();
 sg13g2_fill_1 FILLER_77_645 ();
 sg13g2_fill_2 FILLER_77_655 ();
 sg13g2_fill_2 FILLER_77_700 ();
 sg13g2_fill_1 FILLER_77_702 ();
 sg13g2_fill_1 FILLER_77_717 ();
 sg13g2_fill_1 FILLER_77_728 ();
 sg13g2_fill_1 FILLER_77_737 ();
 sg13g2_decap_8 FILLER_77_778 ();
 sg13g2_decap_8 FILLER_77_785 ();
 sg13g2_fill_1 FILLER_77_818 ();
 sg13g2_fill_1 FILLER_77_835 ();
 sg13g2_fill_2 FILLER_77_842 ();
 sg13g2_fill_2 FILLER_77_871 ();
 sg13g2_fill_1 FILLER_77_873 ();
 sg13g2_fill_2 FILLER_77_888 ();
 sg13g2_decap_8 FILLER_77_898 ();
 sg13g2_decap_8 FILLER_77_905 ();
 sg13g2_fill_1 FILLER_77_912 ();
 sg13g2_decap_8 FILLER_77_922 ();
 sg13g2_fill_2 FILLER_77_929 ();
 sg13g2_fill_1 FILLER_77_931 ();
 sg13g2_fill_1 FILLER_77_940 ();
 sg13g2_fill_1 FILLER_77_948 ();
 sg13g2_fill_2 FILLER_77_961 ();
 sg13g2_fill_1 FILLER_77_963 ();
 sg13g2_fill_2 FILLER_77_981 ();
 sg13g2_fill_1 FILLER_77_983 ();
 sg13g2_fill_2 FILLER_77_989 ();
 sg13g2_fill_1 FILLER_77_991 ();
 sg13g2_decap_8 FILLER_77_998 ();
 sg13g2_fill_2 FILLER_77_1005 ();
 sg13g2_fill_2 FILLER_77_1014 ();
 sg13g2_fill_1 FILLER_77_1016 ();
 sg13g2_decap_4 FILLER_77_1032 ();
 sg13g2_fill_1 FILLER_77_1036 ();
 sg13g2_fill_1 FILLER_77_1095 ();
 sg13g2_fill_1 FILLER_77_1113 ();
 sg13g2_fill_2 FILLER_77_1150 ();
 sg13g2_fill_1 FILLER_77_1152 ();
 sg13g2_fill_1 FILLER_77_1228 ();
 sg13g2_decap_8 FILLER_77_1232 ();
 sg13g2_fill_2 FILLER_77_1239 ();
 sg13g2_fill_1 FILLER_77_1241 ();
 sg13g2_fill_2 FILLER_77_1247 ();
 sg13g2_fill_1 FILLER_77_1249 ();
 sg13g2_decap_4 FILLER_77_1254 ();
 sg13g2_fill_1 FILLER_77_1258 ();
 sg13g2_fill_1 FILLER_77_1263 ();
 sg13g2_fill_2 FILLER_77_1269 ();
 sg13g2_fill_1 FILLER_77_1271 ();
 sg13g2_fill_2 FILLER_77_1293 ();
 sg13g2_fill_2 FILLER_77_1300 ();
 sg13g2_fill_1 FILLER_77_1319 ();
 sg13g2_fill_1 FILLER_77_1331 ();
 sg13g2_decap_8 FILLER_77_1336 ();
 sg13g2_fill_2 FILLER_77_1343 ();
 sg13g2_fill_1 FILLER_77_1345 ();
 sg13g2_decap_8 FILLER_77_1363 ();
 sg13g2_decap_8 FILLER_77_1370 ();
 sg13g2_fill_2 FILLER_77_1377 ();
 sg13g2_fill_1 FILLER_77_1379 ();
 sg13g2_decap_4 FILLER_77_1406 ();
 sg13g2_fill_1 FILLER_77_1410 ();
 sg13g2_fill_2 FILLER_77_1428 ();
 sg13g2_fill_2 FILLER_77_1434 ();
 sg13g2_decap_4 FILLER_77_1445 ();
 sg13g2_decap_8 FILLER_77_1453 ();
 sg13g2_decap_8 FILLER_77_1460 ();
 sg13g2_decap_8 FILLER_77_1467 ();
 sg13g2_decap_8 FILLER_77_1474 ();
 sg13g2_decap_8 FILLER_77_1481 ();
 sg13g2_decap_8 FILLER_77_1488 ();
 sg13g2_decap_8 FILLER_77_1495 ();
 sg13g2_decap_8 FILLER_77_1506 ();
 sg13g2_fill_2 FILLER_77_1513 ();
 sg13g2_fill_1 FILLER_77_1515 ();
 sg13g2_fill_2 FILLER_77_1532 ();
 sg13g2_fill_2 FILLER_77_1539 ();
 sg13g2_decap_8 FILLER_77_1552 ();
 sg13g2_fill_2 FILLER_77_1559 ();
 sg13g2_fill_1 FILLER_77_1561 ();
 sg13g2_fill_2 FILLER_77_1570 ();
 sg13g2_fill_1 FILLER_77_1572 ();
 sg13g2_fill_1 FILLER_77_1593 ();
 sg13g2_decap_8 FILLER_77_1611 ();
 sg13g2_decap_8 FILLER_77_1618 ();
 sg13g2_decap_4 FILLER_77_1625 ();
 sg13g2_fill_1 FILLER_77_1629 ();
 sg13g2_fill_2 FILLER_77_1634 ();
 sg13g2_fill_1 FILLER_77_1636 ();
 sg13g2_fill_1 FILLER_77_1641 ();
 sg13g2_fill_2 FILLER_77_1674 ();
 sg13g2_fill_1 FILLER_77_1676 ();
 sg13g2_decap_8 FILLER_77_1681 ();
 sg13g2_decap_4 FILLER_77_1688 ();
 sg13g2_decap_4 FILLER_77_1701 ();
 sg13g2_fill_1 FILLER_77_1705 ();
 sg13g2_fill_2 FILLER_77_1742 ();
 sg13g2_decap_4 FILLER_77_1770 ();
 sg13g2_fill_1 FILLER_78_26 ();
 sg13g2_decap_8 FILLER_78_40 ();
 sg13g2_decap_8 FILLER_78_47 ();
 sg13g2_decap_8 FILLER_78_54 ();
 sg13g2_decap_8 FILLER_78_96 ();
 sg13g2_fill_1 FILLER_78_123 ();
 sg13g2_fill_1 FILLER_78_128 ();
 sg13g2_fill_1 FILLER_78_134 ();
 sg13g2_fill_2 FILLER_78_140 ();
 sg13g2_decap_4 FILLER_78_178 ();
 sg13g2_fill_2 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_193 ();
 sg13g2_decap_4 FILLER_78_200 ();
 sg13g2_decap_4 FILLER_78_219 ();
 sg13g2_fill_2 FILLER_78_223 ();
 sg13g2_decap_4 FILLER_78_229 ();
 sg13g2_decap_4 FILLER_78_242 ();
 sg13g2_fill_2 FILLER_78_246 ();
 sg13g2_fill_2 FILLER_78_255 ();
 sg13g2_fill_1 FILLER_78_266 ();
 sg13g2_decap_4 FILLER_78_271 ();
 sg13g2_fill_2 FILLER_78_275 ();
 sg13g2_fill_1 FILLER_78_287 ();
 sg13g2_fill_1 FILLER_78_292 ();
 sg13g2_decap_8 FILLER_78_335 ();
 sg13g2_fill_2 FILLER_78_342 ();
 sg13g2_fill_1 FILLER_78_344 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_4 FILLER_78_357 ();
 sg13g2_fill_2 FILLER_78_361 ();
 sg13g2_decap_8 FILLER_78_368 ();
 sg13g2_fill_1 FILLER_78_375 ();
 sg13g2_fill_2 FILLER_78_380 ();
 sg13g2_fill_1 FILLER_78_391 ();
 sg13g2_decap_4 FILLER_78_400 ();
 sg13g2_fill_2 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_422 ();
 sg13g2_fill_1 FILLER_78_428 ();
 sg13g2_fill_1 FILLER_78_433 ();
 sg13g2_decap_4 FILLER_78_437 ();
 sg13g2_fill_1 FILLER_78_445 ();
 sg13g2_fill_1 FILLER_78_451 ();
 sg13g2_fill_1 FILLER_78_461 ();
 sg13g2_fill_2 FILLER_78_468 ();
 sg13g2_fill_1 FILLER_78_474 ();
 sg13g2_fill_2 FILLER_78_480 ();
 sg13g2_fill_2 FILLER_78_497 ();
 sg13g2_fill_1 FILLER_78_499 ();
 sg13g2_fill_1 FILLER_78_508 ();
 sg13g2_decap_8 FILLER_78_514 ();
 sg13g2_decap_4 FILLER_78_521 ();
 sg13g2_fill_2 FILLER_78_530 ();
 sg13g2_decap_8 FILLER_78_542 ();
 sg13g2_decap_8 FILLER_78_577 ();
 sg13g2_decap_8 FILLER_78_584 ();
 sg13g2_decap_8 FILLER_78_591 ();
 sg13g2_decap_8 FILLER_78_598 ();
 sg13g2_fill_2 FILLER_78_605 ();
 sg13g2_fill_1 FILLER_78_607 ();
 sg13g2_fill_2 FILLER_78_613 ();
 sg13g2_decap_8 FILLER_78_620 ();
 sg13g2_fill_2 FILLER_78_627 ();
 sg13g2_decap_4 FILLER_78_633 ();
 sg13g2_fill_1 FILLER_78_637 ();
 sg13g2_decap_4 FILLER_78_686 ();
 sg13g2_fill_2 FILLER_78_690 ();
 sg13g2_fill_1 FILLER_78_706 ();
 sg13g2_fill_2 FILLER_78_715 ();
 sg13g2_fill_1 FILLER_78_722 ();
 sg13g2_fill_1 FILLER_78_735 ();
 sg13g2_decap_4 FILLER_78_778 ();
 sg13g2_fill_2 FILLER_78_782 ();
 sg13g2_fill_2 FILLER_78_817 ();
 sg13g2_fill_2 FILLER_78_840 ();
 sg13g2_fill_1 FILLER_78_850 ();
 sg13g2_fill_1 FILLER_78_862 ();
 sg13g2_fill_2 FILLER_78_884 ();
 sg13g2_decap_8 FILLER_78_894 ();
 sg13g2_fill_2 FILLER_78_901 ();
 sg13g2_fill_1 FILLER_78_903 ();
 sg13g2_fill_2 FILLER_78_908 ();
 sg13g2_decap_4 FILLER_78_914 ();
 sg13g2_fill_2 FILLER_78_918 ();
 sg13g2_fill_1 FILLER_78_924 ();
 sg13g2_fill_2 FILLER_78_930 ();
 sg13g2_decap_4 FILLER_78_937 ();
 sg13g2_fill_1 FILLER_78_941 ();
 sg13g2_decap_4 FILLER_78_965 ();
 sg13g2_decap_8 FILLER_78_974 ();
 sg13g2_decap_8 FILLER_78_981 ();
 sg13g2_decap_8 FILLER_78_988 ();
 sg13g2_decap_8 FILLER_78_995 ();
 sg13g2_fill_2 FILLER_78_1002 ();
 sg13g2_decap_8 FILLER_78_1017 ();
 sg13g2_decap_4 FILLER_78_1024 ();
 sg13g2_fill_1 FILLER_78_1044 ();
 sg13g2_decap_4 FILLER_78_1049 ();
 sg13g2_fill_2 FILLER_78_1053 ();
 sg13g2_fill_2 FILLER_78_1061 ();
 sg13g2_fill_2 FILLER_78_1068 ();
 sg13g2_fill_1 FILLER_78_1070 ();
 sg13g2_fill_2 FILLER_78_1084 ();
 sg13g2_fill_2 FILLER_78_1115 ();
 sg13g2_fill_1 FILLER_78_1117 ();
 sg13g2_decap_8 FILLER_78_1123 ();
 sg13g2_fill_2 FILLER_78_1130 ();
 sg13g2_decap_4 FILLER_78_1136 ();
 sg13g2_fill_2 FILLER_78_1143 ();
 sg13g2_fill_1 FILLER_78_1156 ();
 sg13g2_fill_2 FILLER_78_1166 ();
 sg13g2_fill_1 FILLER_78_1184 ();
 sg13g2_decap_8 FILLER_78_1188 ();
 sg13g2_fill_2 FILLER_78_1195 ();
 sg13g2_decap_8 FILLER_78_1205 ();
 sg13g2_decap_8 FILLER_78_1212 ();
 sg13g2_decap_8 FILLER_78_1253 ();
 sg13g2_decap_8 FILLER_78_1260 ();
 sg13g2_fill_2 FILLER_78_1267 ();
 sg13g2_fill_1 FILLER_78_1269 ();
 sg13g2_fill_2 FILLER_78_1294 ();
 sg13g2_fill_2 FILLER_78_1314 ();
 sg13g2_fill_2 FILLER_78_1324 ();
 sg13g2_decap_8 FILLER_78_1334 ();
 sg13g2_decap_8 FILLER_78_1341 ();
 sg13g2_decap_8 FILLER_78_1348 ();
 sg13g2_decap_8 FILLER_78_1355 ();
 sg13g2_decap_8 FILLER_78_1362 ();
 sg13g2_decap_8 FILLER_78_1369 ();
 sg13g2_decap_8 FILLER_78_1376 ();
 sg13g2_fill_2 FILLER_78_1383 ();
 sg13g2_decap_8 FILLER_78_1389 ();
 sg13g2_decap_8 FILLER_78_1396 ();
 sg13g2_decap_8 FILLER_78_1403 ();
 sg13g2_decap_8 FILLER_78_1410 ();
 sg13g2_decap_8 FILLER_78_1417 ();
 sg13g2_fill_1 FILLER_78_1424 ();
 sg13g2_decap_8 FILLER_78_1428 ();
 sg13g2_decap_8 FILLER_78_1435 ();
 sg13g2_decap_8 FILLER_78_1442 ();
 sg13g2_decap_8 FILLER_78_1449 ();
 sg13g2_decap_8 FILLER_78_1456 ();
 sg13g2_decap_8 FILLER_78_1463 ();
 sg13g2_decap_4 FILLER_78_1470 ();
 sg13g2_fill_1 FILLER_78_1474 ();
 sg13g2_fill_1 FILLER_78_1501 ();
 sg13g2_fill_1 FILLER_78_1506 ();
 sg13g2_decap_4 FILLER_78_1519 ();
 sg13g2_decap_8 FILLER_78_1545 ();
 sg13g2_decap_8 FILLER_78_1552 ();
 sg13g2_decap_4 FILLER_78_1559 ();
 sg13g2_fill_1 FILLER_78_1563 ();
 sg13g2_decap_4 FILLER_78_1581 ();
 sg13g2_fill_2 FILLER_78_1585 ();
 sg13g2_fill_2 FILLER_78_1617 ();
 sg13g2_fill_1 FILLER_78_1619 ();
 sg13g2_fill_2 FILLER_78_1650 ();
 sg13g2_fill_1 FILLER_78_1652 ();
 sg13g2_decap_8 FILLER_78_1657 ();
 sg13g2_decap_8 FILLER_78_1664 ();
 sg13g2_decap_8 FILLER_78_1671 ();
 sg13g2_decap_4 FILLER_78_1678 ();
 sg13g2_fill_2 FILLER_78_1682 ();
 sg13g2_decap_8 FILLER_78_1689 ();
 sg13g2_decap_8 FILLER_78_1696 ();
 sg13g2_decap_4 FILLER_78_1703 ();
 sg13g2_fill_2 FILLER_78_1715 ();
 sg13g2_decap_4 FILLER_78_1721 ();
 sg13g2_fill_2 FILLER_78_1749 ();
 sg13g2_fill_1 FILLER_78_1751 ();
 sg13g2_fill_2 FILLER_78_1756 ();
 sg13g2_fill_1 FILLER_78_1758 ();
 sg13g2_decap_8 FILLER_78_1763 ();
 sg13g2_decap_4 FILLER_78_1770 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_38 ();
 sg13g2_fill_2 FILLER_79_45 ();
 sg13g2_fill_1 FILLER_79_47 ();
 sg13g2_decap_8 FILLER_79_52 ();
 sg13g2_fill_1 FILLER_79_59 ();
 sg13g2_fill_2 FILLER_79_73 ();
 sg13g2_fill_1 FILLER_79_100 ();
 sg13g2_decap_4 FILLER_79_105 ();
 sg13g2_fill_2 FILLER_79_109 ();
 sg13g2_fill_2 FILLER_79_141 ();
 sg13g2_fill_1 FILLER_79_143 ();
 sg13g2_decap_8 FILLER_79_148 ();
 sg13g2_decap_4 FILLER_79_155 ();
 sg13g2_decap_8 FILLER_79_163 ();
 sg13g2_decap_8 FILLER_79_170 ();
 sg13g2_fill_2 FILLER_79_177 ();
 sg13g2_fill_1 FILLER_79_179 ();
 sg13g2_fill_1 FILLER_79_240 ();
 sg13g2_fill_2 FILLER_79_252 ();
 sg13g2_fill_2 FILLER_79_266 ();
 sg13g2_decap_4 FILLER_79_277 ();
 sg13g2_fill_2 FILLER_79_307 ();
 sg13g2_fill_2 FILLER_79_312 ();
 sg13g2_decap_8 FILLER_79_318 ();
 sg13g2_fill_2 FILLER_79_325 ();
 sg13g2_decap_8 FILLER_79_331 ();
 sg13g2_decap_4 FILLER_79_338 ();
 sg13g2_fill_1 FILLER_79_342 ();
 sg13g2_decap_4 FILLER_79_348 ();
 sg13g2_decap_4 FILLER_79_357 ();
 sg13g2_fill_1 FILLER_79_361 ();
 sg13g2_decap_4 FILLER_79_388 ();
 sg13g2_decap_4 FILLER_79_400 ();
 sg13g2_fill_1 FILLER_79_404 ();
 sg13g2_fill_2 FILLER_79_410 ();
 sg13g2_fill_2 FILLER_79_417 ();
 sg13g2_decap_4 FILLER_79_423 ();
 sg13g2_fill_2 FILLER_79_462 ();
 sg13g2_fill_1 FILLER_79_464 ();
 sg13g2_fill_2 FILLER_79_469 ();
 sg13g2_fill_2 FILLER_79_476 ();
 sg13g2_fill_1 FILLER_79_478 ();
 sg13g2_fill_1 FILLER_79_484 ();
 sg13g2_fill_1 FILLER_79_490 ();
 sg13g2_fill_1 FILLER_79_495 ();
 sg13g2_fill_2 FILLER_79_501 ();
 sg13g2_fill_2 FILLER_79_508 ();
 sg13g2_fill_2 FILLER_79_519 ();
 sg13g2_fill_1 FILLER_79_521 ();
 sg13g2_decap_8 FILLER_79_537 ();
 sg13g2_decap_8 FILLER_79_544 ();
 sg13g2_fill_2 FILLER_79_551 ();
 sg13g2_fill_2 FILLER_79_563 ();
 sg13g2_fill_1 FILLER_79_573 ();
 sg13g2_fill_1 FILLER_79_587 ();
 sg13g2_decap_4 FILLER_79_627 ();
 sg13g2_fill_1 FILLER_79_657 ();
 sg13g2_fill_1 FILLER_79_662 ();
 sg13g2_fill_2 FILLER_79_668 ();
 sg13g2_fill_1 FILLER_79_696 ();
 sg13g2_fill_1 FILLER_79_702 ();
 sg13g2_decap_8 FILLER_79_740 ();
 sg13g2_decap_8 FILLER_79_747 ();
 sg13g2_decap_8 FILLER_79_754 ();
 sg13g2_decap_8 FILLER_79_761 ();
 sg13g2_decap_4 FILLER_79_768 ();
 sg13g2_fill_2 FILLER_79_772 ();
 sg13g2_decap_4 FILLER_79_783 ();
 sg13g2_fill_1 FILLER_79_787 ();
 sg13g2_fill_1 FILLER_79_807 ();
 sg13g2_fill_1 FILLER_79_841 ();
 sg13g2_fill_1 FILLER_79_847 ();
 sg13g2_fill_1 FILLER_79_855 ();
 sg13g2_decap_4 FILLER_79_866 ();
 sg13g2_fill_1 FILLER_79_870 ();
 sg13g2_fill_2 FILLER_79_912 ();
 sg13g2_fill_1 FILLER_79_914 ();
 sg13g2_fill_1 FILLER_79_954 ();
 sg13g2_decap_8 FILLER_79_1013 ();
 sg13g2_fill_1 FILLER_79_1020 ();
 sg13g2_fill_1 FILLER_79_1051 ();
 sg13g2_fill_2 FILLER_79_1066 ();
 sg13g2_fill_2 FILLER_79_1083 ();
 sg13g2_fill_1 FILLER_79_1085 ();
 sg13g2_decap_8 FILLER_79_1090 ();
 sg13g2_fill_2 FILLER_79_1097 ();
 sg13g2_decap_8 FILLER_79_1125 ();
 sg13g2_decap_4 FILLER_79_1132 ();
 sg13g2_fill_2 FILLER_79_1136 ();
 sg13g2_fill_1 FILLER_79_1173 ();
 sg13g2_decap_8 FILLER_79_1197 ();
 sg13g2_fill_2 FILLER_79_1204 ();
 sg13g2_fill_1 FILLER_79_1206 ();
 sg13g2_decap_8 FILLER_79_1211 ();
 sg13g2_fill_1 FILLER_79_1218 ();
 sg13g2_decap_8 FILLER_79_1224 ();
 sg13g2_decap_8 FILLER_79_1231 ();
 sg13g2_decap_8 FILLER_79_1238 ();
 sg13g2_decap_8 FILLER_79_1245 ();
 sg13g2_decap_8 FILLER_79_1326 ();
 sg13g2_decap_8 FILLER_79_1333 ();
 sg13g2_decap_8 FILLER_79_1340 ();
 sg13g2_decap_8 FILLER_79_1347 ();
 sg13g2_decap_8 FILLER_79_1354 ();
 sg13g2_decap_8 FILLER_79_1361 ();
 sg13g2_decap_8 FILLER_79_1368 ();
 sg13g2_decap_8 FILLER_79_1375 ();
 sg13g2_decap_8 FILLER_79_1382 ();
 sg13g2_decap_8 FILLER_79_1389 ();
 sg13g2_decap_8 FILLER_79_1396 ();
 sg13g2_decap_8 FILLER_79_1403 ();
 sg13g2_decap_8 FILLER_79_1413 ();
 sg13g2_decap_8 FILLER_79_1420 ();
 sg13g2_decap_8 FILLER_79_1427 ();
 sg13g2_decap_8 FILLER_79_1434 ();
 sg13g2_decap_8 FILLER_79_1441 ();
 sg13g2_decap_8 FILLER_79_1448 ();
 sg13g2_decap_8 FILLER_79_1455 ();
 sg13g2_decap_8 FILLER_79_1462 ();
 sg13g2_decap_8 FILLER_79_1469 ();
 sg13g2_decap_8 FILLER_79_1476 ();
 sg13g2_decap_4 FILLER_79_1487 ();
 sg13g2_fill_1 FILLER_79_1491 ();
 sg13g2_decap_8 FILLER_79_1496 ();
 sg13g2_fill_2 FILLER_79_1503 ();
 sg13g2_fill_1 FILLER_79_1505 ();
 sg13g2_fill_2 FILLER_79_1523 ();
 sg13g2_decap_4 FILLER_79_1534 ();
 sg13g2_fill_2 FILLER_79_1550 ();
 sg13g2_fill_1 FILLER_79_1552 ();
 sg13g2_decap_8 FILLER_79_1557 ();
 sg13g2_decap_4 FILLER_79_1568 ();
 sg13g2_fill_1 FILLER_79_1572 ();
 sg13g2_decap_4 FILLER_79_1585 ();
 sg13g2_decap_8 FILLER_79_1593 ();
 sg13g2_decap_8 FILLER_79_1600 ();
 sg13g2_decap_4 FILLER_79_1607 ();
 sg13g2_decap_8 FILLER_79_1628 ();
 sg13g2_decap_8 FILLER_79_1635 ();
 sg13g2_decap_4 FILLER_79_1642 ();
 sg13g2_decap_8 FILLER_79_1700 ();
 sg13g2_decap_4 FILLER_79_1707 ();
 sg13g2_fill_1 FILLER_79_1711 ();
 sg13g2_decap_8 FILLER_79_1725 ();
 sg13g2_fill_1 FILLER_79_1732 ();
 sg13g2_fill_1 FILLER_79_1737 ();
 sg13g2_decap_8 FILLER_79_1764 ();
 sg13g2_fill_2 FILLER_79_1771 ();
 sg13g2_fill_1 FILLER_79_1773 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_4 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_51 ();
 sg13g2_fill_2 FILLER_80_58 ();
 sg13g2_fill_2 FILLER_80_90 ();
 sg13g2_fill_1 FILLER_80_104 ();
 sg13g2_fill_1 FILLER_80_117 ();
 sg13g2_fill_1 FILLER_80_198 ();
 sg13g2_fill_2 FILLER_80_216 ();
 sg13g2_decap_4 FILLER_80_258 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_284 ();
 sg13g2_decap_4 FILLER_80_291 ();
 sg13g2_decap_8 FILLER_80_302 ();
 sg13g2_decap_4 FILLER_80_309 ();
 sg13g2_fill_2 FILLER_80_313 ();
 sg13g2_decap_4 FILLER_80_319 ();
 sg13g2_fill_1 FILLER_80_323 ();
 sg13g2_fill_2 FILLER_80_345 ();
 sg13g2_fill_1 FILLER_80_347 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_2 FILLER_80_367 ();
 sg13g2_fill_1 FILLER_80_369 ();
 sg13g2_fill_2 FILLER_80_378 ();
 sg13g2_decap_8 FILLER_80_424 ();
 sg13g2_fill_1 FILLER_80_431 ();
 sg13g2_decap_4 FILLER_80_436 ();
 sg13g2_fill_1 FILLER_80_450 ();
 sg13g2_decap_8 FILLER_80_456 ();
 sg13g2_decap_4 FILLER_80_463 ();
 sg13g2_fill_2 FILLER_80_467 ();
 sg13g2_decap_4 FILLER_80_474 ();
 sg13g2_fill_1 FILLER_80_478 ();
 sg13g2_decap_4 FILLER_80_494 ();
 sg13g2_fill_2 FILLER_80_498 ();
 sg13g2_fill_1 FILLER_80_505 ();
 sg13g2_fill_2 FILLER_80_510 ();
 sg13g2_fill_2 FILLER_80_520 ();
 sg13g2_fill_1 FILLER_80_522 ();
 sg13g2_fill_2 FILLER_80_535 ();
 sg13g2_fill_2 FILLER_80_547 ();
 sg13g2_fill_1 FILLER_80_553 ();
 sg13g2_decap_4 FILLER_80_559 ();
 sg13g2_fill_2 FILLER_80_563 ();
 sg13g2_decap_4 FILLER_80_569 ();
 sg13g2_decap_8 FILLER_80_578 ();
 sg13g2_decap_8 FILLER_80_585 ();
 sg13g2_fill_2 FILLER_80_592 ();
 sg13g2_decap_4 FILLER_80_602 ();
 sg13g2_decap_8 FILLER_80_617 ();
 sg13g2_decap_8 FILLER_80_624 ();
 sg13g2_decap_8 FILLER_80_631 ();
 sg13g2_fill_2 FILLER_80_638 ();
 sg13g2_decap_8 FILLER_80_644 ();
 sg13g2_fill_1 FILLER_80_651 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_4 FILLER_80_662 ();
 sg13g2_decap_4 FILLER_80_670 ();
 sg13g2_fill_1 FILLER_80_681 ();
 sg13g2_fill_2 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_733 ();
 sg13g2_decap_8 FILLER_80_740 ();
 sg13g2_decap_8 FILLER_80_747 ();
 sg13g2_decap_8 FILLER_80_754 ();
 sg13g2_decap_8 FILLER_80_761 ();
 sg13g2_decap_8 FILLER_80_768 ();
 sg13g2_decap_8 FILLER_80_775 ();
 sg13g2_decap_8 FILLER_80_782 ();
 sg13g2_decap_8 FILLER_80_789 ();
 sg13g2_decap_8 FILLER_80_796 ();
 sg13g2_decap_8 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_810 ();
 sg13g2_fill_2 FILLER_80_817 ();
 sg13g2_fill_2 FILLER_80_823 ();
 sg13g2_fill_1 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_830 ();
 sg13g2_decap_4 FILLER_80_837 ();
 sg13g2_decap_4 FILLER_80_867 ();
 sg13g2_decap_4 FILLER_80_891 ();
 sg13g2_fill_2 FILLER_80_900 ();
 sg13g2_fill_1 FILLER_80_902 ();
 sg13g2_decap_8 FILLER_80_907 ();
 sg13g2_decap_8 FILLER_80_914 ();
 sg13g2_decap_8 FILLER_80_921 ();
 sg13g2_decap_8 FILLER_80_928 ();
 sg13g2_decap_8 FILLER_80_935 ();
 sg13g2_decap_4 FILLER_80_942 ();
 sg13g2_fill_1 FILLER_80_946 ();
 sg13g2_decap_8 FILLER_80_952 ();
 sg13g2_decap_4 FILLER_80_959 ();
 sg13g2_fill_1 FILLER_80_963 ();
 sg13g2_decap_8 FILLER_80_973 ();
 sg13g2_decap_8 FILLER_80_980 ();
 sg13g2_fill_2 FILLER_80_987 ();
 sg13g2_fill_1 FILLER_80_989 ();
 sg13g2_decap_8 FILLER_80_994 ();
 sg13g2_decap_8 FILLER_80_1001 ();
 sg13g2_decap_4 FILLER_80_1008 ();
 sg13g2_fill_2 FILLER_80_1012 ();
 sg13g2_fill_2 FILLER_80_1049 ();
 sg13g2_fill_1 FILLER_80_1051 ();
 sg13g2_fill_2 FILLER_80_1062 ();
 sg13g2_decap_8 FILLER_80_1077 ();
 sg13g2_decap_8 FILLER_80_1084 ();
 sg13g2_decap_8 FILLER_80_1091 ();
 sg13g2_decap_8 FILLER_80_1098 ();
 sg13g2_fill_1 FILLER_80_1105 ();
 sg13g2_decap_8 FILLER_80_1110 ();
 sg13g2_decap_8 FILLER_80_1117 ();
 sg13g2_decap_8 FILLER_80_1124 ();
 sg13g2_decap_8 FILLER_80_1131 ();
 sg13g2_decap_8 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_decap_8 FILLER_80_1152 ();
 sg13g2_decap_8 FILLER_80_1159 ();
 sg13g2_fill_2 FILLER_80_1166 ();
 sg13g2_fill_1 FILLER_80_1168 ();
 sg13g2_fill_1 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_decap_8 FILLER_80_1186 ();
 sg13g2_decap_4 FILLER_80_1193 ();
 sg13g2_fill_2 FILLER_80_1197 ();
 sg13g2_decap_8 FILLER_80_1225 ();
 sg13g2_decap_8 FILLER_80_1232 ();
 sg13g2_decap_8 FILLER_80_1239 ();
 sg13g2_fill_1 FILLER_80_1286 ();
 sg13g2_decap_8 FILLER_80_1322 ();
 sg13g2_fill_2 FILLER_80_1329 ();
 sg13g2_decap_8 FILLER_80_1336 ();
 sg13g2_decap_8 FILLER_80_1343 ();
 sg13g2_decap_8 FILLER_80_1350 ();
 sg13g2_decap_8 FILLER_80_1357 ();
 sg13g2_decap_8 FILLER_80_1364 ();
 sg13g2_decap_8 FILLER_80_1371 ();
 sg13g2_decap_8 FILLER_80_1378 ();
 sg13g2_decap_8 FILLER_80_1385 ();
 sg13g2_decap_8 FILLER_80_1392 ();
 sg13g2_decap_8 FILLER_80_1399 ();
 sg13g2_decap_8 FILLER_80_1406 ();
 sg13g2_decap_8 FILLER_80_1413 ();
 sg13g2_decap_8 FILLER_80_1420 ();
 sg13g2_decap_8 FILLER_80_1427 ();
 sg13g2_decap_8 FILLER_80_1434 ();
 sg13g2_decap_8 FILLER_80_1441 ();
 sg13g2_decap_8 FILLER_80_1448 ();
 sg13g2_decap_8 FILLER_80_1455 ();
 sg13g2_decap_8 FILLER_80_1462 ();
 sg13g2_decap_8 FILLER_80_1469 ();
 sg13g2_decap_8 FILLER_80_1476 ();
 sg13g2_fill_2 FILLER_80_1483 ();
 sg13g2_decap_8 FILLER_80_1511 ();
 sg13g2_decap_8 FILLER_80_1518 ();
 sg13g2_decap_8 FILLER_80_1525 ();
 sg13g2_decap_8 FILLER_80_1532 ();
 sg13g2_fill_2 FILLER_80_1539 ();
 sg13g2_fill_1 FILLER_80_1541 ();
 sg13g2_decap_8 FILLER_80_1568 ();
 sg13g2_decap_8 FILLER_80_1575 ();
 sg13g2_decap_8 FILLER_80_1608 ();
 sg13g2_decap_8 FILLER_80_1615 ();
 sg13g2_decap_8 FILLER_80_1622 ();
 sg13g2_decap_8 FILLER_80_1629 ();
 sg13g2_decap_8 FILLER_80_1636 ();
 sg13g2_decap_8 FILLER_80_1643 ();
 sg13g2_decap_8 FILLER_80_1650 ();
 sg13g2_fill_1 FILLER_80_1657 ();
 sg13g2_decap_8 FILLER_80_1662 ();
 sg13g2_decap_8 FILLER_80_1669 ();
 sg13g2_fill_2 FILLER_80_1676 ();
 sg13g2_fill_2 FILLER_80_1682 ();
 sg13g2_fill_1 FILLER_80_1684 ();
 sg13g2_fill_2 FILLER_80_1711 ();
 sg13g2_fill_1 FILLER_80_1713 ();
 sg13g2_decap_8 FILLER_80_1740 ();
 sg13g2_decap_8 FILLER_80_1747 ();
 sg13g2_decap_8 FILLER_80_1754 ();
 sg13g2_decap_8 FILLER_80_1761 ();
 sg13g2_decap_4 FILLER_80_1768 ();
 sg13g2_fill_2 FILLER_80_1772 ();
endmodule
