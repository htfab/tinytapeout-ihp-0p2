module tt_um_devinatkin_pulse_width_counter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire clknet_0_clk;
 wire net80;
 wire \mux.data_in[0] ;
 wire \mux.data_in[10] ;
 wire \mux.data_in[11] ;
 wire \mux.data_in[12] ;
 wire \mux.data_in[13] ;
 wire \mux.data_in[14] ;
 wire \mux.data_in[15] ;
 wire \mux.data_in[16] ;
 wire \mux.data_in[17] ;
 wire \mux.data_in[18] ;
 wire \mux.data_in[19] ;
 wire \mux.data_in[1] ;
 wire \mux.data_in[20] ;
 wire \mux.data_in[21] ;
 wire \mux.data_in[22] ;
 wire \mux.data_in[23] ;
 wire \mux.data_in[24] ;
 wire \mux.data_in[25] ;
 wire \mux.data_in[26] ;
 wire \mux.data_in[27] ;
 wire \mux.data_in[28] ;
 wire \mux.data_in[29] ;
 wire \mux.data_in[2] ;
 wire \mux.data_in[30] ;
 wire \mux.data_in[31] ;
 wire \mux.data_in[32] ;
 wire \mux.data_in[33] ;
 wire \mux.data_in[34] ;
 wire \mux.data_in[35] ;
 wire \mux.data_in[36] ;
 wire \mux.data_in[37] ;
 wire \mux.data_in[38] ;
 wire \mux.data_in[39] ;
 wire \mux.data_in[3] ;
 wire \mux.data_in[40] ;
 wire \mux.data_in[41] ;
 wire \mux.data_in[42] ;
 wire \mux.data_in[43] ;
 wire \mux.data_in[44] ;
 wire \mux.data_in[45] ;
 wire \mux.data_in[46] ;
 wire \mux.data_in[47] ;
 wire \mux.data_in[48] ;
 wire \mux.data_in[49] ;
 wire \mux.data_in[4] ;
 wire \mux.data_in[50] ;
 wire \mux.data_in[51] ;
 wire \mux.data_in[52] ;
 wire \mux.data_in[53] ;
 wire \mux.data_in[54] ;
 wire \mux.data_in[55] ;
 wire \mux.data_in[56] ;
 wire \mux.data_in[57] ;
 wire \mux.data_in[58] ;
 wire \mux.data_in[59] ;
 wire \mux.data_in[5] ;
 wire \mux.data_in[60] ;
 wire \mux.data_in[61] ;
 wire \mux.data_in[62] ;
 wire \mux.data_in[63] ;
 wire \mux.data_in[64] ;
 wire \mux.data_in[65] ;
 wire \mux.data_in[66] ;
 wire \mux.data_in[67] ;
 wire \mux.data_in[68] ;
 wire \mux.data_in[69] ;
 wire \mux.data_in[6] ;
 wire \mux.data_in[70] ;
 wire \mux.data_in[71] ;
 wire \mux.data_in[72] ;
 wire \mux.data_in[73] ;
 wire \mux.data_in[74] ;
 wire \mux.data_in[75] ;
 wire \mux.data_in[76] ;
 wire \mux.data_in[77] ;
 wire \mux.data_in[78] ;
 wire \mux.data_in[79] ;
 wire \mux.data_in[7] ;
 wire \mux.data_in[80] ;
 wire \mux.data_in[81] ;
 wire \mux.data_in[82] ;
 wire \mux.data_in[83] ;
 wire \mux.data_in[84] ;
 wire \mux.data_in[85] ;
 wire \mux.data_in[86] ;
 wire \mux.data_in[87] ;
 wire \mux.data_in[88] ;
 wire \mux.data_in[89] ;
 wire \mux.data_in[8] ;
 wire \mux.data_in[90] ;
 wire \mux.data_in[91] ;
 wire \mux.data_in[92] ;
 wire \mux.data_in[93] ;
 wire \mux.data_in[94] ;
 wire \mux.data_in[95] ;
 wire \mux.data_in[9] ;
 wire \pulse_width_counter_module.high_counter[0] ;
 wire \pulse_width_counter_module.high_counter[10] ;
 wire \pulse_width_counter_module.high_counter[11] ;
 wire \pulse_width_counter_module.high_counter[12] ;
 wire \pulse_width_counter_module.high_counter[13] ;
 wire \pulse_width_counter_module.high_counter[14] ;
 wire \pulse_width_counter_module.high_counter[15] ;
 wire \pulse_width_counter_module.high_counter[16] ;
 wire \pulse_width_counter_module.high_counter[17] ;
 wire \pulse_width_counter_module.high_counter[18] ;
 wire \pulse_width_counter_module.high_counter[19] ;
 wire \pulse_width_counter_module.high_counter[1] ;
 wire \pulse_width_counter_module.high_counter[20] ;
 wire \pulse_width_counter_module.high_counter[21] ;
 wire \pulse_width_counter_module.high_counter[22] ;
 wire \pulse_width_counter_module.high_counter[23] ;
 wire \pulse_width_counter_module.high_counter[24] ;
 wire \pulse_width_counter_module.high_counter[25] ;
 wire \pulse_width_counter_module.high_counter[26] ;
 wire \pulse_width_counter_module.high_counter[27] ;
 wire \pulse_width_counter_module.high_counter[28] ;
 wire \pulse_width_counter_module.high_counter[29] ;
 wire \pulse_width_counter_module.high_counter[2] ;
 wire \pulse_width_counter_module.high_counter[30] ;
 wire \pulse_width_counter_module.high_counter[31] ;
 wire \pulse_width_counter_module.high_counter[3] ;
 wire \pulse_width_counter_module.high_counter[4] ;
 wire \pulse_width_counter_module.high_counter[5] ;
 wire \pulse_width_counter_module.high_counter[6] ;
 wire \pulse_width_counter_module.high_counter[7] ;
 wire \pulse_width_counter_module.high_counter[8] ;
 wire \pulse_width_counter_module.high_counter[9] ;
 wire \pulse_width_counter_module.low_counter[0] ;
 wire \pulse_width_counter_module.low_counter[10] ;
 wire \pulse_width_counter_module.low_counter[11] ;
 wire \pulse_width_counter_module.low_counter[12] ;
 wire \pulse_width_counter_module.low_counter[13] ;
 wire \pulse_width_counter_module.low_counter[14] ;
 wire \pulse_width_counter_module.low_counter[15] ;
 wire \pulse_width_counter_module.low_counter[16] ;
 wire \pulse_width_counter_module.low_counter[17] ;
 wire \pulse_width_counter_module.low_counter[18] ;
 wire \pulse_width_counter_module.low_counter[19] ;
 wire \pulse_width_counter_module.low_counter[1] ;
 wire \pulse_width_counter_module.low_counter[20] ;
 wire \pulse_width_counter_module.low_counter[21] ;
 wire \pulse_width_counter_module.low_counter[22] ;
 wire \pulse_width_counter_module.low_counter[23] ;
 wire \pulse_width_counter_module.low_counter[24] ;
 wire \pulse_width_counter_module.low_counter[25] ;
 wire \pulse_width_counter_module.low_counter[26] ;
 wire \pulse_width_counter_module.low_counter[27] ;
 wire \pulse_width_counter_module.low_counter[28] ;
 wire \pulse_width_counter_module.low_counter[29] ;
 wire \pulse_width_counter_module.low_counter[2] ;
 wire \pulse_width_counter_module.low_counter[30] ;
 wire \pulse_width_counter_module.low_counter[31] ;
 wire \pulse_width_counter_module.low_counter[3] ;
 wire \pulse_width_counter_module.low_counter[4] ;
 wire \pulse_width_counter_module.low_counter[5] ;
 wire \pulse_width_counter_module.low_counter[6] ;
 wire \pulse_width_counter_module.low_counter[7] ;
 wire \pulse_width_counter_module.low_counter[8] ;
 wire \pulse_width_counter_module.low_counter[9] ;
 wire \pulse_width_counter_module.previous_freq_in ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_inv_1 _1176_ (.Y(_0445_),
    .A(net1));
 sg13g2_buf_1 _1177_ (.A(_0445_),
    .X(_0446_));
 sg13g2_buf_8 _1178_ (.A(ui_in[0]),
    .X(_0447_));
 sg13g2_buf_2 _1179_ (.A(\pulse_width_counter_module.previous_freq_in ),
    .X(_0448_));
 sg13g2_nor2b_1 _1180_ (.A(_0447_),
    .B_N(_0448_),
    .Y(_0449_));
 sg13g2_buf_2 _1181_ (.A(_0449_),
    .X(_0450_));
 sg13g2_buf_1 _1182_ (.A(_0450_),
    .X(_0451_));
 sg13g2_nor2_1 _1183_ (.A(\mux.data_in[0] ),
    .B(net32),
    .Y(_0452_));
 sg13g2_nand2b_1 _1184_ (.Y(_0453_),
    .B(_0448_),
    .A_N(_0447_));
 sg13g2_buf_1 _1185_ (.A(_0453_),
    .X(_0454_));
 sg13g2_buf_1 _1186_ (.A(_0454_),
    .X(_0455_));
 sg13g2_buf_1 _1187_ (.A(_0455_),
    .X(_0456_));
 sg13g2_xor2_1 _1188_ (.B(\mux.data_in[64] ),
    .A(\mux.data_in[32] ),
    .X(_0457_));
 sg13g2_nor2_1 _1189_ (.A(net16),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_nor3_1 _1190_ (.A(net61),
    .B(_0452_),
    .C(_0458_),
    .Y(_0000_));
 sg13g2_nor2_1 _1191_ (.A(\mux.data_in[10] ),
    .B(net32),
    .Y(_0459_));
 sg13g2_buf_2 _1192_ (.A(\mux.data_in[41] ),
    .X(_0460_));
 sg13g2_buf_2 _1193_ (.A(\mux.data_in[73] ),
    .X(_0461_));
 sg13g2_nor2_1 _1194_ (.A(_0460_),
    .B(_0461_),
    .Y(_0462_));
 sg13g2_buf_1 _1195_ (.A(\mux.data_in[40] ),
    .X(_0463_));
 sg13g2_buf_2 _1196_ (.A(\mux.data_in[72] ),
    .X(_0464_));
 sg13g2_nand2_1 _1197_ (.Y(_0465_),
    .A(_0463_),
    .B(_0464_));
 sg13g2_nand2_1 _1198_ (.Y(_0466_),
    .A(_0460_),
    .B(_0461_));
 sg13g2_buf_2 _1199_ (.A(\mux.data_in[39] ),
    .X(_0467_));
 sg13g2_buf_2 _1200_ (.A(\mux.data_in[71] ),
    .X(_0468_));
 sg13g2_nand3_1 _1201_ (.B(_0467_),
    .C(_0468_),
    .A(_0464_),
    .Y(_0469_));
 sg13g2_nand3_1 _1202_ (.B(_0467_),
    .C(_0468_),
    .A(_0463_),
    .Y(_0470_));
 sg13g2_nand4_1 _1203_ (.B(_0466_),
    .C(_0469_),
    .A(_0465_),
    .Y(_0471_),
    .D(_0470_));
 sg13g2_nand2b_1 _1204_ (.Y(_0472_),
    .B(_0471_),
    .A_N(_0462_));
 sg13g2_xor2_1 _1205_ (.B(_0468_),
    .A(_0467_),
    .X(_0473_));
 sg13g2_xor2_1 _1206_ (.B(_0464_),
    .A(_0463_),
    .X(_0474_));
 sg13g2_xor2_1 _1207_ (.B(_0461_),
    .A(_0460_),
    .X(_0475_));
 sg13g2_nand3_1 _1208_ (.B(_0474_),
    .C(_0475_),
    .A(_0473_),
    .Y(_0476_));
 sg13g2_nor2_1 _1209_ (.A(\mux.data_in[33] ),
    .B(\mux.data_in[65] ),
    .Y(_0477_));
 sg13g2_a22oi_1 _1210_ (.Y(_0478_),
    .B1(\mux.data_in[33] ),
    .B2(\mux.data_in[65] ),
    .A2(\mux.data_in[64] ),
    .A1(\mux.data_in[32] ));
 sg13g2_xnor2_1 _1211_ (.Y(_0479_),
    .A(\mux.data_in[35] ),
    .B(\mux.data_in[67] ));
 sg13g2_buf_2 _1212_ (.A(\mux.data_in[66] ),
    .X(_0480_));
 sg13g2_xnor2_1 _1213_ (.Y(_0481_),
    .A(\mux.data_in[34] ),
    .B(_0480_));
 sg13g2_nor4_2 _1214_ (.A(_0477_),
    .B(_0478_),
    .C(_0479_),
    .Y(_0482_),
    .D(_0481_));
 sg13g2_nor2_1 _1215_ (.A(\mux.data_in[35] ),
    .B(\mux.data_in[67] ),
    .Y(_0483_));
 sg13g2_a22oi_1 _1216_ (.Y(_0484_),
    .B1(\mux.data_in[35] ),
    .B2(\mux.data_in[67] ),
    .A2(_0480_),
    .A1(\mux.data_in[34] ));
 sg13g2_nor2_2 _1217_ (.A(_0483_),
    .B(_0484_),
    .Y(_0485_));
 sg13g2_buf_1 _1218_ (.A(\mux.data_in[36] ),
    .X(_0486_));
 sg13g2_buf_2 _1219_ (.A(\mux.data_in[68] ),
    .X(_0487_));
 sg13g2_and2_1 _1220_ (.A(_0486_),
    .B(_0487_),
    .X(_0488_));
 sg13g2_buf_2 _1221_ (.A(\mux.data_in[70] ),
    .X(_0489_));
 sg13g2_inv_1 _1222_ (.Y(_0490_),
    .A(_0489_));
 sg13g2_buf_2 _1223_ (.A(\mux.data_in[37] ),
    .X(_0491_));
 sg13g2_buf_1 _1224_ (.A(\mux.data_in[69] ),
    .X(_0492_));
 sg13g2_buf_2 _1225_ (.A(\mux.data_in[38] ),
    .X(_0493_));
 sg13g2_nand3_1 _1226_ (.B(net60),
    .C(_0493_),
    .A(_0491_),
    .Y(_0494_));
 sg13g2_a21oi_1 _1227_ (.A1(_0491_),
    .A2(net60),
    .Y(_0495_),
    .B1(_0493_));
 sg13g2_a21oi_1 _1228_ (.A1(_0490_),
    .A2(_0494_),
    .Y(_0496_),
    .B1(_0495_));
 sg13g2_nor4_2 _1229_ (.A(_0482_),
    .B(_0485_),
    .C(_0488_),
    .Y(_0497_),
    .D(_0496_));
 sg13g2_inv_1 _1230_ (.Y(_0498_),
    .A(_0493_));
 sg13g2_nand2_1 _1231_ (.Y(_0499_),
    .A(_0491_),
    .B(net60));
 sg13g2_nor2_1 _1232_ (.A(_0486_),
    .B(_0487_),
    .Y(_0500_));
 sg13g2_nor2_1 _1233_ (.A(_0491_),
    .B(net60),
    .Y(_0501_));
 sg13g2_a221oi_1 _1234_ (.B2(_0500_),
    .C1(_0501_),
    .B1(_0499_),
    .A1(_0498_),
    .Y(_0502_),
    .A2(_0490_));
 sg13g2_a21oi_2 _1235_ (.B1(_0502_),
    .Y(_0503_),
    .A2(_0489_),
    .A1(_0493_));
 sg13g2_or3_1 _1236_ (.A(_0476_),
    .B(_0497_),
    .C(_0503_),
    .X(_0504_));
 sg13g2_nand2_1 _1237_ (.Y(_0505_),
    .A(_0472_),
    .B(_0504_));
 sg13g2_buf_2 _1238_ (.A(\mux.data_in[42] ),
    .X(_0506_));
 sg13g2_buf_2 _1239_ (.A(\mux.data_in[74] ),
    .X(_0507_));
 sg13g2_xor2_1 _1240_ (.B(_0507_),
    .A(_0506_),
    .X(_0508_));
 sg13g2_xor2_1 _1241_ (.B(_0508_),
    .A(_0505_),
    .X(_0509_));
 sg13g2_nor2_1 _1242_ (.A(net16),
    .B(_0509_),
    .Y(_0510_));
 sg13g2_nor3_1 _1243_ (.A(net61),
    .B(_0459_),
    .C(_0510_),
    .Y(_0001_));
 sg13g2_nand2_1 _1244_ (.Y(_0511_),
    .A(\mux.data_in[11] ),
    .B(net16));
 sg13g2_buf_1 _1245_ (.A(_0450_),
    .X(_0512_));
 sg13g2_buf_1 _1246_ (.A(net30),
    .X(_0513_));
 sg13g2_inv_1 _1247_ (.Y(_0514_),
    .A(_0506_));
 sg13g2_inv_1 _1248_ (.Y(_0515_),
    .A(_0507_));
 sg13g2_a22oi_1 _1249_ (.Y(_0516_),
    .B1(_0472_),
    .B2(_0504_),
    .A2(_0515_),
    .A1(_0514_));
 sg13g2_nor2_1 _1250_ (.A(_0514_),
    .B(_0515_),
    .Y(_0517_));
 sg13g2_nor2_1 _1251_ (.A(_0516_),
    .B(_0517_),
    .Y(_0518_));
 sg13g2_buf_2 _1252_ (.A(\mux.data_in[43] ),
    .X(_0519_));
 sg13g2_buf_2 _1253_ (.A(\mux.data_in[75] ),
    .X(_0520_));
 sg13g2_xor2_1 _1254_ (.B(_0520_),
    .A(_0519_),
    .X(_0521_));
 sg13g2_xnor2_1 _1255_ (.Y(_0522_),
    .A(_0518_),
    .B(_0521_));
 sg13g2_nand2_1 _1256_ (.Y(_0523_),
    .A(net15),
    .B(_0522_));
 sg13g2_buf_1 _1257_ (.A(_0445_),
    .X(_0524_));
 sg13g2_buf_1 _1258_ (.A(net59),
    .X(_0525_));
 sg13g2_a21oi_1 _1259_ (.A1(_0511_),
    .A2(_0523_),
    .Y(_0002_),
    .B1(_0525_));
 sg13g2_buf_1 _1260_ (.A(net1),
    .X(_0526_));
 sg13g2_nand2_1 _1261_ (.Y(_0527_),
    .A(_0526_),
    .B(_0450_));
 sg13g2_buf_1 _1262_ (.A(_0527_),
    .X(_0528_));
 sg13g2_inv_1 _1263_ (.Y(_0529_),
    .A(_0519_));
 sg13g2_o21ai_1 _1264_ (.B1(_0520_),
    .Y(_0530_),
    .A1(_0516_),
    .A2(_0517_));
 sg13g2_nor3_1 _1265_ (.A(_0520_),
    .B(_0516_),
    .C(_0517_),
    .Y(_0531_));
 sg13g2_a21oi_1 _1266_ (.A1(_0529_),
    .A2(_0530_),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_buf_2 _1267_ (.A(\mux.data_in[44] ),
    .X(_0533_));
 sg13g2_buf_2 _1268_ (.A(\mux.data_in[76] ),
    .X(_0534_));
 sg13g2_xor2_1 _1269_ (.B(_0534_),
    .A(_0533_),
    .X(_0535_));
 sg13g2_xnor2_1 _1270_ (.Y(_0536_),
    .A(_0532_),
    .B(_0535_));
 sg13g2_nor2_1 _1271_ (.A(_0445_),
    .B(_0450_),
    .Y(_0537_));
 sg13g2_buf_1 _1272_ (.A(_0537_),
    .X(_0538_));
 sg13g2_nand2_1 _1273_ (.Y(_0539_),
    .A(\mux.data_in[12] ),
    .B(net13));
 sg13g2_o21ai_1 _1274_ (.B1(_0539_),
    .Y(_0003_),
    .A1(net14),
    .A2(_0536_));
 sg13g2_nor2_1 _1275_ (.A(\mux.data_in[13] ),
    .B(net32),
    .Y(_0540_));
 sg13g2_buf_1 _1276_ (.A(net31),
    .X(_0541_));
 sg13g2_nand3_1 _1277_ (.B(_0521_),
    .C(_0535_),
    .A(_0508_),
    .Y(_0542_));
 sg13g2_nor4_2 _1278_ (.A(_0476_),
    .B(_0497_),
    .C(_0503_),
    .Y(_0543_),
    .D(_0542_));
 sg13g2_nor2_1 _1279_ (.A(_0533_),
    .B(_0534_),
    .Y(_0544_));
 sg13g2_a22oi_1 _1280_ (.Y(_0545_),
    .B1(_0533_),
    .B2(_0534_),
    .A2(_0520_),
    .A1(_0519_));
 sg13g2_a22oi_1 _1281_ (.Y(_0546_),
    .B1(_0506_),
    .B2(_0507_),
    .A2(_0461_),
    .A1(_0460_));
 sg13g2_nand4_1 _1282_ (.B(_0469_),
    .C(_0470_),
    .A(_0465_),
    .Y(_0547_),
    .D(_0546_));
 sg13g2_nand2_1 _1283_ (.Y(_0548_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_nor2_1 _1284_ (.A(_0506_),
    .B(_0507_),
    .Y(_0549_));
 sg13g2_a21oi_1 _1285_ (.A1(_0462_),
    .A2(_0548_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_nand4_1 _1286_ (.B(_0535_),
    .C(_0547_),
    .A(_0521_),
    .Y(_0551_),
    .D(_0550_));
 sg13g2_o21ai_1 _1287_ (.B1(_0551_),
    .Y(_0552_),
    .A1(_0544_),
    .A2(_0545_));
 sg13g2_nor2_1 _1288_ (.A(_0543_),
    .B(_0552_),
    .Y(_0553_));
 sg13g2_buf_2 _1289_ (.A(\mux.data_in[45] ),
    .X(_0554_));
 sg13g2_buf_2 _1290_ (.A(\mux.data_in[77] ),
    .X(_0555_));
 sg13g2_xnor2_1 _1291_ (.Y(_0556_),
    .A(_0554_),
    .B(_0555_));
 sg13g2_xor2_1 _1292_ (.B(_0556_),
    .A(_0553_),
    .X(_0557_));
 sg13g2_nor2_1 _1293_ (.A(net12),
    .B(_0557_),
    .Y(_0558_));
 sg13g2_nor3_1 _1294_ (.A(net61),
    .B(_0540_),
    .C(_0558_),
    .Y(_0004_));
 sg13g2_inv_1 _1295_ (.Y(_0559_),
    .A(_0554_));
 sg13g2_nor3_1 _1296_ (.A(_0555_),
    .B(_0543_),
    .C(_0552_),
    .Y(_0560_));
 sg13g2_o21ai_1 _1297_ (.B1(_0555_),
    .Y(_0561_),
    .A1(_0543_),
    .A2(_0552_));
 sg13g2_o21ai_1 _1298_ (.B1(_0561_),
    .Y(_0562_),
    .A1(_0559_),
    .A2(_0560_));
 sg13g2_buf_2 _1299_ (.A(\mux.data_in[46] ),
    .X(_0563_));
 sg13g2_buf_2 _1300_ (.A(\mux.data_in[78] ),
    .X(_0564_));
 sg13g2_xor2_1 _1301_ (.B(_0564_),
    .A(_0563_),
    .X(_0565_));
 sg13g2_xnor2_1 _1302_ (.Y(_0566_),
    .A(_0562_),
    .B(_0565_));
 sg13g2_nand2_1 _1303_ (.Y(_0567_),
    .A(\mux.data_in[14] ),
    .B(net13));
 sg13g2_o21ai_1 _1304_ (.B1(_0567_),
    .Y(_0005_),
    .A1(net14),
    .A2(_0566_));
 sg13g2_buf_1 _1305_ (.A(net63),
    .X(_0568_));
 sg13g2_buf_1 _1306_ (.A(_0454_),
    .X(_0569_));
 sg13g2_buf_2 _1307_ (.A(\mux.data_in[47] ),
    .X(_0570_));
 sg13g2_buf_2 _1308_ (.A(\mux.data_in[79] ),
    .X(_0571_));
 sg13g2_xor2_1 _1309_ (.B(_0571_),
    .A(_0570_),
    .X(_0572_));
 sg13g2_nor2_1 _1310_ (.A(_0563_),
    .B(_0564_),
    .Y(_0573_));
 sg13g2_a22oi_1 _1311_ (.Y(_0574_),
    .B1(_0563_),
    .B2(_0564_),
    .A2(_0555_),
    .A1(_0554_));
 sg13g2_nor2b_1 _1312_ (.A(_0556_),
    .B_N(_0565_),
    .Y(_0575_));
 sg13g2_o21ai_1 _1313_ (.B1(_0575_),
    .Y(_0576_),
    .A1(_0543_),
    .A2(_0552_));
 sg13g2_o21ai_1 _1314_ (.B1(_0576_),
    .Y(_0577_),
    .A1(_0573_),
    .A2(_0574_));
 sg13g2_xnor2_1 _1315_ (.Y(_0578_),
    .A(_0572_),
    .B(_0577_));
 sg13g2_buf_1 _1316_ (.A(_0454_),
    .X(_0579_));
 sg13g2_nand2_1 _1317_ (.Y(_0580_),
    .A(\mux.data_in[15] ),
    .B(net28));
 sg13g2_o21ai_1 _1318_ (.B1(_0580_),
    .Y(_0581_),
    .A1(net29),
    .A2(_0578_));
 sg13g2_and2_1 _1319_ (.A(_0568_),
    .B(_0581_),
    .X(_0006_));
 sg13g2_buf_2 _1320_ (.A(\mux.data_in[48] ),
    .X(_0582_));
 sg13g2_buf_1 _1321_ (.A(\mux.data_in[80] ),
    .X(_0583_));
 sg13g2_xor2_1 _1322_ (.B(net57),
    .A(_0582_),
    .X(_0584_));
 sg13g2_and2_1 _1323_ (.A(_0565_),
    .B(_0572_),
    .X(_0585_));
 sg13g2_nor2_1 _1324_ (.A(_0570_),
    .B(_0571_),
    .Y(_0586_));
 sg13g2_and2_1 _1325_ (.A(_0570_),
    .B(_0571_),
    .X(_0587_));
 sg13g2_a21oi_1 _1326_ (.A1(_0563_),
    .A2(_0564_),
    .Y(_0588_),
    .B1(_0587_));
 sg13g2_nor2_1 _1327_ (.A(_0586_),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_a21oi_1 _1328_ (.A1(_0562_),
    .A2(_0585_),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_xor2_1 _1329_ (.B(_0590_),
    .A(_0584_),
    .X(_0591_));
 sg13g2_buf_1 _1330_ (.A(net63),
    .X(_0592_));
 sg13g2_o21ai_1 _1331_ (.B1(net56),
    .Y(_0593_),
    .A1(\mux.data_in[16] ),
    .A2(net30));
 sg13g2_a21oi_1 _1332_ (.A1(net15),
    .A2(_0591_),
    .Y(_0007_),
    .B1(_0593_));
 sg13g2_nor2_1 _1333_ (.A(\mux.data_in[17] ),
    .B(net32),
    .Y(_0594_));
 sg13g2_nand2_1 _1334_ (.Y(_0595_),
    .A(_0572_),
    .B(_0584_));
 sg13g2_nand2_1 _1335_ (.Y(_0596_),
    .A(_0582_),
    .B(net57));
 sg13g2_nor2_1 _1336_ (.A(_0573_),
    .B(_0574_),
    .Y(_0597_));
 sg13g2_nand2_1 _1337_ (.Y(_0598_),
    .A(_0571_),
    .B(_0597_));
 sg13g2_o21ai_1 _1338_ (.B1(_0570_),
    .Y(_0599_),
    .A1(_0571_),
    .A2(_0597_));
 sg13g2_nand3_1 _1339_ (.B(_0598_),
    .C(_0599_),
    .A(_0596_),
    .Y(_0600_));
 sg13g2_o21ai_1 _1340_ (.B1(_0600_),
    .Y(_0601_),
    .A1(_0582_),
    .A2(net57));
 sg13g2_o21ai_1 _1341_ (.B1(_0601_),
    .Y(_0602_),
    .A1(_0576_),
    .A2(_0595_));
 sg13g2_buf_2 _1342_ (.A(\mux.data_in[49] ),
    .X(_0603_));
 sg13g2_buf_1 _1343_ (.A(\mux.data_in[81] ),
    .X(_0604_));
 sg13g2_xor2_1 _1344_ (.B(net55),
    .A(_0603_),
    .X(_0605_));
 sg13g2_xor2_1 _1345_ (.B(_0605_),
    .A(_0602_),
    .X(_0606_));
 sg13g2_nor2_1 _1346_ (.A(net12),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_nor3_1 _1347_ (.A(net61),
    .B(_0594_),
    .C(_0607_),
    .Y(_0008_));
 sg13g2_nor2_1 _1348_ (.A(_0603_),
    .B(net55),
    .Y(_0608_));
 sg13g2_nand2_1 _1349_ (.Y(_0609_),
    .A(_0533_),
    .B(_0534_));
 sg13g2_nor2_1 _1350_ (.A(_0519_),
    .B(_0520_),
    .Y(_0610_));
 sg13g2_a22oi_1 _1351_ (.Y(_0611_),
    .B1(_0519_),
    .B2(_0520_),
    .A2(_0507_),
    .A1(_0506_));
 sg13g2_or3_1 _1352_ (.A(_0544_),
    .B(_0610_),
    .C(_0611_),
    .X(_0612_));
 sg13g2_inv_1 _1353_ (.Y(_0613_),
    .A(_0555_));
 sg13g2_a21oi_1 _1354_ (.A1(_0609_),
    .A2(_0612_),
    .Y(_0614_),
    .B1(_0613_));
 sg13g2_nand3_1 _1355_ (.B(_0609_),
    .C(_0612_),
    .A(_0613_),
    .Y(_0615_));
 sg13g2_and2_1 _1356_ (.A(_0554_),
    .B(_0585_),
    .X(_0616_));
 sg13g2_a221oi_1 _1357_ (.B2(_0616_),
    .C1(_0589_),
    .B1(_0615_),
    .A1(_0585_),
    .Y(_0617_),
    .A2(_0614_));
 sg13g2_nand2b_1 _1358_ (.Y(_0618_),
    .B(_0617_),
    .A_N(net57));
 sg13g2_nor2b_1 _1359_ (.A(_0617_),
    .B_N(_0583_),
    .Y(_0619_));
 sg13g2_a221oi_1 _1360_ (.B2(_0582_),
    .C1(_0619_),
    .B1(_0618_),
    .A1(_0603_),
    .Y(_0620_),
    .A2(_0604_));
 sg13g2_nand3_1 _1361_ (.B(_0585_),
    .C(_0605_),
    .A(_0584_),
    .Y(_0621_));
 sg13g2_nor3_1 _1362_ (.A(_0542_),
    .B(_0556_),
    .C(_0621_),
    .Y(_0622_));
 sg13g2_nand2_1 _1363_ (.Y(_0623_),
    .A(_0505_),
    .B(_0622_));
 sg13g2_o21ai_1 _1364_ (.B1(_0623_),
    .Y(_0624_),
    .A1(_0608_),
    .A2(_0620_));
 sg13g2_buf_1 _1365_ (.A(\mux.data_in[82] ),
    .X(_0625_));
 sg13g2_xor2_1 _1366_ (.B(_0625_),
    .A(\mux.data_in[50] ),
    .X(_0626_));
 sg13g2_xnor2_1 _1367_ (.Y(_0627_),
    .A(_0624_),
    .B(_0626_));
 sg13g2_nand2_1 _1368_ (.Y(_0628_),
    .A(\mux.data_in[18] ),
    .B(net13));
 sg13g2_o21ai_1 _1369_ (.B1(_0628_),
    .Y(_0009_),
    .A1(net14),
    .A2(_0627_));
 sg13g2_nor2_1 _1370_ (.A(\mux.data_in[19] ),
    .B(_0451_),
    .Y(_0629_));
 sg13g2_or4_1 _1371_ (.A(_0476_),
    .B(_0497_),
    .C(_0503_),
    .D(_0542_),
    .X(_0630_));
 sg13g2_or2_1 _1372_ (.X(_0631_),
    .B(_0625_),
    .A(\mux.data_in[50] ));
 sg13g2_buf_1 _1373_ (.A(_0631_),
    .X(_0632_));
 sg13g2_and3_1 _1374_ (.X(_0633_),
    .A(_0583_),
    .B(_0587_),
    .C(_0632_));
 sg13g2_a21o_1 _1375_ (.A2(_0571_),
    .A1(_0570_),
    .B1(net57),
    .X(_0634_));
 sg13g2_and3_1 _1376_ (.X(_0635_),
    .A(_0582_),
    .B(_0632_),
    .C(_0634_));
 sg13g2_o21ai_1 _1377_ (.B1(_0603_),
    .Y(_0636_),
    .A1(_0633_),
    .A2(_0635_));
 sg13g2_nand4_1 _1378_ (.B(net55),
    .C(_0587_),
    .A(net57),
    .Y(_0637_),
    .D(_0632_));
 sg13g2_nand4_1 _1379_ (.B(net55),
    .C(_0632_),
    .A(_0582_),
    .Y(_0638_),
    .D(_0634_));
 sg13g2_nand3_1 _1380_ (.B(net55),
    .C(_0625_),
    .A(_0603_),
    .Y(_0639_));
 sg13g2_a21oi_1 _1381_ (.A1(_0603_),
    .A2(net55),
    .Y(_0640_),
    .B1(_0625_));
 sg13g2_nand2b_1 _1382_ (.Y(_0641_),
    .B(\mux.data_in[50] ),
    .A_N(_0640_));
 sg13g2_and4_1 _1383_ (.A(_0637_),
    .B(_0638_),
    .C(_0639_),
    .D(_0641_),
    .X(_0642_));
 sg13g2_nor2_1 _1384_ (.A(_0544_),
    .B(_0545_),
    .Y(_0643_));
 sg13g2_nor2_1 _1385_ (.A(_0643_),
    .B(_0597_),
    .Y(_0644_));
 sg13g2_and4_1 _1386_ (.A(_0551_),
    .B(_0636_),
    .C(_0642_),
    .D(_0644_),
    .X(_0645_));
 sg13g2_and4_1 _1387_ (.A(_0572_),
    .B(_0584_),
    .C(_0605_),
    .D(_0626_),
    .X(_0646_));
 sg13g2_o21ai_1 _1388_ (.B1(_0646_),
    .Y(_0647_),
    .A1(_0575_),
    .A2(_0597_));
 sg13g2_and3_1 _1389_ (.X(_0648_),
    .A(_0636_),
    .B(_0642_),
    .C(_0647_));
 sg13g2_a21oi_2 _1390_ (.B1(_0648_),
    .Y(_0649_),
    .A2(_0645_),
    .A1(_0630_));
 sg13g2_buf_2 _1391_ (.A(\mux.data_in[51] ),
    .X(_0650_));
 sg13g2_buf_2 _1392_ (.A(\mux.data_in[83] ),
    .X(_0651_));
 sg13g2_xnor2_1 _1393_ (.Y(_0652_),
    .A(_0650_),
    .B(_0651_));
 sg13g2_xnor2_1 _1394_ (.Y(_0653_),
    .A(_0649_),
    .B(_0652_));
 sg13g2_nor2_1 _1395_ (.A(net12),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_nor3_1 _1396_ (.A(net61),
    .B(_0629_),
    .C(_0654_),
    .Y(_0010_));
 sg13g2_nand2_1 _1397_ (.Y(_0655_),
    .A(\mux.data_in[1] ),
    .B(net16));
 sg13g2_nand2_1 _1398_ (.Y(_0656_),
    .A(\mux.data_in[32] ),
    .B(\mux.data_in[64] ));
 sg13g2_xor2_1 _1399_ (.B(\mux.data_in[65] ),
    .A(\mux.data_in[33] ),
    .X(_0657_));
 sg13g2_xnor2_1 _1400_ (.Y(_0658_),
    .A(_0656_),
    .B(_0657_));
 sg13g2_nand2_1 _1401_ (.Y(_0659_),
    .A(net15),
    .B(_0658_));
 sg13g2_a21oi_1 _1402_ (.A1(_0655_),
    .A2(_0659_),
    .Y(_0011_),
    .B1(net45));
 sg13g2_a21o_1 _1403_ (.A2(_0649_),
    .A1(_0651_),
    .B1(_0650_),
    .X(_0660_));
 sg13g2_o21ai_1 _1404_ (.B1(_0660_),
    .Y(_0661_),
    .A1(_0651_),
    .A2(_0649_));
 sg13g2_buf_2 _1405_ (.A(\mux.data_in[52] ),
    .X(_0662_));
 sg13g2_buf_2 _1406_ (.A(\mux.data_in[84] ),
    .X(_0663_));
 sg13g2_xor2_1 _1407_ (.B(_0663_),
    .A(_0662_),
    .X(_0664_));
 sg13g2_xor2_1 _1408_ (.B(_0664_),
    .A(_0661_),
    .X(_0665_));
 sg13g2_o21ai_1 _1409_ (.B1(net56),
    .Y(_0666_),
    .A1(\mux.data_in[20] ),
    .A2(net30));
 sg13g2_a21oi_1 _1410_ (.A1(net15),
    .A2(_0665_),
    .Y(_0012_),
    .B1(_0666_));
 sg13g2_nor2b_1 _1411_ (.A(_0652_),
    .B_N(_0664_),
    .Y(_0667_));
 sg13g2_nor2_1 _1412_ (.A(_0662_),
    .B(_0663_),
    .Y(_0668_));
 sg13g2_a22oi_1 _1413_ (.Y(_0669_),
    .B1(_0662_),
    .B2(_0663_),
    .A2(_0651_),
    .A1(_0650_));
 sg13g2_nor2_1 _1414_ (.A(_0668_),
    .B(_0669_),
    .Y(_0670_));
 sg13g2_a21oi_1 _1415_ (.A1(_0649_),
    .A2(_0667_),
    .Y(_0671_),
    .B1(_0670_));
 sg13g2_buf_2 _1416_ (.A(\mux.data_in[53] ),
    .X(_0672_));
 sg13g2_buf_2 _1417_ (.A(\mux.data_in[85] ),
    .X(_0673_));
 sg13g2_xor2_1 _1418_ (.B(_0673_),
    .A(_0672_),
    .X(_0674_));
 sg13g2_xor2_1 _1419_ (.B(_0674_),
    .A(_0671_),
    .X(_0675_));
 sg13g2_o21ai_1 _1420_ (.B1(net56),
    .Y(_0676_),
    .A1(\mux.data_in[21] ),
    .A2(net30));
 sg13g2_a21oi_1 _1421_ (.A1(net15),
    .A2(_0675_),
    .Y(_0013_),
    .B1(_0676_));
 sg13g2_buf_2 _1422_ (.A(\mux.data_in[54] ),
    .X(_0677_));
 sg13g2_xnor2_1 _1423_ (.Y(_0678_),
    .A(_0677_),
    .B(\mux.data_in[86] ));
 sg13g2_nand2_1 _1424_ (.Y(_0679_),
    .A(_0664_),
    .B(_0674_));
 sg13g2_nor2_1 _1425_ (.A(_0652_),
    .B(_0679_),
    .Y(_0680_));
 sg13g2_nor2_1 _1426_ (.A(_0672_),
    .B(_0673_),
    .Y(_0681_));
 sg13g2_nand2_1 _1427_ (.Y(_0682_),
    .A(_0672_),
    .B(_0673_));
 sg13g2_o21ai_1 _1428_ (.B1(_0682_),
    .Y(_0683_),
    .A1(_0668_),
    .A2(_0669_));
 sg13g2_nor2b_1 _1429_ (.A(_0681_),
    .B_N(_0683_),
    .Y(_0684_));
 sg13g2_a21oi_1 _1430_ (.A1(_0649_),
    .A2(_0680_),
    .Y(_0685_),
    .B1(_0684_));
 sg13g2_xnor2_1 _1431_ (.Y(_0686_),
    .A(_0678_),
    .B(_0685_));
 sg13g2_o21ai_1 _1432_ (.B1(net56),
    .Y(_0687_),
    .A1(\mux.data_in[22] ),
    .A2(net30));
 sg13g2_a21oi_1 _1433_ (.A1(_0513_),
    .A2(_0686_),
    .Y(_0014_),
    .B1(_0687_));
 sg13g2_and2_1 _1434_ (.A(_0636_),
    .B(_0642_),
    .X(_0688_));
 sg13g2_or3_1 _1435_ (.A(_0652_),
    .B(_0678_),
    .C(_0679_),
    .X(_0689_));
 sg13g2_a221oi_1 _1436_ (.B2(_0630_),
    .C1(_0689_),
    .B1(_0645_),
    .A1(_0688_),
    .Y(_0690_),
    .A2(_0647_));
 sg13g2_buf_1 _1437_ (.A(_0690_),
    .X(_0691_));
 sg13g2_inv_1 _1438_ (.Y(_0692_),
    .A(_0677_));
 sg13g2_inv_1 _1439_ (.Y(_0693_),
    .A(\mux.data_in[86] ));
 sg13g2_nor2_1 _1440_ (.A(_0692_),
    .B(_0693_),
    .Y(_0694_));
 sg13g2_o21ai_1 _1441_ (.B1(_0684_),
    .Y(_0695_),
    .A1(_0677_),
    .A2(\mux.data_in[86] ));
 sg13g2_nand2b_2 _1442_ (.Y(_0696_),
    .B(_0695_),
    .A_N(_0694_));
 sg13g2_nor2_1 _1443_ (.A(_0691_),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_buf_1 _1444_ (.A(\mux.data_in[55] ),
    .X(_0698_));
 sg13g2_buf_1 _1445_ (.A(\mux.data_in[87] ),
    .X(_0699_));
 sg13g2_xnor2_1 _1446_ (.Y(_0700_),
    .A(net54),
    .B(net53));
 sg13g2_xnor2_1 _1447_ (.Y(_0701_),
    .A(_0697_),
    .B(_0700_));
 sg13g2_o21ai_1 _1448_ (.B1(net56),
    .Y(_0702_),
    .A1(\mux.data_in[23] ),
    .A2(net30));
 sg13g2_a21oi_1 _1449_ (.A1(_0513_),
    .A2(_0701_),
    .Y(_0015_),
    .B1(_0702_));
 sg13g2_buf_2 _1450_ (.A(\mux.data_in[56] ),
    .X(_0703_));
 sg13g2_buf_1 _1451_ (.A(\mux.data_in[88] ),
    .X(_0704_));
 sg13g2_xor2_1 _1452_ (.B(net52),
    .A(_0703_),
    .X(_0705_));
 sg13g2_inv_1 _1453_ (.Y(_0706_),
    .A(net53));
 sg13g2_o21ai_1 _1454_ (.B1(net54),
    .Y(_0707_),
    .A1(_0691_),
    .A2(_0696_));
 sg13g2_nor3_1 _1455_ (.A(net54),
    .B(_0691_),
    .C(_0696_),
    .Y(_0708_));
 sg13g2_a21oi_1 _1456_ (.A1(_0706_),
    .A2(_0707_),
    .Y(_0709_),
    .B1(_0708_));
 sg13g2_xnor2_1 _1457_ (.Y(_0710_),
    .A(_0705_),
    .B(_0709_));
 sg13g2_nand2_1 _1458_ (.Y(_0711_),
    .A(\mux.data_in[24] ),
    .B(net13));
 sg13g2_o21ai_1 _1459_ (.B1(_0711_),
    .Y(_0016_),
    .A1(net14),
    .A2(_0710_));
 sg13g2_or2_1 _1460_ (.X(_0712_),
    .B(_0696_),
    .A(_0691_));
 sg13g2_a221oi_1 _1461_ (.B2(_0712_),
    .C1(net54),
    .B1(net53),
    .A1(_0703_),
    .Y(_0713_),
    .A2(net52));
 sg13g2_a21oi_1 _1462_ (.A1(_0703_),
    .A2(net52),
    .Y(_0714_),
    .B1(net53));
 sg13g2_nor2_1 _1463_ (.A(_0703_),
    .B(net52),
    .Y(_0715_));
 sg13g2_a21o_1 _1464_ (.A2(_0714_),
    .A1(_0697_),
    .B1(_0715_),
    .X(_0716_));
 sg13g2_buf_2 _1465_ (.A(\mux.data_in[57] ),
    .X(_0717_));
 sg13g2_buf_2 _1466_ (.A(\mux.data_in[89] ),
    .X(_0718_));
 sg13g2_xor2_1 _1467_ (.B(_0718_),
    .A(_0717_),
    .X(_0719_));
 sg13g2_nor2b_1 _1468_ (.A(net14),
    .B_N(_0719_),
    .Y(_0720_));
 sg13g2_o21ai_1 _1469_ (.B1(_0720_),
    .Y(_0721_),
    .A1(_0713_),
    .A2(_0716_));
 sg13g2_or4_1 _1470_ (.A(net14),
    .B(_0713_),
    .C(_0716_),
    .D(_0719_),
    .X(_0722_));
 sg13g2_nand2_1 _1471_ (.Y(_0723_),
    .A(\mux.data_in[25] ),
    .B(net13));
 sg13g2_nand3_1 _1472_ (.B(_0722_),
    .C(_0723_),
    .A(_0721_),
    .Y(_0017_));
 sg13g2_buf_1 _1473_ (.A(_0454_),
    .X(_0724_));
 sg13g2_nor2_1 _1474_ (.A(_0717_),
    .B(_0718_),
    .Y(_0725_));
 sg13g2_a21oi_1 _1475_ (.A1(net54),
    .A2(net53),
    .Y(_0726_),
    .B1(net52));
 sg13g2_nand3_1 _1476_ (.B(net54),
    .C(net53),
    .A(net52),
    .Y(_0727_));
 sg13g2_nor2b_1 _1477_ (.A(_0703_),
    .B_N(_0727_),
    .Y(_0728_));
 sg13g2_nor3_1 _1478_ (.A(_0725_),
    .B(_0726_),
    .C(_0728_),
    .Y(_0729_));
 sg13g2_a21oi_1 _1479_ (.A1(_0717_),
    .A2(_0718_),
    .Y(_0730_),
    .B1(_0729_));
 sg13g2_nand2_1 _1480_ (.Y(_0731_),
    .A(_0705_),
    .B(_0719_));
 sg13g2_nor2_1 _1481_ (.A(_0700_),
    .B(_0731_),
    .Y(_0732_));
 sg13g2_o21ai_1 _1482_ (.B1(_0732_),
    .Y(_0733_),
    .A1(_0691_),
    .A2(_0696_));
 sg13g2_buf_2 _1483_ (.A(\mux.data_in[58] ),
    .X(_0734_));
 sg13g2_buf_2 _1484_ (.A(\mux.data_in[90] ),
    .X(_0735_));
 sg13g2_xor2_1 _1485_ (.B(_0735_),
    .A(_0734_),
    .X(_0736_));
 sg13g2_a21oi_1 _1486_ (.A1(_0730_),
    .A2(_0733_),
    .Y(_0737_),
    .B1(_0736_));
 sg13g2_and3_1 _1487_ (.X(_0738_),
    .A(_0736_),
    .B(_0730_),
    .C(_0733_));
 sg13g2_nor3_1 _1488_ (.A(_0724_),
    .B(_0737_),
    .C(_0738_),
    .Y(_0739_));
 sg13g2_o21ai_1 _1489_ (.B1(_0592_),
    .Y(_0740_),
    .A1(\mux.data_in[26] ),
    .A2(_0451_));
 sg13g2_nor2_1 _1490_ (.A(_0739_),
    .B(_0740_),
    .Y(_0018_));
 sg13g2_nand2_1 _1491_ (.Y(_0741_),
    .A(\mux.data_in[27] ),
    .B(net13));
 sg13g2_inv_1 _1492_ (.Y(_0742_),
    .A(_0734_));
 sg13g2_inv_1 _1493_ (.Y(_0743_),
    .A(_0735_));
 sg13g2_a22oi_1 _1494_ (.Y(_0744_),
    .B1(_0730_),
    .B2(_0733_),
    .A2(_0743_),
    .A1(_0742_));
 sg13g2_nor2_1 _1495_ (.A(_0742_),
    .B(_0743_),
    .Y(_0745_));
 sg13g2_xor2_1 _1496_ (.B(\mux.data_in[91] ),
    .A(\mux.data_in[59] ),
    .X(_0746_));
 sg13g2_inv_1 _1497_ (.Y(_0747_),
    .A(_0746_));
 sg13g2_or4_1 _1498_ (.A(_0527_),
    .B(_0744_),
    .C(_0745_),
    .D(_0747_),
    .X(_0748_));
 sg13g2_nor2_1 _1499_ (.A(net14),
    .B(_0746_),
    .Y(_0749_));
 sg13g2_o21ai_1 _1500_ (.B1(_0749_),
    .Y(_0750_),
    .A1(_0744_),
    .A2(_0745_));
 sg13g2_nand3_1 _1501_ (.B(_0748_),
    .C(_0750_),
    .A(_0741_),
    .Y(_0019_));
 sg13g2_nor2_1 _1502_ (.A(\mux.data_in[28] ),
    .B(net30),
    .Y(_0751_));
 sg13g2_nor4_2 _1503_ (.A(_0678_),
    .B(_0679_),
    .C(_0700_),
    .Y(_0752_),
    .D(_0731_));
 sg13g2_and2_1 _1504_ (.A(_0736_),
    .B(_0746_),
    .X(_0753_));
 sg13g2_and3_1 _1505_ (.X(_0754_),
    .A(_0650_),
    .B(_0651_),
    .C(_0753_));
 sg13g2_a22oi_1 _1506_ (.Y(_0755_),
    .B1(_0717_),
    .B2(_0718_),
    .A2(net52),
    .A1(_0703_));
 sg13g2_nor2_1 _1507_ (.A(_0725_),
    .B(_0755_),
    .Y(_0756_));
 sg13g2_and2_1 _1508_ (.A(\mux.data_in[59] ),
    .B(\mux.data_in[91] ),
    .X(_0757_));
 sg13g2_nor3_1 _1509_ (.A(_0735_),
    .B(_0756_),
    .C(_0757_),
    .Y(_0758_));
 sg13g2_nor3_1 _1510_ (.A(_0734_),
    .B(_0756_),
    .C(_0757_),
    .Y(_0759_));
 sg13g2_a22oi_1 _1511_ (.Y(_0760_),
    .B1(_0672_),
    .B2(_0673_),
    .A2(_0663_),
    .A1(_0662_));
 sg13g2_nor3_1 _1512_ (.A(_0693_),
    .B(_0681_),
    .C(_0760_),
    .Y(_0761_));
 sg13g2_nor3_1 _1513_ (.A(_0692_),
    .B(_0681_),
    .C(_0760_),
    .Y(_0762_));
 sg13g2_or4_1 _1514_ (.A(net53),
    .B(_0694_),
    .C(_0761_),
    .D(_0762_),
    .X(_0763_));
 sg13g2_and3_1 _1515_ (.X(_0764_),
    .A(_0698_),
    .B(_0705_),
    .C(_0719_));
 sg13g2_nor2_1 _1516_ (.A(_0706_),
    .B(_0731_),
    .Y(_0765_));
 sg13g2_o21ai_1 _1517_ (.B1(_0693_),
    .Y(_0766_),
    .A1(_0681_),
    .A2(_0760_));
 sg13g2_a21o_1 _1518_ (.A2(_0766_),
    .A1(_0677_),
    .B1(_0761_),
    .X(_0767_));
 sg13g2_a22oi_1 _1519_ (.Y(_0768_),
    .B1(_0765_),
    .B2(_0767_),
    .A2(_0764_),
    .A1(_0763_));
 sg13g2_o21ai_1 _1520_ (.B1(_0768_),
    .Y(_0769_),
    .A1(_0758_),
    .A2(_0759_));
 sg13g2_nor2_1 _1521_ (.A(\mux.data_in[59] ),
    .B(\mux.data_in[91] ),
    .Y(_0770_));
 sg13g2_nor3_1 _1522_ (.A(_0734_),
    .B(_0735_),
    .C(_0757_),
    .Y(_0771_));
 sg13g2_nor2_1 _1523_ (.A(_0770_),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_nand3_1 _1524_ (.B(_0752_),
    .C(_0753_),
    .A(_0651_),
    .Y(_0773_));
 sg13g2_nand3_1 _1525_ (.B(_0752_),
    .C(_0753_),
    .A(_0650_),
    .Y(_0774_));
 sg13g2_a221oi_1 _1526_ (.B2(_0774_),
    .C1(_0648_),
    .B1(_0773_),
    .A1(_0630_),
    .Y(_0775_),
    .A2(_0645_));
 sg13g2_a221oi_1 _1527_ (.B2(_0772_),
    .C1(_0775_),
    .B1(_0769_),
    .A1(_0752_),
    .Y(_0776_),
    .A2(_0754_));
 sg13g2_xor2_1 _1528_ (.B(\mux.data_in[92] ),
    .A(\mux.data_in[60] ),
    .X(_0777_));
 sg13g2_xnor2_1 _1529_ (.Y(_0778_),
    .A(_0776_),
    .B(_0777_));
 sg13g2_nor2_1 _1530_ (.A(_0541_),
    .B(_0778_),
    .Y(_0779_));
 sg13g2_nor3_1 _1531_ (.A(_0446_),
    .B(_0751_),
    .C(_0779_),
    .Y(_0020_));
 sg13g2_inv_1 _1532_ (.Y(_0780_),
    .A(\mux.data_in[92] ));
 sg13g2_nor2_1 _1533_ (.A(_0780_),
    .B(_0776_),
    .Y(_0781_));
 sg13g2_inv_1 _1534_ (.Y(_0782_),
    .A(\mux.data_in[60] ));
 sg13g2_a21oi_1 _1535_ (.A1(_0780_),
    .A2(_0776_),
    .Y(_0783_),
    .B1(_0782_));
 sg13g2_xor2_1 _1536_ (.B(\mux.data_in[93] ),
    .A(\mux.data_in[61] ),
    .X(_0784_));
 sg13g2_nand3_1 _1537_ (.B(_0512_),
    .C(_0784_),
    .A(_0526_),
    .Y(_0785_));
 sg13g2_nor3_1 _1538_ (.A(_0781_),
    .B(_0783_),
    .C(_0785_),
    .Y(_0786_));
 sg13g2_nor2_1 _1539_ (.A(_0528_),
    .B(_0784_),
    .Y(_0787_));
 sg13g2_o21ai_1 _1540_ (.B1(_0787_),
    .Y(_0788_),
    .A1(_0781_),
    .A2(_0783_));
 sg13g2_nand2_1 _1541_ (.Y(_0789_),
    .A(\mux.data_in[29] ),
    .B(net13));
 sg13g2_nand3b_1 _1542_ (.B(_0788_),
    .C(_0789_),
    .Y(_0021_),
    .A_N(_0786_));
 sg13g2_nand2_1 _1543_ (.Y(_0790_),
    .A(\mux.data_in[2] ),
    .B(net16));
 sg13g2_nor2_1 _1544_ (.A(_0477_),
    .B(_0478_),
    .Y(_0791_));
 sg13g2_xnor2_1 _1545_ (.Y(_0792_),
    .A(_0791_),
    .B(_0481_));
 sg13g2_nand2_1 _1546_ (.Y(_0793_),
    .A(net15),
    .B(_0792_));
 sg13g2_a21oi_1 _1547_ (.A1(_0790_),
    .A2(_0793_),
    .Y(_0022_),
    .B1(net45));
 sg13g2_nand2_1 _1548_ (.Y(_0794_),
    .A(\mux.data_in[30] ),
    .B(_0538_));
 sg13g2_inv_1 _1549_ (.Y(_0795_),
    .A(\mux.data_in[61] ));
 sg13g2_inv_1 _1550_ (.Y(_0796_),
    .A(\mux.data_in[93] ));
 sg13g2_a221oi_1 _1551_ (.B2(_0796_),
    .C1(_0776_),
    .B1(_0795_),
    .A1(_0782_),
    .Y(_0797_),
    .A2(_0780_));
 sg13g2_nor2_1 _1552_ (.A(_0782_),
    .B(_0780_),
    .Y(_0798_));
 sg13g2_o21ai_1 _1553_ (.B1(_0798_),
    .Y(_0799_),
    .A1(\mux.data_in[61] ),
    .A2(\mux.data_in[93] ));
 sg13g2_o21ai_1 _1554_ (.B1(_0799_),
    .Y(_0800_),
    .A1(_0795_),
    .A2(_0796_));
 sg13g2_xnor2_1 _1555_ (.Y(_0801_),
    .A(\mux.data_in[62] ),
    .B(\mux.data_in[94] ));
 sg13g2_or4_1 _1556_ (.A(_0527_),
    .B(_0797_),
    .C(_0800_),
    .D(_0801_),
    .X(_0802_));
 sg13g2_nor2b_1 _1557_ (.A(net14),
    .B_N(_0801_),
    .Y(_0803_));
 sg13g2_o21ai_1 _1558_ (.B1(_0803_),
    .Y(_0804_),
    .A1(_0797_),
    .A2(_0800_));
 sg13g2_nand3_1 _1559_ (.B(_0802_),
    .C(_0804_),
    .A(_0794_),
    .Y(_0023_));
 sg13g2_nand2_1 _1560_ (.Y(_0805_),
    .A(\mux.data_in[62] ),
    .B(\mux.data_in[94] ));
 sg13g2_xor2_1 _1561_ (.B(\mux.data_in[95] ),
    .A(\mux.data_in[63] ),
    .X(_0806_));
 sg13g2_nor2b_1 _1562_ (.A(_0527_),
    .B_N(_0806_),
    .Y(_0807_));
 sg13g2_nand2_1 _1563_ (.Y(_0808_),
    .A(_0805_),
    .B(_0807_));
 sg13g2_nor3_1 _1564_ (.A(_0797_),
    .B(_0800_),
    .C(_0808_),
    .Y(_0809_));
 sg13g2_nor2_1 _1565_ (.A(\mux.data_in[62] ),
    .B(\mux.data_in[94] ),
    .Y(_0810_));
 sg13g2_nor3_1 _1566_ (.A(_0528_),
    .B(_0806_),
    .C(_0810_),
    .Y(_0811_));
 sg13g2_o21ai_1 _1567_ (.B1(_0811_),
    .Y(_0812_),
    .A1(_0797_),
    .A2(_0800_));
 sg13g2_nor3_1 _1568_ (.A(_0527_),
    .B(_0806_),
    .C(_0805_),
    .Y(_0813_));
 sg13g2_a221oi_1 _1569_ (.B2(_0810_),
    .C1(_0813_),
    .B1(_0807_),
    .A1(\mux.data_in[31] ),
    .Y(_0814_),
    .A2(_0538_));
 sg13g2_nand3b_1 _1570_ (.B(_0812_),
    .C(_0814_),
    .Y(_0024_),
    .A_N(_0809_));
 sg13g2_nand2_1 _1571_ (.Y(_0815_),
    .A(\mux.data_in[3] ),
    .B(net16));
 sg13g2_a21oi_1 _1572_ (.A1(_0480_),
    .A2(_0791_),
    .Y(_0816_),
    .B1(\mux.data_in[34] ));
 sg13g2_nor2_1 _1573_ (.A(_0480_),
    .B(_0791_),
    .Y(_0817_));
 sg13g2_nor2_1 _1574_ (.A(_0816_),
    .B(_0817_),
    .Y(_0818_));
 sg13g2_xnor2_1 _1575_ (.Y(_0819_),
    .A(_0479_),
    .B(_0818_));
 sg13g2_nand2_1 _1576_ (.Y(_0820_),
    .A(net15),
    .B(_0819_));
 sg13g2_buf_1 _1577_ (.A(net59),
    .X(_0821_));
 sg13g2_a21oi_1 _1578_ (.A1(_0815_),
    .A2(_0820_),
    .Y(_0025_),
    .B1(net44));
 sg13g2_nor2_1 _1579_ (.A(\mux.data_in[4] ),
    .B(net30),
    .Y(_0822_));
 sg13g2_nor2_1 _1580_ (.A(_0482_),
    .B(_0485_),
    .Y(_0823_));
 sg13g2_xor2_1 _1581_ (.B(_0487_),
    .A(_0486_),
    .X(_0824_));
 sg13g2_xnor2_1 _1582_ (.Y(_0825_),
    .A(_0823_),
    .B(_0824_));
 sg13g2_nor2_1 _1583_ (.A(_0541_),
    .B(_0825_),
    .Y(_0826_));
 sg13g2_nor3_1 _1584_ (.A(_0446_),
    .B(_0822_),
    .C(_0826_),
    .Y(_0026_));
 sg13g2_nand2_1 _1585_ (.Y(_0827_),
    .A(\mux.data_in[5] ),
    .B(net16));
 sg13g2_inv_1 _1586_ (.Y(_0828_),
    .A(_0486_));
 sg13g2_nor3_1 _1587_ (.A(_0487_),
    .B(_0482_),
    .C(_0485_),
    .Y(_0829_));
 sg13g2_o21ai_1 _1588_ (.B1(_0487_),
    .Y(_0830_),
    .A1(_0482_),
    .A2(_0485_));
 sg13g2_o21ai_1 _1589_ (.B1(_0830_),
    .Y(_0831_),
    .A1(_0828_),
    .A2(_0829_));
 sg13g2_xnor2_1 _1590_ (.Y(_0832_),
    .A(_0491_),
    .B(net60));
 sg13g2_xnor2_1 _1591_ (.Y(_0833_),
    .A(_0831_),
    .B(_0832_));
 sg13g2_nand2_1 _1592_ (.Y(_0834_),
    .A(net15),
    .B(_0833_));
 sg13g2_a21oi_1 _1593_ (.A1(_0827_),
    .A2(_0834_),
    .Y(_0027_),
    .B1(net44));
 sg13g2_nand2_1 _1594_ (.Y(_0835_),
    .A(\mux.data_in[6] ),
    .B(_0456_));
 sg13g2_buf_1 _1595_ (.A(_0450_),
    .X(_0836_));
 sg13g2_a21o_1 _1596_ (.A2(_0831_),
    .A1(net60),
    .B1(_0491_),
    .X(_0837_));
 sg13g2_o21ai_1 _1597_ (.B1(_0837_),
    .Y(_0838_),
    .A1(net60),
    .A2(_0831_));
 sg13g2_xor2_1 _1598_ (.B(_0489_),
    .A(_0493_),
    .X(_0839_));
 sg13g2_xnor2_1 _1599_ (.Y(_0840_),
    .A(_0838_),
    .B(_0839_));
 sg13g2_nand2_1 _1600_ (.Y(_0841_),
    .A(_0836_),
    .B(_0840_));
 sg13g2_a21oi_1 _1601_ (.A1(_0835_),
    .A2(_0841_),
    .Y(_0028_),
    .B1(_0821_));
 sg13g2_nand2_1 _1602_ (.Y(_0842_),
    .A(\mux.data_in[7] ),
    .B(_0456_));
 sg13g2_nor2_1 _1603_ (.A(_0497_),
    .B(_0503_),
    .Y(_0843_));
 sg13g2_xor2_1 _1604_ (.B(_0843_),
    .A(_0473_),
    .X(_0844_));
 sg13g2_nand2_1 _1605_ (.Y(_0845_),
    .A(_0836_),
    .B(_0844_));
 sg13g2_a21oi_1 _1606_ (.A1(_0842_),
    .A2(_0845_),
    .Y(_0029_),
    .B1(_0821_));
 sg13g2_buf_1 _1607_ (.A(net61),
    .X(_0846_));
 sg13g2_inv_1 _1608_ (.Y(_0847_),
    .A(_0468_));
 sg13g2_o21ai_1 _1609_ (.B1(_0847_),
    .Y(_0848_),
    .A1(_0497_),
    .A2(_0503_));
 sg13g2_nor3_1 _1610_ (.A(_0847_),
    .B(_0497_),
    .C(_0503_),
    .Y(_0849_));
 sg13g2_a21o_1 _1611_ (.A2(_0848_),
    .A1(_0467_),
    .B1(_0849_),
    .X(_0850_));
 sg13g2_xnor2_1 _1612_ (.Y(_0851_),
    .A(_0474_),
    .B(_0850_));
 sg13g2_nor2_1 _1613_ (.A(net29),
    .B(_0851_),
    .Y(_0852_));
 sg13g2_a21oi_1 _1614_ (.A1(\mux.data_in[8] ),
    .A2(net12),
    .Y(_0853_),
    .B1(_0852_));
 sg13g2_nor2_1 _1615_ (.A(net43),
    .B(_0853_),
    .Y(_0030_));
 sg13g2_nand2_1 _1616_ (.Y(_0854_),
    .A(\mux.data_in[9] ),
    .B(net16));
 sg13g2_a21oi_1 _1617_ (.A1(_0464_),
    .A2(_0850_),
    .Y(_0855_),
    .B1(_0463_));
 sg13g2_nor2_1 _1618_ (.A(_0464_),
    .B(_0850_),
    .Y(_0856_));
 sg13g2_o21ai_1 _1619_ (.B1(_0475_),
    .Y(_0857_),
    .A1(_0855_),
    .A2(_0856_));
 sg13g2_or3_1 _1620_ (.A(_0475_),
    .B(_0855_),
    .C(_0856_),
    .X(_0858_));
 sg13g2_a21o_1 _1621_ (.A2(_0858_),
    .A1(_0857_),
    .B1(net29),
    .X(_0859_));
 sg13g2_a21oi_1 _1622_ (.A1(_0854_),
    .A2(_0859_),
    .Y(_0031_),
    .B1(net44));
 sg13g2_nand2_1 _1623_ (.Y(_0860_),
    .A(\pulse_width_counter_module.high_counter[0] ),
    .B(net26));
 sg13g2_nand2_1 _1624_ (.Y(_0861_),
    .A(\mux.data_in[64] ),
    .B(net12));
 sg13g2_a21oi_1 _1625_ (.A1(_0860_),
    .A2(_0861_),
    .Y(_0032_),
    .B1(net44));
 sg13g2_nand2_1 _1626_ (.Y(_0862_),
    .A(\pulse_width_counter_module.high_counter[10] ),
    .B(net26));
 sg13g2_nand2_1 _1627_ (.Y(_0863_),
    .A(_0507_),
    .B(net12));
 sg13g2_a21oi_1 _1628_ (.A1(_0862_),
    .A2(_0863_),
    .Y(_0033_),
    .B1(net44));
 sg13g2_nand2_1 _1629_ (.Y(_0864_),
    .A(\pulse_width_counter_module.high_counter[11] ),
    .B(net26));
 sg13g2_nand2_1 _1630_ (.Y(_0865_),
    .A(_0520_),
    .B(net12));
 sg13g2_a21oi_1 _1631_ (.A1(_0864_),
    .A2(_0865_),
    .Y(_0034_),
    .B1(net44));
 sg13g2_nand2_1 _1632_ (.Y(_0866_),
    .A(\pulse_width_counter_module.high_counter[12] ),
    .B(net26));
 sg13g2_nand2_1 _1633_ (.Y(_0867_),
    .A(_0534_),
    .B(net12));
 sg13g2_a21oi_1 _1634_ (.A1(_0866_),
    .A2(_0867_),
    .Y(_0035_),
    .B1(net44));
 sg13g2_nand2_1 _1635_ (.Y(_0868_),
    .A(\pulse_width_counter_module.high_counter[13] ),
    .B(net26));
 sg13g2_buf_1 _1636_ (.A(_0455_),
    .X(_0869_));
 sg13g2_nand2_1 _1637_ (.Y(_0870_),
    .A(_0555_),
    .B(net11));
 sg13g2_a21oi_1 _1638_ (.A1(_0868_),
    .A2(_0870_),
    .Y(_0036_),
    .B1(net44));
 sg13g2_nand2_1 _1639_ (.Y(_0871_),
    .A(\pulse_width_counter_module.high_counter[14] ),
    .B(net26));
 sg13g2_nand2_1 _1640_ (.Y(_0872_),
    .A(_0564_),
    .B(net11));
 sg13g2_buf_1 _1641_ (.A(_0524_),
    .X(_0873_));
 sg13g2_a21oi_1 _1642_ (.A1(_0871_),
    .A2(_0872_),
    .Y(_0037_),
    .B1(net42));
 sg13g2_nand2_1 _1643_ (.Y(_0874_),
    .A(\pulse_width_counter_module.high_counter[15] ),
    .B(net26));
 sg13g2_nand2_1 _1644_ (.Y(_0875_),
    .A(_0571_),
    .B(net11));
 sg13g2_a21oi_1 _1645_ (.A1(_0874_),
    .A2(_0875_),
    .Y(_0038_),
    .B1(net42));
 sg13g2_buf_2 _1646_ (.A(\pulse_width_counter_module.high_counter[16] ),
    .X(_0876_));
 sg13g2_nand2_1 _1647_ (.Y(_0877_),
    .A(_0876_),
    .B(net26));
 sg13g2_nand2_1 _1648_ (.Y(_0878_),
    .A(net57),
    .B(net11));
 sg13g2_a21oi_1 _1649_ (.A1(_0877_),
    .A2(_0878_),
    .Y(_0039_),
    .B1(net42));
 sg13g2_buf_1 _1650_ (.A(\pulse_width_counter_module.high_counter[17] ),
    .X(_0879_));
 sg13g2_buf_1 _1651_ (.A(_0450_),
    .X(_0880_));
 sg13g2_nand2_1 _1652_ (.Y(_0881_),
    .A(_0879_),
    .B(net25));
 sg13g2_nand2_1 _1653_ (.Y(_0882_),
    .A(net55),
    .B(net11));
 sg13g2_a21oi_1 _1654_ (.A1(_0881_),
    .A2(_0882_),
    .Y(_0040_),
    .B1(net42));
 sg13g2_nand2_1 _1655_ (.Y(_0883_),
    .A(\pulse_width_counter_module.high_counter[18] ),
    .B(net25));
 sg13g2_nand2_1 _1656_ (.Y(_0884_),
    .A(_0625_),
    .B(_0869_));
 sg13g2_a21oi_1 _1657_ (.A1(_0883_),
    .A2(_0884_),
    .Y(_0041_),
    .B1(_0873_));
 sg13g2_nand2_1 _1658_ (.Y(_0885_),
    .A(\pulse_width_counter_module.high_counter[19] ),
    .B(_0880_));
 sg13g2_nand2_1 _1659_ (.Y(_0886_),
    .A(_0651_),
    .B(net11));
 sg13g2_a21oi_1 _1660_ (.A1(_0885_),
    .A2(_0886_),
    .Y(_0042_),
    .B1(_0873_));
 sg13g2_nand2_1 _1661_ (.Y(_0887_),
    .A(\pulse_width_counter_module.high_counter[1] ),
    .B(net25));
 sg13g2_nand2_1 _1662_ (.Y(_0888_),
    .A(\mux.data_in[65] ),
    .B(net11));
 sg13g2_a21oi_1 _1663_ (.A1(_0887_),
    .A2(_0888_),
    .Y(_0043_),
    .B1(net42));
 sg13g2_nand2_1 _1664_ (.Y(_0889_),
    .A(\pulse_width_counter_module.high_counter[20] ),
    .B(net25));
 sg13g2_nand2_1 _1665_ (.Y(_0890_),
    .A(_0663_),
    .B(net11));
 sg13g2_a21oi_1 _1666_ (.A1(_0889_),
    .A2(_0890_),
    .Y(_0044_),
    .B1(net42));
 sg13g2_nand2_1 _1667_ (.Y(_0891_),
    .A(\pulse_width_counter_module.high_counter[21] ),
    .B(net25));
 sg13g2_nand2_1 _1668_ (.Y(_0892_),
    .A(_0673_),
    .B(_0869_));
 sg13g2_a21oi_1 _1669_ (.A1(_0891_),
    .A2(_0892_),
    .Y(_0045_),
    .B1(net42));
 sg13g2_nand2_1 _1670_ (.Y(_0893_),
    .A(\pulse_width_counter_module.high_counter[22] ),
    .B(net25));
 sg13g2_buf_1 _1671_ (.A(net31),
    .X(_0894_));
 sg13g2_nand2_1 _1672_ (.Y(_0895_),
    .A(\mux.data_in[86] ),
    .B(net10));
 sg13g2_a21oi_1 _1673_ (.A1(_0893_),
    .A2(_0895_),
    .Y(_0046_),
    .B1(net42));
 sg13g2_nand2_1 _1674_ (.Y(_0896_),
    .A(\pulse_width_counter_module.high_counter[23] ),
    .B(net25));
 sg13g2_nand2_1 _1675_ (.Y(_0897_),
    .A(net53),
    .B(net10));
 sg13g2_buf_1 _1676_ (.A(_0524_),
    .X(_0898_));
 sg13g2_a21oi_1 _1677_ (.A1(_0896_),
    .A2(_0897_),
    .Y(_0047_),
    .B1(net41));
 sg13g2_nand2_1 _1678_ (.Y(_0899_),
    .A(\pulse_width_counter_module.high_counter[24] ),
    .B(_0880_));
 sg13g2_nand2_1 _1679_ (.Y(_0900_),
    .A(_0704_),
    .B(net10));
 sg13g2_a21oi_1 _1680_ (.A1(_0899_),
    .A2(_0900_),
    .Y(_0048_),
    .B1(_0898_));
 sg13g2_nand2_1 _1681_ (.Y(_0901_),
    .A(\pulse_width_counter_module.high_counter[25] ),
    .B(net25));
 sg13g2_nand2_1 _1682_ (.Y(_0902_),
    .A(_0718_),
    .B(net10));
 sg13g2_a21oi_1 _1683_ (.A1(_0901_),
    .A2(_0902_),
    .Y(_0049_),
    .B1(net41));
 sg13g2_buf_1 _1684_ (.A(_0450_),
    .X(_0903_));
 sg13g2_nand2_1 _1685_ (.Y(_0904_),
    .A(\pulse_width_counter_module.high_counter[26] ),
    .B(net24));
 sg13g2_nand2_1 _1686_ (.Y(_0905_),
    .A(_0735_),
    .B(_0894_));
 sg13g2_a21oi_1 _1687_ (.A1(_0904_),
    .A2(_0905_),
    .Y(_0050_),
    .B1(net41));
 sg13g2_nand2_1 _1688_ (.Y(_0906_),
    .A(\pulse_width_counter_module.high_counter[27] ),
    .B(net24));
 sg13g2_nand2_1 _1689_ (.Y(_0907_),
    .A(\mux.data_in[91] ),
    .B(net10));
 sg13g2_a21oi_1 _1690_ (.A1(_0906_),
    .A2(_0907_),
    .Y(_0051_),
    .B1(net41));
 sg13g2_nand2_1 _1691_ (.Y(_0908_),
    .A(\pulse_width_counter_module.high_counter[28] ),
    .B(net24));
 sg13g2_nand2_1 _1692_ (.Y(_0909_),
    .A(\mux.data_in[92] ),
    .B(net10));
 sg13g2_a21oi_1 _1693_ (.A1(_0908_),
    .A2(_0909_),
    .Y(_0052_),
    .B1(net41));
 sg13g2_nand2_1 _1694_ (.Y(_0910_),
    .A(\pulse_width_counter_module.high_counter[29] ),
    .B(net24));
 sg13g2_nand2_1 _1695_ (.Y(_0911_),
    .A(\mux.data_in[93] ),
    .B(net10));
 sg13g2_a21oi_1 _1696_ (.A1(_0910_),
    .A2(_0911_),
    .Y(_0053_),
    .B1(net41));
 sg13g2_nand2_1 _1697_ (.Y(_0912_),
    .A(\pulse_width_counter_module.high_counter[2] ),
    .B(net24));
 sg13g2_nand2_1 _1698_ (.Y(_0913_),
    .A(_0480_),
    .B(net10));
 sg13g2_a21oi_1 _1699_ (.A1(_0912_),
    .A2(_0913_),
    .Y(_0054_),
    .B1(net41));
 sg13g2_nand2_1 _1700_ (.Y(_0914_),
    .A(\pulse_width_counter_module.high_counter[30] ),
    .B(_0903_));
 sg13g2_nand2_1 _1701_ (.Y(_0915_),
    .A(\mux.data_in[94] ),
    .B(_0894_));
 sg13g2_a21oi_1 _1702_ (.A1(_0914_),
    .A2(_0915_),
    .Y(_0055_),
    .B1(net41));
 sg13g2_nand2_1 _1703_ (.Y(_0916_),
    .A(\pulse_width_counter_module.high_counter[31] ),
    .B(_0903_));
 sg13g2_nand2_1 _1704_ (.Y(_0917_),
    .A(\mux.data_in[95] ),
    .B(_0724_));
 sg13g2_a21oi_1 _1705_ (.A1(_0916_),
    .A2(_0917_),
    .Y(_0056_),
    .B1(_0898_));
 sg13g2_nand2_1 _1706_ (.Y(_0918_),
    .A(\pulse_width_counter_module.high_counter[3] ),
    .B(net24));
 sg13g2_nand2_1 _1707_ (.Y(_0919_),
    .A(\mux.data_in[67] ),
    .B(net27));
 sg13g2_buf_1 _1708_ (.A(net59),
    .X(_0920_));
 sg13g2_a21oi_1 _1709_ (.A1(_0918_),
    .A2(_0919_),
    .Y(_0057_),
    .B1(net40));
 sg13g2_nand2_1 _1710_ (.Y(_0921_),
    .A(\pulse_width_counter_module.high_counter[4] ),
    .B(net24));
 sg13g2_nand2_1 _1711_ (.Y(_0922_),
    .A(_0487_),
    .B(net27));
 sg13g2_a21oi_1 _1712_ (.A1(_0921_),
    .A2(_0922_),
    .Y(_0058_),
    .B1(net40));
 sg13g2_nand2_1 _1713_ (.Y(_0923_),
    .A(\pulse_width_counter_module.high_counter[5] ),
    .B(net24));
 sg13g2_nand2_1 _1714_ (.Y(_0924_),
    .A(net60),
    .B(net27));
 sg13g2_a21oi_1 _1715_ (.A1(_0923_),
    .A2(_0924_),
    .Y(_0059_),
    .B1(net40));
 sg13g2_nand2_1 _1716_ (.Y(_0925_),
    .A(\pulse_width_counter_module.high_counter[6] ),
    .B(net32));
 sg13g2_nand2_1 _1717_ (.Y(_0926_),
    .A(_0489_),
    .B(net27));
 sg13g2_a21oi_1 _1718_ (.A1(_0925_),
    .A2(_0926_),
    .Y(_0060_),
    .B1(net40));
 sg13g2_nand2_1 _1719_ (.Y(_0927_),
    .A(\pulse_width_counter_module.high_counter[7] ),
    .B(net32));
 sg13g2_nand2_1 _1720_ (.Y(_0928_),
    .A(_0468_),
    .B(net27));
 sg13g2_a21oi_1 _1721_ (.A1(_0927_),
    .A2(_0928_),
    .Y(_0061_),
    .B1(net40));
 sg13g2_nand2_1 _1722_ (.Y(_0929_),
    .A(\pulse_width_counter_module.high_counter[8] ),
    .B(net32));
 sg13g2_nand2_1 _1723_ (.Y(_0930_),
    .A(_0464_),
    .B(net27));
 sg13g2_a21oi_1 _1724_ (.A1(_0929_),
    .A2(_0930_),
    .Y(_0062_),
    .B1(_0920_));
 sg13g2_nand2_1 _1725_ (.Y(_0931_),
    .A(\pulse_width_counter_module.high_counter[9] ),
    .B(net32));
 sg13g2_nand2_1 _1726_ (.Y(_0932_),
    .A(_0461_),
    .B(net27));
 sg13g2_a21oi_1 _1727_ (.A1(_0931_),
    .A2(_0932_),
    .Y(_0063_),
    .B1(net40));
 sg13g2_nor2b_1 _1728_ (.A(_0448_),
    .B_N(_0447_),
    .Y(_0933_));
 sg13g2_buf_2 _1729_ (.A(_0933_),
    .X(_0934_));
 sg13g2_buf_1 _1730_ (.A(_0934_),
    .X(_0935_));
 sg13g2_nand2_1 _1731_ (.Y(_0936_),
    .A(\pulse_width_counter_module.low_counter[0] ),
    .B(_0935_));
 sg13g2_buf_1 _1732_ (.A(_0447_),
    .X(_0937_));
 sg13g2_nand2b_1 _1733_ (.Y(_0938_),
    .B(net51),
    .A_N(_0448_));
 sg13g2_buf_1 _1734_ (.A(_0938_),
    .X(_0939_));
 sg13g2_buf_1 _1735_ (.A(net34),
    .X(_0940_));
 sg13g2_nand2_1 _1736_ (.Y(_0941_),
    .A(\mux.data_in[32] ),
    .B(net22));
 sg13g2_a21oi_1 _1737_ (.A1(_0936_),
    .A2(_0941_),
    .Y(_0064_),
    .B1(net40));
 sg13g2_nand2_1 _1738_ (.Y(_0942_),
    .A(\pulse_width_counter_module.low_counter[10] ),
    .B(net23));
 sg13g2_nand2_1 _1739_ (.Y(_0943_),
    .A(_0506_),
    .B(_0940_));
 sg13g2_a21oi_1 _1740_ (.A1(_0942_),
    .A2(_0943_),
    .Y(_0065_),
    .B1(net40));
 sg13g2_nand2_1 _1741_ (.Y(_0944_),
    .A(\pulse_width_counter_module.low_counter[11] ),
    .B(net23));
 sg13g2_nand2_1 _1742_ (.Y(_0945_),
    .A(_0519_),
    .B(_0940_));
 sg13g2_a21oi_1 _1743_ (.A1(_0944_),
    .A2(_0945_),
    .Y(_0066_),
    .B1(_0920_));
 sg13g2_nand2_1 _1744_ (.Y(_0946_),
    .A(\pulse_width_counter_module.low_counter[12] ),
    .B(net23));
 sg13g2_nand2_1 _1745_ (.Y(_0947_),
    .A(_0533_),
    .B(net22));
 sg13g2_buf_1 _1746_ (.A(net59),
    .X(_0948_));
 sg13g2_a21oi_1 _1747_ (.A1(_0946_),
    .A2(_0947_),
    .Y(_0067_),
    .B1(net39));
 sg13g2_nand2_1 _1748_ (.Y(_0949_),
    .A(\pulse_width_counter_module.low_counter[13] ),
    .B(net23));
 sg13g2_nand2_1 _1749_ (.Y(_0950_),
    .A(_0554_),
    .B(net22));
 sg13g2_a21oi_1 _1750_ (.A1(_0949_),
    .A2(_0950_),
    .Y(_0068_),
    .B1(net39));
 sg13g2_nand2_1 _1751_ (.Y(_0951_),
    .A(\pulse_width_counter_module.low_counter[14] ),
    .B(net23));
 sg13g2_nand2_1 _1752_ (.Y(_0952_),
    .A(_0563_),
    .B(net22));
 sg13g2_a21oi_1 _1753_ (.A1(_0951_),
    .A2(_0952_),
    .Y(_0069_),
    .B1(net39));
 sg13g2_buf_1 _1754_ (.A(\pulse_width_counter_module.low_counter[15] ),
    .X(_0953_));
 sg13g2_nand2_1 _1755_ (.Y(_0954_),
    .A(_0953_),
    .B(net23));
 sg13g2_nand2_1 _1756_ (.Y(_0955_),
    .A(_0570_),
    .B(net22));
 sg13g2_a21oi_1 _1757_ (.A1(_0954_),
    .A2(_0955_),
    .Y(_0070_),
    .B1(net39));
 sg13g2_nand2_1 _1758_ (.Y(_0956_),
    .A(\pulse_width_counter_module.low_counter[16] ),
    .B(net23));
 sg13g2_nand2_1 _1759_ (.Y(_0957_),
    .A(_0582_),
    .B(net22));
 sg13g2_a21oi_1 _1760_ (.A1(_0956_),
    .A2(_0957_),
    .Y(_0071_),
    .B1(net39));
 sg13g2_nand2_1 _1761_ (.Y(_0958_),
    .A(\pulse_width_counter_module.low_counter[17] ),
    .B(_0935_));
 sg13g2_nand2_1 _1762_ (.Y(_0959_),
    .A(_0603_),
    .B(net22));
 sg13g2_a21oi_1 _1763_ (.A1(_0958_),
    .A2(_0959_),
    .Y(_0072_),
    .B1(net39));
 sg13g2_nand2_1 _1764_ (.Y(_0960_),
    .A(\pulse_width_counter_module.low_counter[18] ),
    .B(net23));
 sg13g2_nand2_1 _1765_ (.Y(_0961_),
    .A(\mux.data_in[50] ),
    .B(net22));
 sg13g2_a21oi_1 _1766_ (.A1(_0960_),
    .A2(_0961_),
    .Y(_0073_),
    .B1(net39));
 sg13g2_buf_1 _1767_ (.A(_0934_),
    .X(_0962_));
 sg13g2_nand2_1 _1768_ (.Y(_0963_),
    .A(\pulse_width_counter_module.low_counter[19] ),
    .B(net21));
 sg13g2_buf_1 _1769_ (.A(net34),
    .X(_0964_));
 sg13g2_nand2_1 _1770_ (.Y(_0965_),
    .A(_0650_),
    .B(net20));
 sg13g2_a21oi_1 _1771_ (.A1(_0963_),
    .A2(_0965_),
    .Y(_0074_),
    .B1(net39));
 sg13g2_nand2_1 _1772_ (.Y(_0966_),
    .A(\pulse_width_counter_module.low_counter[1] ),
    .B(net21));
 sg13g2_nand2_1 _1773_ (.Y(_0967_),
    .A(\mux.data_in[33] ),
    .B(net20));
 sg13g2_a21oi_1 _1774_ (.A1(_0966_),
    .A2(_0967_),
    .Y(_0075_),
    .B1(_0948_));
 sg13g2_nand2_1 _1775_ (.Y(_0968_),
    .A(\pulse_width_counter_module.low_counter[20] ),
    .B(net21));
 sg13g2_nand2_1 _1776_ (.Y(_0969_),
    .A(_0662_),
    .B(net20));
 sg13g2_a21oi_1 _1777_ (.A1(_0968_),
    .A2(_0969_),
    .Y(_0076_),
    .B1(_0948_));
 sg13g2_buf_1 _1778_ (.A(\pulse_width_counter_module.low_counter[21] ),
    .X(_0970_));
 sg13g2_nand2_1 _1779_ (.Y(_0971_),
    .A(_0970_),
    .B(net21));
 sg13g2_nand2_1 _1780_ (.Y(_0972_),
    .A(_0672_),
    .B(net20));
 sg13g2_buf_1 _1781_ (.A(net59),
    .X(_0973_));
 sg13g2_a21oi_1 _1782_ (.A1(_0971_),
    .A2(_0972_),
    .Y(_0077_),
    .B1(net38));
 sg13g2_nand2_1 _1783_ (.Y(_0974_),
    .A(\pulse_width_counter_module.low_counter[22] ),
    .B(net21));
 sg13g2_nand2_1 _1784_ (.Y(_0975_),
    .A(_0677_),
    .B(net20));
 sg13g2_a21oi_1 _1785_ (.A1(_0974_),
    .A2(_0975_),
    .Y(_0078_),
    .B1(net38));
 sg13g2_nand2_1 _1786_ (.Y(_0976_),
    .A(\pulse_width_counter_module.low_counter[23] ),
    .B(net21));
 sg13g2_nand2_1 _1787_ (.Y(_0977_),
    .A(net54),
    .B(net20));
 sg13g2_a21oi_1 _1788_ (.A1(_0976_),
    .A2(_0977_),
    .Y(_0079_),
    .B1(net38));
 sg13g2_nand2_1 _1789_ (.Y(_0978_),
    .A(\pulse_width_counter_module.low_counter[24] ),
    .B(net21));
 sg13g2_nand2_1 _1790_ (.Y(_0979_),
    .A(_0703_),
    .B(net20));
 sg13g2_a21oi_1 _1791_ (.A1(_0978_),
    .A2(_0979_),
    .Y(_0080_),
    .B1(net38));
 sg13g2_nand2_1 _1792_ (.Y(_0980_),
    .A(\pulse_width_counter_module.low_counter[25] ),
    .B(net21));
 sg13g2_nand2_1 _1793_ (.Y(_0981_),
    .A(_0717_),
    .B(net20));
 sg13g2_a21oi_1 _1794_ (.A1(_0980_),
    .A2(_0981_),
    .Y(_0081_),
    .B1(net38));
 sg13g2_nand2_1 _1795_ (.Y(_0982_),
    .A(\pulse_width_counter_module.low_counter[26] ),
    .B(_0962_));
 sg13g2_nand2_1 _1796_ (.Y(_0983_),
    .A(_0734_),
    .B(_0964_));
 sg13g2_a21oi_1 _1797_ (.A1(_0982_),
    .A2(_0983_),
    .Y(_0082_),
    .B1(_0973_));
 sg13g2_nand2_1 _1798_ (.Y(_0984_),
    .A(\pulse_width_counter_module.low_counter[27] ),
    .B(_0962_));
 sg13g2_nand2_1 _1799_ (.Y(_0985_),
    .A(\mux.data_in[59] ),
    .B(_0964_));
 sg13g2_a21oi_1 _1800_ (.A1(_0984_),
    .A2(_0985_),
    .Y(_0083_),
    .B1(net38));
 sg13g2_buf_1 _1801_ (.A(_0934_),
    .X(_0986_));
 sg13g2_nand2_1 _1802_ (.Y(_0987_),
    .A(\pulse_width_counter_module.low_counter[28] ),
    .B(net19));
 sg13g2_buf_1 _1803_ (.A(net34),
    .X(_0988_));
 sg13g2_nand2_1 _1804_ (.Y(_0989_),
    .A(\mux.data_in[60] ),
    .B(net18));
 sg13g2_a21oi_1 _1805_ (.A1(_0987_),
    .A2(_0989_),
    .Y(_0084_),
    .B1(net38));
 sg13g2_nand2_1 _1806_ (.Y(_0990_),
    .A(\pulse_width_counter_module.low_counter[29] ),
    .B(net19));
 sg13g2_nand2_1 _1807_ (.Y(_0991_),
    .A(\mux.data_in[61] ),
    .B(net18));
 sg13g2_a21oi_1 _1808_ (.A1(_0990_),
    .A2(_0991_),
    .Y(_0085_),
    .B1(_0973_));
 sg13g2_nand2_1 _1809_ (.Y(_0992_),
    .A(\pulse_width_counter_module.low_counter[2] ),
    .B(net19));
 sg13g2_nand2_1 _1810_ (.Y(_0993_),
    .A(\mux.data_in[34] ),
    .B(net18));
 sg13g2_a21oi_1 _1811_ (.A1(_0992_),
    .A2(_0993_),
    .Y(_0086_),
    .B1(net38));
 sg13g2_nand2_1 _1812_ (.Y(_0994_),
    .A(\pulse_width_counter_module.low_counter[30] ),
    .B(_0986_));
 sg13g2_nand2_1 _1813_ (.Y(_0995_),
    .A(\mux.data_in[62] ),
    .B(_0988_));
 sg13g2_buf_1 _1814_ (.A(net59),
    .X(_0996_));
 sg13g2_a21oi_1 _1815_ (.A1(_0994_),
    .A2(_0995_),
    .Y(_0087_),
    .B1(net37));
 sg13g2_nand2_1 _1816_ (.Y(_0997_),
    .A(\pulse_width_counter_module.low_counter[31] ),
    .B(net19));
 sg13g2_nand2_1 _1817_ (.Y(_0998_),
    .A(\mux.data_in[63] ),
    .B(net18));
 sg13g2_a21oi_1 _1818_ (.A1(_0997_),
    .A2(_0998_),
    .Y(_0088_),
    .B1(net37));
 sg13g2_nand2_1 _1819_ (.Y(_0999_),
    .A(\pulse_width_counter_module.low_counter[3] ),
    .B(net19));
 sg13g2_nand2_1 _1820_ (.Y(_1000_),
    .A(\mux.data_in[35] ),
    .B(net18));
 sg13g2_a21oi_1 _1821_ (.A1(_0999_),
    .A2(_1000_),
    .Y(_0089_),
    .B1(net37));
 sg13g2_nand2_1 _1822_ (.Y(_1001_),
    .A(\pulse_width_counter_module.low_counter[4] ),
    .B(net19));
 sg13g2_nand2_1 _1823_ (.Y(_1002_),
    .A(_0486_),
    .B(net18));
 sg13g2_a21oi_1 _1824_ (.A1(_1001_),
    .A2(_1002_),
    .Y(_0090_),
    .B1(net37));
 sg13g2_nand2_1 _1825_ (.Y(_1003_),
    .A(\pulse_width_counter_module.low_counter[5] ),
    .B(_0986_));
 sg13g2_nand2_1 _1826_ (.Y(_1004_),
    .A(_0491_),
    .B(_0988_));
 sg13g2_a21oi_1 _1827_ (.A1(_1003_),
    .A2(_1004_),
    .Y(_0091_),
    .B1(_0996_));
 sg13g2_nand2_1 _1828_ (.Y(_1005_),
    .A(\pulse_width_counter_module.low_counter[6] ),
    .B(net19));
 sg13g2_nand2_1 _1829_ (.Y(_1006_),
    .A(_0493_),
    .B(net18));
 sg13g2_a21oi_1 _1830_ (.A1(_1005_),
    .A2(_1006_),
    .Y(_0092_),
    .B1(_0996_));
 sg13g2_nand2_1 _1831_ (.Y(_1007_),
    .A(\pulse_width_counter_module.low_counter[7] ),
    .B(net19));
 sg13g2_nand2_1 _1832_ (.Y(_1008_),
    .A(_0467_),
    .B(net18));
 sg13g2_a21oi_1 _1833_ (.A1(_1007_),
    .A2(_1008_),
    .Y(_0093_),
    .B1(net37));
 sg13g2_nand2_1 _1834_ (.Y(_1009_),
    .A(\pulse_width_counter_module.low_counter[8] ),
    .B(_0934_));
 sg13g2_buf_1 _1835_ (.A(net34),
    .X(_1010_));
 sg13g2_nand2_1 _1836_ (.Y(_1011_),
    .A(_0463_),
    .B(net17));
 sg13g2_a21oi_1 _1837_ (.A1(_1009_),
    .A2(_1011_),
    .Y(_0094_),
    .B1(net37));
 sg13g2_nand2_1 _1838_ (.Y(_1012_),
    .A(\pulse_width_counter_module.low_counter[9] ),
    .B(_0934_));
 sg13g2_nand2_1 _1839_ (.Y(_0161_),
    .A(_0460_),
    .B(net17));
 sg13g2_a21oi_1 _1840_ (.A1(_1012_),
    .A2(_0161_),
    .Y(_0095_),
    .B1(net37));
 sg13g2_nand2_2 _1841_ (.Y(_0162_),
    .A(net63),
    .B(net29));
 sg13g2_xnor2_1 _1842_ (.Y(_0163_),
    .A(net51),
    .B(\pulse_width_counter_module.high_counter[0] ));
 sg13g2_nor2_1 _1843_ (.A(_0162_),
    .B(_0163_),
    .Y(_0096_));
 sg13g2_nand2_1 _1844_ (.Y(_0164_),
    .A(\pulse_width_counter_module.high_counter[10] ),
    .B(net28));
 sg13g2_and4_1 _1845_ (.A(_0447_),
    .B(\pulse_width_counter_module.high_counter[0] ),
    .C(\pulse_width_counter_module.high_counter[1] ),
    .D(\pulse_width_counter_module.high_counter[2] ),
    .X(_0165_));
 sg13g2_buf_1 _1846_ (.A(_0165_),
    .X(_0166_));
 sg13g2_and4_1 _1847_ (.A(\pulse_width_counter_module.high_counter[3] ),
    .B(\pulse_width_counter_module.high_counter[4] ),
    .C(\pulse_width_counter_module.high_counter[5] ),
    .D(_0166_),
    .X(_0167_));
 sg13g2_and2_1 _1848_ (.A(\pulse_width_counter_module.high_counter[6] ),
    .B(_0167_),
    .X(_0168_));
 sg13g2_buf_1 _1849_ (.A(_0168_),
    .X(_0169_));
 sg13g2_and3_1 _1850_ (.X(_0170_),
    .A(\pulse_width_counter_module.high_counter[7] ),
    .B(\pulse_width_counter_module.high_counter[8] ),
    .C(\pulse_width_counter_module.high_counter[9] ));
 sg13g2_nand2_1 _1851_ (.Y(_0171_),
    .A(_0169_),
    .B(_0170_));
 sg13g2_mux2_1 _1852_ (.A0(\pulse_width_counter_module.high_counter[10] ),
    .A1(_0164_),
    .S(_0171_),
    .X(_0172_));
 sg13g2_nor2_1 _1853_ (.A(net43),
    .B(_0172_),
    .Y(_0097_));
 sg13g2_nand4_1 _1854_ (.B(\pulse_width_counter_module.high_counter[10] ),
    .C(_0167_),
    .A(\pulse_width_counter_module.high_counter[6] ),
    .Y(_0173_),
    .D(_0170_));
 sg13g2_buf_2 _1855_ (.A(_0173_),
    .X(_0174_));
 sg13g2_nand3_1 _1856_ (.B(net27),
    .C(_0174_),
    .A(\pulse_width_counter_module.high_counter[11] ),
    .Y(_0175_));
 sg13g2_inv_1 _1857_ (.Y(_0176_),
    .A(\pulse_width_counter_module.high_counter[11] ));
 sg13g2_nand2b_1 _1858_ (.Y(_0177_),
    .B(_0176_),
    .A_N(_0174_));
 sg13g2_a21oi_1 _1859_ (.A1(_0175_),
    .A2(_0177_),
    .Y(_0098_),
    .B1(net37));
 sg13g2_nor2_1 _1860_ (.A(_0176_),
    .B(_0174_),
    .Y(_0178_));
 sg13g2_xnor2_1 _1861_ (.Y(_0179_),
    .A(\pulse_width_counter_module.high_counter[12] ),
    .B(_0178_));
 sg13g2_nor2_1 _1862_ (.A(_0162_),
    .B(_0179_),
    .Y(_0099_));
 sg13g2_nand2_1 _1863_ (.Y(_0180_),
    .A(\pulse_width_counter_module.high_counter[13] ),
    .B(net28));
 sg13g2_nand2_1 _1864_ (.Y(_0181_),
    .A(\pulse_width_counter_module.high_counter[11] ),
    .B(\pulse_width_counter_module.high_counter[12] ));
 sg13g2_nor2_1 _1865_ (.A(_0174_),
    .B(_0181_),
    .Y(_0182_));
 sg13g2_mux2_1 _1866_ (.A0(_0180_),
    .A1(\pulse_width_counter_module.high_counter[13] ),
    .S(_0182_),
    .X(_0183_));
 sg13g2_nor2_1 _1867_ (.A(net43),
    .B(_0183_),
    .Y(_0100_));
 sg13g2_nand2_1 _1868_ (.Y(_0184_),
    .A(\pulse_width_counter_module.high_counter[14] ),
    .B(net28));
 sg13g2_nand2_1 _1869_ (.Y(_0185_),
    .A(\pulse_width_counter_module.high_counter[13] ),
    .B(_0182_));
 sg13g2_mux2_1 _1870_ (.A0(\pulse_width_counter_module.high_counter[14] ),
    .A1(_0184_),
    .S(_0185_),
    .X(_0186_));
 sg13g2_nor2_1 _1871_ (.A(net43),
    .B(_0186_),
    .Y(_0101_));
 sg13g2_inv_1 _1872_ (.Y(_0187_),
    .A(\pulse_width_counter_module.high_counter[15] ));
 sg13g2_nand2_1 _1873_ (.Y(_0188_),
    .A(\pulse_width_counter_module.high_counter[13] ),
    .B(\pulse_width_counter_module.high_counter[14] ));
 sg13g2_nor3_1 _1874_ (.A(_0174_),
    .B(_0181_),
    .C(_0188_),
    .Y(_0189_));
 sg13g2_nor3_1 _1875_ (.A(_0187_),
    .B(_0512_),
    .C(_0189_),
    .Y(_0190_));
 sg13g2_a21oi_1 _1876_ (.A1(_0187_),
    .A2(_0189_),
    .Y(_0191_),
    .B1(_0190_));
 sg13g2_nor2_1 _1877_ (.A(net43),
    .B(_0191_),
    .Y(_0102_));
 sg13g2_nor4_2 _1878_ (.A(_0187_),
    .B(_0174_),
    .C(_0181_),
    .Y(_0192_),
    .D(_0188_));
 sg13g2_nand3b_1 _1879_ (.B(_0876_),
    .C(net29),
    .Y(_0193_),
    .A_N(_0192_));
 sg13g2_nand2b_1 _1880_ (.Y(_0194_),
    .B(_0192_),
    .A_N(_0876_));
 sg13g2_buf_1 _1881_ (.A(net59),
    .X(_0195_));
 sg13g2_a21oi_1 _1882_ (.A1(_0193_),
    .A2(_0194_),
    .Y(_0103_),
    .B1(net36));
 sg13g2_nand2_1 _1883_ (.Y(_0196_),
    .A(_0876_),
    .B(_0192_));
 sg13g2_nand3_1 _1884_ (.B(net31),
    .C(_0196_),
    .A(_0879_),
    .Y(_0197_));
 sg13g2_o21ai_1 _1885_ (.B1(_0197_),
    .Y(_0198_),
    .A1(_0879_),
    .A2(_0196_));
 sg13g2_and2_1 _1886_ (.A(_0568_),
    .B(_0198_),
    .X(_0104_));
 sg13g2_nand3_1 _1887_ (.B(_0879_),
    .C(_0192_),
    .A(_0876_),
    .Y(_0199_));
 sg13g2_buf_2 _1888_ (.A(_0199_),
    .X(_0200_));
 sg13g2_nand3_1 _1889_ (.B(net31),
    .C(_0200_),
    .A(\pulse_width_counter_module.high_counter[18] ),
    .Y(_0201_));
 sg13g2_o21ai_1 _1890_ (.B1(_0201_),
    .Y(_0202_),
    .A1(\pulse_width_counter_module.high_counter[18] ),
    .A2(_0200_));
 sg13g2_and2_1 _1891_ (.A(net58),
    .B(_0202_),
    .X(_0105_));
 sg13g2_nand2_1 _1892_ (.Y(_0203_),
    .A(\pulse_width_counter_module.high_counter[19] ),
    .B(net28));
 sg13g2_nand4_1 _1893_ (.B(_0879_),
    .C(\pulse_width_counter_module.high_counter[18] ),
    .A(_0876_),
    .Y(_0204_),
    .D(_0192_));
 sg13g2_mux2_1 _1894_ (.A0(\pulse_width_counter_module.high_counter[19] ),
    .A1(_0203_),
    .S(_0204_),
    .X(_0205_));
 sg13g2_nor2_1 _1895_ (.A(net43),
    .B(_0205_),
    .Y(_0106_));
 sg13g2_nand2_1 _1896_ (.Y(_0206_),
    .A(net51),
    .B(\pulse_width_counter_module.high_counter[0] ));
 sg13g2_xor2_1 _1897_ (.B(_0206_),
    .A(\pulse_width_counter_module.high_counter[1] ),
    .X(_0207_));
 sg13g2_nor2_1 _1898_ (.A(_0162_),
    .B(_0207_),
    .Y(_0107_));
 sg13g2_nand2_1 _1899_ (.Y(_0208_),
    .A(\pulse_width_counter_module.high_counter[20] ),
    .B(net28));
 sg13g2_nand2_1 _1900_ (.Y(_0209_),
    .A(\pulse_width_counter_module.high_counter[18] ),
    .B(\pulse_width_counter_module.high_counter[19] ));
 sg13g2_nor2_1 _1901_ (.A(_0200_),
    .B(_0209_),
    .Y(_0210_));
 sg13g2_mux2_1 _1902_ (.A0(_0208_),
    .A1(\pulse_width_counter_module.high_counter[20] ),
    .S(_0210_),
    .X(_0211_));
 sg13g2_nor2_1 _1903_ (.A(net43),
    .B(_0211_),
    .Y(_0108_));
 sg13g2_nand2_1 _1904_ (.Y(_0212_),
    .A(\pulse_width_counter_module.high_counter[20] ),
    .B(_0210_));
 sg13g2_nand3_1 _1905_ (.B(net29),
    .C(_0212_),
    .A(\pulse_width_counter_module.high_counter[21] ),
    .Y(_0213_));
 sg13g2_or2_1 _1906_ (.X(_0214_),
    .B(_0212_),
    .A(\pulse_width_counter_module.high_counter[21] ));
 sg13g2_a21oi_1 _1907_ (.A1(_0213_),
    .A2(_0214_),
    .Y(_0109_),
    .B1(net36));
 sg13g2_nand2_1 _1908_ (.Y(_0215_),
    .A(\pulse_width_counter_module.high_counter[22] ),
    .B(net28));
 sg13g2_nand3_1 _1909_ (.B(\pulse_width_counter_module.high_counter[21] ),
    .C(_0210_),
    .A(\pulse_width_counter_module.high_counter[20] ),
    .Y(_0216_));
 sg13g2_mux2_1 _1910_ (.A0(\pulse_width_counter_module.high_counter[22] ),
    .A1(_0215_),
    .S(_0216_),
    .X(_0217_));
 sg13g2_nor2_1 _1911_ (.A(net43),
    .B(_0217_),
    .Y(_0110_));
 sg13g2_nand3_1 _1912_ (.B(\pulse_width_counter_module.high_counter[21] ),
    .C(\pulse_width_counter_module.high_counter[22] ),
    .A(\pulse_width_counter_module.high_counter[20] ),
    .Y(_0218_));
 sg13g2_or2_1 _1913_ (.X(_0219_),
    .B(_0218_),
    .A(_0209_));
 sg13g2_and2_1 _1914_ (.A(\pulse_width_counter_module.high_counter[23] ),
    .B(_0454_),
    .X(_0220_));
 sg13g2_o21ai_1 _1915_ (.B1(_0220_),
    .Y(_0221_),
    .A1(_0200_),
    .A2(_0219_));
 sg13g2_or3_1 _1916_ (.A(\pulse_width_counter_module.high_counter[23] ),
    .B(_0200_),
    .C(_0219_),
    .X(_0222_));
 sg13g2_a21oi_1 _1917_ (.A1(_0221_),
    .A2(_0222_),
    .Y(_0111_),
    .B1(net36));
 sg13g2_nand2_1 _1918_ (.Y(_0223_),
    .A(\pulse_width_counter_module.high_counter[24] ),
    .B(net31));
 sg13g2_nand2_1 _1919_ (.Y(_0224_),
    .A(_0879_),
    .B(\pulse_width_counter_module.high_counter[23] ));
 sg13g2_nor2_1 _1920_ (.A(_0219_),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_nand3_1 _1921_ (.B(_0192_),
    .C(_0225_),
    .A(_0876_),
    .Y(_0226_));
 sg13g2_mux2_1 _1922_ (.A0(\pulse_width_counter_module.high_counter[24] ),
    .A1(_0223_),
    .S(_0226_),
    .X(_0227_));
 sg13g2_nor2_1 _1923_ (.A(_0846_),
    .B(_0227_),
    .Y(_0112_));
 sg13g2_nand4_1 _1924_ (.B(\pulse_width_counter_module.high_counter[24] ),
    .C(_0192_),
    .A(_0876_),
    .Y(_0228_),
    .D(_0225_));
 sg13g2_buf_2 _1925_ (.A(_0228_),
    .X(_0229_));
 sg13g2_nand3_1 _1926_ (.B(net29),
    .C(_0229_),
    .A(\pulse_width_counter_module.high_counter[25] ),
    .Y(_0230_));
 sg13g2_or2_1 _1927_ (.X(_0231_),
    .B(_0229_),
    .A(\pulse_width_counter_module.high_counter[25] ));
 sg13g2_a21oi_1 _1928_ (.A1(_0230_),
    .A2(_0231_),
    .Y(_0113_),
    .B1(net36));
 sg13g2_inv_1 _1929_ (.Y(_0232_),
    .A(_0229_));
 sg13g2_nand2_1 _1930_ (.Y(_0233_),
    .A(\pulse_width_counter_module.high_counter[25] ),
    .B(_0232_));
 sg13g2_nand3_1 _1931_ (.B(net29),
    .C(_0233_),
    .A(\pulse_width_counter_module.high_counter[26] ),
    .Y(_0234_));
 sg13g2_or2_1 _1932_ (.X(_0235_),
    .B(_0233_),
    .A(\pulse_width_counter_module.high_counter[26] ));
 sg13g2_a21oi_1 _1933_ (.A1(_0234_),
    .A2(_0235_),
    .Y(_0114_),
    .B1(net36));
 sg13g2_nand2_1 _1934_ (.Y(_0236_),
    .A(\pulse_width_counter_module.high_counter[27] ),
    .B(_0579_));
 sg13g2_nand2_1 _1935_ (.Y(_0237_),
    .A(\pulse_width_counter_module.high_counter[25] ),
    .B(\pulse_width_counter_module.high_counter[26] ));
 sg13g2_nor2_1 _1936_ (.A(_0229_),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_mux2_1 _1937_ (.A0(_0236_),
    .A1(\pulse_width_counter_module.high_counter[27] ),
    .S(_0238_),
    .X(_0239_));
 sg13g2_nor2_1 _1938_ (.A(_0846_),
    .B(_0239_),
    .Y(_0115_));
 sg13g2_nand2_1 _1939_ (.Y(_0240_),
    .A(\pulse_width_counter_module.high_counter[27] ),
    .B(_0238_));
 sg13g2_nand3_1 _1940_ (.B(_0569_),
    .C(_0240_),
    .A(\pulse_width_counter_module.high_counter[28] ),
    .Y(_0241_));
 sg13g2_or2_1 _1941_ (.X(_0242_),
    .B(_0240_),
    .A(\pulse_width_counter_module.high_counter[28] ));
 sg13g2_a21oi_1 _1942_ (.A1(_0241_),
    .A2(_0242_),
    .Y(_0116_),
    .B1(_0195_));
 sg13g2_nand2_1 _1943_ (.Y(_0243_),
    .A(\pulse_width_counter_module.high_counter[29] ),
    .B(_0579_));
 sg13g2_nand2_1 _1944_ (.Y(_0244_),
    .A(\pulse_width_counter_module.high_counter[27] ),
    .B(\pulse_width_counter_module.high_counter[28] ));
 sg13g2_nor3_2 _1945_ (.A(_0229_),
    .B(_0237_),
    .C(_0244_),
    .Y(_0245_));
 sg13g2_mux2_1 _1946_ (.A0(_0243_),
    .A1(\pulse_width_counter_module.high_counter[29] ),
    .S(_0245_),
    .X(_0246_));
 sg13g2_nor2_1 _1947_ (.A(_0525_),
    .B(_0246_),
    .Y(_0117_));
 sg13g2_nand2_1 _1948_ (.Y(_0247_),
    .A(\pulse_width_counter_module.high_counter[0] ),
    .B(\pulse_width_counter_module.high_counter[1] ));
 sg13g2_xnor2_1 _1949_ (.Y(_0248_),
    .A(\pulse_width_counter_module.high_counter[2] ),
    .B(_0247_));
 sg13g2_nor2_1 _1950_ (.A(_0448_),
    .B(_0937_),
    .Y(_0249_));
 sg13g2_a22oi_1 _1951_ (.Y(_0250_),
    .B1(_0249_),
    .B2(\pulse_width_counter_module.high_counter[2] ),
    .A2(_0248_),
    .A1(_0937_));
 sg13g2_nor2_1 _1952_ (.A(net45),
    .B(_0250_),
    .Y(_0118_));
 sg13g2_nand2_1 _1953_ (.Y(_0251_),
    .A(\pulse_width_counter_module.high_counter[29] ),
    .B(_0245_));
 sg13g2_nand3_1 _1954_ (.B(_0569_),
    .C(_0251_),
    .A(\pulse_width_counter_module.high_counter[30] ),
    .Y(_0252_));
 sg13g2_or2_1 _1955_ (.X(_0253_),
    .B(_0251_),
    .A(\pulse_width_counter_module.high_counter[30] ));
 sg13g2_a21oi_1 _1956_ (.A1(_0252_),
    .A2(_0253_),
    .Y(_0119_),
    .B1(_0195_));
 sg13g2_nand3_1 _1957_ (.B(\pulse_width_counter_module.high_counter[30] ),
    .C(_0245_),
    .A(\pulse_width_counter_module.high_counter[29] ),
    .Y(_0254_));
 sg13g2_nand2b_1 _1958_ (.Y(_0255_),
    .B(_0592_),
    .A_N(\pulse_width_counter_module.high_counter[31] ));
 sg13g2_nand3_1 _1959_ (.B(net13),
    .C(_0254_),
    .A(\pulse_width_counter_module.high_counter[31] ),
    .Y(_0256_));
 sg13g2_o21ai_1 _1960_ (.B1(_0256_),
    .Y(_0120_),
    .A1(_0254_),
    .A2(_0255_));
 sg13g2_xnor2_1 _1961_ (.Y(_0257_),
    .A(\pulse_width_counter_module.high_counter[3] ),
    .B(_0166_));
 sg13g2_nor2_1 _1962_ (.A(_0162_),
    .B(_0257_),
    .Y(_0121_));
 sg13g2_nand2_1 _1963_ (.Y(_0258_),
    .A(\pulse_width_counter_module.high_counter[3] ),
    .B(_0166_));
 sg13g2_nand3_1 _1964_ (.B(net31),
    .C(_0258_),
    .A(\pulse_width_counter_module.high_counter[4] ),
    .Y(_0259_));
 sg13g2_o21ai_1 _1965_ (.B1(_0259_),
    .Y(_0260_),
    .A1(\pulse_width_counter_module.high_counter[4] ),
    .A2(_0258_));
 sg13g2_and2_1 _1966_ (.A(net58),
    .B(_0260_),
    .X(_0122_));
 sg13g2_nand3_1 _1967_ (.B(\pulse_width_counter_module.high_counter[4] ),
    .C(_0166_),
    .A(\pulse_width_counter_module.high_counter[3] ),
    .Y(_0261_));
 sg13g2_nand3_1 _1968_ (.B(net31),
    .C(_0261_),
    .A(\pulse_width_counter_module.high_counter[5] ),
    .Y(_0262_));
 sg13g2_o21ai_1 _1969_ (.B1(_0262_),
    .Y(_0263_),
    .A1(\pulse_width_counter_module.high_counter[5] ),
    .A2(_0261_));
 sg13g2_and2_1 _1970_ (.A(net58),
    .B(_0263_),
    .X(_0123_));
 sg13g2_xnor2_1 _1971_ (.Y(_0264_),
    .A(\pulse_width_counter_module.high_counter[6] ),
    .B(_0167_));
 sg13g2_nor2_1 _1972_ (.A(_0162_),
    .B(_0264_),
    .Y(_0124_));
 sg13g2_nand2_1 _1973_ (.Y(_0265_),
    .A(\pulse_width_counter_module.high_counter[7] ),
    .B(net28));
 sg13g2_mux2_1 _1974_ (.A0(_0265_),
    .A1(\pulse_width_counter_module.high_counter[7] ),
    .S(_0169_),
    .X(_0266_));
 sg13g2_nor2_1 _1975_ (.A(net45),
    .B(_0266_),
    .Y(_0125_));
 sg13g2_nand2_1 _1976_ (.Y(_0267_),
    .A(\pulse_width_counter_module.high_counter[7] ),
    .B(_0169_));
 sg13g2_nand3_1 _1977_ (.B(net31),
    .C(_0267_),
    .A(\pulse_width_counter_module.high_counter[8] ),
    .Y(_0268_));
 sg13g2_o21ai_1 _1978_ (.B1(_0268_),
    .Y(_0269_),
    .A1(\pulse_width_counter_module.high_counter[8] ),
    .A2(_0267_));
 sg13g2_and2_1 _1979_ (.A(net58),
    .B(_0269_),
    .X(_0126_));
 sg13g2_nand3_1 _1980_ (.B(\pulse_width_counter_module.high_counter[8] ),
    .C(_0169_),
    .A(\pulse_width_counter_module.high_counter[7] ),
    .Y(_0270_));
 sg13g2_xor2_1 _1981_ (.B(_0270_),
    .A(\pulse_width_counter_module.high_counter[9] ),
    .X(_0271_));
 sg13g2_nor2_1 _1982_ (.A(_0162_),
    .B(_0271_),
    .Y(_0127_));
 sg13g2_nand3_1 _1983_ (.B(net51),
    .C(\pulse_width_counter_module.low_counter[0] ),
    .A(_0448_),
    .Y(_0272_));
 sg13g2_or2_1 _1984_ (.X(_0273_),
    .B(\pulse_width_counter_module.low_counter[0] ),
    .A(net51));
 sg13g2_a21oi_1 _1985_ (.A1(_0272_),
    .A2(_0273_),
    .Y(_0128_),
    .B1(net36));
 sg13g2_inv_1 _1986_ (.Y(_0274_),
    .A(\pulse_width_counter_module.low_counter[5] ));
 sg13g2_inv_1 _1987_ (.Y(_0275_),
    .A(\pulse_width_counter_module.low_counter[2] ));
 sg13g2_inv_1 _1988_ (.Y(_0276_),
    .A(\pulse_width_counter_module.low_counter[3] ));
 sg13g2_inv_1 _1989_ (.Y(_0277_),
    .A(\pulse_width_counter_module.low_counter[4] ));
 sg13g2_nand3b_1 _1990_ (.B(\pulse_width_counter_module.low_counter[0] ),
    .C(\pulse_width_counter_module.low_counter[1] ),
    .Y(_0278_),
    .A_N(_0447_));
 sg13g2_or4_1 _1991_ (.A(_0275_),
    .B(_0276_),
    .C(_0277_),
    .D(_0278_),
    .X(_0279_));
 sg13g2_buf_1 _1992_ (.A(_0279_),
    .X(_0280_));
 sg13g2_nor2_1 _1993_ (.A(_0274_),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_nand3_1 _1994_ (.B(\pulse_width_counter_module.low_counter[7] ),
    .C(_0281_),
    .A(\pulse_width_counter_module.low_counter[6] ),
    .Y(_0282_));
 sg13g2_and2_1 _1995_ (.A(\pulse_width_counter_module.low_counter[8] ),
    .B(\pulse_width_counter_module.low_counter[9] ),
    .X(_0283_));
 sg13g2_nor2b_1 _1996_ (.A(_0282_),
    .B_N(_0283_),
    .Y(_0284_));
 sg13g2_buf_1 _1997_ (.A(_0938_),
    .X(_0285_));
 sg13g2_nand3b_1 _1998_ (.B(\pulse_width_counter_module.low_counter[10] ),
    .C(net33),
    .Y(_0286_),
    .A_N(_0284_));
 sg13g2_nand2b_1 _1999_ (.Y(_0287_),
    .B(_0284_),
    .A_N(\pulse_width_counter_module.low_counter[10] ));
 sg13g2_a21oi_1 _2000_ (.A1(_0286_),
    .A2(_0287_),
    .Y(_0129_),
    .B1(net36));
 sg13g2_nand2_1 _2001_ (.Y(_0288_),
    .A(\pulse_width_counter_module.low_counter[10] ),
    .B(_0284_));
 sg13g2_nand3_1 _2002_ (.B(net17),
    .C(_0288_),
    .A(\pulse_width_counter_module.low_counter[11] ),
    .Y(_0289_));
 sg13g2_or2_1 _2003_ (.X(_0290_),
    .B(_0288_),
    .A(\pulse_width_counter_module.low_counter[11] ));
 sg13g2_a21oi_1 _2004_ (.A1(_0289_),
    .A2(_0290_),
    .Y(_0130_),
    .B1(net36));
 sg13g2_nand2_2 _2005_ (.Y(_0291_),
    .A(net63),
    .B(_0285_));
 sg13g2_inv_1 _2006_ (.Y(_0292_),
    .A(\pulse_width_counter_module.low_counter[12] ));
 sg13g2_inv_1 _2007_ (.Y(_0293_),
    .A(\pulse_width_counter_module.low_counter[6] ));
 sg13g2_nand4_1 _2008_ (.B(\pulse_width_counter_module.low_counter[10] ),
    .C(\pulse_width_counter_module.low_counter[11] ),
    .A(\pulse_width_counter_module.low_counter[7] ),
    .Y(_0294_),
    .D(_0283_));
 sg13g2_or4_1 _2009_ (.A(_0274_),
    .B(_0293_),
    .C(_0280_),
    .D(_0294_),
    .X(_0295_));
 sg13g2_xnor2_1 _2010_ (.Y(_0296_),
    .A(_0292_),
    .B(_0295_));
 sg13g2_nor2_1 _2011_ (.A(_0291_),
    .B(_0296_),
    .Y(_0131_));
 sg13g2_inv_1 _2012_ (.Y(_0297_),
    .A(\pulse_width_counter_module.low_counter[13] ));
 sg13g2_nor2_1 _2013_ (.A(_0292_),
    .B(_0295_),
    .Y(_0298_));
 sg13g2_nor3_1 _2014_ (.A(_0297_),
    .B(_0934_),
    .C(_0298_),
    .Y(_0299_));
 sg13g2_a21oi_1 _2015_ (.A1(_0297_),
    .A2(_0298_),
    .Y(_0300_),
    .B1(_0299_));
 sg13g2_nor2_1 _2016_ (.A(net45),
    .B(_0300_),
    .Y(_0132_));
 sg13g2_inv_1 _2017_ (.Y(_0301_),
    .A(\pulse_width_counter_module.low_counter[14] ));
 sg13g2_and2_1 _2018_ (.A(\pulse_width_counter_module.low_counter[13] ),
    .B(_0298_),
    .X(_0302_));
 sg13g2_buf_2 _2019_ (.A(_0302_),
    .X(_0303_));
 sg13g2_nor3_1 _2020_ (.A(_0301_),
    .B(_0934_),
    .C(_0303_),
    .Y(_0304_));
 sg13g2_a21oi_1 _2021_ (.A1(_0301_),
    .A2(_0303_),
    .Y(_0305_),
    .B1(_0304_));
 sg13g2_nor2_1 _2022_ (.A(net45),
    .B(_0305_),
    .Y(_0133_));
 sg13g2_nand2_1 _2023_ (.Y(_0306_),
    .A(\pulse_width_counter_module.low_counter[14] ),
    .B(_0303_));
 sg13g2_nand3_1 _2024_ (.B(net34),
    .C(_0306_),
    .A(_0953_),
    .Y(_0307_));
 sg13g2_o21ai_1 _2025_ (.B1(_0307_),
    .Y(_0308_),
    .A1(_0953_),
    .A2(_0306_));
 sg13g2_and2_1 _2026_ (.A(net58),
    .B(_0308_),
    .X(_0134_));
 sg13g2_nand3_1 _2027_ (.B(_0953_),
    .C(_0303_),
    .A(\pulse_width_counter_module.low_counter[14] ),
    .Y(_0309_));
 sg13g2_nand3_1 _2028_ (.B(net34),
    .C(_0309_),
    .A(\pulse_width_counter_module.low_counter[16] ),
    .Y(_0310_));
 sg13g2_o21ai_1 _2029_ (.B1(_0310_),
    .Y(_0311_),
    .A1(\pulse_width_counter_module.low_counter[16] ),
    .A2(_0309_));
 sg13g2_and2_1 _2030_ (.A(net58),
    .B(_0311_),
    .X(_0135_));
 sg13g2_nand4_1 _2031_ (.B(_0953_),
    .C(\pulse_width_counter_module.low_counter[16] ),
    .A(\pulse_width_counter_module.low_counter[14] ),
    .Y(_0312_),
    .D(_0303_));
 sg13g2_nand3_1 _2032_ (.B(net34),
    .C(_0312_),
    .A(\pulse_width_counter_module.low_counter[17] ),
    .Y(_0313_));
 sg13g2_o21ai_1 _2033_ (.B1(_0313_),
    .Y(_0314_),
    .A1(\pulse_width_counter_module.low_counter[17] ),
    .A2(_0312_));
 sg13g2_and2_1 _2034_ (.A(net58),
    .B(_0314_),
    .X(_0136_));
 sg13g2_and4_1 _2035_ (.A(\pulse_width_counter_module.low_counter[14] ),
    .B(_0953_),
    .C(\pulse_width_counter_module.low_counter[16] ),
    .D(\pulse_width_counter_module.low_counter[17] ),
    .X(_0315_));
 sg13g2_nand2_1 _2036_ (.Y(_0316_),
    .A(_0303_),
    .B(_0315_));
 sg13g2_nand3_1 _2037_ (.B(net17),
    .C(_0316_),
    .A(\pulse_width_counter_module.low_counter[18] ),
    .Y(_0317_));
 sg13g2_or2_1 _2038_ (.X(_0318_),
    .B(_0316_),
    .A(\pulse_width_counter_module.low_counter[18] ));
 sg13g2_buf_1 _2039_ (.A(net59),
    .X(_0319_));
 sg13g2_a21oi_1 _2040_ (.A1(_0317_),
    .A2(_0318_),
    .Y(_0137_),
    .B1(net35));
 sg13g2_and2_1 _2041_ (.A(\pulse_width_counter_module.low_counter[18] ),
    .B(_0315_),
    .X(_0320_));
 sg13g2_nand2_1 _2042_ (.Y(_0321_),
    .A(_0303_),
    .B(_0320_));
 sg13g2_nand3_1 _2043_ (.B(net17),
    .C(_0321_),
    .A(\pulse_width_counter_module.low_counter[19] ),
    .Y(_0322_));
 sg13g2_or2_1 _2044_ (.X(_0323_),
    .B(_0321_),
    .A(\pulse_width_counter_module.low_counter[19] ));
 sg13g2_a21oi_1 _2045_ (.A1(_0322_),
    .A2(_0323_),
    .Y(_0138_),
    .B1(net35));
 sg13g2_xnor2_1 _2046_ (.Y(_0324_),
    .A(\pulse_width_counter_module.low_counter[0] ),
    .B(\pulse_width_counter_module.low_counter[1] ));
 sg13g2_nand3_1 _2047_ (.B(net51),
    .C(\pulse_width_counter_module.low_counter[1] ),
    .A(_0448_),
    .Y(_0325_));
 sg13g2_o21ai_1 _2048_ (.B1(_0325_),
    .Y(_0326_),
    .A1(net51),
    .A2(_0324_));
 sg13g2_and2_1 _2049_ (.A(net58),
    .B(_0326_),
    .X(_0139_));
 sg13g2_nand3_1 _2050_ (.B(_0303_),
    .C(_0320_),
    .A(\pulse_width_counter_module.low_counter[19] ),
    .Y(_0327_));
 sg13g2_nand3_1 _2051_ (.B(net17),
    .C(_0327_),
    .A(\pulse_width_counter_module.low_counter[20] ),
    .Y(_0328_));
 sg13g2_inv_1 _2052_ (.Y(_0329_),
    .A(\pulse_width_counter_module.low_counter[20] ));
 sg13g2_nand2b_1 _2053_ (.Y(_0330_),
    .B(_0329_),
    .A_N(_0327_));
 sg13g2_a21oi_1 _2054_ (.A1(_0328_),
    .A2(_0330_),
    .Y(_0140_),
    .B1(net35));
 sg13g2_nand3_1 _2055_ (.B(\pulse_width_counter_module.low_counter[19] ),
    .C(_0320_),
    .A(\pulse_width_counter_module.low_counter[13] ),
    .Y(_0331_));
 sg13g2_nor4_2 _2056_ (.A(_0292_),
    .B(_0329_),
    .C(_0295_),
    .Y(_0332_),
    .D(_0331_));
 sg13g2_nand3b_1 _2057_ (.B(_0970_),
    .C(net33),
    .Y(_0333_),
    .A_N(_0332_));
 sg13g2_nand2b_1 _2058_ (.Y(_0334_),
    .B(_0332_),
    .A_N(_0970_));
 sg13g2_a21oi_1 _2059_ (.A1(_0333_),
    .A2(_0334_),
    .Y(_0141_),
    .B1(net35));
 sg13g2_nand2_1 _2060_ (.Y(_0335_),
    .A(_0970_),
    .B(_0332_));
 sg13g2_nand3_1 _2061_ (.B(net17),
    .C(_0335_),
    .A(\pulse_width_counter_module.low_counter[22] ),
    .Y(_0336_));
 sg13g2_or2_1 _2062_ (.X(_0337_),
    .B(_0335_),
    .A(\pulse_width_counter_module.low_counter[22] ));
 sg13g2_a21oi_1 _2063_ (.A1(_0336_),
    .A2(_0337_),
    .Y(_0142_),
    .B1(_0319_));
 sg13g2_nand2_1 _2064_ (.Y(_0338_),
    .A(\pulse_width_counter_module.low_counter[23] ),
    .B(net34));
 sg13g2_nand3_1 _2065_ (.B(\pulse_width_counter_module.low_counter[22] ),
    .C(_0332_),
    .A(_0970_),
    .Y(_0339_));
 sg13g2_mux2_1 _2066_ (.A0(\pulse_width_counter_module.low_counter[23] ),
    .A1(_0338_),
    .S(_0339_),
    .X(_0340_));
 sg13g2_nor2_1 _2067_ (.A(net45),
    .B(_0340_),
    .Y(_0143_));
 sg13g2_nand4_1 _2068_ (.B(\pulse_width_counter_module.low_counter[22] ),
    .C(\pulse_width_counter_module.low_counter[23] ),
    .A(_0970_),
    .Y(_0341_),
    .D(_0332_));
 sg13g2_nand3_1 _2069_ (.B(_1010_),
    .C(_0341_),
    .A(\pulse_width_counter_module.low_counter[24] ),
    .Y(_0342_));
 sg13g2_or2_1 _2070_ (.X(_0343_),
    .B(_0341_),
    .A(\pulse_width_counter_module.low_counter[24] ));
 sg13g2_a21oi_1 _2071_ (.A1(_0342_),
    .A2(_0343_),
    .Y(_0144_),
    .B1(net35));
 sg13g2_and2_1 _2072_ (.A(\pulse_width_counter_module.low_counter[22] ),
    .B(\pulse_width_counter_module.low_counter[23] ),
    .X(_0344_));
 sg13g2_and4_1 _2073_ (.A(_0970_),
    .B(\pulse_width_counter_module.low_counter[24] ),
    .C(_0332_),
    .D(_0344_),
    .X(_0345_));
 sg13g2_buf_1 _2074_ (.A(_0345_),
    .X(_0346_));
 sg13g2_nand3b_1 _2075_ (.B(\pulse_width_counter_module.low_counter[25] ),
    .C(net33),
    .Y(_0347_),
    .A_N(_0346_));
 sg13g2_nand2b_1 _2076_ (.Y(_0348_),
    .B(_0346_),
    .A_N(\pulse_width_counter_module.low_counter[25] ));
 sg13g2_a21oi_1 _2077_ (.A1(_0347_),
    .A2(_0348_),
    .Y(_0145_),
    .B1(net35));
 sg13g2_nand2_1 _2078_ (.Y(_0349_),
    .A(\pulse_width_counter_module.low_counter[25] ),
    .B(_0346_));
 sg13g2_nand3_1 _2079_ (.B(_1010_),
    .C(_0349_),
    .A(\pulse_width_counter_module.low_counter[26] ),
    .Y(_0350_));
 sg13g2_or2_1 _2080_ (.X(_0351_),
    .B(_0349_),
    .A(\pulse_width_counter_module.low_counter[26] ));
 sg13g2_a21oi_1 _2081_ (.A1(_0350_),
    .A2(_0351_),
    .Y(_0146_),
    .B1(net35));
 sg13g2_nand2_1 _2082_ (.Y(_0352_),
    .A(\pulse_width_counter_module.low_counter[27] ),
    .B(_0939_));
 sg13g2_and3_1 _2083_ (.X(_0353_),
    .A(\pulse_width_counter_module.low_counter[25] ),
    .B(\pulse_width_counter_module.low_counter[26] ),
    .C(_0346_));
 sg13g2_mux2_1 _2084_ (.A0(_0352_),
    .A1(\pulse_width_counter_module.low_counter[27] ),
    .S(_0353_),
    .X(_0354_));
 sg13g2_nor2_1 _2085_ (.A(net45),
    .B(_0354_),
    .Y(_0147_));
 sg13g2_nand2_1 _2086_ (.Y(_0355_),
    .A(\pulse_width_counter_module.low_counter[27] ),
    .B(_0353_));
 sg13g2_nand2b_1 _2087_ (.Y(_0356_),
    .B(net56),
    .A_N(\pulse_width_counter_module.low_counter[28] ));
 sg13g2_nand4_1 _2088_ (.B(net63),
    .C(net33),
    .A(\pulse_width_counter_module.low_counter[28] ),
    .Y(_0357_),
    .D(_0355_));
 sg13g2_o21ai_1 _2089_ (.B1(_0357_),
    .Y(_0148_),
    .A1(_0355_),
    .A2(_0356_));
 sg13g2_nand3_1 _2090_ (.B(\pulse_width_counter_module.low_counter[28] ),
    .C(_0353_),
    .A(\pulse_width_counter_module.low_counter[27] ),
    .Y(_0358_));
 sg13g2_nand2b_1 _2091_ (.Y(_0359_),
    .B(net63),
    .A_N(\pulse_width_counter_module.low_counter[29] ));
 sg13g2_nand4_1 _2092_ (.B(net63),
    .C(net33),
    .A(\pulse_width_counter_module.low_counter[29] ),
    .Y(_0360_),
    .D(_0358_));
 sg13g2_o21ai_1 _2093_ (.B1(_0360_),
    .Y(_0149_),
    .A1(_0358_),
    .A2(_0359_));
 sg13g2_xnor2_1 _2094_ (.Y(_0361_),
    .A(_0275_),
    .B(_0278_));
 sg13g2_nor2_1 _2095_ (.A(_0291_),
    .B(_0361_),
    .Y(_0150_));
 sg13g2_nand4_1 _2096_ (.B(\pulse_width_counter_module.low_counter[27] ),
    .C(\pulse_width_counter_module.low_counter[28] ),
    .A(\pulse_width_counter_module.low_counter[26] ),
    .Y(_0362_),
    .D(\pulse_width_counter_module.low_counter[29] ));
 sg13g2_nor2_1 _2097_ (.A(_0349_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_nand3b_1 _2098_ (.B(\pulse_width_counter_module.low_counter[30] ),
    .C(net33),
    .Y(_0364_),
    .A_N(_0363_));
 sg13g2_nand2b_1 _2099_ (.Y(_0365_),
    .B(_0363_),
    .A_N(\pulse_width_counter_module.low_counter[30] ));
 sg13g2_a21oi_1 _2100_ (.A1(_0364_),
    .A2(_0365_),
    .Y(_0151_),
    .B1(net35));
 sg13g2_nand3_1 _2101_ (.B(net63),
    .C(net33),
    .A(\pulse_width_counter_module.low_counter[31] ),
    .Y(_0366_));
 sg13g2_a21oi_1 _2102_ (.A1(\pulse_width_counter_module.low_counter[30] ),
    .A2(_0363_),
    .Y(_0367_),
    .B1(_0366_));
 sg13g2_nor2_1 _2103_ (.A(\pulse_width_counter_module.low_counter[31] ),
    .B(_0445_),
    .Y(_0368_));
 sg13g2_nand3_1 _2104_ (.B(_0363_),
    .C(_0368_),
    .A(\pulse_width_counter_module.low_counter[30] ),
    .Y(_0369_));
 sg13g2_nand2b_1 _2105_ (.Y(_0152_),
    .B(_0369_),
    .A_N(_0367_));
 sg13g2_nor2_1 _2106_ (.A(_0275_),
    .B(_0278_),
    .Y(_0370_));
 sg13g2_xnor2_1 _2107_ (.Y(_0371_),
    .A(\pulse_width_counter_module.low_counter[3] ),
    .B(_0370_));
 sg13g2_nor2_1 _2108_ (.A(_0291_),
    .B(_0371_),
    .Y(_0153_));
 sg13g2_nor3_1 _2109_ (.A(_0275_),
    .B(_0276_),
    .C(_0278_),
    .Y(_0372_));
 sg13g2_nand3b_1 _2110_ (.B(\pulse_width_counter_module.low_counter[4] ),
    .C(_0285_),
    .Y(_0373_),
    .A_N(_0372_));
 sg13g2_nand2_1 _2111_ (.Y(_0374_),
    .A(_0277_),
    .B(_0372_));
 sg13g2_a21oi_1 _2112_ (.A1(_0373_),
    .A2(_0374_),
    .Y(_0154_),
    .B1(_0319_));
 sg13g2_nand3_1 _2113_ (.B(_0939_),
    .C(_0280_),
    .A(\pulse_width_counter_module.low_counter[5] ),
    .Y(_0375_));
 sg13g2_o21ai_1 _2114_ (.B1(_0375_),
    .Y(_0376_),
    .A1(\pulse_width_counter_module.low_counter[5] ),
    .A2(_0280_));
 sg13g2_and2_1 _2115_ (.A(net56),
    .B(_0376_),
    .X(_0155_));
 sg13g2_xnor2_1 _2116_ (.Y(_0377_),
    .A(\pulse_width_counter_module.low_counter[6] ),
    .B(_0281_));
 sg13g2_nor2_1 _2117_ (.A(_0291_),
    .B(_0377_),
    .Y(_0156_));
 sg13g2_nand2_1 _2118_ (.Y(_0378_),
    .A(\pulse_width_counter_module.low_counter[6] ),
    .B(_0281_));
 sg13g2_nand3_1 _2119_ (.B(net17),
    .C(_0378_),
    .A(\pulse_width_counter_module.low_counter[7] ),
    .Y(_0379_));
 sg13g2_or2_1 _2120_ (.X(_0380_),
    .B(_0378_),
    .A(\pulse_width_counter_module.low_counter[7] ));
 sg13g2_a21oi_1 _2121_ (.A1(_0379_),
    .A2(_0380_),
    .Y(_0157_),
    .B1(net61));
 sg13g2_nand3_1 _2122_ (.B(net33),
    .C(_0282_),
    .A(\pulse_width_counter_module.low_counter[8] ),
    .Y(_0381_));
 sg13g2_inv_1 _2123_ (.Y(_0382_),
    .A(\pulse_width_counter_module.low_counter[8] ));
 sg13g2_nand2b_1 _2124_ (.Y(_0383_),
    .B(_0382_),
    .A_N(_0282_));
 sg13g2_a21oi_1 _2125_ (.A1(_0381_),
    .A2(_0383_),
    .Y(_0158_),
    .B1(net61));
 sg13g2_nor2_1 _2126_ (.A(_0382_),
    .B(_0282_),
    .Y(_0384_));
 sg13g2_xnor2_1 _2127_ (.Y(_0385_),
    .A(\pulse_width_counter_module.low_counter[9] ),
    .B(_0384_));
 sg13g2_nor2_1 _2128_ (.A(_0291_),
    .B(_0385_),
    .Y(_0159_));
 sg13g2_and2_1 _2129_ (.A(net51),
    .B(net56),
    .X(_0160_));
 sg13g2_buf_1 _2130_ (.A(ui_in[3]),
    .X(_0386_));
 sg13g2_buf_2 _2131_ (.A(ui_in[4]),
    .X(_0387_));
 sg13g2_buf_1 _2132_ (.A(_0387_),
    .X(_0388_));
 sg13g2_buf_4 _2133_ (.X(_0389_),
    .A(ui_in[1]));
 sg13g2_buf_2 _2134_ (.A(_0389_),
    .X(_0390_));
 sg13g2_buf_2 _2135_ (.A(ui_in[2]),
    .X(_0391_));
 sg13g2_buf_1 _2136_ (.A(_0391_),
    .X(_0392_));
 sg13g2_mux4_1 _2137_ (.S0(net49),
    .A0(\mux.data_in[64] ),
    .A1(_0464_),
    .A2(net57),
    .A3(net52),
    .S1(net48),
    .X(_0393_));
 sg13g2_buf_2 _2138_ (.A(_0389_),
    .X(_0394_));
 sg13g2_buf_1 _2139_ (.A(_0391_),
    .X(_0395_));
 sg13g2_mux4_1 _2140_ (.S0(net47),
    .A0(\mux.data_in[0] ),
    .A1(\mux.data_in[8] ),
    .A2(\mux.data_in[16] ),
    .A3(\mux.data_in[24] ),
    .S1(net46),
    .X(_0396_));
 sg13g2_nor2b_1 _2141_ (.A(net50),
    .B_N(_0396_),
    .Y(_0397_));
 sg13g2_a21oi_1 _2142_ (.A1(net50),
    .A2(_0393_),
    .Y(_0398_),
    .B1(_0397_));
 sg13g2_mux4_1 _2143_ (.S0(net49),
    .A0(\mux.data_in[32] ),
    .A1(_0463_),
    .A2(_0582_),
    .A3(_0703_),
    .S1(net48),
    .X(_0399_));
 sg13g2_nor2b_1 _2144_ (.A(_0387_),
    .B_N(net62),
    .Y(_0400_));
 sg13g2_buf_2 _2145_ (.A(_0400_),
    .X(_0401_));
 sg13g2_nand2_1 _2146_ (.Y(_0402_),
    .A(_0399_),
    .B(_0401_));
 sg13g2_o21ai_1 _2147_ (.B1(_0402_),
    .Y(net2),
    .A1(net62),
    .A2(_0398_));
 sg13g2_mux4_1 _2148_ (.S0(net49),
    .A0(\mux.data_in[65] ),
    .A1(_0461_),
    .A2(net55),
    .A3(_0718_),
    .S1(net48),
    .X(_0403_));
 sg13g2_mux4_1 _2149_ (.S0(net47),
    .A0(\mux.data_in[1] ),
    .A1(\mux.data_in[9] ),
    .A2(\mux.data_in[17] ),
    .A3(\mux.data_in[25] ),
    .S1(net46),
    .X(_0404_));
 sg13g2_nor2b_1 _2150_ (.A(net50),
    .B_N(_0404_),
    .Y(_0405_));
 sg13g2_a21oi_1 _2151_ (.A1(net50),
    .A2(_0403_),
    .Y(_0406_),
    .B1(_0405_));
 sg13g2_mux4_1 _2152_ (.S0(net49),
    .A0(\mux.data_in[33] ),
    .A1(_0460_),
    .A2(_0603_),
    .A3(_0717_),
    .S1(net48),
    .X(_0407_));
 sg13g2_nand2_1 _2153_ (.Y(_0408_),
    .A(_0401_),
    .B(_0407_));
 sg13g2_o21ai_1 _2154_ (.B1(_0408_),
    .Y(net3),
    .A1(net62),
    .A2(_0406_));
 sg13g2_mux4_1 _2155_ (.S0(net47),
    .A0(_0480_),
    .A1(_0507_),
    .A2(_0625_),
    .A3(_0735_),
    .S1(net46),
    .X(_0409_));
 sg13g2_mux4_1 _2156_ (.S0(net47),
    .A0(\mux.data_in[2] ),
    .A1(\mux.data_in[10] ),
    .A2(\mux.data_in[18] ),
    .A3(\mux.data_in[26] ),
    .S1(net46),
    .X(_0410_));
 sg13g2_nor2b_1 _2157_ (.A(_0387_),
    .B_N(_0410_),
    .Y(_0411_));
 sg13g2_a21oi_1 _2158_ (.A1(net50),
    .A2(_0409_),
    .Y(_0412_),
    .B1(_0411_));
 sg13g2_mux4_1 _2159_ (.S0(net49),
    .A0(\mux.data_in[34] ),
    .A1(_0506_),
    .A2(\mux.data_in[50] ),
    .A3(_0734_),
    .S1(net48),
    .X(_0413_));
 sg13g2_nand2_1 _2160_ (.Y(_0414_),
    .A(_0401_),
    .B(_0413_));
 sg13g2_o21ai_1 _2161_ (.B1(_0414_),
    .Y(net4),
    .A1(net62),
    .A2(_0412_));
 sg13g2_mux4_1 _2162_ (.S0(_0394_),
    .A0(\mux.data_in[67] ),
    .A1(_0520_),
    .A2(_0651_),
    .A3(\mux.data_in[91] ),
    .S1(_0395_),
    .X(_0415_));
 sg13g2_mux4_1 _2163_ (.S0(_0394_),
    .A0(\mux.data_in[3] ),
    .A1(\mux.data_in[11] ),
    .A2(\mux.data_in[19] ),
    .A3(\mux.data_in[27] ),
    .S1(_0395_),
    .X(_0416_));
 sg13g2_nor2b_1 _2164_ (.A(_0387_),
    .B_N(_0416_),
    .Y(_0417_));
 sg13g2_a21oi_1 _2165_ (.A1(net50),
    .A2(_0415_),
    .Y(_0418_),
    .B1(_0417_));
 sg13g2_mux4_1 _2166_ (.S0(net49),
    .A0(\mux.data_in[35] ),
    .A1(_0519_),
    .A2(_0650_),
    .A3(\mux.data_in[59] ),
    .S1(net48),
    .X(_0419_));
 sg13g2_nand2_1 _2167_ (.Y(_0420_),
    .A(_0401_),
    .B(_0419_));
 sg13g2_o21ai_1 _2168_ (.B1(_0420_),
    .Y(net5),
    .A1(net62),
    .A2(_0418_));
 sg13g2_mux4_1 _2169_ (.S0(net47),
    .A0(_0487_),
    .A1(_0534_),
    .A2(_0663_),
    .A3(\mux.data_in[92] ),
    .S1(net46),
    .X(_0421_));
 sg13g2_mux4_1 _2170_ (.S0(_0389_),
    .A0(\mux.data_in[4] ),
    .A1(\mux.data_in[12] ),
    .A2(\mux.data_in[20] ),
    .A3(\mux.data_in[28] ),
    .S1(_0391_),
    .X(_0422_));
 sg13g2_nor2b_1 _2171_ (.A(_0387_),
    .B_N(_0422_),
    .Y(_0423_));
 sg13g2_a21oi_1 _2172_ (.A1(net50),
    .A2(_0421_),
    .Y(_0424_),
    .B1(_0423_));
 sg13g2_mux4_1 _2173_ (.S0(net49),
    .A0(_0486_),
    .A1(_0533_),
    .A2(_0662_),
    .A3(\mux.data_in[60] ),
    .S1(net48),
    .X(_0425_));
 sg13g2_nand2_1 _2174_ (.Y(_0426_),
    .A(_0401_),
    .B(_0425_));
 sg13g2_o21ai_1 _2175_ (.B1(_0426_),
    .Y(net6),
    .A1(net62),
    .A2(_0424_));
 sg13g2_mux4_1 _2176_ (.S0(net47),
    .A0(_0492_),
    .A1(_0555_),
    .A2(_0673_),
    .A3(\mux.data_in[93] ),
    .S1(net46),
    .X(_0427_));
 sg13g2_mux4_1 _2177_ (.S0(_0389_),
    .A0(\mux.data_in[5] ),
    .A1(\mux.data_in[13] ),
    .A2(\mux.data_in[21] ),
    .A3(\mux.data_in[29] ),
    .S1(_0391_),
    .X(_0428_));
 sg13g2_nor2b_1 _2178_ (.A(_0387_),
    .B_N(_0428_),
    .Y(_0429_));
 sg13g2_a21oi_1 _2179_ (.A1(_0388_),
    .A2(_0427_),
    .Y(_0430_),
    .B1(_0429_));
 sg13g2_mux4_1 _2180_ (.S0(_0390_),
    .A0(_0491_),
    .A1(_0554_),
    .A2(_0672_),
    .A3(\mux.data_in[61] ),
    .S1(_0392_),
    .X(_0431_));
 sg13g2_nand2_1 _2181_ (.Y(_0432_),
    .A(_0401_),
    .B(_0431_));
 sg13g2_o21ai_1 _2182_ (.B1(_0432_),
    .Y(net7),
    .A1(net62),
    .A2(_0430_));
 sg13g2_mux4_1 _2183_ (.S0(net47),
    .A0(_0489_),
    .A1(_0564_),
    .A2(\mux.data_in[86] ),
    .A3(\mux.data_in[94] ),
    .S1(net46),
    .X(_0433_));
 sg13g2_mux4_1 _2184_ (.S0(_0389_),
    .A0(\mux.data_in[6] ),
    .A1(\mux.data_in[14] ),
    .A2(\mux.data_in[22] ),
    .A3(\mux.data_in[30] ),
    .S1(_0391_),
    .X(_0434_));
 sg13g2_nor2b_1 _2185_ (.A(_0387_),
    .B_N(_0434_),
    .Y(_0435_));
 sg13g2_a21oi_1 _2186_ (.A1(_0388_),
    .A2(_0433_),
    .Y(_0436_),
    .B1(_0435_));
 sg13g2_mux4_1 _2187_ (.S0(_0390_),
    .A0(_0493_),
    .A1(_0563_),
    .A2(_0677_),
    .A3(\mux.data_in[62] ),
    .S1(_0392_),
    .X(_0437_));
 sg13g2_nand2_1 _2188_ (.Y(_0438_),
    .A(_0401_),
    .B(_0437_));
 sg13g2_o21ai_1 _2189_ (.B1(_0438_),
    .Y(net8),
    .A1(_0386_),
    .A2(_0436_));
 sg13g2_mux4_1 _2190_ (.S0(net47),
    .A0(_0468_),
    .A1(_0571_),
    .A2(_0699_),
    .A3(\mux.data_in[95] ),
    .S1(net46),
    .X(_0439_));
 sg13g2_mux4_1 _2191_ (.S0(_0389_),
    .A0(\mux.data_in[7] ),
    .A1(\mux.data_in[15] ),
    .A2(\mux.data_in[23] ),
    .A3(\mux.data_in[31] ),
    .S1(_0391_),
    .X(_0440_));
 sg13g2_nor2b_1 _2192_ (.A(_0387_),
    .B_N(_0440_),
    .Y(_0441_));
 sg13g2_a21oi_1 _2193_ (.A1(net50),
    .A2(_0439_),
    .Y(_0442_),
    .B1(_0441_));
 sg13g2_mux4_1 _2194_ (.S0(net49),
    .A0(_0467_),
    .A1(_0570_),
    .A2(net54),
    .A3(\mux.data_in[63] ),
    .S1(net48),
    .X(_0443_));
 sg13g2_nand2_1 _2195_ (.Y(_0444_),
    .A(_0401_),
    .B(_0443_));
 sg13g2_o21ai_1 _2196_ (.B1(_0444_),
    .Y(net9),
    .A1(net62),
    .A2(_0442_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[0]$_SDFFE_PN0P__80  (.L_HI(net80));
 sg13g2_buf_1 _2199_ (.A(net64),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2200_ (.A(net65),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2201_ (.A(net66),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2202_ (.A(net67),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2203_ (.A(net68),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2204_ (.A(net69),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2205_ (.A(net70),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2206_ (.A(net71),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2207_ (.A(net72),
    .X(uio_out[0]));
 sg13g2_buf_1 _2208_ (.A(net73),
    .X(uio_out[1]));
 sg13g2_buf_1 _2209_ (.A(net74),
    .X(uio_out[2]));
 sg13g2_buf_1 _2210_ (.A(net75),
    .X(uio_out[3]));
 sg13g2_buf_1 _2211_ (.A(net76),
    .X(uio_out[4]));
 sg13g2_buf_1 _2212_ (.A(net77),
    .X(uio_out[5]));
 sg13g2_buf_1 _2213_ (.A(net78),
    .X(uio_out[6]));
 sg13g2_buf_1 _2214_ (.A(net79),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[0]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net80),
    .D(_0000_),
    .Q_N(_1173_),
    .Q(\mux.data_in[0] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[10]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net81),
    .D(_0001_),
    .Q_N(_1172_),
    .Q(\mux.data_in[10] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[11]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net82),
    .D(_0002_),
    .Q_N(_1171_),
    .Q(\mux.data_in[11] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[12]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net83),
    .D(_0003_),
    .Q_N(_1170_),
    .Q(\mux.data_in[12] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[13]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net84),
    .D(_0004_),
    .Q_N(_1169_),
    .Q(\mux.data_in[13] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[14]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net85),
    .D(_0005_),
    .Q_N(_1168_),
    .Q(\mux.data_in[14] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[15]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net86),
    .D(_0006_),
    .Q_N(_1167_),
    .Q(\mux.data_in[15] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[16]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net87),
    .D(_0007_),
    .Q_N(_1166_),
    .Q(\mux.data_in[16] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[17]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net88),
    .D(_0008_),
    .Q_N(_1165_),
    .Q(\mux.data_in[17] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[18]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net89),
    .D(_0009_),
    .Q_N(_1164_),
    .Q(\mux.data_in[18] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[19]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net90),
    .D(_0010_),
    .Q_N(_1163_),
    .Q(\mux.data_in[19] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[1]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net91),
    .D(_0011_),
    .Q_N(_1162_),
    .Q(\mux.data_in[1] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[20]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net92),
    .D(_0012_),
    .Q_N(_1161_),
    .Q(\mux.data_in[20] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[21]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net93),
    .D(_0013_),
    .Q_N(_1160_),
    .Q(\mux.data_in[21] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[22]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net94),
    .D(_0014_),
    .Q_N(_1159_),
    .Q(\mux.data_in[22] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[23]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net95),
    .D(_0015_),
    .Q_N(_1158_),
    .Q(\mux.data_in[23] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[24]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net96),
    .D(_0016_),
    .Q_N(_1157_),
    .Q(\mux.data_in[24] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[25]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net97),
    .D(_0017_),
    .Q_N(_1156_),
    .Q(\mux.data_in[25] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[26]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net98),
    .D(_0018_),
    .Q_N(_1155_),
    .Q(\mux.data_in[26] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[27]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net99),
    .D(_0019_),
    .Q_N(_1154_),
    .Q(\mux.data_in[27] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[28]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net100),
    .D(_0020_),
    .Q_N(_1153_),
    .Q(\mux.data_in[28] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[29]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net101),
    .D(_0021_),
    .Q_N(_1152_),
    .Q(\mux.data_in[29] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[2]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net102),
    .D(_0022_),
    .Q_N(_1151_),
    .Q(\mux.data_in[2] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[30]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net103),
    .D(_0023_),
    .Q_N(_1150_),
    .Q(\mux.data_in[30] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[31]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net104),
    .D(_0024_),
    .Q_N(_1149_),
    .Q(\mux.data_in[31] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[3]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net105),
    .D(_0025_),
    .Q_N(_1148_),
    .Q(\mux.data_in[3] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[4]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net106),
    .D(_0026_),
    .Q_N(_1147_),
    .Q(\mux.data_in[4] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[5]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net107),
    .D(_0027_),
    .Q_N(_1146_),
    .Q(\mux.data_in[5] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[6]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net108),
    .D(_0028_),
    .Q_N(_1145_),
    .Q(\mux.data_in[6] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[7]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net109),
    .D(_0029_),
    .Q_N(_1144_),
    .Q(\mux.data_in[7] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[8]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net110),
    .D(_0030_),
    .Q_N(_1143_),
    .Q(\mux.data_in[8] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.PERIOD[9]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net111),
    .D(_0031_),
    .Q_N(_1142_),
    .Q(\mux.data_in[9] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[0]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net112),
    .D(_0032_),
    .Q_N(_1141_),
    .Q(\mux.data_in[64] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[10]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net113),
    .D(_0033_),
    .Q_N(_1140_),
    .Q(\mux.data_in[74] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[11]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net114),
    .D(_0034_),
    .Q_N(_1139_),
    .Q(\mux.data_in[75] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[12]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net115),
    .D(_0035_),
    .Q_N(_1138_),
    .Q(\mux.data_in[76] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[13]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net116),
    .D(_0036_),
    .Q_N(_1137_),
    .Q(\mux.data_in[77] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[14]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net117),
    .D(_0037_),
    .Q_N(_1136_),
    .Q(\mux.data_in[78] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[15]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net118),
    .D(_0038_),
    .Q_N(_1135_),
    .Q(\mux.data_in[79] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[16]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net119),
    .D(_0039_),
    .Q_N(_1134_),
    .Q(\mux.data_in[80] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[17]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net120),
    .D(_0040_),
    .Q_N(_1133_),
    .Q(\mux.data_in[81] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[18]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net121),
    .D(_0041_),
    .Q_N(_1132_),
    .Q(\mux.data_in[82] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[19]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net122),
    .D(_0042_),
    .Q_N(_1131_),
    .Q(\mux.data_in[83] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[1]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net123),
    .D(_0043_),
    .Q_N(_1130_),
    .Q(\mux.data_in[65] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[20]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net124),
    .D(_0044_),
    .Q_N(_1129_),
    .Q(\mux.data_in[84] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[21]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net125),
    .D(_0045_),
    .Q_N(_1128_),
    .Q(\mux.data_in[85] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[22]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net126),
    .D(_0046_),
    .Q_N(_1127_),
    .Q(\mux.data_in[86] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[23]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net127),
    .D(_0047_),
    .Q_N(_1126_),
    .Q(\mux.data_in[87] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[24]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net128),
    .D(_0048_),
    .Q_N(_1125_),
    .Q(\mux.data_in[88] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[25]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net129),
    .D(_0049_),
    .Q_N(_1124_),
    .Q(\mux.data_in[89] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[26]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net130),
    .D(_0050_),
    .Q_N(_1123_),
    .Q(\mux.data_in[90] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[27]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net131),
    .D(_0051_),
    .Q_N(_1122_),
    .Q(\mux.data_in[91] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[28]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net132),
    .D(_0052_),
    .Q_N(_1121_),
    .Q(\mux.data_in[92] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[29]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net133),
    .D(_0053_),
    .Q_N(_1120_),
    .Q(\mux.data_in[93] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[2]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net134),
    .D(_0054_),
    .Q_N(_1119_),
    .Q(\mux.data_in[66] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[30]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net135),
    .D(_0055_),
    .Q_N(_1118_),
    .Q(\mux.data_in[94] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[31]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net136),
    .D(_0056_),
    .Q_N(_1117_),
    .Q(\mux.data_in[95] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[3]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net137),
    .D(_0057_),
    .Q_N(_1116_),
    .Q(\mux.data_in[67] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[4]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net138),
    .D(_0058_),
    .Q_N(_1115_),
    .Q(\mux.data_in[68] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[5]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net139),
    .D(_0059_),
    .Q_N(_1114_),
    .Q(\mux.data_in[69] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[6]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net140),
    .D(_0060_),
    .Q_N(_1113_),
    .Q(\mux.data_in[70] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[7]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net141),
    .D(_0061_),
    .Q_N(_1112_),
    .Q(\mux.data_in[71] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[8]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net142),
    .D(_0062_),
    .Q_N(_1111_),
    .Q(\mux.data_in[72] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_HIGH[9]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net143),
    .D(_0063_),
    .Q_N(_1110_),
    .Q(\mux.data_in[73] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[0]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net144),
    .D(_0064_),
    .Q_N(_1109_),
    .Q(\mux.data_in[32] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[10]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net145),
    .D(_0065_),
    .Q_N(_1108_),
    .Q(\mux.data_in[42] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[11]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net146),
    .D(_0066_),
    .Q_N(_1107_),
    .Q(\mux.data_in[43] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[12]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net147),
    .D(_0067_),
    .Q_N(_1106_),
    .Q(\mux.data_in[44] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[13]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net148),
    .D(_0068_),
    .Q_N(_1105_),
    .Q(\mux.data_in[45] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[14]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net149),
    .D(_0069_),
    .Q_N(_1104_),
    .Q(\mux.data_in[46] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[15]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net150),
    .D(_0070_),
    .Q_N(_1103_),
    .Q(\mux.data_in[47] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[16]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net151),
    .D(_0071_),
    .Q_N(_1102_),
    .Q(\mux.data_in[48] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[17]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net152),
    .D(_0072_),
    .Q_N(_1101_),
    .Q(\mux.data_in[49] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[18]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net153),
    .D(_0073_),
    .Q_N(_1100_),
    .Q(\mux.data_in[50] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[19]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net154),
    .D(_0074_),
    .Q_N(_1099_),
    .Q(\mux.data_in[51] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[1]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net155),
    .D(_0075_),
    .Q_N(_1098_),
    .Q(\mux.data_in[33] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[20]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net156),
    .D(_0076_),
    .Q_N(_1097_),
    .Q(\mux.data_in[52] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[21]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net157),
    .D(_0077_),
    .Q_N(_1096_),
    .Q(\mux.data_in[53] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[22]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net158),
    .D(_0078_),
    .Q_N(_1095_),
    .Q(\mux.data_in[54] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[23]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net159),
    .D(_0079_),
    .Q_N(_1094_),
    .Q(\mux.data_in[55] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[24]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net160),
    .D(_0080_),
    .Q_N(_1093_),
    .Q(\mux.data_in[56] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[25]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net161),
    .D(_0081_),
    .Q_N(_1092_),
    .Q(\mux.data_in[57] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[26]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net162),
    .D(_0082_),
    .Q_N(_1091_),
    .Q(\mux.data_in[58] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[27]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net163),
    .D(_0083_),
    .Q_N(_1090_),
    .Q(\mux.data_in[59] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[28]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net164),
    .D(_0084_),
    .Q_N(_1089_),
    .Q(\mux.data_in[60] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[29]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net165),
    .D(_0085_),
    .Q_N(_1088_),
    .Q(\mux.data_in[61] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[2]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net166),
    .D(_0086_),
    .Q_N(_1087_),
    .Q(\mux.data_in[34] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[30]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net167),
    .D(_0087_),
    .Q_N(_1086_),
    .Q(\mux.data_in[62] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[31]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net168),
    .D(_0088_),
    .Q_N(_1085_),
    .Q(\mux.data_in[63] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[3]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net169),
    .D(_0089_),
    .Q_N(_1084_),
    .Q(\mux.data_in[35] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[4]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net170),
    .D(_0090_),
    .Q_N(_1083_),
    .Q(\mux.data_in[36] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[5]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net171),
    .D(_0091_),
    .Q_N(_1082_),
    .Q(\mux.data_in[37] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[6]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net172),
    .D(_0092_),
    .Q_N(_1081_),
    .Q(\mux.data_in[38] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[7]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net173),
    .D(_0093_),
    .Q_N(_1080_),
    .Q(\mux.data_in[39] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[8]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net174),
    .D(_0094_),
    .Q_N(_1079_),
    .Q(\mux.data_in[40] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.TIME_LOW[9]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net175),
    .D(_0095_),
    .Q_N(_1078_),
    .Q(\mux.data_in[41] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net176),
    .D(_0096_),
    .Q_N(_1077_),
    .Q(\pulse_width_counter_module.high_counter[0] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[10]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net177),
    .D(_0097_),
    .Q_N(_1076_),
    .Q(\pulse_width_counter_module.high_counter[10] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[11]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net178),
    .D(_0098_),
    .Q_N(_1075_),
    .Q(\pulse_width_counter_module.high_counter[11] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[12]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net179),
    .D(_0099_),
    .Q_N(_1074_),
    .Q(\pulse_width_counter_module.high_counter[12] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[13]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net180),
    .D(_0100_),
    .Q_N(_1073_),
    .Q(\pulse_width_counter_module.high_counter[13] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[14]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net181),
    .D(_0101_),
    .Q_N(_1072_),
    .Q(\pulse_width_counter_module.high_counter[14] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[15]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net182),
    .D(_0102_),
    .Q_N(_1071_),
    .Q(\pulse_width_counter_module.high_counter[15] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[16]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net183),
    .D(_0103_),
    .Q_N(_1070_),
    .Q(\pulse_width_counter_module.high_counter[16] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[17]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net184),
    .D(_0104_),
    .Q_N(_1069_),
    .Q(\pulse_width_counter_module.high_counter[17] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[18]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net185),
    .D(_0105_),
    .Q_N(_1068_),
    .Q(\pulse_width_counter_module.high_counter[18] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[19]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net186),
    .D(_0106_),
    .Q_N(_1067_),
    .Q(\pulse_width_counter_module.high_counter[19] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net187),
    .D(_0107_),
    .Q_N(_1066_),
    .Q(\pulse_width_counter_module.high_counter[1] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[20]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net188),
    .D(_0108_),
    .Q_N(_1065_),
    .Q(\pulse_width_counter_module.high_counter[20] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[21]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net189),
    .D(_0109_),
    .Q_N(_1064_),
    .Q(\pulse_width_counter_module.high_counter[21] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[22]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net190),
    .D(_0110_),
    .Q_N(_1063_),
    .Q(\pulse_width_counter_module.high_counter[22] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[23]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net191),
    .D(_0111_),
    .Q_N(_1062_),
    .Q(\pulse_width_counter_module.high_counter[23] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[24]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net192),
    .D(_0112_),
    .Q_N(_1061_),
    .Q(\pulse_width_counter_module.high_counter[24] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[25]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net193),
    .D(_0113_),
    .Q_N(_1060_),
    .Q(\pulse_width_counter_module.high_counter[25] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[26]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net194),
    .D(_0114_),
    .Q_N(_1059_),
    .Q(\pulse_width_counter_module.high_counter[26] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[27]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net195),
    .D(_0115_),
    .Q_N(_1058_),
    .Q(\pulse_width_counter_module.high_counter[27] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[28]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net196),
    .D(_0116_),
    .Q_N(_1057_),
    .Q(\pulse_width_counter_module.high_counter[28] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[29]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net197),
    .D(_0117_),
    .Q_N(_1056_),
    .Q(\pulse_width_counter_module.high_counter[29] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net198),
    .D(_0118_),
    .Q_N(_1055_),
    .Q(\pulse_width_counter_module.high_counter[2] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[30]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net199),
    .D(_0119_),
    .Q_N(_1054_),
    .Q(\pulse_width_counter_module.high_counter[30] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[31]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net200),
    .D(_0120_),
    .Q_N(_1053_),
    .Q(\pulse_width_counter_module.high_counter[31] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net201),
    .D(_0121_),
    .Q_N(_1052_),
    .Q(\pulse_width_counter_module.high_counter[3] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net202),
    .D(_0122_),
    .Q_N(_1051_),
    .Q(\pulse_width_counter_module.high_counter[4] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net203),
    .D(_0123_),
    .Q_N(_1050_),
    .Q(\pulse_width_counter_module.high_counter[5] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net204),
    .D(_0124_),
    .Q_N(_1049_),
    .Q(\pulse_width_counter_module.high_counter[6] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[7]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net205),
    .D(_0125_),
    .Q_N(_1048_),
    .Q(\pulse_width_counter_module.high_counter[7] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[8]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net206),
    .D(_0126_),
    .Q_N(_1047_),
    .Q(\pulse_width_counter_module.high_counter[8] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.high_counter[9]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net207),
    .D(_0127_),
    .Q_N(_1046_),
    .Q(\pulse_width_counter_module.high_counter[9] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net208),
    .D(_0128_),
    .Q_N(_1045_),
    .Q(\pulse_width_counter_module.low_counter[0] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[10]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net209),
    .D(_0129_),
    .Q_N(_1044_),
    .Q(\pulse_width_counter_module.low_counter[10] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[11]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net210),
    .D(_0130_),
    .Q_N(_1043_),
    .Q(\pulse_width_counter_module.low_counter[11] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[12]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net211),
    .D(_0131_),
    .Q_N(_1042_),
    .Q(\pulse_width_counter_module.low_counter[12] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[13]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net212),
    .D(_0132_),
    .Q_N(_1041_),
    .Q(\pulse_width_counter_module.low_counter[13] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[14]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net213),
    .D(_0133_),
    .Q_N(_1040_),
    .Q(\pulse_width_counter_module.low_counter[14] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[15]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net214),
    .D(_0134_),
    .Q_N(_1039_),
    .Q(\pulse_width_counter_module.low_counter[15] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[16]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net215),
    .D(_0135_),
    .Q_N(_1038_),
    .Q(\pulse_width_counter_module.low_counter[16] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[17]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net216),
    .D(_0136_),
    .Q_N(_1037_),
    .Q(\pulse_width_counter_module.low_counter[17] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[18]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net217),
    .D(_0137_),
    .Q_N(_1036_),
    .Q(\pulse_width_counter_module.low_counter[18] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[19]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net218),
    .D(_0138_),
    .Q_N(_1035_),
    .Q(\pulse_width_counter_module.low_counter[19] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net219),
    .D(_0139_),
    .Q_N(_1034_),
    .Q(\pulse_width_counter_module.low_counter[1] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[20]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net220),
    .D(_0140_),
    .Q_N(_1033_),
    .Q(\pulse_width_counter_module.low_counter[20] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[21]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net221),
    .D(_0141_),
    .Q_N(_1032_),
    .Q(\pulse_width_counter_module.low_counter[21] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[22]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net222),
    .D(_0142_),
    .Q_N(_1031_),
    .Q(\pulse_width_counter_module.low_counter[22] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[23]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net223),
    .D(_0143_),
    .Q_N(_1030_),
    .Q(\pulse_width_counter_module.low_counter[23] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[24]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net224),
    .D(_0144_),
    .Q_N(_1029_),
    .Q(\pulse_width_counter_module.low_counter[24] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[25]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net225),
    .D(_0145_),
    .Q_N(_1028_),
    .Q(\pulse_width_counter_module.low_counter[25] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[26]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net226),
    .D(_0146_),
    .Q_N(_1027_),
    .Q(\pulse_width_counter_module.low_counter[26] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[27]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net227),
    .D(_0147_),
    .Q_N(_1026_),
    .Q(\pulse_width_counter_module.low_counter[27] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[28]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net228),
    .D(_0148_),
    .Q_N(_1025_),
    .Q(\pulse_width_counter_module.low_counter[28] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[29]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net229),
    .D(_0149_),
    .Q_N(_1024_),
    .Q(\pulse_width_counter_module.low_counter[29] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net230),
    .D(_0150_),
    .Q_N(_1023_),
    .Q(\pulse_width_counter_module.low_counter[2] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[30]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net231),
    .D(_0151_),
    .Q_N(_1022_),
    .Q(\pulse_width_counter_module.low_counter[30] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[31]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net232),
    .D(_0152_),
    .Q_N(_1021_),
    .Q(\pulse_width_counter_module.low_counter[31] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net233),
    .D(_0153_),
    .Q_N(_1020_),
    .Q(\pulse_width_counter_module.low_counter[3] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net234),
    .D(_0154_),
    .Q_N(_1019_),
    .Q(\pulse_width_counter_module.low_counter[4] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net235),
    .D(_0155_),
    .Q_N(_1018_),
    .Q(\pulse_width_counter_module.low_counter[5] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net236),
    .D(_0156_),
    .Q_N(_1017_),
    .Q(\pulse_width_counter_module.low_counter[6] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[7]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net237),
    .D(_0157_),
    .Q_N(_1016_),
    .Q(\pulse_width_counter_module.low_counter[7] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[8]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net238),
    .D(_0158_),
    .Q_N(_1015_),
    .Q(\pulse_width_counter_module.low_counter[8] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.low_counter[9]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net239),
    .D(_0159_),
    .Q_N(_1014_),
    .Q(\pulse_width_counter_module.low_counter[9] ));
 sg13g2_dfrbp_1 \pulse_width_counter_module.previous_freq_in$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net240),
    .D(_0160_),
    .Q_N(_1013_),
    .Q(\pulse_width_counter_module.previous_freq_in ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout10 (.A(_0894_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_0869_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0541_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0538_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0528_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0513_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0456_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_1010_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0988_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0986_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0964_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0962_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0940_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0935_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0903_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0880_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0836_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0724_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0579_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0569_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0512_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0455_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0451_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0285_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0939_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0319_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0195_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0996_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0973_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0948_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0920_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0898_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0873_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0846_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0821_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0525_),
    .X(net45));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(_0395_));
 sg13g2_buf_4 fanout47 (.X(net47),
    .A(_0394_));
 sg13g2_buf_4 fanout48 (.X(net48),
    .A(_0392_));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(_0390_));
 sg13g2_buf_2 fanout50 (.A(_0388_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0937_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0704_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0699_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0698_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0604_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0592_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0583_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0568_),
    .X(net58));
 sg13g2_buf_1 fanout59 (.A(_0524_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0492_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0446_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0386_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0526_),
    .X(net63));
 sg13g2_tielo _2199__64 (.L_LO(net64));
 sg13g2_tielo _2200__65 (.L_LO(net65));
 sg13g2_tielo _2201__66 (.L_LO(net66));
 sg13g2_tielo _2202__67 (.L_LO(net67));
 sg13g2_tielo _2203__68 (.L_LO(net68));
 sg13g2_tielo _2204__69 (.L_LO(net69));
 sg13g2_tielo _2205__70 (.L_LO(net70));
 sg13g2_tielo _2206__71 (.L_LO(net71));
 sg13g2_tielo _2207__72 (.L_LO(net72));
 sg13g2_tielo _2208__73 (.L_LO(net73));
 sg13g2_tielo _2209__74 (.L_LO(net74));
 sg13g2_tielo _2210__75 (.L_LO(net75));
 sg13g2_tielo _2211__76 (.L_LO(net76));
 sg13g2_tielo _2212__77 (.L_LO(net77));
 sg13g2_tielo _2213__78 (.L_LO(net78));
 sg13g2_tielo _2214__79 (.L_LO(net79));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[10]$_SDFFE_PN0P__81  (.L_HI(net81));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[11]$_SDFFE_PN0P__82  (.L_HI(net82));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[12]$_SDFFE_PN0P__83  (.L_HI(net83));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[13]$_SDFFE_PN0P__84  (.L_HI(net84));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[14]$_SDFFE_PN0P__85  (.L_HI(net85));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[15]$_SDFFE_PN0P__86  (.L_HI(net86));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[16]$_SDFFE_PN0P__87  (.L_HI(net87));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[17]$_SDFFE_PN0P__88  (.L_HI(net88));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[18]$_SDFFE_PN0P__89  (.L_HI(net89));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[19]$_SDFFE_PN0P__90  (.L_HI(net90));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[1]$_SDFFE_PN0P__91  (.L_HI(net91));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[20]$_SDFFE_PN0P__92  (.L_HI(net92));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[21]$_SDFFE_PN0P__93  (.L_HI(net93));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[22]$_SDFFE_PN0P__94  (.L_HI(net94));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[23]$_SDFFE_PN0P__95  (.L_HI(net95));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[24]$_SDFFE_PN0P__96  (.L_HI(net96));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[25]$_SDFFE_PN0P__97  (.L_HI(net97));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[26]$_SDFFE_PN0P__98  (.L_HI(net98));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[27]$_SDFFE_PN0P__99  (.L_HI(net99));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[28]$_SDFFE_PN0P__100  (.L_HI(net100));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[29]$_SDFFE_PN0P__101  (.L_HI(net101));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[2]$_SDFFE_PN0P__102  (.L_HI(net102));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[30]$_SDFFE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[31]$_SDFFE_PN0P__104  (.L_HI(net104));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[3]$_SDFFE_PN0P__105  (.L_HI(net105));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[4]$_SDFFE_PN0P__106  (.L_HI(net106));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[5]$_SDFFE_PN0P__107  (.L_HI(net107));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[6]$_SDFFE_PN0P__108  (.L_HI(net108));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[7]$_SDFFE_PN0P__109  (.L_HI(net109));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[8]$_SDFFE_PN0P__110  (.L_HI(net110));
 sg13g2_tiehi \pulse_width_counter_module.PERIOD[9]$_SDFFE_PN0P__111  (.L_HI(net111));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[0]$_SDFFE_PN0P__112  (.L_HI(net112));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[10]$_SDFFE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[11]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[12]$_SDFFE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[13]$_SDFFE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[14]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[15]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[16]$_SDFFE_PN0P__119  (.L_HI(net119));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[17]$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[18]$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[19]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[1]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[20]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[21]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[22]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[23]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[24]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[25]$_SDFFE_PN0P__129  (.L_HI(net129));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[26]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[27]$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[28]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[29]$_SDFFE_PN0P__133  (.L_HI(net133));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[2]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[30]$_SDFFE_PN0P__135  (.L_HI(net135));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[31]$_SDFFE_PN0P__136  (.L_HI(net136));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[3]$_SDFFE_PN0P__137  (.L_HI(net137));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[4]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[5]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[6]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[7]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[8]$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \pulse_width_counter_module.TIME_HIGH[9]$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[0]$_SDFFE_PN0P__144  (.L_HI(net144));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[10]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[11]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[12]$_SDFFE_PN0P__147  (.L_HI(net147));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[13]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[14]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[15]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[16]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[17]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[18]$_SDFFE_PN0P__153  (.L_HI(net153));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[19]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[1]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[20]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[21]$_SDFFE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[22]$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[23]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[24]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[25]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[26]$_SDFFE_PN0P__162  (.L_HI(net162));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[27]$_SDFFE_PN0P__163  (.L_HI(net163));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[28]$_SDFFE_PN0P__164  (.L_HI(net164));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[29]$_SDFFE_PN0P__165  (.L_HI(net165));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[2]$_SDFFE_PN0P__166  (.L_HI(net166));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[30]$_SDFFE_PN0P__167  (.L_HI(net167));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[31]$_SDFFE_PN0P__168  (.L_HI(net168));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[3]$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[4]$_SDFFE_PN0P__170  (.L_HI(net170));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[5]$_SDFFE_PN0P__171  (.L_HI(net171));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[6]$_SDFFE_PN0P__172  (.L_HI(net172));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[7]$_SDFFE_PN0P__173  (.L_HI(net173));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[8]$_SDFFE_PN0P__174  (.L_HI(net174));
 sg13g2_tiehi \pulse_width_counter_module.TIME_LOW[9]$_SDFFE_PN0P__175  (.L_HI(net175));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[0]$_SDFFE_PN0P__176  (.L_HI(net176));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[10]$_SDFFE_PN0P__177  (.L_HI(net177));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[11]$_SDFFE_PN0P__178  (.L_HI(net178));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[12]$_SDFFE_PN0P__179  (.L_HI(net179));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[13]$_SDFFE_PN0P__180  (.L_HI(net180));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[14]$_SDFFE_PN0P__181  (.L_HI(net181));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[15]$_SDFFE_PN0P__182  (.L_HI(net182));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[16]$_SDFFE_PN0P__183  (.L_HI(net183));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[17]$_SDFFE_PN0P__184  (.L_HI(net184));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[18]$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[19]$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[1]$_SDFFE_PN0P__187  (.L_HI(net187));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[20]$_SDFFE_PN0P__188  (.L_HI(net188));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[21]$_SDFFE_PN0P__189  (.L_HI(net189));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[22]$_SDFFE_PN0P__190  (.L_HI(net190));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[23]$_SDFFE_PN0P__191  (.L_HI(net191));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[24]$_SDFFE_PN0P__192  (.L_HI(net192));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[25]$_SDFFE_PN0P__193  (.L_HI(net193));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[26]$_SDFFE_PN0P__194  (.L_HI(net194));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[27]$_SDFFE_PN0P__195  (.L_HI(net195));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[28]$_SDFFE_PN0P__196  (.L_HI(net196));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[29]$_SDFFE_PN0P__197  (.L_HI(net197));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[2]$_SDFFE_PN0P__198  (.L_HI(net198));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[30]$_SDFFE_PN0P__199  (.L_HI(net199));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[31]$_SDFFE_PN0P__200  (.L_HI(net200));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[3]$_SDFFE_PN0P__201  (.L_HI(net201));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[4]$_SDFFE_PN0P__202  (.L_HI(net202));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[5]$_SDFFE_PN0P__203  (.L_HI(net203));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[6]$_SDFFE_PN0P__204  (.L_HI(net204));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[7]$_SDFFE_PN0P__205  (.L_HI(net205));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[8]$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \pulse_width_counter_module.high_counter[9]$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[0]$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[10]$_SDFFE_PN0P__209  (.L_HI(net209));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[11]$_SDFFE_PN0P__210  (.L_HI(net210));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[12]$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[13]$_SDFFE_PN0P__212  (.L_HI(net212));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[14]$_SDFFE_PN0P__213  (.L_HI(net213));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[15]$_SDFFE_PN0P__214  (.L_HI(net214));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[16]$_SDFFE_PN0P__215  (.L_HI(net215));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[17]$_SDFFE_PN0P__216  (.L_HI(net216));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[18]$_SDFFE_PN0P__217  (.L_HI(net217));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[19]$_SDFFE_PN0P__218  (.L_HI(net218));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[1]$_SDFFE_PN0P__219  (.L_HI(net219));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[20]$_SDFFE_PN0P__220  (.L_HI(net220));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[21]$_SDFFE_PN0P__221  (.L_HI(net221));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[22]$_SDFFE_PN0P__222  (.L_HI(net222));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[23]$_SDFFE_PN0P__223  (.L_HI(net223));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[24]$_SDFFE_PN0P__224  (.L_HI(net224));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[25]$_SDFFE_PN0P__225  (.L_HI(net225));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[26]$_SDFFE_PN0P__226  (.L_HI(net226));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[27]$_SDFFE_PN0P__227  (.L_HI(net227));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[28]$_SDFFE_PN0P__228  (.L_HI(net228));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[29]$_SDFFE_PN0P__229  (.L_HI(net229));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[2]$_SDFFE_PN0P__230  (.L_HI(net230));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[30]$_SDFFE_PN0P__231  (.L_HI(net231));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[31]$_SDFFE_PN0P__232  (.L_HI(net232));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[3]$_SDFFE_PN0P__233  (.L_HI(net233));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[4]$_SDFFE_PN0P__234  (.L_HI(net234));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[5]$_SDFFE_PN0P__235  (.L_HI(net235));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[6]$_SDFFE_PN0P__236  (.L_HI(net236));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[7]$_SDFFE_PN0P__237  (.L_HI(net237));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[8]$_SDFFE_PN0P__238  (.L_HI(net238));
 sg13g2_tiehi \pulse_width_counter_module.low_counter[9]$_SDFFE_PN0P__239  (.L_HI(net239));
 sg13g2_tiehi \pulse_width_counter_module.previous_freq_in$_SDFF_PN0__240  (.L_HI(net240));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_117 ();
 sg13g2_fill_2 FILLER_0_124 ();
 sg13g2_fill_1 FILLER_0_126 ();
 sg13g2_fill_2 FILLER_0_153 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_4 FILLER_0_166 ();
 sg13g2_fill_2 FILLER_0_206 ();
 sg13g2_fill_1 FILLER_0_208 ();
 sg13g2_fill_2 FILLER_0_239 ();
 sg13g2_fill_1 FILLER_0_241 ();
 sg13g2_fill_2 FILLER_0_272 ();
 sg13g2_fill_1 FILLER_0_300 ();
 sg13g2_fill_1 FILLER_0_305 ();
 sg13g2_fill_1 FILLER_0_332 ();
 sg13g2_fill_2 FILLER_0_337 ();
 sg13g2_decap_4 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_8 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_0_414 ();
 sg13g2_decap_8 FILLER_0_421 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_fill_2 FILLER_1_104 ();
 sg13g2_fill_1 FILLER_1_106 ();
 sg13g2_decap_4 FILLER_1_117 ();
 sg13g2_fill_2 FILLER_1_121 ();
 sg13g2_fill_1 FILLER_1_133 ();
 sg13g2_decap_4 FILLER_1_138 ();
 sg13g2_fill_1 FILLER_1_142 ();
 sg13g2_decap_8 FILLER_1_195 ();
 sg13g2_decap_4 FILLER_1_202 ();
 sg13g2_fill_1 FILLER_1_206 ();
 sg13g2_decap_8 FILLER_1_225 ();
 sg13g2_decap_8 FILLER_1_232 ();
 sg13g2_fill_2 FILLER_1_239 ();
 sg13g2_decap_4 FILLER_1_251 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_fill_2 FILLER_1_273 ();
 sg13g2_fill_1 FILLER_1_275 ();
 sg13g2_decap_4 FILLER_1_285 ();
 sg13g2_fill_2 FILLER_1_289 ();
 sg13g2_fill_1 FILLER_1_296 ();
 sg13g2_fill_2 FILLER_1_301 ();
 sg13g2_fill_1 FILLER_1_308 ();
 sg13g2_fill_2 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_321 ();
 sg13g2_fill_2 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_decap_8 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_1_415 ();
 sg13g2_decap_8 FILLER_1_422 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_fill_1 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_fill_1 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_134 ();
 sg13g2_fill_2 FILLER_2_141 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_4 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_166 ();
 sg13g2_decap_4 FILLER_2_173 ();
 sg13g2_fill_2 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_188 ();
 sg13g2_decap_8 FILLER_2_195 ();
 sg13g2_decap_8 FILLER_2_202 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_4 FILLER_2_235 ();
 sg13g2_fill_1 FILLER_2_239 ();
 sg13g2_decap_8 FILLER_2_278 ();
 sg13g2_decap_4 FILLER_2_285 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_fill_2 FILLER_2_312 ();
 sg13g2_decap_4 FILLER_2_319 ();
 sg13g2_fill_2 FILLER_2_323 ();
 sg13g2_decap_4 FILLER_2_331 ();
 sg13g2_fill_1 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_4 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_8 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_2_412 ();
 sg13g2_decap_8 FILLER_2_419 ();
 sg13g2_decap_4 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_79 ();
 sg13g2_fill_1 FILLER_3_81 ();
 sg13g2_fill_2 FILLER_3_86 ();
 sg13g2_fill_1 FILLER_3_88 ();
 sg13g2_fill_2 FILLER_3_93 ();
 sg13g2_fill_1 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_100 ();
 sg13g2_decap_8 FILLER_3_107 ();
 sg13g2_decap_8 FILLER_3_118 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_167 ();
 sg13g2_fill_2 FILLER_3_200 ();
 sg13g2_fill_2 FILLER_3_238 ();
 sg13g2_fill_1 FILLER_3_240 ();
 sg13g2_fill_1 FILLER_3_259 ();
 sg13g2_decap_4 FILLER_3_264 ();
 sg13g2_fill_2 FILLER_3_268 ();
 sg13g2_fill_2 FILLER_3_300 ();
 sg13g2_fill_1 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_325 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_fill_2 FILLER_3_358 ();
 sg13g2_fill_1 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_fill_2 FILLER_4_35 ();
 sg13g2_fill_1 FILLER_4_37 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_4 FILLER_4_49 ();
 sg13g2_fill_1 FILLER_4_62 ();
 sg13g2_fill_1 FILLER_4_68 ();
 sg13g2_fill_1 FILLER_4_74 ();
 sg13g2_fill_1 FILLER_4_80 ();
 sg13g2_fill_1 FILLER_4_89 ();
 sg13g2_fill_1 FILLER_4_116 ();
 sg13g2_fill_1 FILLER_4_121 ();
 sg13g2_decap_4 FILLER_4_126 ();
 sg13g2_fill_1 FILLER_4_134 ();
 sg13g2_decap_8 FILLER_4_139 ();
 sg13g2_fill_2 FILLER_4_146 ();
 sg13g2_fill_2 FILLER_4_152 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_fill_2 FILLER_4_165 ();
 sg13g2_fill_1 FILLER_4_167 ();
 sg13g2_decap_8 FILLER_4_181 ();
 sg13g2_fill_1 FILLER_4_188 ();
 sg13g2_decap_4 FILLER_4_194 ();
 sg13g2_fill_2 FILLER_4_198 ();
 sg13g2_fill_2 FILLER_4_208 ();
 sg13g2_fill_1 FILLER_4_210 ();
 sg13g2_decap_4 FILLER_4_215 ();
 sg13g2_decap_8 FILLER_4_223 ();
 sg13g2_decap_8 FILLER_4_230 ();
 sg13g2_fill_2 FILLER_4_237 ();
 sg13g2_decap_8 FILLER_4_243 ();
 sg13g2_fill_2 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_270 ();
 sg13g2_fill_1 FILLER_4_277 ();
 sg13g2_fill_1 FILLER_4_288 ();
 sg13g2_fill_2 FILLER_4_293 ();
 sg13g2_fill_1 FILLER_4_295 ();
 sg13g2_fill_2 FILLER_4_301 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_fill_2 FILLER_4_314 ();
 sg13g2_fill_2 FILLER_4_323 ();
 sg13g2_decap_4 FILLER_4_351 ();
 sg13g2_fill_1 FILLER_4_355 ();
 sg13g2_fill_1 FILLER_4_361 ();
 sg13g2_fill_2 FILLER_4_366 ();
 sg13g2_fill_2 FILLER_4_378 ();
 sg13g2_fill_2 FILLER_4_384 ();
 sg13g2_fill_1 FILLER_4_386 ();
 sg13g2_fill_2 FILLER_4_391 ();
 sg13g2_fill_1 FILLER_4_393 ();
 sg13g2_decap_4 FILLER_4_425 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_4 FILLER_5_25 ();
 sg13g2_fill_2 FILLER_5_29 ();
 sg13g2_decap_4 FILLER_5_57 ();
 sg13g2_fill_1 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_80 ();
 sg13g2_decap_8 FILLER_5_87 ();
 sg13g2_decap_4 FILLER_5_98 ();
 sg13g2_fill_1 FILLER_5_102 ();
 sg13g2_decap_4 FILLER_5_107 ();
 sg13g2_fill_2 FILLER_5_119 ();
 sg13g2_fill_1 FILLER_5_121 ();
 sg13g2_fill_2 FILLER_5_162 ();
 sg13g2_fill_2 FILLER_5_190 ();
 sg13g2_fill_1 FILLER_5_192 ();
 sg13g2_fill_2 FILLER_5_202 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_fill_2 FILLER_5_237 ();
 sg13g2_fill_1 FILLER_5_239 ();
 sg13g2_decap_8 FILLER_5_262 ();
 sg13g2_decap_4 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_273 ();
 sg13g2_fill_2 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_fill_1 FILLER_5_299 ();
 sg13g2_fill_2 FILLER_5_304 ();
 sg13g2_fill_1 FILLER_5_306 ();
 sg13g2_fill_1 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_fill_2 FILLER_5_372 ();
 sg13g2_fill_1 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_fill_1 FILLER_5_393 ();
 sg13g2_fill_2 FILLER_5_404 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_4 FILLER_5_424 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_40 ();
 sg13g2_decap_8 FILLER_6_47 ();
 sg13g2_fill_1 FILLER_6_54 ();
 sg13g2_decap_8 FILLER_6_59 ();
 sg13g2_fill_2 FILLER_6_66 ();
 sg13g2_fill_2 FILLER_6_73 ();
 sg13g2_fill_1 FILLER_6_83 ();
 sg13g2_decap_8 FILLER_6_122 ();
 sg13g2_fill_2 FILLER_6_129 ();
 sg13g2_fill_1 FILLER_6_131 ();
 sg13g2_fill_2 FILLER_6_141 ();
 sg13g2_fill_1 FILLER_6_143 ();
 sg13g2_decap_8 FILLER_6_148 ();
 sg13g2_fill_2 FILLER_6_155 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_fill_2 FILLER_6_168 ();
 sg13g2_fill_1 FILLER_6_170 ();
 sg13g2_decap_4 FILLER_6_179 ();
 sg13g2_fill_2 FILLER_6_188 ();
 sg13g2_fill_2 FILLER_6_193 ();
 sg13g2_fill_1 FILLER_6_195 ();
 sg13g2_decap_4 FILLER_6_204 ();
 sg13g2_fill_2 FILLER_6_208 ();
 sg13g2_fill_1 FILLER_6_219 ();
 sg13g2_fill_2 FILLER_6_224 ();
 sg13g2_decap_4 FILLER_6_231 ();
 sg13g2_fill_2 FILLER_6_235 ();
 sg13g2_decap_4 FILLER_6_241 ();
 sg13g2_fill_2 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_285 ();
 sg13g2_decap_4 FILLER_6_292 ();
 sg13g2_fill_1 FILLER_6_309 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_4 FILLER_6_334 ();
 sg13g2_fill_1 FILLER_6_338 ();
 sg13g2_fill_1 FILLER_6_343 ();
 sg13g2_decap_4 FILLER_6_352 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_fill_1 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_2 FILLER_6_408 ();
 sg13g2_fill_1 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_11 ();
 sg13g2_decap_8 FILLER_7_18 ();
 sg13g2_fill_2 FILLER_7_40 ();
 sg13g2_fill_1 FILLER_7_42 ();
 sg13g2_decap_4 FILLER_7_104 ();
 sg13g2_fill_2 FILLER_7_108 ();
 sg13g2_decap_8 FILLER_7_114 ();
 sg13g2_decap_8 FILLER_7_121 ();
 sg13g2_decap_4 FILLER_7_128 ();
 sg13g2_fill_1 FILLER_7_132 ();
 sg13g2_fill_2 FILLER_7_169 ();
 sg13g2_fill_2 FILLER_7_180 ();
 sg13g2_fill_1 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_193 ();
 sg13g2_fill_1 FILLER_7_202 ();
 sg13g2_fill_1 FILLER_7_255 ();
 sg13g2_decap_8 FILLER_7_269 ();
 sg13g2_fill_2 FILLER_7_276 ();
 sg13g2_decap_4 FILLER_7_287 ();
 sg13g2_fill_2 FILLER_7_291 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_4 FILLER_7_304 ();
 sg13g2_fill_1 FILLER_7_308 ();
 sg13g2_fill_1 FILLER_7_314 ();
 sg13g2_decap_4 FILLER_7_323 ();
 sg13g2_fill_2 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_338 ();
 sg13g2_fill_1 FILLER_7_344 ();
 sg13g2_fill_2 FILLER_7_350 ();
 sg13g2_decap_4 FILLER_7_386 ();
 sg13g2_fill_2 FILLER_7_395 ();
 sg13g2_fill_2 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_fill_2 FILLER_8_79 ();
 sg13g2_decap_4 FILLER_8_99 ();
 sg13g2_decap_8 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_136 ();
 sg13g2_decap_8 FILLER_8_146 ();
 sg13g2_fill_2 FILLER_8_153 ();
 sg13g2_fill_2 FILLER_8_190 ();
 sg13g2_fill_1 FILLER_8_192 ();
 sg13g2_decap_4 FILLER_8_206 ();
 sg13g2_fill_2 FILLER_8_210 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_decap_8 FILLER_8_235 ();
 sg13g2_decap_4 FILLER_8_264 ();
 sg13g2_fill_2 FILLER_8_277 ();
 sg13g2_fill_1 FILLER_8_340 ();
 sg13g2_fill_2 FILLER_8_367 ();
 sg13g2_fill_2 FILLER_8_374 ();
 sg13g2_fill_1 FILLER_8_376 ();
 sg13g2_decap_4 FILLER_8_385 ();
 sg13g2_fill_2 FILLER_8_389 ();
 sg13g2_fill_1 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_8_409 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_4 ();
 sg13g2_fill_2 FILLER_9_82 ();
 sg13g2_fill_1 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_89 ();
 sg13g2_decap_8 FILLER_9_96 ();
 sg13g2_decap_8 FILLER_9_103 ();
 sg13g2_decap_8 FILLER_9_110 ();
 sg13g2_decap_8 FILLER_9_117 ();
 sg13g2_fill_2 FILLER_9_124 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_172 ();
 sg13g2_fill_2 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_185 ();
 sg13g2_fill_1 FILLER_9_187 ();
 sg13g2_decap_4 FILLER_9_192 ();
 sg13g2_fill_1 FILLER_9_196 ();
 sg13g2_fill_2 FILLER_9_223 ();
 sg13g2_decap_8 FILLER_9_251 ();
 sg13g2_decap_4 FILLER_9_258 ();
 sg13g2_decap_4 FILLER_9_267 ();
 sg13g2_fill_1 FILLER_9_280 ();
 sg13g2_fill_2 FILLER_9_285 ();
 sg13g2_fill_2 FILLER_9_292 ();
 sg13g2_decap_4 FILLER_9_298 ();
 sg13g2_fill_1 FILLER_9_302 ();
 sg13g2_fill_2 FILLER_9_311 ();
 sg13g2_decap_4 FILLER_9_317 ();
 sg13g2_fill_2 FILLER_9_326 ();
 sg13g2_decap_4 FILLER_9_332 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_fill_2 FILLER_9_370 ();
 sg13g2_fill_1 FILLER_9_372 ();
 sg13g2_decap_4 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_11 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_44 ();
 sg13g2_fill_2 FILLER_10_51 ();
 sg13g2_decap_4 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_65 ();
 sg13g2_fill_2 FILLER_10_75 ();
 sg13g2_fill_1 FILLER_10_77 ();
 sg13g2_fill_1 FILLER_10_104 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_4 FILLER_10_158 ();
 sg13g2_fill_2 FILLER_10_162 ();
 sg13g2_decap_8 FILLER_10_195 ();
 sg13g2_fill_1 FILLER_10_202 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_2 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_239 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_decap_4 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_fill_1 FILLER_10_330 ();
 sg13g2_fill_1 FILLER_10_336 ();
 sg13g2_fill_2 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_391 ();
 sg13g2_fill_1 FILLER_10_396 ();
 sg13g2_fill_1 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_4 FILLER_11_31 ();
 sg13g2_fill_2 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_fill_1 FILLER_11_87 ();
 sg13g2_decap_4 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_109 ();
 sg13g2_fill_2 FILLER_11_116 ();
 sg13g2_decap_4 FILLER_11_122 ();
 sg13g2_fill_2 FILLER_11_130 ();
 sg13g2_fill_1 FILLER_11_137 ();
 sg13g2_fill_2 FILLER_11_142 ();
 sg13g2_decap_8 FILLER_11_156 ();
 sg13g2_decap_4 FILLER_11_167 ();
 sg13g2_fill_2 FILLER_11_171 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_fill_2 FILLER_11_184 ();
 sg13g2_decap_4 FILLER_11_217 ();
 sg13g2_decap_4 FILLER_11_247 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_1 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_263 ();
 sg13g2_fill_2 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_279 ();
 sg13g2_decap_4 FILLER_11_291 ();
 sg13g2_fill_2 FILLER_11_295 ();
 sg13g2_fill_2 FILLER_11_331 ();
 sg13g2_fill_1 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_4 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_361 ();
 sg13g2_fill_1 FILLER_11_367 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_fill_1 FILLER_11_397 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_11_409 ();
 sg13g2_decap_8 FILLER_11_416 ();
 sg13g2_decap_8 FILLER_11_423 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_4 FILLER_12_18 ();
 sg13g2_fill_2 FILLER_12_31 ();
 sg13g2_decap_4 FILLER_12_37 ();
 sg13g2_fill_2 FILLER_12_54 ();
 sg13g2_fill_1 FILLER_12_56 ();
 sg13g2_fill_1 FILLER_12_62 ();
 sg13g2_decap_4 FILLER_12_79 ();
 sg13g2_fill_2 FILLER_12_83 ();
 sg13g2_decap_4 FILLER_12_116 ();
 sg13g2_fill_2 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_160 ();
 sg13g2_fill_1 FILLER_12_162 ();
 sg13g2_decap_4 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_176 ();
 sg13g2_fill_2 FILLER_12_196 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_fill_1 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_233 ();
 sg13g2_decap_4 FILLER_12_240 ();
 sg13g2_decap_4 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_253 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_fill_1 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_4 FILLER_12_380 ();
 sg13g2_decap_4 FILLER_12_389 ();
 sg13g2_fill_2 FILLER_12_393 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_2 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_414 ();
 sg13g2_decap_8 FILLER_12_421 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_fill_1 FILLER_13_31 ();
 sg13g2_fill_1 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_79 ();
 sg13g2_decap_4 FILLER_13_84 ();
 sg13g2_fill_2 FILLER_13_88 ();
 sg13g2_fill_2 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_104 ();
 sg13g2_fill_1 FILLER_13_141 ();
 sg13g2_fill_2 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_194 ();
 sg13g2_fill_2 FILLER_13_200 ();
 sg13g2_decap_4 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_fill_2 FILLER_13_261 ();
 sg13g2_fill_1 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_268 ();
 sg13g2_fill_2 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_decap_4 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_297 ();
 sg13g2_fill_2 FILLER_13_302 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_315 ();
 sg13g2_fill_2 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_decap_4 FILLER_13_350 ();
 sg13g2_fill_2 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_fill_1 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_37 ();
 sg13g2_decap_4 FILLER_14_44 ();
 sg13g2_decap_8 FILLER_14_52 ();
 sg13g2_fill_1 FILLER_14_59 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_decap_4 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_121 ();
 sg13g2_decap_8 FILLER_14_131 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_fill_2 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_decap_4 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_179 ();
 sg13g2_fill_2 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_225 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_fill_2 FILLER_14_241 ();
 sg13g2_fill_1 FILLER_14_248 ();
 sg13g2_decap_4 FILLER_14_283 ();
 sg13g2_fill_2 FILLER_14_287 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_307 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_decap_4 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_372 ();
 sg13g2_decap_8 FILLER_14_379 ();
 sg13g2_decap_4 FILLER_14_386 ();
 sg13g2_fill_1 FILLER_15_26 ();
 sg13g2_fill_2 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_44 ();
 sg13g2_fill_2 FILLER_15_81 ();
 sg13g2_fill_1 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_110 ();
 sg13g2_decap_4 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_145 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_180 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_209 ();
 sg13g2_fill_2 FILLER_15_214 ();
 sg13g2_decap_4 FILLER_15_225 ();
 sg13g2_decap_4 FILLER_15_235 ();
 sg13g2_fill_2 FILLER_15_243 ();
 sg13g2_decap_4 FILLER_15_250 ();
 sg13g2_fill_2 FILLER_15_254 ();
 sg13g2_fill_2 FILLER_15_274 ();
 sg13g2_fill_1 FILLER_15_281 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_fill_1 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_298 ();
 sg13g2_decap_4 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_309 ();
 sg13g2_fill_2 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_341 ();
 sg13g2_decap_4 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_404 ();
 sg13g2_decap_8 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_11 ();
 sg13g2_fill_2 FILLER_16_29 ();
 sg13g2_fill_1 FILLER_16_31 ();
 sg13g2_decap_8 FILLER_16_37 ();
 sg13g2_decap_8 FILLER_16_44 ();
 sg13g2_fill_1 FILLER_16_51 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_4 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_71 ();
 sg13g2_fill_2 FILLER_16_77 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_121 ();
 sg13g2_decap_4 FILLER_16_128 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_fill_2 FILLER_16_148 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_160 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_decap_8 FILLER_16_174 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_decap_4 FILLER_16_194 ();
 sg13g2_fill_1 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_205 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_decap_4 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_253 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_4 FILLER_16_283 ();
 sg13g2_fill_2 FILLER_16_292 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_fill_2 FILLER_16_346 ();
 sg13g2_fill_2 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_8 FILLER_16_404 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_41 ();
 sg13g2_decap_8 FILLER_17_47 ();
 sg13g2_fill_2 FILLER_17_54 ();
 sg13g2_fill_1 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_60 ();
 sg13g2_decap_8 FILLER_17_65 ();
 sg13g2_fill_2 FILLER_17_72 ();
 sg13g2_fill_1 FILLER_17_74 ();
 sg13g2_fill_2 FILLER_17_86 ();
 sg13g2_fill_2 FILLER_17_93 ();
 sg13g2_decap_4 FILLER_17_103 ();
 sg13g2_decap_8 FILLER_17_172 ();
 sg13g2_fill_2 FILLER_17_193 ();
 sg13g2_decap_4 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_207 ();
 sg13g2_fill_1 FILLER_17_212 ();
 sg13g2_decap_4 FILLER_17_217 ();
 sg13g2_fill_1 FILLER_17_221 ();
 sg13g2_fill_2 FILLER_17_227 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_4 FILLER_17_245 ();
 sg13g2_fill_2 FILLER_17_249 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_fill_2 FILLER_17_289 ();
 sg13g2_fill_1 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_fill_2 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_17_386 ();
 sg13g2_fill_1 FILLER_17_388 ();
 sg13g2_decap_4 FILLER_18_26 ();
 sg13g2_fill_1 FILLER_18_34 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_fill_2 FILLER_18_100 ();
 sg13g2_decap_4 FILLER_18_107 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_122 ();
 sg13g2_decap_4 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_137 ();
 sg13g2_fill_2 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_153 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_decap_8 FILLER_18_166 ();
 sg13g2_decap_8 FILLER_18_173 ();
 sg13g2_decap_4 FILLER_18_180 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_decap_4 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_fill_1 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_decap_4 FILLER_18_358 ();
 sg13g2_fill_1 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_4 FILLER_18_374 ();
 sg13g2_fill_2 FILLER_18_412 ();
 sg13g2_decap_8 FILLER_18_419 ();
 sg13g2_decap_4 FILLER_18_426 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_15 ();
 sg13g2_decap_4 FILLER_19_22 ();
 sg13g2_decap_8 FILLER_19_38 ();
 sg13g2_decap_8 FILLER_19_45 ();
 sg13g2_decap_8 FILLER_19_52 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_fill_1 FILLER_19_66 ();
 sg13g2_fill_2 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_85 ();
 sg13g2_decap_4 FILLER_19_90 ();
 sg13g2_fill_2 FILLER_19_94 ();
 sg13g2_decap_4 FILLER_19_101 ();
 sg13g2_fill_2 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_164 ();
 sg13g2_decap_8 FILLER_19_178 ();
 sg13g2_decap_4 FILLER_19_185 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_fill_1 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_215 ();
 sg13g2_decap_4 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_229 ();
 sg13g2_decap_8 FILLER_19_236 ();
 sg13g2_decap_8 FILLER_19_243 ();
 sg13g2_decap_4 FILLER_19_254 ();
 sg13g2_fill_1 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_267 ();
 sg13g2_fill_1 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_decap_4 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_fill_2 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_fill_1 FILLER_19_359 ();
 sg13g2_fill_1 FILLER_19_364 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_fill_1 FILLER_19_374 ();
 sg13g2_fill_2 FILLER_19_380 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_387 ();
 sg13g2_fill_2 FILLER_19_392 ();
 sg13g2_fill_1 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_20_34 ();
 sg13g2_fill_2 FILLER_20_41 ();
 sg13g2_fill_1 FILLER_20_47 ();
 sg13g2_decap_8 FILLER_20_113 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_8 FILLER_20_138 ();
 sg13g2_decap_8 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_157 ();
 sg13g2_decap_8 FILLER_20_164 ();
 sg13g2_fill_2 FILLER_20_171 ();
 sg13g2_fill_1 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_183 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_decap_4 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_205 ();
 sg13g2_decap_8 FILLER_20_243 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_fill_1 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_decap_8 FILLER_20_327 ();
 sg13g2_decap_4 FILLER_20_334 ();
 sg13g2_fill_1 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_354 ();
 sg13g2_decap_4 FILLER_20_385 ();
 sg13g2_fill_1 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_fill_2 FILLER_20_402 ();
 sg13g2_fill_2 FILLER_20_409 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_21 ();
 sg13g2_fill_1 FILLER_21_27 ();
 sg13g2_fill_2 FILLER_21_33 ();
 sg13g2_fill_1 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_40 ();
 sg13g2_decap_4 FILLER_21_47 ();
 sg13g2_fill_2 FILLER_21_51 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_104 ();
 sg13g2_decap_4 FILLER_21_109 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_decap_4 FILLER_21_124 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_2 FILLER_21_186 ();
 sg13g2_fill_1 FILLER_21_188 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_4 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_4 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_342 ();
 sg13g2_decap_4 FILLER_21_352 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_fill_2 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_370 ();
 sg13g2_fill_1 FILLER_21_377 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_65 ();
 sg13g2_fill_2 FILLER_22_92 ();
 sg13g2_decap_4 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_fill_1 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_195 ();
 sg13g2_decap_8 FILLER_22_202 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_229 ();
 sg13g2_decap_4 FILLER_22_236 ();
 sg13g2_decap_4 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_270 ();
 sg13g2_decap_4 FILLER_22_292 ();
 sg13g2_decap_4 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_305 ();
 sg13g2_decap_4 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_4 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_22_414 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_18 ();
 sg13g2_fill_2 FILLER_23_34 ();
 sg13g2_fill_1 FILLER_23_36 ();
 sg13g2_fill_2 FILLER_23_58 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_decap_4 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_decap_4 FILLER_23_82 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_114 ();
 sg13g2_fill_2 FILLER_23_120 ();
 sg13g2_decap_8 FILLER_23_148 ();
 sg13g2_decap_8 FILLER_23_155 ();
 sg13g2_fill_2 FILLER_23_170 ();
 sg13g2_decap_4 FILLER_23_180 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_fill_2 FILLER_23_251 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_fill_2 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_352 ();
 sg13g2_decap_4 FILLER_23_359 ();
 sg13g2_fill_2 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_370 ();
 sg13g2_decap_4 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_389 ();
 sg13g2_decap_4 FILLER_23_399 ();
 sg13g2_fill_1 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_24_26 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_72 ();
 sg13g2_fill_2 FILLER_24_79 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_2 FILLER_24_115 ();
 sg13g2_decap_8 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_132 ();
 sg13g2_decap_8 FILLER_24_138 ();
 sg13g2_decap_8 FILLER_24_150 ();
 sg13g2_fill_2 FILLER_24_157 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_183 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_222 ();
 sg13g2_decap_4 FILLER_24_226 ();
 sg13g2_fill_2 FILLER_24_230 ();
 sg13g2_decap_4 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_decap_4 FILLER_24_305 ();
 sg13g2_fill_2 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_4 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_402 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_fill_2 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_33 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_44 ();
 sg13g2_fill_2 FILLER_25_51 ();
 sg13g2_decap_4 FILLER_25_57 ();
 sg13g2_decap_4 FILLER_25_90 ();
 sg13g2_fill_2 FILLER_25_94 ();
 sg13g2_decap_8 FILLER_25_100 ();
 sg13g2_decap_4 FILLER_25_107 ();
 sg13g2_fill_2 FILLER_25_120 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_decap_4 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_132 ();
 sg13g2_decap_4 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_156 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_229 ();
 sg13g2_decap_8 FILLER_25_267 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_fill_2 FILLER_25_330 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_fill_1 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_16 ();
 sg13g2_decap_8 FILLER_26_36 ();
 sg13g2_decap_8 FILLER_26_43 ();
 sg13g2_decap_8 FILLER_26_50 ();
 sg13g2_decap_8 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_64 ();
 sg13g2_fill_1 FILLER_26_83 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_decap_8 FILLER_26_92 ();
 sg13g2_decap_8 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_110 ();
 sg13g2_decap_4 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_160 ();
 sg13g2_decap_8 FILLER_26_173 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_193 ();
 sg13g2_decap_4 FILLER_26_200 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_237 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_decap_4 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_299 ();
 sg13g2_decap_4 FILLER_26_306 ();
 sg13g2_fill_2 FILLER_26_310 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_fill_2 FILLER_26_354 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_decap_4 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_371 ();
 sg13g2_fill_1 FILLER_26_376 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_27_71 ();
 sg13g2_fill_1 FILLER_27_73 ();
 sg13g2_decap_4 FILLER_27_124 ();
 sg13g2_decap_8 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_decap_4 FILLER_27_158 ();
 sg13g2_fill_1 FILLER_27_162 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_decap_8 FILLER_27_176 ();
 sg13g2_decap_4 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_207 ();
 sg13g2_decap_4 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_218 ();
 sg13g2_fill_2 FILLER_27_241 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_275 ();
 sg13g2_fill_2 FILLER_27_290 ();
 sg13g2_fill_1 FILLER_27_292 ();
 sg13g2_fill_1 FILLER_27_307 ();
 sg13g2_decap_4 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_338 ();
 sg13g2_fill_2 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_decap_4 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_decap_4 FILLER_27_397 ();
 sg13g2_fill_1 FILLER_27_401 ();
 sg13g2_decap_8 FILLER_27_414 ();
 sg13g2_decap_8 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_9 ();
 sg13g2_fill_2 FILLER_28_16 ();
 sg13g2_fill_1 FILLER_28_18 ();
 sg13g2_fill_1 FILLER_28_24 ();
 sg13g2_decap_4 FILLER_28_40 ();
 sg13g2_fill_2 FILLER_28_44 ();
 sg13g2_decap_4 FILLER_28_50 ();
 sg13g2_fill_1 FILLER_28_54 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_4 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_decap_4 FILLER_28_109 ();
 sg13g2_fill_2 FILLER_28_113 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_121 ();
 sg13g2_fill_2 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_154 ();
 sg13g2_fill_2 FILLER_28_163 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_4 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_201 ();
 sg13g2_fill_2 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_237 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_decap_4 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_276 ();
 sg13g2_decap_4 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_308 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_fill_2 FILLER_28_342 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_372 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_decap_4 FILLER_28_385 ();
 sg13g2_fill_2 FILLER_28_389 ();
 sg13g2_decap_4 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_416 ();
 sg13g2_decap_8 FILLER_28_423 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_34 ();
 sg13g2_fill_2 FILLER_29_41 ();
 sg13g2_fill_1 FILLER_29_43 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_decap_4 FILLER_29_86 ();
 sg13g2_fill_2 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_99 ();
 sg13g2_decap_8 FILLER_29_104 ();
 sg13g2_decap_8 FILLER_29_111 ();
 sg13g2_decap_4 FILLER_29_118 ();
 sg13g2_fill_1 FILLER_29_122 ();
 sg13g2_decap_8 FILLER_29_128 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_fill_2 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_205 ();
 sg13g2_decap_8 FILLER_29_212 ();
 sg13g2_decap_4 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_223 ();
 sg13g2_decap_4 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_237 ();
 sg13g2_decap_4 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_decap_8 FILLER_29_275 ();
 sg13g2_decap_4 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_4 FILLER_29_371 ();
 sg13g2_fill_2 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_2 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_52 ();
 sg13g2_decap_4 FILLER_30_57 ();
 sg13g2_decap_8 FILLER_30_79 ();
 sg13g2_decap_8 FILLER_30_86 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_185 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_decap_4 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_216 ();
 sg13g2_decap_4 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_299 ();
 sg13g2_decap_8 FILLER_30_306 ();
 sg13g2_decap_4 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_327 ();
 sg13g2_decap_4 FILLER_30_334 ();
 sg13g2_decap_8 FILLER_30_351 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_365 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_fill_2 FILLER_30_385 ();
 sg13g2_fill_1 FILLER_30_392 ();
 sg13g2_decap_4 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_30_414 ();
 sg13g2_decap_8 FILLER_30_421 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_decap_8 FILLER_31_9 ();
 sg13g2_decap_8 FILLER_31_16 ();
 sg13g2_decap_4 FILLER_31_23 ();
 sg13g2_decap_8 FILLER_31_31 ();
 sg13g2_decap_4 FILLER_31_38 ();
 sg13g2_fill_1 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_58 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_114 ();
 sg13g2_decap_8 FILLER_31_121 ();
 sg13g2_decap_4 FILLER_31_128 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_218 ();
 sg13g2_decap_4 FILLER_31_225 ();
 sg13g2_decap_4 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_242 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_289 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_decap_4 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_decap_4 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_decap_4 FILLER_31_355 ();
 sg13g2_fill_2 FILLER_31_385 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_fill_2 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_12 ();
 sg13g2_fill_1 FILLER_32_16 ();
 sg13g2_fill_1 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_71 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_88 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_decap_4 FILLER_32_131 ();
 sg13g2_fill_1 FILLER_32_135 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_4 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_decap_4 FILLER_32_173 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_234 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_294 ();
 sg13g2_decap_4 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_4 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_32_377 ();
 sg13g2_fill_1 FILLER_32_384 ();
 sg13g2_decap_4 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_fill_2 FILLER_33_26 ();
 sg13g2_fill_2 FILLER_33_32 ();
 sg13g2_fill_1 FILLER_33_34 ();
 sg13g2_fill_1 FILLER_33_53 ();
 sg13g2_fill_2 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_fill_2 FILLER_33_92 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_decap_8 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_106 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_decap_8 FILLER_33_164 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_185 ();
 sg13g2_decap_8 FILLER_33_192 ();
 sg13g2_decap_4 FILLER_33_199 ();
 sg13g2_fill_2 FILLER_33_207 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_4 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_262 ();
 sg13g2_decap_8 FILLER_33_269 ();
 sg13g2_decap_8 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_decap_8 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_decap_4 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_2 FILLER_33_378 ();
 sg13g2_fill_1 FILLER_33_380 ();
 sg13g2_fill_1 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_29 ();
 sg13g2_decap_4 FILLER_34_36 ();
 sg13g2_fill_1 FILLER_34_46 ();
 sg13g2_fill_1 FILLER_34_52 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_decap_8 FILLER_34_67 ();
 sg13g2_decap_8 FILLER_34_74 ();
 sg13g2_decap_4 FILLER_34_81 ();
 sg13g2_decap_4 FILLER_34_94 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_134 ();
 sg13g2_decap_8 FILLER_34_139 ();
 sg13g2_decap_8 FILLER_34_146 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_decap_8 FILLER_34_160 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_decap_4 FILLER_34_200 ();
 sg13g2_decap_4 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_decap_8 FILLER_34_241 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_decap_4 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_296 ();
 sg13g2_decap_8 FILLER_34_324 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_decap_8 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_345 ();
 sg13g2_decap_4 FILLER_34_352 ();
 sg13g2_fill_1 FILLER_34_364 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_fill_2 FILLER_34_374 ();
 sg13g2_fill_2 FILLER_34_384 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_fill_2 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_415 ();
 sg13g2_decap_8 FILLER_34_422 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_11 ();
 sg13g2_fill_1 FILLER_35_29 ();
 sg13g2_decap_4 FILLER_35_34 ();
 sg13g2_fill_1 FILLER_35_38 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_107 ();
 sg13g2_fill_2 FILLER_35_113 ();
 sg13g2_fill_2 FILLER_35_119 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_131 ();
 sg13g2_fill_1 FILLER_35_133 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_decap_4 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_183 ();
 sg13g2_decap_8 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_decap_4 FILLER_35_202 ();
 sg13g2_decap_8 FILLER_35_263 ();
 sg13g2_decap_4 FILLER_35_280 ();
 sg13g2_fill_2 FILLER_35_284 ();
 sg13g2_decap_4 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_304 ();
 sg13g2_decap_8 FILLER_35_311 ();
 sg13g2_decap_4 FILLER_35_318 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_4 FILLER_35_365 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_388 ();
 sg13g2_fill_1 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_418 ();
 sg13g2_decap_4 FILLER_35_425 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_fill_2 FILLER_36_31 ();
 sg13g2_fill_2 FILLER_36_38 ();
 sg13g2_fill_1 FILLER_36_40 ();
 sg13g2_fill_2 FILLER_36_45 ();
 sg13g2_fill_1 FILLER_36_47 ();
 sg13g2_fill_2 FILLER_36_54 ();
 sg13g2_fill_1 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_64 ();
 sg13g2_decap_4 FILLER_36_71 ();
 sg13g2_decap_8 FILLER_36_79 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_fill_2 FILLER_36_116 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_fill_2 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_fill_2 FILLER_36_131 ();
 sg13g2_fill_1 FILLER_36_133 ();
 sg13g2_fill_1 FILLER_36_139 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_decap_8 FILLER_36_150 ();
 sg13g2_decap_8 FILLER_36_157 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_230 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_243 ();
 sg13g2_decap_4 FILLER_36_250 ();
 sg13g2_decap_8 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_fill_1 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_15 ();
 sg13g2_fill_1 FILLER_37_22 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_4 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_decap_8 FILLER_37_54 ();
 sg13g2_decap_8 FILLER_37_92 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_decap_4 FILLER_37_131 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_4 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_181 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_212 ();
 sg13g2_decap_4 FILLER_37_219 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_fill_2 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_282 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_298 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_305 ();
 sg13g2_fill_1 FILLER_37_343 ();
 sg13g2_decap_4 FILLER_37_379 ();
 sg13g2_fill_2 FILLER_37_388 ();
 sg13g2_fill_1 FILLER_37_397 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_decap_8 FILLER_38_29 ();
 sg13g2_fill_1 FILLER_38_36 ();
 sg13g2_fill_2 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_decap_4 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_decap_4 FILLER_38_280 ();
 sg13g2_decap_4 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_314 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_decap_4 FILLER_38_334 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_344 ();
 sg13g2_decap_4 FILLER_38_351 ();
 sg13g2_fill_2 FILLER_38_355 ();
 sg13g2_fill_2 FILLER_38_361 ();
 sg13g2_decap_4 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
