module tt_um_gray_sobel (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire LFSR_enable_i_sync;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire clknet_leaf_0_clk;
 wire net202;
 wire \gray_sobel0.gray_scale0.nreset_i ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[0] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[1] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[2] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[3] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[4] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[5] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[6] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[7] ;
 wire \gray_sobel0.gray_scale0.px_rdy_i ;
 wire \gray_sobel0.gray_scale0.px_rdy_o ;
 wire \gray_sobel0.out_px_sobel[0] ;
 wire \gray_sobel0.out_px_sobel[1] ;
 wire \gray_sobel0.out_px_sobel[2] ;
 wire \gray_sobel0.out_px_sobel[3] ;
 wire \gray_sobel0.out_px_sobel[4] ;
 wire \gray_sobel0.out_px_sobel[5] ;
 wire \gray_sobel0.out_px_sobel[6] ;
 wire \gray_sobel0.out_px_sobel[7] ;
 wire \gray_sobel0.px_rdy_o_sobel ;
 wire \gray_sobel0.sobel0.counter_pixels[0] ;
 wire \gray_sobel0.sobel0.counter_pixels[10] ;
 wire \gray_sobel0.sobel0.counter_pixels[11] ;
 wire \gray_sobel0.sobel0.counter_pixels[12] ;
 wire \gray_sobel0.sobel0.counter_pixels[13] ;
 wire \gray_sobel0.sobel0.counter_pixels[14] ;
 wire \gray_sobel0.sobel0.counter_pixels[15] ;
 wire \gray_sobel0.sobel0.counter_pixels[16] ;
 wire \gray_sobel0.sobel0.counter_pixels[17] ;
 wire \gray_sobel0.sobel0.counter_pixels[18] ;
 wire \gray_sobel0.sobel0.counter_pixels[19] ;
 wire \gray_sobel0.sobel0.counter_pixels[1] ;
 wire \gray_sobel0.sobel0.counter_pixels[20] ;
 wire \gray_sobel0.sobel0.counter_pixels[21] ;
 wire \gray_sobel0.sobel0.counter_pixels[22] ;
 wire \gray_sobel0.sobel0.counter_pixels[23] ;
 wire \gray_sobel0.sobel0.counter_pixels[2] ;
 wire \gray_sobel0.sobel0.counter_pixels[3] ;
 wire \gray_sobel0.sobel0.counter_pixels[4] ;
 wire \gray_sobel0.sobel0.counter_pixels[5] ;
 wire \gray_sobel0.sobel0.counter_pixels[6] ;
 wire \gray_sobel0.sobel0.counter_pixels[7] ;
 wire \gray_sobel0.sobel0.counter_pixels[8] ;
 wire \gray_sobel0.sobel0.counter_pixels[9] ;
 wire \gray_sobel0.sobel0.counter_sobel[0] ;
 wire \gray_sobel0.sobel0.counter_sobel[1] ;
 wire \gray_sobel0.sobel0.counter_sobel[2] ;
 wire \gray_sobel0.sobel0.counter_sobel[3] ;
 wire \gray_sobel0.sobel0.fsm_state[0] ;
 wire \gray_sobel0.sobel0.fsm_state[1] ;
 wire \gray_sobel0.sobel0.next[0] ;
 wire \gray_sobel0.sobel0.next[1] ;
 wire \gray_sobel0.sobel0.px_ready ;
 wire \gray_sobel0.sobel0.sobel.pix0_0[0] ;
 wire \gray_sobel0.sobel0.sobel.pix0_0[1] ;
 wire \gray_sobel0.sobel0.sobel.pix0_0[2] ;
 wire \gray_sobel0.sobel0.sobel.pix0_0[3] ;
 wire \gray_sobel0.sobel0.sobel.pix0_0[4] ;
 wire \gray_sobel0.sobel0.sobel.pix0_0[5] ;
 wire \gray_sobel0.sobel0.sobel.pix0_0[6] ;
 wire \gray_sobel0.sobel0.sobel.pix0_0[7] ;
 wire \gray_sobel0.sobel0.sobel.pix0_1[0] ;
 wire \gray_sobel0.sobel0.sobel.pix0_1[1] ;
 wire \gray_sobel0.sobel0.sobel.pix0_1[2] ;
 wire \gray_sobel0.sobel0.sobel.pix0_1[3] ;
 wire \gray_sobel0.sobel0.sobel.pix0_1[4] ;
 wire \gray_sobel0.sobel0.sobel.pix0_1[5] ;
 wire \gray_sobel0.sobel0.sobel.pix0_1[6] ;
 wire \gray_sobel0.sobel0.sobel.pix0_1[7] ;
 wire \gray_sobel0.sobel0.sobel.pix0_2[0] ;
 wire \gray_sobel0.sobel0.sobel.pix0_2[1] ;
 wire \gray_sobel0.sobel0.sobel.pix0_2[2] ;
 wire \gray_sobel0.sobel0.sobel.pix0_2[3] ;
 wire \gray_sobel0.sobel0.sobel.pix0_2[4] ;
 wire \gray_sobel0.sobel0.sobel.pix0_2[5] ;
 wire \gray_sobel0.sobel0.sobel.pix0_2[6] ;
 wire \gray_sobel0.sobel0.sobel.pix0_2[7] ;
 wire \gray_sobel0.sobel0.sobel.pix1_0[0] ;
 wire \gray_sobel0.sobel0.sobel.pix1_0[1] ;
 wire \gray_sobel0.sobel0.sobel.pix1_0[2] ;
 wire \gray_sobel0.sobel0.sobel.pix1_0[3] ;
 wire \gray_sobel0.sobel0.sobel.pix1_0[4] ;
 wire \gray_sobel0.sobel0.sobel.pix1_0[5] ;
 wire \gray_sobel0.sobel0.sobel.pix1_0[6] ;
 wire \gray_sobel0.sobel0.sobel.pix1_0[7] ;
 wire \gray_sobel0.sobel0.sobel.pix1_1[0] ;
 wire \gray_sobel0.sobel0.sobel.pix1_1[1] ;
 wire \gray_sobel0.sobel0.sobel.pix1_1[2] ;
 wire \gray_sobel0.sobel0.sobel.pix1_1[3] ;
 wire \gray_sobel0.sobel0.sobel.pix1_1[4] ;
 wire \gray_sobel0.sobel0.sobel.pix1_1[5] ;
 wire \gray_sobel0.sobel0.sobel.pix1_1[6] ;
 wire \gray_sobel0.sobel0.sobel.pix1_1[7] ;
 wire \gray_sobel0.sobel0.sobel.pix1_2[0] ;
 wire \gray_sobel0.sobel0.sobel.pix1_2[1] ;
 wire \gray_sobel0.sobel0.sobel.pix1_2[2] ;
 wire \gray_sobel0.sobel0.sobel.pix1_2[3] ;
 wire \gray_sobel0.sobel0.sobel.pix1_2[4] ;
 wire \gray_sobel0.sobel0.sobel.pix1_2[5] ;
 wire \gray_sobel0.sobel0.sobel.pix1_2[6] ;
 wire \gray_sobel0.sobel0.sobel.pix1_2[7] ;
 wire \gray_sobel0.sobel0.sobel.pix2_0[0] ;
 wire \gray_sobel0.sobel0.sobel.pix2_0[1] ;
 wire \gray_sobel0.sobel0.sobel.pix2_0[2] ;
 wire \gray_sobel0.sobel0.sobel.pix2_0[3] ;
 wire \gray_sobel0.sobel0.sobel.pix2_0[4] ;
 wire \gray_sobel0.sobel0.sobel.pix2_0[5] ;
 wire \gray_sobel0.sobel0.sobel.pix2_0[6] ;
 wire \gray_sobel0.sobel0.sobel.pix2_0[7] ;
 wire \gray_sobel0.sobel0.sobel.pix2_1[0] ;
 wire \gray_sobel0.sobel0.sobel.pix2_1[1] ;
 wire \gray_sobel0.sobel0.sobel.pix2_1[2] ;
 wire \gray_sobel0.sobel0.sobel.pix2_1[3] ;
 wire \gray_sobel0.sobel0.sobel.pix2_1[4] ;
 wire \gray_sobel0.sobel0.sobel.pix2_1[5] ;
 wire \gray_sobel0.sobel0.sobel.pix2_1[6] ;
 wire \gray_sobel0.sobel0.sobel.pix2_1[7] ;
 wire \gray_sobel0.sobel0.sobel.pix2_2[0] ;
 wire \gray_sobel0.sobel0.sobel.pix2_2[1] ;
 wire \gray_sobel0.sobel0.sobel.pix2_2[2] ;
 wire \gray_sobel0.sobel0.sobel.pix2_2[3] ;
 wire \gray_sobel0.sobel0.sobel.pix2_2[4] ;
 wire \gray_sobel0.sobel0.sobel.pix2_2[5] ;
 wire \gray_sobel0.sobel0.sobel.pix2_2[6] ;
 wire \gray_sobel0.sobel0.sobel.pix2_2[7] ;
 wire in_data_rdy;
 wire in_lfsr_rdy;
 wire \input_data[0] ;
 wire \input_data[10] ;
 wire \input_data[11] ;
 wire \input_data[12] ;
 wire \input_data[13] ;
 wire \input_data[14] ;
 wire \input_data[15] ;
 wire \input_data[16] ;
 wire \input_data[17] ;
 wire \input_data[18] ;
 wire \input_data[19] ;
 wire \input_data[1] ;
 wire \input_data[20] ;
 wire \input_data[21] ;
 wire \input_data[22] ;
 wire \input_data[23] ;
 wire \input_data[2] ;
 wire \input_data[3] ;
 wire \input_data[4] ;
 wire \input_data[5] ;
 wire \input_data[6] ;
 wire \input_data[7] ;
 wire \input_data[8] ;
 wire \input_data[9] ;
 wire \lfsr0.config_done_o ;
 wire \lfsr0.config_i ;
 wire \lfsr0.lfsr_done ;
 wire \lfsr0.lfsr_en_i ;
 wire \lfsr0.lfsr_out[0] ;
 wire \lfsr0.lfsr_out[10] ;
 wire \lfsr0.lfsr_out[11] ;
 wire \lfsr0.lfsr_out[12] ;
 wire \lfsr0.lfsr_out[13] ;
 wire \lfsr0.lfsr_out[14] ;
 wire \lfsr0.lfsr_out[15] ;
 wire \lfsr0.lfsr_out[16] ;
 wire \lfsr0.lfsr_out[17] ;
 wire \lfsr0.lfsr_out[18] ;
 wire \lfsr0.lfsr_out[19] ;
 wire \lfsr0.lfsr_out[1] ;
 wire \lfsr0.lfsr_out[20] ;
 wire \lfsr0.lfsr_out[21] ;
 wire \lfsr0.lfsr_out[22] ;
 wire \lfsr0.lfsr_out[23] ;
 wire \lfsr0.lfsr_out[2] ;
 wire \lfsr0.lfsr_out[3] ;
 wire \lfsr0.lfsr_out[4] ;
 wire \lfsr0.lfsr_out[5] ;
 wire \lfsr0.lfsr_out[6] ;
 wire \lfsr0.lfsr_out[7] ;
 wire \lfsr0.lfsr_out[8] ;
 wire \lfsr0.lfsr_out[9] ;
 wire \lfsr0.lfsr_rdy_o ;
 wire \lfsr0.seed_reg[0] ;
 wire \lfsr0.seed_reg[10] ;
 wire \lfsr0.seed_reg[11] ;
 wire \lfsr0.seed_reg[12] ;
 wire \lfsr0.seed_reg[13] ;
 wire \lfsr0.seed_reg[14] ;
 wire \lfsr0.seed_reg[15] ;
 wire \lfsr0.seed_reg[16] ;
 wire \lfsr0.seed_reg[17] ;
 wire \lfsr0.seed_reg[18] ;
 wire \lfsr0.seed_reg[19] ;
 wire \lfsr0.seed_reg[1] ;
 wire \lfsr0.seed_reg[20] ;
 wire \lfsr0.seed_reg[21] ;
 wire \lfsr0.seed_reg[22] ;
 wire \lfsr0.seed_reg[23] ;
 wire \lfsr0.seed_reg[2] ;
 wire \lfsr0.seed_reg[3] ;
 wire \lfsr0.seed_reg[4] ;
 wire \lfsr0.seed_reg[5] ;
 wire \lfsr0.seed_reg[6] ;
 wire \lfsr0.seed_reg[7] ;
 wire \lfsr0.seed_reg[8] ;
 wire \lfsr0.seed_reg[9] ;
 wire \lfsr0.stop_reg[0] ;
 wire \lfsr0.stop_reg[10] ;
 wire \lfsr0.stop_reg[11] ;
 wire \lfsr0.stop_reg[12] ;
 wire \lfsr0.stop_reg[13] ;
 wire \lfsr0.stop_reg[14] ;
 wire \lfsr0.stop_reg[15] ;
 wire \lfsr0.stop_reg[16] ;
 wire \lfsr0.stop_reg[17] ;
 wire \lfsr0.stop_reg[18] ;
 wire \lfsr0.stop_reg[19] ;
 wire \lfsr0.stop_reg[1] ;
 wire \lfsr0.stop_reg[20] ;
 wire \lfsr0.stop_reg[21] ;
 wire \lfsr0.stop_reg[22] ;
 wire \lfsr0.stop_reg[23] ;
 wire \lfsr0.stop_reg[2] ;
 wire \lfsr0.stop_reg[3] ;
 wire \lfsr0.stop_reg[4] ;
 wire \lfsr0.stop_reg[5] ;
 wire \lfsr0.stop_reg[6] ;
 wire \lfsr0.stop_reg[7] ;
 wire \lfsr0.stop_reg[8] ;
 wire \lfsr0.stop_reg[9] ;
 wire \nreset_sync0.r_sync ;
 wire \sgnl_sync0.signal_sync ;
 wire \sgnl_sync1.signal_sync ;
 wire \sgnl_sync2.signal_sync ;
 wire \spi0.data_tx[0] ;
 wire \spi0.data_tx[10] ;
 wire \spi0.data_tx[11] ;
 wire \spi0.data_tx[12] ;
 wire \spi0.data_tx[13] ;
 wire \spi0.data_tx[14] ;
 wire \spi0.data_tx[15] ;
 wire \spi0.data_tx[16] ;
 wire \spi0.data_tx[17] ;
 wire \spi0.data_tx[18] ;
 wire \spi0.data_tx[19] ;
 wire \spi0.data_tx[1] ;
 wire \spi0.data_tx[20] ;
 wire \spi0.data_tx[21] ;
 wire \spi0.data_tx[22] ;
 wire \spi0.data_tx[23] ;
 wire \spi0.data_tx[2] ;
 wire \spi0.data_tx[3] ;
 wire \spi0.data_tx[4] ;
 wire \spi0.data_tx[5] ;
 wire \spi0.data_tx[6] ;
 wire \spi0.data_tx[7] ;
 wire \spi0.data_tx[8] ;
 wire \spi0.data_tx[9] ;
 wire \spi0.rxtx_done ;
 wire \spi0.rxtx_done_reg ;
 wire \spi0.rxtx_done_rising ;
 wire \spi0.signal_sync1.async_signal_i ;
 wire \spi0.signal_sync1.signal_sync ;
 wire \spi0.spi0.counter[0] ;
 wire \spi0.spi0.counter[1] ;
 wire \spi0.spi0.counter[2] ;
 wire \spi0.spi0.counter[3] ;
 wire \spi0.spi0.counter[4] ;
 wire \spi0.spi0.counter[5] ;
 wire \spi0.spi0.data_rx_o[0] ;
 wire \spi0.spi0.data_rx_o[10] ;
 wire \spi0.spi0.data_rx_o[11] ;
 wire \spi0.spi0.data_rx_o[12] ;
 wire \spi0.spi0.data_rx_o[13] ;
 wire \spi0.spi0.data_rx_o[14] ;
 wire \spi0.spi0.data_rx_o[15] ;
 wire \spi0.spi0.data_rx_o[16] ;
 wire \spi0.spi0.data_rx_o[17] ;
 wire \spi0.spi0.data_rx_o[18] ;
 wire \spi0.spi0.data_rx_o[19] ;
 wire \spi0.spi0.data_rx_o[1] ;
 wire \spi0.spi0.data_rx_o[20] ;
 wire \spi0.spi0.data_rx_o[21] ;
 wire \spi0.spi0.data_rx_o[22] ;
 wire \spi0.spi0.data_rx_o[23] ;
 wire \spi0.spi0.data_rx_o[2] ;
 wire \spi0.spi0.data_rx_o[3] ;
 wire \spi0.spi0.data_rx_o[4] ;
 wire \spi0.spi0.data_rx_o[5] ;
 wire \spi0.spi0.data_rx_o[6] ;
 wire \spi0.spi0.data_rx_o[7] ;
 wire \spi0.spi0.data_rx_o[8] ;
 wire \spi0.spi0.data_rx_o[9] ;
 wire \spi0.spi0.sdo_o ;
 wire \spi0.spi0.sdo_register[0] ;
 wire \spi0.spi0.sdo_register[10] ;
 wire \spi0.spi0.sdo_register[11] ;
 wire \spi0.spi0.sdo_register[12] ;
 wire \spi0.spi0.sdo_register[13] ;
 wire \spi0.spi0.sdo_register[14] ;
 wire \spi0.spi0.sdo_register[15] ;
 wire \spi0.spi0.sdo_register[16] ;
 wire \spi0.spi0.sdo_register[17] ;
 wire \spi0.spi0.sdo_register[18] ;
 wire \spi0.spi0.sdo_register[19] ;
 wire \spi0.spi0.sdo_register[1] ;
 wire \spi0.spi0.sdo_register[20] ;
 wire \spi0.spi0.sdo_register[21] ;
 wire \spi0.spi0.sdo_register[22] ;
 wire \spi0.spi0.sdo_register[2] ;
 wire \spi0.spi0.sdo_register[3] ;
 wire \spi0.spi0.sdo_register[4] ;
 wire \spi0.spi0.sdo_register[5] ;
 wire \spi0.spi0.sdo_register[6] ;
 wire \spi0.spi0.sdo_register[7] ;
 wire \spi0.spi0.sdo_register[8] ;
 wire \spi0.spi0.sdo_register[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_2 _2498_ (.A(\lfsr0.lfsr_out[4] ),
    .X(_1828_));
 sg13g2_xnor2_1 _2499_ (.Y(_1829_),
    .A(\lfsr0.stop_reg[4] ),
    .B(_1828_));
 sg13g2_xnor2_1 _2500_ (.Y(_1830_),
    .A(\lfsr0.stop_reg[19] ),
    .B(\lfsr0.lfsr_out[19] ));
 sg13g2_buf_1 _2501_ (.A(\lfsr0.lfsr_out[9] ),
    .X(_1831_));
 sg13g2_xnor2_1 _2502_ (.Y(_1832_),
    .A(\lfsr0.stop_reg[9] ),
    .B(_1831_));
 sg13g2_xnor2_1 _2503_ (.Y(_1833_),
    .A(\lfsr0.stop_reg[0] ),
    .B(\lfsr0.lfsr_out[0] ));
 sg13g2_nand4_1 _2504_ (.B(_1830_),
    .C(_1832_),
    .A(_1829_),
    .Y(_1834_),
    .D(_1833_));
 sg13g2_buf_1 _2505_ (.A(\lfsr0.lfsr_out[3] ),
    .X(_1835_));
 sg13g2_xnor2_1 _2506_ (.Y(_1836_),
    .A(\lfsr0.stop_reg[3] ),
    .B(_1835_));
 sg13g2_xnor2_1 _2507_ (.Y(_1837_),
    .A(\lfsr0.stop_reg[16] ),
    .B(\lfsr0.lfsr_out[16] ));
 sg13g2_xnor2_1 _2508_ (.Y(_1838_),
    .A(\lfsr0.stop_reg[13] ),
    .B(\lfsr0.lfsr_out[13] ));
 sg13g2_buf_1 _2509_ (.A(\lfsr0.lfsr_out[6] ),
    .X(_1839_));
 sg13g2_xnor2_1 _2510_ (.Y(_1840_),
    .A(\lfsr0.stop_reg[6] ),
    .B(net119));
 sg13g2_nand4_1 _2511_ (.B(_1837_),
    .C(_1838_),
    .A(_1836_),
    .Y(_1841_),
    .D(_1840_));
 sg13g2_buf_1 _2512_ (.A(\lfsr0.lfsr_out[12] ),
    .X(_1842_));
 sg13g2_xnor2_1 _2513_ (.Y(_1843_),
    .A(\lfsr0.stop_reg[12] ),
    .B(_1842_));
 sg13g2_xnor2_1 _2514_ (.Y(_1844_),
    .A(\lfsr0.stop_reg[1] ),
    .B(\lfsr0.lfsr_out[1] ));
 sg13g2_xnor2_1 _2515_ (.Y(_1845_),
    .A(\lfsr0.lfsr_out[23] ),
    .B(\lfsr0.stop_reg[23] ));
 sg13g2_buf_1 _2516_ (.A(\lfsr0.lfsr_out[18] ),
    .X(_1846_));
 sg13g2_xnor2_1 _2517_ (.Y(_1847_),
    .A(\lfsr0.stop_reg[18] ),
    .B(_1846_));
 sg13g2_nand4_1 _2518_ (.B(_1844_),
    .C(_1845_),
    .A(_1843_),
    .Y(_1848_),
    .D(_1847_));
 sg13g2_xnor2_1 _2519_ (.Y(_1849_),
    .A(\lfsr0.stop_reg[10] ),
    .B(\lfsr0.lfsr_out[10] ));
 sg13g2_buf_1 _2520_ (.A(\lfsr0.lfsr_out[5] ),
    .X(_1850_));
 sg13g2_xnor2_1 _2521_ (.Y(_1851_),
    .A(\lfsr0.stop_reg[5] ),
    .B(net117));
 sg13g2_xnor2_1 _2522_ (.Y(_1852_),
    .A(\lfsr0.stop_reg[22] ),
    .B(\lfsr0.lfsr_out[22] ));
 sg13g2_buf_1 _2523_ (.A(\lfsr0.lfsr_out[7] ),
    .X(_1853_));
 sg13g2_xnor2_1 _2524_ (.Y(_1854_),
    .A(\lfsr0.stop_reg[7] ),
    .B(net116));
 sg13g2_nand4_1 _2525_ (.B(_1851_),
    .C(_1852_),
    .A(_1849_),
    .Y(_1855_),
    .D(_1854_));
 sg13g2_nor4_1 _2526_ (.A(_1834_),
    .B(_1841_),
    .C(_1848_),
    .D(_1855_),
    .Y(_1856_));
 sg13g2_xor2_1 _2527_ (.B(\lfsr0.lfsr_out[2] ),
    .A(\lfsr0.stop_reg[2] ),
    .X(_1857_));
 sg13g2_xor2_1 _2528_ (.B(\lfsr0.lfsr_out[20] ),
    .A(\lfsr0.stop_reg[20] ),
    .X(_1858_));
 sg13g2_xor2_1 _2529_ (.B(\lfsr0.lfsr_out[8] ),
    .A(\lfsr0.stop_reg[8] ),
    .X(_1859_));
 sg13g2_xor2_1 _2530_ (.B(\lfsr0.lfsr_out[14] ),
    .A(\lfsr0.stop_reg[14] ),
    .X(_1860_));
 sg13g2_nor4_1 _2531_ (.A(_1857_),
    .B(_1858_),
    .C(_1859_),
    .D(_1860_),
    .Y(_1861_));
 sg13g2_xor2_1 _2532_ (.B(\lfsr0.lfsr_out[17] ),
    .A(\lfsr0.stop_reg[17] ),
    .X(_1862_));
 sg13g2_xor2_1 _2533_ (.B(\lfsr0.lfsr_out[15] ),
    .A(\lfsr0.stop_reg[15] ),
    .X(_1863_));
 sg13g2_xor2_1 _2534_ (.B(\lfsr0.lfsr_out[11] ),
    .A(\lfsr0.stop_reg[11] ),
    .X(_1864_));
 sg13g2_buf_2 _2535_ (.A(\lfsr0.lfsr_out[21] ),
    .X(_1865_));
 sg13g2_xor2_1 _2536_ (.B(_1865_),
    .A(\lfsr0.stop_reg[21] ),
    .X(_1866_));
 sg13g2_nor4_1 _2537_ (.A(_1862_),
    .B(_1863_),
    .C(_1864_),
    .D(_1866_),
    .Y(_1867_));
 sg13g2_nand3_1 _2538_ (.B(_1861_),
    .C(_1867_),
    .A(_1856_),
    .Y(_1868_));
 sg13g2_buf_1 _2539_ (.A(_1868_),
    .X(_1869_));
 sg13g2_buf_1 _2540_ (.A(_1869_),
    .X(_1870_));
 sg13g2_inv_1 _2541_ (.Y(\lfsr0.lfsr_done ),
    .A(net64));
 sg13g2_buf_1 _2542_ (.A(\lfsr0.lfsr_en_i ),
    .X(_1871_));
 sg13g2_buf_1 _2543_ (.A(_1871_),
    .X(_1872_));
 sg13g2_buf_1 _2544_ (.A(net94),
    .X(_1873_));
 sg13g2_buf_1 _2545_ (.A(_1869_),
    .X(_1874_));
 sg13g2_and2_1 _2546_ (.A(net79),
    .B(net63),
    .X(_0000_));
 sg13g2_nor2b_1 _2547_ (.A(\gray_sobel0.sobel0.fsm_state[0] ),
    .B_N(net6),
    .Y(_1875_));
 sg13g2_buf_1 _2548_ (.A(\gray_sobel0.sobel0.counter_pixels[17] ),
    .X(_1876_));
 sg13g2_buf_1 _2549_ (.A(\gray_sobel0.sobel0.counter_pixels[16] ),
    .X(_1877_));
 sg13g2_buf_1 _2550_ (.A(\gray_sobel0.sobel0.counter_pixels[19] ),
    .X(_1878_));
 sg13g2_buf_1 _2551_ (.A(\gray_sobel0.sobel0.counter_pixels[18] ),
    .X(_1879_));
 sg13g2_nor4_1 _2552_ (.A(_1876_),
    .B(_1877_),
    .C(_1878_),
    .D(_1879_),
    .Y(_1880_));
 sg13g2_buf_1 _2553_ (.A(\gray_sobel0.sobel0.counter_pixels[21] ),
    .X(_1881_));
 sg13g2_buf_1 _2554_ (.A(\gray_sobel0.sobel0.counter_pixels[20] ),
    .X(_1882_));
 sg13g2_buf_1 _2555_ (.A(\gray_sobel0.sobel0.counter_pixels[22] ),
    .X(_1883_));
 sg13g2_nor4_1 _2556_ (.A(_1881_),
    .B(_1882_),
    .C(\gray_sobel0.sobel0.counter_pixels[23] ),
    .D(_1883_),
    .Y(_1884_));
 sg13g2_buf_1 _2557_ (.A(\gray_sobel0.sobel0.counter_pixels[4] ),
    .X(_1885_));
 sg13g2_buf_1 _2558_ (.A(\gray_sobel0.sobel0.counter_pixels[7] ),
    .X(_1886_));
 sg13g2_nor4_1 _2559_ (.A(\gray_sobel0.sobel0.counter_pixels[5] ),
    .B(_1885_),
    .C(_1886_),
    .D(\gray_sobel0.sobel0.counter_pixels[6] ),
    .Y(_1887_));
 sg13g2_buf_1 _2560_ (.A(\gray_sobel0.sobel0.counter_pixels[15] ),
    .X(_1888_));
 sg13g2_buf_1 _2561_ (.A(\gray_sobel0.sobel0.counter_pixels[14] ),
    .X(_1889_));
 sg13g2_nor4_1 _2562_ (.A(\gray_sobel0.sobel0.counter_pixels[3] ),
    .B(\gray_sobel0.sobel0.counter_pixels[2] ),
    .C(_1888_),
    .D(_1889_),
    .Y(_1890_));
 sg13g2_nand4_1 _2563_ (.B(_1884_),
    .C(_1887_),
    .A(_1880_),
    .Y(_1891_),
    .D(_1890_));
 sg13g2_buf_1 _2564_ (.A(\gray_sobel0.sobel0.counter_pixels[8] ),
    .X(_1892_));
 sg13g2_buf_1 _2565_ (.A(\gray_sobel0.sobel0.counter_pixels[11] ),
    .X(_1893_));
 sg13g2_buf_1 _2566_ (.A(\gray_sobel0.sobel0.counter_pixels[10] ),
    .X(_1894_));
 sg13g2_buf_1 _2567_ (.A(\gray_sobel0.sobel0.counter_pixels[12] ),
    .X(_1895_));
 sg13g2_nor4_1 _2568_ (.A(_1892_),
    .B(_1893_),
    .C(_1894_),
    .D(_1895_),
    .Y(_1896_));
 sg13g2_buf_1 _2569_ (.A(\gray_sobel0.sobel0.counter_pixels[9] ),
    .X(_1897_));
 sg13g2_buf_1 _2570_ (.A(\gray_sobel0.sobel0.counter_pixels[13] ),
    .X(_1898_));
 sg13g2_buf_1 _2571_ (.A(\gray_sobel0.sobel0.counter_pixels[1] ),
    .X(_1899_));
 sg13g2_buf_2 _2572_ (.A(\gray_sobel0.sobel0.counter_pixels[0] ),
    .X(_1900_));
 sg13g2_nand2b_1 _2573_ (.Y(_1901_),
    .B(_1900_),
    .A_N(_1899_));
 sg13g2_nor3_1 _2574_ (.A(_1897_),
    .B(_1898_),
    .C(_1901_),
    .Y(_1902_));
 sg13g2_nand2_1 _2575_ (.Y(_1903_),
    .A(_1896_),
    .B(_1902_));
 sg13g2_nor2_1 _2576_ (.A(_1891_),
    .B(_1903_),
    .Y(_1904_));
 sg13g2_nor2b_1 _2577_ (.A(\gray_sobel0.sobel0.fsm_state[1] ),
    .B_N(\gray_sobel0.sobel0.fsm_state[0] ),
    .Y(_1905_));
 sg13g2_a22oi_1 _2578_ (.Y(_1906_),
    .B1(_1904_),
    .B2(_1905_),
    .A2(_1875_),
    .A1(\gray_sobel0.sobel0.fsm_state[1] ));
 sg13g2_buf_1 _2579_ (.A(_1906_),
    .X(_1907_));
 sg13g2_inv_2 _2580_ (.Y(_1908_),
    .A(_1907_));
 sg13g2_buf_1 _2581_ (.A(_1908_),
    .X(\gray_sobel0.sobel0.next[1] ));
 sg13g2_xnor2_1 _2582_ (.Y(_1909_),
    .A(net6),
    .B(\gray_sobel0.sobel0.fsm_state[1] ));
 sg13g2_o21ai_1 _2583_ (.B1(_1905_),
    .Y(_1910_),
    .A1(_1891_),
    .A2(_1903_));
 sg13g2_o21ai_1 _2584_ (.B1(_1910_),
    .Y(_1911_),
    .A1(\gray_sobel0.sobel0.fsm_state[0] ),
    .A2(_1909_));
 sg13g2_buf_1 _2585_ (.A(_1911_),
    .X(\gray_sobel0.sobel0.next[0] ));
 sg13g2_buf_2 _2586_ (.A(LFSR_enable_i_sync),
    .X(_1912_));
 sg13g2_buf_1 _2587_ (.A(_1912_),
    .X(_1913_));
 sg13g2_buf_1 _2588_ (.A(_1913_),
    .X(_1914_));
 sg13g2_mux2_1 _2589_ (.A0(in_data_rdy),
    .A1(\lfsr0.lfsr_rdy_o ),
    .S(_1914_),
    .X(\gray_sobel0.gray_scale0.px_rdy_i ));
 sg13g2_buf_1 _2590_ (.A(net78),
    .X(_1915_));
 sg13g2_buf_1 _2591_ (.A(net71),
    .X(_1916_));
 sg13g2_buf_1 _2592_ (.A(_1916_),
    .X(_1917_));
 sg13g2_and2_1 _2593_ (.A(_1917_),
    .B(in_data_rdy),
    .X(_1918_));
 sg13g2_buf_1 _2594_ (.A(_1918_),
    .X(in_lfsr_rdy));
 sg13g2_buf_1 _2595_ (.A(\spi0.spi0.counter[0] ),
    .X(_1919_));
 sg13g2_buf_1 _2596_ (.A(\spi0.spi0.counter[2] ),
    .X(_1920_));
 sg13g2_nor3_1 _2597_ (.A(_1919_),
    .B(_1920_),
    .C(\spi0.spi0.counter[5] ),
    .Y(_1921_));
 sg13g2_buf_1 _2598_ (.A(\spi0.spi0.counter[1] ),
    .X(_1922_));
 sg13g2_buf_1 _2599_ (.A(\spi0.spi0.counter[3] ),
    .X(_1923_));
 sg13g2_nand2_1 _2600_ (.Y(_1924_),
    .A(_1923_),
    .B(\spi0.spi0.counter[4] ));
 sg13g2_nor2_1 _2601_ (.A(_1922_),
    .B(_1924_),
    .Y(_1925_));
 sg13g2_and2_1 _2602_ (.A(_1921_),
    .B(_1925_),
    .X(_1926_));
 sg13g2_buf_2 _2603_ (.A(_1926_),
    .X(_1927_));
 sg13g2_buf_1 _2604_ (.A(_1927_),
    .X(_0008_));
 sg13g2_and2_1 _2605_ (.A(\spi0.data_tx[16] ),
    .B(net61),
    .X(_0009_));
 sg13g2_mux2_1 _2606_ (.A0(\spi0.spi0.sdo_register[0] ),
    .A1(\spi0.data_tx[17] ),
    .S(net61),
    .X(_0020_));
 sg13g2_mux2_1 _2607_ (.A0(\spi0.spi0.sdo_register[1] ),
    .A1(\spi0.data_tx[18] ),
    .S(net61),
    .X(_0025_));
 sg13g2_mux2_1 _2608_ (.A0(\spi0.spi0.sdo_register[2] ),
    .A1(\spi0.data_tx[19] ),
    .S(net61),
    .X(_0026_));
 sg13g2_mux2_1 _2609_ (.A0(\spi0.spi0.sdo_register[3] ),
    .A1(\spi0.data_tx[20] ),
    .S(net61),
    .X(_0027_));
 sg13g2_mux2_1 _2610_ (.A0(\spi0.spi0.sdo_register[4] ),
    .A1(\spi0.data_tx[21] ),
    .S(net61),
    .X(_0028_));
 sg13g2_mux2_1 _2611_ (.A0(\spi0.spi0.sdo_register[5] ),
    .A1(\spi0.data_tx[22] ),
    .S(_0008_),
    .X(_0029_));
 sg13g2_mux2_1 _2612_ (.A0(\spi0.spi0.sdo_register[6] ),
    .A1(\spi0.data_tx[23] ),
    .S(net61),
    .X(_0030_));
 sg13g2_buf_1 _2613_ (.A(_1927_),
    .X(_1928_));
 sg13g2_mux2_1 _2614_ (.A0(\spi0.spi0.sdo_register[7] ),
    .A1(\spi0.data_tx[8] ),
    .S(net60),
    .X(_0031_));
 sg13g2_mux2_1 _2615_ (.A0(\spi0.spi0.sdo_register[8] ),
    .A1(\spi0.data_tx[9] ),
    .S(net60),
    .X(_0032_));
 sg13g2_mux2_1 _2616_ (.A0(\spi0.spi0.sdo_register[9] ),
    .A1(\spi0.data_tx[10] ),
    .S(net60),
    .X(_0010_));
 sg13g2_mux2_1 _2617_ (.A0(\spi0.spi0.sdo_register[10] ),
    .A1(\spi0.data_tx[11] ),
    .S(net60),
    .X(_0011_));
 sg13g2_mux2_1 _2618_ (.A0(\spi0.spi0.sdo_register[11] ),
    .A1(\spi0.data_tx[12] ),
    .S(net60),
    .X(_0012_));
 sg13g2_mux2_1 _2619_ (.A0(\spi0.spi0.sdo_register[12] ),
    .A1(\spi0.data_tx[13] ),
    .S(_1928_),
    .X(_0013_));
 sg13g2_mux2_1 _2620_ (.A0(\spi0.spi0.sdo_register[13] ),
    .A1(\spi0.data_tx[14] ),
    .S(net60),
    .X(_0014_));
 sg13g2_mux2_1 _2621_ (.A0(\spi0.spi0.sdo_register[14] ),
    .A1(\spi0.data_tx[15] ),
    .S(_1928_),
    .X(_0015_));
 sg13g2_mux2_1 _2622_ (.A0(\spi0.spi0.sdo_register[15] ),
    .A1(\spi0.data_tx[0] ),
    .S(net60),
    .X(_0016_));
 sg13g2_mux2_1 _2623_ (.A0(\spi0.spi0.sdo_register[16] ),
    .A1(\spi0.data_tx[1] ),
    .S(net60),
    .X(_0017_));
 sg13g2_mux2_1 _2624_ (.A0(\spi0.spi0.sdo_register[17] ),
    .A1(\spi0.data_tx[2] ),
    .S(_1927_),
    .X(_0018_));
 sg13g2_mux2_1 _2625_ (.A0(\spi0.spi0.sdo_register[18] ),
    .A1(\spi0.data_tx[3] ),
    .S(_1927_),
    .X(_0019_));
 sg13g2_mux2_1 _2626_ (.A0(\spi0.spi0.sdo_register[19] ),
    .A1(\spi0.data_tx[4] ),
    .S(_1927_),
    .X(_0021_));
 sg13g2_mux2_1 _2627_ (.A0(\spi0.spi0.sdo_register[20] ),
    .A1(\spi0.data_tx[5] ),
    .S(_1927_),
    .X(_0022_));
 sg13g2_mux2_1 _2628_ (.A0(\spi0.spi0.sdo_register[21] ),
    .A1(\spi0.data_tx[6] ),
    .S(_1927_),
    .X(_0023_));
 sg13g2_mux2_1 _2629_ (.A0(\spi0.spi0.sdo_register[22] ),
    .A1(\spi0.data_tx[7] ),
    .S(_1927_),
    .X(_0024_));
 sg13g2_inv_1 _2630_ (.Y(_0002_),
    .A(_1919_));
 sg13g2_xor2_1 _2631_ (.B(_1919_),
    .A(_1922_),
    .X(_0003_));
 sg13g2_nand2_1 _2632_ (.Y(_1929_),
    .A(_1922_),
    .B(_1919_));
 sg13g2_xnor2_1 _2633_ (.Y(_0004_),
    .A(_1920_),
    .B(_1929_));
 sg13g2_nand3_1 _2634_ (.B(_1919_),
    .C(_1920_),
    .A(_1922_),
    .Y(_1930_));
 sg13g2_xor2_1 _2635_ (.B(_1930_),
    .A(_1923_),
    .X(_1931_));
 sg13g2_nor2_1 _2636_ (.A(_0008_),
    .B(_1931_),
    .Y(_0005_));
 sg13g2_nor2_1 _2637_ (.A(_1924_),
    .B(_1930_),
    .Y(_1932_));
 sg13g2_nand3_1 _2638_ (.B(_1923_),
    .C(_1920_),
    .A(_1919_),
    .Y(_1933_));
 sg13g2_nor2b_1 _2639_ (.A(\spi0.spi0.counter[4] ),
    .B_N(_1933_),
    .Y(_1934_));
 sg13g2_nand2_1 _2640_ (.Y(_1935_),
    .A(_1923_),
    .B(_1921_));
 sg13g2_a21oi_1 _2641_ (.A1(\spi0.spi0.counter[4] ),
    .A2(_1935_),
    .Y(_1936_),
    .B1(_1922_));
 sg13g2_nor3_1 _2642_ (.A(_1932_),
    .B(_1934_),
    .C(_1936_),
    .Y(_0006_));
 sg13g2_xor2_1 _2643_ (.B(_1932_),
    .A(\spi0.spi0.counter[5] ),
    .X(_0007_));
 sg13g2_nor2_2 _2644_ (.A(_1908_),
    .B(net62),
    .Y(_1937_));
 sg13g2_buf_1 _2645_ (.A(\gray_sobel0.sobel0.counter_sobel[1] ),
    .X(_1938_));
 sg13g2_buf_2 _2646_ (.A(\gray_sobel0.sobel0.counter_sobel[3] ),
    .X(_1939_));
 sg13g2_buf_2 _2647_ (.A(\gray_sobel0.sobel0.counter_sobel[2] ),
    .X(_1940_));
 sg13g2_nor2_1 _2648_ (.A(\gray_sobel0.sobel0.counter_sobel[0] ),
    .B(_1940_),
    .Y(_1941_));
 sg13g2_nand3b_1 _2649_ (.B(_1939_),
    .C(_1941_),
    .Y(_1942_),
    .A_N(_1938_));
 sg13g2_a21oi_1 _2650_ (.A1(net62),
    .A2(_1942_),
    .Y(_1943_),
    .B1(_1908_));
 sg13g2_nand3b_1 _2651_ (.B(_1941_),
    .C(_1938_),
    .Y(_1944_),
    .A_N(_1939_));
 sg13g2_buf_1 _2652_ (.A(ui_in[3]),
    .X(_1945_));
 sg13g2_mux2_1 _2653_ (.A0(\gray_sobel0.gray_scale0.px_rdy_o ),
    .A1(\gray_sobel0.gray_scale0.px_rdy_i ),
    .S(_1945_),
    .X(_1946_));
 sg13g2_nor2b_1 _2654_ (.A(net5),
    .B_N(_1946_),
    .Y(_1947_));
 sg13g2_buf_1 _2655_ (.A(_1947_),
    .X(_1948_));
 sg13g2_o21ai_1 _2656_ (.B1(_1948_),
    .Y(_1949_),
    .A1(net62),
    .A2(_1944_));
 sg13g2_nor2_1 _2657_ (.A(_1943_),
    .B(_1949_),
    .Y(_1950_));
 sg13g2_nor2_2 _2658_ (.A(_1937_),
    .B(_1948_),
    .Y(_1951_));
 sg13g2_or2_1 _2659_ (.X(_1952_),
    .B(_1951_),
    .A(_1950_));
 sg13g2_buf_1 _2660_ (.A(_1952_),
    .X(_1953_));
 sg13g2_or2_1 _2661_ (.X(_1954_),
    .B(_1953_),
    .A(_1937_));
 sg13g2_buf_1 _2662_ (.A(_1954_),
    .X(_1955_));
 sg13g2_inv_1 _2663_ (.Y(_1956_),
    .A(_1955_));
 sg13g2_buf_1 _2664_ (.A(_1956_),
    .X(_1957_));
 sg13g2_buf_1 _2665_ (.A(net24),
    .X(_0001_));
 sg13g2_buf_1 _2666_ (.A(\input_data[18] ),
    .X(_1958_));
 sg13g2_buf_2 _2667_ (.A(\input_data[21] ),
    .X(_1959_));
 sg13g2_xnor2_1 _2668_ (.Y(_1960_),
    .A(_1958_),
    .B(_1959_));
 sg13g2_xor2_1 _2669_ (.B(_1865_),
    .A(_1846_),
    .X(_1961_));
 sg13g2_nand2_1 _2670_ (.Y(_1962_),
    .A(net93),
    .B(_1961_));
 sg13g2_o21ai_1 _2671_ (.B1(_1962_),
    .Y(_1963_),
    .A1(net93),
    .A2(_1960_));
 sg13g2_buf_1 _2672_ (.A(_1963_),
    .X(_1964_));
 sg13g2_xor2_1 _2673_ (.B(net117),
    .A(_1828_),
    .X(_1965_));
 sg13g2_buf_2 _2674_ (.A(\input_data[4] ),
    .X(_1966_));
 sg13g2_buf_1 _2675_ (.A(\input_data[5] ),
    .X(_1967_));
 sg13g2_xnor2_1 _2676_ (.Y(_1968_),
    .A(_1966_),
    .B(net115));
 sg13g2_nor2_1 _2677_ (.A(net93),
    .B(_1968_),
    .Y(_1969_));
 sg13g2_a21oi_1 _2678_ (.A1(net93),
    .A2(_1965_),
    .Y(_1970_),
    .B1(_1969_));
 sg13g2_xnor2_1 _2679_ (.Y(_1971_),
    .A(_1964_),
    .B(_1970_));
 sg13g2_buf_1 _2680_ (.A(_1917_),
    .X(_1972_));
 sg13g2_buf_1 _2681_ (.A(net59),
    .X(_1973_));
 sg13g2_xor2_1 _2682_ (.B(net118),
    .A(_1831_),
    .X(_1974_));
 sg13g2_buf_2 _2683_ (.A(\input_data[9] ),
    .X(_1975_));
 sg13g2_buf_1 _2684_ (.A(\input_data[12] ),
    .X(_1976_));
 sg13g2_xnor2_1 _2685_ (.Y(_1977_),
    .A(_1975_),
    .B(net114));
 sg13g2_nor2_1 _2686_ (.A(net59),
    .B(_1977_),
    .Y(_1978_));
 sg13g2_a21oi_1 _2687_ (.A1(net55),
    .A2(_1974_),
    .Y(_1979_),
    .B1(_1978_));
 sg13g2_xnor2_1 _2688_ (.Y(_0033_),
    .A(_1971_),
    .B(_1979_));
 sg13g2_buf_1 _2689_ (.A(\input_data[14] ),
    .X(_1980_));
 sg13g2_mux2_1 _2690_ (.A0(_1980_),
    .A1(\lfsr0.lfsr_out[14] ),
    .S(_1915_),
    .X(_1981_));
 sg13g2_buf_2 _2691_ (.A(_1981_),
    .X(_1982_));
 sg13g2_and2_1 _2692_ (.A(_1846_),
    .B(_1865_),
    .X(_1983_));
 sg13g2_nor2b_1 _2693_ (.A(_1912_),
    .B_N(_1958_),
    .Y(_1984_));
 sg13g2_a22oi_1 _2694_ (.Y(_1985_),
    .B1(_1984_),
    .B2(_1959_),
    .A2(_1983_),
    .A1(_1912_));
 sg13g2_buf_1 _2695_ (.A(\input_data[22] ),
    .X(_1986_));
 sg13g2_mux2_1 _2696_ (.A0(_1986_),
    .A1(\lfsr0.lfsr_out[22] ),
    .S(_1912_),
    .X(_1987_));
 sg13g2_buf_1 _2697_ (.A(_1987_),
    .X(_1988_));
 sg13g2_buf_1 _2698_ (.A(_1988_),
    .X(_1989_));
 sg13g2_buf_1 _2699_ (.A(\input_data[19] ),
    .X(_1990_));
 sg13g2_mux2_1 _2700_ (.A0(_1990_),
    .A1(\lfsr0.lfsr_out[19] ),
    .S(_1912_),
    .X(_1991_));
 sg13g2_xor2_1 _2701_ (.B(_1991_),
    .A(_1989_),
    .X(_1992_));
 sg13g2_xnor2_1 _2702_ (.Y(_1993_),
    .A(_1985_),
    .B(_1992_));
 sg13g2_a21oi_1 _2703_ (.A1(net119),
    .A2(_1993_),
    .Y(_1994_),
    .B1(net117));
 sg13g2_nor2_1 _2704_ (.A(net119),
    .B(_1993_),
    .Y(_1995_));
 sg13g2_nor2_1 _2705_ (.A(_1994_),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_buf_1 _2706_ (.A(\input_data[6] ),
    .X(_1997_));
 sg13g2_a21oi_1 _2707_ (.A1(net113),
    .A2(_1993_),
    .Y(_1998_),
    .B1(net115));
 sg13g2_nor2_1 _2708_ (.A(net113),
    .B(_1993_),
    .Y(_1999_));
 sg13g2_nor3_1 _2709_ (.A(net78),
    .B(_1998_),
    .C(_1999_),
    .Y(_2000_));
 sg13g2_a21oi_1 _2710_ (.A1(net71),
    .A2(_1996_),
    .Y(_2001_),
    .B1(_2000_));
 sg13g2_nor2_1 _2711_ (.A(_1988_),
    .B(_1991_),
    .Y(_2002_));
 sg13g2_nor2_1 _2712_ (.A(_1985_),
    .B(_2002_),
    .Y(_2003_));
 sg13g2_a21oi_1 _2713_ (.A1(_1989_),
    .A2(_1991_),
    .Y(_2004_),
    .B1(_2003_));
 sg13g2_buf_1 _2714_ (.A(\input_data[23] ),
    .X(_2005_));
 sg13g2_mux2_1 _2715_ (.A0(_2005_),
    .A1(\lfsr0.lfsr_out[23] ),
    .S(_1912_),
    .X(_2006_));
 sg13g2_buf_2 _2716_ (.A(_2006_),
    .X(_2007_));
 sg13g2_buf_1 _2717_ (.A(\input_data[20] ),
    .X(_2008_));
 sg13g2_mux2_1 _2718_ (.A0(_2008_),
    .A1(\lfsr0.lfsr_out[20] ),
    .S(net93),
    .X(_2009_));
 sg13g2_xor2_1 _2719_ (.B(_2009_),
    .A(_2007_),
    .X(_2010_));
 sg13g2_xnor2_1 _2720_ (.Y(_2011_),
    .A(_2004_),
    .B(_2010_));
 sg13g2_xor2_1 _2721_ (.B(net116),
    .A(net119),
    .X(_2012_));
 sg13g2_buf_1 _2722_ (.A(\input_data[7] ),
    .X(_2013_));
 sg13g2_xnor2_1 _2723_ (.Y(_2014_),
    .A(net113),
    .B(net112));
 sg13g2_nor2_1 _2724_ (.A(net93),
    .B(_2014_),
    .Y(_2015_));
 sg13g2_a21oi_1 _2725_ (.A1(net93),
    .A2(_2012_),
    .Y(_2016_),
    .B1(_2015_));
 sg13g2_xnor2_1 _2726_ (.Y(_2017_),
    .A(_2011_),
    .B(_2016_));
 sg13g2_buf_1 _2727_ (.A(\input_data[11] ),
    .X(_2018_));
 sg13g2_mux2_1 _2728_ (.A0(_2018_),
    .A1(\lfsr0.lfsr_out[11] ),
    .S(net78),
    .X(_2019_));
 sg13g2_xnor2_1 _2729_ (.Y(_2020_),
    .A(_2017_),
    .B(_2019_));
 sg13g2_xnor2_1 _2730_ (.Y(_2021_),
    .A(_2001_),
    .B(_2020_));
 sg13g2_xor2_1 _2731_ (.B(net119),
    .A(net117),
    .X(_2022_));
 sg13g2_xnor2_1 _2732_ (.Y(_2023_),
    .A(net115),
    .B(net113));
 sg13g2_nor2_1 _2733_ (.A(net93),
    .B(_2023_),
    .Y(_2024_));
 sg13g2_a21oi_1 _2734_ (.A1(net78),
    .A2(_2022_),
    .Y(_2025_),
    .B1(_2024_));
 sg13g2_xnor2_1 _2735_ (.Y(_2026_),
    .A(_1993_),
    .B(_2025_));
 sg13g2_buf_1 _2736_ (.A(\input_data[10] ),
    .X(_2027_));
 sg13g2_mux2_1 _2737_ (.A0(_2027_),
    .A1(\lfsr0.lfsr_out[10] ),
    .S(net78),
    .X(_2028_));
 sg13g2_nor2_1 _2738_ (.A(_2026_),
    .B(_2028_),
    .Y(_2029_));
 sg13g2_nand2_1 _2739_ (.Y(_2030_),
    .A(_2026_),
    .B(_2028_));
 sg13g2_a21oi_1 _2740_ (.A1(net117),
    .A2(_1964_),
    .Y(_2031_),
    .B1(_1828_));
 sg13g2_nor2_1 _2741_ (.A(net117),
    .B(_1964_),
    .Y(_2032_));
 sg13g2_nor2_1 _2742_ (.A(_2031_),
    .B(_2032_),
    .Y(_2033_));
 sg13g2_a21oi_1 _2743_ (.A1(net115),
    .A2(_1964_),
    .Y(_2034_),
    .B1(_1966_));
 sg13g2_nor2_1 _2744_ (.A(net115),
    .B(_1964_),
    .Y(_2035_));
 sg13g2_nor3_1 _2745_ (.A(net78),
    .B(_2034_),
    .C(_2035_),
    .Y(_2036_));
 sg13g2_a21oi_1 _2746_ (.A1(net71),
    .A2(_2033_),
    .Y(_2037_),
    .B1(_2036_));
 sg13g2_nand2_1 _2747_ (.Y(_2038_),
    .A(_2030_),
    .B(_2037_));
 sg13g2_nand2b_1 _2748_ (.Y(_2039_),
    .B(_2038_),
    .A_N(_2029_));
 sg13g2_xnor2_1 _2749_ (.Y(_2040_),
    .A(_2021_),
    .B(_2039_));
 sg13g2_xnor2_1 _2750_ (.Y(_2041_),
    .A(_1982_),
    .B(_2040_));
 sg13g2_buf_1 _2751_ (.A(\input_data[13] ),
    .X(_2042_));
 sg13g2_mux2_1 _2752_ (.A0(_2042_),
    .A1(\lfsr0.lfsr_out[13] ),
    .S(_1915_),
    .X(_2043_));
 sg13g2_buf_1 _2753_ (.A(_2043_),
    .X(_2044_));
 sg13g2_a21oi_1 _2754_ (.A1(net118),
    .A2(_1971_),
    .Y(_2045_),
    .B1(_1831_));
 sg13g2_nor2_1 _2755_ (.A(net118),
    .B(_1971_),
    .Y(_2046_));
 sg13g2_nor2_1 _2756_ (.A(_2045_),
    .B(_2046_),
    .Y(_2047_));
 sg13g2_a21oi_1 _2757_ (.A1(net114),
    .A2(_1971_),
    .Y(_2048_),
    .B1(_1975_));
 sg13g2_nor2_1 _2758_ (.A(net114),
    .B(_1971_),
    .Y(_2049_));
 sg13g2_nor3_1 _2759_ (.A(net71),
    .B(_2048_),
    .C(_2049_),
    .Y(_2050_));
 sg13g2_a21oi_1 _2760_ (.A1(net71),
    .A2(_2047_),
    .Y(_2051_),
    .B1(_2050_));
 sg13g2_inv_1 _2761_ (.Y(_2052_),
    .A(_2051_));
 sg13g2_nor2_1 _2762_ (.A(net66),
    .B(_2052_),
    .Y(_2053_));
 sg13g2_nand2b_1 _2763_ (.Y(_2054_),
    .B(_2030_),
    .A_N(_2029_));
 sg13g2_xnor2_1 _2764_ (.Y(_2055_),
    .A(_2037_),
    .B(_2054_));
 sg13g2_nand2_1 _2765_ (.Y(_2056_),
    .A(net66),
    .B(_2052_));
 sg13g2_o21ai_1 _2766_ (.B1(_2056_),
    .Y(_2057_),
    .A1(_2053_),
    .A2(_2055_));
 sg13g2_xor2_1 _2767_ (.B(_2057_),
    .A(_2041_),
    .X(_0035_));
 sg13g2_a21oi_1 _2768_ (.A1(net116),
    .A2(_2011_),
    .Y(_2058_),
    .B1(net119));
 sg13g2_nor2_1 _2769_ (.A(net116),
    .B(_2011_),
    .Y(_2059_));
 sg13g2_nor2_1 _2770_ (.A(_2058_),
    .B(_2059_),
    .Y(_2060_));
 sg13g2_a21oi_1 _2771_ (.A1(net112),
    .A2(_2011_),
    .Y(_2061_),
    .B1(net113));
 sg13g2_nor2_1 _2772_ (.A(net112),
    .B(_2011_),
    .Y(_2062_));
 sg13g2_nor3_1 _2773_ (.A(net71),
    .B(_2061_),
    .C(_2062_),
    .Y(_2063_));
 sg13g2_a21oi_1 _2774_ (.A1(net71),
    .A2(_2060_),
    .Y(_2064_),
    .B1(_2063_));
 sg13g2_nor2_1 _2775_ (.A(_2007_),
    .B(_2009_),
    .Y(_2065_));
 sg13g2_nand2_1 _2776_ (.Y(_2066_),
    .A(_2007_),
    .B(_2009_));
 sg13g2_o21ai_1 _2777_ (.B1(_2066_),
    .Y(_2067_),
    .A1(_2004_),
    .A2(_2065_));
 sg13g2_mux2_1 _2778_ (.A0(_1959_),
    .A1(_1865_),
    .S(_1913_),
    .X(_2068_));
 sg13g2_buf_1 _2779_ (.A(_2068_),
    .X(_2069_));
 sg13g2_xor2_1 _2780_ (.B(_2069_),
    .A(_2067_),
    .X(_2070_));
 sg13g2_xor2_1 _2781_ (.B(net118),
    .A(net116),
    .X(_2071_));
 sg13g2_xnor2_1 _2782_ (.Y(_2072_),
    .A(net112),
    .B(net114));
 sg13g2_nor2_1 _2783_ (.A(net78),
    .B(_2072_),
    .Y(_2073_));
 sg13g2_a21oi_1 _2784_ (.A1(net78),
    .A2(_2071_),
    .Y(_2074_),
    .B1(_2073_));
 sg13g2_xnor2_1 _2785_ (.Y(_2075_),
    .A(_2070_),
    .B(_2074_));
 sg13g2_buf_1 _2786_ (.A(\input_data[15] ),
    .X(_2076_));
 sg13g2_mux2_1 _2787_ (.A0(_2076_),
    .A1(\lfsr0.lfsr_out[15] ),
    .S(_1914_),
    .X(_2077_));
 sg13g2_buf_1 _2788_ (.A(_2077_),
    .X(_2078_));
 sg13g2_xnor2_1 _2789_ (.Y(_2079_),
    .A(_2075_),
    .B(_2078_));
 sg13g2_xnor2_1 _2790_ (.Y(_2080_),
    .A(_2064_),
    .B(_2079_));
 sg13g2_nor2_1 _2791_ (.A(_2017_),
    .B(_2019_),
    .Y(_2081_));
 sg13g2_nand2_1 _2792_ (.Y(_2082_),
    .A(_2017_),
    .B(_2019_));
 sg13g2_o21ai_1 _2793_ (.B1(_2082_),
    .Y(_2083_),
    .A1(_2001_),
    .A2(_2081_));
 sg13g2_xnor2_1 _2794_ (.Y(_2084_),
    .A(_2080_),
    .B(_2083_));
 sg13g2_nand2_1 _2795_ (.Y(_2085_),
    .A(_2041_),
    .B(_2057_));
 sg13g2_nor2_1 _2796_ (.A(_2021_),
    .B(_2039_),
    .Y(_2086_));
 sg13g2_nand2_1 _2797_ (.Y(_2087_),
    .A(_2021_),
    .B(_2039_));
 sg13g2_o21ai_1 _2798_ (.B1(_2087_),
    .Y(_2088_),
    .A1(_1982_),
    .A2(_2086_));
 sg13g2_xnor2_1 _2799_ (.Y(_2089_),
    .A(_2085_),
    .B(_2088_));
 sg13g2_xnor2_1 _2800_ (.Y(_0036_),
    .A(_2084_),
    .B(_2089_));
 sg13g2_nand2b_1 _2801_ (.Y(_2090_),
    .B(_2088_),
    .A_N(_2084_));
 sg13g2_nand2b_1 _2802_ (.Y(_2091_),
    .B(_2084_),
    .A_N(_2088_));
 sg13g2_nand2_1 _2803_ (.Y(_2092_),
    .A(_2085_),
    .B(_2091_));
 sg13g2_nand2_1 _2804_ (.Y(_2093_),
    .A(_2090_),
    .B(_2092_));
 sg13g2_nor2b_1 _2805_ (.A(_2080_),
    .B_N(_2083_),
    .Y(_2094_));
 sg13g2_nor2_1 _2806_ (.A(_2075_),
    .B(_2078_),
    .Y(_2095_));
 sg13g2_nand2_1 _2807_ (.Y(_2096_),
    .A(_2075_),
    .B(_2078_));
 sg13g2_o21ai_1 _2808_ (.B1(_2096_),
    .Y(_2097_),
    .A1(_2064_),
    .A2(_2095_));
 sg13g2_a21oi_1 _2809_ (.A1(net118),
    .A2(_2070_),
    .Y(_2098_),
    .B1(net116));
 sg13g2_nor2_1 _2810_ (.A(net118),
    .B(_2070_),
    .Y(_2099_));
 sg13g2_nor2_1 _2811_ (.A(_2098_),
    .B(_2099_),
    .Y(_2100_));
 sg13g2_a21oi_1 _2812_ (.A1(net114),
    .A2(_2070_),
    .Y(_2101_),
    .B1(net112));
 sg13g2_nor2_1 _2813_ (.A(net114),
    .B(_2070_),
    .Y(_2102_));
 sg13g2_nor3_1 _2814_ (.A(net71),
    .B(_2101_),
    .C(_2102_),
    .Y(_2103_));
 sg13g2_a21oi_1 _2815_ (.A1(net69),
    .A2(_2100_),
    .Y(_2104_),
    .B1(_2103_));
 sg13g2_buf_2 _2816_ (.A(_2104_),
    .X(_2105_));
 sg13g2_nand2_2 _2817_ (.Y(_2106_),
    .A(_2067_),
    .B(_2069_));
 sg13g2_xnor2_1 _2818_ (.Y(_2107_),
    .A(net70),
    .B(_2106_));
 sg13g2_xor2_1 _2819_ (.B(_2107_),
    .A(net66),
    .X(_2108_));
 sg13g2_xnor2_1 _2820_ (.Y(_2109_),
    .A(_2105_),
    .B(_2108_));
 sg13g2_xnor2_1 _2821_ (.Y(_2110_),
    .A(_2097_),
    .B(_2109_));
 sg13g2_xnor2_1 _2822_ (.Y(_2111_),
    .A(_2094_),
    .B(_2110_));
 sg13g2_xnor2_1 _2823_ (.Y(_0037_),
    .A(_2093_),
    .B(_2111_));
 sg13g2_nor2_1 _2824_ (.A(_2093_),
    .B(_2110_),
    .Y(_2112_));
 sg13g2_nand2_1 _2825_ (.Y(_2113_),
    .A(_2093_),
    .B(_2110_));
 sg13g2_o21ai_1 _2826_ (.B1(_2113_),
    .Y(_2114_),
    .A1(_2094_),
    .A2(_2112_));
 sg13g2_nand2_1 _2827_ (.Y(_2115_),
    .A(_2097_),
    .B(_2109_));
 sg13g2_xor2_1 _2828_ (.B(_2007_),
    .A(_1982_),
    .X(_2116_));
 sg13g2_nor2_1 _2829_ (.A(_2106_),
    .B(_2105_),
    .Y(_2117_));
 sg13g2_nor2_1 _2830_ (.A(net66),
    .B(_2117_),
    .Y(_2118_));
 sg13g2_a21oi_1 _2831_ (.A1(_2106_),
    .A2(_2105_),
    .Y(_2119_),
    .B1(_2118_));
 sg13g2_nand4_1 _2832_ (.B(net66),
    .C(_2067_),
    .A(net70),
    .Y(_2120_),
    .D(_2069_));
 sg13g2_nand2b_1 _2833_ (.Y(_2121_),
    .B(_2106_),
    .A_N(net66));
 sg13g2_mux2_1 _2834_ (.A0(_2120_),
    .A1(_2121_),
    .S(_2105_),
    .X(_2122_));
 sg13g2_o21ai_1 _2835_ (.B1(_2122_),
    .Y(_2123_),
    .A1(net70),
    .A2(_2119_));
 sg13g2_xor2_1 _2836_ (.B(_2123_),
    .A(_2116_),
    .X(_2124_));
 sg13g2_xor2_1 _2837_ (.B(_2124_),
    .A(_2115_),
    .X(_2125_));
 sg13g2_xnor2_1 _2838_ (.Y(_0038_),
    .A(_2114_),
    .B(_2125_));
 sg13g2_nand2_1 _2839_ (.Y(_2126_),
    .A(_2124_),
    .B(_2114_));
 sg13g2_o21ai_1 _2840_ (.B1(_2115_),
    .Y(_2127_),
    .A1(_2124_),
    .A2(_2114_));
 sg13g2_nand2_1 _2841_ (.Y(_2128_),
    .A(_2126_),
    .B(_2127_));
 sg13g2_nand2b_1 _2842_ (.Y(_2129_),
    .B(net66),
    .A_N(net70));
 sg13g2_inv_1 _2843_ (.Y(_2130_),
    .A(_2105_));
 sg13g2_o21ai_1 _2844_ (.B1(_2107_),
    .Y(_2131_),
    .A1(_2044_),
    .A2(_2130_));
 sg13g2_o21ai_1 _2845_ (.B1(_2131_),
    .Y(_2132_),
    .A1(_2105_),
    .A2(_2129_));
 sg13g2_nor2_1 _2846_ (.A(_2116_),
    .B(_2120_),
    .Y(_2133_));
 sg13g2_a22oi_1 _2847_ (.Y(_2134_),
    .B1(_2133_),
    .B2(_2130_),
    .A2(_2132_),
    .A1(_2116_));
 sg13g2_nor2b_1 _2848_ (.A(_2106_),
    .B_N(net70),
    .Y(_2135_));
 sg13g2_a21o_1 _2849_ (.A2(_2135_),
    .A1(_2007_),
    .B1(_1982_),
    .X(_2136_));
 sg13g2_o21ai_1 _2850_ (.B1(_2136_),
    .Y(_2137_),
    .A1(_2007_),
    .A2(_2135_));
 sg13g2_xnor2_1 _2851_ (.Y(_2138_),
    .A(_2078_),
    .B(_2137_));
 sg13g2_xnor2_1 _2852_ (.Y(_2139_),
    .A(_2134_),
    .B(_2138_));
 sg13g2_xnor2_1 _2853_ (.Y(_0039_),
    .A(_2128_),
    .B(_2139_));
 sg13g2_nor2b_1 _2854_ (.A(_2106_),
    .B_N(_2044_),
    .Y(_2140_));
 sg13g2_nand2b_1 _2855_ (.Y(_2141_),
    .B(_2121_),
    .A_N(_2140_));
 sg13g2_nand2b_1 _2856_ (.Y(_2142_),
    .B(net70),
    .A_N(_2121_));
 sg13g2_o21ai_1 _2857_ (.B1(_2142_),
    .Y(_2143_),
    .A1(net70),
    .A2(_2141_));
 sg13g2_a21oi_1 _2858_ (.A1(_2116_),
    .A2(_2143_),
    .Y(_2144_),
    .B1(_2133_));
 sg13g2_or2_1 _2859_ (.X(_2145_),
    .B(_2144_),
    .A(_2105_));
 sg13g2_a221oi_1 _2860_ (.B2(net70),
    .C1(_2140_),
    .B1(_2121_),
    .A1(_1982_),
    .Y(_2146_),
    .A2(_2007_));
 sg13g2_inv_1 _2861_ (.Y(_2147_),
    .A(_2146_));
 sg13g2_o21ai_1 _2862_ (.B1(_2147_),
    .Y(_2148_),
    .A1(_1982_),
    .A2(_2007_));
 sg13g2_nand2_1 _2863_ (.Y(_2149_),
    .A(_2145_),
    .B(_2148_));
 sg13g2_o21ai_1 _2864_ (.B1(_2128_),
    .Y(_2150_),
    .A1(_2145_),
    .A2(_2148_));
 sg13g2_a21oi_1 _2865_ (.A1(_2149_),
    .A2(_2150_),
    .Y(_2151_),
    .B1(_2078_));
 sg13g2_nand2b_1 _2866_ (.Y(_2152_),
    .B(_2128_),
    .A_N(_2149_));
 sg13g2_nor2b_1 _2867_ (.A(_2151_),
    .B_N(_2152_),
    .Y(_0040_));
 sg13g2_xnor2_1 _2868_ (.Y(_2153_),
    .A(_2051_),
    .B(_2055_));
 sg13g2_xnor2_1 _2869_ (.Y(_0034_),
    .A(net66),
    .B(_2153_));
 sg13g2_inv_1 _2870_ (.Y(_0042_),
    .A(net185));
 sg13g2_inv_1 _2871_ (.Y(_0041_),
    .A(net3));
 sg13g2_buf_1 _2872_ (.A(_1955_),
    .X(_2154_));
 sg13g2_buf_1 _2873_ (.A(_1953_),
    .X(_2155_));
 sg13g2_nand2_1 _2874_ (.Y(_2156_),
    .A(_1900_),
    .B(net33));
 sg13g2_o21ai_1 _2875_ (.B1(_2156_),
    .Y(_0043_),
    .A1(_1900_),
    .A2(net30));
 sg13g2_buf_1 _2876_ (.A(net24),
    .X(_2157_));
 sg13g2_inv_1 _2877_ (.Y(_2158_),
    .A(\gray_sobel0.sobel0.counter_pixels[3] ));
 sg13g2_nand3_1 _2878_ (.B(_1899_),
    .C(\gray_sobel0.sobel0.counter_pixels[2] ),
    .A(_1900_),
    .Y(_2159_));
 sg13g2_nor2_2 _2879_ (.A(_2158_),
    .B(_2159_),
    .Y(_2160_));
 sg13g2_and3_1 _2880_ (.X(_2161_),
    .A(\gray_sobel0.sobel0.counter_pixels[5] ),
    .B(_1885_),
    .C(_2160_));
 sg13g2_buf_1 _2881_ (.A(_2161_),
    .X(_2162_));
 sg13g2_and2_1 _2882_ (.A(\gray_sobel0.sobel0.counter_pixels[6] ),
    .B(_2162_),
    .X(_2163_));
 sg13g2_buf_1 _2883_ (.A(_2163_),
    .X(_2164_));
 sg13g2_and2_1 _2884_ (.A(_1886_),
    .B(_2164_),
    .X(_2165_));
 sg13g2_buf_1 _2885_ (.A(_2165_),
    .X(_2166_));
 sg13g2_and3_1 _2886_ (.X(_2167_),
    .A(_1897_),
    .B(_1892_),
    .C(_2166_));
 sg13g2_buf_1 _2887_ (.A(_2167_),
    .X(_2168_));
 sg13g2_nand2_1 _2888_ (.Y(_2169_),
    .A(net21),
    .B(_2168_));
 sg13g2_nor2_1 _2889_ (.A(net30),
    .B(_2168_),
    .Y(_2170_));
 sg13g2_o21ai_1 _2890_ (.B1(_1894_),
    .Y(_2171_),
    .A1(net33),
    .A2(_2170_));
 sg13g2_o21ai_1 _2891_ (.B1(_2171_),
    .Y(_0044_),
    .A1(_1894_),
    .A2(_2169_));
 sg13g2_and2_1 _2892_ (.A(_1894_),
    .B(_2168_),
    .X(_2172_));
 sg13g2_buf_1 _2893_ (.A(_2172_),
    .X(_2173_));
 sg13g2_nand2_1 _2894_ (.Y(_2174_),
    .A(_2157_),
    .B(_2173_));
 sg13g2_nor2_1 _2895_ (.A(net30),
    .B(_2173_),
    .Y(_2175_));
 sg13g2_o21ai_1 _2896_ (.B1(_1893_),
    .Y(_2176_),
    .A1(net33),
    .A2(_2175_));
 sg13g2_o21ai_1 _2897_ (.B1(_2176_),
    .Y(_0045_),
    .A1(_1893_),
    .A2(_2174_));
 sg13g2_buf_1 _2898_ (.A(_1956_),
    .X(_2177_));
 sg13g2_nand3_1 _2899_ (.B(net23),
    .C(_2173_),
    .A(_1893_),
    .Y(_2178_));
 sg13g2_buf_1 _2900_ (.A(_1955_),
    .X(_2179_));
 sg13g2_a21oi_1 _2901_ (.A1(_1893_),
    .A2(_2173_),
    .Y(_2180_),
    .B1(net29));
 sg13g2_o21ai_1 _2902_ (.B1(_1895_),
    .Y(_2181_),
    .A1(_2155_),
    .A2(_2180_));
 sg13g2_o21ai_1 _2903_ (.B1(_2181_),
    .Y(_0046_),
    .A1(_1895_),
    .A2(_2178_));
 sg13g2_and4_1 _2904_ (.A(_1886_),
    .B(_1897_),
    .C(_1892_),
    .D(_1894_),
    .X(_2182_));
 sg13g2_and4_1 _2905_ (.A(_1893_),
    .B(_1895_),
    .C(_2164_),
    .D(_2182_),
    .X(_2183_));
 sg13g2_buf_1 _2906_ (.A(_2183_),
    .X(_2184_));
 sg13g2_nor2_1 _2907_ (.A(_2154_),
    .B(_2184_),
    .Y(_2185_));
 sg13g2_o21ai_1 _2908_ (.B1(_1898_),
    .Y(_0271_),
    .A1(_2155_),
    .A2(_2185_));
 sg13g2_nand3b_1 _2909_ (.B(_2157_),
    .C(_2184_),
    .Y(_0272_),
    .A_N(_1898_));
 sg13g2_nand2_1 _2910_ (.Y(_0047_),
    .A(_0271_),
    .B(_0272_));
 sg13g2_nand2_1 _2911_ (.Y(_0273_),
    .A(_1898_),
    .B(_2184_));
 sg13g2_a21o_1 _2912_ (.A2(_0273_),
    .A1(_1957_),
    .B1(_1953_),
    .X(_0274_));
 sg13g2_nor3_1 _2913_ (.A(_1889_),
    .B(net30),
    .C(_0273_),
    .Y(_0275_));
 sg13g2_a21o_1 _2914_ (.A2(_0274_),
    .A1(_1889_),
    .B1(_0275_),
    .X(_0048_));
 sg13g2_and4_1 _2915_ (.A(_1893_),
    .B(_1898_),
    .C(_1895_),
    .D(_2173_),
    .X(_0276_));
 sg13g2_nand3_1 _2916_ (.B(net23),
    .C(_0276_),
    .A(_1889_),
    .Y(_0277_));
 sg13g2_and3_1 _2917_ (.X(_0278_),
    .A(_1898_),
    .B(_1889_),
    .C(_2184_));
 sg13g2_buf_1 _2918_ (.A(_0278_),
    .X(_0279_));
 sg13g2_nor2_1 _2919_ (.A(net30),
    .B(_0279_),
    .Y(_0280_));
 sg13g2_o21ai_1 _2920_ (.B1(_1888_),
    .Y(_0281_),
    .A1(net33),
    .A2(_0280_));
 sg13g2_o21ai_1 _2921_ (.B1(_0281_),
    .Y(_0049_),
    .A1(_1888_),
    .A2(_0277_));
 sg13g2_nand3_1 _2922_ (.B(net24),
    .C(_0279_),
    .A(_1888_),
    .Y(_0282_));
 sg13g2_a21oi_1 _2923_ (.A1(_1888_),
    .A2(_0279_),
    .Y(_0283_),
    .B1(_2179_));
 sg13g2_o21ai_1 _2924_ (.B1(_1877_),
    .Y(_0284_),
    .A1(net33),
    .A2(_0283_));
 sg13g2_o21ai_1 _2925_ (.B1(_0284_),
    .Y(_0050_),
    .A1(_1877_),
    .A2(_0282_));
 sg13g2_and4_1 _2926_ (.A(_1888_),
    .B(_1889_),
    .C(_1877_),
    .D(_0276_),
    .X(_0285_));
 sg13g2_buf_1 _2927_ (.A(_0285_),
    .X(_0286_));
 sg13g2_nand2_1 _2928_ (.Y(_0287_),
    .A(_2177_),
    .B(_0286_));
 sg13g2_nor2_1 _2929_ (.A(net30),
    .B(_0286_),
    .Y(_0288_));
 sg13g2_o21ai_1 _2930_ (.B1(_1876_),
    .Y(_0289_),
    .A1(net33),
    .A2(_0288_));
 sg13g2_o21ai_1 _2931_ (.B1(_0289_),
    .Y(_0051_),
    .A1(_1876_),
    .A2(_0287_));
 sg13g2_and2_1 _2932_ (.A(_1876_),
    .B(_0286_),
    .X(_0290_));
 sg13g2_nand2_1 _2933_ (.Y(_0291_),
    .A(_2177_),
    .B(_0290_));
 sg13g2_and4_1 _2934_ (.A(_1888_),
    .B(_1876_),
    .C(_1877_),
    .D(_0279_),
    .X(_0292_));
 sg13g2_nor2_1 _2935_ (.A(_2179_),
    .B(_0292_),
    .Y(_0293_));
 sg13g2_o21ai_1 _2936_ (.B1(_1879_),
    .Y(_0294_),
    .A1(net33),
    .A2(_0293_));
 sg13g2_o21ai_1 _2937_ (.B1(_0294_),
    .Y(_0052_),
    .A1(_1879_),
    .A2(_0291_));
 sg13g2_nand3_1 _2938_ (.B(net24),
    .C(_0290_),
    .A(_1879_),
    .Y(_0295_));
 sg13g2_buf_1 _2939_ (.A(_1953_),
    .X(_0296_));
 sg13g2_and2_1 _2940_ (.A(_1879_),
    .B(_0292_),
    .X(_0297_));
 sg13g2_nor2_1 _2941_ (.A(net29),
    .B(_0297_),
    .Y(_0298_));
 sg13g2_o21ai_1 _2942_ (.B1(_1878_),
    .Y(_0299_),
    .A1(net32),
    .A2(_0298_));
 sg13g2_o21ai_1 _2943_ (.B1(_0299_),
    .Y(_0053_),
    .A1(_1878_),
    .A2(_0295_));
 sg13g2_nor2_1 _2944_ (.A(_1900_),
    .B(_1937_),
    .Y(_0300_));
 sg13g2_o21ai_1 _2945_ (.B1(_1899_),
    .Y(_0301_),
    .A1(net32),
    .A2(_0300_));
 sg13g2_o21ai_1 _2946_ (.B1(_0301_),
    .Y(_0054_),
    .A1(_1901_),
    .A2(_2154_));
 sg13g2_and3_1 _2947_ (.X(_0302_),
    .A(_1878_),
    .B(_1879_),
    .C(_0290_));
 sg13g2_buf_1 _2948_ (.A(_0302_),
    .X(_0303_));
 sg13g2_nand2_1 _2949_ (.Y(_0304_),
    .A(net23),
    .B(_0303_));
 sg13g2_nor2_1 _2950_ (.A(net29),
    .B(_0303_),
    .Y(_0305_));
 sg13g2_o21ai_1 _2951_ (.B1(_1882_),
    .Y(_0306_),
    .A1(net32),
    .A2(_0305_));
 sg13g2_o21ai_1 _2952_ (.B1(_0306_),
    .Y(_0055_),
    .A1(_1882_),
    .A2(_0304_));
 sg13g2_and2_1 _2953_ (.A(_1882_),
    .B(_0303_),
    .X(_0307_));
 sg13g2_buf_1 _2954_ (.A(_0307_),
    .X(_0308_));
 sg13g2_nand2_1 _2955_ (.Y(_0309_),
    .A(net23),
    .B(_0308_));
 sg13g2_nor2_1 _2956_ (.A(net29),
    .B(_0308_),
    .Y(_0310_));
 sg13g2_o21ai_1 _2957_ (.B1(_1881_),
    .Y(_0311_),
    .A1(net32),
    .A2(_0310_));
 sg13g2_o21ai_1 _2958_ (.B1(_0311_),
    .Y(_0056_),
    .A1(_1881_),
    .A2(_0309_));
 sg13g2_nand4_1 _2959_ (.B(_1881_),
    .C(_1882_),
    .A(_1878_),
    .Y(_0312_),
    .D(_0297_));
 sg13g2_a21o_1 _2960_ (.A2(_0312_),
    .A1(net24),
    .B1(_1953_),
    .X(_0313_));
 sg13g2_nor3_1 _2961_ (.A(_1883_),
    .B(net30),
    .C(_0312_),
    .Y(_0314_));
 sg13g2_a21o_1 _2962_ (.A2(_0313_),
    .A1(_1883_),
    .B1(_0314_),
    .X(_0057_));
 sg13g2_nand4_1 _2963_ (.B(_1883_),
    .C(net24),
    .A(_1881_),
    .Y(_0315_),
    .D(_0308_));
 sg13g2_inv_1 _2964_ (.Y(_0316_),
    .A(_0312_));
 sg13g2_a21oi_1 _2965_ (.A1(_1883_),
    .A2(_0316_),
    .Y(_0317_),
    .B1(_1955_));
 sg13g2_o21ai_1 _2966_ (.B1(\gray_sobel0.sobel0.counter_pixels[23] ),
    .Y(_0318_),
    .A1(net32),
    .A2(_0317_));
 sg13g2_o21ai_1 _2967_ (.B1(_0318_),
    .Y(_0058_),
    .A1(\gray_sobel0.sobel0.counter_pixels[23] ),
    .A2(_0315_));
 sg13g2_nand3_1 _2968_ (.B(_1899_),
    .C(net24),
    .A(_1900_),
    .Y(_0319_));
 sg13g2_a21oi_1 _2969_ (.A1(_1900_),
    .A2(_1899_),
    .Y(_0320_),
    .B1(_1955_));
 sg13g2_o21ai_1 _2970_ (.B1(\gray_sobel0.sobel0.counter_pixels[2] ),
    .Y(_0321_),
    .A1(_0296_),
    .A2(_0320_));
 sg13g2_o21ai_1 _2971_ (.B1(_0321_),
    .Y(_0059_),
    .A1(\gray_sobel0.sobel0.counter_pixels[2] ),
    .A2(_0319_));
 sg13g2_xnor2_1 _2972_ (.Y(_0322_),
    .A(_2158_),
    .B(_2159_));
 sg13g2_nand2_1 _2973_ (.Y(_0323_),
    .A(\gray_sobel0.sobel0.counter_pixels[3] ),
    .B(net33));
 sg13g2_o21ai_1 _2974_ (.B1(_0323_),
    .Y(_0060_),
    .A1(net30),
    .A2(_0322_));
 sg13g2_nand2_1 _2975_ (.Y(_0324_),
    .A(net23),
    .B(_2160_));
 sg13g2_nor2_1 _2976_ (.A(net29),
    .B(_2160_),
    .Y(_0325_));
 sg13g2_o21ai_1 _2977_ (.B1(_1885_),
    .Y(_0326_),
    .A1(net32),
    .A2(_0325_));
 sg13g2_o21ai_1 _2978_ (.B1(_0326_),
    .Y(_0061_),
    .A1(_1885_),
    .A2(_0324_));
 sg13g2_nand3_1 _2979_ (.B(net24),
    .C(_2160_),
    .A(_1885_),
    .Y(_0327_));
 sg13g2_a21oi_1 _2980_ (.A1(_1885_),
    .A2(_2160_),
    .Y(_0328_),
    .B1(_1955_));
 sg13g2_o21ai_1 _2981_ (.B1(\gray_sobel0.sobel0.counter_pixels[5] ),
    .Y(_0329_),
    .A1(_0296_),
    .A2(_0328_));
 sg13g2_o21ai_1 _2982_ (.B1(_0329_),
    .Y(_0062_),
    .A1(\gray_sobel0.sobel0.counter_pixels[5] ),
    .A2(_0327_));
 sg13g2_nand2_1 _2983_ (.Y(_0330_),
    .A(net23),
    .B(_2162_));
 sg13g2_nor2_1 _2984_ (.A(net29),
    .B(_2162_),
    .Y(_0331_));
 sg13g2_o21ai_1 _2985_ (.B1(\gray_sobel0.sobel0.counter_pixels[6] ),
    .Y(_0332_),
    .A1(net32),
    .A2(_0331_));
 sg13g2_o21ai_1 _2986_ (.B1(_0332_),
    .Y(_0063_),
    .A1(\gray_sobel0.sobel0.counter_pixels[6] ),
    .A2(_0330_));
 sg13g2_nand2_1 _2987_ (.Y(_0333_),
    .A(net23),
    .B(_2164_));
 sg13g2_nor2_1 _2988_ (.A(net29),
    .B(_2164_),
    .Y(_0334_));
 sg13g2_o21ai_1 _2989_ (.B1(_1886_),
    .Y(_0335_),
    .A1(net32),
    .A2(_0334_));
 sg13g2_o21ai_1 _2990_ (.B1(_0335_),
    .Y(_0064_),
    .A1(_1886_),
    .A2(_0333_));
 sg13g2_nand2_1 _2991_ (.Y(_0336_),
    .A(net23),
    .B(_2166_));
 sg13g2_nor2_1 _2992_ (.A(net29),
    .B(_2166_),
    .Y(_0337_));
 sg13g2_o21ai_1 _2993_ (.B1(_1892_),
    .Y(_0338_),
    .A1(_1953_),
    .A2(_0337_));
 sg13g2_o21ai_1 _2994_ (.B1(_0338_),
    .Y(_0065_),
    .A1(_1892_),
    .A2(_0336_));
 sg13g2_nand3_1 _2995_ (.B(_1957_),
    .C(_2166_),
    .A(_1892_),
    .Y(_0339_));
 sg13g2_a21oi_1 _2996_ (.A1(_1892_),
    .A2(_2166_),
    .Y(_0340_),
    .B1(_1955_));
 sg13g2_o21ai_1 _2997_ (.B1(_1897_),
    .Y(_0341_),
    .A1(_1953_),
    .A2(_0340_));
 sg13g2_o21ai_1 _2998_ (.B1(_0341_),
    .Y(_0066_),
    .A1(_1897_),
    .A2(_0339_));
 sg13g2_buf_1 _2999_ (.A(\gray_sobel0.sobel0.counter_sobel[0] ),
    .X(_0342_));
 sg13g2_inv_1 _3000_ (.Y(_0343_),
    .A(_1950_));
 sg13g2_nand2_1 _3001_ (.Y(_0344_),
    .A(net111),
    .B(_1951_));
 sg13g2_o21ai_1 _3002_ (.B1(_0344_),
    .Y(_0067_),
    .A1(net111),
    .A2(_0343_));
 sg13g2_buf_1 _3003_ (.A(_1938_),
    .X(_0345_));
 sg13g2_nor2_1 _3004_ (.A(_1940_),
    .B(_1939_),
    .Y(_0346_));
 sg13g2_nor2b_1 _3005_ (.A(net62),
    .B_N(_0346_),
    .Y(_0347_));
 sg13g2_o21ai_1 _3006_ (.B1(_1948_),
    .Y(_0348_),
    .A1(net111),
    .A2(_0347_));
 sg13g2_nand2_1 _3007_ (.Y(_0349_),
    .A(net111),
    .B(_1948_));
 sg13g2_nor2_1 _3008_ (.A(net92),
    .B(_0349_),
    .Y(_0350_));
 sg13g2_a21oi_1 _3009_ (.A1(net92),
    .A2(_0348_),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_nor2_1 _3010_ (.A(_1937_),
    .B(_0351_),
    .Y(_0068_));
 sg13g2_nand3_1 _3011_ (.B(net111),
    .C(_1950_),
    .A(_0345_),
    .Y(_0352_));
 sg13g2_a21oi_1 _3012_ (.A1(_0345_),
    .A2(_0342_),
    .Y(_0353_),
    .B1(_0343_));
 sg13g2_o21ai_1 _3013_ (.B1(_1940_),
    .Y(_0354_),
    .A1(_1951_),
    .A2(_0353_));
 sg13g2_o21ai_1 _3014_ (.B1(_0354_),
    .Y(_0069_),
    .A1(_1940_),
    .A2(_0352_));
 sg13g2_nand3_1 _3015_ (.B(_0342_),
    .C(_1940_),
    .A(net92),
    .Y(_0355_));
 sg13g2_nor3_1 _3016_ (.A(_1939_),
    .B(_1951_),
    .C(_0355_),
    .Y(_0356_));
 sg13g2_a21oi_1 _3017_ (.A1(_1939_),
    .A2(_0355_),
    .Y(_0357_),
    .B1(_0356_));
 sg13g2_nand2_1 _3018_ (.Y(_0358_),
    .A(_1939_),
    .B(_1951_));
 sg13g2_o21ai_1 _3019_ (.B1(_0358_),
    .Y(_0070_),
    .A1(_1943_),
    .A2(_0357_));
 sg13g2_inv_1 _3020_ (.Y(_0359_),
    .A(\gray_sobel0.out_px_sobel[0] ));
 sg13g2_inv_1 _3021_ (.Y(_0360_),
    .A(\gray_sobel0.sobel0.px_ready ));
 sg13g2_buf_1 _3022_ (.A(\gray_sobel0.sobel0.sobel.pix2_2[6] ),
    .X(_0361_));
 sg13g2_buf_2 _3023_ (.A(\gray_sobel0.sobel0.sobel.pix0_0[6] ),
    .X(_0362_));
 sg13g2_buf_1 _3024_ (.A(\gray_sobel0.sobel0.sobel.pix0_2[6] ),
    .X(_0363_));
 sg13g2_xor2_1 _3025_ (.B(_0363_),
    .A(_0362_),
    .X(_0364_));
 sg13g2_buf_8 _3026_ (.A(\gray_sobel0.sobel0.sobel.pix0_0[4] ),
    .X(_0365_));
 sg13g2_buf_8 _3027_ (.A(\gray_sobel0.sobel0.sobel.pix0_2[4] ),
    .X(_0366_));
 sg13g2_nor2b_1 _3028_ (.A(_0365_),
    .B_N(_0366_),
    .Y(_0367_));
 sg13g2_buf_1 _3029_ (.A(\gray_sobel0.sobel0.sobel.pix0_0[5] ),
    .X(_0368_));
 sg13g2_buf_1 _3030_ (.A(\gray_sobel0.sobel0.sobel.pix0_2[5] ),
    .X(_0369_));
 sg13g2_nor2b_1 _3031_ (.A(net107),
    .B_N(net106),
    .Y(_0370_));
 sg13g2_nand2b_1 _3032_ (.Y(_0371_),
    .B(net107),
    .A_N(net106));
 sg13g2_o21ai_1 _3033_ (.B1(_0371_),
    .Y(_0372_),
    .A1(_0367_),
    .A2(_0370_));
 sg13g2_buf_2 _3034_ (.A(_0372_),
    .X(_0373_));
 sg13g2_buf_1 _3035_ (.A(\gray_sobel0.sobel0.sobel.pix0_2[1] ),
    .X(_0374_));
 sg13g2_buf_2 _3036_ (.A(\gray_sobel0.sobel0.sobel.pix0_0[1] ),
    .X(_0375_));
 sg13g2_nand2b_1 _3037_ (.Y(_0376_),
    .B(_0375_),
    .A_N(_0374_));
 sg13g2_buf_8 _3038_ (.A(\gray_sobel0.sobel0.sobel.pix0_0[0] ),
    .X(_0377_));
 sg13g2_nand2b_1 _3039_ (.Y(_0378_),
    .B(_0377_),
    .A_N(\gray_sobel0.sobel0.sobel.pix0_2[0] ));
 sg13g2_buf_2 _3040_ (.A(_0378_),
    .X(_0379_));
 sg13g2_nor2b_1 _3041_ (.A(_0375_),
    .B_N(_0374_),
    .Y(_0380_));
 sg13g2_a21o_1 _3042_ (.A2(_0379_),
    .A1(_0376_),
    .B1(_0380_),
    .X(_0381_));
 sg13g2_buf_1 _3043_ (.A(\gray_sobel0.sobel0.sobel.pix0_2[3] ),
    .X(_0382_));
 sg13g2_nor2b_1 _3044_ (.A(net105),
    .B_N(\gray_sobel0.sobel0.sobel.pix0_0[3] ),
    .Y(_0383_));
 sg13g2_buf_1 _3045_ (.A(\gray_sobel0.sobel0.sobel.pix0_2[2] ),
    .X(_0384_));
 sg13g2_buf_1 _3046_ (.A(\gray_sobel0.sobel0.sobel.pix0_0[2] ),
    .X(_0385_));
 sg13g2_nor2b_1 _3047_ (.A(net104),
    .B_N(net103),
    .Y(_0386_));
 sg13g2_buf_2 _3048_ (.A(_0386_),
    .X(_0387_));
 sg13g2_nor2_1 _3049_ (.A(_0383_),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_nand2b_1 _3050_ (.Y(_0389_),
    .B(net104),
    .A_N(net103));
 sg13g2_buf_1 _3051_ (.A(\gray_sobel0.sobel0.sobel.pix0_0[3] ),
    .X(_0390_));
 sg13g2_nand2b_1 _3052_ (.Y(_0391_),
    .B(net105),
    .A_N(_0390_));
 sg13g2_o21ai_1 _3053_ (.B1(_0391_),
    .Y(_0392_),
    .A1(_0383_),
    .A2(_0389_));
 sg13g2_a21oi_1 _3054_ (.A1(_0381_),
    .A2(_0388_),
    .Y(_0393_),
    .B1(_0392_));
 sg13g2_buf_1 _3055_ (.A(_0393_),
    .X(_0394_));
 sg13g2_nand2b_1 _3056_ (.Y(_0395_),
    .B(_0365_),
    .A_N(_0366_));
 sg13g2_o21ai_1 _3057_ (.B1(_0371_),
    .Y(_0396_),
    .A1(_0395_),
    .A2(_0370_));
 sg13g2_a21oi_1 _3058_ (.A1(_0373_),
    .A2(net65),
    .Y(_0397_),
    .B1(_0396_));
 sg13g2_xnor2_1 _3059_ (.Y(_0398_),
    .A(_0364_),
    .B(_0397_));
 sg13g2_nand2_1 _3060_ (.Y(_0399_),
    .A(net109),
    .B(_0398_));
 sg13g2_buf_2 _3061_ (.A(\gray_sobel0.sobel0.sobel.pix2_0[6] ),
    .X(_0400_));
 sg13g2_inv_1 _3062_ (.Y(_0401_),
    .A(_0400_));
 sg13g2_o21ai_1 _3063_ (.B1(_0401_),
    .Y(_0402_),
    .A1(net109),
    .A2(_0398_));
 sg13g2_nand2_1 _3064_ (.Y(_0403_),
    .A(_0399_),
    .B(_0402_));
 sg13g2_buf_1 _3065_ (.A(\gray_sobel0.sobel0.sobel.pix2_2[7] ),
    .X(_0404_));
 sg13g2_xnor2_1 _3066_ (.Y(_0405_),
    .A(net101),
    .B(\gray_sobel0.sobel0.sobel.pix0_0[7] ));
 sg13g2_buf_2 _3067_ (.A(\gray_sobel0.sobel0.sobel.pix2_0[7] ),
    .X(_0406_));
 sg13g2_xor2_1 _3068_ (.B(\gray_sobel0.sobel0.sobel.pix0_2[7] ),
    .A(_0406_),
    .X(_0407_));
 sg13g2_xnor2_1 _3069_ (.Y(_0408_),
    .A(_0405_),
    .B(_0407_));
 sg13g2_buf_2 _3070_ (.A(_0408_),
    .X(_0409_));
 sg13g2_inv_1 _3071_ (.Y(_0410_),
    .A(\gray_sobel0.sobel0.sobel.pix0_2[6] ));
 sg13g2_and2_1 _3072_ (.A(_0410_),
    .B(_0373_),
    .X(_0411_));
 sg13g2_nor2b_1 _3073_ (.A(_0366_),
    .B_N(_0365_),
    .Y(_0412_));
 sg13g2_nand2b_1 _3074_ (.Y(_0413_),
    .B(net106),
    .A_N(net107));
 sg13g2_nor2b_1 _3075_ (.A(net106),
    .B_N(net107),
    .Y(_0414_));
 sg13g2_a21oi_1 _3076_ (.A1(_0412_),
    .A2(_0413_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_inv_1 _3077_ (.Y(_0416_),
    .A(_0362_));
 sg13g2_o21ai_1 _3078_ (.B1(_0416_),
    .Y(_0417_),
    .A1(net108),
    .A2(_0415_));
 sg13g2_a21oi_2 _3079_ (.B1(_0417_),
    .Y(_0418_),
    .A2(net65),
    .A1(_0411_));
 sg13g2_nand2_1 _3080_ (.Y(_0419_),
    .A(net108),
    .B(_0415_));
 sg13g2_a21oi_2 _3081_ (.B1(_0419_),
    .Y(_0420_),
    .A2(net65),
    .A1(_0373_));
 sg13g2_nor2_1 _3082_ (.A(_0418_),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_xnor2_1 _3083_ (.Y(_0422_),
    .A(_0409_),
    .B(_0421_));
 sg13g2_inv_1 _3084_ (.Y(_0423_),
    .A(\gray_sobel0.sobel0.sobel.pix1_2[5] ));
 sg13g2_nand2b_1 _3085_ (.Y(_0424_),
    .B(\gray_sobel0.sobel0.sobel.pix1_0[4] ),
    .A_N(\gray_sobel0.sobel0.sobel.pix1_2[4] ));
 sg13g2_nor2b_1 _3086_ (.A(\gray_sobel0.sobel0.sobel.pix1_0[2] ),
    .B_N(\gray_sobel0.sobel0.sobel.pix1_2[2] ),
    .Y(_0425_));
 sg13g2_buf_1 _3087_ (.A(\gray_sobel0.sobel0.sobel.pix1_0[3] ),
    .X(_0426_));
 sg13g2_nand2b_1 _3088_ (.Y(_0427_),
    .B(_0426_),
    .A_N(\gray_sobel0.sobel0.sobel.pix1_2[3] ));
 sg13g2_nor2b_1 _3089_ (.A(_0426_),
    .B_N(\gray_sobel0.sobel0.sobel.pix1_2[3] ),
    .Y(_0428_));
 sg13g2_a21o_1 _3090_ (.A2(_0427_),
    .A1(_0425_),
    .B1(_0428_),
    .X(_0429_));
 sg13g2_inv_1 _3091_ (.Y(_0430_),
    .A(\gray_sobel0.sobel0.sobel.pix1_2[3] ));
 sg13g2_inv_1 _3092_ (.Y(_0431_),
    .A(\gray_sobel0.sobel0.sobel.pix1_2[4] ));
 sg13g2_nor2b_1 _3093_ (.A(\gray_sobel0.sobel0.sobel.pix1_2[2] ),
    .B_N(\gray_sobel0.sobel0.sobel.pix1_0[2] ),
    .Y(_0432_));
 sg13g2_buf_1 _3094_ (.A(_0432_),
    .X(_0433_));
 sg13g2_a221oi_1 _3095_ (.B2(\gray_sobel0.sobel0.sobel.pix1_0[4] ),
    .C1(_0433_),
    .B1(_0431_),
    .A1(_0426_),
    .Y(_0434_),
    .A2(_0430_));
 sg13g2_buf_1 _3096_ (.A(\gray_sobel0.sobel0.sobel.pix1_0[1] ),
    .X(_0435_));
 sg13g2_buf_1 _3097_ (.A(\gray_sobel0.sobel0.sobel.pix1_2[1] ),
    .X(_0436_));
 sg13g2_nand2b_1 _3098_ (.Y(_0437_),
    .B(_0436_),
    .A_N(_0435_));
 sg13g2_buf_2 _3099_ (.A(\gray_sobel0.sobel0.sobel.pix1_2[0] ),
    .X(_0438_));
 sg13g2_buf_2 _3100_ (.A(\gray_sobel0.sobel0.sobel.pix1_0[0] ),
    .X(_0439_));
 sg13g2_nor2b_1 _3101_ (.A(_0438_),
    .B_N(_0439_),
    .Y(_0440_));
 sg13g2_nor2b_1 _3102_ (.A(_0436_),
    .B_N(_0435_),
    .Y(_0441_));
 sg13g2_a21oi_2 _3103_ (.B1(_0441_),
    .Y(_0442_),
    .A2(_0440_),
    .A1(_0437_));
 sg13g2_nand2b_1 _3104_ (.Y(_0443_),
    .B(\gray_sobel0.sobel0.sobel.pix1_2[4] ),
    .A_N(\gray_sobel0.sobel0.sobel.pix1_0[4] ));
 sg13g2_inv_1 _3105_ (.Y(_0444_),
    .A(_0443_));
 sg13g2_a221oi_1 _3106_ (.B2(_0442_),
    .C1(_0444_),
    .B1(_0434_),
    .A1(_0424_),
    .Y(_0445_),
    .A2(_0429_));
 sg13g2_buf_2 _3107_ (.A(_0445_),
    .X(_0446_));
 sg13g2_nor2_1 _3108_ (.A(_0423_),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_buf_1 _3109_ (.A(\gray_sobel0.sobel0.sobel.pix1_0[5] ),
    .X(_0448_));
 sg13g2_a21oi_1 _3110_ (.A1(_0423_),
    .A2(_0446_),
    .Y(_0449_),
    .B1(_0448_));
 sg13g2_nor2_1 _3111_ (.A(_0447_),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_nand2b_1 _3112_ (.Y(_0451_),
    .B(\gray_sobel0.sobel0.sobel.pix1_2[6] ),
    .A_N(\gray_sobel0.sobel0.sobel.pix1_0[6] ));
 sg13g2_inv_1 _3113_ (.Y(_0452_),
    .A(\gray_sobel0.sobel0.sobel.pix1_2[6] ));
 sg13g2_nand2_1 _3114_ (.Y(_0453_),
    .A(\gray_sobel0.sobel0.sobel.pix1_0[6] ),
    .B(_0452_));
 sg13g2_nand2_1 _3115_ (.Y(_0454_),
    .A(_0451_),
    .B(_0453_));
 sg13g2_xnor2_1 _3116_ (.Y(_0455_),
    .A(_0450_),
    .B(_0454_));
 sg13g2_xor2_1 _3117_ (.B(_0455_),
    .A(_0422_),
    .X(_0456_));
 sg13g2_xor2_1 _3118_ (.B(_0456_),
    .A(_0403_),
    .X(_0457_));
 sg13g2_buf_1 _3119_ (.A(\gray_sobel0.sobel0.sobel.pix2_2[0] ),
    .X(_0458_));
 sg13g2_xor2_1 _3120_ (.B(\gray_sobel0.sobel0.sobel.pix0_2[0] ),
    .A(_0377_),
    .X(_0459_));
 sg13g2_buf_1 _3121_ (.A(_0459_),
    .X(_0460_));
 sg13g2_nand2_1 _3122_ (.Y(_0461_),
    .A(net100),
    .B(net77));
 sg13g2_xnor2_1 _3123_ (.Y(_0462_),
    .A(_0439_),
    .B(_0438_));
 sg13g2_xnor2_1 _3124_ (.Y(_0463_),
    .A(_0375_),
    .B(_0374_));
 sg13g2_buf_2 _3125_ (.A(_0463_),
    .X(_0464_));
 sg13g2_xor2_1 _3126_ (.B(_0379_),
    .A(_0464_),
    .X(_0465_));
 sg13g2_buf_2 _3127_ (.A(_0465_),
    .X(_0466_));
 sg13g2_buf_1 _3128_ (.A(\gray_sobel0.sobel0.sobel.pix2_0[1] ),
    .X(_0467_));
 sg13g2_buf_1 _3129_ (.A(\gray_sobel0.sobel0.sobel.pix2_2[1] ),
    .X(_0468_));
 sg13g2_xnor2_1 _3130_ (.Y(_0469_),
    .A(_0467_),
    .B(_0468_));
 sg13g2_xnor2_1 _3131_ (.Y(_0470_),
    .A(_0466_),
    .B(_0469_));
 sg13g2_and3_1 _3132_ (.X(_0471_),
    .A(_0461_),
    .B(_0462_),
    .C(_0470_));
 sg13g2_xor2_1 _3133_ (.B(_0438_),
    .A(_0439_),
    .X(_0472_));
 sg13g2_nor3_1 _3134_ (.A(_0466_),
    .B(_0472_),
    .C(_0469_),
    .Y(_0473_));
 sg13g2_nor2b_1 _3135_ (.A(_0469_),
    .B_N(_0464_),
    .Y(_0474_));
 sg13g2_nor2_1 _3136_ (.A(net100),
    .B(_0460_),
    .Y(_0475_));
 sg13g2_o21ai_1 _3137_ (.B1(_0475_),
    .Y(_0476_),
    .A1(_0462_),
    .A2(_0474_));
 sg13g2_nor2b_1 _3138_ (.A(_0473_),
    .B_N(_0476_),
    .Y(_0477_));
 sg13g2_nor3_1 _3139_ (.A(net100),
    .B(_0464_),
    .C(_0460_),
    .Y(_0478_));
 sg13g2_a21oi_1 _3140_ (.A1(_0466_),
    .A2(_0462_),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_nand2b_1 _3141_ (.Y(_0480_),
    .B(_0469_),
    .A_N(_0479_));
 sg13g2_buf_1 _3142_ (.A(\gray_sobel0.sobel0.sobel.pix2_0[0] ),
    .X(_0481_));
 sg13g2_buf_1 _3143_ (.A(_0481_),
    .X(_0482_));
 sg13g2_inv_1 _3144_ (.Y(_0483_),
    .A(net91));
 sg13g2_a21oi_1 _3145_ (.A1(_0477_),
    .A2(_0480_),
    .Y(_0484_),
    .B1(net76));
 sg13g2_xor2_1 _3146_ (.B(_0469_),
    .A(_0466_),
    .X(_0485_));
 sg13g2_nor3_1 _3147_ (.A(_0481_),
    .B(_0461_),
    .C(_0462_),
    .Y(_0486_));
 sg13g2_buf_8 _3148_ (.A(\gray_sobel0.sobel0.sobel.pix2_2[2] ),
    .X(_0487_));
 sg13g2_xnor2_1 _3149_ (.Y(_0488_),
    .A(\gray_sobel0.sobel0.sobel.pix2_0[2] ),
    .B(_0487_));
 sg13g2_xnor2_1 _3150_ (.Y(_0489_),
    .A(net103),
    .B(_0384_));
 sg13g2_buf_1 _3151_ (.A(_0489_),
    .X(_0490_));
 sg13g2_nand2b_1 _3152_ (.Y(_0491_),
    .B(net75),
    .A_N(_0488_));
 sg13g2_nand2b_1 _3153_ (.Y(_0492_),
    .B(_0488_),
    .A_N(net75));
 sg13g2_a21oi_2 _3154_ (.B1(_0380_),
    .Y(_0493_),
    .A2(_0379_),
    .A1(_0376_));
 sg13g2_a21oi_1 _3155_ (.A1(_0491_),
    .A2(_0492_),
    .Y(_0494_),
    .B1(_0493_));
 sg13g2_or2_1 _3156_ (.X(_0495_),
    .B(_0488_),
    .A(net75));
 sg13g2_nand2_1 _3157_ (.Y(_0496_),
    .A(_0490_),
    .B(_0488_));
 sg13g2_a21oi_1 _3158_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0497_),
    .B1(_0381_));
 sg13g2_nand2b_1 _3159_ (.Y(_0498_),
    .B(_0439_),
    .A_N(_0438_));
 sg13g2_nor2b_1 _3160_ (.A(_0435_),
    .B_N(_0436_),
    .Y(_0499_));
 sg13g2_nor2_1 _3161_ (.A(_0499_),
    .B(_0441_),
    .Y(_0500_));
 sg13g2_xnor2_1 _3162_ (.Y(_0501_),
    .A(_0498_),
    .B(_0500_));
 sg13g2_o21ai_1 _3163_ (.B1(_0501_),
    .Y(_0502_),
    .A1(_0494_),
    .A2(_0497_));
 sg13g2_buf_1 _3164_ (.A(_0502_),
    .X(_0503_));
 sg13g2_or3_1 _3165_ (.A(_0501_),
    .B(_0494_),
    .C(_0497_),
    .X(_0504_));
 sg13g2_buf_1 _3166_ (.A(_0504_),
    .X(_0505_));
 sg13g2_buf_1 _3167_ (.A(_0468_),
    .X(_0506_));
 sg13g2_nand2_1 _3168_ (.Y(_0507_),
    .A(_0506_),
    .B(_0466_));
 sg13g2_inv_1 _3169_ (.Y(_0508_),
    .A(_0467_));
 sg13g2_o21ai_1 _3170_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0468_),
    .A2(_0466_));
 sg13g2_nand2_1 _3171_ (.Y(_0510_),
    .A(_0507_),
    .B(_0509_));
 sg13g2_a221oi_1 _3172_ (.B2(_0505_),
    .C1(_0510_),
    .B1(_0503_),
    .A1(_0485_),
    .Y(_0511_),
    .A2(_0486_));
 sg13g2_nand2_1 _3173_ (.Y(_0512_),
    .A(_0485_),
    .B(_0486_));
 sg13g2_and4_1 _3174_ (.A(_0510_),
    .B(_0512_),
    .C(_0503_),
    .D(_0505_),
    .X(_0513_));
 sg13g2_or4_1 _3175_ (.A(_0471_),
    .B(_0484_),
    .C(_0511_),
    .D(_0513_),
    .X(_0514_));
 sg13g2_buf_2 _3176_ (.A(_0514_),
    .X(_0515_));
 sg13g2_nand3_1 _3177_ (.B(_0509_),
    .C(_0501_),
    .A(_0507_),
    .Y(_0516_));
 sg13g2_nor2_1 _3178_ (.A(_0494_),
    .B(_0497_),
    .Y(_0517_));
 sg13g2_a21oi_1 _3179_ (.A1(_0507_),
    .A2(_0509_),
    .Y(_0518_),
    .B1(_0501_));
 sg13g2_a21o_1 _3180_ (.A2(_0517_),
    .A1(_0516_),
    .B1(_0518_),
    .X(_0519_));
 sg13g2_inv_1 _3181_ (.Y(_0520_),
    .A(net103));
 sg13g2_a221oi_1 _3182_ (.B2(_0379_),
    .C1(_0380_),
    .B1(_0376_),
    .A1(_0520_),
    .Y(_0521_),
    .A2(net104));
 sg13g2_buf_2 _3183_ (.A(_0521_),
    .X(_0522_));
 sg13g2_xnor2_1 _3184_ (.Y(_0523_),
    .A(\gray_sobel0.sobel0.sobel.pix0_0[3] ),
    .B(net105));
 sg13g2_buf_2 _3185_ (.A(_0523_),
    .X(_0524_));
 sg13g2_buf_1 _3186_ (.A(\gray_sobel0.sobel0.sobel.pix2_0[3] ),
    .X(_0525_));
 sg13g2_buf_2 _3187_ (.A(\gray_sobel0.sobel0.sobel.pix2_2[3] ),
    .X(_0526_));
 sg13g2_xnor2_1 _3188_ (.Y(_0527_),
    .A(_0525_),
    .B(_0526_));
 sg13g2_xnor2_1 _3189_ (.Y(_0528_),
    .A(_0524_),
    .B(_0527_));
 sg13g2_o21ai_1 _3190_ (.B1(_0528_),
    .Y(_0529_),
    .A1(_0387_),
    .A2(_0522_));
 sg13g2_buf_1 _3191_ (.A(_0529_),
    .X(_0530_));
 sg13g2_or3_1 _3192_ (.A(_0387_),
    .B(_0528_),
    .C(_0522_),
    .X(_0531_));
 sg13g2_buf_1 _3193_ (.A(_0531_),
    .X(_0532_));
 sg13g2_nor2_1 _3194_ (.A(_0425_),
    .B(_0433_),
    .Y(_0533_));
 sg13g2_xor2_1 _3195_ (.B(_0533_),
    .A(_0442_),
    .X(_0534_));
 sg13g2_a21oi_1 _3196_ (.A1(_0530_),
    .A2(_0532_),
    .Y(_0535_),
    .B1(_0534_));
 sg13g2_and3_1 _3197_ (.X(_0536_),
    .A(_0534_),
    .B(_0530_),
    .C(_0532_));
 sg13g2_inv_1 _3198_ (.Y(_0537_),
    .A(\gray_sobel0.sobel0.sobel.pix2_0[2] ));
 sg13g2_inv_1 _3199_ (.Y(_0538_),
    .A(_0487_));
 sg13g2_nand2_1 _3200_ (.Y(_0539_),
    .A(_0538_),
    .B(net75));
 sg13g2_or2_1 _3201_ (.X(_0540_),
    .B(net75),
    .A(_0487_));
 sg13g2_mux2_1 _3202_ (.A0(_0539_),
    .A1(_0540_),
    .S(_0493_),
    .X(_0541_));
 sg13g2_nor2_1 _3203_ (.A(_0538_),
    .B(net75),
    .Y(_0542_));
 sg13g2_and2_1 _3204_ (.A(_0487_),
    .B(net75),
    .X(_0543_));
 sg13g2_mux2_1 _3205_ (.A0(_0542_),
    .A1(_0543_),
    .S(_0493_),
    .X(_0544_));
 sg13g2_a21oi_1 _3206_ (.A1(_0537_),
    .A2(_0541_),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_o21ai_1 _3207_ (.B1(_0545_),
    .Y(_0546_),
    .A1(_0535_),
    .A2(_0536_));
 sg13g2_a21o_1 _3208_ (.A2(_0541_),
    .A1(_0537_),
    .B1(_0544_),
    .X(_0547_));
 sg13g2_a21o_1 _3209_ (.A2(_0532_),
    .A1(_0530_),
    .B1(_0534_),
    .X(_0548_));
 sg13g2_nand3_1 _3210_ (.B(_0530_),
    .C(_0532_),
    .A(_0534_),
    .Y(_0549_));
 sg13g2_nand3_1 _3211_ (.B(_0548_),
    .C(_0549_),
    .A(_0547_),
    .Y(_0550_));
 sg13g2_nand3_1 _3212_ (.B(_0546_),
    .C(_0550_),
    .A(_0519_),
    .Y(_0551_));
 sg13g2_buf_1 _3213_ (.A(_0551_),
    .X(_0552_));
 sg13g2_a21oi_1 _3214_ (.A1(_0546_),
    .A2(_0550_),
    .Y(_0553_),
    .B1(_0519_));
 sg13g2_a21oi_1 _3215_ (.A1(_0515_),
    .A2(_0552_),
    .Y(_0554_),
    .B1(_0553_));
 sg13g2_buf_2 _3216_ (.A(\gray_sobel0.sobel0.sobel.pix2_0[4] ),
    .X(_0555_));
 sg13g2_inv_1 _3217_ (.Y(_0556_),
    .A(_0555_));
 sg13g2_buf_1 _3218_ (.A(\gray_sobel0.sobel0.sobel.pix2_2[4] ),
    .X(_0557_));
 sg13g2_xnor2_1 _3219_ (.Y(_0558_),
    .A(_0365_),
    .B(_0366_));
 sg13g2_xnor2_1 _3220_ (.Y(_0559_),
    .A(_0557_),
    .B(_0558_));
 sg13g2_xnor2_1 _3221_ (.Y(_0560_),
    .A(_0556_),
    .B(_0559_));
 sg13g2_buf_2 _3222_ (.A(_0560_),
    .X(_0561_));
 sg13g2_xnor2_1 _3223_ (.Y(_0562_),
    .A(_0561_),
    .B(net65));
 sg13g2_inv_1 _3224_ (.Y(_0563_),
    .A(\gray_sobel0.sobel0.sobel.pix1_0[2] ));
 sg13g2_nand2b_1 _3225_ (.Y(_0564_),
    .B(_0435_),
    .A_N(_0436_));
 sg13g2_a221oi_1 _3226_ (.B2(_0498_),
    .C1(_0499_),
    .B1(_0564_),
    .A1(_0563_),
    .Y(_0565_),
    .A2(\gray_sobel0.sobel0.sobel.pix1_2[2] ));
 sg13g2_or2_1 _3227_ (.X(_0566_),
    .B(_0565_),
    .A(_0433_));
 sg13g2_nor2b_1 _3228_ (.A(_0428_),
    .B_N(_0427_),
    .Y(_0567_));
 sg13g2_xnor2_1 _3229_ (.Y(_0568_),
    .A(_0566_),
    .B(_0567_));
 sg13g2_or2_1 _3230_ (.X(_0569_),
    .B(_0568_),
    .A(_0562_));
 sg13g2_buf_1 _3231_ (.A(_0569_),
    .X(_0570_));
 sg13g2_nor2_1 _3232_ (.A(_0526_),
    .B(_0524_),
    .Y(_0571_));
 sg13g2_or2_1 _3233_ (.X(_0572_),
    .B(_0522_),
    .A(_0387_));
 sg13g2_nand2b_1 _3234_ (.Y(_0573_),
    .B(_0385_),
    .A_N(_0384_));
 sg13g2_nand3b_1 _3235_ (.B(_0573_),
    .C(_0526_),
    .Y(_0574_),
    .A_N(_0524_));
 sg13g2_nand2_1 _3236_ (.Y(_0575_),
    .A(_0526_),
    .B(_0524_));
 sg13g2_mux2_1 _3237_ (.A0(_0574_),
    .A1(_0575_),
    .S(_0522_),
    .X(_0576_));
 sg13g2_inv_1 _3238_ (.Y(_0577_),
    .A(_0526_));
 sg13g2_nor2_1 _3239_ (.A(net89),
    .B(_0573_),
    .Y(_0578_));
 sg13g2_inv_2 _3240_ (.Y(_0579_),
    .A(_0525_));
 sg13g2_a21oi_1 _3241_ (.A1(_0524_),
    .A2(_0578_),
    .Y(_0580_),
    .B1(_0579_));
 sg13g2_nand2_1 _3242_ (.Y(_0581_),
    .A(_0577_),
    .B(_0524_));
 sg13g2_nor3_1 _3243_ (.A(_0387_),
    .B(_0522_),
    .C(_0581_),
    .Y(_0582_));
 sg13g2_a221oi_1 _3244_ (.B2(_0580_),
    .C1(_0582_),
    .B1(_0576_),
    .A1(_0571_),
    .Y(_0583_),
    .A2(_0572_));
 sg13g2_buf_1 _3245_ (.A(_0583_),
    .X(_0584_));
 sg13g2_nor2_1 _3246_ (.A(_0570_),
    .B(_0584_),
    .Y(_0585_));
 sg13g2_a21o_1 _3247_ (.A2(_0568_),
    .A1(_0562_),
    .B1(_0584_),
    .X(_0586_));
 sg13g2_a21oi_1 _3248_ (.A1(_0545_),
    .A2(_0549_),
    .Y(_0587_),
    .B1(_0535_));
 sg13g2_a21oi_1 _3249_ (.A1(_0570_),
    .A2(_0586_),
    .Y(_0588_),
    .B1(_0587_));
 sg13g2_nor2_1 _3250_ (.A(_0585_),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_nor2_1 _3251_ (.A(_0554_),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_inv_1 _3252_ (.Y(_0591_),
    .A(_0557_));
 sg13g2_nand2_1 _3253_ (.Y(_0592_),
    .A(_0555_),
    .B(_0591_));
 sg13g2_nand2b_1 _3254_ (.Y(_0593_),
    .B(_0592_),
    .A_N(_0558_));
 sg13g2_nand2_1 _3255_ (.Y(_0594_),
    .A(_0558_),
    .B(_0592_));
 sg13g2_mux2_1 _3256_ (.A0(_0593_),
    .A1(_0594_),
    .S(net65),
    .X(_0595_));
 sg13g2_nand2_1 _3257_ (.Y(_0596_),
    .A(_0556_),
    .B(_0557_));
 sg13g2_and2_1 _3258_ (.A(_0595_),
    .B(_0596_),
    .X(_0597_));
 sg13g2_a21o_1 _3259_ (.A2(_0388_),
    .A1(_0381_),
    .B1(_0392_),
    .X(_0598_));
 sg13g2_a21oi_2 _3260_ (.B1(_0367_),
    .Y(_0599_),
    .A2(_0598_),
    .A1(_0395_));
 sg13g2_o21ai_1 _3261_ (.B1(_0430_),
    .Y(_0600_),
    .A1(_0433_),
    .A2(_0565_));
 sg13g2_buf_1 _3262_ (.A(_0600_),
    .X(_0601_));
 sg13g2_nand2b_1 _3263_ (.Y(_0602_),
    .B(\gray_sobel0.sobel0.sobel.pix1_2[3] ),
    .A_N(_0433_));
 sg13g2_o21ai_1 _3264_ (.B1(_0426_),
    .Y(_0603_),
    .A1(_0565_),
    .A2(_0602_));
 sg13g2_buf_1 _3265_ (.A(_0603_),
    .X(_0604_));
 sg13g2_buf_1 _3266_ (.A(\gray_sobel0.sobel0.sobel.pix2_2[5] ),
    .X(_0605_));
 sg13g2_buf_1 _3267_ (.A(\gray_sobel0.sobel0.sobel.pix2_0[5] ),
    .X(_0606_));
 sg13g2_nand2b_1 _3268_ (.Y(_0607_),
    .B(_0606_),
    .A_N(_0605_));
 sg13g2_buf_1 _3269_ (.A(_0605_),
    .X(_0608_));
 sg13g2_nand2b_1 _3270_ (.Y(_0609_),
    .B(net88),
    .A_N(net99));
 sg13g2_xnor2_1 _3271_ (.Y(_0610_),
    .A(net107),
    .B(net106));
 sg13g2_a21oi_1 _3272_ (.A1(_0607_),
    .A2(_0609_),
    .Y(_0611_),
    .B1(_0610_));
 sg13g2_or2_1 _3273_ (.X(_0612_),
    .B(_0605_),
    .A(_0606_));
 sg13g2_nand2_1 _3274_ (.Y(_0613_),
    .A(net99),
    .B(net88));
 sg13g2_xor2_1 _3275_ (.B(net106),
    .A(net107),
    .X(_0614_));
 sg13g2_a21oi_1 _3276_ (.A1(_0612_),
    .A2(_0613_),
    .Y(_0615_),
    .B1(_0614_));
 sg13g2_nand2_1 _3277_ (.Y(_0616_),
    .A(_0443_),
    .B(_0424_));
 sg13g2_o21ai_1 _3278_ (.B1(_0616_),
    .Y(_0617_),
    .A1(_0611_),
    .A2(_0615_));
 sg13g2_or3_1 _3279_ (.A(_0611_),
    .B(_0615_),
    .C(_0616_),
    .X(_0618_));
 sg13g2_and4_1 _3280_ (.A(_0601_),
    .B(_0604_),
    .C(_0617_),
    .D(_0618_),
    .X(_0619_));
 sg13g2_a22oi_1 _3281_ (.Y(_0620_),
    .B1(_0617_),
    .B2(_0618_),
    .A2(_0604_),
    .A1(_0601_));
 sg13g2_or3_1 _3282_ (.A(_0599_),
    .B(_0619_),
    .C(_0620_),
    .X(_0621_));
 sg13g2_o21ai_1 _3283_ (.B1(_0599_),
    .Y(_0622_),
    .A1(_0619_),
    .A2(_0620_));
 sg13g2_nand3_1 _3284_ (.B(_0621_),
    .C(_0622_),
    .A(_0597_),
    .Y(_0623_));
 sg13g2_a21o_1 _3285_ (.A2(_0622_),
    .A1(_0621_),
    .B1(_0597_),
    .X(_0624_));
 sg13g2_xnor2_1 _3286_ (.Y(_0625_),
    .A(_0555_),
    .B(_0559_));
 sg13g2_buf_2 _3287_ (.A(_0625_),
    .X(_0626_));
 sg13g2_nand2_1 _3288_ (.Y(_0627_),
    .A(_0626_),
    .B(net65));
 sg13g2_nand2_1 _3289_ (.Y(_0628_),
    .A(_0561_),
    .B(_0598_));
 sg13g2_a221oi_1 _3290_ (.B2(_0628_),
    .C1(_0536_),
    .B1(_0627_),
    .A1(_0547_),
    .Y(_0629_),
    .A2(_0548_));
 sg13g2_nor2_1 _3291_ (.A(_0568_),
    .B(_0584_),
    .Y(_0630_));
 sg13g2_and2_1 _3292_ (.A(_0629_),
    .B(_0630_),
    .X(_0631_));
 sg13g2_a21oi_1 _3293_ (.A1(_0623_),
    .A2(_0624_),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_or2_1 _3294_ (.X(_0633_),
    .B(_0615_),
    .A(_0611_));
 sg13g2_xor2_1 _3295_ (.B(_0599_),
    .A(_0633_),
    .X(_0634_));
 sg13g2_a21o_1 _3296_ (.A2(_0604_),
    .A1(_0601_),
    .B1(_0616_),
    .X(_0635_));
 sg13g2_nand3_1 _3297_ (.B(_0604_),
    .C(_0616_),
    .A(_0601_),
    .Y(_0636_));
 sg13g2_nand4_1 _3298_ (.B(_0596_),
    .C(_0635_),
    .A(_0595_),
    .Y(_0637_),
    .D(_0636_));
 sg13g2_a22oi_1 _3299_ (.Y(_0638_),
    .B1(_0635_),
    .B2(_0636_),
    .A2(_0596_),
    .A1(_0595_));
 sg13g2_a21o_1 _3300_ (.A2(_0637_),
    .A1(_0634_),
    .B1(_0638_),
    .X(_0639_));
 sg13g2_buf_1 _3301_ (.A(_0639_),
    .X(_0640_));
 sg13g2_xor2_1 _3302_ (.B(net109),
    .A(_0400_),
    .X(_0641_));
 sg13g2_xnor2_1 _3303_ (.Y(_0642_),
    .A(_0364_),
    .B(_0641_));
 sg13g2_xnor2_1 _3304_ (.Y(_0643_),
    .A(_0642_),
    .B(_0397_));
 sg13g2_buf_1 _3305_ (.A(_0643_),
    .X(_0644_));
 sg13g2_xor2_1 _3306_ (.B(\gray_sobel0.sobel0.sobel.pix1_2[5] ),
    .A(_0448_),
    .X(_0645_));
 sg13g2_nand2b_1 _3307_ (.Y(_0646_),
    .B(_0645_),
    .A_N(_0446_));
 sg13g2_inv_1 _3308_ (.Y(_0647_),
    .A(_0645_));
 sg13g2_nand2_1 _3309_ (.Y(_0648_),
    .A(_0446_),
    .B(_0647_));
 sg13g2_and2_1 _3310_ (.A(_0646_),
    .B(_0648_),
    .X(_0649_));
 sg13g2_nor2_1 _3311_ (.A(net88),
    .B(_0614_),
    .Y(_0650_));
 sg13g2_nor2_1 _3312_ (.A(net88),
    .B(_0610_),
    .Y(_0651_));
 sg13g2_mux2_1 _3313_ (.A0(_0650_),
    .A1(_0651_),
    .S(_0599_),
    .X(_0652_));
 sg13g2_inv_1 _3314_ (.Y(_0653_),
    .A(net99));
 sg13g2_xnor2_1 _3315_ (.Y(_0654_),
    .A(_0446_),
    .B(_0647_));
 sg13g2_nor2_1 _3316_ (.A(_0653_),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_nand2_1 _3317_ (.Y(_0656_),
    .A(net88),
    .B(_0614_));
 sg13g2_nand2_1 _3318_ (.Y(_0657_),
    .A(net88),
    .B(_0610_));
 sg13g2_mux2_1 _3319_ (.A0(_0656_),
    .A1(_0657_),
    .S(_0599_),
    .X(_0658_));
 sg13g2_a22oi_1 _3320_ (.Y(_0659_),
    .B1(_0655_),
    .B2(_0658_),
    .A2(_0652_),
    .A1(_0649_));
 sg13g2_buf_1 _3321_ (.A(_0659_),
    .X(_0660_));
 sg13g2_and3_1 _3322_ (.X(_0661_),
    .A(_0640_),
    .B(net50),
    .C(_0660_));
 sg13g2_nand2_1 _3323_ (.Y(_0662_),
    .A(_0632_),
    .B(_0661_));
 sg13g2_nand3_1 _3324_ (.B(_0568_),
    .C(_0584_),
    .A(_0562_),
    .Y(_0663_));
 sg13g2_nand3_1 _3325_ (.B(_0570_),
    .C(_0586_),
    .A(_0587_),
    .Y(_0664_));
 sg13g2_a221oi_1 _3326_ (.B2(_0664_),
    .C1(_0553_),
    .B1(_0663_),
    .A1(_0515_),
    .Y(_0665_),
    .A2(_0552_));
 sg13g2_buf_1 _3327_ (.A(_0665_),
    .X(_0666_));
 sg13g2_and2_1 _3328_ (.A(_0587_),
    .B(_0562_),
    .X(_0667_));
 sg13g2_buf_1 _3329_ (.A(_0667_),
    .X(_0668_));
 sg13g2_and2_1 _3330_ (.A(_0568_),
    .B(_0584_),
    .X(_0669_));
 sg13g2_buf_1 _3331_ (.A(_0669_),
    .X(_0670_));
 sg13g2_and2_1 _3332_ (.A(_0668_),
    .B(_0670_),
    .X(_0671_));
 sg13g2_buf_1 _3333_ (.A(_0671_),
    .X(_0672_));
 sg13g2_o21ai_1 _3334_ (.B1(_0661_),
    .Y(_0673_),
    .A1(_0666_),
    .A2(_0672_));
 sg13g2_o21ai_1 _3335_ (.B1(_0673_),
    .Y(_0674_),
    .A1(_0590_),
    .A2(_0662_));
 sg13g2_nor3_1 _3336_ (.A(_0640_),
    .B(net50),
    .C(_0660_),
    .Y(_0675_));
 sg13g2_o21ai_1 _3337_ (.B1(_0632_),
    .Y(_0676_),
    .A1(_0554_),
    .A2(_0589_));
 sg13g2_buf_1 _3338_ (.A(_0676_),
    .X(_0677_));
 sg13g2_nor2_1 _3339_ (.A(_0666_),
    .B(_0672_),
    .Y(_0678_));
 sg13g2_a21oi_2 _3340_ (.B1(_0638_),
    .Y(_0679_),
    .A2(_0637_),
    .A1(_0634_));
 sg13g2_a221oi_1 _3341_ (.B2(_0648_),
    .C1(_0652_),
    .B1(_0646_),
    .A1(net99),
    .Y(_0680_),
    .A2(_0658_));
 sg13g2_o21ai_1 _3342_ (.B1(_0660_),
    .Y(_0681_),
    .A1(_0680_),
    .A2(net50));
 sg13g2_nor2_1 _3343_ (.A(net50),
    .B(_0660_),
    .Y(_0682_));
 sg13g2_a21o_1 _3344_ (.A2(_0681_),
    .A1(_0679_),
    .B1(_0682_),
    .X(_0683_));
 sg13g2_and3_1 _3345_ (.X(_0684_),
    .A(_0677_),
    .B(_0678_),
    .C(_0683_));
 sg13g2_a221oi_1 _3346_ (.B2(_0640_),
    .C1(_0666_),
    .B1(net50),
    .A1(_0668_),
    .Y(_0685_),
    .A2(_0670_));
 sg13g2_o21ai_1 _3347_ (.B1(_0680_),
    .Y(_0686_),
    .A1(_0640_),
    .A2(net50));
 sg13g2_a21oi_1 _3348_ (.A1(_0677_),
    .A2(_0685_),
    .Y(_0687_),
    .B1(_0686_));
 sg13g2_or4_1 _3349_ (.A(_0674_),
    .B(_0675_),
    .C(_0684_),
    .D(_0687_),
    .X(_0688_));
 sg13g2_xnor2_1 _3350_ (.Y(_0689_),
    .A(_0457_),
    .B(_0688_));
 sg13g2_nand2_1 _3351_ (.Y(_0690_),
    .A(_0677_),
    .B(_0678_));
 sg13g2_a21oi_1 _3352_ (.A1(net99),
    .A2(_0658_),
    .Y(_0691_),
    .B1(_0652_));
 sg13g2_xnor2_1 _3353_ (.Y(_0692_),
    .A(_0654_),
    .B(net50));
 sg13g2_xnor2_1 _3354_ (.Y(_0693_),
    .A(_0679_),
    .B(_0692_));
 sg13g2_xnor2_1 _3355_ (.Y(_0694_),
    .A(_0691_),
    .B(_0693_));
 sg13g2_xor2_1 _3356_ (.B(_0694_),
    .A(_0690_),
    .X(_0695_));
 sg13g2_buf_2 _3357_ (.A(_0695_),
    .X(_0696_));
 sg13g2_nor2b_1 _3358_ (.A(_0553_),
    .B_N(_0552_),
    .Y(_0697_));
 sg13g2_xnor2_1 _3359_ (.Y(_0698_),
    .A(_0472_),
    .B(_0470_));
 sg13g2_buf_2 _3360_ (.A(_0698_),
    .X(_0699_));
 sg13g2_inv_2 _3361_ (.Y(_0700_),
    .A(net100));
 sg13g2_xnor2_1 _3362_ (.Y(_0701_),
    .A(_0700_),
    .B(net77));
 sg13g2_buf_1 _3363_ (.A(_0701_),
    .X(_0702_));
 sg13g2_and2_1 _3364_ (.A(_0481_),
    .B(net68),
    .X(_0703_));
 sg13g2_a21o_1 _3365_ (.A2(_0475_),
    .A1(net76),
    .B1(_0703_),
    .X(_0704_));
 sg13g2_nor3_1 _3366_ (.A(net91),
    .B(_0461_),
    .C(_0699_),
    .Y(_0705_));
 sg13g2_a21oi_1 _3367_ (.A1(_0699_),
    .A2(_0704_),
    .Y(_0706_),
    .B1(_0705_));
 sg13g2_a21oi_1 _3368_ (.A1(_0503_),
    .A2(_0505_),
    .Y(_0707_),
    .B1(_0510_));
 sg13g2_nand3_1 _3369_ (.B(_0503_),
    .C(_0505_),
    .A(_0510_),
    .Y(_0708_));
 sg13g2_nand2b_1 _3370_ (.Y(_0709_),
    .B(_0708_),
    .A_N(_0707_));
 sg13g2_and2_1 _3371_ (.A(_0485_),
    .B(_0486_),
    .X(_0710_));
 sg13g2_nor3_1 _3372_ (.A(_0710_),
    .B(_0471_),
    .C(_0484_),
    .Y(_0711_));
 sg13g2_xnor2_1 _3373_ (.Y(_0712_),
    .A(_0709_),
    .B(_0711_));
 sg13g2_nor2_1 _3374_ (.A(_0706_),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_nand2_1 _3375_ (.Y(_0714_),
    .A(_0697_),
    .B(_0713_));
 sg13g2_nor2_1 _3376_ (.A(_0629_),
    .B(_0668_),
    .Y(_0715_));
 sg13g2_and2_1 _3377_ (.A(_0623_),
    .B(_0624_),
    .X(_0716_));
 sg13g2_buf_1 _3378_ (.A(_0716_),
    .X(_0717_));
 sg13g2_mux2_1 _3379_ (.A0(_0630_),
    .A1(_0670_),
    .S(_0717_),
    .X(_0718_));
 sg13g2_nor2_1 _3380_ (.A(_0630_),
    .B(_0670_),
    .Y(_0719_));
 sg13g2_mux2_1 _3381_ (.A0(_0629_),
    .A1(_0668_),
    .S(_0717_),
    .X(_0720_));
 sg13g2_a21o_1 _3382_ (.A2(_0552_),
    .A1(_0515_),
    .B1(_0553_),
    .X(_0721_));
 sg13g2_a221oi_1 _3383_ (.B2(_0720_),
    .C1(_0721_),
    .B1(_0719_),
    .A1(_0715_),
    .Y(_0722_),
    .A2(_0718_));
 sg13g2_or2_1 _3384_ (.X(_0723_),
    .B(_0722_),
    .A(_0714_));
 sg13g2_buf_1 _3385_ (.A(_0723_),
    .X(_0724_));
 sg13g2_nor2_1 _3386_ (.A(_0696_),
    .B(_0724_),
    .Y(_0725_));
 sg13g2_and2_1 _3387_ (.A(_0689_),
    .B(_0725_),
    .X(_0726_));
 sg13g2_nand2_1 _3388_ (.Y(_0727_),
    .A(_0654_),
    .B(_0691_));
 sg13g2_nand4_1 _3389_ (.B(_0679_),
    .C(_0677_),
    .A(_0727_),
    .Y(_0728_),
    .D(_0678_));
 sg13g2_xnor2_1 _3390_ (.Y(_0729_),
    .A(_0403_),
    .B(_0456_));
 sg13g2_and2_1 _3391_ (.A(_0729_),
    .B(_0660_),
    .X(_0730_));
 sg13g2_nand3_1 _3392_ (.B(_0677_),
    .C(_0678_),
    .A(_0457_),
    .Y(_0731_));
 sg13g2_nand2_1 _3393_ (.Y(_0732_),
    .A(net50),
    .B(_0660_));
 sg13g2_a21oi_1 _3394_ (.A1(_0457_),
    .A2(_0679_),
    .Y(_0733_),
    .B1(_0732_));
 sg13g2_nor2_1 _3395_ (.A(_0640_),
    .B(_0644_),
    .Y(_0734_));
 sg13g2_a221oi_1 _3396_ (.B2(_0685_),
    .C1(_0734_),
    .B1(_0677_),
    .A1(_0727_),
    .Y(_0735_),
    .A2(_0457_));
 sg13g2_a221oi_1 _3397_ (.B2(_0733_),
    .C1(_0735_),
    .B1(_0731_),
    .A1(_0728_),
    .Y(_0736_),
    .A2(_0730_));
 sg13g2_buf_2 _3398_ (.A(_0736_),
    .X(_0737_));
 sg13g2_nand3_1 _3399_ (.B(_0443_),
    .C(_0451_),
    .A(_0423_),
    .Y(_0738_));
 sg13g2_a221oi_1 _3400_ (.B2(_0442_),
    .C1(_0738_),
    .B1(_0434_),
    .A1(_0424_),
    .Y(_0739_),
    .A2(_0429_));
 sg13g2_nand3_1 _3401_ (.B(_0443_),
    .C(_0451_),
    .A(_0448_),
    .Y(_0740_));
 sg13g2_a221oi_1 _3402_ (.B2(_0442_),
    .C1(_0740_),
    .B1(_0434_),
    .A1(_0424_),
    .Y(_0741_),
    .A2(_0429_));
 sg13g2_nand3_1 _3403_ (.B(_0423_),
    .C(_0451_),
    .A(_0448_),
    .Y(_0742_));
 sg13g2_nand2_1 _3404_ (.Y(_0743_),
    .A(_0453_),
    .B(_0742_));
 sg13g2_nor3_2 _3405_ (.A(_0739_),
    .B(_0741_),
    .C(_0743_),
    .Y(_0744_));
 sg13g2_inv_1 _3406_ (.Y(_0745_),
    .A(\gray_sobel0.sobel0.sobel.pix1_0[7] ));
 sg13g2_nand2_1 _3407_ (.Y(_0746_),
    .A(_0745_),
    .B(\gray_sobel0.sobel0.sobel.pix1_2[7] ));
 sg13g2_nor2_1 _3408_ (.A(_0745_),
    .B(\gray_sobel0.sobel0.sobel.pix1_2[7] ),
    .Y(_0747_));
 sg13g2_a21oi_2 _3409_ (.B1(_0747_),
    .Y(_0748_),
    .A2(_0746_),
    .A1(_0744_));
 sg13g2_inv_2 _3410_ (.Y(_0749_),
    .A(_0406_));
 sg13g2_buf_1 _3411_ (.A(\gray_sobel0.sobel0.sobel.pix0_2[7] ),
    .X(_0750_));
 sg13g2_inv_1 _3412_ (.Y(_0751_),
    .A(_0750_));
 sg13g2_nor3_2 _3413_ (.A(net87),
    .B(_0418_),
    .C(_0420_),
    .Y(_0752_));
 sg13g2_nor2_1 _3414_ (.A(net98),
    .B(_0362_),
    .Y(_0753_));
 sg13g2_a22oi_1 _3415_ (.Y(_0754_),
    .B1(_0396_),
    .B2(_0410_),
    .A2(net65),
    .A1(_0411_));
 sg13g2_buf_1 _3416_ (.A(\gray_sobel0.sobel0.sobel.pix0_0[7] ),
    .X(_0755_));
 sg13g2_a221oi_1 _3417_ (.B2(_0754_),
    .C1(net97),
    .B1(_0753_),
    .A1(net87),
    .Y(_0756_),
    .A2(_0420_));
 sg13g2_buf_1 _3418_ (.A(_0756_),
    .X(_0757_));
 sg13g2_or4_1 _3419_ (.A(_0749_),
    .B(net101),
    .C(_0752_),
    .D(_0757_),
    .X(_0758_));
 sg13g2_buf_1 _3420_ (.A(_0758_),
    .X(_0759_));
 sg13g2_nor2_1 _3421_ (.A(_0748_),
    .B(_0759_),
    .Y(_0760_));
 sg13g2_inv_1 _3422_ (.Y(_0761_),
    .A(_0760_));
 sg13g2_inv_1 _3423_ (.Y(_0762_),
    .A(_0404_));
 sg13g2_buf_1 _3424_ (.A(_0762_),
    .X(_0763_));
 sg13g2_nor2_1 _3425_ (.A(_0406_),
    .B(net74),
    .Y(_0764_));
 sg13g2_o21ai_1 _3426_ (.B1(_0764_),
    .Y(_0765_),
    .A1(_0752_),
    .A2(_0757_));
 sg13g2_a21oi_1 _3427_ (.A1(_0759_),
    .A2(_0765_),
    .Y(_0766_),
    .B1(_0748_));
 sg13g2_nand3_1 _3428_ (.B(_0759_),
    .C(_0765_),
    .A(_0748_),
    .Y(_0767_));
 sg13g2_nor2b_2 _3429_ (.A(_0766_),
    .B_N(_0767_),
    .Y(_0768_));
 sg13g2_nor3_1 _3430_ (.A(net101),
    .B(_0752_),
    .C(_0757_),
    .Y(_0769_));
 sg13g2_a21o_1 _3431_ (.A2(net65),
    .A1(_0411_),
    .B1(_0417_),
    .X(_0770_));
 sg13g2_a21o_1 _3432_ (.A2(_0394_),
    .A1(_0373_),
    .B1(_0419_),
    .X(_0771_));
 sg13g2_a21oi_1 _3433_ (.A1(_0770_),
    .A2(_0771_),
    .Y(_0772_),
    .B1(net98));
 sg13g2_nor2b_1 _3434_ (.A(_0747_),
    .B_N(_0746_),
    .Y(_0773_));
 sg13g2_xor2_1 _3435_ (.B(_0773_),
    .A(_0744_),
    .X(_0774_));
 sg13g2_a21oi_1 _3436_ (.A1(net97),
    .A2(_0772_),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_buf_1 _3437_ (.A(_0406_),
    .X(_0776_));
 sg13g2_o21ai_1 _3438_ (.B1(net86),
    .Y(_0777_),
    .A1(_0769_),
    .A2(_0775_));
 sg13g2_nand3_1 _3439_ (.B(_0770_),
    .C(_0771_),
    .A(net98),
    .Y(_0778_));
 sg13g2_nor3_1 _3440_ (.A(_0749_),
    .B(net97),
    .C(_0778_),
    .Y(_0779_));
 sg13g2_nor4_1 _3441_ (.A(net86),
    .B(_0752_),
    .C(_0757_),
    .D(_0774_),
    .Y(_0780_));
 sg13g2_o21ai_1 _3442_ (.B1(net101),
    .Y(_0781_),
    .A1(_0779_),
    .A2(_0780_));
 sg13g2_nor3_1 _3443_ (.A(_0406_),
    .B(net97),
    .C(net87),
    .Y(_0782_));
 sg13g2_and2_1 _3444_ (.A(_0421_),
    .B(_0782_),
    .X(_0783_));
 sg13g2_o21ai_1 _3445_ (.B1(net74),
    .Y(_0784_),
    .A1(_0775_),
    .A2(_0783_));
 sg13g2_nand3_1 _3446_ (.B(_0781_),
    .C(_0784_),
    .A(_0777_),
    .Y(_0785_));
 sg13g2_buf_1 _3447_ (.A(_0785_),
    .X(_0786_));
 sg13g2_nand3_1 _3448_ (.B(net97),
    .C(_0772_),
    .A(net86),
    .Y(_0787_));
 sg13g2_nor3_1 _3449_ (.A(_0406_),
    .B(net74),
    .C(net87),
    .Y(_0788_));
 sg13g2_o21ai_1 _3450_ (.B1(_0421_),
    .Y(_0789_),
    .A1(_0782_),
    .A2(_0788_));
 sg13g2_nor2b_1 _3451_ (.A(net101),
    .B_N(\gray_sobel0.sobel0.sobel.pix0_0[7] ),
    .Y(_0790_));
 sg13g2_inv_1 _3452_ (.Y(_0791_),
    .A(net97));
 sg13g2_nand2_1 _3453_ (.Y(_0792_),
    .A(net101),
    .B(_0791_));
 sg13g2_nor4_1 _3454_ (.A(net87),
    .B(_0792_),
    .C(_0418_),
    .D(_0420_),
    .Y(_0793_));
 sg13g2_a221oi_1 _3455_ (.B2(_0764_),
    .C1(_0793_),
    .B1(_0757_),
    .A1(_0790_),
    .Y(_0794_),
    .A2(_0772_));
 sg13g2_nand4_1 _3456_ (.B(_0787_),
    .C(_0789_),
    .A(_0759_),
    .Y(_0795_),
    .D(_0794_));
 sg13g2_xor2_1 _3457_ (.B(_0795_),
    .A(_0774_),
    .X(_0796_));
 sg13g2_buf_2 _3458_ (.A(_0796_),
    .X(_0797_));
 sg13g2_nand3_1 _3459_ (.B(_0402_),
    .C(_0455_),
    .A(_0399_),
    .Y(_0798_));
 sg13g2_a21oi_1 _3460_ (.A1(_0399_),
    .A2(_0402_),
    .Y(_0799_),
    .B1(_0455_));
 sg13g2_a21oi_1 _3461_ (.A1(_0422_),
    .A2(_0798_),
    .Y(_0800_),
    .B1(_0799_));
 sg13g2_buf_1 _3462_ (.A(_0800_),
    .X(_0801_));
 sg13g2_nor3_1 _3463_ (.A(_0786_),
    .B(_0797_),
    .C(net35),
    .Y(_0802_));
 sg13g2_o21ai_1 _3464_ (.B1(_0786_),
    .Y(_0803_),
    .A1(_0797_),
    .A2(net35));
 sg13g2_o21ai_1 _3465_ (.B1(_0803_),
    .Y(_0804_),
    .A1(_0768_),
    .A2(_0802_));
 sg13g2_nand3_1 _3466_ (.B(_0761_),
    .C(_0804_),
    .A(_0737_),
    .Y(_0805_));
 sg13g2_buf_2 _3467_ (.A(_0805_),
    .X(_0806_));
 sg13g2_nand3_1 _3468_ (.B(_0797_),
    .C(net35),
    .A(_0786_),
    .Y(_0807_));
 sg13g2_a21oi_1 _3469_ (.A1(_0797_),
    .A2(_0801_),
    .Y(_0808_),
    .B1(_0786_));
 sg13g2_a21oi_1 _3470_ (.A1(_0768_),
    .A2(_0807_),
    .Y(_0809_),
    .B1(_0808_));
 sg13g2_o21ai_1 _3471_ (.B1(_0748_),
    .Y(_0810_),
    .A1(_0752_),
    .A2(_0757_));
 sg13g2_nor3_2 _3472_ (.A(net86),
    .B(net74),
    .C(_0810_),
    .Y(_0811_));
 sg13g2_a21oi_1 _3473_ (.A1(_0761_),
    .A2(_0809_),
    .Y(_0812_),
    .B1(_0811_));
 sg13g2_buf_1 _3474_ (.A(_0812_),
    .X(_0813_));
 sg13g2_nand2_1 _3475_ (.Y(_0814_),
    .A(_0806_),
    .B(_0813_));
 sg13g2_buf_2 _3476_ (.A(_0814_),
    .X(_0815_));
 sg13g2_nor2b_1 _3477_ (.A(_0726_),
    .B_N(_0815_),
    .Y(_0816_));
 sg13g2_xnor2_1 _3478_ (.Y(_0817_),
    .A(_0797_),
    .B(net35));
 sg13g2_xnor2_1 _3479_ (.Y(_0818_),
    .A(_0737_),
    .B(_0817_));
 sg13g2_xnor2_1 _3480_ (.Y(_0819_),
    .A(_0816_),
    .B(_0818_));
 sg13g2_xnor2_1 _3481_ (.Y(_0820_),
    .A(_0729_),
    .B(_0688_));
 sg13g2_nor2_1 _3482_ (.A(net109),
    .B(_0416_),
    .Y(_0821_));
 sg13g2_nor2_1 _3483_ (.A(net107),
    .B(net106),
    .Y(_0822_));
 sg13g2_nand2_1 _3484_ (.Y(_0823_),
    .A(_0368_),
    .B(_0369_));
 sg13g2_o21ai_1 _3485_ (.B1(_0823_),
    .Y(_0824_),
    .A1(_0608_),
    .A2(_0822_));
 sg13g2_buf_1 _3486_ (.A(_0824_),
    .X(_0825_));
 sg13g2_and2_1 _3487_ (.A(net108),
    .B(_0825_),
    .X(_0826_));
 sg13g2_or2_1 _3488_ (.X(_0827_),
    .B(_0825_),
    .A(net108));
 sg13g2_nor2_1 _3489_ (.A(_0400_),
    .B(net109),
    .Y(_0828_));
 sg13g2_and2_1 _3490_ (.A(_0362_),
    .B(_0828_),
    .X(_0829_));
 sg13g2_or2_1 _3491_ (.X(_0830_),
    .B(_0369_),
    .A(_0368_));
 sg13g2_nand2_1 _3492_ (.Y(_0831_),
    .A(_0608_),
    .B(_0823_));
 sg13g2_nand2_1 _3493_ (.Y(_0832_),
    .A(net109),
    .B(_0416_));
 sg13g2_nand2_1 _3494_ (.Y(_0833_),
    .A(_0400_),
    .B(_0416_));
 sg13g2_a221oi_1 _3495_ (.B2(_0833_),
    .C1(net108),
    .B1(_0832_),
    .A1(_0830_),
    .Y(_0834_),
    .A2(_0831_));
 sg13g2_a221oi_1 _3496_ (.B2(_0829_),
    .C1(_0834_),
    .B1(_0827_),
    .A1(_0821_),
    .Y(_0835_),
    .A2(_0826_));
 sg13g2_nand2_1 _3497_ (.Y(_0836_),
    .A(net108),
    .B(_0825_));
 sg13g2_nand2_1 _3498_ (.Y(_0837_),
    .A(_0400_),
    .B(net109));
 sg13g2_nor2_1 _3499_ (.A(_0362_),
    .B(_0837_),
    .Y(_0838_));
 sg13g2_nor3_1 _3500_ (.A(net108),
    .B(_0825_),
    .C(_0837_),
    .Y(_0839_));
 sg13g2_a21oi_1 _3501_ (.A1(_0836_),
    .A2(_0838_),
    .Y(_0840_),
    .B1(_0839_));
 sg13g2_nor2_1 _3502_ (.A(_0400_),
    .B(_0416_),
    .Y(_0841_));
 sg13g2_o21ai_1 _3503_ (.B1(_0826_),
    .Y(_0842_),
    .A1(_0828_),
    .A2(_0841_));
 sg13g2_nand3_1 _3504_ (.B(_0840_),
    .C(_0842_),
    .A(_0835_),
    .Y(_0843_));
 sg13g2_xor2_1 _3505_ (.B(_0843_),
    .A(_0409_),
    .X(_0844_));
 sg13g2_buf_1 _3506_ (.A(\gray_sobel0.sobel0.sobel.pix2_1[5] ),
    .X(_0845_));
 sg13g2_nor2b_1 _3507_ (.A(\gray_sobel0.sobel0.sobel.pix0_1[5] ),
    .B_N(_0845_),
    .Y(_0846_));
 sg13g2_buf_1 _3508_ (.A(\gray_sobel0.sobel0.sobel.pix2_1[4] ),
    .X(_0847_));
 sg13g2_inv_1 _3509_ (.Y(_0848_),
    .A(_0847_));
 sg13g2_buf_1 _3510_ (.A(\gray_sobel0.sobel0.sobel.pix0_1[4] ),
    .X(_0849_));
 sg13g2_nor2_1 _3511_ (.A(_0848_),
    .B(_0849_),
    .Y(_0850_));
 sg13g2_nor2_1 _3512_ (.A(_0846_),
    .B(_0850_),
    .Y(_0851_));
 sg13g2_buf_2 _3513_ (.A(\gray_sobel0.sobel0.sobel.pix2_1[3] ),
    .X(_0852_));
 sg13g2_nor2b_1 _3514_ (.A(\gray_sobel0.sobel0.sobel.pix0_1[2] ),
    .B_N(\gray_sobel0.sobel0.sobel.pix2_1[2] ),
    .Y(_0853_));
 sg13g2_buf_1 _3515_ (.A(\gray_sobel0.sobel0.sobel.pix2_1[1] ),
    .X(_0854_));
 sg13g2_nor2b_1 _3516_ (.A(\gray_sobel0.sobel0.sobel.pix0_1[1] ),
    .B_N(_0854_),
    .Y(_0855_));
 sg13g2_nand2b_1 _3517_ (.Y(_0856_),
    .B(\gray_sobel0.sobel0.sobel.pix0_1[0] ),
    .A_N(\gray_sobel0.sobel0.sobel.pix2_1[0] ));
 sg13g2_nor3_2 _3518_ (.A(_0853_),
    .B(_0855_),
    .C(_0856_),
    .Y(_0857_));
 sg13g2_nand2b_1 _3519_ (.Y(_0858_),
    .B(\gray_sobel0.sobel0.sobel.pix0_1[1] ),
    .A_N(_0854_));
 sg13g2_nand2b_1 _3520_ (.Y(_0859_),
    .B(\gray_sobel0.sobel0.sobel.pix0_1[2] ),
    .A_N(\gray_sobel0.sobel0.sobel.pix2_1[2] ));
 sg13g2_o21ai_1 _3521_ (.B1(_0859_),
    .Y(_0860_),
    .A1(_0853_),
    .A2(_0858_));
 sg13g2_buf_1 _3522_ (.A(_0860_),
    .X(_0861_));
 sg13g2_buf_1 _3523_ (.A(\gray_sobel0.sobel0.sobel.pix0_1[3] ),
    .X(_0862_));
 sg13g2_o21ai_1 _3524_ (.B1(_0862_),
    .Y(_0863_),
    .A1(_0857_),
    .A2(_0861_));
 sg13g2_nor3_1 _3525_ (.A(_0862_),
    .B(_0857_),
    .C(_0861_),
    .Y(_0864_));
 sg13g2_a21oi_2 _3526_ (.B1(_0864_),
    .Y(_0865_),
    .A2(_0863_),
    .A1(_0852_));
 sg13g2_nand2b_1 _3527_ (.Y(_0866_),
    .B(_0849_),
    .A_N(_0847_));
 sg13g2_nand2b_1 _3528_ (.Y(_0867_),
    .B(\gray_sobel0.sobel0.sobel.pix0_1[5] ),
    .A_N(_0845_));
 sg13g2_a21oi_1 _3529_ (.A1(_0866_),
    .A2(_0867_),
    .Y(_0868_),
    .B1(_0846_));
 sg13g2_a21o_1 _3530_ (.A2(_0865_),
    .A1(_0851_),
    .B1(_0868_),
    .X(_0869_));
 sg13g2_buf_1 _3531_ (.A(_0869_),
    .X(_0870_));
 sg13g2_buf_1 _3532_ (.A(\gray_sobel0.sobel0.sobel.pix2_1[6] ),
    .X(_0871_));
 sg13g2_buf_1 _3533_ (.A(\gray_sobel0.sobel0.sobel.pix0_1[6] ),
    .X(_0872_));
 sg13g2_xor2_1 _3534_ (.B(_0872_),
    .A(_0871_),
    .X(_0873_));
 sg13g2_xnor2_1 _3535_ (.Y(_0874_),
    .A(_0870_),
    .B(_0873_));
 sg13g2_xnor2_1 _3536_ (.Y(_0875_),
    .A(_0844_),
    .B(_0874_));
 sg13g2_inv_1 _3537_ (.Y(_0876_),
    .A(_0852_));
 sg13g2_or2_1 _3538_ (.X(_0877_),
    .B(_0861_),
    .A(_0857_));
 sg13g2_a221oi_1 _3539_ (.B2(_0876_),
    .C1(_0877_),
    .B1(_0862_),
    .A1(_0848_),
    .Y(_0878_),
    .A2(_0849_));
 sg13g2_nand2b_1 _3540_ (.Y(_0879_),
    .B(_0852_),
    .A_N(_0862_));
 sg13g2_a21oi_1 _3541_ (.A1(_0848_),
    .A2(_0849_),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_nor3_2 _3542_ (.A(_0850_),
    .B(_0878_),
    .C(_0880_),
    .Y(_0881_));
 sg13g2_nor2b_1 _3543_ (.A(_0845_),
    .B_N(\gray_sobel0.sobel0.sobel.pix0_1[5] ),
    .Y(_0882_));
 sg13g2_nor2_1 _3544_ (.A(_0846_),
    .B(_0882_),
    .Y(_0883_));
 sg13g2_xor2_1 _3545_ (.B(_0883_),
    .A(_0881_),
    .X(_0884_));
 sg13g2_nor2_1 _3546_ (.A(_0365_),
    .B(_0366_),
    .Y(_0885_));
 sg13g2_nand2_1 _3547_ (.Y(_0886_),
    .A(_0365_),
    .B(_0366_));
 sg13g2_o21ai_1 _3548_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0557_),
    .A2(_0885_));
 sg13g2_xnor2_1 _3549_ (.Y(_0888_),
    .A(net88),
    .B(_0610_));
 sg13g2_nand2_1 _3550_ (.Y(_0889_),
    .A(net99),
    .B(_0888_));
 sg13g2_nor2_1 _3551_ (.A(net99),
    .B(_0888_),
    .Y(_0890_));
 sg13g2_a21oi_1 _3552_ (.A1(_0887_),
    .A2(_0889_),
    .Y(_0891_),
    .B1(_0890_));
 sg13g2_buf_1 _3553_ (.A(_0891_),
    .X(_0892_));
 sg13g2_inv_1 _3554_ (.Y(_0893_),
    .A(_0892_));
 sg13g2_xnor2_1 _3555_ (.Y(_0894_),
    .A(_0881_),
    .B(_0883_));
 sg13g2_nand2b_1 _3556_ (.Y(_0895_),
    .B(_0642_),
    .A_N(_0825_));
 sg13g2_nand3b_1 _3557_ (.B(_0831_),
    .C(_0830_),
    .Y(_0896_),
    .A_N(_0642_));
 sg13g2_nand2_2 _3558_ (.Y(_0897_),
    .A(_0895_),
    .B(_0896_));
 sg13g2_o21ai_1 _3559_ (.B1(_0897_),
    .Y(_0898_),
    .A1(_0894_),
    .A2(_0892_));
 sg13g2_o21ai_1 _3560_ (.B1(_0898_),
    .Y(_0899_),
    .A1(_0884_),
    .A2(_0893_));
 sg13g2_xor2_1 _3561_ (.B(_0899_),
    .A(_0875_),
    .X(_0900_));
 sg13g2_inv_1 _3562_ (.Y(_0901_),
    .A(_0900_));
 sg13g2_or2_1 _3563_ (.X(_0902_),
    .B(net104),
    .A(net103));
 sg13g2_and2_1 _3564_ (.A(net103),
    .B(net104),
    .X(_0903_));
 sg13g2_a21o_1 _3565_ (.A2(_0902_),
    .A1(_0538_),
    .B1(_0903_),
    .X(_0904_));
 sg13g2_and2_1 _3566_ (.A(_0579_),
    .B(_0904_),
    .X(_0905_));
 sg13g2_and2_1 _3567_ (.A(net102),
    .B(net105),
    .X(_0906_));
 sg13g2_nor2_1 _3568_ (.A(net102),
    .B(_0382_),
    .Y(_0907_));
 sg13g2_mux2_1 _3569_ (.A0(_0906_),
    .A1(_0907_),
    .S(_0626_),
    .X(_0908_));
 sg13g2_a22oi_1 _3570_ (.Y(_0909_),
    .B1(_0571_),
    .B2(_0561_),
    .A2(_0908_),
    .A1(_0526_));
 sg13g2_nor2_1 _3571_ (.A(net89),
    .B(_0906_),
    .Y(_0910_));
 sg13g2_nor2_1 _3572_ (.A(_0907_),
    .B(_0910_),
    .Y(_0911_));
 sg13g2_nand2_1 _3573_ (.Y(_0912_),
    .A(net89),
    .B(net102));
 sg13g2_mux2_1 _3574_ (.A0(_0911_),
    .A1(_0912_),
    .S(_0561_),
    .X(_0913_));
 sg13g2_or3_1 _3575_ (.A(_0579_),
    .B(_0904_),
    .C(_0913_),
    .X(_0914_));
 sg13g2_o21ai_1 _3576_ (.B1(_0914_),
    .Y(_0915_),
    .A1(_0905_),
    .A2(_0909_));
 sg13g2_buf_1 _3577_ (.A(_0915_),
    .X(_0916_));
 sg13g2_nor2b_1 _3578_ (.A(_0487_),
    .B_N(net105),
    .Y(_0917_));
 sg13g2_a22oi_1 _3579_ (.Y(_0918_),
    .B1(_0917_),
    .B2(_0902_),
    .A2(_0903_),
    .A1(net105));
 sg13g2_nor2_1 _3580_ (.A(_0912_),
    .B(_0918_),
    .Y(_0919_));
 sg13g2_nor2_1 _3581_ (.A(net103),
    .B(net104),
    .Y(_0920_));
 sg13g2_a21oi_1 _3582_ (.A1(net103),
    .A2(net104),
    .Y(_0921_),
    .B1(net105));
 sg13g2_o21ai_1 _3583_ (.B1(_0921_),
    .Y(_0922_),
    .A1(_0487_),
    .A2(_0920_));
 sg13g2_buf_1 _3584_ (.A(_0922_),
    .X(_0923_));
 sg13g2_nor3_1 _3585_ (.A(net89),
    .B(net102),
    .C(_0923_),
    .Y(_0924_));
 sg13g2_and4_1 _3586_ (.A(_0579_),
    .B(net89),
    .C(net102),
    .D(_0923_),
    .X(_0925_));
 sg13g2_nor3_1 _3587_ (.A(_0579_),
    .B(net102),
    .C(_0923_),
    .Y(_0926_));
 sg13g2_nor4_2 _3588_ (.A(_0919_),
    .B(_0924_),
    .C(_0925_),
    .Y(_0927_),
    .D(_0926_));
 sg13g2_nand2_1 _3589_ (.Y(_0928_),
    .A(_0525_),
    .B(_0526_));
 sg13g2_nor2_1 _3590_ (.A(_0923_),
    .B(_0928_),
    .Y(_0929_));
 sg13g2_nor2_1 _3591_ (.A(net102),
    .B(_0928_),
    .Y(_0930_));
 sg13g2_and2_1 _3592_ (.A(_0918_),
    .B(_0930_),
    .X(_0931_));
 sg13g2_nand2_1 _3593_ (.Y(_0932_),
    .A(_0579_),
    .B(net89));
 sg13g2_nand2_1 _3594_ (.Y(_0933_),
    .A(_0579_),
    .B(net102));
 sg13g2_a21oi_1 _3595_ (.A1(_0932_),
    .A2(_0933_),
    .Y(_0934_),
    .B1(_0918_));
 sg13g2_nor3_2 _3596_ (.A(_0929_),
    .B(_0931_),
    .C(_0934_),
    .Y(_0935_));
 sg13g2_and2_1 _3597_ (.A(_0927_),
    .B(_0935_),
    .X(_0936_));
 sg13g2_xnor2_1 _3598_ (.Y(_0937_),
    .A(_0561_),
    .B(_0936_));
 sg13g2_nand2_1 _3599_ (.Y(_0938_),
    .A(_0375_),
    .B(_0374_));
 sg13g2_xnor2_1 _3600_ (.Y(_0939_),
    .A(_0487_),
    .B(net75));
 sg13g2_nor2_1 _3601_ (.A(_0938_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_a21oi_1 _3602_ (.A1(_0938_),
    .A2(_0939_),
    .Y(_0941_),
    .B1(\gray_sobel0.sobel0.sobel.pix2_0[2] ));
 sg13g2_xnor2_1 _3603_ (.Y(_0942_),
    .A(_0904_),
    .B(_0528_));
 sg13g2_o21ai_1 _3604_ (.B1(_0942_),
    .Y(_0943_),
    .A1(_0940_),
    .A2(_0941_));
 sg13g2_a21oi_1 _3605_ (.A1(_0856_),
    .A2(_0858_),
    .Y(_0944_),
    .B1(_0855_));
 sg13g2_nor2b_1 _3606_ (.A(_0853_),
    .B_N(_0859_),
    .Y(_0945_));
 sg13g2_xnor2_1 _3607_ (.Y(_0946_),
    .A(_0944_),
    .B(_0945_));
 sg13g2_nor3_1 _3608_ (.A(_0940_),
    .B(_0941_),
    .C(_0942_),
    .Y(_0947_));
 sg13g2_a21oi_2 _3609_ (.B1(_0947_),
    .Y(_0948_),
    .A2(_0946_),
    .A1(_0943_));
 sg13g2_inv_2 _3610_ (.Y(_0949_),
    .A(_0948_));
 sg13g2_nor2_1 _3611_ (.A(_0467_),
    .B(_0464_),
    .Y(_0950_));
 sg13g2_nand2b_1 _3612_ (.Y(_0951_),
    .B(_0377_),
    .A_N(net100));
 sg13g2_inv_1 _3613_ (.Y(_0952_),
    .A(\gray_sobel0.sobel0.sobel.pix0_2[0] ));
 sg13g2_nor2b_1 _3614_ (.A(_0377_),
    .B_N(_0458_),
    .Y(_0953_));
 sg13g2_a221oi_1 _3615_ (.B2(_0952_),
    .C1(_0953_),
    .B1(_0951_),
    .A1(_0467_),
    .Y(_0954_),
    .A2(_0464_));
 sg13g2_nor2_1 _3616_ (.A(_0950_),
    .B(_0954_),
    .Y(_0955_));
 sg13g2_xnor2_1 _3617_ (.Y(_0956_),
    .A(_0938_),
    .B(_0488_));
 sg13g2_xnor2_1 _3618_ (.Y(_0957_),
    .A(_0490_),
    .B(_0956_));
 sg13g2_nor2_1 _3619_ (.A(_0955_),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_xor2_1 _3620_ (.B(\gray_sobel0.sobel0.sobel.pix0_1[1] ),
    .A(_0854_),
    .X(_0959_));
 sg13g2_xnor2_1 _3621_ (.Y(_0960_),
    .A(_0856_),
    .B(_0959_));
 sg13g2_a21o_1 _3622_ (.A2(_0957_),
    .A1(_0955_),
    .B1(_0960_),
    .X(_0961_));
 sg13g2_nand2b_1 _3623_ (.Y(_0962_),
    .B(_0961_),
    .A_N(_0958_));
 sg13g2_nor2_1 _3624_ (.A(_0940_),
    .B(_0941_),
    .Y(_0963_));
 sg13g2_xnor2_1 _3625_ (.Y(_0964_),
    .A(_0942_),
    .B(_0946_));
 sg13g2_xnor2_1 _3626_ (.Y(_0965_),
    .A(_0963_),
    .B(_0964_));
 sg13g2_buf_2 _3627_ (.A(_0965_),
    .X(_0966_));
 sg13g2_nor2_1 _3628_ (.A(_0962_),
    .B(_0966_),
    .Y(_0967_));
 sg13g2_a21oi_1 _3629_ (.A1(_0962_),
    .A2(_0966_),
    .Y(_0968_),
    .B1(_0948_));
 sg13g2_xor2_1 _3630_ (.B(\gray_sobel0.sobel0.sobel.pix0_1[0] ),
    .A(\gray_sobel0.sobel0.sobel.pix2_1[0] ),
    .X(_0969_));
 sg13g2_a21oi_1 _3631_ (.A1(_0952_),
    .A2(_0951_),
    .Y(_0970_),
    .B1(_0953_));
 sg13g2_xnor2_1 _3632_ (.Y(_0971_),
    .A(_0508_),
    .B(_0464_));
 sg13g2_xnor2_1 _3633_ (.Y(_0972_),
    .A(_0970_),
    .B(_0971_));
 sg13g2_and2_1 _3634_ (.A(_0969_),
    .B(_0972_),
    .X(_0973_));
 sg13g2_buf_2 _3635_ (.A(_0973_),
    .X(_0974_));
 sg13g2_o21ai_1 _3636_ (.B1(_0960_),
    .Y(_0975_),
    .A1(_0950_),
    .A2(_0954_));
 sg13g2_or3_1 _3637_ (.A(_0950_),
    .B(_0954_),
    .C(_0960_),
    .X(_0976_));
 sg13g2_a21o_1 _3638_ (.A2(_0976_),
    .A1(_0975_),
    .B1(_0957_),
    .X(_0977_));
 sg13g2_nand3_1 _3639_ (.B(_0975_),
    .C(_0976_),
    .A(_0957_),
    .Y(_0978_));
 sg13g2_nand2_1 _3640_ (.Y(_0979_),
    .A(net90),
    .B(_0703_));
 sg13g2_nand3_1 _3641_ (.B(_0978_),
    .C(_0979_),
    .A(_0977_),
    .Y(_0980_));
 sg13g2_a21o_1 _3642_ (.A2(_0702_),
    .A1(_0481_),
    .B1(_0969_),
    .X(_0981_));
 sg13g2_o21ai_1 _3643_ (.B1(net90),
    .Y(_0982_),
    .A1(_0972_),
    .A2(_0981_));
 sg13g2_o21ai_1 _3644_ (.B1(_0703_),
    .Y(_0983_),
    .A1(_0969_),
    .A2(_0972_));
 sg13g2_a22oi_1 _3645_ (.Y(_0984_),
    .B1(_0982_),
    .B2(_0983_),
    .A2(_0978_),
    .A1(_0977_));
 sg13g2_a21o_1 _3646_ (.A2(_0980_),
    .A1(_0974_),
    .B1(_0984_),
    .X(_0985_));
 sg13g2_buf_8 _3647_ (.A(_0985_),
    .X(_0986_));
 sg13g2_xor2_1 _3648_ (.B(_0862_),
    .A(_0852_),
    .X(_0987_));
 sg13g2_or3_1 _3649_ (.A(_0857_),
    .B(_0861_),
    .C(_0987_),
    .X(_0988_));
 sg13g2_buf_1 _3650_ (.A(_0988_),
    .X(_0989_));
 sg13g2_o21ai_1 _3651_ (.B1(_0987_),
    .Y(_0990_),
    .A1(_0857_),
    .A2(_0861_));
 sg13g2_buf_1 _3652_ (.A(_0990_),
    .X(_0991_));
 sg13g2_and2_1 _3653_ (.A(_0989_),
    .B(_0991_),
    .X(_0992_));
 sg13g2_buf_2 _3654_ (.A(_0992_),
    .X(_0993_));
 sg13g2_a221oi_1 _3655_ (.B2(_0986_),
    .C1(_0993_),
    .B1(_0968_),
    .A1(_0949_),
    .Y(_0994_),
    .A2(_0967_));
 sg13g2_nand3b_1 _3656_ (.B(_0937_),
    .C(_0994_),
    .Y(_0995_),
    .A_N(net49));
 sg13g2_xor2_1 _3657_ (.B(_0849_),
    .A(_0847_),
    .X(_0996_));
 sg13g2_xnor2_1 _3658_ (.Y(_0997_),
    .A(_0865_),
    .B(_0996_));
 sg13g2_xor2_1 _3659_ (.B(_0633_),
    .A(_0887_),
    .X(_0998_));
 sg13g2_nor2_1 _3660_ (.A(_0555_),
    .B(_0559_),
    .Y(_0999_));
 sg13g2_nand2_1 _3661_ (.Y(_1000_),
    .A(_0555_),
    .B(_0559_));
 sg13g2_o21ai_1 _3662_ (.B1(_1000_),
    .Y(_1001_),
    .A1(_0911_),
    .A2(_0999_));
 sg13g2_xor2_1 _3663_ (.B(_1001_),
    .A(_0998_),
    .X(_1002_));
 sg13g2_xor2_1 _3664_ (.B(_1002_),
    .A(_0997_),
    .X(_1003_));
 sg13g2_buf_2 _3665_ (.A(_1003_),
    .X(_1004_));
 sg13g2_or2_1 _3666_ (.X(_1005_),
    .B(_0946_),
    .A(_0947_));
 sg13g2_nand2_1 _3667_ (.Y(_1006_),
    .A(_0962_),
    .B(_0966_));
 sg13g2_a221oi_1 _3668_ (.B2(_0986_),
    .C1(_0967_),
    .B1(_1006_),
    .A1(_0943_),
    .Y(_1007_),
    .A2(_1005_));
 sg13g2_buf_1 _3669_ (.A(_1007_),
    .X(_1008_));
 sg13g2_xnor2_1 _3670_ (.Y(_1009_),
    .A(_0626_),
    .B(_0936_));
 sg13g2_buf_2 _3671_ (.A(_1009_),
    .X(_1010_));
 sg13g2_a21oi_1 _3672_ (.A1(_0993_),
    .A2(_1010_),
    .Y(_1011_),
    .B1(net49));
 sg13g2_o21ai_1 _3673_ (.B1(_1011_),
    .Y(_1012_),
    .A1(_1004_),
    .A2(_1008_));
 sg13g2_nand3_1 _3674_ (.B(_0989_),
    .C(_0991_),
    .A(_0626_),
    .Y(_1013_));
 sg13g2_a21o_1 _3675_ (.A2(_0935_),
    .A1(_0927_),
    .B1(_1013_),
    .X(_1014_));
 sg13g2_nand4_1 _3676_ (.B(_0993_),
    .C(_0927_),
    .A(_0561_),
    .Y(_1015_),
    .D(_0935_));
 sg13g2_a21o_1 _3677_ (.A2(_0991_),
    .A1(_0989_),
    .B1(_0626_),
    .X(_1016_));
 sg13g2_a21o_1 _3678_ (.A2(_0935_),
    .A1(_0927_),
    .B1(_1016_),
    .X(_1017_));
 sg13g2_nand2_1 _3679_ (.Y(_1018_),
    .A(_0989_),
    .B(_0991_));
 sg13g2_nand4_1 _3680_ (.B(_1018_),
    .C(_0927_),
    .A(_0626_),
    .Y(_1019_),
    .D(_0935_));
 sg13g2_nand4_1 _3681_ (.B(_1015_),
    .C(_1017_),
    .A(_1014_),
    .Y(_1020_),
    .D(_1019_));
 sg13g2_buf_1 _3682_ (.A(_1020_),
    .X(_1021_));
 sg13g2_nor2_1 _3683_ (.A(_0949_),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_a221oi_1 _3684_ (.B2(_0949_),
    .C1(_0967_),
    .B1(_1021_),
    .A1(_1006_),
    .Y(_1023_),
    .A2(_0986_));
 sg13g2_o21ai_1 _3685_ (.B1(_1004_),
    .Y(_1024_),
    .A1(_1022_),
    .A2(_1023_));
 sg13g2_and3_1 _3686_ (.X(_1025_),
    .A(_0995_),
    .B(_1012_),
    .C(_1024_));
 sg13g2_buf_8 _3687_ (.A(_1025_),
    .X(_1026_));
 sg13g2_nand2_1 _3688_ (.Y(_1027_),
    .A(_0998_),
    .B(_1001_));
 sg13g2_nor2_1 _3689_ (.A(_0998_),
    .B(_1001_),
    .Y(_1028_));
 sg13g2_a21o_1 _3690_ (.A2(_1027_),
    .A1(_0997_),
    .B1(_1028_),
    .X(_1029_));
 sg13g2_buf_2 _3691_ (.A(_1029_),
    .X(_1030_));
 sg13g2_xor2_1 _3692_ (.B(_0892_),
    .A(_0897_),
    .X(_1031_));
 sg13g2_xnor2_1 _3693_ (.Y(_1032_),
    .A(_0894_),
    .B(_1031_));
 sg13g2_or2_1 _3694_ (.X(_1033_),
    .B(_1032_),
    .A(_1030_));
 sg13g2_inv_1 _3695_ (.Y(_1034_),
    .A(_1033_));
 sg13g2_nand2_1 _3696_ (.Y(_1035_),
    .A(_1030_),
    .B(_1032_));
 sg13g2_o21ai_1 _3697_ (.B1(_1035_),
    .Y(_1036_),
    .A1(_1026_),
    .A2(_1034_));
 sg13g2_buf_1 _3698_ (.A(_1036_),
    .X(_1037_));
 sg13g2_nor2b_1 _3699_ (.A(_0958_),
    .B_N(_0961_),
    .Y(_1038_));
 sg13g2_buf_2 _3700_ (.A(_1038_),
    .X(_1039_));
 sg13g2_xor2_1 _3701_ (.B(_0964_),
    .A(_0963_),
    .X(_1040_));
 sg13g2_a21oi_1 _3702_ (.A1(_0974_),
    .A2(_0980_),
    .Y(_1041_),
    .B1(_0984_));
 sg13g2_xnor2_1 _3703_ (.Y(_1042_),
    .A(_1040_),
    .B(_1041_));
 sg13g2_nor2_1 _3704_ (.A(_1039_),
    .B(_0966_),
    .Y(_1043_));
 sg13g2_xnor2_1 _3705_ (.Y(_1044_),
    .A(_0949_),
    .B(_1021_));
 sg13g2_a221oi_1 _3706_ (.B2(_0986_),
    .C1(_1044_),
    .B1(_1043_),
    .A1(_1039_),
    .Y(_1045_),
    .A2(_1042_));
 sg13g2_nor2_1 _3707_ (.A(_1039_),
    .B(_1040_),
    .Y(_1046_));
 sg13g2_nand2_1 _3708_ (.Y(_1047_),
    .A(_1046_),
    .B(_1041_));
 sg13g2_and2_1 _3709_ (.A(_0977_),
    .B(_0978_),
    .X(_1048_));
 sg13g2_buf_1 _3710_ (.A(_1048_),
    .X(_1049_));
 sg13g2_nand2_1 _3711_ (.Y(_1050_),
    .A(net90),
    .B(net68));
 sg13g2_nor2_1 _3712_ (.A(net76),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_nor2_1 _3713_ (.A(_0969_),
    .B(_0972_),
    .Y(_1052_));
 sg13g2_nor3_1 _3714_ (.A(net91),
    .B(_0506_),
    .C(net68),
    .Y(_1053_));
 sg13g2_a22oi_1 _3715_ (.Y(_1054_),
    .B1(_1053_),
    .B2(_0974_),
    .A2(_1052_),
    .A1(_1051_));
 sg13g2_xor2_1 _3716_ (.B(_0972_),
    .A(_0969_),
    .X(_1055_));
 sg13g2_nand2b_1 _3717_ (.Y(_1056_),
    .B(net90),
    .A_N(net68));
 sg13g2_inv_1 _3718_ (.Y(_1057_),
    .A(net90));
 sg13g2_nand3_1 _3719_ (.B(_1057_),
    .C(net68),
    .A(_0482_),
    .Y(_1058_));
 sg13g2_o21ai_1 _3720_ (.B1(_1058_),
    .Y(_1059_),
    .A1(net91),
    .A2(_1056_));
 sg13g2_nand2_1 _3721_ (.Y(_1060_),
    .A(_1055_),
    .B(_1059_));
 sg13g2_nand2_1 _3722_ (.Y(_1061_),
    .A(_1054_),
    .B(_1060_));
 sg13g2_a22oi_1 _3723_ (.Y(_1062_),
    .B1(_1052_),
    .B2(_1053_),
    .A2(_1051_),
    .A1(_0974_));
 sg13g2_nand2_1 _3724_ (.Y(_1063_),
    .A(_1049_),
    .B(_1062_));
 sg13g2_o21ai_1 _3725_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_1049_),
    .A2(_1061_));
 sg13g2_buf_1 _3726_ (.A(_1064_),
    .X(_1065_));
 sg13g2_a21oi_1 _3727_ (.A1(_1044_),
    .A2(_1047_),
    .Y(_1066_),
    .B1(_1065_));
 sg13g2_nand2b_1 _3728_ (.Y(_1067_),
    .B(_1066_),
    .A_N(_1045_));
 sg13g2_a221oi_1 _3729_ (.B2(_0980_),
    .C1(_0984_),
    .B1(_0974_),
    .A1(_1039_),
    .Y(_1068_),
    .A2(_1040_));
 sg13g2_o21ai_1 _3730_ (.B1(_0948_),
    .Y(_1069_),
    .A1(_1046_),
    .A2(_1068_));
 sg13g2_or4_1 _3731_ (.A(_0916_),
    .B(_1004_),
    .C(_1069_),
    .D(_1010_),
    .X(_1070_));
 sg13g2_nand4_1 _3732_ (.B(_1018_),
    .C(_1004_),
    .A(net49),
    .Y(_1071_),
    .D(_0937_));
 sg13g2_or4_1 _3733_ (.A(_0916_),
    .B(_0993_),
    .C(_1004_),
    .D(_1010_),
    .X(_1072_));
 sg13g2_nor3_2 _3734_ (.A(_0948_),
    .B(_1046_),
    .C(_1068_),
    .Y(_1073_));
 sg13g2_a21o_1 _3735_ (.A2(_1072_),
    .A1(_1071_),
    .B1(_1073_),
    .X(_1074_));
 sg13g2_xnor2_1 _3736_ (.Y(_1075_),
    .A(_0997_),
    .B(_1002_));
 sg13g2_nand3_1 _3737_ (.B(_1075_),
    .C(_1073_),
    .A(net49),
    .Y(_1076_));
 sg13g2_nand3_1 _3738_ (.B(_1004_),
    .C(_1010_),
    .A(_0993_),
    .Y(_1077_));
 sg13g2_nand3_1 _3739_ (.B(_1075_),
    .C(_1010_),
    .A(_0993_),
    .Y(_1078_));
 sg13g2_mux2_1 _3740_ (.A0(_1077_),
    .A1(_1078_),
    .S(_1073_),
    .X(_1079_));
 sg13g2_nand4_1 _3741_ (.B(_1074_),
    .C(_1076_),
    .A(_1070_),
    .Y(_1080_),
    .D(_1079_));
 sg13g2_buf_1 _3742_ (.A(_1080_),
    .X(_1081_));
 sg13g2_nor3_1 _3743_ (.A(net49),
    .B(_1075_),
    .C(_1010_),
    .Y(_1082_));
 sg13g2_and4_1 _3744_ (.A(net49),
    .B(_0993_),
    .C(_1075_),
    .D(_0937_),
    .X(_1083_));
 sg13g2_a22oi_1 _3745_ (.Y(_1084_),
    .B1(_1083_),
    .B2(_1069_),
    .A2(_1082_),
    .A1(_1073_));
 sg13g2_nor4_1 _3746_ (.A(net49),
    .B(_1018_),
    .C(_1075_),
    .D(_1010_),
    .Y(_1085_));
 sg13g2_nand2_1 _3747_ (.Y(_1086_),
    .A(_1069_),
    .B(_1085_));
 sg13g2_nand2_1 _3748_ (.Y(_1087_),
    .A(_1017_),
    .B(_1019_));
 sg13g2_nand2_1 _3749_ (.Y(_1088_),
    .A(_1004_),
    .B(_1087_));
 sg13g2_nand2_1 _3750_ (.Y(_1089_),
    .A(net49),
    .B(_1004_));
 sg13g2_mux2_1 _3751_ (.A0(_1088_),
    .A1(_1089_),
    .S(_1008_),
    .X(_1090_));
 sg13g2_nand3_1 _3752_ (.B(_1008_),
    .C(_1087_),
    .A(_1075_),
    .Y(_1091_));
 sg13g2_nand4_1 _3753_ (.B(_1086_),
    .C(_1090_),
    .A(_1084_),
    .Y(_1092_),
    .D(_1091_));
 sg13g2_buf_1 _3754_ (.A(_1092_),
    .X(_1093_));
 sg13g2_inv_1 _3755_ (.Y(_1094_),
    .A(_1032_));
 sg13g2_nor4_1 _3756_ (.A(_1067_),
    .B(_1081_),
    .C(_1093_),
    .D(_1094_),
    .Y(_1095_));
 sg13g2_a21oi_2 _3757_ (.B1(_1028_),
    .Y(_1096_),
    .A2(_1027_),
    .A1(_0997_));
 sg13g2_nor4_1 _3758_ (.A(_1096_),
    .B(_1067_),
    .C(_1081_),
    .D(_1093_),
    .Y(_1097_));
 sg13g2_nor3_1 _3759_ (.A(_1037_),
    .B(_1095_),
    .C(_1097_),
    .Y(_1098_));
 sg13g2_nand2b_1 _3760_ (.Y(_1099_),
    .B(\gray_sobel0.sobel0.sobel.pix2_1[7] ),
    .A_N(\gray_sobel0.sobel0.sobel.pix0_1[7] ));
 sg13g2_buf_1 _3761_ (.A(_1099_),
    .X(_1100_));
 sg13g2_nand2_1 _3762_ (.Y(_1101_),
    .A(_0872_),
    .B(_0870_));
 sg13g2_inv_1 _3763_ (.Y(_1102_),
    .A(_0871_));
 sg13g2_o21ai_1 _3764_ (.B1(_1102_),
    .Y(_1103_),
    .A1(_0872_),
    .A2(_0870_));
 sg13g2_and2_1 _3765_ (.A(_1101_),
    .B(_1103_),
    .X(_1104_));
 sg13g2_nor2b_1 _3766_ (.A(\gray_sobel0.sobel0.sobel.pix2_1[7] ),
    .B_N(\gray_sobel0.sobel0.sobel.pix0_1[7] ),
    .Y(_1105_));
 sg13g2_a21oi_1 _3767_ (.A1(_1100_),
    .A2(_1104_),
    .Y(_1106_),
    .B1(_1105_));
 sg13g2_nand3_1 _3768_ (.B(net98),
    .C(_0790_),
    .A(_0749_),
    .Y(_1107_));
 sg13g2_inv_1 _3769_ (.Y(_1108_),
    .A(_1107_));
 sg13g2_nand2b_1 _3770_ (.Y(_1109_),
    .B(_1108_),
    .A_N(_1106_));
 sg13g2_inv_1 _3771_ (.Y(_1110_),
    .A(\gray_sobel0.sobel0.sobel.pix2_1[7] ));
 sg13g2_nor4_1 _3772_ (.A(_0749_),
    .B(_0762_),
    .C(net97),
    .D(net98),
    .Y(_1111_));
 sg13g2_or2_1 _3773_ (.X(_1112_),
    .B(_1111_),
    .A(_1108_));
 sg13g2_inv_1 _3774_ (.Y(_1113_),
    .A(_1112_));
 sg13g2_a221oi_1 _3775_ (.B2(_1103_),
    .C1(_1113_),
    .B1(_1101_),
    .A1(_1110_),
    .Y(_1114_),
    .A2(\gray_sobel0.sobel0.sobel.pix0_1[7] ));
 sg13g2_and4_1 _3776_ (.A(_1100_),
    .B(_1101_),
    .C(_1103_),
    .D(_1113_),
    .X(_1115_));
 sg13g2_nand2_1 _3777_ (.Y(_1116_),
    .A(_1105_),
    .B(_1113_));
 sg13g2_o21ai_1 _3778_ (.B1(_1116_),
    .Y(_1117_),
    .A1(_1100_),
    .A2(_1113_));
 sg13g2_nor3_2 _3779_ (.A(_1114_),
    .B(_1115_),
    .C(_1117_),
    .Y(_1118_));
 sg13g2_nand2b_1 _3780_ (.Y(_1119_),
    .B(_1100_),
    .A_N(_1105_));
 sg13g2_nand2b_1 _3781_ (.Y(_1120_),
    .B(_0871_),
    .A_N(_0872_));
 sg13g2_nand4_1 _3782_ (.B(_0851_),
    .C(_1120_),
    .A(_1119_),
    .Y(_1121_),
    .D(_0865_));
 sg13g2_a21o_1 _3783_ (.A2(_0863_),
    .A1(_0852_),
    .B1(_0864_),
    .X(_1122_));
 sg13g2_nor2b_1 _3784_ (.A(_0871_),
    .B_N(_0872_),
    .Y(_1123_));
 sg13g2_nor2_1 _3785_ (.A(_1119_),
    .B(_1123_),
    .Y(_1124_));
 sg13g2_and3_1 _3786_ (.X(_1125_),
    .A(_0866_),
    .B(_0867_),
    .C(_1124_));
 sg13g2_nor2_1 _3787_ (.A(_0882_),
    .B(_0851_),
    .Y(_1126_));
 sg13g2_nor2b_1 _3788_ (.A(_1105_),
    .B_N(_1100_),
    .Y(_1127_));
 sg13g2_nand2_1 _3789_ (.Y(_1128_),
    .A(_0868_),
    .B(_1120_));
 sg13g2_nor2_1 _3790_ (.A(_1127_),
    .B(_1123_),
    .Y(_1129_));
 sg13g2_a22oi_1 _3791_ (.Y(_1130_),
    .B1(_1128_),
    .B2(_1129_),
    .A2(_1120_),
    .A1(_1127_));
 sg13g2_a221oi_1 _3792_ (.B2(_1124_),
    .C1(_1130_),
    .B1(_1126_),
    .A1(_1122_),
    .Y(_1131_),
    .A2(_1125_));
 sg13g2_nand2_1 _3793_ (.Y(_1132_),
    .A(_1121_),
    .B(_1131_));
 sg13g2_inv_1 _3794_ (.Y(_1133_),
    .A(net109));
 sg13g2_or2_1 _3795_ (.X(_1134_),
    .B(_0363_),
    .A(_0362_));
 sg13g2_and2_1 _3796_ (.A(_0362_),
    .B(\gray_sobel0.sobel0.sobel.pix0_2[6] ),
    .X(_1135_));
 sg13g2_buf_1 _3797_ (.A(_1135_),
    .X(_1136_));
 sg13g2_a21o_1 _3798_ (.A2(_1134_),
    .A1(_1133_),
    .B1(_1136_),
    .X(_1137_));
 sg13g2_nor2_1 _3799_ (.A(net87),
    .B(_1137_),
    .Y(_1138_));
 sg13g2_a21oi_2 _3800_ (.B1(_1136_),
    .Y(_1139_),
    .A2(_1134_),
    .A1(_1133_));
 sg13g2_nor2_1 _3801_ (.A(net98),
    .B(_1139_),
    .Y(_1140_));
 sg13g2_a21oi_1 _3802_ (.A1(net98),
    .A2(_1139_),
    .Y(_1141_),
    .B1(_0755_));
 sg13g2_nor2_1 _3803_ (.A(_1140_),
    .B(_1141_),
    .Y(_1142_));
 sg13g2_a221oi_1 _3804_ (.B2(net74),
    .C1(_0406_),
    .B1(_1142_),
    .A1(_0755_),
    .Y(_1143_),
    .A2(_1138_));
 sg13g2_or2_1 _3805_ (.X(_1144_),
    .B(_1141_),
    .A(_1140_));
 sg13g2_a221oi_1 _3806_ (.B2(net101),
    .C1(_0749_),
    .B1(_1144_),
    .A1(_0791_),
    .Y(_1145_),
    .A2(_1140_));
 sg13g2_nor3_1 _3807_ (.A(net98),
    .B(_1139_),
    .C(_0792_),
    .Y(_1146_));
 sg13g2_a21oi_1 _3808_ (.A1(_0790_),
    .A2(_1138_),
    .Y(_1147_),
    .B1(_1146_));
 sg13g2_o21ai_1 _3809_ (.B1(_1147_),
    .Y(_1148_),
    .A1(_1143_),
    .A2(_1145_));
 sg13g2_xor2_1 _3810_ (.B(_1148_),
    .A(_1132_),
    .X(_1149_));
 sg13g2_nand2_1 _3811_ (.Y(_1150_),
    .A(_0409_),
    .B(_0821_));
 sg13g2_o21ai_1 _3812_ (.B1(_1150_),
    .Y(_1151_),
    .A1(_1137_),
    .A2(_0409_));
 sg13g2_nor2_1 _3813_ (.A(_0401_),
    .B(_0825_),
    .Y(_1152_));
 sg13g2_nor2_1 _3814_ (.A(_0362_),
    .B(net108),
    .Y(_1153_));
 sg13g2_mux2_1 _3815_ (.A0(_1153_),
    .A1(_1136_),
    .S(_0409_),
    .X(_1154_));
 sg13g2_and2_1 _3816_ (.A(_1133_),
    .B(_0364_),
    .X(_1155_));
 sg13g2_a22oi_1 _3817_ (.Y(_1156_),
    .B1(_1155_),
    .B2(_0409_),
    .A2(_1154_),
    .A1(_0361_));
 sg13g2_a21oi_1 _3818_ (.A1(_0401_),
    .A2(_0825_),
    .Y(_1157_),
    .B1(_1156_));
 sg13g2_a21oi_1 _3819_ (.A1(_1151_),
    .A2(_1152_),
    .Y(_1158_),
    .B1(_1157_));
 sg13g2_o21ai_1 _3820_ (.B1(_1158_),
    .Y(_1159_),
    .A1(_0844_),
    .A2(_0874_));
 sg13g2_buf_1 _3821_ (.A(_1159_),
    .X(_1160_));
 sg13g2_nor2_1 _3822_ (.A(_1149_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_nor4_1 _3823_ (.A(_0749_),
    .B(_0763_),
    .C(net87),
    .D(_1139_),
    .Y(_1162_));
 sg13g2_nand2_1 _3824_ (.Y(_1163_),
    .A(_0749_),
    .B(_0751_));
 sg13g2_a21oi_1 _3825_ (.A1(_1121_),
    .A2(_1131_),
    .Y(_1164_),
    .B1(_1163_));
 sg13g2_o21ai_1 _3826_ (.B1(_0791_),
    .Y(_1165_),
    .A1(_1162_),
    .A2(_1164_));
 sg13g2_nand2_1 _3827_ (.Y(_1166_),
    .A(net101),
    .B(_0751_));
 sg13g2_nand2_1 _3828_ (.Y(_1167_),
    .A(_0763_),
    .B(_0750_));
 sg13g2_and3_1 _3829_ (.X(_1168_),
    .A(net86),
    .B(_1166_),
    .C(_1167_));
 sg13g2_a22oi_1 _3830_ (.Y(_1169_),
    .B1(_1139_),
    .B2(_1166_),
    .A2(_0404_),
    .A1(net86));
 sg13g2_o21ai_1 _3831_ (.B1(_1132_),
    .Y(_1170_),
    .A1(_1168_),
    .A2(_1169_));
 sg13g2_nand2_1 _3832_ (.Y(_1171_),
    .A(_0776_),
    .B(_0405_));
 sg13g2_o21ai_1 _3833_ (.B1(_1171_),
    .Y(_1172_),
    .A1(net86),
    .A2(_0792_));
 sg13g2_o21ai_1 _3834_ (.B1(_1172_),
    .Y(_1173_),
    .A1(_1132_),
    .A2(_1140_));
 sg13g2_nand4_1 _3835_ (.B(_1107_),
    .C(_1170_),
    .A(_1165_),
    .Y(_1174_),
    .D(_1173_));
 sg13g2_buf_1 _3836_ (.A(_1174_),
    .X(_1175_));
 sg13g2_a21oi_1 _3837_ (.A1(_1118_),
    .A2(_1161_),
    .Y(_1176_),
    .B1(_1175_));
 sg13g2_nor2_1 _3838_ (.A(_1118_),
    .B(_1161_),
    .Y(_1177_));
 sg13g2_nand2_1 _3839_ (.Y(_1178_),
    .A(_1106_),
    .B(_1111_));
 sg13g2_o21ai_1 _3840_ (.B1(_1178_),
    .Y(_1179_),
    .A1(_1176_),
    .A2(_1177_));
 sg13g2_nor3_1 _3841_ (.A(_0897_),
    .B(_1096_),
    .C(_0892_),
    .Y(_1180_));
 sg13g2_nand2b_1 _3842_ (.Y(_1181_),
    .B(_0894_),
    .A_N(_1180_));
 sg13g2_nor2_1 _3843_ (.A(_1030_),
    .B(_0893_),
    .Y(_1182_));
 sg13g2_nand2_1 _3844_ (.Y(_1183_),
    .A(_1030_),
    .B(_0893_));
 sg13g2_o21ai_1 _3845_ (.B1(_1183_),
    .Y(_1184_),
    .A1(_0897_),
    .A2(_1182_));
 sg13g2_a21oi_1 _3846_ (.A1(_1181_),
    .A2(_1184_),
    .Y(_1185_),
    .B1(_0875_));
 sg13g2_a21oi_1 _3847_ (.A1(_0884_),
    .A2(_1180_),
    .Y(_1186_),
    .B1(_0875_));
 sg13g2_nand4_1 _3848_ (.B(_1012_),
    .C(_1024_),
    .A(_0995_),
    .Y(_1187_),
    .D(_1186_));
 sg13g2_nor2b_1 _3849_ (.A(_1185_),
    .B_N(_1187_),
    .Y(_1188_));
 sg13g2_nand2_1 _3850_ (.Y(_1189_),
    .A(_1149_),
    .B(_1160_));
 sg13g2_a21oi_1 _3851_ (.A1(_1175_),
    .A2(_1189_),
    .Y(_1190_),
    .B1(_1118_));
 sg13g2_nor2_1 _3852_ (.A(_1175_),
    .B(_1189_),
    .Y(_1191_));
 sg13g2_a221oi_1 _3853_ (.B2(_0893_),
    .C1(_0884_),
    .B1(_1030_),
    .A1(_0895_),
    .Y(_1192_),
    .A2(_0896_));
 sg13g2_nand3_1 _3854_ (.B(_1096_),
    .C(_0892_),
    .A(_0897_),
    .Y(_1193_));
 sg13g2_nand3_1 _3855_ (.B(_1096_),
    .C(_0892_),
    .A(_0894_),
    .Y(_1194_));
 sg13g2_nand3b_1 _3856_ (.B(_1193_),
    .C(_1194_),
    .Y(_1195_),
    .A_N(_1192_));
 sg13g2_and4_1 _3857_ (.A(_0995_),
    .B(_1012_),
    .C(_1024_),
    .D(_1195_),
    .X(_1196_));
 sg13g2_nand3_1 _3858_ (.B(_0897_),
    .C(_1182_),
    .A(_0894_),
    .Y(_1197_));
 sg13g2_o21ai_1 _3859_ (.B1(_1197_),
    .Y(_1198_),
    .A1(_1107_),
    .A2(_1106_));
 sg13g2_nor4_1 _3860_ (.A(_1190_),
    .B(_1191_),
    .C(_1196_),
    .D(_1198_),
    .Y(_1199_));
 sg13g2_a22oi_1 _3861_ (.Y(_1200_),
    .B1(_1188_),
    .B2(_1199_),
    .A2(_1179_),
    .A1(_1109_));
 sg13g2_buf_1 _3862_ (.A(_1200_),
    .X(_1201_));
 sg13g2_mux2_1 _3863_ (.A0(_1098_),
    .A1(_1037_),
    .S(net20),
    .X(_1202_));
 sg13g2_xnor2_1 _3864_ (.Y(_1203_),
    .A(_0901_),
    .B(_1202_));
 sg13g2_nand2b_1 _3865_ (.Y(_1204_),
    .B(_0815_),
    .A_N(_0725_));
 sg13g2_nand3_1 _3866_ (.B(_1203_),
    .C(_1204_),
    .A(_0820_),
    .Y(_1205_));
 sg13g2_nor3_1 _3867_ (.A(_1067_),
    .B(_1081_),
    .C(_1093_),
    .Y(_1206_));
 sg13g2_xnor2_1 _3868_ (.Y(_1207_),
    .A(_1030_),
    .B(_1032_));
 sg13g2_xor2_1 _3869_ (.B(_1207_),
    .A(_1026_),
    .X(_1208_));
 sg13g2_o21ai_1 _3870_ (.B1(_1208_),
    .Y(_1209_),
    .A1(net20),
    .A2(_1206_));
 sg13g2_buf_2 _3871_ (.A(_1209_),
    .X(_1210_));
 sg13g2_or3_1 _3872_ (.A(net20),
    .B(_1206_),
    .C(_1208_),
    .X(_1211_));
 sg13g2_buf_2 _3873_ (.A(_1211_),
    .X(_1212_));
 sg13g2_and3_1 _3874_ (.X(_1213_),
    .A(_0696_),
    .B(_1210_),
    .C(_1212_));
 sg13g2_nand3_1 _3875_ (.B(_0806_),
    .C(net19),
    .A(_0820_),
    .Y(_1214_));
 sg13g2_buf_1 _3876_ (.A(net20),
    .X(_1215_));
 sg13g2_nor2_1 _3877_ (.A(_0900_),
    .B(_0724_),
    .Y(_1216_));
 sg13g2_nand3b_1 _3878_ (.B(_1098_),
    .C(_1216_),
    .Y(_1217_),
    .A_N(net18));
 sg13g2_or4_1 _3879_ (.A(net20),
    .B(_0901_),
    .C(_0724_),
    .D(_1098_),
    .X(_1218_));
 sg13g2_nor2_1 _3880_ (.A(_0714_),
    .B(_0722_),
    .Y(_1219_));
 sg13g2_and3_1 _3881_ (.X(_1220_),
    .A(_0901_),
    .B(_1219_),
    .C(_1037_));
 sg13g2_nor3_1 _3882_ (.A(_0901_),
    .B(_0724_),
    .C(_1037_),
    .Y(_1221_));
 sg13g2_o21ai_1 _3883_ (.B1(net18),
    .Y(_1222_),
    .A1(_1220_),
    .A2(_1221_));
 sg13g2_nand4_1 _3884_ (.B(_1217_),
    .C(_1218_),
    .A(_1214_),
    .Y(_1223_),
    .D(_1222_));
 sg13g2_inv_1 _3885_ (.Y(_1224_),
    .A(_0696_));
 sg13g2_and4_1 _3886_ (.A(_0820_),
    .B(_1224_),
    .C(_1210_),
    .D(_1212_),
    .X(_1225_));
 sg13g2_a22oi_1 _3887_ (.Y(_1226_),
    .B1(_1225_),
    .B2(_1203_),
    .A2(_1223_),
    .A1(_1213_));
 sg13g2_and4_1 _3888_ (.A(_0689_),
    .B(_0696_),
    .C(_1210_),
    .D(_1212_),
    .X(_1227_));
 sg13g2_a21oi_1 _3889_ (.A1(_0806_),
    .A2(net19),
    .Y(_1228_),
    .B1(_0820_));
 sg13g2_and3_1 _3890_ (.X(_1229_),
    .A(_1210_),
    .B(_1212_),
    .C(_1228_));
 sg13g2_nor2_1 _3891_ (.A(_1224_),
    .B(_0724_),
    .Y(_1230_));
 sg13g2_nor2_1 _3892_ (.A(_0696_),
    .B(_1219_),
    .Y(_1231_));
 sg13g2_and4_1 _3893_ (.A(_1210_),
    .B(_1212_),
    .C(_1228_),
    .D(_1231_),
    .X(_1232_));
 sg13g2_a221oi_1 _3894_ (.B2(_1230_),
    .C1(_1232_),
    .B1(_1229_),
    .A1(_1203_),
    .Y(_1233_),
    .A2(_1227_));
 sg13g2_and2_1 _3895_ (.A(_0724_),
    .B(_1228_),
    .X(_1234_));
 sg13g2_and2_1 _3896_ (.A(_0696_),
    .B(_1228_),
    .X(_1235_));
 sg13g2_o21ai_1 _3897_ (.B1(_1203_),
    .Y(_1236_),
    .A1(_1234_),
    .A2(_1235_));
 sg13g2_nand4_1 _3898_ (.B(_1226_),
    .C(_1233_),
    .A(_1205_),
    .Y(_1237_),
    .D(_1236_));
 sg13g2_buf_1 _3899_ (.A(_1237_),
    .X(_1238_));
 sg13g2_inv_1 _3900_ (.Y(_1239_),
    .A(net20));
 sg13g2_mux2_1 _3901_ (.A0(_1033_),
    .A1(_1207_),
    .S(_1026_),
    .X(_1240_));
 sg13g2_nor2_1 _3902_ (.A(_0900_),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_nor3_1 _3903_ (.A(_1026_),
    .B(_0901_),
    .C(_1035_),
    .Y(_1242_));
 sg13g2_o21ai_1 _3904_ (.B1(_1206_),
    .Y(_1243_),
    .A1(_1241_),
    .A2(_1242_));
 sg13g2_nand2_1 _3905_ (.Y(_1244_),
    .A(_1239_),
    .B(_1243_));
 sg13g2_nand3b_1 _3906_ (.B(_1197_),
    .C(_1188_),
    .Y(_1245_),
    .A_N(_1196_));
 sg13g2_buf_1 _3907_ (.A(_1245_),
    .X(_1246_));
 sg13g2_xnor2_1 _3908_ (.Y(_1247_),
    .A(_1149_),
    .B(_1160_));
 sg13g2_xnor2_1 _3909_ (.Y(_1248_),
    .A(_1246_),
    .B(_1247_));
 sg13g2_xnor2_1 _3910_ (.Y(_1249_),
    .A(_1244_),
    .B(_1248_));
 sg13g2_a21oi_1 _3911_ (.A1(_0819_),
    .A2(_1238_),
    .Y(_1250_),
    .B1(_1249_));
 sg13g2_nor2_1 _3912_ (.A(_0819_),
    .B(_1238_),
    .Y(_1251_));
 sg13g2_xnor2_1 _3913_ (.Y(_1252_),
    .A(_1175_),
    .B(_1118_));
 sg13g2_or2_1 _3914_ (.X(_1253_),
    .B(net18),
    .A(_1189_));
 sg13g2_a21oi_1 _3915_ (.A1(_1160_),
    .A2(_1246_),
    .Y(_1254_),
    .B1(_1149_));
 sg13g2_nor2_1 _3916_ (.A(_1160_),
    .B(_1246_),
    .Y(_1255_));
 sg13g2_o21ai_1 _3917_ (.B1(net18),
    .Y(_1256_),
    .A1(_1254_),
    .A2(_1255_));
 sg13g2_inv_1 _3918_ (.Y(_1257_),
    .A(_1161_));
 sg13g2_nand4_1 _3919_ (.B(_1246_),
    .C(_1239_),
    .A(_1257_),
    .Y(_1258_),
    .D(_1243_));
 sg13g2_and4_1 _3920_ (.A(_1252_),
    .B(_1253_),
    .C(_1256_),
    .D(_1258_),
    .X(_1259_));
 sg13g2_buf_1 _3921_ (.A(_1259_),
    .X(_1260_));
 sg13g2_xnor2_1 _3922_ (.Y(_1261_),
    .A(_0768_),
    .B(_0786_));
 sg13g2_a21oi_1 _3923_ (.A1(net35),
    .A2(_0737_),
    .Y(_1262_),
    .B1(_0797_));
 sg13g2_nand3_1 _3924_ (.B(_0689_),
    .C(_0725_),
    .A(net35),
    .Y(_1263_));
 sg13g2_and3_1 _3925_ (.X(_1264_),
    .A(_1262_),
    .B(_1263_),
    .C(_0815_));
 sg13g2_nor4_1 _3926_ (.A(net35),
    .B(_0737_),
    .C(_0726_),
    .D(net19),
    .Y(_1265_));
 sg13g2_nor2_1 _3927_ (.A(net35),
    .B(_0737_),
    .Y(_1266_));
 sg13g2_nor3_1 _3928_ (.A(_1262_),
    .B(_0815_),
    .C(_1266_),
    .Y(_1267_));
 sg13g2_or4_1 _3929_ (.A(_1261_),
    .B(_1264_),
    .C(_1265_),
    .D(_1267_),
    .X(_1268_));
 sg13g2_buf_1 _3930_ (.A(_1268_),
    .X(_1269_));
 sg13g2_inv_1 _3931_ (.Y(_1270_),
    .A(_1269_));
 sg13g2_nand2_1 _3932_ (.Y(_1271_),
    .A(_1260_),
    .B(_1270_));
 sg13g2_o21ai_1 _3933_ (.B1(_1271_),
    .Y(_1272_),
    .A1(_1250_),
    .A2(_1251_));
 sg13g2_nand2b_1 _3934_ (.Y(_1273_),
    .B(_1269_),
    .A_N(_1260_));
 sg13g2_a21oi_1 _3935_ (.A1(_1272_),
    .A2(_1273_),
    .Y(_1274_),
    .B1(net110));
 sg13g2_nand2_2 _3936_ (.Y(_1275_),
    .A(_1210_),
    .B(_1212_));
 sg13g2_a21oi_1 _3937_ (.A1(_0806_),
    .A2(net19),
    .Y(_1276_),
    .B1(_1219_));
 sg13g2_xnor2_1 _3938_ (.Y(_1277_),
    .A(_1224_),
    .B(_1276_));
 sg13g2_xnor2_1 _3939_ (.Y(_1278_),
    .A(_1275_),
    .B(_1277_));
 sg13g2_xnor2_1 _3940_ (.Y(_1279_),
    .A(_0689_),
    .B(_1203_));
 sg13g2_xnor2_1 _3941_ (.Y(_1280_),
    .A(_1204_),
    .B(_1279_));
 sg13g2_xnor2_1 _3942_ (.Y(_1281_),
    .A(_0715_),
    .B(_0719_));
 sg13g2_xnor2_1 _3943_ (.Y(_1282_),
    .A(_0721_),
    .B(_1281_));
 sg13g2_inv_1 _3944_ (.Y(_1283_),
    .A(_0714_));
 sg13g2_a22oi_1 _3945_ (.Y(_1284_),
    .B1(_1282_),
    .B2(_1283_),
    .A2(net19),
    .A1(_0806_));
 sg13g2_or4_1 _3946_ (.A(_0590_),
    .B(_0631_),
    .C(_0666_),
    .D(_0672_),
    .X(_1285_));
 sg13g2_xnor2_1 _3947_ (.Y(_1286_),
    .A(_0717_),
    .B(_1285_));
 sg13g2_xnor2_1 _3948_ (.Y(_1287_),
    .A(_1284_),
    .B(_1286_));
 sg13g2_nor2_1 _3949_ (.A(_1081_),
    .B(_1093_),
    .Y(_1288_));
 sg13g2_nor2b_1 _3950_ (.A(net18),
    .B_N(_1067_),
    .Y(_1289_));
 sg13g2_xnor2_1 _3951_ (.Y(_1290_),
    .A(_1288_),
    .B(_1289_));
 sg13g2_nor2_2 _3952_ (.A(_1287_),
    .B(_1290_),
    .Y(_1291_));
 sg13g2_nand2_1 _3953_ (.Y(_1292_),
    .A(_0714_),
    .B(_0815_));
 sg13g2_xnor2_1 _3954_ (.Y(_1293_),
    .A(_1282_),
    .B(_1292_));
 sg13g2_buf_2 _3955_ (.A(_1293_),
    .X(_1294_));
 sg13g2_nor2_1 _3956_ (.A(_1291_),
    .B(_1294_),
    .Y(_1295_));
 sg13g2_nand3_1 _3957_ (.B(_1280_),
    .C(_1295_),
    .A(_1278_),
    .Y(_1296_));
 sg13g2_inv_1 _3958_ (.Y(_1297_),
    .A(_1291_));
 sg13g2_nand2_1 _3959_ (.Y(_1298_),
    .A(_1041_),
    .B(net20));
 sg13g2_nor2_1 _3960_ (.A(_0986_),
    .B(_1065_),
    .Y(_1299_));
 sg13g2_o21ai_1 _3961_ (.B1(_0966_),
    .Y(_1300_),
    .A1(net18),
    .A2(_1299_));
 sg13g2_a21oi_1 _3962_ (.A1(_1298_),
    .A2(_1300_),
    .Y(_1301_),
    .B1(_1039_));
 sg13g2_nand2_1 _3963_ (.Y(_1302_),
    .A(_0986_),
    .B(_1065_));
 sg13g2_o21ai_1 _3964_ (.B1(_1302_),
    .Y(_1303_),
    .A1(_0966_),
    .A2(_1299_));
 sg13g2_nand2_1 _3965_ (.Y(_1304_),
    .A(_1039_),
    .B(_1303_));
 sg13g2_o21ai_1 _3966_ (.B1(_1304_),
    .Y(_1305_),
    .A1(_0966_),
    .A2(_1302_));
 sg13g2_nand2b_1 _3967_ (.Y(_1306_),
    .B(_1305_),
    .A_N(net18));
 sg13g2_o21ai_1 _3968_ (.B1(_1306_),
    .Y(_1307_),
    .A1(_1040_),
    .A2(_1298_));
 sg13g2_xnor2_1 _3969_ (.Y(_1308_),
    .A(_0948_),
    .B(_1021_));
 sg13g2_o21ai_1 _3970_ (.B1(_1308_),
    .Y(_1309_),
    .A1(_1301_),
    .A2(_1307_));
 sg13g2_or3_1 _3971_ (.A(_1308_),
    .B(_1301_),
    .C(_1307_),
    .X(_1310_));
 sg13g2_nand2_2 _3972_ (.Y(_1311_),
    .A(_1309_),
    .B(_1310_));
 sg13g2_nand4_1 _3973_ (.B(_1280_),
    .C(_1297_),
    .A(_1278_),
    .Y(_1312_),
    .D(_1311_));
 sg13g2_nand2b_1 _3974_ (.Y(_1313_),
    .B(_1065_),
    .A_N(net18));
 sg13g2_xnor2_1 _3975_ (.Y(_1314_),
    .A(_1039_),
    .B(_1042_));
 sg13g2_xnor2_1 _3976_ (.Y(_1315_),
    .A(_1313_),
    .B(_1314_));
 sg13g2_a21oi_1 _3977_ (.A1(_0806_),
    .A2(net19),
    .Y(_1316_),
    .B1(_0713_));
 sg13g2_xnor2_1 _3978_ (.Y(_1317_),
    .A(_0515_),
    .B(_0697_));
 sg13g2_xnor2_1 _3979_ (.Y(_1318_),
    .A(_1316_),
    .B(_1317_));
 sg13g2_nand2_1 _3980_ (.Y(_1319_),
    .A(_1315_),
    .B(_1318_));
 sg13g2_inv_1 _3981_ (.Y(_1320_),
    .A(_0706_));
 sg13g2_a21oi_1 _3982_ (.A1(_0806_),
    .A2(net19),
    .Y(_1321_),
    .B1(_1320_));
 sg13g2_xor2_1 _3983_ (.B(_1321_),
    .A(_0712_),
    .X(_1322_));
 sg13g2_o21ai_1 _3984_ (.B1(net91),
    .Y(_1323_),
    .A1(net90),
    .A2(net68));
 sg13g2_nand2_1 _3985_ (.Y(_1324_),
    .A(_1050_),
    .B(_1323_));
 sg13g2_xnor2_1 _3986_ (.Y(_1325_),
    .A(_1055_),
    .B(_1324_));
 sg13g2_xnor2_1 _3987_ (.Y(_1326_),
    .A(net20),
    .B(_1325_));
 sg13g2_nand2b_1 _3988_ (.Y(_1327_),
    .B(net91),
    .A_N(net68));
 sg13g2_nand2_1 _3989_ (.Y(_1328_),
    .A(net76),
    .B(net68));
 sg13g2_xnor2_1 _3990_ (.Y(_1329_),
    .A(_0699_),
    .B(_0760_));
 sg13g2_and2_1 _3991_ (.A(net76),
    .B(net77),
    .X(_1330_));
 sg13g2_nor2_1 _3992_ (.A(_0483_),
    .B(net100),
    .Y(_1331_));
 sg13g2_a21oi_1 _3993_ (.A1(_0699_),
    .A2(_1330_),
    .Y(_1332_),
    .B1(_1331_));
 sg13g2_or3_1 _3994_ (.A(net76),
    .B(net77),
    .C(_0699_),
    .X(_1333_));
 sg13g2_nand2_1 _3995_ (.Y(_1334_),
    .A(net91),
    .B(_0699_));
 sg13g2_nand2_1 _3996_ (.Y(_1335_),
    .A(net76),
    .B(_0699_));
 sg13g2_mux2_1 _3997_ (.A0(_1334_),
    .A1(_1335_),
    .S(_0760_),
    .X(_1336_));
 sg13g2_o21ai_1 _3998_ (.B1(_1336_),
    .Y(_1337_),
    .A1(_0761_),
    .A2(_1333_));
 sg13g2_a22oi_1 _3999_ (.Y(_1338_),
    .B1(_1337_),
    .B2(_0700_),
    .A2(_1332_),
    .A1(_1329_));
 sg13g2_a21o_1 _4000_ (.A2(_0804_),
    .A1(_0737_),
    .B1(_0809_),
    .X(_1339_));
 sg13g2_nand2_1 _4001_ (.Y(_1340_),
    .A(_0768_),
    .B(_0807_));
 sg13g2_a21o_1 _4002_ (.A2(_0801_),
    .A1(_0797_),
    .B1(_0786_),
    .X(_1341_));
 sg13g2_inv_1 _4003_ (.Y(_1342_),
    .A(_0699_));
 sg13g2_nor2_1 _4004_ (.A(_1342_),
    .B(_0811_),
    .Y(_1343_));
 sg13g2_nand2_1 _4005_ (.Y(_1344_),
    .A(_0483_),
    .B(net77));
 sg13g2_and2_1 _4006_ (.A(_1342_),
    .B(_0811_),
    .X(_1345_));
 sg13g2_a21oi_1 _4007_ (.A1(_1343_),
    .A2(_1344_),
    .Y(_1346_),
    .B1(_1345_));
 sg13g2_a21oi_1 _4008_ (.A1(_1333_),
    .A2(_1335_),
    .Y(_1347_),
    .B1(_0811_));
 sg13g2_nor4_1 _4009_ (.A(net86),
    .B(net74),
    .C(_0810_),
    .D(_1334_),
    .Y(_1348_));
 sg13g2_o21ai_1 _4010_ (.B1(_0700_),
    .Y(_1349_),
    .A1(_1347_),
    .A2(_1348_));
 sg13g2_o21ai_1 _4011_ (.B1(_1349_),
    .Y(_1350_),
    .A1(_1331_),
    .A2(_1346_));
 sg13g2_a221oi_1 _4012_ (.B2(_1341_),
    .C1(_1350_),
    .B1(_1340_),
    .A1(_0737_),
    .Y(_1351_),
    .A2(_0804_));
 sg13g2_a221oi_1 _4013_ (.B2(_1339_),
    .C1(_1351_),
    .B1(_1338_),
    .A1(_1327_),
    .Y(_1352_),
    .A2(_1328_));
 sg13g2_nand2_2 _4014_ (.Y(_1353_),
    .A(_1327_),
    .B(_1328_));
 sg13g2_xnor2_1 _4015_ (.Y(_1354_),
    .A(net90),
    .B(_1325_));
 sg13g2_o21ai_1 _4016_ (.B1(_0706_),
    .Y(_1355_),
    .A1(_1353_),
    .A2(_1354_));
 sg13g2_a21oi_2 _4017_ (.B1(_1355_),
    .Y(_1356_),
    .A2(_1352_),
    .A1(_1326_));
 sg13g2_nor2_1 _4018_ (.A(_1322_),
    .B(_1356_),
    .Y(_1357_));
 sg13g2_o21ai_1 _4019_ (.B1(_1201_),
    .Y(_1358_),
    .A1(_1353_),
    .A2(_1325_));
 sg13g2_nand2_1 _4020_ (.Y(_1359_),
    .A(net90),
    .B(_1358_));
 sg13g2_inv_1 _4021_ (.Y(_1360_),
    .A(_1052_));
 sg13g2_a21oi_1 _4022_ (.A1(_1360_),
    .A2(_1324_),
    .Y(_1361_),
    .B1(_0974_));
 sg13g2_xnor2_1 _4023_ (.Y(_1362_),
    .A(_1049_),
    .B(_1361_));
 sg13g2_nor2b_1 _4024_ (.A(_1353_),
    .B_N(_1325_),
    .Y(_1363_));
 sg13g2_nor2_1 _4025_ (.A(_1215_),
    .B(_1363_),
    .Y(_1364_));
 sg13g2_nor2_1 _4026_ (.A(_1362_),
    .B(_1364_),
    .Y(_1365_));
 sg13g2_o21ai_1 _4027_ (.B1(_1057_),
    .Y(_1366_),
    .A1(_1215_),
    .A2(_1363_));
 sg13g2_and3_1 _4028_ (.X(_1367_),
    .A(_1362_),
    .B(_1358_),
    .C(_1366_));
 sg13g2_a221oi_1 _4029_ (.B2(_1365_),
    .C1(_1367_),
    .B1(_1359_),
    .A1(_1322_),
    .Y(_1368_),
    .A2(_1356_));
 sg13g2_or2_1 _4030_ (.X(_1369_),
    .B(_1318_),
    .A(_1315_));
 sg13g2_o21ai_1 _4031_ (.B1(_1369_),
    .Y(_1370_),
    .A1(_1357_),
    .A2(_1368_));
 sg13g2_nand2_2 _4032_ (.Y(_1371_),
    .A(_1319_),
    .B(_1370_));
 sg13g2_a21oi_1 _4033_ (.A1(_1296_),
    .A2(_1312_),
    .Y(_1372_),
    .B1(_1371_));
 sg13g2_nand2_2 _4034_ (.Y(_1373_),
    .A(_1287_),
    .B(_1290_));
 sg13g2_nand2_1 _4035_ (.Y(_1374_),
    .A(_1311_),
    .B(_1295_));
 sg13g2_nand2_1 _4036_ (.Y(_1375_),
    .A(_1278_),
    .B(_1280_));
 sg13g2_a21oi_1 _4037_ (.A1(_1373_),
    .A2(_1374_),
    .Y(_1376_),
    .B1(_1375_));
 sg13g2_or2_1 _4038_ (.X(_1377_),
    .B(_0819_),
    .A(_1249_));
 sg13g2_nand2_1 _4039_ (.Y(_1378_),
    .A(_1249_),
    .B(_0819_));
 sg13g2_xnor2_1 _4040_ (.Y(_1379_),
    .A(_1260_),
    .B(_1269_));
 sg13g2_mux2_1 _4041_ (.A0(_1377_),
    .A1(_1378_),
    .S(_1379_),
    .X(_1380_));
 sg13g2_nor4_1 _4042_ (.A(_1238_),
    .B(_1372_),
    .C(_1376_),
    .D(_1380_),
    .Y(_1381_));
 sg13g2_and2_1 _4043_ (.A(_1274_),
    .B(_1381_),
    .X(_1382_));
 sg13g2_buf_8 _4044_ (.A(_1382_),
    .X(_1383_));
 sg13g2_a21oi_1 _4045_ (.A1(_0359_),
    .A2(net110),
    .Y(_0071_),
    .B1(_1383_));
 sg13g2_inv_1 _4046_ (.Y(_1384_),
    .A(\gray_sobel0.out_px_sobel[1] ));
 sg13g2_nand2b_1 _4047_ (.Y(_1385_),
    .B(_0815_),
    .A_N(net77));
 sg13g2_nor2b_1 _4048_ (.A(_0815_),
    .B_N(net77),
    .Y(_1386_));
 sg13g2_a21oi_1 _4049_ (.A1(net100),
    .A2(_1385_),
    .Y(_1387_),
    .B1(_1386_));
 sg13g2_a21oi_1 _4050_ (.A1(_0806_),
    .A2(net19),
    .Y(_1388_),
    .B1(net77));
 sg13g2_a22oi_1 _4051_ (.Y(_1389_),
    .B1(_1388_),
    .B2(_1331_),
    .A2(_1386_),
    .A1(net100));
 sg13g2_o21ai_1 _4052_ (.B1(_1389_),
    .Y(_1390_),
    .A1(net91),
    .A2(_1387_));
 sg13g2_nor2_1 _4053_ (.A(_1057_),
    .B(_1353_),
    .Y(_1391_));
 sg13g2_a21oi_1 _4054_ (.A1(_1239_),
    .A2(_1353_),
    .Y(_1392_),
    .B1(_1391_));
 sg13g2_xnor2_1 _4055_ (.Y(_1393_),
    .A(_1342_),
    .B(_1325_));
 sg13g2_xnor2_1 _4056_ (.Y(_1394_),
    .A(_1392_),
    .B(_1393_));
 sg13g2_xnor2_1 _4057_ (.Y(_1395_),
    .A(_1390_),
    .B(_1394_));
 sg13g2_a22oi_1 _4058_ (.Y(_0072_),
    .B1(_1383_),
    .B2(_1395_),
    .A2(_1384_),
    .A1(net110));
 sg13g2_inv_1 _4059_ (.Y(_1396_),
    .A(\gray_sobel0.out_px_sobel[2] ));
 sg13g2_a21oi_1 _4060_ (.A1(_1359_),
    .A2(_1365_),
    .Y(_1397_),
    .B1(_1367_));
 sg13g2_xnor2_1 _4061_ (.Y(_1398_),
    .A(_1356_),
    .B(_1397_));
 sg13g2_xnor2_1 _4062_ (.Y(_1399_),
    .A(_1322_),
    .B(_1398_));
 sg13g2_a22oi_1 _4063_ (.Y(_0073_),
    .B1(_1383_),
    .B2(_1399_),
    .A2(_1396_),
    .A1(net110));
 sg13g2_inv_1 _4064_ (.Y(_1400_),
    .A(\gray_sobel0.out_px_sobel[3] ));
 sg13g2_nor2_1 _4065_ (.A(_1357_),
    .B(_1368_),
    .Y(_1401_));
 sg13g2_and2_1 _4066_ (.A(_1319_),
    .B(_1369_),
    .X(_1402_));
 sg13g2_xnor2_1 _4067_ (.Y(_1403_),
    .A(_1401_),
    .B(_1402_));
 sg13g2_a22oi_1 _4068_ (.Y(_0074_),
    .B1(_1383_),
    .B2(_1403_),
    .A2(_1400_),
    .A1(_0360_));
 sg13g2_inv_1 _4069_ (.Y(_1404_),
    .A(\gray_sobel0.out_px_sobel[4] ));
 sg13g2_and4_1 _4070_ (.A(_1238_),
    .B(_1379_),
    .C(_1378_),
    .D(_1377_),
    .X(_1405_));
 sg13g2_or2_1 _4071_ (.X(_1406_),
    .B(_1405_),
    .A(_1381_));
 sg13g2_xor2_1 _4072_ (.B(_1311_),
    .A(_1294_),
    .X(_1407_));
 sg13g2_xnor2_1 _4073_ (.Y(_1408_),
    .A(_1371_),
    .B(_1407_));
 sg13g2_and2_1 _4074_ (.A(_1274_),
    .B(_1408_),
    .X(_1409_));
 sg13g2_a22oi_1 _4075_ (.Y(_0075_),
    .B1(_1406_),
    .B2(_1409_),
    .A2(_1404_),
    .A1(net110));
 sg13g2_inv_1 _4076_ (.Y(_1410_),
    .A(\gray_sobel0.out_px_sobel[5] ));
 sg13g2_nand2_1 _4077_ (.Y(_1411_),
    .A(_1371_),
    .B(_1294_));
 sg13g2_inv_1 _4078_ (.Y(_1412_),
    .A(_1311_));
 sg13g2_o21ai_1 _4079_ (.B1(_1412_),
    .Y(_1413_),
    .A1(_1371_),
    .A2(_1294_));
 sg13g2_nand2_1 _4080_ (.Y(_1414_),
    .A(_1411_),
    .B(_1413_));
 sg13g2_nand2_1 _4081_ (.Y(_1415_),
    .A(_1373_),
    .B(_1297_));
 sg13g2_xnor2_1 _4082_ (.Y(_1416_),
    .A(_1414_),
    .B(_1415_));
 sg13g2_a22oi_1 _4083_ (.Y(_0076_),
    .B1(_1383_),
    .B2(_1416_),
    .A2(net110),
    .A1(_1410_));
 sg13g2_inv_1 _4084_ (.Y(_1417_),
    .A(\gray_sobel0.out_px_sobel[6] ));
 sg13g2_and2_1 _4085_ (.A(_1210_),
    .B(_1212_),
    .X(_1418_));
 sg13g2_buf_1 _4086_ (.A(_1418_),
    .X(_1419_));
 sg13g2_xnor2_1 _4087_ (.Y(_1420_),
    .A(_1419_),
    .B(_1277_));
 sg13g2_nand2_1 _4088_ (.Y(_1421_),
    .A(_1420_),
    .B(_1373_));
 sg13g2_or2_1 _4089_ (.X(_1422_),
    .B(_1421_),
    .A(_1413_));
 sg13g2_nand4_1 _4090_ (.B(_1297_),
    .C(_1411_),
    .A(_1278_),
    .Y(_1423_),
    .D(_1413_));
 sg13g2_or2_1 _4091_ (.X(_1424_),
    .B(_1421_),
    .A(_1411_));
 sg13g2_nor2_1 _4092_ (.A(_1420_),
    .B(_1373_),
    .Y(_1425_));
 sg13g2_a21oi_1 _4093_ (.A1(_1420_),
    .A2(_1291_),
    .Y(_1426_),
    .B1(_1425_));
 sg13g2_nand4_1 _4094_ (.B(_1423_),
    .C(_1424_),
    .A(_1422_),
    .Y(_1427_),
    .D(_1426_));
 sg13g2_a22oi_1 _4095_ (.Y(_0077_),
    .B1(_1383_),
    .B2(_1427_),
    .A2(net110),
    .A1(_1417_));
 sg13g2_inv_1 _4096_ (.Y(_1428_),
    .A(\gray_sobel0.out_px_sobel[7] ));
 sg13g2_xnor2_1 _4097_ (.Y(_1429_),
    .A(_0696_),
    .B(_1276_));
 sg13g2_nand3_1 _4098_ (.B(_1373_),
    .C(_1294_),
    .A(_1275_),
    .Y(_1430_));
 sg13g2_nand4_1 _4099_ (.B(_1373_),
    .C(_1309_),
    .A(_1275_),
    .Y(_1431_),
    .D(_1310_));
 sg13g2_a22oi_1 _4100_ (.Y(_1432_),
    .B1(_1430_),
    .B2(_1431_),
    .A2(_1370_),
    .A1(_1319_));
 sg13g2_nand2_1 _4101_ (.Y(_1433_),
    .A(_1275_),
    .B(_1291_));
 sg13g2_o21ai_1 _4102_ (.B1(_1433_),
    .Y(_1434_),
    .A1(_1311_),
    .A2(_1430_));
 sg13g2_nor3_1 _4103_ (.A(_1429_),
    .B(_1432_),
    .C(_1434_),
    .Y(_1435_));
 sg13g2_or3_1 _4104_ (.A(_1275_),
    .B(_1291_),
    .C(_1294_),
    .X(_1436_));
 sg13g2_nand3_1 _4105_ (.B(_1297_),
    .C(_1311_),
    .A(_1419_),
    .Y(_1437_));
 sg13g2_a21oi_1 _4106_ (.A1(_1436_),
    .A2(_1437_),
    .Y(_1438_),
    .B1(_1371_));
 sg13g2_nand3_1 _4107_ (.B(_1287_),
    .C(_1290_),
    .A(_1419_),
    .Y(_1439_));
 sg13g2_o21ai_1 _4108_ (.B1(_1439_),
    .Y(_1440_),
    .A1(_1412_),
    .A2(_1436_));
 sg13g2_nor3_1 _4109_ (.A(_1435_),
    .B(_1438_),
    .C(_1440_),
    .Y(_1441_));
 sg13g2_xor2_1 _4110_ (.B(_1441_),
    .A(_1280_),
    .X(_1442_));
 sg13g2_a22oi_1 _4111_ (.Y(_0078_),
    .B1(_1383_),
    .B2(_1442_),
    .A2(net110),
    .A1(_1428_));
 sg13g2_buf_1 _4112_ (.A(net180),
    .X(_1443_));
 sg13g2_nor2b_1 _4113_ (.A(net69),
    .B_N(\input_data[0] ),
    .Y(_1444_));
 sg13g2_a21oi_1 _4114_ (.A1(\lfsr0.lfsr_out[0] ),
    .A2(net67),
    .Y(_1445_),
    .B1(_1444_));
 sg13g2_nor2_1 _4115_ (.A(net180),
    .B(\gray_sobel0.gray_scale0.out_px_gray_o[0] ),
    .Y(_1446_));
 sg13g2_a21oi_2 _4116_ (.B1(_1446_),
    .Y(_1447_),
    .A2(_1445_),
    .A1(net96));
 sg13g2_nand2_1 _4117_ (.Y(_1448_),
    .A(net22),
    .B(_1447_));
 sg13g2_o21ai_1 _4118_ (.B1(_1448_),
    .Y(_0079_),
    .A1(_0700_),
    .A2(net22));
 sg13g2_nor2b_1 _4119_ (.A(_1916_),
    .B_N(\input_data[2] ),
    .Y(_1449_));
 sg13g2_a21oi_1 _4120_ (.A1(\lfsr0.lfsr_out[2] ),
    .A2(net67),
    .Y(_1450_),
    .B1(_1449_));
 sg13g2_nor2_1 _4121_ (.A(net180),
    .B(\gray_sobel0.gray_scale0.out_px_gray_o[2] ),
    .Y(_1451_));
 sg13g2_a21oi_2 _4122_ (.B1(_1451_),
    .Y(_1452_),
    .A2(_1450_),
    .A1(net96));
 sg13g2_and3_1 _4123_ (.X(_1453_),
    .A(net92),
    .B(_1940_),
    .C(net62));
 sg13g2_buf_1 _4124_ (.A(_1907_),
    .X(_1454_));
 sg13g2_nor3_1 _4125_ (.A(net92),
    .B(_1940_),
    .C(_1454_),
    .Y(_1455_));
 sg13g2_nor2_1 _4126_ (.A(_1939_),
    .B(_0349_),
    .Y(_1456_));
 sg13g2_o21ai_1 _4127_ (.B1(_1456_),
    .Y(_1457_),
    .A1(_1453_),
    .A2(_1455_));
 sg13g2_buf_4 _4128_ (.X(_1458_),
    .A(_1457_));
 sg13g2_mux2_1 _4129_ (.A0(_1452_),
    .A1(\gray_sobel0.sobel0.sobel.pix2_1[2] ),
    .S(_1458_),
    .X(_0080_));
 sg13g2_nor2b_1 _4130_ (.A(net69),
    .B_N(\input_data[3] ),
    .Y(_1459_));
 sg13g2_a21oi_1 _4131_ (.A1(_1835_),
    .A2(net67),
    .Y(_1460_),
    .B1(_1459_));
 sg13g2_nor2_1 _4132_ (.A(net180),
    .B(\gray_sobel0.gray_scale0.out_px_gray_o[3] ),
    .Y(_1461_));
 sg13g2_a21oi_2 _4133_ (.B1(_1461_),
    .Y(_1462_),
    .A2(_1460_),
    .A1(net96));
 sg13g2_mux2_1 _4134_ (.A0(_1462_),
    .A1(_0852_),
    .S(_1458_),
    .X(_0081_));
 sg13g2_nor2b_1 _4135_ (.A(net69),
    .B_N(_1966_),
    .Y(_1463_));
 sg13g2_a21oi_1 _4136_ (.A1(_1828_),
    .A2(net67),
    .Y(_1464_),
    .B1(_1463_));
 sg13g2_nor2_1 _4137_ (.A(net180),
    .B(\gray_sobel0.gray_scale0.out_px_gray_o[4] ),
    .Y(_1465_));
 sg13g2_a21oi_2 _4138_ (.B1(_1465_),
    .Y(_1466_),
    .A2(_1464_),
    .A1(net96));
 sg13g2_mux2_1 _4139_ (.A0(_1466_),
    .A1(_0847_),
    .S(_1458_),
    .X(_0082_));
 sg13g2_nor2b_1 _4140_ (.A(net69),
    .B_N(net115),
    .Y(_1467_));
 sg13g2_a21oi_1 _4141_ (.A1(net117),
    .A2(net67),
    .Y(_1468_),
    .B1(_1467_));
 sg13g2_nor2_1 _4142_ (.A(net96),
    .B(\gray_sobel0.gray_scale0.out_px_gray_o[5] ),
    .Y(_1469_));
 sg13g2_a21oi_2 _4143_ (.B1(_1469_),
    .Y(_1470_),
    .A2(_1468_),
    .A1(net96));
 sg13g2_mux2_1 _4144_ (.A0(_1470_),
    .A1(_0845_),
    .S(_1458_),
    .X(_0083_));
 sg13g2_nor2b_1 _4145_ (.A(net69),
    .B_N(net113),
    .Y(_1471_));
 sg13g2_a21oi_1 _4146_ (.A1(net119),
    .A2(net67),
    .Y(_1472_),
    .B1(_1471_));
 sg13g2_nor2_1 _4147_ (.A(net180),
    .B(\gray_sobel0.gray_scale0.out_px_gray_o[6] ),
    .Y(_1473_));
 sg13g2_a21oi_2 _4148_ (.B1(_1473_),
    .Y(_1474_),
    .A2(_1472_),
    .A1(net96));
 sg13g2_mux2_1 _4149_ (.A0(_1474_),
    .A1(_0871_),
    .S(_1458_),
    .X(_0084_));
 sg13g2_nor2b_1 _4150_ (.A(net69),
    .B_N(net112),
    .Y(_1475_));
 sg13g2_a21oi_1 _4151_ (.A1(net116),
    .A2(net67),
    .Y(_1476_),
    .B1(_1475_));
 sg13g2_nor2_1 _4152_ (.A(net180),
    .B(\gray_sobel0.gray_scale0.out_px_gray_o[7] ),
    .Y(_1477_));
 sg13g2_a21oi_2 _4153_ (.B1(_1477_),
    .Y(_1478_),
    .A2(_1476_),
    .A1(net96));
 sg13g2_mux2_1 _4154_ (.A0(_1478_),
    .A1(\gray_sobel0.sobel0.sobel.pix2_1[7] ),
    .S(_1458_),
    .X(_0085_));
 sg13g2_and2_1 _4155_ (.A(\gray_sobel0.sobel0.next[0] ),
    .B(_1948_),
    .X(_1479_));
 sg13g2_buf_1 _4156_ (.A(_1479_),
    .X(_1480_));
 sg13g2_nor2b_1 _4157_ (.A(_1939_),
    .B_N(_1940_),
    .Y(_1481_));
 sg13g2_nand3b_1 _4158_ (.B(_1481_),
    .C(net92),
    .Y(_1482_),
    .A_N(net111));
 sg13g2_nor2_1 _4159_ (.A(_1938_),
    .B(\gray_sobel0.sobel0.counter_sobel[0] ),
    .Y(_1483_));
 sg13g2_and2_1 _4160_ (.A(_0346_),
    .B(_1483_),
    .X(_1484_));
 sg13g2_nor2b_1 _4161_ (.A(_1937_),
    .B_N(_1948_),
    .Y(_1485_));
 sg13g2_o21ai_1 _4162_ (.B1(_1485_),
    .Y(_1486_),
    .A1(_1454_),
    .A2(_1484_));
 sg13g2_buf_1 _4163_ (.A(_1486_),
    .X(_1487_));
 sg13g2_a21o_1 _4164_ (.A2(_1482_),
    .A1(_1480_),
    .B1(_1487_),
    .X(_1488_));
 sg13g2_buf_4 _4165_ (.X(_1489_),
    .A(_1488_));
 sg13g2_mux2_1 _4166_ (.A0(_1447_),
    .A1(_0482_),
    .S(_1489_),
    .X(_0086_));
 sg13g2_nor2b_1 _4167_ (.A(net69),
    .B_N(\input_data[1] ),
    .Y(_1490_));
 sg13g2_a21oi_1 _4168_ (.A1(\lfsr0.lfsr_out[1] ),
    .A2(net67),
    .Y(_1491_),
    .B1(_1490_));
 sg13g2_nor2_1 _4169_ (.A(net180),
    .B(\gray_sobel0.gray_scale0.out_px_gray_o[1] ),
    .Y(_1492_));
 sg13g2_a21oi_2 _4170_ (.B1(_1492_),
    .Y(_1493_),
    .A2(_1491_),
    .A1(_1443_));
 sg13g2_mux2_1 _4171_ (.A0(_1493_),
    .A1(_0467_),
    .S(_1489_),
    .X(_0087_));
 sg13g2_mux2_1 _4172_ (.A0(_1452_),
    .A1(\gray_sobel0.sobel0.sobel.pix2_0[2] ),
    .S(_1489_),
    .X(_0088_));
 sg13g2_mux2_1 _4173_ (.A0(_1462_),
    .A1(_0525_),
    .S(_1489_),
    .X(_0089_));
 sg13g2_nand2_1 _4174_ (.Y(_1494_),
    .A(net21),
    .B(_1493_));
 sg13g2_o21ai_1 _4175_ (.B1(_1494_),
    .Y(_0090_),
    .A1(_1057_),
    .A2(net22));
 sg13g2_mux2_1 _4176_ (.A0(_1466_),
    .A1(_0555_),
    .S(_1489_),
    .X(_0091_));
 sg13g2_mux2_1 _4177_ (.A0(_1470_),
    .A1(net99),
    .S(_1489_),
    .X(_0092_));
 sg13g2_mux2_1 _4178_ (.A0(_1474_),
    .A1(_0400_),
    .S(_1489_),
    .X(_0093_));
 sg13g2_mux2_1 _4179_ (.A0(_1478_),
    .A1(_0776_),
    .S(_1489_),
    .X(_0094_));
 sg13g2_inv_1 _4180_ (.Y(_1495_),
    .A(_0438_));
 sg13g2_nor2b_1 _4181_ (.A(net92),
    .B_N(net111),
    .Y(_1496_));
 sg13g2_nand2_1 _4182_ (.Y(_1497_),
    .A(_1481_),
    .B(_1496_));
 sg13g2_a21o_1 _4183_ (.A2(_1497_),
    .A1(_1480_),
    .B1(_1487_),
    .X(_1498_));
 sg13g2_buf_2 _4184_ (.A(_1498_),
    .X(_1499_));
 sg13g2_buf_1 _4185_ (.A(_1499_),
    .X(_1500_));
 sg13g2_buf_1 _4186_ (.A(net54),
    .X(_1501_));
 sg13g2_buf_1 _4187_ (.A(net48),
    .X(_1502_));
 sg13g2_nand2_2 _4188_ (.Y(_1503_),
    .A(_1501_),
    .B(_1447_));
 sg13g2_o21ai_1 _4189_ (.B1(_1503_),
    .Y(_1504_),
    .A1(_0700_),
    .A2(_1502_));
 sg13g2_nor2_1 _4190_ (.A(net28),
    .B(_1504_),
    .Y(_1505_));
 sg13g2_a21oi_1 _4191_ (.A1(_1495_),
    .A2(net28),
    .Y(_0095_),
    .B1(_1505_));
 sg13g2_inv_1 _4192_ (.Y(_1506_),
    .A(_0436_));
 sg13g2_nand2_2 _4193_ (.Y(_1507_),
    .A(net54),
    .B(_1493_));
 sg13g2_o21ai_1 _4194_ (.B1(_1507_),
    .Y(_1508_),
    .A1(_1057_),
    .A2(_1502_));
 sg13g2_nor2_1 _4195_ (.A(_1500_),
    .B(_1508_),
    .Y(_1509_));
 sg13g2_a21oi_1 _4196_ (.A1(_1506_),
    .A2(_1500_),
    .Y(_0096_),
    .B1(_1509_));
 sg13g2_inv_1 _4197_ (.Y(_1510_),
    .A(\gray_sobel0.sobel0.sobel.pix1_2[2] ));
 sg13g2_nand2_2 _4198_ (.Y(_1511_),
    .A(net54),
    .B(_1452_));
 sg13g2_o21ai_1 _4199_ (.B1(_1511_),
    .Y(_1512_),
    .A1(_0538_),
    .A2(net47));
 sg13g2_nor2_1 _4200_ (.A(_1499_),
    .B(_1512_),
    .Y(_1513_));
 sg13g2_a21oi_1 _4201_ (.A1(_1510_),
    .A2(net28),
    .Y(_0097_),
    .B1(_1513_));
 sg13g2_nand2_2 _4202_ (.Y(_1514_),
    .A(net54),
    .B(_1462_));
 sg13g2_o21ai_1 _4203_ (.B1(_1514_),
    .Y(_1515_),
    .A1(net89),
    .A2(net47));
 sg13g2_nor2_1 _4204_ (.A(_1499_),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_a21oi_1 _4205_ (.A1(_0430_),
    .A2(net28),
    .Y(_0098_),
    .B1(_1516_));
 sg13g2_nand2_2 _4206_ (.Y(_1517_),
    .A(net54),
    .B(_1466_));
 sg13g2_o21ai_1 _4207_ (.B1(_1517_),
    .Y(_1518_),
    .A1(_0591_),
    .A2(net47));
 sg13g2_nor2_1 _4208_ (.A(_1499_),
    .B(_1518_),
    .Y(_1519_));
 sg13g2_a21oi_1 _4209_ (.A1(_0431_),
    .A2(net28),
    .Y(_0099_),
    .B1(_1519_));
 sg13g2_inv_1 _4210_ (.Y(_1520_),
    .A(net88));
 sg13g2_buf_1 _4211_ (.A(net48),
    .X(_1521_));
 sg13g2_nand2_2 _4212_ (.Y(_1522_),
    .A(net54),
    .B(_1470_));
 sg13g2_o21ai_1 _4213_ (.B1(_1522_),
    .Y(_1523_),
    .A1(_1520_),
    .A2(net46));
 sg13g2_nor2_1 _4214_ (.A(_1499_),
    .B(_1523_),
    .Y(_1524_));
 sg13g2_a21oi_1 _4215_ (.A1(_0423_),
    .A2(net28),
    .Y(_0100_),
    .B1(_1524_));
 sg13g2_nand2_1 _4216_ (.Y(_1525_),
    .A(net21),
    .B(_1452_));
 sg13g2_o21ai_1 _4217_ (.B1(_1525_),
    .Y(_0101_),
    .A1(_0538_),
    .A2(net22));
 sg13g2_nand2_2 _4218_ (.Y(_1526_),
    .A(net54),
    .B(_1474_));
 sg13g2_o21ai_1 _4219_ (.B1(_1526_),
    .Y(_1527_),
    .A1(_1133_),
    .A2(net46));
 sg13g2_nor2_1 _4220_ (.A(_1499_),
    .B(_1527_),
    .Y(_1528_));
 sg13g2_a21oi_1 _4221_ (.A1(_0452_),
    .A2(net28),
    .Y(_0102_),
    .B1(_1528_));
 sg13g2_inv_1 _4222_ (.Y(_1529_),
    .A(\gray_sobel0.sobel0.sobel.pix1_2[7] ));
 sg13g2_nand2_2 _4223_ (.Y(_1530_),
    .A(net54),
    .B(_1478_));
 sg13g2_o21ai_1 _4224_ (.B1(_1530_),
    .Y(_1531_),
    .A1(net74),
    .A2(net46));
 sg13g2_nor2_1 _4225_ (.A(_1499_),
    .B(_1531_),
    .Y(_1532_));
 sg13g2_a21oi_1 _4226_ (.A1(_1529_),
    .A2(net28),
    .Y(_0103_),
    .B1(_1532_));
 sg13g2_nand2_1 _4227_ (.Y(_1533_),
    .A(_1481_),
    .B(_1483_));
 sg13g2_a21o_1 _4228_ (.A2(_1533_),
    .A1(_1480_),
    .B1(_1487_),
    .X(_1534_));
 sg13g2_buf_1 _4229_ (.A(_1534_),
    .X(_1535_));
 sg13g2_buf_1 _4230_ (.A(_1535_),
    .X(_1536_));
 sg13g2_nand2_1 _4231_ (.Y(_1537_),
    .A(\gray_sobel0.sobel0.sobel.pix2_1[0] ),
    .B(net51));
 sg13g2_a21oi_1 _4232_ (.A1(_1503_),
    .A2(_1537_),
    .Y(_1538_),
    .B1(net27));
 sg13g2_a21o_1 _4233_ (.A2(net27),
    .A1(\gray_sobel0.sobel0.sobel.pix1_1[0] ),
    .B1(_1538_),
    .X(_0104_));
 sg13g2_nand2_1 _4234_ (.Y(_1539_),
    .A(_0854_),
    .B(net51));
 sg13g2_a21oi_1 _4235_ (.A1(_1507_),
    .A2(_1539_),
    .Y(_1540_),
    .B1(_1536_));
 sg13g2_a21o_1 _4236_ (.A2(_1536_),
    .A1(\gray_sobel0.sobel0.sobel.pix1_1[1] ),
    .B1(_1540_),
    .X(_0105_));
 sg13g2_nand2_1 _4237_ (.Y(_1541_),
    .A(\gray_sobel0.sobel0.sobel.pix2_1[2] ),
    .B(net51));
 sg13g2_a21oi_1 _4238_ (.A1(_1511_),
    .A2(_1541_),
    .Y(_1542_),
    .B1(_1535_));
 sg13g2_a21o_1 _4239_ (.A2(net27),
    .A1(\gray_sobel0.sobel0.sobel.pix1_1[2] ),
    .B1(_1542_),
    .X(_0106_));
 sg13g2_buf_1 _4240_ (.A(net48),
    .X(_1543_));
 sg13g2_o21ai_1 _4241_ (.B1(_1514_),
    .Y(_1544_),
    .A1(_0876_),
    .A2(net45));
 sg13g2_mux2_1 _4242_ (.A0(_1544_),
    .A1(\gray_sobel0.sobel0.sobel.pix1_1[3] ),
    .S(net27),
    .X(_0107_));
 sg13g2_o21ai_1 _4243_ (.B1(_1517_),
    .Y(_1545_),
    .A1(_0848_),
    .A2(net45));
 sg13g2_mux2_1 _4244_ (.A0(_1545_),
    .A1(\gray_sobel0.sobel0.sobel.pix1_1[4] ),
    .S(net27),
    .X(_0108_));
 sg13g2_nand2_1 _4245_ (.Y(_1546_),
    .A(_0845_),
    .B(net51));
 sg13g2_a21oi_1 _4246_ (.A1(_1522_),
    .A2(_1546_),
    .Y(_1547_),
    .B1(_1535_));
 sg13g2_a21o_1 _4247_ (.A2(net27),
    .A1(\gray_sobel0.sobel0.sobel.pix1_1[5] ),
    .B1(_1547_),
    .X(_0109_));
 sg13g2_o21ai_1 _4248_ (.B1(_1526_),
    .Y(_1548_),
    .A1(_1102_),
    .A2(_1543_));
 sg13g2_mux2_1 _4249_ (.A0(_1548_),
    .A1(\gray_sobel0.sobel0.sobel.pix1_1[6] ),
    .S(net27),
    .X(_0110_));
 sg13g2_o21ai_1 _4250_ (.B1(_1530_),
    .Y(_1549_),
    .A1(_1110_),
    .A2(_1543_));
 sg13g2_mux2_1 _4251_ (.A0(_1549_),
    .A1(\gray_sobel0.sobel0.sobel.pix1_1[7] ),
    .S(net27),
    .X(_0111_));
 sg13g2_nand2_1 _4252_ (.Y(_1550_),
    .A(net21),
    .B(_1462_));
 sg13g2_o21ai_1 _4253_ (.B1(_1550_),
    .Y(_0112_),
    .A1(net89),
    .A2(net22));
 sg13g2_inv_1 _4254_ (.Y(_1551_),
    .A(_0439_));
 sg13g2_nand3_1 _4255_ (.B(net111),
    .C(_0346_),
    .A(net92),
    .Y(_1552_));
 sg13g2_a21oi_1 _4256_ (.A1(net62),
    .A2(_1552_),
    .Y(_1553_),
    .B1(_1487_));
 sg13g2_buf_2 _4257_ (.A(_1553_),
    .X(_1554_));
 sg13g2_buf_1 _4258_ (.A(_1554_),
    .X(_1555_));
 sg13g2_o21ai_1 _4259_ (.B1(_1503_),
    .Y(_1556_),
    .A1(net76),
    .A2(_1521_));
 sg13g2_nand2_1 _4260_ (.Y(_1557_),
    .A(net26),
    .B(_1556_));
 sg13g2_o21ai_1 _4261_ (.B1(_1557_),
    .Y(_0113_),
    .A1(_1551_),
    .A2(net26));
 sg13g2_inv_1 _4262_ (.Y(_1558_),
    .A(_0435_));
 sg13g2_o21ai_1 _4263_ (.B1(_1507_),
    .Y(_1559_),
    .A1(_0508_),
    .A2(_1521_));
 sg13g2_nand2_1 _4264_ (.Y(_1560_),
    .A(net26),
    .B(_1559_));
 sg13g2_o21ai_1 _4265_ (.B1(_1560_),
    .Y(_0114_),
    .A1(_1558_),
    .A2(net26));
 sg13g2_o21ai_1 _4266_ (.B1(_1511_),
    .Y(_1561_),
    .A1(_0537_),
    .A2(net46));
 sg13g2_nand2_1 _4267_ (.Y(_1562_),
    .A(_1554_),
    .B(_1561_));
 sg13g2_o21ai_1 _4268_ (.B1(_1562_),
    .Y(_0115_),
    .A1(_0563_),
    .A2(_1555_));
 sg13g2_inv_1 _4269_ (.Y(_1563_),
    .A(_0426_));
 sg13g2_o21ai_1 _4270_ (.B1(_1514_),
    .Y(_1564_),
    .A1(_0579_),
    .A2(net46));
 sg13g2_nand2_1 _4271_ (.Y(_1565_),
    .A(_1554_),
    .B(_1564_));
 sg13g2_o21ai_1 _4272_ (.B1(_1565_),
    .Y(_0116_),
    .A1(_1563_),
    .A2(net26));
 sg13g2_inv_1 _4273_ (.Y(_1566_),
    .A(\gray_sobel0.sobel0.sobel.pix1_0[4] ));
 sg13g2_o21ai_1 _4274_ (.B1(_1517_),
    .Y(_1567_),
    .A1(_0556_),
    .A2(net46));
 sg13g2_nand2_1 _4275_ (.Y(_1568_),
    .A(_1554_),
    .B(_1567_));
 sg13g2_o21ai_1 _4276_ (.B1(_1568_),
    .Y(_0117_),
    .A1(_1566_),
    .A2(net26));
 sg13g2_inv_1 _4277_ (.Y(_1569_),
    .A(_0448_));
 sg13g2_o21ai_1 _4278_ (.B1(_1522_),
    .Y(_1570_),
    .A1(_0653_),
    .A2(net46));
 sg13g2_nand2_1 _4279_ (.Y(_1571_),
    .A(_1554_),
    .B(_1570_));
 sg13g2_o21ai_1 _4280_ (.B1(_1571_),
    .Y(_0118_),
    .A1(_1569_),
    .A2(net26));
 sg13g2_inv_1 _4281_ (.Y(_1572_),
    .A(\gray_sobel0.sobel0.sobel.pix1_0[6] ));
 sg13g2_o21ai_1 _4282_ (.B1(_1526_),
    .Y(_1573_),
    .A1(_0401_),
    .A2(net46));
 sg13g2_nand2_1 _4283_ (.Y(_1574_),
    .A(_1554_),
    .B(_1573_));
 sg13g2_o21ai_1 _4284_ (.B1(_1574_),
    .Y(_0119_),
    .A1(_1572_),
    .A2(_1555_));
 sg13g2_o21ai_1 _4285_ (.B1(_1530_),
    .Y(_1575_),
    .A1(_0749_),
    .A2(net48));
 sg13g2_nand2_1 _4286_ (.Y(_1576_),
    .A(_1554_),
    .B(_1575_));
 sg13g2_o21ai_1 _4287_ (.B1(_1576_),
    .Y(_0120_),
    .A1(_0745_),
    .A2(net26));
 sg13g2_a21oi_1 _4288_ (.A1(net62),
    .A2(_1944_),
    .Y(_1577_),
    .B1(_1487_));
 sg13g2_buf_1 _4289_ (.A(_1577_),
    .X(_1578_));
 sg13g2_o21ai_1 _4290_ (.B1(_1503_),
    .Y(_1579_),
    .A1(_1495_),
    .A2(_1501_));
 sg13g2_nand2_1 _4291_ (.Y(_1580_),
    .A(net31),
    .B(_1579_));
 sg13g2_o21ai_1 _4292_ (.B1(_1580_),
    .Y(_0121_),
    .A1(_0952_),
    .A2(net31));
 sg13g2_o21ai_1 _4293_ (.B1(_1507_),
    .Y(_1581_),
    .A1(_1506_),
    .A2(net45));
 sg13g2_mux2_1 _4294_ (.A0(_0374_),
    .A1(_1581_),
    .S(net31),
    .X(_0122_));
 sg13g2_nand2_1 _4295_ (.Y(_1582_),
    .A(net21),
    .B(_1466_));
 sg13g2_o21ai_1 _4296_ (.B1(_1582_),
    .Y(_0123_),
    .A1(_0591_),
    .A2(net22));
 sg13g2_o21ai_1 _4297_ (.B1(_1511_),
    .Y(_1583_),
    .A1(_1510_),
    .A2(net45));
 sg13g2_mux2_1 _4298_ (.A0(net104),
    .A1(_1583_),
    .S(net31),
    .X(_0124_));
 sg13g2_o21ai_1 _4299_ (.B1(_1514_),
    .Y(_1584_),
    .A1(_0430_),
    .A2(net45));
 sg13g2_mux2_1 _4300_ (.A0(net105),
    .A1(_1584_),
    .S(net31),
    .X(_0125_));
 sg13g2_o21ai_1 _4301_ (.B1(_1517_),
    .Y(_1585_),
    .A1(_0431_),
    .A2(net45));
 sg13g2_mux2_1 _4302_ (.A0(_0366_),
    .A1(_1585_),
    .S(net31),
    .X(_0126_));
 sg13g2_o21ai_1 _4303_ (.B1(_1522_),
    .Y(_1586_),
    .A1(_0423_),
    .A2(net45));
 sg13g2_mux2_1 _4304_ (.A0(net106),
    .A1(_1586_),
    .S(net31),
    .X(_0127_));
 sg13g2_o21ai_1 _4305_ (.B1(_1526_),
    .Y(_1587_),
    .A1(_0452_),
    .A2(net48));
 sg13g2_nand2_1 _4306_ (.Y(_1588_),
    .A(_1578_),
    .B(_1587_));
 sg13g2_o21ai_1 _4307_ (.B1(_1588_),
    .Y(_0128_),
    .A1(_0410_),
    .A2(net31));
 sg13g2_o21ai_1 _4308_ (.B1(_1530_),
    .Y(_1589_),
    .A1(_1529_),
    .A2(net48));
 sg13g2_nand2_1 _4309_ (.Y(_1590_),
    .A(_1577_),
    .B(_1589_));
 sg13g2_o21ai_1 _4310_ (.B1(_1590_),
    .Y(_0129_),
    .A1(net87),
    .A2(_1578_));
 sg13g2_nand2_1 _4311_ (.Y(_1591_),
    .A(_0346_),
    .B(_1496_));
 sg13g2_a21o_1 _4312_ (.A2(_1591_),
    .A1(_1480_),
    .B1(_1487_),
    .X(_1592_));
 sg13g2_buf_1 _4313_ (.A(_1592_),
    .X(_1593_));
 sg13g2_buf_1 _4314_ (.A(_1593_),
    .X(_1594_));
 sg13g2_nand2_1 _4315_ (.Y(_1595_),
    .A(\gray_sobel0.sobel0.sobel.pix1_1[0] ),
    .B(\gray_sobel0.sobel0.next[1] ));
 sg13g2_a21oi_1 _4316_ (.A1(_1503_),
    .A2(_1595_),
    .Y(_1596_),
    .B1(net25));
 sg13g2_a21o_1 _4317_ (.A2(net25),
    .A1(\gray_sobel0.sobel0.sobel.pix0_1[0] ),
    .B1(_1596_),
    .X(_0130_));
 sg13g2_nand2_1 _4318_ (.Y(_1597_),
    .A(\gray_sobel0.sobel0.sobel.pix1_1[1] ),
    .B(net51));
 sg13g2_a21oi_1 _4319_ (.A1(_1507_),
    .A2(_1597_),
    .Y(_1598_),
    .B1(_1594_));
 sg13g2_a21o_1 _4320_ (.A2(net25),
    .A1(\gray_sobel0.sobel0.sobel.pix0_1[1] ),
    .B1(_1598_),
    .X(_0131_));
 sg13g2_nand2_1 _4321_ (.Y(_1599_),
    .A(\gray_sobel0.sobel0.sobel.pix1_1[2] ),
    .B(net51));
 sg13g2_a21oi_1 _4322_ (.A1(_1511_),
    .A2(_1599_),
    .Y(_1600_),
    .B1(_1593_));
 sg13g2_a21o_1 _4323_ (.A2(net25),
    .A1(\gray_sobel0.sobel0.sobel.pix0_1[2] ),
    .B1(_1600_),
    .X(_0132_));
 sg13g2_nand2_1 _4324_ (.Y(_1601_),
    .A(\gray_sobel0.sobel0.sobel.pix1_1[3] ),
    .B(net51));
 sg13g2_a21oi_1 _4325_ (.A1(_1514_),
    .A2(_1601_),
    .Y(_1602_),
    .B1(_1593_));
 sg13g2_a21o_1 _4326_ (.A2(_1594_),
    .A1(_0862_),
    .B1(_1602_),
    .X(_0133_));
 sg13g2_nand2_1 _4327_ (.Y(_1603_),
    .A(net21),
    .B(_1470_));
 sg13g2_o21ai_1 _4328_ (.B1(_1603_),
    .Y(_0134_),
    .A1(_1520_),
    .A2(net22));
 sg13g2_nand2_1 _4329_ (.Y(_1604_),
    .A(\gray_sobel0.sobel0.sobel.pix1_1[4] ),
    .B(net51));
 sg13g2_a21oi_1 _4330_ (.A1(_1517_),
    .A2(_1604_),
    .Y(_1605_),
    .B1(_1593_));
 sg13g2_a21o_1 _4331_ (.A2(net25),
    .A1(_0849_),
    .B1(_1605_),
    .X(_0135_));
 sg13g2_nand2_1 _4332_ (.Y(_1606_),
    .A(\gray_sobel0.sobel0.sobel.pix1_1[5] ),
    .B(_1908_));
 sg13g2_a21oi_1 _4333_ (.A1(_1522_),
    .A2(_1606_),
    .Y(_1607_),
    .B1(_1593_));
 sg13g2_a21o_1 _4334_ (.A2(net25),
    .A1(\gray_sobel0.sobel0.sobel.pix0_1[5] ),
    .B1(_1607_),
    .X(_0136_));
 sg13g2_nand2_1 _4335_ (.Y(_1608_),
    .A(\gray_sobel0.sobel0.sobel.pix1_1[6] ),
    .B(_1908_));
 sg13g2_a21oi_1 _4336_ (.A1(_1526_),
    .A2(_1608_),
    .Y(_1609_),
    .B1(_1593_));
 sg13g2_a21o_1 _4337_ (.A2(net25),
    .A1(_0872_),
    .B1(_1609_),
    .X(_0137_));
 sg13g2_nand2_1 _4338_ (.Y(_1610_),
    .A(\gray_sobel0.sobel0.sobel.pix1_1[7] ),
    .B(_1908_));
 sg13g2_a21oi_1 _4339_ (.A1(_1530_),
    .A2(_1610_),
    .Y(_1611_),
    .B1(_1593_));
 sg13g2_a21o_1 _4340_ (.A2(net25),
    .A1(\gray_sobel0.sobel0.sobel.pix0_1[7] ),
    .B1(_1611_),
    .X(_0138_));
 sg13g2_o21ai_1 _4341_ (.B1(_1503_),
    .Y(_1612_),
    .A1(_1551_),
    .A2(net45));
 sg13g2_and2_1 _4342_ (.A(_1485_),
    .B(_1484_),
    .X(_1613_));
 sg13g2_buf_1 _4343_ (.A(_1613_),
    .X(_1614_));
 sg13g2_mux2_1 _4344_ (.A0(_0377_),
    .A1(_1612_),
    .S(_1614_),
    .X(_0139_));
 sg13g2_o21ai_1 _4345_ (.B1(_1507_),
    .Y(_1615_),
    .A1(_1558_),
    .A2(net47));
 sg13g2_mux2_1 _4346_ (.A0(_0375_),
    .A1(_1615_),
    .S(net34),
    .X(_0140_));
 sg13g2_o21ai_1 _4347_ (.B1(_1511_),
    .Y(_1616_),
    .A1(_0563_),
    .A2(net48));
 sg13g2_nand2_1 _4348_ (.Y(_1617_),
    .A(net34),
    .B(_1616_));
 sg13g2_o21ai_1 _4349_ (.B1(_1617_),
    .Y(_0141_),
    .A1(_0520_),
    .A2(_1614_));
 sg13g2_o21ai_1 _4350_ (.B1(_1514_),
    .Y(_1618_),
    .A1(_1563_),
    .A2(net47));
 sg13g2_mux2_1 _4351_ (.A0(_0390_),
    .A1(_1618_),
    .S(net34),
    .X(_0142_));
 sg13g2_o21ai_1 _4352_ (.B1(_1517_),
    .Y(_1619_),
    .A1(_1566_),
    .A2(net47));
 sg13g2_mux2_1 _4353_ (.A0(_0365_),
    .A1(_1619_),
    .S(net34),
    .X(_0143_));
 sg13g2_o21ai_1 _4354_ (.B1(_1522_),
    .Y(_1620_),
    .A1(_1569_),
    .A2(net47));
 sg13g2_mux2_1 _4355_ (.A0(net107),
    .A1(_1620_),
    .S(net34),
    .X(_0144_));
 sg13g2_nand2_1 _4356_ (.Y(_1621_),
    .A(net21),
    .B(_1474_));
 sg13g2_o21ai_1 _4357_ (.B1(_1621_),
    .Y(_0145_),
    .A1(_1133_),
    .A2(net22));
 sg13g2_o21ai_1 _4358_ (.B1(_1526_),
    .Y(_1622_),
    .A1(_1572_),
    .A2(net48));
 sg13g2_nand2_1 _4359_ (.Y(_1623_),
    .A(net34),
    .B(_1622_));
 sg13g2_o21ai_1 _4360_ (.B1(_1623_),
    .Y(_0146_),
    .A1(_0416_),
    .A2(net34));
 sg13g2_o21ai_1 _4361_ (.B1(_1530_),
    .Y(_1624_),
    .A1(_0745_),
    .A2(net47));
 sg13g2_mux2_1 _4362_ (.A0(net97),
    .A1(_1624_),
    .S(net34),
    .X(_0147_));
 sg13g2_nand2_1 _4363_ (.Y(_1625_),
    .A(net21),
    .B(_1478_));
 sg13g2_o21ai_1 _4364_ (.B1(_1625_),
    .Y(_0148_),
    .A1(net74),
    .A2(_0001_));
 sg13g2_mux2_1 _4365_ (.A0(_1447_),
    .A1(\gray_sobel0.sobel0.sobel.pix2_1[0] ),
    .S(_1458_),
    .X(_0149_));
 sg13g2_mux2_1 _4366_ (.A0(_1493_),
    .A1(_0854_),
    .S(_1458_),
    .X(_0150_));
 sg13g2_xnor2_1 _4367_ (.Y(_1626_),
    .A(_1835_),
    .B(net118));
 sg13g2_buf_1 _4368_ (.A(_1871_),
    .X(_1627_));
 sg13g2_nor2b_1 _4369_ (.A(net85),
    .B_N(\lfsr0.seed_reg[0] ),
    .Y(_1628_));
 sg13g2_a21oi_1 _4370_ (.A1(net79),
    .A2(_1626_),
    .Y(_1629_),
    .B1(_1628_));
 sg13g2_nor2_1 _4371_ (.A(\lfsr0.lfsr_out[0] ),
    .B(net63),
    .Y(_1630_));
 sg13g2_a21oi_1 _4372_ (.A1(net64),
    .A2(_1629_),
    .Y(_0151_),
    .B1(_1630_));
 sg13g2_nor2b_1 _4373_ (.A(net85),
    .B_N(\lfsr0.seed_reg[10] ),
    .Y(_1631_));
 sg13g2_a21oi_1 _4374_ (.A1(_1831_),
    .A2(net79),
    .Y(_1632_),
    .B1(_1631_));
 sg13g2_nor2_1 _4375_ (.A(\lfsr0.lfsr_out[10] ),
    .B(net63),
    .Y(_1633_));
 sg13g2_a21oi_1 _4376_ (.A1(net64),
    .A2(_1632_),
    .Y(_0152_),
    .B1(_1633_));
 sg13g2_nor2b_1 _4377_ (.A(net85),
    .B_N(\lfsr0.seed_reg[11] ),
    .Y(_1634_));
 sg13g2_a21oi_1 _4378_ (.A1(\lfsr0.lfsr_out[10] ),
    .A2(net79),
    .Y(_1635_),
    .B1(_1634_));
 sg13g2_nor2_1 _4379_ (.A(\lfsr0.lfsr_out[11] ),
    .B(net63),
    .Y(_1636_));
 sg13g2_a21oi_1 _4380_ (.A1(net64),
    .A2(_1635_),
    .Y(_0153_),
    .B1(_1636_));
 sg13g2_nor2b_1 _4381_ (.A(net85),
    .B_N(\lfsr0.seed_reg[12] ),
    .Y(_1637_));
 sg13g2_a21oi_1 _4382_ (.A1(\lfsr0.lfsr_out[11] ),
    .A2(net79),
    .Y(_1638_),
    .B1(_1637_));
 sg13g2_nor2_1 _4383_ (.A(net118),
    .B(_1874_),
    .Y(_1639_));
 sg13g2_a21oi_1 _4384_ (.A1(_1870_),
    .A2(_1638_),
    .Y(_0154_),
    .B1(_1639_));
 sg13g2_nor2b_1 _4385_ (.A(_1627_),
    .B_N(\lfsr0.seed_reg[13] ),
    .Y(_1640_));
 sg13g2_a21oi_1 _4386_ (.A1(_1842_),
    .A2(net79),
    .Y(_1641_),
    .B1(_1640_));
 sg13g2_buf_1 _4387_ (.A(_1869_),
    .X(_1642_));
 sg13g2_nor2_1 _4388_ (.A(\lfsr0.lfsr_out[13] ),
    .B(net58),
    .Y(_1643_));
 sg13g2_a21oi_1 _4389_ (.A1(net64),
    .A2(_1641_),
    .Y(_0155_),
    .B1(_1643_));
 sg13g2_buf_1 _4390_ (.A(_1871_),
    .X(_1644_));
 sg13g2_nor2b_1 _4391_ (.A(net84),
    .B_N(\lfsr0.seed_reg[14] ),
    .Y(_1645_));
 sg13g2_a21oi_1 _4392_ (.A1(\lfsr0.lfsr_out[13] ),
    .A2(net79),
    .Y(_1646_),
    .B1(_1645_));
 sg13g2_nor2_1 _4393_ (.A(\lfsr0.lfsr_out[14] ),
    .B(net58),
    .Y(_1647_));
 sg13g2_a21oi_1 _4394_ (.A1(net64),
    .A2(_1646_),
    .Y(_0156_),
    .B1(_1647_));
 sg13g2_nor2b_1 _4395_ (.A(net84),
    .B_N(\lfsr0.seed_reg[15] ),
    .Y(_1648_));
 sg13g2_a21oi_1 _4396_ (.A1(\lfsr0.lfsr_out[14] ),
    .A2(net79),
    .Y(_1649_),
    .B1(_1648_));
 sg13g2_nor2_1 _4397_ (.A(\lfsr0.lfsr_out[15] ),
    .B(net58),
    .Y(_1650_));
 sg13g2_a21oi_1 _4398_ (.A1(net64),
    .A2(_1649_),
    .Y(_0157_),
    .B1(_1650_));
 sg13g2_nor2b_1 _4399_ (.A(_1644_),
    .B_N(\lfsr0.seed_reg[16] ),
    .Y(_1651_));
 sg13g2_a21oi_1 _4400_ (.A1(\lfsr0.lfsr_out[15] ),
    .A2(_1873_),
    .Y(_1652_),
    .B1(_1651_));
 sg13g2_nor2_1 _4401_ (.A(\lfsr0.lfsr_out[16] ),
    .B(_1642_),
    .Y(_1653_));
 sg13g2_a21oi_1 _4402_ (.A1(net64),
    .A2(_1652_),
    .Y(_0158_),
    .B1(_1653_));
 sg13g2_nor2b_1 _4403_ (.A(_1644_),
    .B_N(\lfsr0.seed_reg[17] ),
    .Y(_1654_));
 sg13g2_a21oi_1 _4404_ (.A1(\lfsr0.lfsr_out[16] ),
    .A2(_1873_),
    .Y(_1655_),
    .B1(_1654_));
 sg13g2_nor2_1 _4405_ (.A(\lfsr0.lfsr_out[17] ),
    .B(_1642_),
    .Y(_1656_));
 sg13g2_a21oi_1 _4406_ (.A1(_1870_),
    .A2(_1655_),
    .Y(_0159_),
    .B1(_1656_));
 sg13g2_buf_1 _4407_ (.A(_1869_),
    .X(_1657_));
 sg13g2_buf_1 _4408_ (.A(_1871_),
    .X(_1658_));
 sg13g2_nor2b_1 _4409_ (.A(net84),
    .B_N(\lfsr0.seed_reg[18] ),
    .Y(_1659_));
 sg13g2_a21oi_1 _4410_ (.A1(\lfsr0.lfsr_out[17] ),
    .A2(net83),
    .Y(_1660_),
    .B1(_1659_));
 sg13g2_nor2_1 _4411_ (.A(_1846_),
    .B(net58),
    .Y(_1661_));
 sg13g2_a21oi_1 _4412_ (.A1(net57),
    .A2(_1660_),
    .Y(_0160_),
    .B1(_1661_));
 sg13g2_nor2b_1 _4413_ (.A(net84),
    .B_N(\lfsr0.seed_reg[19] ),
    .Y(_1662_));
 sg13g2_a21oi_1 _4414_ (.A1(_1846_),
    .A2(net83),
    .Y(_1663_),
    .B1(_1662_));
 sg13g2_nor2_1 _4415_ (.A(\lfsr0.lfsr_out[19] ),
    .B(net58),
    .Y(_1664_));
 sg13g2_a21oi_1 _4416_ (.A1(net57),
    .A2(_1663_),
    .Y(_0161_),
    .B1(_1664_));
 sg13g2_nor2b_1 _4417_ (.A(net84),
    .B_N(\lfsr0.seed_reg[1] ),
    .Y(_1665_));
 sg13g2_a21oi_1 _4418_ (.A1(\lfsr0.lfsr_out[0] ),
    .A2(net83),
    .Y(_1666_),
    .B1(_1665_));
 sg13g2_nor2_1 _4419_ (.A(\lfsr0.lfsr_out[1] ),
    .B(net58),
    .Y(_1667_));
 sg13g2_a21oi_1 _4420_ (.A1(net57),
    .A2(_1666_),
    .Y(_0162_),
    .B1(_1667_));
 sg13g2_nor2b_1 _4421_ (.A(net84),
    .B_N(\lfsr0.seed_reg[20] ),
    .Y(_1668_));
 sg13g2_a21oi_1 _4422_ (.A1(\lfsr0.lfsr_out[19] ),
    .A2(net83),
    .Y(_1669_),
    .B1(_1668_));
 sg13g2_nor2_1 _4423_ (.A(\lfsr0.lfsr_out[20] ),
    .B(net58),
    .Y(_1670_));
 sg13g2_a21oi_1 _4424_ (.A1(net57),
    .A2(_1669_),
    .Y(_0163_),
    .B1(_1670_));
 sg13g2_nor2b_1 _4425_ (.A(net84),
    .B_N(\lfsr0.seed_reg[21] ),
    .Y(_1671_));
 sg13g2_a21oi_1 _4426_ (.A1(\lfsr0.lfsr_out[20] ),
    .A2(_1658_),
    .Y(_1672_),
    .B1(_1671_));
 sg13g2_nor2_1 _4427_ (.A(_1865_),
    .B(net58),
    .Y(_1673_));
 sg13g2_a21oi_1 _4428_ (.A1(_1657_),
    .A2(_1672_),
    .Y(_0164_),
    .B1(_1673_));
 sg13g2_nor2b_1 _4429_ (.A(net84),
    .B_N(\lfsr0.seed_reg[22] ),
    .Y(_1674_));
 sg13g2_a21oi_1 _4430_ (.A1(_1865_),
    .A2(_1658_),
    .Y(_1675_),
    .B1(_1674_));
 sg13g2_buf_1 _4431_ (.A(_1869_),
    .X(_1676_));
 sg13g2_nor2_1 _4432_ (.A(\lfsr0.lfsr_out[22] ),
    .B(net56),
    .Y(_1677_));
 sg13g2_a21oi_1 _4433_ (.A1(_1657_),
    .A2(_1675_),
    .Y(_0165_),
    .B1(_1677_));
 sg13g2_nor2b_1 _4434_ (.A(net94),
    .B_N(\lfsr0.seed_reg[23] ),
    .Y(_1678_));
 sg13g2_a21oi_1 _4435_ (.A1(\lfsr0.lfsr_out[22] ),
    .A2(net83),
    .Y(_1679_),
    .B1(_1678_));
 sg13g2_nor2_1 _4436_ (.A(\lfsr0.lfsr_out[23] ),
    .B(net56),
    .Y(_1680_));
 sg13g2_a21oi_1 _4437_ (.A1(net57),
    .A2(_1679_),
    .Y(_0166_),
    .B1(_1680_));
 sg13g2_nor2b_1 _4438_ (.A(net94),
    .B_N(\lfsr0.seed_reg[2] ),
    .Y(_1681_));
 sg13g2_a21oi_1 _4439_ (.A1(\lfsr0.lfsr_out[1] ),
    .A2(net83),
    .Y(_1682_),
    .B1(_1681_));
 sg13g2_nor2_1 _4440_ (.A(\lfsr0.lfsr_out[2] ),
    .B(net56),
    .Y(_1683_));
 sg13g2_a21oi_1 _4441_ (.A1(net57),
    .A2(_1682_),
    .Y(_0167_),
    .B1(_1683_));
 sg13g2_nor2b_1 _4442_ (.A(net94),
    .B_N(\lfsr0.seed_reg[3] ),
    .Y(_1684_));
 sg13g2_a21oi_1 _4443_ (.A1(\lfsr0.lfsr_out[2] ),
    .A2(net83),
    .Y(_1685_),
    .B1(_1684_));
 sg13g2_nor2_1 _4444_ (.A(_1835_),
    .B(_1676_),
    .Y(_1686_));
 sg13g2_a21oi_1 _4445_ (.A1(net57),
    .A2(_1685_),
    .Y(_0168_),
    .B1(_1686_));
 sg13g2_nor2b_1 _4446_ (.A(net94),
    .B_N(\lfsr0.seed_reg[4] ),
    .Y(_1687_));
 sg13g2_a21oi_1 _4447_ (.A1(_1835_),
    .A2(net83),
    .Y(_1688_),
    .B1(_1687_));
 sg13g2_nor2_1 _4448_ (.A(_1828_),
    .B(net56),
    .Y(_1689_));
 sg13g2_a21oi_1 _4449_ (.A1(net57),
    .A2(_1688_),
    .Y(_0169_),
    .B1(_1689_));
 sg13g2_nor2b_1 _4450_ (.A(net94),
    .B_N(\lfsr0.seed_reg[5] ),
    .Y(_1690_));
 sg13g2_a21oi_1 _4451_ (.A1(_1828_),
    .A2(net85),
    .Y(_1691_),
    .B1(_1690_));
 sg13g2_nor2_1 _4452_ (.A(net117),
    .B(net56),
    .Y(_1692_));
 sg13g2_a21oi_1 _4453_ (.A1(net63),
    .A2(_1691_),
    .Y(_0170_),
    .B1(_1692_));
 sg13g2_nor2b_1 _4454_ (.A(_1872_),
    .B_N(\lfsr0.seed_reg[6] ),
    .Y(_1693_));
 sg13g2_a21oi_1 _4455_ (.A1(_1850_),
    .A2(net85),
    .Y(_1694_),
    .B1(_1693_));
 sg13g2_nor2_1 _4456_ (.A(net119),
    .B(net56),
    .Y(_1695_));
 sg13g2_a21oi_1 _4457_ (.A1(net63),
    .A2(_1694_),
    .Y(_0171_),
    .B1(_1695_));
 sg13g2_nor2b_1 _4458_ (.A(_1872_),
    .B_N(\lfsr0.seed_reg[7] ),
    .Y(_1696_));
 sg13g2_a21oi_1 _4459_ (.A1(_1839_),
    .A2(net85),
    .Y(_1697_),
    .B1(_1696_));
 sg13g2_nor2_1 _4460_ (.A(net116),
    .B(_1676_),
    .Y(_1698_));
 sg13g2_a21oi_1 _4461_ (.A1(net63),
    .A2(_1697_),
    .Y(_0172_),
    .B1(_1698_));
 sg13g2_nor2b_1 _4462_ (.A(net94),
    .B_N(\lfsr0.seed_reg[8] ),
    .Y(_1699_));
 sg13g2_a21oi_1 _4463_ (.A1(_1853_),
    .A2(_1627_),
    .Y(_1700_),
    .B1(_1699_));
 sg13g2_nor2_1 _4464_ (.A(\lfsr0.lfsr_out[8] ),
    .B(net56),
    .Y(_1701_));
 sg13g2_a21oi_1 _4465_ (.A1(net63),
    .A2(_1700_),
    .Y(_0173_),
    .B1(_1701_));
 sg13g2_nor2b_1 _4466_ (.A(net94),
    .B_N(\lfsr0.seed_reg[9] ),
    .Y(_1702_));
 sg13g2_a21oi_1 _4467_ (.A1(\lfsr0.lfsr_out[8] ),
    .A2(net85),
    .Y(_1703_),
    .B1(_1702_));
 sg13g2_nor2_1 _4468_ (.A(_1831_),
    .B(net56),
    .Y(_1704_));
 sg13g2_a21oi_1 _4469_ (.A1(_1874_),
    .A2(_1703_),
    .Y(_0174_),
    .B1(_1704_));
 sg13g2_nor2b_1 _4470_ (.A(\spi0.rxtx_done_reg ),
    .B_N(\spi0.rxtx_done ),
    .Y(_1705_));
 sg13g2_buf_2 _4471_ (.A(_1705_),
    .X(_1706_));
 sg13g2_buf_1 _4472_ (.A(_1706_),
    .X(\spi0.rxtx_done_rising ));
 sg13g2_mux2_1 _4473_ (.A0(\input_data[0] ),
    .A1(\spi0.spi0.data_rx_o[16] ),
    .S(net73),
    .X(_0223_));
 sg13g2_mux2_1 _4474_ (.A0(_2027_),
    .A1(\spi0.spi0.data_rx_o[10] ),
    .S(net73),
    .X(_0224_));
 sg13g2_mux2_1 _4475_ (.A0(_2018_),
    .A1(\spi0.spi0.data_rx_o[11] ),
    .S(net73),
    .X(_0225_));
 sg13g2_mux2_1 _4476_ (.A0(net114),
    .A1(\spi0.spi0.data_rx_o[12] ),
    .S(net73),
    .X(_0226_));
 sg13g2_mux2_1 _4477_ (.A0(_2042_),
    .A1(\spi0.spi0.data_rx_o[13] ),
    .S(net73),
    .X(_0227_));
 sg13g2_mux2_1 _4478_ (.A0(_1980_),
    .A1(\spi0.spi0.data_rx_o[14] ),
    .S(net73),
    .X(_0228_));
 sg13g2_mux2_1 _4479_ (.A0(_2076_),
    .A1(\spi0.spi0.data_rx_o[15] ),
    .S(net73),
    .X(_0229_));
 sg13g2_mux2_1 _4480_ (.A0(\input_data[16] ),
    .A1(\spi0.spi0.data_rx_o[0] ),
    .S(\spi0.rxtx_done_rising ),
    .X(_0230_));
 sg13g2_mux2_1 _4481_ (.A0(\input_data[17] ),
    .A1(\spi0.spi0.data_rx_o[1] ),
    .S(net73),
    .X(_0231_));
 sg13g2_buf_1 _4482_ (.A(_1706_),
    .X(_1707_));
 sg13g2_mux2_1 _4483_ (.A0(_1958_),
    .A1(\spi0.spi0.data_rx_o[2] ),
    .S(net72),
    .X(_0232_));
 sg13g2_mux2_1 _4484_ (.A0(_1990_),
    .A1(\spi0.spi0.data_rx_o[3] ),
    .S(net72),
    .X(_0233_));
 sg13g2_mux2_1 _4485_ (.A0(\input_data[1] ),
    .A1(\spi0.spi0.data_rx_o[17] ),
    .S(net72),
    .X(_0234_));
 sg13g2_mux2_1 _4486_ (.A0(_2008_),
    .A1(\spi0.spi0.data_rx_o[4] ),
    .S(net72),
    .X(_0235_));
 sg13g2_mux2_1 _4487_ (.A0(_1959_),
    .A1(\spi0.spi0.data_rx_o[5] ),
    .S(net72),
    .X(_0236_));
 sg13g2_mux2_1 _4488_ (.A0(_1986_),
    .A1(\spi0.spi0.data_rx_o[6] ),
    .S(_1707_),
    .X(_0237_));
 sg13g2_mux2_1 _4489_ (.A0(_2005_),
    .A1(\spi0.spi0.data_rx_o[7] ),
    .S(_1707_),
    .X(_0238_));
 sg13g2_mux2_1 _4490_ (.A0(\input_data[2] ),
    .A1(\spi0.spi0.data_rx_o[18] ),
    .S(net72),
    .X(_0239_));
 sg13g2_mux2_1 _4491_ (.A0(\input_data[3] ),
    .A1(\spi0.spi0.data_rx_o[19] ),
    .S(net72),
    .X(_0240_));
 sg13g2_mux2_1 _4492_ (.A0(_1966_),
    .A1(\spi0.spi0.data_rx_o[20] ),
    .S(net72),
    .X(_0241_));
 sg13g2_mux2_1 _4493_ (.A0(net115),
    .A1(\spi0.spi0.data_rx_o[21] ),
    .S(_1706_),
    .X(_0242_));
 sg13g2_mux2_1 _4494_ (.A0(net113),
    .A1(\spi0.spi0.data_rx_o[22] ),
    .S(_1706_),
    .X(_0243_));
 sg13g2_mux2_1 _4495_ (.A0(net112),
    .A1(\spi0.spi0.data_rx_o[23] ),
    .S(_1706_),
    .X(_0244_));
 sg13g2_mux2_1 _4496_ (.A0(\input_data[8] ),
    .A1(\spi0.spi0.data_rx_o[8] ),
    .S(_1706_),
    .X(_0245_));
 sg13g2_mux2_1 _4497_ (.A0(_1975_),
    .A1(\spi0.spi0.data_rx_o[9] ),
    .S(_1706_),
    .X(_0246_));
 sg13g2_buf_1 _4498_ (.A(net59),
    .X(_1708_));
 sg13g2_buf_1 _4499_ (.A(\lfsr0.config_i ),
    .X(_1709_));
 sg13g2_buf_1 _4500_ (.A(_1709_),
    .X(_1710_));
 sg13g2_buf_1 _4501_ (.A(_1709_),
    .X(_1711_));
 sg13g2_nand2b_1 _4502_ (.Y(_1712_),
    .B(net81),
    .A_N(\lfsr0.stop_reg[0] ));
 sg13g2_o21ai_1 _4503_ (.B1(_1712_),
    .Y(_1713_),
    .A1(net82),
    .A2(\lfsr0.seed_reg[0] ));
 sg13g2_buf_1 _4504_ (.A(net5),
    .X(_1714_));
 sg13g2_buf_1 _4505_ (.A(net164),
    .X(_1715_));
 sg13g2_nand2_1 _4506_ (.Y(_1716_),
    .A(_1714_),
    .B(_1447_));
 sg13g2_o21ai_1 _4507_ (.B1(_1716_),
    .Y(net13),
    .A1(_1715_),
    .A2(_0359_));
 sg13g2_nor2_1 _4508_ (.A(_1973_),
    .B(net13),
    .Y(_1717_));
 sg13g2_a21oi_1 _4509_ (.A1(net53),
    .A2(_1713_),
    .Y(_1718_),
    .B1(_1717_));
 sg13g2_nor2b_1 _4510_ (.A(net164),
    .B_N(\gray_sobel0.px_rdy_o_sobel ),
    .Y(_1719_));
 sg13g2_a21oi_1 _4511_ (.A1(net164),
    .A2(_1946_),
    .Y(_1720_),
    .B1(_1719_));
 sg13g2_nand2_1 _4512_ (.Y(_1721_),
    .A(net59),
    .B(\lfsr0.config_done_o ));
 sg13g2_o21ai_1 _4513_ (.B1(_1721_),
    .Y(_1722_),
    .A1(net59),
    .A2(_1720_));
 sg13g2_buf_1 _4514_ (.A(_1722_),
    .X(_1723_));
 sg13g2_buf_1 _4515_ (.A(_1723_),
    .X(_1724_));
 sg13g2_mux2_1 _4516_ (.A0(\spi0.data_tx[0] ),
    .A1(_1718_),
    .S(net43),
    .X(_0247_));
 sg13g2_buf_1 _4517_ (.A(_1723_),
    .X(_1725_));
 sg13g2_nand2_1 _4518_ (.Y(_1726_),
    .A(net164),
    .B(_1443_));
 sg13g2_nor2_1 _4519_ (.A(net59),
    .B(_1726_),
    .Y(_1727_));
 sg13g2_buf_2 _4520_ (.A(_1727_),
    .X(_1728_));
 sg13g2_buf_1 _4521_ (.A(_1728_),
    .X(_1729_));
 sg13g2_mux2_1 _4522_ (.A0(\lfsr0.seed_reg[10] ),
    .A1(\lfsr0.stop_reg[10] ),
    .S(_1710_),
    .X(_1730_));
 sg13g2_buf_1 _4523_ (.A(net59),
    .X(_1731_));
 sg13g2_a22oi_1 _4524_ (.Y(_1732_),
    .B1(_1730_),
    .B2(net52),
    .A2(net44),
    .A1(_2027_));
 sg13g2_buf_1 _4525_ (.A(_1723_),
    .X(_1733_));
 sg13g2_nor2_1 _4526_ (.A(\spi0.data_tx[10] ),
    .B(net41),
    .Y(_1734_));
 sg13g2_a21oi_1 _4527_ (.A1(net42),
    .A2(_1732_),
    .Y(_0248_),
    .B1(_1734_));
 sg13g2_mux2_1 _4528_ (.A0(\lfsr0.seed_reg[11] ),
    .A1(\lfsr0.stop_reg[11] ),
    .S(net82),
    .X(_1735_));
 sg13g2_a22oi_1 _4529_ (.Y(_1736_),
    .B1(_1735_),
    .B2(net52),
    .A2(net44),
    .A1(_2018_));
 sg13g2_nor2_1 _4530_ (.A(\spi0.data_tx[11] ),
    .B(net41),
    .Y(_1737_));
 sg13g2_a21oi_1 _4531_ (.A1(net42),
    .A2(_1736_),
    .Y(_0249_),
    .B1(_1737_));
 sg13g2_buf_1 _4532_ (.A(_1709_),
    .X(_1738_));
 sg13g2_mux2_1 _4533_ (.A0(\lfsr0.seed_reg[12] ),
    .A1(\lfsr0.stop_reg[12] ),
    .S(net80),
    .X(_1739_));
 sg13g2_a22oi_1 _4534_ (.Y(_1740_),
    .B1(_1739_),
    .B2(net52),
    .A2(net44),
    .A1(net114));
 sg13g2_nor2_1 _4535_ (.A(\spi0.data_tx[12] ),
    .B(net41),
    .Y(_1741_));
 sg13g2_a21oi_1 _4536_ (.A1(net42),
    .A2(_1740_),
    .Y(_0250_),
    .B1(_1741_));
 sg13g2_mux2_1 _4537_ (.A0(\lfsr0.seed_reg[13] ),
    .A1(\lfsr0.stop_reg[13] ),
    .S(net80),
    .X(_1742_));
 sg13g2_a22oi_1 _4538_ (.Y(_1743_),
    .B1(_1742_),
    .B2(net52),
    .A2(net44),
    .A1(_2042_));
 sg13g2_nor2_1 _4539_ (.A(\spi0.data_tx[13] ),
    .B(net41),
    .Y(_1744_));
 sg13g2_a21oi_1 _4540_ (.A1(net42),
    .A2(_1743_),
    .Y(_0251_),
    .B1(_1744_));
 sg13g2_mux2_1 _4541_ (.A0(\lfsr0.seed_reg[14] ),
    .A1(\lfsr0.stop_reg[14] ),
    .S(net80),
    .X(_1745_));
 sg13g2_a22oi_1 _4542_ (.Y(_1746_),
    .B1(_1745_),
    .B2(net52),
    .A2(net44),
    .A1(_1980_));
 sg13g2_nor2_1 _4543_ (.A(\spi0.data_tx[14] ),
    .B(_1733_),
    .Y(_1747_));
 sg13g2_a21oi_1 _4544_ (.A1(net42),
    .A2(_1746_),
    .Y(_0252_),
    .B1(_1747_));
 sg13g2_mux2_1 _4545_ (.A0(\lfsr0.seed_reg[15] ),
    .A1(\lfsr0.stop_reg[15] ),
    .S(_1738_),
    .X(_1748_));
 sg13g2_a22oi_1 _4546_ (.Y(_1749_),
    .B1(_1748_),
    .B2(net52),
    .A2(net44),
    .A1(_2076_));
 sg13g2_nor2_1 _4547_ (.A(\spi0.data_tx[15] ),
    .B(_1733_),
    .Y(_1750_));
 sg13g2_a21oi_1 _4548_ (.A1(net42),
    .A2(_1749_),
    .Y(_0253_),
    .B1(_1750_));
 sg13g2_mux2_1 _4549_ (.A0(\lfsr0.seed_reg[16] ),
    .A1(\lfsr0.stop_reg[16] ),
    .S(net80),
    .X(_1751_));
 sg13g2_a22oi_1 _4550_ (.Y(_1752_),
    .B1(_1751_),
    .B2(_1731_),
    .A2(_1729_),
    .A1(\input_data[16] ));
 sg13g2_buf_1 _4551_ (.A(_1723_),
    .X(_1753_));
 sg13g2_nor2_1 _4552_ (.A(\spi0.data_tx[16] ),
    .B(net40),
    .Y(_1754_));
 sg13g2_a21oi_1 _4553_ (.A1(net42),
    .A2(_1752_),
    .Y(_0254_),
    .B1(_1754_));
 sg13g2_mux2_1 _4554_ (.A0(\lfsr0.seed_reg[17] ),
    .A1(\lfsr0.stop_reg[17] ),
    .S(_1738_),
    .X(_1755_));
 sg13g2_a22oi_1 _4555_ (.Y(_1756_),
    .B1(_1755_),
    .B2(_1731_),
    .A2(_1729_),
    .A1(\input_data[17] ));
 sg13g2_nor2_1 _4556_ (.A(\spi0.data_tx[17] ),
    .B(net40),
    .Y(_1757_));
 sg13g2_a21oi_1 _4557_ (.A1(net42),
    .A2(_1756_),
    .Y(_0255_),
    .B1(_1757_));
 sg13g2_mux2_1 _4558_ (.A0(\lfsr0.seed_reg[18] ),
    .A1(\lfsr0.stop_reg[18] ),
    .S(net80),
    .X(_1758_));
 sg13g2_a22oi_1 _4559_ (.Y(_1759_),
    .B1(_1758_),
    .B2(net52),
    .A2(net44),
    .A1(_1958_));
 sg13g2_nor2_1 _4560_ (.A(\spi0.data_tx[18] ),
    .B(net40),
    .Y(_1760_));
 sg13g2_a21oi_1 _4561_ (.A1(_1725_),
    .A2(_1759_),
    .Y(_0256_),
    .B1(_1760_));
 sg13g2_mux2_1 _4562_ (.A0(\lfsr0.seed_reg[19] ),
    .A1(\lfsr0.stop_reg[19] ),
    .S(net80),
    .X(_1761_));
 sg13g2_a22oi_1 _4563_ (.Y(_1762_),
    .B1(_1761_),
    .B2(net52),
    .A2(net44),
    .A1(_1990_));
 sg13g2_nor2_1 _4564_ (.A(\spi0.data_tx[19] ),
    .B(net40),
    .Y(_1763_));
 sg13g2_a21oi_1 _4565_ (.A1(_1725_),
    .A2(_1762_),
    .Y(_0257_),
    .B1(_1763_));
 sg13g2_nand2b_1 _4566_ (.Y(_1764_),
    .B(net81),
    .A_N(\lfsr0.stop_reg[1] ));
 sg13g2_o21ai_1 _4567_ (.B1(_1764_),
    .Y(_1765_),
    .A1(net82),
    .A2(\lfsr0.seed_reg[1] ));
 sg13g2_nand2_1 _4568_ (.Y(_1766_),
    .A(net164),
    .B(_1493_));
 sg13g2_o21ai_1 _4569_ (.B1(_1766_),
    .Y(net14),
    .A1(net95),
    .A2(_1384_));
 sg13g2_nor2_1 _4570_ (.A(_1973_),
    .B(net14),
    .Y(_1767_));
 sg13g2_a21oi_1 _4571_ (.A1(net53),
    .A2(_1765_),
    .Y(_1768_),
    .B1(_1767_));
 sg13g2_mux2_1 _4572_ (.A0(\spi0.data_tx[1] ),
    .A1(_1768_),
    .S(net43),
    .X(_0258_));
 sg13g2_mux2_1 _4573_ (.A0(\lfsr0.seed_reg[20] ),
    .A1(\lfsr0.stop_reg[20] ),
    .S(net80),
    .X(_1769_));
 sg13g2_a22oi_1 _4574_ (.Y(_1770_),
    .B1(_1769_),
    .B2(net53),
    .A2(_1728_),
    .A1(_2008_));
 sg13g2_nor2_1 _4575_ (.A(\spi0.data_tx[20] ),
    .B(net40),
    .Y(_1771_));
 sg13g2_a21oi_1 _4576_ (.A1(net43),
    .A2(_1770_),
    .Y(_0259_),
    .B1(_1771_));
 sg13g2_mux2_1 _4577_ (.A0(\lfsr0.seed_reg[21] ),
    .A1(\lfsr0.stop_reg[21] ),
    .S(net80),
    .X(_1772_));
 sg13g2_a22oi_1 _4578_ (.Y(_1773_),
    .B1(_1772_),
    .B2(net53),
    .A2(_1728_),
    .A1(_1959_));
 sg13g2_nor2_1 _4579_ (.A(\spi0.data_tx[21] ),
    .B(_1753_),
    .Y(_1774_));
 sg13g2_a21oi_1 _4580_ (.A1(net43),
    .A2(_1773_),
    .Y(_0260_),
    .B1(_1774_));
 sg13g2_mux2_1 _4581_ (.A0(\lfsr0.seed_reg[22] ),
    .A1(\lfsr0.stop_reg[22] ),
    .S(net81),
    .X(_1775_));
 sg13g2_a22oi_1 _4582_ (.Y(_1776_),
    .B1(_1775_),
    .B2(net53),
    .A2(_1728_),
    .A1(_1986_));
 sg13g2_nor2_1 _4583_ (.A(\spi0.data_tx[22] ),
    .B(_1753_),
    .Y(_1777_));
 sg13g2_a21oi_1 _4584_ (.A1(net43),
    .A2(_1776_),
    .Y(_0261_),
    .B1(_1777_));
 sg13g2_mux2_1 _4585_ (.A0(\lfsr0.seed_reg[23] ),
    .A1(\lfsr0.stop_reg[23] ),
    .S(net81),
    .X(_1778_));
 sg13g2_a22oi_1 _4586_ (.Y(_1779_),
    .B1(_1778_),
    .B2(net53),
    .A2(_1728_),
    .A1(_2005_));
 sg13g2_nor2_1 _4587_ (.A(\spi0.data_tx[23] ),
    .B(net40),
    .Y(_1780_));
 sg13g2_a21oi_1 _4588_ (.A1(_1724_),
    .A2(_1779_),
    .Y(_0262_),
    .B1(_1780_));
 sg13g2_nand2b_1 _4589_ (.Y(_1781_),
    .B(net81),
    .A_N(\lfsr0.stop_reg[2] ));
 sg13g2_o21ai_1 _4590_ (.B1(_1781_),
    .Y(_1782_),
    .A1(net82),
    .A2(\lfsr0.seed_reg[2] ));
 sg13g2_nand2_1 _4591_ (.Y(_1783_),
    .A(_1714_),
    .B(_1452_));
 sg13g2_o21ai_1 _4592_ (.B1(_1783_),
    .Y(net15),
    .A1(_1715_),
    .A2(_1396_));
 sg13g2_nor2_1 _4593_ (.A(net55),
    .B(net15),
    .Y(_1784_));
 sg13g2_a21oi_1 _4594_ (.A1(_1708_),
    .A2(_1782_),
    .Y(_1785_),
    .B1(_1784_));
 sg13g2_mux2_1 _4595_ (.A0(\spi0.data_tx[2] ),
    .A1(_1785_),
    .S(net43),
    .X(_0263_));
 sg13g2_nand2b_1 _4596_ (.Y(_1786_),
    .B(net81),
    .A_N(\lfsr0.stop_reg[3] ));
 sg13g2_o21ai_1 _4597_ (.B1(_1786_),
    .Y(_1787_),
    .A1(net82),
    .A2(\lfsr0.seed_reg[3] ));
 sg13g2_nand2_1 _4598_ (.Y(_1788_),
    .A(net164),
    .B(_1462_));
 sg13g2_o21ai_1 _4599_ (.B1(_1788_),
    .Y(net16),
    .A1(net95),
    .A2(_1400_));
 sg13g2_nor2_1 _4600_ (.A(net55),
    .B(net16),
    .Y(_1789_));
 sg13g2_a21oi_1 _4601_ (.A1(_1708_),
    .A2(_1787_),
    .Y(_1790_),
    .B1(_1789_));
 sg13g2_mux2_1 _4602_ (.A0(\spi0.data_tx[3] ),
    .A1(_1790_),
    .S(net43),
    .X(_0264_));
 sg13g2_nand2b_1 _4603_ (.Y(_1791_),
    .B(net81),
    .A_N(\lfsr0.stop_reg[4] ));
 sg13g2_o21ai_1 _4604_ (.B1(_1791_),
    .Y(_1792_),
    .A1(net82),
    .A2(\lfsr0.seed_reg[4] ));
 sg13g2_nand2_1 _4605_ (.Y(_1793_),
    .A(net164),
    .B(_1466_));
 sg13g2_o21ai_1 _4606_ (.B1(_1793_),
    .Y(net17),
    .A1(net164),
    .A2(_1404_));
 sg13g2_nor2_1 _4607_ (.A(net55),
    .B(net17),
    .Y(_1794_));
 sg13g2_a21oi_1 _4608_ (.A1(net55),
    .A2(_1792_),
    .Y(_1795_),
    .B1(_1794_));
 sg13g2_mux2_1 _4609_ (.A0(\spi0.data_tx[4] ),
    .A1(_1795_),
    .S(net41),
    .X(_0265_));
 sg13g2_nand2b_1 _4610_ (.Y(_1796_),
    .B(net81),
    .A_N(\lfsr0.stop_reg[5] ));
 sg13g2_o21ai_1 _4611_ (.B1(_1796_),
    .Y(_1797_),
    .A1(net82),
    .A2(\lfsr0.seed_reg[5] ));
 sg13g2_nand2_1 _4612_ (.Y(_1798_),
    .A(net95),
    .B(_1470_));
 sg13g2_o21ai_1 _4613_ (.B1(_1798_),
    .Y(_1799_),
    .A1(net95),
    .A2(_1410_));
 sg13g2_nor2_1 _4614_ (.A(_1972_),
    .B(_1799_),
    .Y(_1800_));
 sg13g2_a21oi_1 _4615_ (.A1(net55),
    .A2(_1797_),
    .Y(_1801_),
    .B1(_1800_));
 sg13g2_mux2_1 _4616_ (.A0(\spi0.data_tx[5] ),
    .A1(_1801_),
    .S(net41),
    .X(_0266_));
 sg13g2_nand2b_1 _4617_ (.Y(_1802_),
    .B(_1709_),
    .A_N(\lfsr0.stop_reg[6] ));
 sg13g2_o21ai_1 _4618_ (.B1(_1802_),
    .Y(_1803_),
    .A1(_1710_),
    .A2(\lfsr0.seed_reg[6] ));
 sg13g2_nand2_1 _4619_ (.Y(_1804_),
    .A(net95),
    .B(_1474_));
 sg13g2_o21ai_1 _4620_ (.B1(_1804_),
    .Y(_1805_),
    .A1(net95),
    .A2(_1417_));
 sg13g2_nor2_1 _4621_ (.A(net59),
    .B(_1805_),
    .Y(_1806_));
 sg13g2_a21oi_1 _4622_ (.A1(net55),
    .A2(_1803_),
    .Y(_1807_),
    .B1(_1806_));
 sg13g2_mux2_1 _4623_ (.A0(\spi0.data_tx[6] ),
    .A1(_1807_),
    .S(net41),
    .X(_0267_));
 sg13g2_nand2b_1 _4624_ (.Y(_1808_),
    .B(_1709_),
    .A_N(\lfsr0.stop_reg[7] ));
 sg13g2_o21ai_1 _4625_ (.B1(_1808_),
    .Y(_1809_),
    .A1(net82),
    .A2(\lfsr0.seed_reg[7] ));
 sg13g2_nand2_1 _4626_ (.Y(_1810_),
    .A(net95),
    .B(_1478_));
 sg13g2_o21ai_1 _4627_ (.B1(_1810_),
    .Y(_1811_),
    .A1(net95),
    .A2(_1428_));
 sg13g2_nor2_1 _4628_ (.A(_1972_),
    .B(_1811_),
    .Y(_1812_));
 sg13g2_a21oi_1 _4629_ (.A1(net55),
    .A2(_1809_),
    .Y(_1813_),
    .B1(_1812_));
 sg13g2_mux2_1 _4630_ (.A0(\spi0.data_tx[7] ),
    .A1(_1813_),
    .S(net41),
    .X(_0268_));
 sg13g2_mux2_1 _4631_ (.A0(\lfsr0.seed_reg[8] ),
    .A1(\lfsr0.stop_reg[8] ),
    .S(_1711_),
    .X(_1814_));
 sg13g2_a22oi_1 _4632_ (.Y(_1815_),
    .B1(_1814_),
    .B2(net53),
    .A2(_1728_),
    .A1(\input_data[8] ));
 sg13g2_nor2_1 _4633_ (.A(\spi0.data_tx[8] ),
    .B(net40),
    .Y(_1816_));
 sg13g2_a21oi_1 _4634_ (.A1(_1724_),
    .A2(_1815_),
    .Y(_0269_),
    .B1(_1816_));
 sg13g2_mux2_1 _4635_ (.A0(\lfsr0.seed_reg[9] ),
    .A1(\lfsr0.stop_reg[9] ),
    .S(_1711_),
    .X(_1817_));
 sg13g2_a22oi_1 _4636_ (.Y(_1818_),
    .B1(_1817_),
    .B2(net53),
    .A2(_1728_),
    .A1(_1975_));
 sg13g2_nor2_1 _4637_ (.A(\spi0.data_tx[9] ),
    .B(net40),
    .Y(_1819_));
 sg13g2_a21oi_1 _4638_ (.A1(net43),
    .A2(_1818_),
    .Y(_0270_),
    .B1(_1819_));
 sg13g2_nor2b_1 _4639_ (.A(_1709_),
    .B_N(in_lfsr_rdy),
    .Y(_1820_));
 sg13g2_buf_2 _4640_ (.A(_1820_),
    .X(_1821_));
 sg13g2_buf_1 _4641_ (.A(_1821_),
    .X(_1822_));
 sg13g2_mux2_1 _4642_ (.A0(\lfsr0.seed_reg[0] ),
    .A1(\input_data[0] ),
    .S(net39),
    .X(_0175_));
 sg13g2_mux2_1 _4643_ (.A0(\lfsr0.seed_reg[10] ),
    .A1(_2027_),
    .S(net39),
    .X(_0176_));
 sg13g2_mux2_1 _4644_ (.A0(\lfsr0.seed_reg[11] ),
    .A1(_2018_),
    .S(net39),
    .X(_0177_));
 sg13g2_mux2_1 _4645_ (.A0(\lfsr0.seed_reg[12] ),
    .A1(_1976_),
    .S(_1822_),
    .X(_0178_));
 sg13g2_mux2_1 _4646_ (.A0(\lfsr0.seed_reg[13] ),
    .A1(_2042_),
    .S(net39),
    .X(_0179_));
 sg13g2_mux2_1 _4647_ (.A0(\lfsr0.seed_reg[14] ),
    .A1(_1980_),
    .S(net39),
    .X(_0180_));
 sg13g2_mux2_1 _4648_ (.A0(\lfsr0.seed_reg[15] ),
    .A1(_2076_),
    .S(net39),
    .X(_0181_));
 sg13g2_mux2_1 _4649_ (.A0(\lfsr0.seed_reg[16] ),
    .A1(\input_data[16] ),
    .S(net39),
    .X(_0182_));
 sg13g2_mux2_1 _4650_ (.A0(\lfsr0.seed_reg[17] ),
    .A1(\input_data[17] ),
    .S(_1822_),
    .X(_0183_));
 sg13g2_mux2_1 _4651_ (.A0(\lfsr0.seed_reg[18] ),
    .A1(_1958_),
    .S(net39),
    .X(_0184_));
 sg13g2_buf_1 _4652_ (.A(_1821_),
    .X(_1823_));
 sg13g2_mux2_1 _4653_ (.A0(\lfsr0.seed_reg[19] ),
    .A1(_1990_),
    .S(net38),
    .X(_0185_));
 sg13g2_mux2_1 _4654_ (.A0(\lfsr0.seed_reg[1] ),
    .A1(\input_data[1] ),
    .S(net38),
    .X(_0186_));
 sg13g2_mux2_1 _4655_ (.A0(\lfsr0.seed_reg[20] ),
    .A1(_2008_),
    .S(net38),
    .X(_0187_));
 sg13g2_mux2_1 _4656_ (.A0(\lfsr0.seed_reg[21] ),
    .A1(_1959_),
    .S(net38),
    .X(_0188_));
 sg13g2_mux2_1 _4657_ (.A0(\lfsr0.seed_reg[22] ),
    .A1(_1986_),
    .S(net38),
    .X(_0189_));
 sg13g2_mux2_1 _4658_ (.A0(\lfsr0.seed_reg[23] ),
    .A1(_2005_),
    .S(net38),
    .X(_0190_));
 sg13g2_mux2_1 _4659_ (.A0(\lfsr0.seed_reg[2] ),
    .A1(\input_data[2] ),
    .S(net38),
    .X(_0191_));
 sg13g2_mux2_1 _4660_ (.A0(\lfsr0.seed_reg[3] ),
    .A1(\input_data[3] ),
    .S(net38),
    .X(_0192_));
 sg13g2_mux2_1 _4661_ (.A0(\lfsr0.seed_reg[4] ),
    .A1(_1966_),
    .S(_1823_),
    .X(_0193_));
 sg13g2_mux2_1 _4662_ (.A0(\lfsr0.seed_reg[5] ),
    .A1(net115),
    .S(_1823_),
    .X(_0194_));
 sg13g2_mux2_1 _4663_ (.A0(\lfsr0.seed_reg[6] ),
    .A1(net113),
    .S(_1821_),
    .X(_0195_));
 sg13g2_mux2_1 _4664_ (.A0(\lfsr0.seed_reg[7] ),
    .A1(net112),
    .S(_1821_),
    .X(_0196_));
 sg13g2_mux2_1 _4665_ (.A0(\lfsr0.seed_reg[8] ),
    .A1(\input_data[8] ),
    .S(_1821_),
    .X(_0197_));
 sg13g2_mux2_1 _4666_ (.A0(\lfsr0.seed_reg[9] ),
    .A1(_1975_),
    .S(_1821_),
    .X(_0198_));
 sg13g2_nand2_1 _4667_ (.Y(_1824_),
    .A(_1709_),
    .B(in_lfsr_rdy));
 sg13g2_buf_2 _4668_ (.A(_1824_),
    .X(_1825_));
 sg13g2_buf_1 _4669_ (.A(_1825_),
    .X(_1826_));
 sg13g2_mux2_1 _4670_ (.A0(\input_data[0] ),
    .A1(\lfsr0.stop_reg[0] ),
    .S(net37),
    .X(_0199_));
 sg13g2_mux2_1 _4671_ (.A0(_2027_),
    .A1(\lfsr0.stop_reg[10] ),
    .S(net37),
    .X(_0200_));
 sg13g2_mux2_1 _4672_ (.A0(_2018_),
    .A1(\lfsr0.stop_reg[11] ),
    .S(net37),
    .X(_0201_));
 sg13g2_mux2_1 _4673_ (.A0(_1976_),
    .A1(\lfsr0.stop_reg[12] ),
    .S(net37),
    .X(_0202_));
 sg13g2_mux2_1 _4674_ (.A0(_2042_),
    .A1(\lfsr0.stop_reg[13] ),
    .S(net37),
    .X(_0203_));
 sg13g2_mux2_1 _4675_ (.A0(_1980_),
    .A1(\lfsr0.stop_reg[14] ),
    .S(net37),
    .X(_0204_));
 sg13g2_mux2_1 _4676_ (.A0(_2076_),
    .A1(\lfsr0.stop_reg[15] ),
    .S(net37),
    .X(_0205_));
 sg13g2_mux2_1 _4677_ (.A0(\input_data[16] ),
    .A1(\lfsr0.stop_reg[16] ),
    .S(_1826_),
    .X(_0206_));
 sg13g2_mux2_1 _4678_ (.A0(\input_data[17] ),
    .A1(\lfsr0.stop_reg[17] ),
    .S(_1826_),
    .X(_0207_));
 sg13g2_mux2_1 _4679_ (.A0(_1958_),
    .A1(\lfsr0.stop_reg[18] ),
    .S(net37),
    .X(_0208_));
 sg13g2_buf_1 _4680_ (.A(_1825_),
    .X(_1827_));
 sg13g2_mux2_1 _4681_ (.A0(_1990_),
    .A1(\lfsr0.stop_reg[19] ),
    .S(net36),
    .X(_0209_));
 sg13g2_mux2_1 _4682_ (.A0(\input_data[1] ),
    .A1(\lfsr0.stop_reg[1] ),
    .S(net36),
    .X(_0210_));
 sg13g2_mux2_1 _4683_ (.A0(_2008_),
    .A1(\lfsr0.stop_reg[20] ),
    .S(net36),
    .X(_0211_));
 sg13g2_mux2_1 _4684_ (.A0(_1959_),
    .A1(\lfsr0.stop_reg[21] ),
    .S(net36),
    .X(_0212_));
 sg13g2_mux2_1 _4685_ (.A0(_1986_),
    .A1(\lfsr0.stop_reg[22] ),
    .S(_1827_),
    .X(_0213_));
 sg13g2_mux2_1 _4686_ (.A0(_2005_),
    .A1(\lfsr0.stop_reg[23] ),
    .S(_1827_),
    .X(_0214_));
 sg13g2_mux2_1 _4687_ (.A0(\input_data[2] ),
    .A1(\lfsr0.stop_reg[2] ),
    .S(net36),
    .X(_0215_));
 sg13g2_mux2_1 _4688_ (.A0(\input_data[3] ),
    .A1(\lfsr0.stop_reg[3] ),
    .S(net36),
    .X(_0216_));
 sg13g2_mux2_1 _4689_ (.A0(_1966_),
    .A1(\lfsr0.stop_reg[4] ),
    .S(net36),
    .X(_0217_));
 sg13g2_mux2_1 _4690_ (.A0(_1967_),
    .A1(\lfsr0.stop_reg[5] ),
    .S(net36),
    .X(_0218_));
 sg13g2_mux2_1 _4691_ (.A0(_1997_),
    .A1(\lfsr0.stop_reg[6] ),
    .S(_1825_),
    .X(_0219_));
 sg13g2_mux2_1 _4692_ (.A0(_2013_),
    .A1(\lfsr0.stop_reg[7] ),
    .S(_1825_),
    .X(_0220_));
 sg13g2_mux2_1 _4693_ (.A0(\input_data[8] ),
    .A1(\lfsr0.stop_reg[8] ),
    .S(_1825_),
    .X(_0221_));
 sg13g2_mux2_1 _4694_ (.A0(_1975_),
    .A1(\lfsr0.stop_reg[9] ),
    .S(_1825_),
    .X(_0222_));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi \nreset_sync0.r_sync$_DFF_PN0__202  (.L_HI(net202));
 sg13g2_buf_1 _4697_ (.A(net186),
    .X(uio_oe[0]));
 sg13g2_buf_1 _4698_ (.A(net187),
    .X(uio_oe[1]));
 sg13g2_buf_1 _4699_ (.A(net188),
    .X(uio_oe[2]));
 sg13g2_buf_1 _4700_ (.A(net189),
    .X(uio_oe[3]));
 sg13g2_buf_1 _4701_ (.A(net190),
    .X(uio_oe[4]));
 sg13g2_buf_1 _4702_ (.A(net191),
    .X(uio_oe[5]));
 sg13g2_buf_1 _4703_ (.A(net192),
    .X(uio_oe[6]));
 sg13g2_buf_1 _4704_ (.A(net193),
    .X(uio_oe[7]));
 sg13g2_buf_1 _4705_ (.A(net194),
    .X(uio_out[0]));
 sg13g2_buf_1 _4706_ (.A(net195),
    .X(uio_out[1]));
 sg13g2_buf_1 _4707_ (.A(net196),
    .X(uio_out[2]));
 sg13g2_buf_1 _4708_ (.A(net197),
    .X(uio_out[3]));
 sg13g2_buf_1 _4709_ (.A(net198),
    .X(uio_out[4]));
 sg13g2_buf_1 _4710_ (.A(net199),
    .X(uio_out[5]));
 sg13g2_buf_1 _4711_ (.A(net200),
    .X(uio_out[6]));
 sg13g2_buf_1 _4712_ (.A(net201),
    .X(uio_out[7]));
 sg13g2_buf_1 _4713_ (.A(\spi0.spi0.sdo_o ),
    .X(net10));
 sg13g2_buf_1 _4714_ (.A(\lfsr0.lfsr_done ),
    .X(net11));
 sg13g2_buf_1 _4715_ (.A(ena),
    .X(net12));
 sg13g2_dfrbp_1 \gray_sobel0.gray_scale0.out_px_gray_o[0]$_DFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net132),
    .D(_0033_),
    .Q_N(_2470_),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.gray_scale0.out_px_gray_o[1]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net127),
    .D(_0034_),
    .Q_N(_2471_),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.gray_scale0.out_px_gray_o[2]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net127),
    .D(_0035_),
    .Q_N(_2472_),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.gray_scale0.out_px_gray_o[3]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net127),
    .D(_0036_),
    .Q_N(_2473_),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.gray_scale0.out_px_gray_o[4]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net127),
    .D(_0037_),
    .Q_N(_2474_),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.gray_scale0.out_px_gray_o[5]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net127),
    .D(_0038_),
    .Q_N(_2475_),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.gray_scale0.out_px_gray_o[6]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net128),
    .D(_0039_),
    .Q_N(_2476_),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.gray_scale0.out_px_gray_o[7]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net127),
    .D(_0040_),
    .Q_N(_2477_),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.gray_scale0.px_rdy_o$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net159),
    .D(\gray_sobel0.gray_scale0.px_rdy_i ),
    .Q_N(_2469_),
    .Q(\gray_sobel0.gray_scale0.px_rdy_o ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net141),
    .D(_0043_),
    .Q_N(_2468_),
    .Q(\gray_sobel0.sobel0.counter_pixels[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net146),
    .D(_0044_),
    .Q_N(_2467_),
    .Q(\gray_sobel0.sobel0.counter_pixels[10] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net147),
    .D(_0045_),
    .Q_N(_2466_),
    .Q(\gray_sobel0.sobel0.counter_pixels[11] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(_0046_),
    .Q_N(_2465_),
    .Q(\gray_sobel0.sobel0.counter_pixels[12] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net142),
    .D(_0047_),
    .Q_N(_2464_),
    .Q(\gray_sobel0.sobel0.counter_pixels[13] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net142),
    .D(_0048_),
    .Q_N(_2463_),
    .Q(\gray_sobel0.sobel0.counter_pixels[14] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net141),
    .D(_0049_),
    .Q_N(_2462_),
    .Q(\gray_sobel0.sobel0.counter_pixels[15] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net141),
    .D(_0050_),
    .Q_N(_2461_),
    .Q(\gray_sobel0.sobel0.counter_pixels[16] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net141),
    .D(_0051_),
    .Q_N(_2460_),
    .Q(\gray_sobel0.sobel0.counter_pixels[17] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net141),
    .D(_0052_),
    .Q_N(_2459_),
    .Q(\gray_sobel0.sobel0.counter_pixels[18] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net141),
    .D(_0053_),
    .Q_N(_2458_),
    .Q(\gray_sobel0.sobel0.counter_pixels[19] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net141),
    .D(_0054_),
    .Q_N(_2457_),
    .Q(\gray_sobel0.sobel0.counter_pixels[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net139),
    .D(_0055_),
    .Q_N(_2456_),
    .Q(\gray_sobel0.sobel0.counter_pixels[20] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net139),
    .D(_0056_),
    .Q_N(_2455_),
    .Q(\gray_sobel0.sobel0.counter_pixels[21] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net139),
    .D(_0057_),
    .Q_N(_2454_),
    .Q(\gray_sobel0.sobel0.counter_pixels[22] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net139),
    .D(_0058_),
    .Q_N(_2453_),
    .Q(\gray_sobel0.sobel0.counter_pixels[23] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net142),
    .D(_0059_),
    .Q_N(_2452_),
    .Q(\gray_sobel0.sobel0.counter_pixels[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net141),
    .D(_0060_),
    .Q_N(_2451_),
    .Q(\gray_sobel0.sobel0.counter_pixels[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net139),
    .D(_0061_),
    .Q_N(_2450_),
    .Q(\gray_sobel0.sobel0.counter_pixels[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net139),
    .D(_0062_),
    .Q_N(_2449_),
    .Q(\gray_sobel0.sobel0.counter_pixels[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net140),
    .D(_0063_),
    .Q_N(_2448_),
    .Q(\gray_sobel0.sobel0.counter_pixels[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net140),
    .D(_0064_),
    .Q_N(_2447_),
    .Q(\gray_sobel0.sobel0.counter_pixels[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net146),
    .D(_0065_),
    .Q_N(_2446_),
    .Q(\gray_sobel0.sobel0.counter_pixels[8] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_pixels[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net142),
    .D(_0066_),
    .Q_N(_2445_),
    .Q(\gray_sobel0.sobel0.counter_pixels[9] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_sobel[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(_0067_),
    .Q_N(_2444_),
    .Q(\gray_sobel0.sobel0.counter_sobel[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_sobel[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net158),
    .D(_0068_),
    .Q_N(_2443_),
    .Q(\gray_sobel0.sobel0.counter_sobel[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_sobel[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net158),
    .D(_0069_),
    .Q_N(_2442_),
    .Q(\gray_sobel0.sobel0.counter_sobel[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.counter_sobel[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net158),
    .D(_0070_),
    .Q_N(_2478_),
    .Q(\gray_sobel0.sobel0.counter_sobel[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.fsm_state[0]$_DFF_PN0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(net62),
    .Q_N(_2479_),
    .Q(\gray_sobel0.sobel0.fsm_state[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.fsm_state[1]$_DFF_PN0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net147),
    .D(\gray_sobel0.sobel0.next[1] ),
    .Q_N(_2441_),
    .Q(\gray_sobel0.sobel0.fsm_state[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.out_sobel[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net157),
    .D(_0071_),
    .Q_N(_2440_),
    .Q(\gray_sobel0.out_px_sobel[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.out_sobel[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net150),
    .D(_0072_),
    .Q_N(_2439_),
    .Q(\gray_sobel0.out_px_sobel[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.out_sobel[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net157),
    .D(_0073_),
    .Q_N(_2438_),
    .Q(\gray_sobel0.out_px_sobel[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.out_sobel[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net150),
    .D(_0074_),
    .Q_N(_2437_),
    .Q(\gray_sobel0.out_px_sobel[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.out_sobel[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net148),
    .D(_0075_),
    .Q_N(_2436_),
    .Q(\gray_sobel0.out_px_sobel[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.out_sobel[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net139),
    .D(_0076_),
    .Q_N(_2435_),
    .Q(\gray_sobel0.out_px_sobel[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.out_sobel[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net148),
    .D(_0077_),
    .Q_N(_2434_),
    .Q(\gray_sobel0.out_px_sobel[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.out_sobel[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net148),
    .D(_0078_),
    .Q_N(_2480_),
    .Q(\gray_sobel0.out_px_sobel[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.px_rdy_o$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net157),
    .D(\gray_sobel0.sobel0.px_ready ),
    .Q_N(_2481_),
    .Q(\gray_sobel0.px_rdy_o_sobel ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.px_ready$_DFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net157),
    .D(_0001_),
    .Q_N(_2433_),
    .Q(\gray_sobel0.sobel0.px_ready ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net132),
    .D(_0079_),
    .Q_N(_2432_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_2[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net150),
    .D(_0080_),
    .Q_N(_2431_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_1[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net148),
    .D(_0081_),
    .Q_N(_2430_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_1[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net148),
    .D(_0082_),
    .Q_N(_2429_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_1[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net144),
    .D(_0083_),
    .Q_N(_2428_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_1[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net148),
    .D(_0084_),
    .Q_N(_2427_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_1[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net140),
    .D(_0085_),
    .Q_N(_2426_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_1[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net132),
    .D(_0086_),
    .Q_N(_2425_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_0[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net132),
    .D(_0087_),
    .Q_N(_2424_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_0[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net127),
    .D(_0088_),
    .Q_N(_2423_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_0[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net125),
    .D(_0089_),
    .Q_N(_2422_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_0[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net132),
    .D(_0090_),
    .Q_N(_2421_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_2[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net127),
    .D(_0091_),
    .Q_N(_2420_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_0[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net120),
    .D(_0092_),
    .Q_N(_2419_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_0[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net122),
    .D(_0093_),
    .Q_N(_2418_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_0[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net122),
    .D(_0094_),
    .Q_N(_2417_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_0[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net123),
    .D(_0095_),
    .Q_N(_2416_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_2[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net123),
    .D(_0096_),
    .Q_N(_2415_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_2[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net121),
    .D(_0097_),
    .Q_N(_2414_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_2[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net121),
    .D(_0098_),
    .Q_N(_2413_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_2[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net124),
    .D(_0099_),
    .Q_N(_2412_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_2[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net120),
    .D(_0100_),
    .Q_N(_2411_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_2[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net125),
    .D(_0101_),
    .Q_N(_2410_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_2[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net122),
    .D(_0102_),
    .Q_N(_2409_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_2[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net123),
    .D(_0103_),
    .Q_N(_2408_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_2[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[32]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0104_),
    .Q_N(_2407_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_1[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[33]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net144),
    .D(_0105_),
    .Q_N(_2406_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_1[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[34]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0106_),
    .Q_N(_2405_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_1[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[35]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net144),
    .D(_0107_),
    .Q_N(_2404_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_1[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[36]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net144),
    .D(_0108_),
    .Q_N(_2403_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_1[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[37]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net146),
    .D(_0109_),
    .Q_N(_2402_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_1[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[38]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net144),
    .D(_0110_),
    .Q_N(_2401_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_1[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[39]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net144),
    .D(_0111_),
    .Q_N(_2400_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_1[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net125),
    .D(_0112_),
    .Q_N(_2399_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_2[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[40]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net123),
    .D(_0113_),
    .Q_N(_2398_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_0[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[41]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net123),
    .D(_0114_),
    .Q_N(_2397_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_0[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[42]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net121),
    .D(_0115_),
    .Q_N(_2396_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_0[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[43]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net121),
    .D(_0116_),
    .Q_N(_2395_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_0[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[44]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net124),
    .D(_0117_),
    .Q_N(_2394_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_0[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[45]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net120),
    .D(_0118_),
    .Q_N(_2393_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_0[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[46]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net122),
    .D(_0119_),
    .Q_N(_2392_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_0[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[47]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net123),
    .D(_0120_),
    .Q_N(_2391_),
    .Q(\gray_sobel0.sobel0.sobel.pix1_0[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[48]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net134),
    .D(_0121_),
    .Q_N(_2390_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_2[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[49]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net134),
    .D(_0122_),
    .Q_N(_2389_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_2[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net121),
    .D(_0123_),
    .Q_N(_2388_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_2[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[50]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net125),
    .D(_0124_),
    .Q_N(_2387_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_2[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[51]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net121),
    .D(_0125_),
    .Q_N(_2386_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_2[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[52]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net120),
    .D(_0126_),
    .Q_N(_2385_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_2[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[53]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net120),
    .D(_0127_),
    .Q_N(_2384_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_2[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[54]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net122),
    .D(_0128_),
    .Q_N(_2383_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_2[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[55]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net123),
    .D(_0129_),
    .Q_N(_2382_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_2[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[56]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0130_),
    .Q_N(_2381_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_1[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[57]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0131_),
    .Q_N(_2380_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_1[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[58]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0132_),
    .Q_N(_2379_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_1[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[59]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net145),
    .D(_0133_),
    .Q_N(_2378_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_1[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net120),
    .D(_0134_),
    .Q_N(_2377_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_2[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[60]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net144),
    .D(_0135_),
    .Q_N(_2376_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_1[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[61]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net144),
    .D(_0136_),
    .Q_N(_2375_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_1[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[62]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net139),
    .D(_0137_),
    .Q_N(_2374_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_1[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[63]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net140),
    .D(_0138_),
    .Q_N(_2373_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_1[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[64]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net134),
    .D(_0139_),
    .Q_N(_2372_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_0[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[65]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net134),
    .D(_0140_),
    .Q_N(_2371_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_0[1] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[66]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net125),
    .D(_0141_),
    .Q_N(_2370_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_0[2] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[67]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net121),
    .D(_0142_),
    .Q_N(_2369_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_0[3] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[68]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net120),
    .D(_0143_),
    .Q_N(_2368_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_0[4] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[69]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net120),
    .D(_0144_),
    .Q_N(_2367_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_0[5] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net122),
    .D(_0145_),
    .Q_N(_2366_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_2[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[70]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net122),
    .D(_0146_),
    .Q_N(_2365_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_0[6] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[71]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net122),
    .D(_0147_),
    .Q_N(_2364_),
    .Q(\gray_sobel0.sobel0.sobel.pix0_0[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net148),
    .D(_0148_),
    .Q_N(_2363_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_2[7] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net157),
    .D(_0149_),
    .Q_N(_2362_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_1[0] ));
 sg13g2_dfrbp_1 \gray_sobel0.sobel0.sobel_pixels[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net150),
    .D(_0150_),
    .Q_N(_2482_),
    .Q(\gray_sobel0.sobel0.sobel.pix2_1[1] ));
 sg13g2_dfrbp_1 \lfsr0.config_done_o$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net159),
    .D(in_lfsr_rdy),
    .Q_N(_2361_),
    .Q(\lfsr0.config_done_o ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net151),
    .D(_0151_),
    .Q_N(_2360_),
    .Q(\lfsr0.lfsr_out[0] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net149),
    .D(_0152_),
    .Q_N(_2359_),
    .Q(\lfsr0.lfsr_out[10] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net152),
    .D(_0153_),
    .Q_N(_2358_),
    .Q(\lfsr0.lfsr_out[11] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net152),
    .D(_0154_),
    .Q_N(_2357_),
    .Q(\lfsr0.lfsr_out[12] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net152),
    .D(_0155_),
    .Q_N(_2356_),
    .Q(\lfsr0.lfsr_out[13] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net152),
    .D(_0156_),
    .Q_N(_2355_),
    .Q(\lfsr0.lfsr_out[14] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net153),
    .D(_0157_),
    .Q_N(_2354_),
    .Q(\lfsr0.lfsr_out[15] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net152),
    .D(_0158_),
    .Q_N(_2353_),
    .Q(\lfsr0.lfsr_out[16] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net152),
    .D(_0159_),
    .Q_N(_2352_),
    .Q(\lfsr0.lfsr_out[17] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net136),
    .D(_0160_),
    .Q_N(_2351_),
    .Q(\lfsr0.lfsr_out[18] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net137),
    .D(_0161_),
    .Q_N(_2350_),
    .Q(\lfsr0.lfsr_out[19] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net133),
    .D(_0162_),
    .Q_N(_2349_),
    .Q(\lfsr0.lfsr_out[1] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net135),
    .D(_0163_),
    .Q_N(_2348_),
    .Q(\lfsr0.lfsr_out[20] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net135),
    .D(_0164_),
    .Q_N(_2347_),
    .Q(\lfsr0.lfsr_out[21] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net135),
    .D(_0165_),
    .Q_N(_2346_),
    .Q(\lfsr0.lfsr_out[22] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net135),
    .D(_0166_),
    .Q_N(_2345_),
    .Q(\lfsr0.lfsr_out[23] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net134),
    .D(_0167_),
    .Q_N(_2344_),
    .Q(\lfsr0.lfsr_out[2] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net151),
    .D(_0168_),
    .Q_N(_2343_),
    .Q(\lfsr0.lfsr_out[3] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net133),
    .D(_0169_),
    .Q_N(_2342_),
    .Q(\lfsr0.lfsr_out[4] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net149),
    .D(_0170_),
    .Q_N(_2341_),
    .Q(\lfsr0.lfsr_out[5] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net149),
    .D(_0171_),
    .Q_N(_2340_),
    .Q(\lfsr0.lfsr_out[6] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net151),
    .D(_0172_),
    .Q_N(_2339_),
    .Q(\lfsr0.lfsr_out[7] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net152),
    .D(_0173_),
    .Q_N(_2338_),
    .Q(\lfsr0.lfsr_out[8] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_out[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net149),
    .D(_0174_),
    .Q_N(_2483_),
    .Q(\lfsr0.lfsr_out[9] ));
 sg13g2_dfrbp_1 \lfsr0.lfsr_rdy_o$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net151),
    .D(_0000_),
    .Q_N(_2337_),
    .Q(\lfsr0.lfsr_rdy_o ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net133),
    .D(_0175_),
    .Q_N(_2336_),
    .Q(\lfsr0.seed_reg[0] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net154),
    .D(_0176_),
    .Q_N(_2335_),
    .Q(\lfsr0.seed_reg[10] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net136),
    .D(_0177_),
    .Q_N(_2334_),
    .Q(\lfsr0.seed_reg[11] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net154),
    .D(_0178_),
    .Q_N(_2333_),
    .Q(\lfsr0.seed_reg[12] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net154),
    .D(_0179_),
    .Q_N(_2332_),
    .Q(\lfsr0.seed_reg[13] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net153),
    .D(_0180_),
    .Q_N(_2331_),
    .Q(\lfsr0.seed_reg[14] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net153),
    .D(_0181_),
    .Q_N(_2330_),
    .Q(\lfsr0.seed_reg[15] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net155),
    .D(_0182_),
    .Q_N(_2329_),
    .Q(\lfsr0.seed_reg[16] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net153),
    .D(_0183_),
    .Q_N(_2328_),
    .Q(\lfsr0.seed_reg[17] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net136),
    .D(_0184_),
    .Q_N(_2327_),
    .Q(\lfsr0.seed_reg[18] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net135),
    .D(_0185_),
    .Q_N(_2326_),
    .Q(\lfsr0.seed_reg[19] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net133),
    .D(_0186_),
    .Q_N(_2325_),
    .Q(\lfsr0.seed_reg[1] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net135),
    .D(_0187_),
    .Q_N(_2324_),
    .Q(\lfsr0.seed_reg[20] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net135),
    .D(_0188_),
    .Q_N(_2323_),
    .Q(\lfsr0.seed_reg[21] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net137),
    .D(_0189_),
    .Q_N(_2322_),
    .Q(\lfsr0.seed_reg[22] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net135),
    .D(_0190_),
    .Q_N(_2321_),
    .Q(\lfsr0.seed_reg[23] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net134),
    .D(_0191_),
    .Q_N(_2320_),
    .Q(\lfsr0.seed_reg[2] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net149),
    .D(_0192_),
    .Q_N(_2319_),
    .Q(\lfsr0.seed_reg[3] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net132),
    .D(_0193_),
    .Q_N(_2318_),
    .Q(\lfsr0.seed_reg[4] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net149),
    .D(_0194_),
    .Q_N(_2317_),
    .Q(\lfsr0.seed_reg[5] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net150),
    .D(_0195_),
    .Q_N(_2316_),
    .Q(\lfsr0.seed_reg[6] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net150),
    .D(_0196_),
    .Q_N(_2315_),
    .Q(\lfsr0.seed_reg[7] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net154),
    .D(_0197_),
    .Q_N(_2314_),
    .Q(\lfsr0.seed_reg[8] ));
 sg13g2_dfrbp_1 \lfsr0.seed_reg[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net159),
    .D(_0198_),
    .Q_N(_2313_),
    .Q(\lfsr0.seed_reg[9] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net133),
    .D(_0199_),
    .Q_N(_2312_),
    .Q(\lfsr0.stop_reg[0] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net154),
    .D(_0200_),
    .Q_N(_2311_),
    .Q(\lfsr0.stop_reg[10] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net136),
    .D(_0201_),
    .Q_N(_2310_),
    .Q(\lfsr0.stop_reg[11] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net154),
    .D(_0202_),
    .Q_N(_2309_),
    .Q(\lfsr0.stop_reg[12] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net155),
    .D(_0203_),
    .Q_N(_2308_),
    .Q(\lfsr0.stop_reg[13] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net136),
    .D(_0204_),
    .Q_N(_2307_),
    .Q(\lfsr0.stop_reg[14] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net153),
    .D(_0205_),
    .Q_N(_2306_),
    .Q(\lfsr0.stop_reg[15] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net155),
    .D(_0206_),
    .Q_N(_2305_),
    .Q(\lfsr0.stop_reg[16] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net152),
    .D(_0207_),
    .Q_N(_2304_),
    .Q(\lfsr0.stop_reg[17] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net136),
    .D(_0208_),
    .Q_N(_2303_),
    .Q(\lfsr0.stop_reg[18] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net137),
    .D(_0209_),
    .Q_N(_2302_),
    .Q(\lfsr0.stop_reg[19] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net133),
    .D(_0210_),
    .Q_N(_2301_),
    .Q(\lfsr0.stop_reg[1] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net137),
    .D(_0211_),
    .Q_N(_2300_),
    .Q(\lfsr0.stop_reg[20] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net137),
    .D(_0212_),
    .Q_N(_2299_),
    .Q(\lfsr0.stop_reg[21] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net136),
    .D(_0213_),
    .Q_N(_2298_),
    .Q(\lfsr0.stop_reg[22] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net136),
    .D(_0214_),
    .Q_N(_2297_),
    .Q(\lfsr0.stop_reg[23] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net132),
    .D(_0215_),
    .Q_N(_2296_),
    .Q(\lfsr0.stop_reg[2] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net149),
    .D(_0216_),
    .Q_N(_2295_),
    .Q(\lfsr0.stop_reg[3] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net132),
    .D(_0217_),
    .Q_N(_2294_),
    .Q(\lfsr0.stop_reg[4] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net149),
    .D(_0218_),
    .Q_N(_2293_),
    .Q(\lfsr0.stop_reg[5] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net151),
    .D(_0219_),
    .Q_N(_2292_),
    .Q(\lfsr0.stop_reg[6] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net150),
    .D(_0220_),
    .Q_N(_2291_),
    .Q(\lfsr0.stop_reg[7] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net154),
    .D(_0221_),
    .Q_N(_2290_),
    .Q(\lfsr0.stop_reg[8] ));
 sg13g2_dfrbp_1 \lfsr0.stop_reg[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net151),
    .D(_0222_),
    .Q_N(_2484_),
    .Q(\lfsr0.stop_reg[9] ));
 sg13g2_dfrbp_1 \nreset_sync0.nreset_o$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1),
    .D(\nreset_sync0.r_sync ),
    .Q_N(_2485_),
    .Q(\gray_sobel0.gray_scale0.nreset_i ));
 sg13g2_dfrbp_1 \nreset_sync0.r_sync$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1),
    .D(net202),
    .Q_N(_2486_),
    .Q(\nreset_sync0.r_sync ));
 sg13g2_dfrbp_1 \sgnl_sync0.signal_o$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net160),
    .D(\sgnl_sync0.signal_sync ),
    .Q_N(_2487_),
    .Q(LFSR_enable_i_sync));
 sg13g2_dfrbp_1 \sgnl_sync0.signal_sync$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net160),
    .D(net7),
    .Q_N(_2488_),
    .Q(\sgnl_sync0.signal_sync ));
 sg13g2_dfrbp_1 \sgnl_sync1.signal_o$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net160),
    .D(\sgnl_sync1.signal_sync ),
    .Q_N(_2489_),
    .Q(\lfsr0.config_i ));
 sg13g2_dfrbp_1 \sgnl_sync1.signal_sync$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net160),
    .D(net8),
    .Q_N(_2490_),
    .Q(\sgnl_sync1.signal_sync ));
 sg13g2_dfrbp_1 \sgnl_sync2.signal_o$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net160),
    .D(\sgnl_sync2.signal_sync ),
    .Q_N(_2491_),
    .Q(\lfsr0.lfsr_en_i ));
 sg13g2_dfrbp_1 \sgnl_sync2.signal_sync$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net158),
    .D(net9),
    .Q_N(_2289_),
    .Q(\sgnl_sync2.signal_sync ));
 sg13g2_dfrbp_1 \spi0.data_rx[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net128),
    .D(_0223_),
    .Q_N(_2288_),
    .Q(\input_data[0] ));
 sg13g2_dfrbp_1 \spi0.data_rx[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net126),
    .D(_0224_),
    .Q_N(_2287_),
    .Q(\input_data[10] ));
 sg13g2_dfrbp_1 \spi0.data_rx[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net129),
    .D(_0225_),
    .Q_N(_2286_),
    .Q(\input_data[11] ));
 sg13g2_dfrbp_1 \spi0.data_rx[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net129),
    .D(_0226_),
    .Q_N(_2285_),
    .Q(\input_data[12] ));
 sg13g2_dfrbp_1 \spi0.data_rx[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net129),
    .D(_0227_),
    .Q_N(_2284_),
    .Q(\input_data[13] ));
 sg13g2_dfrbp_1 \spi0.data_rx[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0228_),
    .Q_N(_2283_),
    .Q(\input_data[14] ));
 sg13g2_dfrbp_1 \spi0.data_rx[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0229_),
    .Q_N(_2282_),
    .Q(\input_data[15] ));
 sg13g2_dfrbp_1 \spi0.data_rx[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net154),
    .D(_0230_),
    .Q_N(_2281_),
    .Q(\input_data[16] ));
 sg13g2_dfrbp_1 \spi0.data_rx[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net155),
    .D(_0231_),
    .Q_N(_2280_),
    .Q(\input_data[17] ));
 sg13g2_dfrbp_1 \spi0.data_rx[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net129),
    .D(_0232_),
    .Q_N(_2279_),
    .Q(\input_data[18] ));
 sg13g2_dfrbp_1 \spi0.data_rx[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net130),
    .D(_0233_),
    .Q_N(_2278_),
    .Q(\input_data[19] ));
 sg13g2_dfrbp_1 \spi0.data_rx[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net126),
    .D(_0234_),
    .Q_N(_2277_),
    .Q(\input_data[1] ));
 sg13g2_dfrbp_1 \spi0.data_rx[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net130),
    .D(_0235_),
    .Q_N(_2276_),
    .Q(\input_data[20] ));
 sg13g2_dfrbp_1 \spi0.data_rx[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net130),
    .D(_0236_),
    .Q_N(_2275_),
    .Q(\input_data[21] ));
 sg13g2_dfrbp_1 \spi0.data_rx[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net129),
    .D(_0237_),
    .Q_N(_2274_),
    .Q(\input_data[22] ));
 sg13g2_dfrbp_1 \spi0.data_rx[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net129),
    .D(_0238_),
    .Q_N(_2273_),
    .Q(\input_data[23] ));
 sg13g2_dfrbp_1 \spi0.data_rx[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net125),
    .D(_0239_),
    .Q_N(_2272_),
    .Q(\input_data[2] ));
 sg13g2_dfrbp_1 \spi0.data_rx[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net125),
    .D(_0240_),
    .Q_N(_2271_),
    .Q(\input_data[3] ));
 sg13g2_dfrbp_1 \spi0.data_rx[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net125),
    .D(_0241_),
    .Q_N(_2270_),
    .Q(\input_data[4] ));
 sg13g2_dfrbp_1 \spi0.data_rx[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net126),
    .D(_0242_),
    .Q_N(_2269_),
    .Q(\input_data[5] ));
 sg13g2_dfrbp_1 \spi0.data_rx[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net126),
    .D(_0243_),
    .Q_N(_2268_),
    .Q(\input_data[6] ));
 sg13g2_dfrbp_1 \spi0.data_rx[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net129),
    .D(_0244_),
    .Q_N(_2267_),
    .Q(\input_data[7] ));
 sg13g2_dfrbp_1 \spi0.data_rx[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net129),
    .D(_0245_),
    .Q_N(_2266_),
    .Q(\input_data[8] ));
 sg13g2_dfrbp_1 \spi0.data_rx[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net126),
    .D(_0246_),
    .Q_N(_2265_),
    .Q(\input_data[9] ));
 sg13g2_dfrbp_1 \spi0.data_tx[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net157),
    .D(_0247_),
    .Q_N(_2264_),
    .Q(\spi0.data_tx[0] ));
 sg13g2_dfrbp_1 \spi0.data_tx[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net161),
    .D(_0248_),
    .Q_N(_2263_),
    .Q(\spi0.data_tx[10] ));
 sg13g2_dfrbp_1 \spi0.data_tx[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net161),
    .D(_0249_),
    .Q_N(_2262_),
    .Q(\spi0.data_tx[11] ));
 sg13g2_dfrbp_1 \spi0.data_tx[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net161),
    .D(_0250_),
    .Q_N(_2261_),
    .Q(\spi0.data_tx[12] ));
 sg13g2_dfrbp_1 \spi0.data_tx[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net161),
    .D(_0251_),
    .Q_N(_2260_),
    .Q(\spi0.data_tx[13] ));
 sg13g2_dfrbp_1 \spi0.data_tx[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net161),
    .D(_0252_),
    .Q_N(_2259_),
    .Q(\spi0.data_tx[14] ));
 sg13g2_dfrbp_1 \spi0.data_tx[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net161),
    .D(_0253_),
    .Q_N(_2258_),
    .Q(\spi0.data_tx[15] ));
 sg13g2_dfrbp_1 \spi0.data_tx[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net155),
    .D(_0254_),
    .Q_N(_2257_),
    .Q(\spi0.data_tx[16] ));
 sg13g2_dfrbp_1 \spi0.data_tx[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net155),
    .D(_0255_),
    .Q_N(_2256_),
    .Q(\spi0.data_tx[17] ));
 sg13g2_dfrbp_1 \spi0.data_tx[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net155),
    .D(_0256_),
    .Q_N(_2255_),
    .Q(\spi0.data_tx[18] ));
 sg13g2_dfrbp_1 \spi0.data_tx[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net161),
    .D(_0257_),
    .Q_N(_2254_),
    .Q(\spi0.data_tx[19] ));
 sg13g2_dfrbp_1 \spi0.data_tx[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net157),
    .D(_0258_),
    .Q_N(_2253_),
    .Q(\spi0.data_tx[1] ));
 sg13g2_dfrbp_1 \spi0.data_tx[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net161),
    .D(_0259_),
    .Q_N(_2252_),
    .Q(\spi0.data_tx[20] ));
 sg13g2_dfrbp_1 \spi0.data_tx[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net162),
    .D(_0260_),
    .Q_N(_2251_),
    .Q(\spi0.data_tx[21] ));
 sg13g2_dfrbp_1 \spi0.data_tx[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net160),
    .D(_0261_),
    .Q_N(_2250_),
    .Q(\spi0.data_tx[22] ));
 sg13g2_dfrbp_1 \spi0.data_tx[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net160),
    .D(_0262_),
    .Q_N(_2249_),
    .Q(\spi0.data_tx[23] ));
 sg13g2_dfrbp_1 \spi0.data_tx[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net157),
    .D(_0263_),
    .Q_N(_2248_),
    .Q(\spi0.data_tx[2] ));
 sg13g2_dfrbp_1 \spi0.data_tx[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net158),
    .D(_0264_),
    .Q_N(_2247_),
    .Q(\spi0.data_tx[3] ));
 sg13g2_dfrbp_1 \spi0.data_tx[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net158),
    .D(_0265_),
    .Q_N(_2246_),
    .Q(\spi0.data_tx[4] ));
 sg13g2_dfrbp_1 \spi0.data_tx[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net158),
    .D(_0266_),
    .Q_N(_2245_),
    .Q(\spi0.data_tx[5] ));
 sg13g2_dfrbp_1 \spi0.data_tx[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net158),
    .D(_0267_),
    .Q_N(_2244_),
    .Q(\spi0.data_tx[6] ));
 sg13g2_dfrbp_1 \spi0.data_tx[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net159),
    .D(_0268_),
    .Q_N(_2243_),
    .Q(\spi0.data_tx[7] ));
 sg13g2_dfrbp_1 \spi0.data_tx[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net160),
    .D(_0269_),
    .Q_N(_2242_),
    .Q(\spi0.data_tx[8] ));
 sg13g2_dfrbp_1 \spi0.data_tx[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net159),
    .D(_0270_),
    .Q_N(_2492_),
    .Q(\spi0.data_tx[9] ));
 sg13g2_dfrbp_1 \spi0.px_rdy_i_spi_o$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net150),
    .D(\spi0.rxtx_done_rising ),
    .Q_N(_2493_),
    .Q(in_data_rdy));
 sg13g2_dfrbp_1 \spi0.rxtx_done_reg$_DFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net130),
    .D(\spi0.rxtx_done ),
    .Q_N(_2494_),
    .Q(\spi0.rxtx_done_reg ));
 sg13g2_dfrbp_1 \spi0.signal_sync1.signal_o$_DFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net130),
    .D(\spi0.signal_sync1.signal_sync ),
    .Q_N(_2495_),
    .Q(\spi0.rxtx_done ));
 sg13g2_dfrbp_1 \spi0.signal_sync1.signal_sync$_DFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net131),
    .D(\spi0.signal_sync1.async_signal_i ),
    .Q_N(_2241_),
    .Q(\spi0.signal_sync1.signal_sync ));
 sg13g2_dfrbp_1 \spi0.spi0.counter[0]$_DFF_NP0_  (.CLK(net178),
    .RESET_B(net172),
    .D(_0002_),
    .Q_N(_2240_),
    .Q(\spi0.spi0.counter[0] ));
 sg13g2_dfrbp_1 \spi0.spi0.counter[1]$_DFF_NP0_  (.CLK(net178),
    .RESET_B(net172),
    .D(_0003_),
    .Q_N(_2239_),
    .Q(\spi0.spi0.counter[1] ));
 sg13g2_dfrbp_1 \spi0.spi0.counter[2]$_DFF_NP0_  (.CLK(net178),
    .RESET_B(net172),
    .D(_0004_),
    .Q_N(_2238_),
    .Q(\spi0.spi0.counter[2] ));
 sg13g2_dfrbp_1 \spi0.spi0.counter[3]$_DFF_NP0_  (.CLK(net179),
    .RESET_B(net173),
    .D(_0005_),
    .Q_N(_2237_),
    .Q(\spi0.spi0.counter[3] ));
 sg13g2_dfrbp_1 \spi0.spi0.counter[4]$_DFF_NP0_  (.CLK(net178),
    .RESET_B(net172),
    .D(_0006_),
    .Q_N(_2236_),
    .Q(\spi0.spi0.counter[4] ));
 sg13g2_dfrbp_1 \spi0.spi0.counter[5]$_DFF_NP0_  (.CLK(net179),
    .RESET_B(net172),
    .D(_0007_),
    .Q_N(_2235_),
    .Q(\spi0.spi0.counter[5] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[0]$_DFF_PP0_  (.CLK(net185),
    .RESET_B(net172),
    .D(net4),
    .Q_N(_2234_),
    .Q(\spi0.spi0.data_rx_o[0] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[10]$_DFF_PP0_  (.CLK(net181),
    .RESET_B(net165),
    .D(\spi0.spi0.data_rx_o[9] ),
    .Q_N(_2233_),
    .Q(\spi0.spi0.data_rx_o[10] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[11]$_DFF_PP0_  (.CLK(net182),
    .RESET_B(net166),
    .D(\spi0.spi0.data_rx_o[10] ),
    .Q_N(_2232_),
    .Q(\spi0.spi0.data_rx_o[11] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[12]$_DFF_PP0_  (.CLK(net182),
    .RESET_B(net166),
    .D(\spi0.spi0.data_rx_o[11] ),
    .Q_N(_2231_),
    .Q(\spi0.spi0.data_rx_o[12] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[13]$_DFF_PP0_  (.CLK(net183),
    .RESET_B(net167),
    .D(\spi0.spi0.data_rx_o[12] ),
    .Q_N(_2230_),
    .Q(\spi0.spi0.data_rx_o[13] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[14]$_DFF_PP0_  (.CLK(net183),
    .RESET_B(net168),
    .D(\spi0.spi0.data_rx_o[13] ),
    .Q_N(_2229_),
    .Q(\spi0.spi0.data_rx_o[14] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[15]$_DFF_PP0_  (.CLK(net184),
    .RESET_B(net167),
    .D(\spi0.spi0.data_rx_o[14] ),
    .Q_N(_2228_),
    .Q(\spi0.spi0.data_rx_o[15] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[16]$_DFF_PP0_  (.CLK(net184),
    .RESET_B(net168),
    .D(\spi0.spi0.data_rx_o[15] ),
    .Q_N(_2227_),
    .Q(\spi0.spi0.data_rx_o[16] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[17]$_DFF_PP0_  (.CLK(net181),
    .RESET_B(net165),
    .D(\spi0.spi0.data_rx_o[16] ),
    .Q_N(_2226_),
    .Q(\spi0.spi0.data_rx_o[17] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[18]$_DFF_PP0_  (.CLK(net181),
    .RESET_B(net165),
    .D(\spi0.spi0.data_rx_o[17] ),
    .Q_N(_2225_),
    .Q(\spi0.spi0.data_rx_o[18] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[19]$_DFF_PP0_  (.CLK(net181),
    .RESET_B(net165),
    .D(\spi0.spi0.data_rx_o[18] ),
    .Q_N(_2224_),
    .Q(\spi0.spi0.data_rx_o[19] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[1]$_DFF_PP0_  (.CLK(net185),
    .RESET_B(net174),
    .D(\spi0.spi0.data_rx_o[0] ),
    .Q_N(_2223_),
    .Q(\spi0.spi0.data_rx_o[1] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[20]$_DFF_PP0_  (.CLK(net181),
    .RESET_B(net165),
    .D(\spi0.spi0.data_rx_o[19] ),
    .Q_N(_2222_),
    .Q(\spi0.spi0.data_rx_o[20] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[21]$_DFF_PP0_  (.CLK(net181),
    .RESET_B(net165),
    .D(\spi0.spi0.data_rx_o[20] ),
    .Q_N(_2221_),
    .Q(\spi0.spi0.data_rx_o[21] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[22]$_DFF_PP0_  (.CLK(net181),
    .RESET_B(net165),
    .D(\spi0.spi0.data_rx_o[21] ),
    .Q_N(_2220_),
    .Q(\spi0.spi0.data_rx_o[22] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[23]$_DFF_PP0_  (.CLK(net182),
    .RESET_B(net166),
    .D(\spi0.spi0.data_rx_o[22] ),
    .Q_N(_2219_),
    .Q(\spi0.spi0.data_rx_o[23] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[2]$_DFF_PP0_  (.CLK(net184),
    .RESET_B(net168),
    .D(\spi0.spi0.data_rx_o[1] ),
    .Q_N(_2218_),
    .Q(\spi0.spi0.data_rx_o[2] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[3]$_DFF_PP0_  (.CLK(net183),
    .RESET_B(net167),
    .D(\spi0.spi0.data_rx_o[2] ),
    .Q_N(_2217_),
    .Q(\spi0.spi0.data_rx_o[3] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[4]$_DFF_PP0_  (.CLK(net183),
    .RESET_B(net167),
    .D(\spi0.spi0.data_rx_o[3] ),
    .Q_N(_2216_),
    .Q(\spi0.spi0.data_rx_o[4] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[5]$_DFF_PP0_  (.CLK(net183),
    .RESET_B(net167),
    .D(\spi0.spi0.data_rx_o[4] ),
    .Q_N(_2215_),
    .Q(\spi0.spi0.data_rx_o[5] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[6]$_DFF_PP0_  (.CLK(net183),
    .RESET_B(net167),
    .D(\spi0.spi0.data_rx_o[5] ),
    .Q_N(_2214_),
    .Q(\spi0.spi0.data_rx_o[6] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[7]$_DFF_PP0_  (.CLK(net183),
    .RESET_B(net167),
    .D(\spi0.spi0.data_rx_o[6] ),
    .Q_N(_2213_),
    .Q(\spi0.spi0.data_rx_o[7] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[8]$_DFF_PP0_  (.CLK(net183),
    .RESET_B(net167),
    .D(\spi0.spi0.data_rx_o[7] ),
    .Q_N(_2212_),
    .Q(\spi0.spi0.data_rx_o[8] ));
 sg13g2_dfrbp_1 \spi0.spi0.data_rx_o[9]$_DFF_PP0_  (.CLK(net181),
    .RESET_B(net165),
    .D(\spi0.spi0.data_rx_o[8] ),
    .Q_N(_2211_),
    .Q(\spi0.spi0.data_rx_o[9] ));
 sg13g2_dfrbp_1 \spi0.spi0.rxtx_done_o$_DFF_PP0_  (.CLK(net185),
    .RESET_B(net174),
    .D(net61),
    .Q_N(_2210_),
    .Q(\spi0.signal_sync1.async_signal_i ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[0]$_DFF_NP0_  (.CLK(net177),
    .RESET_B(net171),
    .D(_0009_),
    .Q_N(_2209_),
    .Q(\spi0.spi0.sdo_register[0] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[10]$_DFF_NP0_  (.CLK(net176),
    .RESET_B(net170),
    .D(_0010_),
    .Q_N(_2208_),
    .Q(\spi0.spi0.sdo_register[10] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[11]$_DFF_NP0_  (.CLK(net177),
    .RESET_B(net171),
    .D(_0011_),
    .Q_N(_2207_),
    .Q(\spi0.spi0.sdo_register[11] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[12]$_DFF_NP0_  (.CLK(net177),
    .RESET_B(net171),
    .D(_0012_),
    .Q_N(_2206_),
    .Q(\spi0.spi0.sdo_register[12] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[13]$_DFF_NP0_  (.CLK(net177),
    .RESET_B(net171),
    .D(_0013_),
    .Q_N(_2205_),
    .Q(\spi0.spi0.sdo_register[13] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[14]$_DFF_NP0_  (.CLK(net177),
    .RESET_B(net173),
    .D(_0014_),
    .Q_N(_2204_),
    .Q(\spi0.spi0.sdo_register[14] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[15]$_DFF_NP0_  (.CLK(net176),
    .RESET_B(net170),
    .D(_0015_),
    .Q_N(_2203_),
    .Q(\spi0.spi0.sdo_register[15] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[16]$_DFF_NP0_  (.CLK(net176),
    .RESET_B(net170),
    .D(_0016_),
    .Q_N(_2202_),
    .Q(\spi0.spi0.sdo_register[16] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[17]$_DFF_NP0_  (.CLK(net175),
    .RESET_B(net169),
    .D(_0017_),
    .Q_N(_2201_),
    .Q(\spi0.spi0.sdo_register[17] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[18]$_DFF_NP0_  (.CLK(net175),
    .RESET_B(net169),
    .D(_0018_),
    .Q_N(_2200_),
    .Q(\spi0.spi0.sdo_register[18] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[19]$_DFF_NP0_  (.CLK(net175),
    .RESET_B(net169),
    .D(_0019_),
    .Q_N(_2199_),
    .Q(\spi0.spi0.sdo_register[19] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[1]$_DFF_NP0_  (.CLK(net177),
    .RESET_B(net171),
    .D(_0020_),
    .Q_N(_2198_),
    .Q(\spi0.spi0.sdo_register[1] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[20]$_DFF_NP0_  (.CLK(net175),
    .RESET_B(net169),
    .D(_0021_),
    .Q_N(_2197_),
    .Q(\spi0.spi0.sdo_register[20] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[21]$_DFF_NP0_  (.CLK(net175),
    .RESET_B(net169),
    .D(_0022_),
    .Q_N(_2196_),
    .Q(\spi0.spi0.sdo_register[21] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[22]$_DFF_NP0_  (.CLK(net175),
    .RESET_B(net169),
    .D(_0023_),
    .Q_N(_2195_),
    .Q(\spi0.spi0.sdo_register[22] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[23]$_DFF_NP0_  (.CLK(net175),
    .RESET_B(net169),
    .D(_0024_),
    .Q_N(_2194_),
    .Q(\spi0.spi0.sdo_o ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[2]$_DFF_NP0_  (.CLK(net177),
    .RESET_B(net171),
    .D(_0025_),
    .Q_N(_2193_),
    .Q(\spi0.spi0.sdo_register[2] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[3]$_DFF_NP0_  (.CLK(net177),
    .RESET_B(net171),
    .D(_0026_),
    .Q_N(_2192_),
    .Q(\spi0.spi0.sdo_register[3] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[4]$_DFF_NP0_  (.CLK(net178),
    .RESET_B(net171),
    .D(_0027_),
    .Q_N(_2191_),
    .Q(\spi0.spi0.sdo_register[4] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[5]$_DFF_NP0_  (.CLK(net178),
    .RESET_B(net172),
    .D(_0028_),
    .Q_N(_2190_),
    .Q(\spi0.spi0.sdo_register[5] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[6]$_DFF_NP0_  (.CLK(net178),
    .RESET_B(net172),
    .D(_0029_),
    .Q_N(_2189_),
    .Q(\spi0.spi0.sdo_register[6] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[7]$_DFF_NP0_  (.CLK(net176),
    .RESET_B(net170),
    .D(_0030_),
    .Q_N(_2188_),
    .Q(\spi0.spi0.sdo_register[7] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[8]$_DFF_NP0_  (.CLK(net175),
    .RESET_B(net169),
    .D(_0031_),
    .Q_N(_2187_),
    .Q(\spi0.spi0.sdo_register[8] ));
 sg13g2_dfrbp_1 \spi0.spi0.sdo_register[9]$_DFF_NP0_  (.CLK(net176),
    .RESET_B(net170),
    .D(_0032_),
    .Q_N(_2186_),
    .Q(\spi0.spi0.sdo_register[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[0]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[1]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[2]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[3]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[6]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout18 (.A(_1215_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0813_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_1201_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_2157_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0001_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_2177_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1957_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1594_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1555_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1536_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1500_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_2179_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_2154_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1578_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0296_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_2155_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1614_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0801_),
    .X(net35));
 sg13g2_buf_4 fanout36 (.X(net36),
    .A(_1827_));
 sg13g2_buf_4 fanout37 (.X(net37),
    .A(_1826_));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(_1823_));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(_1822_));
 sg13g2_buf_2 fanout40 (.A(_1753_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1733_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1725_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1724_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1729_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1543_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1521_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1502_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1501_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0916_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0644_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(\gray_sobel0.sobel0.next[1] ),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1731_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1708_),
    .X(net53));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(_1454_));
 sg13g2_buf_2 fanout55 (.A(_1973_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1676_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1657_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1642_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1972_),
    .X(net59));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(_1928_));
 sg13g2_buf_2 fanout61 (.A(_0008_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(\gray_sobel0.sobel0.next[0] ),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1874_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1870_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0394_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_2044_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1917_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0702_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1916_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1989_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1915_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_1707_));
 sg13g2_buf_4 fanout73 (.X(net73),
    .A(\spi0.rxtx_done_rising ));
 sg13g2_buf_2 fanout74 (.A(_0763_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0490_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0483_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0460_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1914_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1873_),
    .X(net79));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_1738_));
 sg13g2_buf_2 fanout81 (.A(_1711_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1710_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1658_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1644_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1627_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0776_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0751_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0608_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0577_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0506_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0482_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0345_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1913_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_1872_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_1715_),
    .X(net95));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(_1443_));
 sg13g2_buf_2 fanout97 (.A(_0755_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0750_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0606_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0458_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0404_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0390_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0385_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0384_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0382_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0369_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0368_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0363_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0361_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_0360_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0342_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_2013_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_1997_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_1976_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_1967_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_1853_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_1850_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_1842_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_1839_),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(net121));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(net124));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(net123));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(net124));
 sg13g2_buf_2 fanout124 (.A(\gray_sobel0.gray_scale0.nreset_i ),
    .X(net124));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(net128));
 sg13g2_buf_2 fanout126 (.A(net128),
    .X(net126));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(net128));
 sg13g2_buf_2 fanout128 (.A(net138),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(net131));
 sg13g2_buf_2 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(net138),
    .X(net131));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(net134));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net138));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net137));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(net137));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net138));
 sg13g2_buf_1 fanout138 (.A(\gray_sobel0.gray_scale0.nreset_i ),
    .X(net138));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net143));
 sg13g2_buf_2 fanout140 (.A(net143),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net143));
 sg13g2_buf_2 fanout142 (.A(net143),
    .X(net142));
 sg13g2_buf_1 fanout143 (.A(net147),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net146));
 sg13g2_buf_2 fanout145 (.A(net146),
    .X(net145));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net147));
 sg13g2_buf_1 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net163));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(net151));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(net151));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(net163));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(net156));
 sg13g2_buf_2 fanout153 (.A(net156),
    .X(net153));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(net156));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(net156));
 sg13g2_buf_1 fanout156 (.A(net163),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(net159));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net159));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(net162));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(net162));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(net162));
 sg13g2_buf_1 fanout162 (.A(net163),
    .X(net162));
 sg13g2_buf_1 fanout163 (.A(\gray_sobel0.gray_scale0.nreset_i ),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_1714_),
    .X(net164));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(net166));
 sg13g2_buf_2 fanout166 (.A(net168),
    .X(net166));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(net168));
 sg13g2_buf_2 fanout168 (.A(_0041_),
    .X(net168));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(net170));
 sg13g2_buf_2 fanout170 (.A(net174),
    .X(net170));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(net173));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(net173));
 sg13g2_buf_2 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_1 fanout174 (.A(_0041_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_1 fanout176 (.A(net179),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_1 fanout179 (.A(_0042_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_1945_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(net182),
    .X(net181));
 sg13g2_buf_1 fanout182 (.A(net184),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_1 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_1 fanout185 (.A(net2),
    .X(net185));
 sg13g2_tielo _4697__186 (.L_LO(net186));
 sg13g2_tielo _4698__187 (.L_LO(net187));
 sg13g2_tielo _4699__188 (.L_LO(net188));
 sg13g2_tielo _4700__189 (.L_LO(net189));
 sg13g2_tielo _4701__190 (.L_LO(net190));
 sg13g2_tielo _4702__191 (.L_LO(net191));
 sg13g2_tielo _4703__192 (.L_LO(net192));
 sg13g2_tielo _4704__193 (.L_LO(net193));
 sg13g2_tielo _4705__194 (.L_LO(net194));
 sg13g2_tielo _4706__195 (.L_LO(net195));
 sg13g2_tielo _4707__196 (.L_LO(net196));
 sg13g2_tielo _4708__197 (.L_LO(net197));
 sg13g2_tielo _4709__198 (.L_LO(net198));
 sg13g2_tielo _4710__199 (.L_LO(net199));
 sg13g2_tielo _4711__200 (.L_LO(net200));
 sg13g2_tielo _4712__201 (.L_LO(net201));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_33_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_34_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_35_clk));
 sg13g2_buf_16 clkload5 (.A(clknet_leaf_36_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_leaf_0_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_32_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_37_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_27_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_29_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_leaf_22_clk));
 sg13g2_buf_16 clkload12 (.A(clknet_leaf_1_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_9_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_7_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_leaf_19_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_13_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_15_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(\spi0.signal_sync1.async_signal_i ));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(\spi0.signal_sync1.async_signal_i ));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_antennanp ANTENNA_7 (.A(\spi0.signal_sync1.async_signal_i ));
 sg13g2_antennanp ANTENNA_8 (.A(\spi0.signal_sync1.async_signal_i ));
 sg13g2_antennanp ANTENNA_9 (.A(\spi0.signal_sync1.async_signal_i ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_fill_2 FILLER_0_343 ();
 sg13g2_fill_1 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_4 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_2 FILLER_1_49 ();
 sg13g2_decap_4 FILLER_1_90 ();
 sg13g2_decap_8 FILLER_1_120 ();
 sg13g2_fill_2 FILLER_1_127 ();
 sg13g2_decap_8 FILLER_1_155 ();
 sg13g2_fill_2 FILLER_1_162 ();
 sg13g2_decap_4 FILLER_1_200 ();
 sg13g2_fill_1 FILLER_1_204 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_283 ();
 sg13g2_decap_8 FILLER_1_290 ();
 sg13g2_decap_8 FILLER_1_297 ();
 sg13g2_decap_4 FILLER_1_304 ();
 sg13g2_fill_2 FILLER_1_308 ();
 sg13g2_decap_4 FILLER_1_346 ();
 sg13g2_fill_1 FILLER_1_350 ();
 sg13g2_decap_4 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_4 FILLER_2_28 ();
 sg13g2_fill_1 FILLER_2_32 ();
 sg13g2_decap_4 FILLER_2_59 ();
 sg13g2_fill_1 FILLER_2_63 ();
 sg13g2_fill_1 FILLER_2_84 ();
 sg13g2_fill_1 FILLER_2_98 ();
 sg13g2_fill_1 FILLER_2_107 ();
 sg13g2_fill_1 FILLER_2_138 ();
 sg13g2_fill_1 FILLER_2_142 ();
 sg13g2_fill_2 FILLER_2_148 ();
 sg13g2_fill_2 FILLER_2_154 ();
 sg13g2_fill_2 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_163 ();
 sg13g2_decap_8 FILLER_2_190 ();
 sg13g2_decap_8 FILLER_2_201 ();
 sg13g2_decap_8 FILLER_2_208 ();
 sg13g2_decap_8 FILLER_2_215 ();
 sg13g2_decap_8 FILLER_2_222 ();
 sg13g2_decap_8 FILLER_2_229 ();
 sg13g2_decap_8 FILLER_2_236 ();
 sg13g2_fill_2 FILLER_2_243 ();
 sg13g2_fill_1 FILLER_2_245 ();
 sg13g2_fill_2 FILLER_2_334 ();
 sg13g2_fill_1 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_decap_8 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_2_414 ();
 sg13g2_decap_8 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_428 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_55 ();
 sg13g2_fill_1 FILLER_3_57 ();
 sg13g2_fill_2 FILLER_3_98 ();
 sg13g2_fill_1 FILLER_3_105 ();
 sg13g2_fill_2 FILLER_3_111 ();
 sg13g2_fill_1 FILLER_3_113 ();
 sg13g2_decap_8 FILLER_3_122 ();
 sg13g2_decap_4 FILLER_3_129 ();
 sg13g2_fill_2 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_171 ();
 sg13g2_fill_2 FILLER_3_182 ();
 sg13g2_fill_2 FILLER_3_192 ();
 sg13g2_fill_1 FILLER_3_194 ();
 sg13g2_fill_1 FILLER_3_225 ();
 sg13g2_decap_8 FILLER_3_230 ();
 sg13g2_decap_4 FILLER_3_237 ();
 sg13g2_fill_2 FILLER_3_241 ();
 sg13g2_decap_8 FILLER_3_269 ();
 sg13g2_fill_1 FILLER_3_276 ();
 sg13g2_decap_4 FILLER_3_313 ();
 sg13g2_fill_2 FILLER_3_317 ();
 sg13g2_decap_4 FILLER_3_324 ();
 sg13g2_fill_1 FILLER_3_328 ();
 sg13g2_fill_2 FILLER_3_339 ();
 sg13g2_fill_1 FILLER_3_341 ();
 sg13g2_fill_1 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_414 ();
 sg13g2_decap_8 FILLER_3_421 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_fill_2 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_66 ();
 sg13g2_decap_8 FILLER_4_73 ();
 sg13g2_decap_8 FILLER_4_80 ();
 sg13g2_decap_8 FILLER_4_87 ();
 sg13g2_decap_8 FILLER_4_94 ();
 sg13g2_decap_4 FILLER_4_101 ();
 sg13g2_fill_1 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_132 ();
 sg13g2_decap_8 FILLER_4_139 ();
 sg13g2_fill_2 FILLER_4_146 ();
 sg13g2_fill_1 FILLER_4_148 ();
 sg13g2_fill_1 FILLER_4_162 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_203 ();
 sg13g2_fill_2 FILLER_4_218 ();
 sg13g2_fill_1 FILLER_4_220 ();
 sg13g2_decap_8 FILLER_4_226 ();
 sg13g2_decap_4 FILLER_4_233 ();
 sg13g2_fill_1 FILLER_4_237 ();
 sg13g2_decap_8 FILLER_4_248 ();
 sg13g2_decap_8 FILLER_4_255 ();
 sg13g2_fill_2 FILLER_4_262 ();
 sg13g2_decap_4 FILLER_4_269 ();
 sg13g2_fill_1 FILLER_4_273 ();
 sg13g2_decap_4 FILLER_4_288 ();
 sg13g2_fill_1 FILLER_4_292 ();
 sg13g2_fill_1 FILLER_4_302 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_decap_8 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_4_415 ();
 sg13g2_decap_8 FILLER_4_422 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_fill_2 FILLER_5_98 ();
 sg13g2_fill_1 FILLER_5_100 ();
 sg13g2_fill_2 FILLER_5_105 ();
 sg13g2_fill_1 FILLER_5_107 ();
 sg13g2_decap_4 FILLER_5_118 ();
 sg13g2_fill_1 FILLER_5_122 ();
 sg13g2_decap_4 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_fill_2 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_218 ();
 sg13g2_decap_8 FILLER_5_225 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_fill_2 FILLER_5_239 ();
 sg13g2_decap_4 FILLER_5_267 ();
 sg13g2_fill_2 FILLER_5_271 ();
 sg13g2_decap_4 FILLER_5_335 ();
 sg13g2_fill_2 FILLER_5_339 ();
 sg13g2_fill_2 FILLER_5_352 ();
 sg13g2_fill_1 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_2 FILLER_6_18 ();
 sg13g2_fill_1 FILLER_6_46 ();
 sg13g2_fill_1 FILLER_6_52 ();
 sg13g2_fill_1 FILLER_6_58 ();
 sg13g2_fill_2 FILLER_6_63 ();
 sg13g2_fill_1 FILLER_6_65 ();
 sg13g2_decap_4 FILLER_6_76 ();
 sg13g2_fill_1 FILLER_6_80 ();
 sg13g2_decap_4 FILLER_6_109 ();
 sg13g2_fill_1 FILLER_6_113 ();
 sg13g2_decap_8 FILLER_6_118 ();
 sg13g2_decap_8 FILLER_6_125 ();
 sg13g2_decap_8 FILLER_6_132 ();
 sg13g2_decap_4 FILLER_6_139 ();
 sg13g2_fill_1 FILLER_6_143 ();
 sg13g2_decap_4 FILLER_6_148 ();
 sg13g2_fill_2 FILLER_6_161 ();
 sg13g2_fill_1 FILLER_6_176 ();
 sg13g2_fill_2 FILLER_6_185 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_279 ();
 sg13g2_decap_8 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_293 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_fill_1 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_419 ();
 sg13g2_decap_4 FILLER_6_426 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_4 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_18 ();
 sg13g2_fill_1 FILLER_7_45 ();
 sg13g2_fill_1 FILLER_7_54 ();
 sg13g2_decap_4 FILLER_7_60 ();
 sg13g2_fill_1 FILLER_7_64 ();
 sg13g2_decap_4 FILLER_7_73 ();
 sg13g2_fill_2 FILLER_7_77 ();
 sg13g2_fill_2 FILLER_7_110 ();
 sg13g2_decap_4 FILLER_7_138 ();
 sg13g2_decap_8 FILLER_7_145 ();
 sg13g2_decap_8 FILLER_7_152 ();
 sg13g2_fill_2 FILLER_7_159 ();
 sg13g2_fill_1 FILLER_7_161 ();
 sg13g2_decap_4 FILLER_7_178 ();
 sg13g2_decap_8 FILLER_7_207 ();
 sg13g2_decap_4 FILLER_7_214 ();
 sg13g2_fill_2 FILLER_7_218 ();
 sg13g2_decap_4 FILLER_7_250 ();
 sg13g2_fill_2 FILLER_7_254 ();
 sg13g2_decap_8 FILLER_7_317 ();
 sg13g2_decap_8 FILLER_7_324 ();
 sg13g2_fill_1 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_8 FILLER_7_344 ();
 sg13g2_decap_4 FILLER_7_351 ();
 sg13g2_fill_1 FILLER_7_355 ();
 sg13g2_decap_4 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_decap_8 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_7_414 ();
 sg13g2_decap_8 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_fill_2 FILLER_8_35 ();
 sg13g2_fill_2 FILLER_8_83 ();
 sg13g2_decap_4 FILLER_8_93 ();
 sg13g2_fill_2 FILLER_8_108 ();
 sg13g2_fill_1 FILLER_8_110 ();
 sg13g2_fill_2 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_4 FILLER_8_161 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_fill_1 FILLER_8_178 ();
 sg13g2_fill_2 FILLER_8_184 ();
 sg13g2_fill_1 FILLER_8_204 ();
 sg13g2_decap_8 FILLER_8_220 ();
 sg13g2_decap_8 FILLER_8_227 ();
 sg13g2_decap_8 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_241 ();
 sg13g2_decap_4 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_264 ();
 sg13g2_decap_8 FILLER_8_271 ();
 sg13g2_fill_2 FILLER_8_278 ();
 sg13g2_fill_2 FILLER_8_332 ();
 sg13g2_fill_1 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_8 FILLER_8_404 ();
 sg13g2_decap_8 FILLER_8_411 ();
 sg13g2_decap_8 FILLER_8_418 ();
 sg13g2_decap_4 FILLER_8_425 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_fill_2 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_37 ();
 sg13g2_decap_4 FILLER_9_44 ();
 sg13g2_fill_2 FILLER_9_48 ();
 sg13g2_decap_8 FILLER_9_64 ();
 sg13g2_decap_8 FILLER_9_71 ();
 sg13g2_decap_4 FILLER_9_82 ();
 sg13g2_fill_2 FILLER_9_86 ();
 sg13g2_fill_1 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_4 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_170 ();
 sg13g2_decap_4 FILLER_9_177 ();
 sg13g2_fill_1 FILLER_9_181 ();
 sg13g2_decap_4 FILLER_9_186 ();
 sg13g2_fill_2 FILLER_9_190 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_213 ();
 sg13g2_fill_2 FILLER_9_220 ();
 sg13g2_decap_4 FILLER_9_227 ();
 sg13g2_fill_2 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_289 ();
 sg13g2_fill_2 FILLER_9_299 ();
 sg13g2_fill_1 FILLER_9_306 ();
 sg13g2_fill_2 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_4 FILLER_9_383 ();
 sg13g2_fill_1 FILLER_9_387 ();
 sg13g2_fill_2 FILLER_9_391 ();
 sg13g2_fill_1 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_31 ();
 sg13g2_fill_2 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_72 ();
 sg13g2_decap_8 FILLER_10_79 ();
 sg13g2_decap_8 FILLER_10_86 ();
 sg13g2_decap_8 FILLER_10_97 ();
 sg13g2_fill_2 FILLER_10_104 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_decap_4 FILLER_10_136 ();
 sg13g2_fill_2 FILLER_10_140 ();
 sg13g2_fill_2 FILLER_10_173 ();
 sg13g2_fill_2 FILLER_10_179 ();
 sg13g2_fill_1 FILLER_10_181 ();
 sg13g2_fill_1 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_fill_2 FILLER_10_238 ();
 sg13g2_decap_4 FILLER_10_244 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_decap_4 FILLER_10_275 ();
 sg13g2_fill_1 FILLER_10_279 ();
 sg13g2_fill_1 FILLER_10_285 ();
 sg13g2_fill_2 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_fill_2 FILLER_10_338 ();
 sg13g2_decap_4 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_32 ();
 sg13g2_fill_2 FILLER_11_59 ();
 sg13g2_fill_1 FILLER_11_61 ();
 sg13g2_decap_4 FILLER_11_82 ();
 sg13g2_decap_8 FILLER_11_90 ();
 sg13g2_decap_8 FILLER_11_97 ();
 sg13g2_decap_8 FILLER_11_104 ();
 sg13g2_fill_1 FILLER_11_111 ();
 sg13g2_decap_8 FILLER_11_117 ();
 sg13g2_decap_4 FILLER_11_124 ();
 sg13g2_fill_2 FILLER_11_128 ();
 sg13g2_decap_8 FILLER_11_146 ();
 sg13g2_decap_8 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_fill_2 FILLER_11_183 ();
 sg13g2_decap_4 FILLER_11_210 ();
 sg13g2_fill_2 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_229 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_fill_2 FILLER_11_264 ();
 sg13g2_fill_1 FILLER_11_266 ();
 sg13g2_decap_4 FILLER_11_293 ();
 sg13g2_fill_1 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_decap_4 FILLER_11_335 ();
 sg13g2_fill_2 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_fill_1 FILLER_11_353 ();
 sg13g2_fill_2 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_416 ();
 sg13g2_decap_8 FILLER_11_423 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_decap_4 FILLER_12_23 ();
 sg13g2_decap_4 FILLER_12_31 ();
 sg13g2_fill_2 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_45 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_fill_1 FILLER_12_86 ();
 sg13g2_decap_4 FILLER_12_92 ();
 sg13g2_decap_4 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_4 FILLER_12_158 ();
 sg13g2_fill_2 FILLER_12_162 ();
 sg13g2_fill_1 FILLER_12_174 ();
 sg13g2_fill_1 FILLER_12_181 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_fill_2 FILLER_12_201 ();
 sg13g2_fill_1 FILLER_12_203 ();
 sg13g2_decap_4 FILLER_12_209 ();
 sg13g2_decap_4 FILLER_12_218 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_decap_8 FILLER_12_241 ();
 sg13g2_decap_8 FILLER_12_248 ();
 sg13g2_decap_8 FILLER_12_255 ();
 sg13g2_decap_8 FILLER_12_262 ();
 sg13g2_decap_8 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_283 ();
 sg13g2_decap_8 FILLER_12_290 ();
 sg13g2_decap_8 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_304 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_4 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_12_411 ();
 sg13g2_decap_8 FILLER_12_417 ();
 sg13g2_decap_4 FILLER_12_424 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_22 ();
 sg13g2_fill_1 FILLER_13_29 ();
 sg13g2_decap_8 FILLER_13_45 ();
 sg13g2_fill_2 FILLER_13_52 ();
 sg13g2_fill_1 FILLER_13_54 ();
 sg13g2_fill_2 FILLER_13_67 ();
 sg13g2_fill_1 FILLER_13_69 ();
 sg13g2_decap_4 FILLER_13_75 ();
 sg13g2_fill_2 FILLER_13_79 ();
 sg13g2_decap_8 FILLER_13_132 ();
 sg13g2_decap_4 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_169 ();
 sg13g2_decap_4 FILLER_13_176 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_205 ();
 sg13g2_decap_8 FILLER_13_248 ();
 sg13g2_decap_8 FILLER_13_255 ();
 sg13g2_decap_8 FILLER_13_262 ();
 sg13g2_decap_4 FILLER_13_269 ();
 sg13g2_decap_4 FILLER_13_309 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_fill_2 FILLER_13_341 ();
 sg13g2_fill_1 FILLER_13_343 ();
 sg13g2_decap_4 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_fill_2 FILLER_13_391 ();
 sg13g2_fill_1 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_31 ();
 sg13g2_decap_8 FILLER_14_38 ();
 sg13g2_decap_8 FILLER_14_45 ();
 sg13g2_fill_2 FILLER_14_52 ();
 sg13g2_decap_8 FILLER_14_71 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_100 ();
 sg13g2_decap_4 FILLER_14_113 ();
 sg13g2_fill_2 FILLER_14_121 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_fill_2 FILLER_14_140 ();
 sg13g2_fill_1 FILLER_14_142 ();
 sg13g2_fill_2 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_157 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_4 FILLER_14_186 ();
 sg13g2_fill_2 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_202 ();
 sg13g2_decap_8 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_223 ();
 sg13g2_decap_8 FILLER_14_230 ();
 sg13g2_fill_2 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_fill_2 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_fill_2 FILLER_14_324 ();
 sg13g2_fill_1 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_decap_4 FILLER_14_338 ();
 sg13g2_fill_1 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_4 FILLER_14_391 ();
 sg13g2_fill_1 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_13 ();
 sg13g2_fill_2 FILLER_15_24 ();
 sg13g2_fill_1 FILLER_15_26 ();
 sg13g2_fill_2 FILLER_15_31 ();
 sg13g2_fill_1 FILLER_15_33 ();
 sg13g2_fill_2 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_55 ();
 sg13g2_decap_8 FILLER_15_62 ();
 sg13g2_fill_1 FILLER_15_69 ();
 sg13g2_decap_8 FILLER_15_83 ();
 sg13g2_decap_8 FILLER_15_90 ();
 sg13g2_decap_8 FILLER_15_97 ();
 sg13g2_decap_8 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_111 ();
 sg13g2_decap_8 FILLER_15_118 ();
 sg13g2_decap_8 FILLER_15_125 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_fill_1 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_decap_8 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_4 FILLER_15_196 ();
 sg13g2_fill_1 FILLER_15_200 ();
 sg13g2_decap_4 FILLER_15_208 ();
 sg13g2_fill_1 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_242 ();
 sg13g2_fill_1 FILLER_15_249 ();
 sg13g2_decap_8 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_283 ();
 sg13g2_fill_2 FILLER_15_307 ();
 sg13g2_fill_2 FILLER_15_337 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_fill_2 FILLER_15_359 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_decap_4 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_16 ();
 sg13g2_fill_2 FILLER_16_31 ();
 sg13g2_fill_2 FILLER_16_37 ();
 sg13g2_fill_1 FILLER_16_44 ();
 sg13g2_fill_2 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_55 ();
 sg13g2_fill_2 FILLER_16_62 ();
 sg13g2_fill_2 FILLER_16_69 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_decap_4 FILLER_16_88 ();
 sg13g2_fill_1 FILLER_16_92 ();
 sg13g2_decap_4 FILLER_16_110 ();
 sg13g2_decap_8 FILLER_16_122 ();
 sg13g2_fill_1 FILLER_16_129 ();
 sg13g2_decap_8 FILLER_16_152 ();
 sg13g2_decap_4 FILLER_16_159 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_4 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_179 ();
 sg13g2_fill_1 FILLER_16_184 ();
 sg13g2_decap_4 FILLER_16_189 ();
 sg13g2_decap_4 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_fill_1 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_279 ();
 sg13g2_fill_2 FILLER_16_289 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_2 FILLER_17_10 ();
 sg13g2_fill_1 FILLER_17_12 ();
 sg13g2_fill_1 FILLER_17_34 ();
 sg13g2_fill_1 FILLER_17_45 ();
 sg13g2_fill_1 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_61 ();
 sg13g2_decap_4 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_113 ();
 sg13g2_fill_1 FILLER_17_115 ();
 sg13g2_decap_8 FILLER_17_121 ();
 sg13g2_fill_2 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_150 ();
 sg13g2_decap_4 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_fill_2 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_246 ();
 sg13g2_fill_2 FILLER_17_291 ();
 sg13g2_fill_1 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_fill_2 FILLER_17_328 ();
 sg13g2_decap_4 FILLER_17_344 ();
 sg13g2_fill_2 FILLER_17_356 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_17_385 ();
 sg13g2_decap_4 FILLER_17_395 ();
 sg13g2_fill_2 FILLER_17_404 ();
 sg13g2_decap_8 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_4 FILLER_17_424 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_fill_1 FILLER_18_29 ();
 sg13g2_fill_1 FILLER_18_58 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_84 ();
 sg13g2_fill_1 FILLER_18_86 ();
 sg13g2_fill_2 FILLER_18_99 ();
 sg13g2_fill_1 FILLER_18_101 ();
 sg13g2_decap_4 FILLER_18_106 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_2 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_141 ();
 sg13g2_decap_4 FILLER_18_163 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_fill_1 FILLER_18_186 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_fill_2 FILLER_18_215 ();
 sg13g2_fill_1 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_4 FILLER_18_244 ();
 sg13g2_fill_1 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_decap_8 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_325 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_2 FILLER_18_338 ();
 sg13g2_fill_2 FILLER_18_348 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_4 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_414 ();
 sg13g2_decap_8 FILLER_18_421 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_decap_8 FILLER_19_27 ();
 sg13g2_decap_8 FILLER_19_34 ();
 sg13g2_fill_1 FILLER_19_41 ();
 sg13g2_decap_8 FILLER_19_50 ();
 sg13g2_decap_8 FILLER_19_57 ();
 sg13g2_decap_8 FILLER_19_64 ();
 sg13g2_decap_4 FILLER_19_71 ();
 sg13g2_fill_2 FILLER_19_75 ();
 sg13g2_decap_8 FILLER_19_82 ();
 sg13g2_decap_4 FILLER_19_89 ();
 sg13g2_fill_2 FILLER_19_93 ();
 sg13g2_fill_2 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_100 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_107 ();
 sg13g2_fill_2 FILLER_19_113 ();
 sg13g2_decap_8 FILLER_19_131 ();
 sg13g2_decap_4 FILLER_19_138 ();
 sg13g2_fill_2 FILLER_19_142 ();
 sg13g2_fill_2 FILLER_19_149 ();
 sg13g2_fill_2 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_158 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_fill_1 FILLER_19_192 ();
 sg13g2_fill_1 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_215 ();
 sg13g2_decap_8 FILLER_19_222 ();
 sg13g2_decap_8 FILLER_19_229 ();
 sg13g2_decap_8 FILLER_19_236 ();
 sg13g2_fill_2 FILLER_19_243 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_344 ();
 sg13g2_decap_4 FILLER_19_379 ();
 sg13g2_fill_2 FILLER_19_383 ();
 sg13g2_fill_2 FILLER_19_389 ();
 sg13g2_fill_1 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_19_409 ();
 sg13g2_decap_8 FILLER_19_416 ();
 sg13g2_decap_8 FILLER_19_423 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_27 ();
 sg13g2_decap_8 FILLER_20_34 ();
 sg13g2_decap_8 FILLER_20_41 ();
 sg13g2_fill_2 FILLER_20_48 ();
 sg13g2_decap_4 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_120 ();
 sg13g2_decap_8 FILLER_20_127 ();
 sg13g2_decap_8 FILLER_20_134 ();
 sg13g2_fill_2 FILLER_20_141 ();
 sg13g2_fill_1 FILLER_20_143 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_decap_4 FILLER_20_169 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_decap_8 FILLER_20_218 ();
 sg13g2_decap_8 FILLER_20_225 ();
 sg13g2_decap_8 FILLER_20_232 ();
 sg13g2_fill_2 FILLER_20_239 ();
 sg13g2_fill_1 FILLER_20_241 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_fill_2 FILLER_20_283 ();
 sg13g2_fill_1 FILLER_20_285 ();
 sg13g2_decap_8 FILLER_20_295 ();
 sg13g2_fill_1 FILLER_20_302 ();
 sg13g2_decap_4 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_4 FILLER_20_342 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_fill_2 FILLER_20_371 ();
 sg13g2_fill_1 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_20_409 ();
 sg13g2_decap_8 FILLER_20_416 ();
 sg13g2_decap_8 FILLER_20_423 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_9 ();
 sg13g2_decap_4 FILLER_21_23 ();
 sg13g2_fill_2 FILLER_21_27 ();
 sg13g2_decap_8 FILLER_21_33 ();
 sg13g2_decap_8 FILLER_21_40 ();
 sg13g2_decap_4 FILLER_21_47 ();
 sg13g2_fill_2 FILLER_21_51 ();
 sg13g2_fill_2 FILLER_21_57 ();
 sg13g2_fill_1 FILLER_21_59 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_decap_4 FILLER_21_72 ();
 sg13g2_fill_1 FILLER_21_76 ();
 sg13g2_decap_8 FILLER_21_108 ();
 sg13g2_decap_8 FILLER_21_115 ();
 sg13g2_decap_8 FILLER_21_122 ();
 sg13g2_decap_4 FILLER_21_129 ();
 sg13g2_decap_4 FILLER_21_137 ();
 sg13g2_fill_2 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_decap_8 FILLER_21_192 ();
 sg13g2_decap_8 FILLER_21_199 ();
 sg13g2_decap_4 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_248 ();
 sg13g2_decap_8 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_decap_4 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_decap_4 FILLER_21_302 ();
 sg13g2_fill_1 FILLER_21_306 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_337 ();
 sg13g2_decap_4 FILLER_21_346 ();
 sg13g2_fill_1 FILLER_21_350 ();
 sg13g2_fill_1 FILLER_21_368 ();
 sg13g2_fill_2 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_414 ();
 sg13g2_decap_8 FILLER_21_421 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_43 ();
 sg13g2_decap_8 FILLER_22_50 ();
 sg13g2_decap_8 FILLER_22_57 ();
 sg13g2_fill_2 FILLER_22_64 ();
 sg13g2_fill_1 FILLER_22_66 ();
 sg13g2_decap_8 FILLER_22_72 ();
 sg13g2_decap_8 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_86 ();
 sg13g2_fill_2 FILLER_22_92 ();
 sg13g2_fill_1 FILLER_22_94 ();
 sg13g2_decap_4 FILLER_22_121 ();
 sg13g2_fill_2 FILLER_22_130 ();
 sg13g2_fill_2 FILLER_22_163 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_decap_4 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_240 ();
 sg13g2_decap_8 FILLER_22_247 ();
 sg13g2_decap_4 FILLER_22_262 ();
 sg13g2_decap_4 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_282 ();
 sg13g2_fill_1 FILLER_22_288 ();
 sg13g2_fill_2 FILLER_22_294 ();
 sg13g2_decap_4 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_333 ();
 sg13g2_decap_4 FILLER_22_347 ();
 sg13g2_fill_2 FILLER_22_359 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_decap_4 FILLER_22_372 ();
 sg13g2_fill_2 FILLER_22_376 ();
 sg13g2_decap_4 FILLER_22_388 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_decap_4 FILLER_22_399 ();
 sg13g2_fill_1 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_2 FILLER_23_19 ();
 sg13g2_fill_2 FILLER_23_25 ();
 sg13g2_decap_4 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_47 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_decap_4 FILLER_23_61 ();
 sg13g2_fill_2 FILLER_23_65 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_107 ();
 sg13g2_decap_4 FILLER_23_114 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_decap_8 FILLER_23_160 ();
 sg13g2_decap_4 FILLER_23_167 ();
 sg13g2_fill_2 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_187 ();
 sg13g2_decap_4 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_198 ();
 sg13g2_fill_2 FILLER_23_204 ();
 sg13g2_decap_8 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_239 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_4 FILLER_23_294 ();
 sg13g2_fill_2 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_decap_4 FILLER_23_368 ();
 sg13g2_decap_4 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_decap_8 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_17 ();
 sg13g2_fill_1 FILLER_24_24 ();
 sg13g2_fill_2 FILLER_24_34 ();
 sg13g2_fill_2 FILLER_24_57 ();
 sg13g2_decap_8 FILLER_24_64 ();
 sg13g2_fill_2 FILLER_24_71 ();
 sg13g2_fill_1 FILLER_24_73 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_106 ();
 sg13g2_fill_1 FILLER_24_108 ();
 sg13g2_decap_4 FILLER_24_135 ();
 sg13g2_fill_2 FILLER_24_143 ();
 sg13g2_fill_2 FILLER_24_150 ();
 sg13g2_fill_1 FILLER_24_152 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_234 ();
 sg13g2_decap_4 FILLER_24_249 ();
 sg13g2_fill_2 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_263 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_4 FILLER_24_285 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_2 FILLER_24_334 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_decap_4 FILLER_24_394 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_27 ();
 sg13g2_fill_1 FILLER_25_34 ();
 sg13g2_fill_2 FILLER_25_57 ();
 sg13g2_fill_2 FILLER_25_64 ();
 sg13g2_decap_8 FILLER_25_82 ();
 sg13g2_decap_8 FILLER_25_93 ();
 sg13g2_decap_8 FILLER_25_100 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_decap_8 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_142 ();
 sg13g2_decap_8 FILLER_25_149 ();
 sg13g2_decap_8 FILLER_25_156 ();
 sg13g2_decap_8 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_235 ();
 sg13g2_fill_2 FILLER_25_242 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_decap_8 FILLER_25_316 ();
 sg13g2_decap_4 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_327 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_decap_4 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_fill_2 FILLER_25_427 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_9 ();
 sg13g2_decap_8 FILLER_26_16 ();
 sg13g2_decap_8 FILLER_26_23 ();
 sg13g2_fill_2 FILLER_26_30 ();
 sg13g2_fill_1 FILLER_26_59 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_65 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_decap_4 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_decap_4 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_170 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_255 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_294 ();
 sg13g2_decap_4 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_347 ();
 sg13g2_fill_2 FILLER_26_354 ();
 sg13g2_decap_4 FILLER_26_371 ();
 sg13g2_decap_4 FILLER_26_388 ();
 sg13g2_fill_1 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_412 ();
 sg13g2_decap_8 FILLER_26_419 ();
 sg13g2_decap_4 FILLER_26_426 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_9 ();
 sg13g2_fill_2 FILLER_27_36 ();
 sg13g2_decap_4 FILLER_27_57 ();
 sg13g2_fill_2 FILLER_27_61 ();
 sg13g2_decap_8 FILLER_27_129 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_decap_8 FILLER_27_143 ();
 sg13g2_fill_1 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_decap_4 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_216 ();
 sg13g2_decap_8 FILLER_27_244 ();
 sg13g2_decap_4 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_255 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_decap_4 FILLER_27_271 ();
 sg13g2_fill_1 FILLER_27_275 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_decap_4 FILLER_27_302 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_324 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_4 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_392 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_36 ();
 sg13g2_fill_1 FILLER_28_38 ();
 sg13g2_decap_4 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_58 ();
 sg13g2_decap_8 FILLER_28_62 ();
 sg13g2_decap_8 FILLER_28_69 ();
 sg13g2_fill_1 FILLER_28_76 ();
 sg13g2_fill_1 FILLER_28_86 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_decap_4 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_103 ();
 sg13g2_fill_2 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_145 ();
 sg13g2_fill_1 FILLER_28_155 ();
 sg13g2_fill_2 FILLER_28_164 ();
 sg13g2_decap_8 FILLER_28_171 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_fill_1 FILLER_28_180 ();
 sg13g2_fill_1 FILLER_28_194 ();
 sg13g2_decap_4 FILLER_28_199 ();
 sg13g2_decap_4 FILLER_28_208 ();
 sg13g2_fill_2 FILLER_28_212 ();
 sg13g2_fill_2 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_decap_8 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_232 ();
 sg13g2_decap_8 FILLER_28_239 ();
 sg13g2_decap_8 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_decap_8 FILLER_28_279 ();
 sg13g2_fill_2 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_fill_2 FILLER_28_310 ();
 sg13g2_decap_8 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_decap_4 FILLER_28_372 ();
 sg13g2_fill_1 FILLER_28_376 ();
 sg13g2_fill_2 FILLER_28_382 ();
 sg13g2_fill_1 FILLER_28_384 ();
 sg13g2_decap_4 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_409 ();
 sg13g2_decap_8 FILLER_28_416 ();
 sg13g2_decap_8 FILLER_28_423 ();
 sg13g2_decap_4 FILLER_29_48 ();
 sg13g2_fill_1 FILLER_29_52 ();
 sg13g2_decap_8 FILLER_29_57 ();
 sg13g2_decap_8 FILLER_29_64 ();
 sg13g2_fill_1 FILLER_29_71 ();
 sg13g2_decap_8 FILLER_29_86 ();
 sg13g2_decap_8 FILLER_29_93 ();
 sg13g2_decap_8 FILLER_29_100 ();
 sg13g2_fill_2 FILLER_29_115 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_174 ();
 sg13g2_decap_8 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_211 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_fill_2 FILLER_29_286 ();
 sg13g2_decap_8 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_29_312 ();
 sg13g2_fill_2 FILLER_29_319 ();
 sg13g2_fill_1 FILLER_29_321 ();
 sg13g2_fill_1 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_fill_2 FILLER_29_368 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_32 ();
 sg13g2_fill_1 FILLER_30_34 ();
 sg13g2_fill_2 FILLER_30_60 ();
 sg13g2_fill_2 FILLER_30_66 ();
 sg13g2_fill_1 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_98 ();
 sg13g2_decap_4 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_116 ();
 sg13g2_decap_8 FILLER_30_134 ();
 sg13g2_decap_8 FILLER_30_141 ();
 sg13g2_decap_8 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_206 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_222 ();
 sg13g2_decap_8 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_262 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_decap_8 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_309 ();
 sg13g2_fill_1 FILLER_30_311 ();
 sg13g2_decap_8 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_341 ();
 sg13g2_decap_8 FILLER_30_348 ();
 sg13g2_decap_4 FILLER_30_355 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_30_412 ();
 sg13g2_decap_8 FILLER_30_419 ();
 sg13g2_decap_4 FILLER_30_426 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_19 ();
 sg13g2_fill_1 FILLER_31_23 ();
 sg13g2_fill_2 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_fill_2 FILLER_31_105 ();
 sg13g2_fill_1 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_125 ();
 sg13g2_decap_8 FILLER_31_132 ();
 sg13g2_decap_4 FILLER_31_139 ();
 sg13g2_decap_4 FILLER_31_151 ();
 sg13g2_fill_1 FILLER_31_155 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_4 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_207 ();
 sg13g2_fill_2 FILLER_31_252 ();
 sg13g2_fill_1 FILLER_31_254 ();
 sg13g2_fill_2 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_31_391 ();
 sg13g2_fill_1 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_16 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_fill_1 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_55 ();
 sg13g2_decap_4 FILLER_32_62 ();
 sg13g2_fill_1 FILLER_32_66 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_fill_1 FILLER_32_102 ();
 sg13g2_fill_1 FILLER_32_118 ();
 sg13g2_fill_1 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_155 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_decap_8 FILLER_32_184 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_226 ();
 sg13g2_decap_8 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_249 ();
 sg13g2_decap_4 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_fill_1 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_404 ();
 sg13g2_decap_8 FILLER_32_411 ();
 sg13g2_decap_8 FILLER_32_418 ();
 sg13g2_decap_4 FILLER_32_425 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_23 ();
 sg13g2_decap_8 FILLER_33_37 ();
 sg13g2_decap_8 FILLER_33_44 ();
 sg13g2_decap_8 FILLER_33_51 ();
 sg13g2_decap_8 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_85 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_118 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_fill_1 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_decap_4 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_2 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_216 ();
 sg13g2_decap_4 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_decap_8 FILLER_33_237 ();
 sg13g2_decap_8 FILLER_33_254 ();
 sg13g2_decap_4 FILLER_33_261 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_decap_4 FILLER_33_375 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_decap_8 FILLER_34_33 ();
 sg13g2_decap_8 FILLER_34_40 ();
 sg13g2_fill_2 FILLER_34_47 ();
 sg13g2_fill_1 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_66 ();
 sg13g2_fill_2 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_89 ();
 sg13g2_fill_2 FILLER_34_96 ();
 sg13g2_fill_1 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_104 ();
 sg13g2_fill_1 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_decap_4 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_197 ();
 sg13g2_decap_8 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_fill_2 FILLER_34_273 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_decap_8 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_307 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_decap_4 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_329 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_372 ();
 sg13g2_fill_2 FILLER_34_384 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_416 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_16 ();
 sg13g2_fill_1 FILLER_35_18 ();
 sg13g2_decap_8 FILLER_35_27 ();
 sg13g2_fill_2 FILLER_35_34 ();
 sg13g2_decap_4 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_fill_1 FILLER_35_109 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_fill_1 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_217 ();
 sg13g2_decap_4 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_227 ();
 sg13g2_decap_4 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_267 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_fill_1 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_fill_2 FILLER_35_390 ();
 sg13g2_fill_1 FILLER_35_392 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_17 ();
 sg13g2_fill_1 FILLER_36_24 ();
 sg13g2_decap_8 FILLER_36_33 ();
 sg13g2_fill_1 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_55 ();
 sg13g2_fill_1 FILLER_36_59 ();
 sg13g2_decap_4 FILLER_36_64 ();
 sg13g2_decap_8 FILLER_36_72 ();
 sg13g2_decap_8 FILLER_36_79 ();
 sg13g2_decap_8 FILLER_36_86 ();
 sg13g2_decap_8 FILLER_36_93 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_decap_8 FILLER_36_107 ();
 sg13g2_decap_8 FILLER_36_114 ();
 sg13g2_decap_8 FILLER_36_137 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_decap_8 FILLER_36_162 ();
 sg13g2_decap_8 FILLER_36_169 ();
 sg13g2_fill_2 FILLER_36_176 ();
 sg13g2_fill_1 FILLER_36_178 ();
 sg13g2_fill_2 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_4 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_233 ();
 sg13g2_decap_8 FILLER_36_240 ();
 sg13g2_fill_2 FILLER_36_251 ();
 sg13g2_decap_4 FILLER_36_268 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_decap_4 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_decap_4 FILLER_36_374 ();
 sg13g2_fill_1 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_36_409 ();
 sg13g2_decap_8 FILLER_36_416 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_22 ();
 sg13g2_decap_4 FILLER_37_29 ();
 sg13g2_fill_1 FILLER_37_33 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_57 ();
 sg13g2_decap_4 FILLER_37_62 ();
 sg13g2_decap_8 FILLER_37_85 ();
 sg13g2_decap_4 FILLER_37_92 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_decap_8 FILLER_37_101 ();
 sg13g2_decap_8 FILLER_37_108 ();
 sg13g2_decap_8 FILLER_37_115 ();
 sg13g2_decap_4 FILLER_37_122 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_141 ();
 sg13g2_decap_4 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_159 ();
 sg13g2_decap_8 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_173 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_fill_2 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_251 ();
 sg13g2_decap_4 FILLER_37_258 ();
 sg13g2_decap_8 FILLER_37_303 ();
 sg13g2_decap_8 FILLER_37_310 ();
 sg13g2_decap_4 FILLER_37_317 ();
 sg13g2_fill_2 FILLER_37_321 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_366 ();
 sg13g2_decap_8 FILLER_37_373 ();
 sg13g2_decap_4 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_384 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_17 ();
 sg13g2_decap_8 FILLER_38_29 ();
 sg13g2_decap_8 FILLER_38_36 ();
 sg13g2_decap_8 FILLER_38_43 ();
 sg13g2_decap_8 FILLER_38_50 ();
 sg13g2_decap_4 FILLER_38_57 ();
 sg13g2_fill_1 FILLER_38_86 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_4 FILLER_38_98 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_decap_8 FILLER_38_111 ();
 sg13g2_decap_8 FILLER_38_118 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_decap_8 FILLER_38_132 ();
 sg13g2_decap_8 FILLER_38_139 ();
 sg13g2_fill_1 FILLER_38_146 ();
 sg13g2_fill_1 FILLER_38_171 ();
 sg13g2_fill_1 FILLER_38_177 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_fill_2 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_decap_8 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_232 ();
 sg13g2_decap_4 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_decap_4 FILLER_38_254 ();
 sg13g2_fill_1 FILLER_38_258 ();
 sg13g2_fill_2 FILLER_38_264 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_302 ();
 sg13g2_decap_8 FILLER_38_309 ();
 sg13g2_fill_1 FILLER_38_316 ();
 sg13g2_decap_4 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_fill_2 FILLER_38_399 ();
 sg13g2_fill_1 FILLER_38_401 ();
 sg13g2_decap_8 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_421 ();
 sg13g2_fill_2 FILLER_38_428 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_18 ();
 sg13g2_fill_1 FILLER_39_20 ();
 sg13g2_decap_4 FILLER_39_29 ();
 sg13g2_fill_2 FILLER_39_33 ();
 sg13g2_decap_4 FILLER_39_40 ();
 sg13g2_fill_1 FILLER_39_44 ();
 sg13g2_fill_2 FILLER_39_80 ();
 sg13g2_fill_1 FILLER_39_123 ();
 sg13g2_decap_4 FILLER_39_132 ();
 sg13g2_fill_2 FILLER_39_136 ();
 sg13g2_fill_2 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_4 FILLER_39_176 ();
 sg13g2_decap_8 FILLER_39_187 ();
 sg13g2_decap_8 FILLER_39_214 ();
 sg13g2_fill_2 FILLER_39_221 ();
 sg13g2_fill_1 FILLER_39_223 ();
 sg13g2_fill_2 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_262 ();
 sg13g2_decap_8 FILLER_39_268 ();
 sg13g2_decap_8 FILLER_39_275 ();
 sg13g2_decap_4 FILLER_39_282 ();
 sg13g2_fill_1 FILLER_39_286 ();
 sg13g2_fill_1 FILLER_39_295 ();
 sg13g2_fill_2 FILLER_39_306 ();
 sg13g2_fill_2 FILLER_39_318 ();
 sg13g2_fill_2 FILLER_39_354 ();
 sg13g2_fill_1 FILLER_39_356 ();
 sg13g2_fill_2 FILLER_39_365 ();
 sg13g2_decap_4 FILLER_39_377 ();
 sg13g2_fill_1 FILLER_39_381 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_decap_4 FILLER_40_30 ();
 sg13g2_decap_4 FILLER_40_55 ();
 sg13g2_fill_1 FILLER_40_59 ();
 sg13g2_fill_1 FILLER_40_82 ();
 sg13g2_fill_1 FILLER_40_106 ();
 sg13g2_fill_2 FILLER_40_111 ();
 sg13g2_decap_8 FILLER_40_118 ();
 sg13g2_fill_2 FILLER_40_154 ();
 sg13g2_fill_1 FILLER_40_156 ();
 sg13g2_decap_8 FILLER_40_166 ();
 sg13g2_decap_4 FILLER_40_173 ();
 sg13g2_fill_2 FILLER_40_177 ();
 sg13g2_fill_2 FILLER_40_200 ();
 sg13g2_fill_1 FILLER_40_205 ();
 sg13g2_fill_1 FILLER_40_219 ();
 sg13g2_fill_2 FILLER_40_259 ();
 sg13g2_fill_2 FILLER_40_271 ();
 sg13g2_decap_4 FILLER_40_281 ();
 sg13g2_decap_4 FILLER_40_289 ();
 sg13g2_fill_1 FILLER_40_293 ();
 sg13g2_fill_2 FILLER_40_304 ();
 sg13g2_decap_4 FILLER_40_320 ();
 sg13g2_fill_2 FILLER_40_324 ();
 sg13g2_decap_8 FILLER_40_338 ();
 sg13g2_fill_1 FILLER_40_345 ();
 sg13g2_decap_4 FILLER_40_355 ();
 sg13g2_decap_4 FILLER_40_363 ();
 sg13g2_decap_4 FILLER_40_377 ();
 sg13g2_fill_1 FILLER_40_392 ();
 sg13g2_fill_1 FILLER_40_403 ();
 sg13g2_decap_8 FILLER_40_412 ();
 sg13g2_decap_8 FILLER_40_419 ();
 sg13g2_decap_4 FILLER_40_426 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_4 ();
 sg13g2_fill_2 FILLER_41_23 ();
 sg13g2_fill_1 FILLER_41_25 ();
 sg13g2_decap_4 FILLER_41_31 ();
 sg13g2_fill_2 FILLER_41_50 ();
 sg13g2_decap_8 FILLER_41_59 ();
 sg13g2_decap_4 FILLER_41_71 ();
 sg13g2_fill_2 FILLER_41_85 ();
 sg13g2_fill_1 FILLER_41_91 ();
 sg13g2_fill_2 FILLER_41_104 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_decap_8 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_129 ();
 sg13g2_fill_1 FILLER_41_136 ();
 sg13g2_fill_2 FILLER_41_145 ();
 sg13g2_fill_1 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_167 ();
 sg13g2_fill_2 FILLER_41_174 ();
 sg13g2_fill_1 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_185 ();
 sg13g2_fill_1 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_fill_1 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_298 ();
 sg13g2_fill_1 FILLER_41_305 ();
 sg13g2_decap_8 FILLER_41_314 ();
 sg13g2_decap_8 FILLER_41_321 ();
 sg13g2_fill_1 FILLER_41_328 ();
 sg13g2_decap_8 FILLER_41_333 ();
 sg13g2_decap_8 FILLER_41_340 ();
 sg13g2_fill_2 FILLER_41_347 ();
 sg13g2_fill_1 FILLER_41_349 ();
 sg13g2_fill_1 FILLER_41_368 ();
 sg13g2_decap_8 FILLER_41_374 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_383 ();
 sg13g2_decap_4 FILLER_41_396 ();
 sg13g2_decap_4 FILLER_41_426 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_9 ();
 sg13g2_fill_2 FILLER_42_13 ();
 sg13g2_fill_2 FILLER_42_19 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_42 ();
 sg13g2_fill_2 FILLER_42_49 ();
 sg13g2_fill_1 FILLER_42_51 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_4 FILLER_42_63 ();
 sg13g2_fill_1 FILLER_42_67 ();
 sg13g2_fill_1 FILLER_42_76 ();
 sg13g2_fill_2 FILLER_42_88 ();
 sg13g2_fill_1 FILLER_42_95 ();
 sg13g2_fill_2 FILLER_42_100 ();
 sg13g2_decap_4 FILLER_42_128 ();
 sg13g2_fill_2 FILLER_42_152 ();
 sg13g2_fill_1 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_170 ();
 sg13g2_decap_8 FILLER_42_177 ();
 sg13g2_fill_2 FILLER_42_184 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_4 FILLER_42_252 ();
 sg13g2_fill_2 FILLER_42_256 ();
 sg13g2_fill_2 FILLER_42_263 ();
 sg13g2_fill_1 FILLER_42_265 ();
 sg13g2_decap_4 FILLER_42_270 ();
 sg13g2_fill_1 FILLER_42_274 ();
 sg13g2_decap_8 FILLER_42_320 ();
 sg13g2_fill_2 FILLER_42_327 ();
 sg13g2_fill_1 FILLER_42_333 ();
 sg13g2_decap_8 FILLER_42_338 ();
 sg13g2_decap_4 FILLER_42_345 ();
 sg13g2_fill_1 FILLER_42_349 ();
 sg13g2_fill_2 FILLER_42_381 ();
 sg13g2_fill_2 FILLER_42_388 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_8 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_42_412 ();
 sg13g2_decap_8 FILLER_42_419 ();
 sg13g2_decap_4 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_11 ();
 sg13g2_decap_4 FILLER_43_28 ();
 sg13g2_fill_2 FILLER_43_32 ();
 sg13g2_decap_8 FILLER_43_39 ();
 sg13g2_decap_4 FILLER_43_46 ();
 sg13g2_fill_2 FILLER_43_53 ();
 sg13g2_fill_1 FILLER_43_60 ();
 sg13g2_decap_8 FILLER_43_65 ();
 sg13g2_decap_8 FILLER_43_76 ();
 sg13g2_decap_8 FILLER_43_83 ();
 sg13g2_decap_8 FILLER_43_90 ();
 sg13g2_decap_8 FILLER_43_97 ();
 sg13g2_decap_8 FILLER_43_104 ();
 sg13g2_decap_8 FILLER_43_111 ();
 sg13g2_decap_8 FILLER_43_118 ();
 sg13g2_fill_1 FILLER_43_125 ();
 sg13g2_fill_1 FILLER_43_152 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_fill_2 FILLER_43_175 ();
 sg13g2_fill_1 FILLER_43_177 ();
 sg13g2_decap_8 FILLER_43_191 ();
 sg13g2_decap_8 FILLER_43_198 ();
 sg13g2_decap_8 FILLER_43_205 ();
 sg13g2_fill_1 FILLER_43_212 ();
 sg13g2_fill_1 FILLER_43_217 ();
 sg13g2_decap_4 FILLER_43_222 ();
 sg13g2_fill_1 FILLER_43_226 ();
 sg13g2_fill_1 FILLER_43_253 ();
 sg13g2_fill_1 FILLER_43_259 ();
 sg13g2_fill_1 FILLER_43_268 ();
 sg13g2_fill_2 FILLER_43_274 ();
 sg13g2_fill_2 FILLER_43_284 ();
 sg13g2_fill_2 FILLER_43_291 ();
 sg13g2_decap_8 FILLER_43_298 ();
 sg13g2_fill_2 FILLER_43_305 ();
 sg13g2_fill_1 FILLER_43_307 ();
 sg13g2_fill_1 FILLER_43_343 ();
 sg13g2_fill_1 FILLER_43_353 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_decap_4 FILLER_43_390 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_4 FILLER_44_21 ();
 sg13g2_fill_1 FILLER_44_25 ();
 sg13g2_decap_8 FILLER_44_31 ();
 sg13g2_fill_1 FILLER_44_38 ();
 sg13g2_fill_2 FILLER_44_44 ();
 sg13g2_fill_1 FILLER_44_60 ();
 sg13g2_decap_8 FILLER_44_69 ();
 sg13g2_decap_4 FILLER_44_76 ();
 sg13g2_fill_2 FILLER_44_80 ();
 sg13g2_decap_8 FILLER_44_85 ();
 sg13g2_decap_8 FILLER_44_92 ();
 sg13g2_decap_8 FILLER_44_99 ();
 sg13g2_fill_2 FILLER_44_114 ();
 sg13g2_decap_8 FILLER_44_124 ();
 sg13g2_fill_2 FILLER_44_131 ();
 sg13g2_decap_4 FILLER_44_138 ();
 sg13g2_fill_1 FILLER_44_142 ();
 sg13g2_decap_8 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_decap_4 FILLER_44_165 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_decap_4 FILLER_44_178 ();
 sg13g2_fill_2 FILLER_44_190 ();
 sg13g2_fill_1 FILLER_44_192 ();
 sg13g2_fill_2 FILLER_44_200 ();
 sg13g2_decap_8 FILLER_44_219 ();
 sg13g2_decap_8 FILLER_44_226 ();
 sg13g2_fill_2 FILLER_44_233 ();
 sg13g2_fill_1 FILLER_44_235 ();
 sg13g2_decap_4 FILLER_44_246 ();
 sg13g2_fill_2 FILLER_44_260 ();
 sg13g2_fill_1 FILLER_44_262 ();
 sg13g2_decap_8 FILLER_44_289 ();
 sg13g2_decap_4 FILLER_44_296 ();
 sg13g2_decap_4 FILLER_44_309 ();
 sg13g2_fill_2 FILLER_44_317 ();
 sg13g2_fill_1 FILLER_44_319 ();
 sg13g2_fill_1 FILLER_44_325 ();
 sg13g2_fill_2 FILLER_44_331 ();
 sg13g2_fill_1 FILLER_44_333 ();
 sg13g2_fill_1 FILLER_44_364 ();
 sg13g2_fill_2 FILLER_44_370 ();
 sg13g2_fill_1 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_23 ();
 sg13g2_fill_1 FILLER_45_29 ();
 sg13g2_fill_1 FILLER_45_65 ();
 sg13g2_decap_4 FILLER_45_70 ();
 sg13g2_fill_1 FILLER_45_74 ();
 sg13g2_fill_1 FILLER_45_86 ();
 sg13g2_fill_2 FILLER_45_96 ();
 sg13g2_fill_1 FILLER_45_98 ();
 sg13g2_fill_1 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_128 ();
 sg13g2_decap_8 FILLER_45_135 ();
 sg13g2_decap_8 FILLER_45_142 ();
 sg13g2_decap_8 FILLER_45_149 ();
 sg13g2_decap_8 FILLER_45_156 ();
 sg13g2_decap_4 FILLER_45_163 ();
 sg13g2_fill_2 FILLER_45_182 ();
 sg13g2_decap_4 FILLER_45_205 ();
 sg13g2_decap_8 FILLER_45_214 ();
 sg13g2_fill_2 FILLER_45_221 ();
 sg13g2_fill_1 FILLER_45_223 ();
 sg13g2_fill_1 FILLER_45_255 ();
 sg13g2_fill_2 FILLER_45_264 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_decap_8 FILLER_45_278 ();
 sg13g2_decap_8 FILLER_45_289 ();
 sg13g2_fill_2 FILLER_45_296 ();
 sg13g2_fill_1 FILLER_45_298 ();
 sg13g2_decap_4 FILLER_45_325 ();
 sg13g2_fill_2 FILLER_45_338 ();
 sg13g2_fill_1 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_355 ();
 sg13g2_decap_8 FILLER_45_362 ();
 sg13g2_fill_2 FILLER_45_369 ();
 sg13g2_fill_1 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_411 ();
 sg13g2_decap_8 FILLER_45_418 ();
 sg13g2_decap_4 FILLER_45_425 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_27 ();
 sg13g2_decap_4 FILLER_46_40 ();
 sg13g2_fill_2 FILLER_46_44 ();
 sg13g2_fill_2 FILLER_46_51 ();
 sg13g2_fill_2 FILLER_46_97 ();
 sg13g2_decap_8 FILLER_46_106 ();
 sg13g2_fill_2 FILLER_46_113 ();
 sg13g2_fill_1 FILLER_46_115 ();
 sg13g2_decap_8 FILLER_46_129 ();
 sg13g2_decap_8 FILLER_46_136 ();
 sg13g2_fill_2 FILLER_46_143 ();
 sg13g2_decap_4 FILLER_46_150 ();
 sg13g2_fill_2 FILLER_46_154 ();
 sg13g2_decap_4 FILLER_46_160 ();
 sg13g2_fill_2 FILLER_46_164 ();
 sg13g2_decap_8 FILLER_46_211 ();
 sg13g2_decap_8 FILLER_46_218 ();
 sg13g2_decap_8 FILLER_46_225 ();
 sg13g2_decap_8 FILLER_46_232 ();
 sg13g2_decap_8 FILLER_46_239 ();
 sg13g2_decap_8 FILLER_46_246 ();
 sg13g2_fill_1 FILLER_46_253 ();
 sg13g2_fill_1 FILLER_46_270 ();
 sg13g2_fill_1 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_286 ();
 sg13g2_decap_8 FILLER_46_293 ();
 sg13g2_decap_8 FILLER_46_300 ();
 sg13g2_fill_1 FILLER_46_307 ();
 sg13g2_decap_4 FILLER_46_313 ();
 sg13g2_fill_2 FILLER_46_317 ();
 sg13g2_fill_2 FILLER_46_327 ();
 sg13g2_decap_4 FILLER_46_335 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_fill_2 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_fill_2 FILLER_46_427 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_40 ();
 sg13g2_fill_2 FILLER_47_44 ();
 sg13g2_fill_2 FILLER_47_65 ();
 sg13g2_fill_1 FILLER_47_67 ();
 sg13g2_fill_2 FILLER_47_74 ();
 sg13g2_fill_1 FILLER_47_76 ();
 sg13g2_fill_1 FILLER_47_82 ();
 sg13g2_fill_1 FILLER_47_97 ();
 sg13g2_fill_2 FILLER_47_111 ();
 sg13g2_fill_1 FILLER_47_113 ();
 sg13g2_decap_4 FILLER_47_129 ();
 sg13g2_fill_2 FILLER_47_162 ();
 sg13g2_decap_8 FILLER_47_197 ();
 sg13g2_decap_4 FILLER_47_204 ();
 sg13g2_decap_8 FILLER_47_212 ();
 sg13g2_decap_4 FILLER_47_219 ();
 sg13g2_fill_2 FILLER_47_223 ();
 sg13g2_decap_4 FILLER_47_251 ();
 sg13g2_fill_2 FILLER_47_255 ();
 sg13g2_fill_1 FILLER_47_298 ();
 sg13g2_decap_8 FILLER_47_303 ();
 sg13g2_decap_4 FILLER_47_323 ();
 sg13g2_fill_1 FILLER_47_327 ();
 sg13g2_fill_1 FILLER_47_333 ();
 sg13g2_fill_2 FILLER_47_344 ();
 sg13g2_fill_2 FILLER_47_382 ();
 sg13g2_fill_1 FILLER_47_389 ();
 sg13g2_decap_8 FILLER_47_395 ();
 sg13g2_fill_2 FILLER_47_402 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_48_7 ();
 sg13g2_fill_2 FILLER_48_11 ();
 sg13g2_fill_2 FILLER_48_26 ();
 sg13g2_decap_8 FILLER_48_33 ();
 sg13g2_fill_2 FILLER_48_40 ();
 sg13g2_decap_8 FILLER_48_54 ();
 sg13g2_decap_4 FILLER_48_61 ();
 sg13g2_decap_8 FILLER_48_73 ();
 sg13g2_decap_4 FILLER_48_80 ();
 sg13g2_fill_2 FILLER_48_84 ();
 sg13g2_fill_1 FILLER_48_105 ();
 sg13g2_decap_4 FILLER_48_145 ();
 sg13g2_decap_8 FILLER_48_157 ();
 sg13g2_decap_8 FILLER_48_164 ();
 sg13g2_fill_2 FILLER_48_171 ();
 sg13g2_fill_1 FILLER_48_173 ();
 sg13g2_decap_8 FILLER_48_188 ();
 sg13g2_decap_4 FILLER_48_195 ();
 sg13g2_fill_1 FILLER_48_199 ();
 sg13g2_decap_4 FILLER_48_250 ();
 sg13g2_fill_1 FILLER_48_254 ();
 sg13g2_fill_2 FILLER_48_265 ();
 sg13g2_fill_1 FILLER_48_276 ();
 sg13g2_decap_4 FILLER_48_286 ();
 sg13g2_fill_2 FILLER_48_298 ();
 sg13g2_fill_1 FILLER_48_300 ();
 sg13g2_fill_1 FILLER_48_323 ();
 sg13g2_fill_2 FILLER_48_329 ();
 sg13g2_fill_2 FILLER_48_337 ();
 sg13g2_fill_1 FILLER_48_339 ();
 sg13g2_fill_1 FILLER_48_344 ();
 sg13g2_fill_2 FILLER_48_350 ();
 sg13g2_fill_2 FILLER_48_360 ();
 sg13g2_fill_1 FILLER_48_362 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_4 ();
 sg13g2_fill_1 FILLER_49_9 ();
 sg13g2_fill_1 FILLER_49_26 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_4 FILLER_49_46 ();
 sg13g2_fill_2 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_57 ();
 sg13g2_decap_8 FILLER_49_66 ();
 sg13g2_decap_4 FILLER_49_73 ();
 sg13g2_fill_2 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_83 ();
 sg13g2_fill_1 FILLER_49_90 ();
 sg13g2_fill_1 FILLER_49_96 ();
 sg13g2_fill_2 FILLER_49_110 ();
 sg13g2_fill_2 FILLER_49_157 ();
 sg13g2_fill_1 FILLER_49_159 ();
 sg13g2_fill_2 FILLER_49_166 ();
 sg13g2_fill_1 FILLER_49_168 ();
 sg13g2_decap_4 FILLER_49_177 ();
 sg13g2_decap_4 FILLER_49_185 ();
 sg13g2_fill_2 FILLER_49_189 ();
 sg13g2_fill_2 FILLER_49_213 ();
 sg13g2_fill_1 FILLER_49_215 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_257 ();
 sg13g2_fill_2 FILLER_49_321 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_fill_2 FILLER_49_364 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_decap_4 FILLER_49_379 ();
 sg13g2_fill_2 FILLER_49_383 ();
 sg13g2_fill_1 FILLER_49_405 ();
 sg13g2_fill_1 FILLER_49_414 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_fill_2 FILLER_49_427 ();
 sg13g2_fill_1 FILLER_49_429 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_fill_1 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_34 ();
 sg13g2_decap_8 FILLER_50_41 ();
 sg13g2_decap_8 FILLER_50_48 ();
 sg13g2_decap_8 FILLER_50_59 ();
 sg13g2_decap_8 FILLER_50_66 ();
 sg13g2_decap_4 FILLER_50_73 ();
 sg13g2_fill_1 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_82 ();
 sg13g2_fill_1 FILLER_50_97 ();
 sg13g2_decap_4 FILLER_50_106 ();
 sg13g2_fill_2 FILLER_50_110 ();
 sg13g2_fill_1 FILLER_50_131 ();
 sg13g2_decap_8 FILLER_50_163 ();
 sg13g2_decap_8 FILLER_50_207 ();
 sg13g2_decap_8 FILLER_50_214 ();
 sg13g2_decap_8 FILLER_50_221 ();
 sg13g2_fill_2 FILLER_50_228 ();
 sg13g2_decap_8 FILLER_50_235 ();
 sg13g2_decap_8 FILLER_50_242 ();
 sg13g2_decap_8 FILLER_50_249 ();
 sg13g2_fill_2 FILLER_50_256 ();
 sg13g2_fill_1 FILLER_50_258 ();
 sg13g2_fill_2 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_274 ();
 sg13g2_decap_4 FILLER_50_285 ();
 sg13g2_fill_1 FILLER_50_289 ();
 sg13g2_fill_1 FILLER_50_302 ();
 sg13g2_decap_4 FILLER_50_308 ();
 sg13g2_fill_2 FILLER_50_317 ();
 sg13g2_decap_8 FILLER_50_356 ();
 sg13g2_decap_8 FILLER_50_363 ();
 sg13g2_decap_8 FILLER_50_370 ();
 sg13g2_decap_8 FILLER_50_377 ();
 sg13g2_decap_8 FILLER_50_384 ();
 sg13g2_fill_2 FILLER_50_391 ();
 sg13g2_fill_1 FILLER_50_393 ();
 sg13g2_decap_8 FILLER_50_404 ();
 sg13g2_decap_8 FILLER_50_411 ();
 sg13g2_decap_8 FILLER_50_418 ();
 sg13g2_decap_4 FILLER_50_425 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_40 ();
 sg13g2_decap_4 FILLER_51_47 ();
 sg13g2_fill_2 FILLER_51_51 ();
 sg13g2_fill_1 FILLER_51_67 ();
 sg13g2_decap_4 FILLER_51_81 ();
 sg13g2_fill_2 FILLER_51_92 ();
 sg13g2_decap_8 FILLER_51_99 ();
 sg13g2_decap_8 FILLER_51_106 ();
 sg13g2_decap_8 FILLER_51_113 ();
 sg13g2_decap_4 FILLER_51_120 ();
 sg13g2_fill_2 FILLER_51_124 ();
 sg13g2_fill_2 FILLER_51_135 ();
 sg13g2_fill_1 FILLER_51_142 ();
 sg13g2_fill_1 FILLER_51_166 ();
 sg13g2_fill_2 FILLER_51_174 ();
 sg13g2_decap_4 FILLER_51_184 ();
 sg13g2_fill_2 FILLER_51_193 ();
 sg13g2_decap_8 FILLER_51_199 ();
 sg13g2_decap_8 FILLER_51_206 ();
 sg13g2_decap_4 FILLER_51_213 ();
 sg13g2_fill_2 FILLER_51_217 ();
 sg13g2_decap_8 FILLER_51_245 ();
 sg13g2_fill_2 FILLER_51_252 ();
 sg13g2_fill_1 FILLER_51_254 ();
 sg13g2_fill_1 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_270 ();
 sg13g2_decap_8 FILLER_51_277 ();
 sg13g2_decap_8 FILLER_51_284 ();
 sg13g2_decap_8 FILLER_51_291 ();
 sg13g2_decap_4 FILLER_51_298 ();
 sg13g2_fill_1 FILLER_51_302 ();
 sg13g2_fill_2 FILLER_51_312 ();
 sg13g2_decap_8 FILLER_51_324 ();
 sg13g2_fill_2 FILLER_51_331 ();
 sg13g2_fill_1 FILLER_51_333 ();
 sg13g2_fill_1 FILLER_51_342 ();
 sg13g2_decap_8 FILLER_51_379 ();
 sg13g2_decap_8 FILLER_51_386 ();
 sg13g2_fill_1 FILLER_51_393 ();
 sg13g2_decap_4 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_2 FILLER_52_21 ();
 sg13g2_fill_1 FILLER_52_23 ();
 sg13g2_decap_8 FILLER_52_32 ();
 sg13g2_decap_8 FILLER_52_39 ();
 sg13g2_decap_4 FILLER_52_46 ();
 sg13g2_fill_2 FILLER_52_58 ();
 sg13g2_decap_4 FILLER_52_100 ();
 sg13g2_fill_2 FILLER_52_104 ();
 sg13g2_decap_8 FILLER_52_122 ();
 sg13g2_decap_8 FILLER_52_129 ();
 sg13g2_decap_8 FILLER_52_136 ();
 sg13g2_decap_8 FILLER_52_143 ();
 sg13g2_decap_4 FILLER_52_150 ();
 sg13g2_decap_4 FILLER_52_175 ();
 sg13g2_fill_2 FILLER_52_179 ();
 sg13g2_decap_4 FILLER_52_185 ();
 sg13g2_decap_8 FILLER_52_195 ();
 sg13g2_decap_8 FILLER_52_202 ();
 sg13g2_decap_4 FILLER_52_209 ();
 sg13g2_fill_2 FILLER_52_213 ();
 sg13g2_decap_8 FILLER_52_267 ();
 sg13g2_decap_4 FILLER_52_274 ();
 sg13g2_fill_1 FILLER_52_278 ();
 sg13g2_fill_2 FILLER_52_341 ();
 sg13g2_fill_1 FILLER_52_343 ();
 sg13g2_decap_8 FILLER_52_390 ();
 sg13g2_decap_8 FILLER_52_397 ();
 sg13g2_decap_8 FILLER_52_404 ();
 sg13g2_decap_8 FILLER_52_411 ();
 sg13g2_decap_8 FILLER_52_418 ();
 sg13g2_decap_4 FILLER_52_425 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_13 ();
 sg13g2_fill_2 FILLER_53_17 ();
 sg13g2_decap_4 FILLER_53_28 ();
 sg13g2_fill_1 FILLER_53_32 ();
 sg13g2_decap_8 FILLER_53_37 ();
 sg13g2_decap_4 FILLER_53_44 ();
 sg13g2_fill_1 FILLER_53_48 ();
 sg13g2_fill_2 FILLER_53_67 ();
 sg13g2_fill_1 FILLER_53_72 ();
 sg13g2_fill_1 FILLER_53_83 ();
 sg13g2_decap_8 FILLER_53_103 ();
 sg13g2_decap_8 FILLER_53_110 ();
 sg13g2_fill_2 FILLER_53_117 ();
 sg13g2_fill_1 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_fill_2 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_141 ();
 sg13g2_decap_8 FILLER_53_148 ();
 sg13g2_fill_1 FILLER_53_155 ();
 sg13g2_decap_4 FILLER_53_160 ();
 sg13g2_fill_1 FILLER_53_164 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_decap_8 FILLER_53_175 ();
 sg13g2_decap_8 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_195 ();
 sg13g2_decap_8 FILLER_53_202 ();
 sg13g2_decap_4 FILLER_53_209 ();
 sg13g2_fill_2 FILLER_53_213 ();
 sg13g2_decap_8 FILLER_53_227 ();
 sg13g2_fill_1 FILLER_53_234 ();
 sg13g2_fill_2 FILLER_53_238 ();
 sg13g2_decap_4 FILLER_53_276 ();
 sg13g2_decap_4 FILLER_53_285 ();
 sg13g2_fill_1 FILLER_53_289 ();
 sg13g2_fill_1 FILLER_53_305 ();
 sg13g2_decap_8 FILLER_53_316 ();
 sg13g2_fill_2 FILLER_53_323 ();
 sg13g2_fill_1 FILLER_53_325 ();
 sg13g2_decap_4 FILLER_53_336 ();
 sg13g2_fill_2 FILLER_53_340 ();
 sg13g2_fill_1 FILLER_53_364 ();
 sg13g2_fill_2 FILLER_53_369 ();
 sg13g2_fill_2 FILLER_53_379 ();
 sg13g2_fill_2 FILLER_53_391 ();
 sg13g2_fill_1 FILLER_53_393 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_4 ();
 sg13g2_decap_4 FILLER_54_12 ();
 sg13g2_fill_1 FILLER_54_16 ();
 sg13g2_decap_8 FILLER_54_32 ();
 sg13g2_decap_8 FILLER_54_39 ();
 sg13g2_decap_4 FILLER_54_46 ();
 sg13g2_decap_8 FILLER_54_58 ();
 sg13g2_decap_4 FILLER_54_65 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_fill_2 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_96 ();
 sg13g2_decap_8 FILLER_54_103 ();
 sg13g2_decap_8 FILLER_54_110 ();
 sg13g2_fill_2 FILLER_54_117 ();
 sg13g2_decap_8 FILLER_54_159 ();
 sg13g2_fill_1 FILLER_54_166 ();
 sg13g2_fill_2 FILLER_54_171 ();
 sg13g2_decap_8 FILLER_54_179 ();
 sg13g2_decap_8 FILLER_54_186 ();
 sg13g2_decap_8 FILLER_54_193 ();
 sg13g2_fill_2 FILLER_54_200 ();
 sg13g2_fill_1 FILLER_54_202 ();
 sg13g2_fill_2 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_241 ();
 sg13g2_decap_8 FILLER_54_245 ();
 sg13g2_decap_8 FILLER_54_252 ();
 sg13g2_decap_4 FILLER_54_259 ();
 sg13g2_fill_2 FILLER_54_263 ();
 sg13g2_fill_1 FILLER_54_275 ();
 sg13g2_fill_1 FILLER_54_281 ();
 sg13g2_fill_1 FILLER_54_308 ();
 sg13g2_fill_2 FILLER_54_335 ();
 sg13g2_fill_1 FILLER_54_337 ();
 sg13g2_decap_4 FILLER_54_348 ();
 sg13g2_decap_4 FILLER_54_378 ();
 sg13g2_fill_1 FILLER_54_382 ();
 sg13g2_fill_1 FILLER_54_393 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_9 ();
 sg13g2_fill_2 FILLER_55_23 ();
 sg13g2_decap_8 FILLER_55_48 ();
 sg13g2_decap_8 FILLER_55_55 ();
 sg13g2_decap_8 FILLER_55_62 ();
 sg13g2_decap_8 FILLER_55_69 ();
 sg13g2_decap_8 FILLER_55_76 ();
 sg13g2_fill_2 FILLER_55_83 ();
 sg13g2_fill_1 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_95 ();
 sg13g2_decap_8 FILLER_55_101 ();
 sg13g2_decap_8 FILLER_55_108 ();
 sg13g2_fill_2 FILLER_55_115 ();
 sg13g2_fill_1 FILLER_55_129 ();
 sg13g2_decap_8 FILLER_55_138 ();
 sg13g2_decap_8 FILLER_55_145 ();
 sg13g2_decap_8 FILLER_55_152 ();
 sg13g2_fill_1 FILLER_55_164 ();
 sg13g2_decap_4 FILLER_55_170 ();
 sg13g2_decap_8 FILLER_55_200 ();
 sg13g2_decap_8 FILLER_55_207 ();
 sg13g2_decap_8 FILLER_55_214 ();
 sg13g2_fill_2 FILLER_55_221 ();
 sg13g2_fill_1 FILLER_55_223 ();
 sg13g2_fill_1 FILLER_55_232 ();
 sg13g2_decap_8 FILLER_55_237 ();
 sg13g2_decap_8 FILLER_55_244 ();
 sg13g2_decap_8 FILLER_55_251 ();
 sg13g2_decap_8 FILLER_55_266 ();
 sg13g2_decap_4 FILLER_55_278 ();
 sg13g2_fill_2 FILLER_55_291 ();
 sg13g2_fill_2 FILLER_55_321 ();
 sg13g2_fill_2 FILLER_55_333 ();
 sg13g2_fill_2 FILLER_55_349 ();
 sg13g2_fill_2 FILLER_55_356 ();
 sg13g2_fill_2 FILLER_55_363 ();
 sg13g2_fill_1 FILLER_55_365 ();
 sg13g2_decap_4 FILLER_55_402 ();
 sg13g2_decap_8 FILLER_55_411 ();
 sg13g2_decap_8 FILLER_55_418 ();
 sg13g2_decap_4 FILLER_55_425 ();
 sg13g2_fill_1 FILLER_55_429 ();
 sg13g2_fill_2 FILLER_56_23 ();
 sg13g2_fill_2 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_67 ();
 sg13g2_fill_2 FILLER_56_88 ();
 sg13g2_fill_1 FILLER_56_90 ();
 sg13g2_fill_2 FILLER_56_100 ();
 sg13g2_fill_2 FILLER_56_107 ();
 sg13g2_fill_2 FILLER_56_126 ();
 sg13g2_fill_1 FILLER_56_128 ();
 sg13g2_decap_4 FILLER_56_134 ();
 sg13g2_fill_1 FILLER_56_138 ();
 sg13g2_decap_4 FILLER_56_185 ();
 sg13g2_decap_4 FILLER_56_194 ();
 sg13g2_decap_4 FILLER_56_206 ();
 sg13g2_decap_4 FILLER_56_218 ();
 sg13g2_fill_2 FILLER_56_222 ();
 sg13g2_decap_8 FILLER_56_233 ();
 sg13g2_decap_8 FILLER_56_240 ();
 sg13g2_decap_8 FILLER_56_247 ();
 sg13g2_decap_8 FILLER_56_254 ();
 sg13g2_decap_8 FILLER_56_261 ();
 sg13g2_decap_8 FILLER_56_268 ();
 sg13g2_decap_8 FILLER_56_275 ();
 sg13g2_decap_8 FILLER_56_282 ();
 sg13g2_decap_8 FILLER_56_289 ();
 sg13g2_decap_8 FILLER_56_296 ();
 sg13g2_decap_8 FILLER_56_303 ();
 sg13g2_decap_8 FILLER_56_310 ();
 sg13g2_decap_8 FILLER_56_317 ();
 sg13g2_decap_8 FILLER_56_324 ();
 sg13g2_decap_8 FILLER_56_331 ();
 sg13g2_decap_8 FILLER_56_364 ();
 sg13g2_decap_8 FILLER_56_371 ();
 sg13g2_decap_4 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_56_415 ();
 sg13g2_decap_8 FILLER_56_422 ();
 sg13g2_fill_1 FILLER_56_429 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_16 ();
 sg13g2_fill_2 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_34 ();
 sg13g2_decap_8 FILLER_57_41 ();
 sg13g2_decap_8 FILLER_57_48 ();
 sg13g2_decap_8 FILLER_57_55 ();
 sg13g2_decap_8 FILLER_57_62 ();
 sg13g2_decap_8 FILLER_57_69 ();
 sg13g2_decap_4 FILLER_57_76 ();
 sg13g2_fill_2 FILLER_57_97 ();
 sg13g2_fill_1 FILLER_57_130 ();
 sg13g2_fill_2 FILLER_57_135 ();
 sg13g2_fill_2 FILLER_57_141 ();
 sg13g2_fill_2 FILLER_57_146 ();
 sg13g2_fill_1 FILLER_57_148 ();
 sg13g2_decap_4 FILLER_57_167 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_182 ();
 sg13g2_fill_2 FILLER_57_188 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_4 FILLER_57_224 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_decap_8 FILLER_57_248 ();
 sg13g2_fill_1 FILLER_57_255 ();
 sg13g2_fill_2 FILLER_57_265 ();
 sg13g2_fill_1 FILLER_57_303 ();
 sg13g2_decap_8 FILLER_57_314 ();
 sg13g2_decap_8 FILLER_57_347 ();
 sg13g2_decap_8 FILLER_57_354 ();
 sg13g2_decap_8 FILLER_57_361 ();
 sg13g2_decap_8 FILLER_57_368 ();
 sg13g2_decap_4 FILLER_57_375 ();
 sg13g2_fill_1 FILLER_57_379 ();
 sg13g2_decap_8 FILLER_57_388 ();
 sg13g2_decap_8 FILLER_57_395 ();
 sg13g2_decap_8 FILLER_57_402 ();
 sg13g2_decap_8 FILLER_57_409 ();
 sg13g2_decap_8 FILLER_57_416 ();
 sg13g2_decap_8 FILLER_57_423 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_4 FILLER_58_14 ();
 sg13g2_fill_1 FILLER_58_18 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_4 FILLER_58_35 ();
 sg13g2_fill_2 FILLER_58_39 ();
 sg13g2_fill_1 FILLER_58_52 ();
 sg13g2_fill_2 FILLER_58_119 ();
 sg13g2_fill_1 FILLER_58_136 ();
 sg13g2_decap_8 FILLER_58_164 ();
 sg13g2_decap_8 FILLER_58_171 ();
 sg13g2_decap_4 FILLER_58_193 ();
 sg13g2_fill_1 FILLER_58_202 ();
 sg13g2_decap_8 FILLER_58_216 ();
 sg13g2_decap_8 FILLER_58_223 ();
 sg13g2_fill_2 FILLER_58_230 ();
 sg13g2_fill_1 FILLER_58_232 ();
 sg13g2_fill_2 FILLER_58_246 ();
 sg13g2_decap_8 FILLER_58_337 ();
 sg13g2_decap_8 FILLER_58_344 ();
 sg13g2_decap_8 FILLER_58_351 ();
 sg13g2_decap_8 FILLER_58_358 ();
 sg13g2_decap_4 FILLER_58_365 ();
 sg13g2_decap_8 FILLER_59_26 ();
 sg13g2_decap_8 FILLER_59_68 ();
 sg13g2_fill_1 FILLER_59_75 ();
 sg13g2_decap_8 FILLER_59_80 ();
 sg13g2_fill_2 FILLER_59_87 ();
 sg13g2_fill_2 FILLER_59_97 ();
 sg13g2_decap_8 FILLER_59_108 ();
 sg13g2_decap_8 FILLER_59_115 ();
 sg13g2_fill_2 FILLER_59_122 ();
 sg13g2_fill_1 FILLER_59_124 ();
 sg13g2_decap_8 FILLER_59_130 ();
 sg13g2_fill_1 FILLER_59_137 ();
 sg13g2_decap_8 FILLER_59_143 ();
 sg13g2_fill_1 FILLER_59_150 ();
 sg13g2_decap_8 FILLER_59_156 ();
 sg13g2_decap_8 FILLER_59_163 ();
 sg13g2_decap_8 FILLER_59_170 ();
 sg13g2_decap_8 FILLER_59_177 ();
 sg13g2_decap_8 FILLER_59_184 ();
 sg13g2_decap_8 FILLER_59_191 ();
 sg13g2_fill_1 FILLER_59_198 ();
 sg13g2_decap_4 FILLER_59_259 ();
 sg13g2_fill_1 FILLER_59_271 ();
 sg13g2_fill_1 FILLER_59_282 ();
 sg13g2_fill_1 FILLER_59_288 ();
 sg13g2_decap_8 FILLER_59_341 ();
 sg13g2_decap_8 FILLER_59_348 ();
 sg13g2_fill_2 FILLER_59_355 ();
 sg13g2_fill_1 FILLER_59_392 ();
 sg13g2_fill_2 FILLER_59_402 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_14 ();
 sg13g2_fill_1 FILLER_60_18 ();
 sg13g2_decap_8 FILLER_60_54 ();
 sg13g2_decap_8 FILLER_60_61 ();
 sg13g2_decap_8 FILLER_60_68 ();
 sg13g2_decap_8 FILLER_60_75 ();
 sg13g2_fill_2 FILLER_60_82 ();
 sg13g2_decap_4 FILLER_60_94 ();
 sg13g2_fill_2 FILLER_60_101 ();
 sg13g2_fill_1 FILLER_60_103 ();
 sg13g2_decap_8 FILLER_60_134 ();
 sg13g2_fill_2 FILLER_60_141 ();
 sg13g2_decap_8 FILLER_60_179 ();
 sg13g2_decap_4 FILLER_60_192 ();
 sg13g2_decap_8 FILLER_60_206 ();
 sg13g2_decap_8 FILLER_60_213 ();
 sg13g2_decap_8 FILLER_60_220 ();
 sg13g2_fill_1 FILLER_60_227 ();
 sg13g2_decap_4 FILLER_60_241 ();
 sg13g2_fill_1 FILLER_60_245 ();
 sg13g2_fill_1 FILLER_60_250 ();
 sg13g2_decap_4 FILLER_60_260 ();
 sg13g2_fill_2 FILLER_60_274 ();
 sg13g2_fill_1 FILLER_60_276 ();
 sg13g2_fill_1 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_324 ();
 sg13g2_decap_8 FILLER_60_331 ();
 sg13g2_decap_8 FILLER_60_338 ();
 sg13g2_decap_8 FILLER_60_345 ();
 sg13g2_decap_4 FILLER_60_352 ();
 sg13g2_fill_1 FILLER_60_356 ();
 sg13g2_decap_8 FILLER_60_361 ();
 sg13g2_fill_2 FILLER_60_368 ();
 sg13g2_fill_1 FILLER_60_370 ();
 sg13g2_decap_4 FILLER_60_424 ();
 sg13g2_fill_2 FILLER_60_428 ();
 sg13g2_decap_8 FILLER_61_26 ();
 sg13g2_decap_8 FILLER_61_33 ();
 sg13g2_decap_8 FILLER_61_40 ();
 sg13g2_decap_8 FILLER_61_47 ();
 sg13g2_decap_8 FILLER_61_54 ();
 sg13g2_decap_4 FILLER_61_61 ();
 sg13g2_fill_1 FILLER_61_65 ();
 sg13g2_decap_8 FILLER_61_92 ();
 sg13g2_decap_8 FILLER_61_99 ();
 sg13g2_decap_8 FILLER_61_106 ();
 sg13g2_decap_8 FILLER_61_113 ();
 sg13g2_decap_4 FILLER_61_120 ();
 sg13g2_fill_1 FILLER_61_124 ();
 sg13g2_fill_1 FILLER_61_151 ();
 sg13g2_fill_1 FILLER_61_183 ();
 sg13g2_fill_1 FILLER_61_191 ();
 sg13g2_fill_2 FILLER_61_199 ();
 sg13g2_decap_4 FILLER_61_205 ();
 sg13g2_fill_2 FILLER_61_209 ();
 sg13g2_fill_2 FILLER_61_237 ();
 sg13g2_decap_8 FILLER_61_243 ();
 sg13g2_decap_8 FILLER_61_250 ();
 sg13g2_decap_8 FILLER_61_257 ();
 sg13g2_fill_1 FILLER_61_264 ();
 sg13g2_decap_8 FILLER_61_270 ();
 sg13g2_decap_4 FILLER_61_277 ();
 sg13g2_fill_1 FILLER_61_281 ();
 sg13g2_decap_8 FILLER_61_290 ();
 sg13g2_decap_8 FILLER_61_297 ();
 sg13g2_decap_8 FILLER_61_304 ();
 sg13g2_decap_8 FILLER_61_311 ();
 sg13g2_decap_4 FILLER_61_344 ();
 sg13g2_fill_2 FILLER_61_348 ();
 sg13g2_decap_4 FILLER_61_381 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_4 FILLER_62_19 ();
 sg13g2_decap_8 FILLER_62_27 ();
 sg13g2_decap_4 FILLER_62_34 ();
 sg13g2_decap_8 FILLER_62_64 ();
 sg13g2_decap_4 FILLER_62_71 ();
 sg13g2_fill_1 FILLER_62_108 ();
 sg13g2_decap_8 FILLER_62_124 ();
 sg13g2_decap_8 FILLER_62_131 ();
 sg13g2_fill_2 FILLER_62_138 ();
 sg13g2_fill_1 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_205 ();
 sg13g2_decap_4 FILLER_62_212 ();
 sg13g2_fill_1 FILLER_62_216 ();
 sg13g2_decap_8 FILLER_62_223 ();
 sg13g2_fill_2 FILLER_62_230 ();
 sg13g2_fill_1 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_242 ();
 sg13g2_fill_2 FILLER_62_256 ();
 sg13g2_decap_8 FILLER_62_262 ();
 sg13g2_decap_4 FILLER_62_269 ();
 sg13g2_fill_1 FILLER_62_273 ();
 sg13g2_decap_8 FILLER_62_300 ();
 sg13g2_decap_8 FILLER_62_307 ();
 sg13g2_fill_2 FILLER_62_314 ();
 sg13g2_fill_1 FILLER_62_316 ();
 sg13g2_decap_8 FILLER_62_325 ();
 sg13g2_decap_4 FILLER_62_332 ();
 sg13g2_fill_2 FILLER_62_336 ();
 sg13g2_decap_4 FILLER_62_373 ();
 sg13g2_decap_8 FILLER_62_382 ();
 sg13g2_decap_8 FILLER_62_389 ();
 sg13g2_decap_8 FILLER_62_406 ();
 sg13g2_decap_8 FILLER_62_413 ();
 sg13g2_decap_8 FILLER_62_420 ();
 sg13g2_fill_2 FILLER_62_427 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_2 ();
 sg13g2_decap_8 FILLER_63_29 ();
 sg13g2_decap_4 FILLER_63_36 ();
 sg13g2_fill_1 FILLER_63_40 ();
 sg13g2_fill_2 FILLER_63_46 ();
 sg13g2_fill_1 FILLER_63_48 ();
 sg13g2_decap_4 FILLER_63_54 ();
 sg13g2_decap_8 FILLER_63_62 ();
 sg13g2_decap_8 FILLER_63_69 ();
 sg13g2_decap_8 FILLER_63_76 ();
 sg13g2_decap_8 FILLER_63_83 ();
 sg13g2_decap_8 FILLER_63_90 ();
 sg13g2_decap_8 FILLER_63_97 ();
 sg13g2_decap_4 FILLER_63_104 ();
 sg13g2_fill_1 FILLER_63_108 ();
 sg13g2_decap_4 FILLER_63_151 ();
 sg13g2_decap_8 FILLER_63_159 ();
 sg13g2_decap_4 FILLER_63_166 ();
 sg13g2_fill_2 FILLER_63_170 ();
 sg13g2_decap_8 FILLER_63_176 ();
 sg13g2_fill_1 FILLER_63_183 ();
 sg13g2_fill_1 FILLER_63_245 ();
 sg13g2_fill_1 FILLER_63_250 ();
 sg13g2_decap_8 FILLER_63_260 ();
 sg13g2_decap_4 FILLER_63_267 ();
 sg13g2_fill_1 FILLER_63_271 ();
 sg13g2_decap_8 FILLER_63_277 ();
 sg13g2_decap_8 FILLER_63_284 ();
 sg13g2_decap_8 FILLER_63_291 ();
 sg13g2_decap_4 FILLER_63_302 ();
 sg13g2_fill_1 FILLER_63_306 ();
 sg13g2_decap_4 FILLER_63_359 ();
 sg13g2_fill_1 FILLER_63_363 ();
 sg13g2_fill_1 FILLER_63_369 ();
 sg13g2_decap_8 FILLER_63_396 ();
 sg13g2_fill_1 FILLER_63_403 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_11 ();
 sg13g2_fill_2 FILLER_64_31 ();
 sg13g2_fill_1 FILLER_64_33 ();
 sg13g2_decap_8 FILLER_64_59 ();
 sg13g2_decap_8 FILLER_64_97 ();
 sg13g2_decap_8 FILLER_64_104 ();
 sg13g2_decap_8 FILLER_64_111 ();
 sg13g2_decap_8 FILLER_64_118 ();
 sg13g2_fill_2 FILLER_64_129 ();
 sg13g2_decap_8 FILLER_64_157 ();
 sg13g2_decap_4 FILLER_64_164 ();
 sg13g2_decap_8 FILLER_64_178 ();
 sg13g2_decap_8 FILLER_64_185 ();
 sg13g2_decap_4 FILLER_64_192 ();
 sg13g2_decap_8 FILLER_64_200 ();
 sg13g2_decap_8 FILLER_64_207 ();
 sg13g2_decap_4 FILLER_64_214 ();
 sg13g2_decap_4 FILLER_64_228 ();
 sg13g2_fill_2 FILLER_64_232 ();
 sg13g2_decap_4 FILLER_64_239 ();
 sg13g2_fill_1 FILLER_64_243 ();
 sg13g2_decap_4 FILLER_64_247 ();
 sg13g2_fill_1 FILLER_64_251 ();
 sg13g2_decap_8 FILLER_64_256 ();
 sg13g2_fill_2 FILLER_64_263 ();
 sg13g2_fill_1 FILLER_64_265 ();
 sg13g2_decap_8 FILLER_64_306 ();
 sg13g2_decap_4 FILLER_64_313 ();
 sg13g2_fill_1 FILLER_64_317 ();
 sg13g2_fill_2 FILLER_64_323 ();
 sg13g2_decap_4 FILLER_64_334 ();
 sg13g2_fill_1 FILLER_64_338 ();
 sg13g2_decap_8 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_358 ();
 sg13g2_decap_8 FILLER_64_365 ();
 sg13g2_fill_2 FILLER_64_372 ();
 sg13g2_fill_1 FILLER_64_374 ();
 sg13g2_decap_8 FILLER_64_379 ();
 sg13g2_fill_2 FILLER_64_386 ();
 sg13g2_fill_1 FILLER_64_388 ();
 sg13g2_decap_4 FILLER_64_424 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_16 ();
 sg13g2_decap_4 FILLER_65_29 ();
 sg13g2_fill_2 FILLER_65_33 ();
 sg13g2_fill_2 FILLER_65_85 ();
 sg13g2_decap_4 FILLER_65_99 ();
 sg13g2_decap_8 FILLER_65_107 ();
 sg13g2_decap_4 FILLER_65_114 ();
 sg13g2_fill_1 FILLER_65_118 ();
 sg13g2_decap_8 FILLER_65_124 ();
 sg13g2_decap_4 FILLER_65_131 ();
 sg13g2_fill_2 FILLER_65_135 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_fill_2 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_177 ();
 sg13g2_fill_1 FILLER_65_184 ();
 sg13g2_decap_8 FILLER_65_200 ();
 sg13g2_decap_8 FILLER_65_207 ();
 sg13g2_decap_8 FILLER_65_214 ();
 sg13g2_decap_4 FILLER_65_221 ();
 sg13g2_fill_1 FILLER_65_225 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_fill_1 FILLER_65_259 ();
 sg13g2_fill_1 FILLER_65_275 ();
 sg13g2_decap_8 FILLER_65_284 ();
 sg13g2_decap_8 FILLER_65_291 ();
 sg13g2_decap_4 FILLER_65_298 ();
 sg13g2_fill_1 FILLER_65_302 ();
 sg13g2_decap_8 FILLER_65_313 ();
 sg13g2_decap_4 FILLER_65_320 ();
 sg13g2_fill_2 FILLER_65_324 ();
 sg13g2_fill_2 FILLER_65_335 ();
 sg13g2_decap_8 FILLER_65_413 ();
 sg13g2_decap_8 FILLER_65_420 ();
 sg13g2_fill_2 FILLER_65_427 ();
 sg13g2_fill_1 FILLER_65_429 ();
 sg13g2_fill_2 FILLER_66_31 ();
 sg13g2_fill_1 FILLER_66_33 ();
 sg13g2_decap_4 FILLER_66_44 ();
 sg13g2_fill_2 FILLER_66_53 ();
 sg13g2_decap_8 FILLER_66_69 ();
 sg13g2_fill_2 FILLER_66_76 ();
 sg13g2_fill_1 FILLER_66_85 ();
 sg13g2_decap_4 FILLER_66_90 ();
 sg13g2_fill_1 FILLER_66_94 ();
 sg13g2_decap_8 FILLER_66_129 ();
 sg13g2_fill_1 FILLER_66_136 ();
 sg13g2_fill_2 FILLER_66_163 ();
 sg13g2_fill_1 FILLER_66_165 ();
 sg13g2_decap_4 FILLER_66_222 ();
 sg13g2_decap_8 FILLER_66_229 ();
 sg13g2_decap_4 FILLER_66_236 ();
 sg13g2_decap_8 FILLER_66_245 ();
 sg13g2_fill_2 FILLER_66_252 ();
 sg13g2_fill_1 FILLER_66_254 ();
 sg13g2_fill_1 FILLER_66_260 ();
 sg13g2_decap_8 FILLER_66_265 ();
 sg13g2_decap_8 FILLER_66_282 ();
 sg13g2_fill_1 FILLER_66_289 ();
 sg13g2_decap_8 FILLER_66_321 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_fill_2 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_341 ();
 sg13g2_decap_8 FILLER_66_352 ();
 sg13g2_decap_8 FILLER_66_369 ();
 sg13g2_fill_2 FILLER_66_376 ();
 sg13g2_decap_8 FILLER_66_393 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_2 ();
 sg13g2_fill_1 FILLER_67_21 ();
 sg13g2_decap_4 FILLER_67_32 ();
 sg13g2_fill_1 FILLER_67_36 ();
 sg13g2_decap_8 FILLER_67_40 ();
 sg13g2_decap_8 FILLER_67_51 ();
 sg13g2_fill_2 FILLER_67_58 ();
 sg13g2_fill_2 FILLER_67_100 ();
 sg13g2_fill_1 FILLER_67_102 ();
 sg13g2_decap_8 FILLER_67_136 ();
 sg13g2_fill_2 FILLER_67_143 ();
 sg13g2_fill_1 FILLER_67_145 ();
 sg13g2_decap_4 FILLER_67_185 ();
 sg13g2_fill_1 FILLER_67_189 ();
 sg13g2_decap_4 FILLER_67_223 ();
 sg13g2_fill_2 FILLER_67_227 ();
 sg13g2_decap_4 FILLER_67_255 ();
 sg13g2_fill_1 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_265 ();
 sg13g2_decap_4 FILLER_67_272 ();
 sg13g2_fill_2 FILLER_67_276 ();
 sg13g2_decap_8 FILLER_67_304 ();
 sg13g2_decap_4 FILLER_67_311 ();
 sg13g2_fill_1 FILLER_67_315 ();
 sg13g2_decap_8 FILLER_67_368 ();
 sg13g2_decap_4 FILLER_67_375 ();
 sg13g2_fill_2 FILLER_67_379 ();
 sg13g2_decap_4 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_67_421 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_4 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_11 ();
 sg13g2_decap_8 FILLER_68_16 ();
 sg13g2_decap_4 FILLER_68_23 ();
 sg13g2_fill_2 FILLER_68_27 ();
 sg13g2_decap_8 FILLER_68_59 ();
 sg13g2_fill_2 FILLER_68_66 ();
 sg13g2_fill_1 FILLER_68_68 ();
 sg13g2_decap_8 FILLER_68_73 ();
 sg13g2_decap_8 FILLER_68_85 ();
 sg13g2_fill_2 FILLER_68_92 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_4 FILLER_68_105 ();
 sg13g2_fill_1 FILLER_68_109 ();
 sg13g2_decap_4 FILLER_68_120 ();
 sg13g2_fill_2 FILLER_68_124 ();
 sg13g2_fill_2 FILLER_68_133 ();
 sg13g2_fill_1 FILLER_68_135 ();
 sg13g2_fill_2 FILLER_68_141 ();
 sg13g2_fill_1 FILLER_68_143 ();
 sg13g2_decap_4 FILLER_68_149 ();
 sg13g2_fill_1 FILLER_68_153 ();
 sg13g2_decap_4 FILLER_68_158 ();
 sg13g2_fill_1 FILLER_68_167 ();
 sg13g2_decap_8 FILLER_68_185 ();
 sg13g2_fill_2 FILLER_68_192 ();
 sg13g2_decap_4 FILLER_68_201 ();
 sg13g2_fill_1 FILLER_68_205 ();
 sg13g2_fill_2 FILLER_68_232 ();
 sg13g2_fill_2 FILLER_68_260 ();
 sg13g2_fill_1 FILLER_68_262 ();
 sg13g2_fill_2 FILLER_68_273 ();
 sg13g2_fill_2 FILLER_68_301 ();
 sg13g2_fill_2 FILLER_68_329 ();
 sg13g2_fill_1 FILLER_68_331 ();
 sg13g2_fill_1 FILLER_68_358 ();
 sg13g2_fill_2 FILLER_68_367 ();
 sg13g2_fill_1 FILLER_68_369 ();
 sg13g2_fill_1 FILLER_68_375 ();
 sg13g2_decap_4 FILLER_68_402 ();
 sg13g2_fill_1 FILLER_68_406 ();
 sg13g2_decap_8 FILLER_68_415 ();
 sg13g2_decap_8 FILLER_68_422 ();
 sg13g2_fill_1 FILLER_68_429 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_decap_4 FILLER_69_30 ();
 sg13g2_fill_1 FILLER_69_34 ();
 sg13g2_fill_2 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_54 ();
 sg13g2_decap_8 FILLER_69_61 ();
 sg13g2_decap_8 FILLER_69_68 ();
 sg13g2_decap_8 FILLER_69_75 ();
 sg13g2_decap_8 FILLER_69_82 ();
 sg13g2_decap_4 FILLER_69_89 ();
 sg13g2_fill_2 FILLER_69_93 ();
 sg13g2_decap_8 FILLER_69_99 ();
 sg13g2_decap_8 FILLER_69_106 ();
 sg13g2_fill_1 FILLER_69_113 ();
 sg13g2_decap_8 FILLER_69_145 ();
 sg13g2_decap_8 FILLER_69_152 ();
 sg13g2_decap_4 FILLER_69_159 ();
 sg13g2_fill_1 FILLER_69_163 ();
 sg13g2_decap_8 FILLER_69_177 ();
 sg13g2_decap_8 FILLER_69_184 ();
 sg13g2_decap_8 FILLER_69_191 ();
 sg13g2_decap_8 FILLER_69_198 ();
 sg13g2_decap_8 FILLER_69_213 ();
 sg13g2_decap_8 FILLER_69_220 ();
 sg13g2_decap_4 FILLER_69_227 ();
 sg13g2_decap_8 FILLER_69_236 ();
 sg13g2_decap_4 FILLER_69_243 ();
 sg13g2_fill_1 FILLER_69_247 ();
 sg13g2_decap_8 FILLER_69_258 ();
 sg13g2_decap_8 FILLER_69_265 ();
 sg13g2_decap_8 FILLER_69_272 ();
 sg13g2_decap_8 FILLER_69_279 ();
 sg13g2_decap_8 FILLER_69_286 ();
 sg13g2_fill_2 FILLER_69_293 ();
 sg13g2_fill_1 FILLER_69_295 ();
 sg13g2_fill_1 FILLER_69_306 ();
 sg13g2_fill_1 FILLER_69_316 ();
 sg13g2_fill_2 FILLER_69_327 ();
 sg13g2_fill_1 FILLER_69_329 ();
 sg13g2_decap_8 FILLER_69_335 ();
 sg13g2_decap_8 FILLER_69_342 ();
 sg13g2_decap_4 FILLER_69_384 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_8 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_69_412 ();
 sg13g2_decap_8 FILLER_69_419 ();
 sg13g2_decap_4 FILLER_69_426 ();
 sg13g2_decap_4 FILLER_70_42 ();
 sg13g2_fill_1 FILLER_70_50 ();
 sg13g2_fill_1 FILLER_70_90 ();
 sg13g2_decap_4 FILLER_70_96 ();
 sg13g2_fill_2 FILLER_70_100 ();
 sg13g2_decap_8 FILLER_70_111 ();
 sg13g2_decap_8 FILLER_70_118 ();
 sg13g2_fill_1 FILLER_70_125 ();
 sg13g2_fill_2 FILLER_70_181 ();
 sg13g2_fill_1 FILLER_70_183 ();
 sg13g2_decap_8 FILLER_70_207 ();
 sg13g2_decap_8 FILLER_70_214 ();
 sg13g2_decap_8 FILLER_70_221 ();
 sg13g2_decap_8 FILLER_70_228 ();
 sg13g2_decap_4 FILLER_70_235 ();
 sg13g2_decap_8 FILLER_70_243 ();
 sg13g2_decap_8 FILLER_70_250 ();
 sg13g2_decap_8 FILLER_70_257 ();
 sg13g2_fill_1 FILLER_70_264 ();
 sg13g2_decap_8 FILLER_70_291 ();
 sg13g2_decap_8 FILLER_70_298 ();
 sg13g2_decap_8 FILLER_70_305 ();
 sg13g2_decap_8 FILLER_70_312 ();
 sg13g2_decap_8 FILLER_70_319 ();
 sg13g2_fill_1 FILLER_70_326 ();
 sg13g2_fill_2 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_347 ();
 sg13g2_decap_8 FILLER_70_354 ();
 sg13g2_decap_8 FILLER_70_361 ();
 sg13g2_fill_2 FILLER_70_368 ();
 sg13g2_decap_8 FILLER_70_379 ();
 sg13g2_decap_8 FILLER_70_386 ();
 sg13g2_decap_8 FILLER_70_393 ();
 sg13g2_decap_8 FILLER_70_400 ();
 sg13g2_decap_8 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_70_414 ();
 sg13g2_decap_8 FILLER_70_421 ();
 sg13g2_fill_2 FILLER_70_428 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_9 ();
 sg13g2_decap_8 FILLER_71_27 ();
 sg13g2_decap_8 FILLER_71_34 ();
 sg13g2_decap_8 FILLER_71_41 ();
 sg13g2_fill_1 FILLER_71_72 ();
 sg13g2_fill_1 FILLER_71_78 ();
 sg13g2_fill_1 FILLER_71_88 ();
 sg13g2_decap_8 FILLER_71_129 ();
 sg13g2_decap_4 FILLER_71_136 ();
 sg13g2_fill_1 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_145 ();
 sg13g2_fill_2 FILLER_71_160 ();
 sg13g2_fill_1 FILLER_71_162 ();
 sg13g2_fill_2 FILLER_71_170 ();
 sg13g2_fill_1 FILLER_71_172 ();
 sg13g2_fill_2 FILLER_71_178 ();
 sg13g2_fill_1 FILLER_71_180 ();
 sg13g2_fill_2 FILLER_71_188 ();
 sg13g2_decap_8 FILLER_71_200 ();
 sg13g2_fill_2 FILLER_71_207 ();
 sg13g2_decap_8 FILLER_71_214 ();
 sg13g2_decap_4 FILLER_71_221 ();
 sg13g2_fill_1 FILLER_71_225 ();
 sg13g2_decap_8 FILLER_71_272 ();
 sg13g2_decap_8 FILLER_71_279 ();
 sg13g2_decap_8 FILLER_71_286 ();
 sg13g2_fill_2 FILLER_71_293 ();
 sg13g2_fill_1 FILLER_71_300 ();
 sg13g2_decap_4 FILLER_71_315 ();
 sg13g2_fill_1 FILLER_71_319 ();
 sg13g2_decap_4 FILLER_71_346 ();
 sg13g2_fill_1 FILLER_71_350 ();
 sg13g2_fill_2 FILLER_71_377 ();
 sg13g2_decap_8 FILLER_71_405 ();
 sg13g2_decap_8 FILLER_71_412 ();
 sg13g2_decap_8 FILLER_71_423 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_4 FILLER_72_7 ();
 sg13g2_decap_4 FILLER_72_16 ();
 sg13g2_fill_1 FILLER_72_20 ();
 sg13g2_fill_2 FILLER_72_26 ();
 sg13g2_decap_8 FILLER_72_32 ();
 sg13g2_decap_4 FILLER_72_39 ();
 sg13g2_fill_2 FILLER_72_62 ();
 sg13g2_fill_2 FILLER_72_90 ();
 sg13g2_fill_2 FILLER_72_97 ();
 sg13g2_fill_1 FILLER_72_99 ();
 sg13g2_fill_1 FILLER_72_104 ();
 sg13g2_fill_2 FILLER_72_110 ();
 sg13g2_fill_1 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_139 ();
 sg13g2_decap_8 FILLER_72_146 ();
 sg13g2_decap_8 FILLER_72_153 ();
 sg13g2_decap_4 FILLER_72_160 ();
 sg13g2_fill_1 FILLER_72_185 ();
 sg13g2_fill_1 FILLER_72_191 ();
 sg13g2_fill_1 FILLER_72_197 ();
 sg13g2_fill_1 FILLER_72_219 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_fill_1 FILLER_72_248 ();
 sg13g2_decap_4 FILLER_72_259 ();
 sg13g2_fill_1 FILLER_72_263 ();
 sg13g2_decap_8 FILLER_72_290 ();
 sg13g2_decap_4 FILLER_72_297 ();
 sg13g2_decap_8 FILLER_72_337 ();
 sg13g2_decap_8 FILLER_72_344 ();
 sg13g2_decap_4 FILLER_72_351 ();
 sg13g2_fill_1 FILLER_72_363 ();
 sg13g2_fill_2 FILLER_72_368 ();
 sg13g2_decap_4 FILLER_72_380 ();
 sg13g2_fill_2 FILLER_72_384 ();
 sg13g2_decap_4 FILLER_72_395 ();
 sg13g2_fill_1 FILLER_72_399 ();
 sg13g2_fill_1 FILLER_73_31 ();
 sg13g2_fill_1 FILLER_73_58 ();
 sg13g2_fill_2 FILLER_73_72 ();
 sg13g2_fill_1 FILLER_73_74 ();
 sg13g2_fill_1 FILLER_73_80 ();
 sg13g2_fill_2 FILLER_73_86 ();
 sg13g2_decap_8 FILLER_73_92 ();
 sg13g2_decap_4 FILLER_73_99 ();
 sg13g2_decap_8 FILLER_73_110 ();
 sg13g2_decap_8 FILLER_73_117 ();
 sg13g2_decap_8 FILLER_73_124 ();
 sg13g2_decap_4 FILLER_73_131 ();
 sg13g2_fill_2 FILLER_73_139 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_169 ();
 sg13g2_fill_2 FILLER_73_176 ();
 sg13g2_decap_8 FILLER_73_187 ();
 sg13g2_fill_1 FILLER_73_194 ();
 sg13g2_decap_4 FILLER_73_199 ();
 sg13g2_fill_2 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_218 ();
 sg13g2_fill_2 FILLER_73_251 ();
 sg13g2_decap_8 FILLER_73_279 ();
 sg13g2_fill_1 FILLER_73_286 ();
 sg13g2_fill_2 FILLER_73_339 ();
 sg13g2_fill_1 FILLER_73_341 ();
 sg13g2_fill_2 FILLER_73_347 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_fill_2 FILLER_73_366 ();
 sg13g2_fill_1 FILLER_73_368 ();
 sg13g2_fill_2 FILLER_73_416 ();
 sg13g2_decap_8 FILLER_73_422 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_fill_1 FILLER_74_11 ();
 sg13g2_decap_4 FILLER_74_16 ();
 sg13g2_decap_4 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_39 ();
 sg13g2_decap_8 FILLER_74_62 ();
 sg13g2_fill_1 FILLER_74_69 ();
 sg13g2_fill_1 FILLER_74_86 ();
 sg13g2_fill_2 FILLER_74_105 ();
 sg13g2_fill_1 FILLER_74_107 ();
 sg13g2_fill_1 FILLER_74_112 ();
 sg13g2_fill_1 FILLER_74_117 ();
 sg13g2_fill_1 FILLER_74_144 ();
 sg13g2_fill_1 FILLER_74_149 ();
 sg13g2_fill_2 FILLER_74_154 ();
 sg13g2_fill_1 FILLER_74_156 ();
 sg13g2_fill_1 FILLER_74_167 ();
 sg13g2_decap_8 FILLER_74_172 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_decap_4 FILLER_74_202 ();
 sg13g2_decap_8 FILLER_74_236 ();
 sg13g2_decap_4 FILLER_74_279 ();
 sg13g2_fill_2 FILLER_74_283 ();
 sg13g2_decap_4 FILLER_74_311 ();
 sg13g2_fill_1 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_342 ();
 sg13g2_decap_8 FILLER_74_349 ();
 sg13g2_decap_8 FILLER_74_356 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_decap_8 FILLER_74_375 ();
 sg13g2_decap_4 FILLER_74_382 ();
 sg13g2_fill_1 FILLER_74_386 ();
 sg13g2_fill_2 FILLER_74_401 ();
 sg13g2_fill_1 FILLER_74_403 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_4 FILLER_75_7 ();
 sg13g2_fill_1 FILLER_75_20 ();
 sg13g2_fill_2 FILLER_75_33 ();
 sg13g2_fill_1 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_41 ();
 sg13g2_decap_8 FILLER_75_48 ();
 sg13g2_fill_2 FILLER_75_55 ();
 sg13g2_fill_1 FILLER_75_57 ();
 sg13g2_decap_8 FILLER_75_67 ();
 sg13g2_decap_4 FILLER_75_74 ();
 sg13g2_fill_1 FILLER_75_78 ();
 sg13g2_fill_1 FILLER_75_84 ();
 sg13g2_decap_4 FILLER_75_89 ();
 sg13g2_fill_1 FILLER_75_101 ();
 sg13g2_fill_2 FILLER_75_121 ();
 sg13g2_fill_2 FILLER_75_129 ();
 sg13g2_fill_1 FILLER_75_131 ();
 sg13g2_fill_2 FILLER_75_136 ();
 sg13g2_fill_1 FILLER_75_138 ();
 sg13g2_decap_8 FILLER_75_170 ();
 sg13g2_decap_8 FILLER_75_177 ();
 sg13g2_decap_8 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_191 ();
 sg13g2_decap_8 FILLER_75_212 ();
 sg13g2_decap_8 FILLER_75_219 ();
 sg13g2_decap_8 FILLER_75_226 ();
 sg13g2_decap_8 FILLER_75_233 ();
 sg13g2_decap_8 FILLER_75_240 ();
 sg13g2_decap_8 FILLER_75_247 ();
 sg13g2_decap_8 FILLER_75_254 ();
 sg13g2_decap_8 FILLER_75_261 ();
 sg13g2_decap_8 FILLER_75_268 ();
 sg13g2_decap_4 FILLER_75_275 ();
 sg13g2_fill_1 FILLER_75_279 ();
 sg13g2_decap_8 FILLER_75_285 ();
 sg13g2_decap_8 FILLER_75_292 ();
 sg13g2_decap_8 FILLER_75_299 ();
 sg13g2_decap_8 FILLER_75_306 ();
 sg13g2_decap_8 FILLER_75_313 ();
 sg13g2_decap_8 FILLER_75_320 ();
 sg13g2_decap_4 FILLER_75_327 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_decap_8 FILLER_75_358 ();
 sg13g2_decap_4 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_369 ();
 sg13g2_fill_1 FILLER_75_396 ();
 sg13g2_fill_1 FILLER_75_402 ();
 sg13g2_decap_8 FILLER_75_418 ();
 sg13g2_decap_4 FILLER_75_425 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_19 ();
 sg13g2_fill_1 FILLER_76_25 ();
 sg13g2_fill_2 FILLER_76_34 ();
 sg13g2_fill_1 FILLER_76_36 ();
 sg13g2_decap_8 FILLER_76_50 ();
 sg13g2_fill_2 FILLER_76_57 ();
 sg13g2_fill_1 FILLER_76_59 ();
 sg13g2_fill_1 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_118 ();
 sg13g2_decap_8 FILLER_76_125 ();
 sg13g2_decap_8 FILLER_76_132 ();
 sg13g2_decap_4 FILLER_76_139 ();
 sg13g2_fill_2 FILLER_76_143 ();
 sg13g2_fill_1 FILLER_76_149 ();
 sg13g2_fill_2 FILLER_76_177 ();
 sg13g2_fill_1 FILLER_76_179 ();
 sg13g2_fill_1 FILLER_76_185 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_fill_2 FILLER_76_238 ();
 sg13g2_decap_4 FILLER_76_260 ();
 sg13g2_fill_1 FILLER_76_264 ();
 sg13g2_fill_1 FILLER_76_275 ();
 sg13g2_decap_8 FILLER_76_305 ();
 sg13g2_decap_8 FILLER_76_312 ();
 sg13g2_decap_8 FILLER_76_319 ();
 sg13g2_decap_8 FILLER_76_326 ();
 sg13g2_decap_8 FILLER_76_333 ();
 sg13g2_decap_4 FILLER_76_344 ();
 sg13g2_fill_2 FILLER_76_348 ();
 sg13g2_decap_8 FILLER_76_354 ();
 sg13g2_decap_8 FILLER_76_361 ();
 sg13g2_decap_4 FILLER_76_368 ();
 sg13g2_decap_4 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_415 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_fill_2 FILLER_77_40 ();
 sg13g2_fill_1 FILLER_77_42 ();
 sg13g2_decap_4 FILLER_77_52 ();
 sg13g2_fill_1 FILLER_77_75 ();
 sg13g2_fill_1 FILLER_77_80 ();
 sg13g2_fill_1 FILLER_77_86 ();
 sg13g2_decap_4 FILLER_77_98 ();
 sg13g2_fill_1 FILLER_77_102 ();
 sg13g2_fill_1 FILLER_77_108 ();
 sg13g2_fill_2 FILLER_77_140 ();
 sg13g2_decap_4 FILLER_77_168 ();
 sg13g2_fill_2 FILLER_77_186 ();
 sg13g2_fill_1 FILLER_77_188 ();
 sg13g2_fill_2 FILLER_77_212 ();
 sg13g2_fill_1 FILLER_77_214 ();
 sg13g2_decap_8 FILLER_77_261 ();
 sg13g2_decap_4 FILLER_77_268 ();
 sg13g2_fill_1 FILLER_77_272 ();
 sg13g2_fill_1 FILLER_77_283 ();
 sg13g2_decap_8 FILLER_77_310 ();
 sg13g2_decap_8 FILLER_77_373 ();
 sg13g2_decap_8 FILLER_77_380 ();
 sg13g2_fill_1 FILLER_77_395 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_27 ();
 sg13g2_fill_2 FILLER_78_33 ();
 sg13g2_decap_8 FILLER_78_40 ();
 sg13g2_fill_2 FILLER_78_47 ();
 sg13g2_fill_2 FILLER_78_53 ();
 sg13g2_fill_1 FILLER_78_55 ();
 sg13g2_decap_4 FILLER_78_63 ();
 sg13g2_fill_1 FILLER_78_67 ();
 sg13g2_fill_1 FILLER_78_76 ();
 sg13g2_fill_1 FILLER_78_85 ();
 sg13g2_fill_2 FILLER_78_95 ();
 sg13g2_fill_1 FILLER_78_101 ();
 sg13g2_fill_1 FILLER_78_107 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_4 FILLER_78_154 ();
 sg13g2_fill_2 FILLER_78_158 ();
 sg13g2_fill_2 FILLER_78_176 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_fill_2 FILLER_78_189 ();
 sg13g2_fill_1 FILLER_78_191 ();
 sg13g2_fill_1 FILLER_78_202 ();
 sg13g2_decap_8 FILLER_78_285 ();
 sg13g2_decap_8 FILLER_78_292 ();
 sg13g2_decap_8 FILLER_78_299 ();
 sg13g2_fill_2 FILLER_78_310 ();
 sg13g2_fill_1 FILLER_78_346 ();
 sg13g2_fill_2 FILLER_78_352 ();
 sg13g2_fill_1 FILLER_78_366 ();
 sg13g2_decap_4 FILLER_78_400 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_51 ();
 sg13g2_fill_2 FILLER_79_78 ();
 sg13g2_fill_2 FILLER_79_106 ();
 sg13g2_fill_1 FILLER_79_108 ();
 sg13g2_decap_8 FILLER_79_117 ();
 sg13g2_decap_8 FILLER_79_124 ();
 sg13g2_decap_4 FILLER_79_131 ();
 sg13g2_decap_4 FILLER_79_139 ();
 sg13g2_decap_8 FILLER_79_151 ();
 sg13g2_fill_1 FILLER_79_158 ();
 sg13g2_decap_4 FILLER_79_163 ();
 sg13g2_fill_2 FILLER_79_167 ();
 sg13g2_fill_1 FILLER_79_173 ();
 sg13g2_fill_1 FILLER_79_204 ();
 sg13g2_decap_4 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_239 ();
 sg13g2_decap_8 FILLER_79_246 ();
 sg13g2_fill_2 FILLER_79_253 ();
 sg13g2_fill_2 FILLER_79_295 ();
 sg13g2_fill_1 FILLER_79_297 ();
 sg13g2_fill_2 FILLER_79_324 ();
 sg13g2_fill_2 FILLER_79_404 ();
 sg13g2_decap_4 FILLER_79_414 ();
 sg13g2_fill_1 FILLER_79_418 ();
 sg13g2_fill_2 FILLER_79_427 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_4 FILLER_80_81 ();
 sg13g2_fill_2 FILLER_80_113 ();
 sg13g2_fill_1 FILLER_80_119 ();
 sg13g2_fill_2 FILLER_80_128 ();
 sg13g2_fill_1 FILLER_80_130 ();
 sg13g2_fill_2 FILLER_80_139 ();
 sg13g2_fill_1 FILLER_80_141 ();
 sg13g2_fill_1 FILLER_80_150 ();
 sg13g2_fill_2 FILLER_80_159 ();
 sg13g2_decap_4 FILLER_80_173 ();
 sg13g2_fill_1 FILLER_80_193 ();
 sg13g2_decap_8 FILLER_80_198 ();
 sg13g2_decap_4 FILLER_80_205 ();
 sg13g2_fill_2 FILLER_80_209 ();
 sg13g2_fill_1 FILLER_80_219 ();
 sg13g2_decap_4 FILLER_80_224 ();
 sg13g2_decap_8 FILLER_80_240 ();
 sg13g2_decap_8 FILLER_80_247 ();
 sg13g2_fill_2 FILLER_80_254 ();
 sg13g2_fill_1 FILLER_80_260 ();
 sg13g2_decap_8 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_280 ();
 sg13g2_fill_1 FILLER_80_310 ();
 sg13g2_fill_2 FILLER_80_323 ();
 sg13g2_decap_4 FILLER_80_329 ();
 sg13g2_fill_1 FILLER_80_333 ();
 sg13g2_decap_8 FILLER_80_354 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_4 FILLER_80_368 ();
 sg13g2_decap_8 FILLER_80_376 ();
 sg13g2_fill_1 FILLER_80_383 ();
 sg13g2_decap_4 FILLER_80_408 ();
 sg13g2_decap_8 FILLER_80_420 ();
 sg13g2_fill_2 FILLER_80_427 ();
 sg13g2_fill_1 FILLER_80_429 ();
endmodule
