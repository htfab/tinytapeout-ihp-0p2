module tt_um_digital_clock_example (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire clknet_0_clk;
 wire net60;
 wire \desk_clock.clk_gen_inst.i_refclk ;
 wire \desk_clock.clk_gen_inst.refclk_div[0] ;
 wire \desk_clock.clk_gen_inst.refclk_div[10] ;
 wire \desk_clock.clk_gen_inst.refclk_div[11] ;
 wire \desk_clock.clk_gen_inst.refclk_div[12] ;
 wire \desk_clock.clk_gen_inst.refclk_div[13] ;
 wire \desk_clock.clk_gen_inst.refclk_div[14] ;
 wire \desk_clock.clk_gen_inst.refclk_div[1] ;
 wire \desk_clock.clk_gen_inst.refclk_div[2] ;
 wire \desk_clock.clk_gen_inst.refclk_div[3] ;
 wire \desk_clock.clk_gen_inst.refclk_div[4] ;
 wire \desk_clock.clk_gen_inst.refclk_div[5] ;
 wire \desk_clock.clk_gen_inst.refclk_div[6] ;
 wire \desk_clock.clk_gen_inst.refclk_div[7] ;
 wire \desk_clock.clk_gen_inst.refclk_div[8] ;
 wire \desk_clock.clk_gen_inst.refclk_div[9] ;
 wire \desk_clock.clk_gen_inst.stb_gen_1hz.sig_hold ;
 wire \desk_clock.clk_gen_inst.stb_gen_debounce_clk.sig_hold ;
 wire \desk_clock.clk_gen_inst.stb_gen_fast_clk.sig_hold ;
 wire \desk_clock.clk_gen_inst.stb_gen_refclk.sig_hold ;
 wire \desk_clock.clk_gen_inst.stb_gen_slow_clk.sig_hold ;
 wire \desk_clock.clk_hours[0] ;
 wire \desk_clock.clk_hours[1] ;
 wire \desk_clock.clk_hours[2] ;
 wire \desk_clock.clk_hours[3] ;
 wire \desk_clock.clk_hours[4] ;
 wire \desk_clock.clk_minutes[0] ;
 wire \desk_clock.clk_minutes[1] ;
 wire \desk_clock.clk_minutes[2] ;
 wire \desk_clock.clk_minutes[3] ;
 wire \desk_clock.clk_minutes[4] ;
 wire \desk_clock.clk_minutes[5] ;
 wire \desk_clock.clk_seconds[0] ;
 wire \desk_clock.clk_seconds[1] ;
 wire \desk_clock.clk_seconds[2] ;
 wire \desk_clock.clk_seconds[3] ;
 wire \desk_clock.clk_seconds[4] ;
 wire \desk_clock.clk_seconds[5] ;
 wire \desk_clock.display_control_inst.display_update ;
 wire \desk_clock.display_control_inst.o_write_config ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[0] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[1] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[2] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[3] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[4] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[0] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[1] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[2] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[3] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[4] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[5] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[0] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[1] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[2] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[3] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[4] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[5] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[0] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[10] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[11] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[12] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[13] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[14] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[15] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[1] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[2] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[3] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[4] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[5] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[6] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[7] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[8] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[9] ;
 wire \desk_clock.display_inst.disp_driver.i_addr[0] ;
 wire \desk_clock.display_inst.disp_driver.i_addr[1] ;
 wire \desk_clock.display_inst.disp_driver.i_addr[2] ;
 wire \desk_clock.display_inst.disp_driver.i_addr[3] ;
 wire \desk_clock.display_inst.disp_driver.i_data[0] ;
 wire \desk_clock.display_inst.disp_driver.i_data[1] ;
 wire \desk_clock.display_inst.disp_driver.i_data[2] ;
 wire \desk_clock.display_inst.disp_driver.i_data[3] ;
 wire \desk_clock.display_inst.disp_driver.i_data[4] ;
 wire \desk_clock.display_inst.disp_driver.i_data[7] ;
 wire \desk_clock.display_inst.disp_driver.o_serial_clk ;
 wire \desk_clock.display_inst.disp_driver.o_serial_load ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[0] ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[1] ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[2] ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[3] ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[4] ;
 wire \desk_clock.display_inst.display_settings.transfer_state[0] ;
 wire \desk_clock.display_inst.display_settings.transfer_state[1] ;
 wire \desk_clock.display_inst.display_settings.transfer_state[2] ;
 wire \desk_clock.display_inst.display_settings.transfer_state[3] ;
 wire \desk_clock.display_inst.display_settings.write_config ;
 wire \desk_clock.display_inst.state[0] ;
 wire \desk_clock.display_inst.state[1] ;
 wire \desk_clock.display_inst.state[2] ;
 wire \desk_clock.display_inst.state[3] ;
 wire \desk_clock.input_debounce.fast_set_reg[0] ;
 wire \desk_clock.input_debounce.fast_set_reg[1] ;
 wire \desk_clock.input_debounce.fast_set_reg[2] ;
 wire \desk_clock.input_debounce.fast_set_reg[3] ;
 wire \desk_clock.input_debounce.fast_set_reg[4] ;
 wire \desk_clock.input_debounce.fast_set_reg[5] ;
 wire \desk_clock.input_debounce.set_hours_reg[0] ;
 wire \desk_clock.input_debounce.set_hours_reg[1] ;
 wire \desk_clock.input_debounce.set_hours_reg[2] ;
 wire \desk_clock.input_debounce.set_hours_reg[3] ;
 wire \desk_clock.input_debounce.set_hours_reg[4] ;
 wire \desk_clock.input_debounce.set_hours_reg[5] ;
 wire \desk_clock.input_debounce.set_minutes_reg[0] ;
 wire \desk_clock.input_debounce.set_minutes_reg[1] ;
 wire \desk_clock.input_debounce.set_minutes_reg[2] ;
 wire \desk_clock.input_debounce.set_minutes_reg[3] ;
 wire \desk_clock.input_debounce.set_minutes_reg[4] ;
 wire \desk_clock.input_debounce.set_minutes_reg[5] ;
 wire \desk_clock.refclk_sync_inst.refclk_sync_reg[0] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_inv_1 _0712_ (.Y(_0121_),
    .A(\desk_clock.display_inst.display_settings.write_config ));
 sg13g2_buf_1 _0713_ (.A(\desk_clock.display_inst.state[1] ),
    .X(_0122_));
 sg13g2_buf_1 _0714_ (.A(\desk_clock.display_inst.state[0] ),
    .X(_0123_));
 sg13g2_or3_1 _0715_ (.A(\desk_clock.display_inst.state[2] ),
    .B(net40),
    .C(net39),
    .X(_0124_));
 sg13g2_buf_1 _0716_ (.A(_0124_),
    .X(_0125_));
 sg13g2_buf_1 _0717_ (.A(\desk_clock.display_inst.state[2] ),
    .X(_0126_));
 sg13g2_nand3_1 _0718_ (.B(_0122_),
    .C(net39),
    .A(_0126_),
    .Y(_0127_));
 sg13g2_buf_1 _0719_ (.A(\desk_clock.display_inst.state[3] ),
    .X(_0128_));
 sg13g2_a21oi_2 _0720_ (.B1(_0128_),
    .Y(_0129_),
    .A2(_0127_),
    .A1(_0125_));
 sg13g2_buf_2 _0721_ (.A(\desk_clock.display_inst.display_settings.transfer_state[3] ),
    .X(_0130_));
 sg13g2_buf_1 _0722_ (.A(\desk_clock.display_inst.display_settings.transfer_state[0] ),
    .X(_0131_));
 sg13g2_nor3_2 _0723_ (.A(\desk_clock.display_inst.display_settings.transfer_state[2] ),
    .B(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .C(net37),
    .Y(_0132_));
 sg13g2_and3_1 _0724_ (.X(_0133_),
    .A(\desk_clock.display_inst.display_settings.transfer_state[2] ),
    .B(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .C(\desk_clock.display_inst.display_settings.transfer_state[0] ));
 sg13g2_nor3_2 _0725_ (.A(_0130_),
    .B(_0132_),
    .C(_0133_),
    .Y(_0134_));
 sg13g2_nor2_2 _0726_ (.A(_0129_),
    .B(_0134_),
    .Y(_0135_));
 sg13g2_nand2_1 _0727_ (.Y(_0136_),
    .A(\desk_clock.display_control_inst.o_write_config ),
    .B(_0135_));
 sg13g2_o21ai_1 _0728_ (.B1(_0136_),
    .Y(_0079_),
    .A1(_0121_),
    .A2(_0135_));
 sg13g2_buf_1 _0729_ (.A(rst_n),
    .X(_0137_));
 sg13g2_inv_2 _0730_ (.Y(_0138_),
    .A(_0137_));
 sg13g2_a21o_1 _0731_ (.A2(\desk_clock.clk_hours[4] ),
    .A1(\desk_clock.clk_hours[3] ),
    .B1(_0138_),
    .X(_0139_));
 sg13g2_and4_1 _0732_ (.A(\desk_clock.input_debounce.set_minutes_reg[0] ),
    .B(\desk_clock.input_debounce.set_minutes_reg[3] ),
    .C(\desk_clock.input_debounce.set_minutes_reg[2] ),
    .D(\desk_clock.input_debounce.set_minutes_reg[4] ),
    .X(_0140_));
 sg13g2_nand2_2 _0733_ (.Y(_0141_),
    .A(\desk_clock.input_debounce.set_minutes_reg[1] ),
    .B(_0140_));
 sg13g2_nor2b_2 _0734_ (.A(\desk_clock.clk_gen_inst.stb_gen_1hz.sig_hold ),
    .B_N(\desk_clock.clk_gen_inst.refclk_div[14] ),
    .Y(_0142_));
 sg13g2_and2_1 _0735_ (.A(\desk_clock.clk_seconds[0] ),
    .B(\desk_clock.clk_seconds[1] ),
    .X(_0143_));
 sg13g2_a21oi_1 _0736_ (.A1(_0142_),
    .A2(_0143_),
    .Y(_0144_),
    .B1(\desk_clock.clk_seconds[2] ));
 sg13g2_nand4_1 _0737_ (.B(\desk_clock.clk_seconds[4] ),
    .C(\desk_clock.clk_seconds[3] ),
    .A(\desk_clock.clk_seconds[5] ),
    .Y(_0145_),
    .D(_0142_));
 sg13g2_buf_2 _0738_ (.A(\desk_clock.clk_minutes[0] ),
    .X(_0146_));
 sg13g2_a21oi_1 _0739_ (.A1(\desk_clock.clk_minutes[1] ),
    .A2(_0146_),
    .Y(_0147_),
    .B1(\desk_clock.clk_minutes[2] ));
 sg13g2_nand3_1 _0740_ (.B(\desk_clock.clk_minutes[4] ),
    .C(\desk_clock.clk_minutes[3] ),
    .A(\desk_clock.clk_minutes[5] ),
    .Y(_0148_));
 sg13g2_nor4_2 _0741_ (.A(_0144_),
    .B(_0145_),
    .C(_0147_),
    .Y(_0149_),
    .D(_0148_));
 sg13g2_inv_1 _0742_ (.Y(_0150_),
    .A(\desk_clock.clk_gen_inst.stb_gen_fast_clk.sig_hold ));
 sg13g2_and4_1 _0743_ (.A(\desk_clock.input_debounce.fast_set_reg[0] ),
    .B(\desk_clock.input_debounce.fast_set_reg[3] ),
    .C(\desk_clock.input_debounce.fast_set_reg[2] ),
    .D(\desk_clock.input_debounce.fast_set_reg[4] ),
    .X(_0151_));
 sg13g2_nand4_1 _0744_ (.B(\desk_clock.clk_gen_inst.refclk_div[11] ),
    .C(_0150_),
    .A(\desk_clock.input_debounce.fast_set_reg[1] ),
    .Y(_0152_),
    .D(_0151_));
 sg13g2_nand2b_1 _0745_ (.Y(_0153_),
    .B(\desk_clock.clk_gen_inst.refclk_div[13] ),
    .A_N(\desk_clock.clk_gen_inst.stb_gen_slow_clk.sig_hold ));
 sg13g2_a21o_1 _0746_ (.A2(_0151_),
    .A1(\desk_clock.input_debounce.fast_set_reg[1] ),
    .B1(_0153_),
    .X(_0154_));
 sg13g2_nand2_1 _0747_ (.Y(_0155_),
    .A(_0152_),
    .B(_0154_));
 sg13g2_inv_1 _0748_ (.Y(_0156_),
    .A(\desk_clock.input_debounce.set_hours_reg[1] ));
 sg13g2_nand4_1 _0749_ (.B(\desk_clock.input_debounce.set_hours_reg[3] ),
    .C(\desk_clock.input_debounce.set_hours_reg[2] ),
    .A(\desk_clock.input_debounce.set_hours_reg[0] ),
    .Y(_0157_),
    .D(\desk_clock.input_debounce.set_hours_reg[4] ));
 sg13g2_nor2_2 _0750_ (.A(_0156_),
    .B(_0157_),
    .Y(_0158_));
 sg13g2_mux2_1 _0751_ (.A0(_0149_),
    .A1(_0155_),
    .S(_0158_),
    .X(_0159_));
 sg13g2_nand2_1 _0752_ (.Y(_0160_),
    .A(_0141_),
    .B(_0159_));
 sg13g2_xor2_1 _0753_ (.B(_0160_),
    .A(\desk_clock.clk_hours[0] ),
    .X(_0161_));
 sg13g2_nor2_1 _0754_ (.A(_0139_),
    .B(_0161_),
    .Y(_0026_));
 sg13g2_nand3_1 _0755_ (.B(_0141_),
    .C(_0159_),
    .A(\desk_clock.clk_hours[0] ),
    .Y(_0162_));
 sg13g2_xor2_1 _0756_ (.B(_0162_),
    .A(\desk_clock.clk_hours[1] ),
    .X(_0163_));
 sg13g2_nor2_1 _0757_ (.A(_0139_),
    .B(_0163_),
    .Y(_0027_));
 sg13g2_and2_1 _0758_ (.A(\desk_clock.clk_hours[1] ),
    .B(\desk_clock.clk_hours[0] ),
    .X(_0164_));
 sg13g2_nand3_1 _0759_ (.B(_0159_),
    .C(_0164_),
    .A(_0141_),
    .Y(_0165_));
 sg13g2_xor2_1 _0760_ (.B(_0165_),
    .A(\desk_clock.clk_hours[2] ),
    .X(_0166_));
 sg13g2_nor2_1 _0761_ (.A(_0139_),
    .B(_0166_),
    .Y(_0028_));
 sg13g2_buf_2 _0762_ (.A(_0137_),
    .X(_0167_));
 sg13g2_buf_8 _0763_ (.A(net36),
    .X(_0168_));
 sg13g2_a21oi_1 _0764_ (.A1(\desk_clock.clk_hours[4] ),
    .A2(_0149_),
    .Y(_0169_),
    .B1(\desk_clock.clk_hours[3] ));
 sg13g2_nor2b_1 _0765_ (.A(\desk_clock.clk_hours[4] ),
    .B_N(\desk_clock.clk_hours[3] ),
    .Y(_0170_));
 sg13g2_nand4_1 _0766_ (.B(_0141_),
    .C(_0159_),
    .A(\desk_clock.clk_hours[2] ),
    .Y(_0171_),
    .D(_0164_));
 sg13g2_mux2_1 _0767_ (.A0(_0169_),
    .A1(_0170_),
    .S(_0171_),
    .X(_0172_));
 sg13g2_and2_1 _0768_ (.A(net33),
    .B(_0172_),
    .X(_0029_));
 sg13g2_nand2_1 _0769_ (.Y(_0173_),
    .A(net36),
    .B(_0170_));
 sg13g2_inv_1 _0770_ (.Y(_0174_),
    .A(_0149_));
 sg13g2_inv_1 _0771_ (.Y(_0175_),
    .A(\desk_clock.clk_hours[4] ));
 sg13g2_nor3_1 _0772_ (.A(_0138_),
    .B(\desk_clock.clk_hours[3] ),
    .C(_0175_),
    .Y(_0176_));
 sg13g2_o21ai_1 _0773_ (.B1(_0176_),
    .Y(_0177_),
    .A1(_0174_),
    .A2(_0171_));
 sg13g2_o21ai_1 _0774_ (.B1(_0177_),
    .Y(_0030_),
    .A1(_0171_),
    .A2(_0173_));
 sg13g2_a21o_1 _0775_ (.A2(_0154_),
    .A1(_0152_),
    .B1(_0141_),
    .X(_0178_));
 sg13g2_and2_1 _0776_ (.A(\desk_clock.input_debounce.set_minutes_reg[1] ),
    .B(_0140_),
    .X(_0179_));
 sg13g2_or3_1 _0777_ (.A(_0179_),
    .B(_0144_),
    .C(_0145_),
    .X(_0180_));
 sg13g2_a21oi_2 _0778_ (.B1(_0158_),
    .Y(_0181_),
    .A2(_0180_),
    .A1(_0178_));
 sg13g2_inv_1 _0779_ (.Y(_0182_),
    .A(\desk_clock.clk_minutes[5] ));
 sg13g2_and2_1 _0780_ (.A(\desk_clock.clk_minutes[3] ),
    .B(\desk_clock.clk_minutes[2] ),
    .X(_0183_));
 sg13g2_nand2_1 _0781_ (.Y(_0184_),
    .A(\desk_clock.clk_minutes[4] ),
    .B(_0183_));
 sg13g2_o21ai_1 _0782_ (.B1(_0137_),
    .Y(_0185_),
    .A1(_0182_),
    .A2(_0184_));
 sg13g2_a21oi_2 _0783_ (.B1(_0185_),
    .Y(_0186_),
    .A2(_0181_),
    .A1(_0149_));
 sg13g2_xor2_1 _0784_ (.B(_0181_),
    .A(_0146_),
    .X(_0187_));
 sg13g2_and2_1 _0785_ (.A(_0186_),
    .B(_0187_),
    .X(_0031_));
 sg13g2_nand2_1 _0786_ (.Y(_0188_),
    .A(_0146_),
    .B(_0181_));
 sg13g2_xor2_1 _0787_ (.B(_0188_),
    .A(\desk_clock.clk_minutes[1] ),
    .X(_0189_));
 sg13g2_nor2b_1 _0788_ (.A(_0189_),
    .B_N(_0186_),
    .Y(_0032_));
 sg13g2_nand3_1 _0789_ (.B(_0146_),
    .C(_0181_),
    .A(\desk_clock.clk_minutes[1] ),
    .Y(_0190_));
 sg13g2_xor2_1 _0790_ (.B(_0190_),
    .A(\desk_clock.clk_minutes[2] ),
    .X(_0191_));
 sg13g2_nor2b_1 _0791_ (.A(_0191_),
    .B_N(_0186_),
    .Y(_0033_));
 sg13g2_nand4_1 _0792_ (.B(\desk_clock.clk_minutes[1] ),
    .C(_0146_),
    .A(\desk_clock.clk_minutes[2] ),
    .Y(_0192_),
    .D(_0181_));
 sg13g2_xor2_1 _0793_ (.B(_0192_),
    .A(\desk_clock.clk_minutes[3] ),
    .X(_0193_));
 sg13g2_nor2b_1 _0794_ (.A(_0193_),
    .B_N(_0186_),
    .Y(_0034_));
 sg13g2_nand4_1 _0795_ (.B(_0146_),
    .C(_0181_),
    .A(\desk_clock.clk_minutes[1] ),
    .Y(_0194_),
    .D(_0183_));
 sg13g2_xor2_1 _0796_ (.B(_0194_),
    .A(\desk_clock.clk_minutes[4] ),
    .X(_0195_));
 sg13g2_nor2b_1 _0797_ (.A(_0195_),
    .B_N(_0186_),
    .Y(_0035_));
 sg13g2_or2_1 _0798_ (.X(_0196_),
    .B(_0190_),
    .A(_0184_));
 sg13g2_a221oi_1 _0799_ (.B2(_0182_),
    .C1(_0185_),
    .B1(_0196_),
    .A1(_0149_),
    .Y(_0036_),
    .A2(_0181_));
 sg13g2_and3_1 _0800_ (.X(_0197_),
    .A(\desk_clock.clk_seconds[4] ),
    .B(\desk_clock.clk_seconds[3] ),
    .C(\desk_clock.clk_seconds[2] ));
 sg13g2_a221oi_1 _0801_ (.B2(\desk_clock.clk_seconds[5] ),
    .C1(_0138_),
    .B1(_0197_),
    .A1(_0179_),
    .Y(_0198_),
    .A2(_0158_));
 sg13g2_or2_1 _0802_ (.X(_0199_),
    .B(_0145_),
    .A(_0144_));
 sg13g2_nand2_1 _0803_ (.Y(_0200_),
    .A(_0142_),
    .B(_0199_));
 sg13g2_nand2b_1 _0804_ (.Y(_0201_),
    .B(\desk_clock.clk_seconds[0] ),
    .A_N(_0142_));
 sg13g2_o21ai_1 _0805_ (.B1(_0201_),
    .Y(_0202_),
    .A1(\desk_clock.clk_seconds[0] ),
    .A2(_0200_));
 sg13g2_and2_1 _0806_ (.A(_0198_),
    .B(_0202_),
    .X(_0037_));
 sg13g2_nand2_2 _0807_ (.Y(_0203_),
    .A(_0199_),
    .B(_0198_));
 sg13g2_nand2_1 _0808_ (.Y(_0204_),
    .A(\desk_clock.clk_seconds[0] ),
    .B(_0142_));
 sg13g2_xor2_1 _0809_ (.B(_0204_),
    .A(\desk_clock.clk_seconds[1] ),
    .X(_0205_));
 sg13g2_nor2_1 _0810_ (.A(_0203_),
    .B(_0205_),
    .Y(_0038_));
 sg13g2_and2_1 _0811_ (.A(_0142_),
    .B(_0143_),
    .X(_0206_));
 sg13g2_buf_1 _0812_ (.A(_0206_),
    .X(_0207_));
 sg13g2_xnor2_1 _0813_ (.Y(_0208_),
    .A(\desk_clock.clk_seconds[2] ),
    .B(_0207_));
 sg13g2_nor2_1 _0814_ (.A(_0203_),
    .B(_0208_),
    .Y(_0039_));
 sg13g2_nand2_1 _0815_ (.Y(_0209_),
    .A(\desk_clock.clk_seconds[2] ),
    .B(_0207_));
 sg13g2_xor2_1 _0816_ (.B(_0209_),
    .A(\desk_clock.clk_seconds[3] ),
    .X(_0210_));
 sg13g2_nor2_1 _0817_ (.A(_0203_),
    .B(_0210_),
    .Y(_0040_));
 sg13g2_nand3_1 _0818_ (.B(\desk_clock.clk_seconds[2] ),
    .C(_0207_),
    .A(\desk_clock.clk_seconds[3] ),
    .Y(_0211_));
 sg13g2_xor2_1 _0819_ (.B(_0211_),
    .A(\desk_clock.clk_seconds[4] ),
    .X(_0212_));
 sg13g2_nor2_1 _0820_ (.A(_0203_),
    .B(_0212_),
    .Y(_0041_));
 sg13g2_a21oi_1 _0821_ (.A1(_0207_),
    .A2(_0197_),
    .Y(_0213_),
    .B1(\desk_clock.clk_seconds[5] ));
 sg13g2_nor2_1 _0822_ (.A(_0203_),
    .B(_0213_),
    .Y(_0042_));
 sg13g2_buf_2 _0823_ (.A(_0000_),
    .X(_0214_));
 sg13g2_nor3_1 _0824_ (.A(_0128_),
    .B(_0214_),
    .C(_0127_),
    .Y(_0215_));
 sg13g2_inv_1 _0825_ (.Y(_0216_),
    .A(\desk_clock.display_control_inst.display_update ));
 sg13g2_nor4_1 _0826_ (.A(_0128_),
    .B(\desk_clock.display_control_inst.o_write_config ),
    .C(_0216_),
    .D(_0127_),
    .Y(_0217_));
 sg13g2_nor2_1 _0827_ (.A(_0179_),
    .B(_0158_),
    .Y(_0218_));
 sg13g2_mux2_1 _0828_ (.A0(_0155_),
    .A1(_0142_),
    .S(_0218_),
    .X(_0219_));
 sg13g2_nand2b_1 _0829_ (.Y(_0220_),
    .B(_0219_),
    .A_N(_0217_));
 sg13g2_nand3b_1 _0830_ (.B(net33),
    .C(_0220_),
    .Y(_0043_),
    .A_N(_0215_));
 sg13g2_buf_1 _0831_ (.A(\desk_clock.display_inst.disp_driver.transfer_state[1] ),
    .X(_0221_));
 sg13g2_nor3_1 _0832_ (.A(\desk_clock.display_inst.disp_driver.transfer_state[3] ),
    .B(\desk_clock.display_inst.disp_driver.transfer_state[2] ),
    .C(_0221_),
    .Y(_0222_));
 sg13g2_nand2_1 _0833_ (.Y(_0223_),
    .A(_0001_),
    .B(_0222_));
 sg13g2_buf_2 _0834_ (.A(\desk_clock.display_inst.disp_driver.transfer_state[0] ),
    .X(_0224_));
 sg13g2_or3_1 _0835_ (.A(\desk_clock.display_inst.disp_driver.transfer_state[3] ),
    .B(\desk_clock.display_inst.disp_driver.transfer_state[2] ),
    .C(_0221_),
    .X(_0225_));
 sg13g2_o21ai_1 _0836_ (.B1(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .Y(_0226_),
    .A1(_0224_),
    .A2(_0225_));
 sg13g2_o21ai_1 _0837_ (.B1(_0226_),
    .Y(_0227_),
    .A1(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .A2(_0223_));
 sg13g2_buf_1 _0838_ (.A(\desk_clock.display_inst.display_settings.transfer_state[2] ),
    .X(_0228_));
 sg13g2_buf_1 _0839_ (.A(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .X(_0229_));
 sg13g2_nor2_1 _0840_ (.A(net35),
    .B(net34),
    .Y(_0230_));
 sg13g2_inv_1 _0841_ (.Y(_0231_),
    .A(_0130_));
 sg13g2_o21ai_1 _0842_ (.B1(_0231_),
    .Y(_0232_),
    .A1(_0230_),
    .A2(_0133_));
 sg13g2_buf_1 _0843_ (.A(_0232_),
    .X(_0233_));
 sg13g2_nand2_2 _0844_ (.Y(_0234_),
    .A(_0227_),
    .B(net19));
 sg13g2_nand2_1 _0845_ (.Y(_0235_),
    .A(net36),
    .B(_0234_));
 sg13g2_nor3_2 _0846_ (.A(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .B(_0224_),
    .C(_0225_),
    .Y(_0236_));
 sg13g2_buf_1 _0847_ (.A(_0236_),
    .X(_0237_));
 sg13g2_buf_1 _0848_ (.A(_0236_),
    .X(_0238_));
 sg13g2_nor2b_1 _0849_ (.A(net17),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[11] ),
    .Y(_0239_));
 sg13g2_a21oi_1 _0850_ (.A1(\desk_clock.display_inst.disp_driver.data_reg[12] ),
    .A2(net18),
    .Y(_0240_),
    .B1(_0239_));
 sg13g2_nor2_1 _0851_ (.A(_0235_),
    .B(_0240_),
    .Y(_0048_));
 sg13g2_nor2b_1 _0852_ (.A(net17),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[12] ),
    .Y(_0241_));
 sg13g2_a21oi_1 _0853_ (.A1(\desk_clock.display_inst.disp_driver.data_reg[13] ),
    .A2(net18),
    .Y(_0242_),
    .B1(_0241_));
 sg13g2_nor2_1 _0854_ (.A(_0235_),
    .B(_0242_),
    .Y(_0049_));
 sg13g2_nor2b_1 _0855_ (.A(_0238_),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[13] ),
    .Y(_0243_));
 sg13g2_a21oi_1 _0856_ (.A1(\desk_clock.display_inst.disp_driver.data_reg[14] ),
    .A2(_0237_),
    .Y(_0244_),
    .B1(_0243_));
 sg13g2_nor2_1 _0857_ (.A(_0235_),
    .B(_0244_),
    .Y(_0050_));
 sg13g2_nor2b_1 _0858_ (.A(net17),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[14] ),
    .Y(_0245_));
 sg13g2_a21oi_1 _0859_ (.A1(\desk_clock.display_inst.disp_driver.data_reg[15] ),
    .A2(net18),
    .Y(_0246_),
    .B1(_0245_));
 sg13g2_nor2_1 _0860_ (.A(_0235_),
    .B(_0246_),
    .Y(_0051_));
 sg13g2_buf_1 _0861_ (.A(_0234_),
    .X(_0247_));
 sg13g2_buf_1 _0862_ (.A(_0167_),
    .X(_0248_));
 sg13g2_nand3_1 _0863_ (.B(_0001_),
    .C(_0226_),
    .A(net32),
    .Y(_0249_));
 sg13g2_a21oi_1 _0864_ (.A1(net12),
    .A2(net18),
    .Y(_0061_),
    .B1(_0249_));
 sg13g2_nand3_1 _0865_ (.B(_0226_),
    .C(_0234_),
    .A(net36),
    .Y(_0250_));
 sg13g2_xnor2_1 _0866_ (.Y(_0251_),
    .A(_0221_),
    .B(_0224_));
 sg13g2_nor2_1 _0867_ (.A(_0250_),
    .B(_0251_),
    .Y(_0062_));
 sg13g2_nand2_1 _0868_ (.Y(_0252_),
    .A(_0221_),
    .B(_0224_));
 sg13g2_xor2_1 _0869_ (.B(_0252_),
    .A(\desk_clock.display_inst.disp_driver.transfer_state[2] ),
    .X(_0253_));
 sg13g2_nor2_1 _0870_ (.A(_0250_),
    .B(_0253_),
    .Y(_0063_));
 sg13g2_nand3_1 _0871_ (.B(_0221_),
    .C(_0224_),
    .A(\desk_clock.display_inst.disp_driver.transfer_state[2] ),
    .Y(_0254_));
 sg13g2_xor2_1 _0872_ (.B(_0254_),
    .A(\desk_clock.display_inst.disp_driver.transfer_state[3] ),
    .X(_0255_));
 sg13g2_nor2_1 _0873_ (.A(_0250_),
    .B(_0255_),
    .Y(_0064_));
 sg13g2_nand4_1 _0874_ (.B(\desk_clock.display_inst.disp_driver.transfer_state[2] ),
    .C(_0221_),
    .A(\desk_clock.display_inst.disp_driver.transfer_state[3] ),
    .Y(_0256_),
    .D(_0224_));
 sg13g2_xor2_1 _0875_ (.B(_0256_),
    .A(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .X(_0257_));
 sg13g2_nor2_1 _0876_ (.A(_0250_),
    .B(_0257_),
    .Y(_0065_));
 sg13g2_buf_1 _0877_ (.A(_0138_),
    .X(_0258_));
 sg13g2_nor3_1 _0878_ (.A(\desk_clock.display_control_inst.o_write_config ),
    .B(_0129_),
    .C(_0134_),
    .Y(_0259_));
 sg13g2_buf_1 _0879_ (.A(_0259_),
    .X(_0260_));
 sg13g2_and2_1 _0880_ (.A(net35),
    .B(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .X(_0261_));
 sg13g2_nand2_1 _0881_ (.Y(_0262_),
    .A(_0231_),
    .B(\desk_clock.display_inst.display_settings.write_config ));
 sg13g2_nor3_2 _0882_ (.A(_0132_),
    .B(_0261_),
    .C(_0262_),
    .Y(_0263_));
 sg13g2_nor2_1 _0883_ (.A(\desk_clock.display_inst.disp_driver.i_data[4] ),
    .B(_0263_),
    .Y(_0264_));
 sg13g2_xnor2_1 _0884_ (.Y(_0265_),
    .A(net35),
    .B(_0229_));
 sg13g2_nor2_1 _0885_ (.A(_0262_),
    .B(_0265_),
    .Y(_0266_));
 sg13g2_nor4_1 _0886_ (.A(net31),
    .B(net11),
    .C(_0264_),
    .D(_0266_),
    .Y(_0074_));
 sg13g2_nor3_1 _0887_ (.A(net35),
    .B(_0130_),
    .C(net34),
    .Y(_0267_));
 sg13g2_nand3_1 _0888_ (.B(_0224_),
    .C(_0222_),
    .A(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .Y(_0268_));
 sg13g2_nand2_1 _0889_ (.Y(_0269_),
    .A(net37),
    .B(_0267_));
 sg13g2_o21ai_1 _0890_ (.B1(_0269_),
    .Y(_0270_),
    .A1(_0267_),
    .A2(_0268_));
 sg13g2_mux2_1 _0891_ (.A0(net37),
    .A1(_0004_),
    .S(_0270_),
    .X(_0271_));
 sg13g2_nor2_1 _0892_ (.A(_0135_),
    .B(_0271_),
    .Y(_0272_));
 sg13g2_nor3_1 _0893_ (.A(_0130_),
    .B(_0138_),
    .C(_0133_),
    .Y(_0273_));
 sg13g2_nand2b_1 _0894_ (.Y(_0274_),
    .B(_0273_),
    .A_N(net11));
 sg13g2_nor2_1 _0895_ (.A(_0272_),
    .B(_0274_),
    .Y(_0076_));
 sg13g2_or2_1 _0896_ (.X(_0275_),
    .B(_0134_),
    .A(_0129_));
 sg13g2_o21ai_1 _0897_ (.B1(_0273_),
    .Y(_0276_),
    .A1(_0214_),
    .A2(_0275_));
 sg13g2_a21o_1 _0898_ (.A2(_0270_),
    .A1(net37),
    .B1(net34),
    .X(_0277_));
 sg13g2_nand3_1 _0899_ (.B(net37),
    .C(_0270_),
    .A(net34),
    .Y(_0278_));
 sg13g2_a21oi_1 _0900_ (.A1(_0277_),
    .A2(_0278_),
    .Y(_0279_),
    .B1(_0135_));
 sg13g2_nor2_1 _0901_ (.A(_0276_),
    .B(_0279_),
    .Y(_0077_));
 sg13g2_xor2_1 _0902_ (.B(_0278_),
    .A(net35),
    .X(_0280_));
 sg13g2_a21oi_1 _0903_ (.A1(_0275_),
    .A2(_0280_),
    .Y(_0078_),
    .B1(_0276_));
 sg13g2_nor2b_1 _0904_ (.A(_0128_),
    .B_N(_0127_),
    .Y(_0281_));
 sg13g2_nand2_1 _0905_ (.Y(_0282_),
    .A(_0137_),
    .B(_0281_));
 sg13g2_a21o_1 _0906_ (.A2(_0281_),
    .A1(_0125_),
    .B1(_0216_),
    .X(_0283_));
 sg13g2_buf_2 _0907_ (.A(_0283_),
    .X(_0284_));
 sg13g2_buf_1 _0908_ (.A(_0284_),
    .X(_0285_));
 sg13g2_nor2_1 _0909_ (.A(_0214_),
    .B(net10),
    .Y(_0286_));
 sg13g2_inv_1 _0910_ (.Y(_0287_),
    .A(net39));
 sg13g2_or2_1 _0911_ (.X(_0288_),
    .B(_0125_),
    .A(_0128_));
 sg13g2_and3_1 _0912_ (.X(_0289_),
    .A(_0231_),
    .B(_0133_),
    .C(_0288_));
 sg13g2_buf_1 _0913_ (.A(_0289_),
    .X(_0290_));
 sg13g2_nand2_1 _0914_ (.Y(_0291_),
    .A(_0002_),
    .B(_0290_));
 sg13g2_o21ai_1 _0915_ (.B1(_0291_),
    .Y(_0292_),
    .A1(_0287_),
    .A2(_0290_));
 sg13g2_nor2b_1 _0916_ (.A(_0292_),
    .B_N(net10),
    .Y(_0293_));
 sg13g2_nor3_1 _0917_ (.A(_0282_),
    .B(_0286_),
    .C(_0293_),
    .Y(_0097_));
 sg13g2_buf_1 _0918_ (.A(net39),
    .X(_0294_));
 sg13g2_a21oi_1 _0919_ (.A1(_0294_),
    .A2(_0290_),
    .Y(_0295_),
    .B1(net40));
 sg13g2_and2_1 _0920_ (.A(\desk_clock.display_inst.state[1] ),
    .B(net39),
    .X(_0296_));
 sg13g2_buf_1 _0921_ (.A(_0296_),
    .X(_0297_));
 sg13g2_nand2_1 _0922_ (.Y(_0298_),
    .A(_0297_),
    .B(_0290_));
 sg13g2_nand2b_1 _0923_ (.Y(_0299_),
    .B(_0298_),
    .A_N(_0295_));
 sg13g2_inv_1 _0924_ (.Y(_0300_),
    .A(_0282_));
 sg13g2_o21ai_1 _0925_ (.B1(_0300_),
    .Y(_0301_),
    .A1(\desk_clock.display_control_inst.o_write_config ),
    .A2(net10));
 sg13g2_a21oi_1 _0926_ (.A1(net10),
    .A2(_0299_),
    .Y(_0098_),
    .B1(_0301_));
 sg13g2_inv_1 _0927_ (.Y(_0302_),
    .A(net38));
 sg13g2_xnor2_1 _0928_ (.Y(_0303_),
    .A(_0302_),
    .B(_0298_));
 sg13g2_a21oi_1 _0929_ (.A1(net10),
    .A2(_0303_),
    .Y(_0099_),
    .B1(_0301_));
 sg13g2_inv_1 _0930_ (.Y(_0304_),
    .A(_0122_));
 sg13g2_nor3_1 _0931_ (.A(_0302_),
    .B(_0304_),
    .C(_0002_),
    .Y(_0305_));
 sg13g2_a21oi_1 _0932_ (.A1(_0290_),
    .A2(_0305_),
    .Y(_0306_),
    .B1(_0128_));
 sg13g2_nand2_1 _0933_ (.Y(_0307_),
    .A(_0300_),
    .B(net10));
 sg13g2_nor2_1 _0934_ (.A(_0306_),
    .B(_0307_),
    .Y(_0100_));
 sg13g2_nand2b_2 _0935_ (.Y(_0308_),
    .B(\desk_clock.clk_gen_inst.i_refclk ),
    .A_N(\desk_clock.clk_gen_inst.stb_gen_refclk.sig_hold ));
 sg13g2_mux2_1 _0936_ (.A0(_0005_),
    .A1(\desk_clock.clk_gen_inst.refclk_div[0] ),
    .S(_0308_),
    .X(_0309_));
 sg13g2_and2_1 _0937_ (.A(net33),
    .B(_0309_),
    .X(_0006_));
 sg13g2_buf_1 _0938_ (.A(_0258_),
    .X(_0310_));
 sg13g2_inv_1 _0939_ (.Y(_0311_),
    .A(\desk_clock.clk_gen_inst.refclk_div[4] ));
 sg13g2_nand4_1 _0940_ (.B(\desk_clock.clk_gen_inst.refclk_div[0] ),
    .C(\desk_clock.clk_gen_inst.refclk_div[2] ),
    .A(\desk_clock.clk_gen_inst.refclk_div[1] ),
    .Y(_0312_),
    .D(\desk_clock.clk_gen_inst.refclk_div[3] ));
 sg13g2_nand4_1 _0941_ (.B(\desk_clock.clk_gen_inst.refclk_div[6] ),
    .C(\desk_clock.clk_gen_inst.refclk_div[7] ),
    .A(\desk_clock.clk_gen_inst.refclk_div[5] ),
    .Y(_0313_),
    .D(\desk_clock.clk_gen_inst.refclk_div[8] ));
 sg13g2_nor4_1 _0942_ (.A(_0311_),
    .B(_0308_),
    .C(_0312_),
    .D(_0313_),
    .Y(_0314_));
 sg13g2_and2_1 _0943_ (.A(\desk_clock.clk_gen_inst.refclk_div[9] ),
    .B(_0314_),
    .X(_0315_));
 sg13g2_buf_1 _0944_ (.A(_0315_),
    .X(_0316_));
 sg13g2_xnor2_1 _0945_ (.Y(_0317_),
    .A(\desk_clock.clk_gen_inst.refclk_div[10] ),
    .B(_0316_));
 sg13g2_nor2_1 _0946_ (.A(net24),
    .B(_0317_),
    .Y(_0007_));
 sg13g2_nand2_1 _0947_ (.Y(_0318_),
    .A(\desk_clock.clk_gen_inst.refclk_div[10] ),
    .B(_0316_));
 sg13g2_xor2_1 _0948_ (.B(_0318_),
    .A(\desk_clock.clk_gen_inst.refclk_div[11] ),
    .X(_0319_));
 sg13g2_nor2_1 _0949_ (.A(net24),
    .B(_0319_),
    .Y(_0008_));
 sg13g2_nand3_1 _0950_ (.B(\desk_clock.clk_gen_inst.refclk_div[10] ),
    .C(_0316_),
    .A(\desk_clock.clk_gen_inst.refclk_div[11] ),
    .Y(_0320_));
 sg13g2_xor2_1 _0951_ (.B(_0320_),
    .A(\desk_clock.clk_gen_inst.refclk_div[12] ),
    .X(_0321_));
 sg13g2_nor2_1 _0952_ (.A(net24),
    .B(_0321_),
    .Y(_0009_));
 sg13g2_inv_1 _0953_ (.Y(_0322_),
    .A(\desk_clock.clk_gen_inst.refclk_div[13] ));
 sg13g2_nand4_1 _0954_ (.B(\desk_clock.clk_gen_inst.refclk_div[10] ),
    .C(\desk_clock.clk_gen_inst.refclk_div[12] ),
    .A(\desk_clock.clk_gen_inst.refclk_div[11] ),
    .Y(_0323_),
    .D(_0316_));
 sg13g2_xnor2_1 _0955_ (.Y(_0324_),
    .A(_0322_),
    .B(_0323_));
 sg13g2_nor2_1 _0956_ (.A(net24),
    .B(_0324_),
    .Y(_0010_));
 sg13g2_nor2_1 _0957_ (.A(_0322_),
    .B(_0323_),
    .Y(_0325_));
 sg13g2_xor2_1 _0958_ (.B(_0325_),
    .A(\desk_clock.clk_gen_inst.refclk_div[14] ),
    .X(_0326_));
 sg13g2_and2_1 _0959_ (.A(net33),
    .B(_0326_),
    .X(_0011_));
 sg13g2_inv_1 _0960_ (.Y(_0327_),
    .A(\desk_clock.clk_gen_inst.refclk_div[1] ));
 sg13g2_nand3b_1 _0961_ (.B(\desk_clock.clk_gen_inst.i_refclk ),
    .C(\desk_clock.clk_gen_inst.refclk_div[0] ),
    .Y(_0328_),
    .A_N(\desk_clock.clk_gen_inst.stb_gen_refclk.sig_hold ));
 sg13g2_xnor2_1 _0962_ (.Y(_0329_),
    .A(_0327_),
    .B(_0328_));
 sg13g2_nor2_1 _0963_ (.A(net24),
    .B(_0329_),
    .Y(_0012_));
 sg13g2_nor2_1 _0964_ (.A(_0327_),
    .B(_0328_),
    .Y(_0330_));
 sg13g2_xnor2_1 _0965_ (.Y(_0331_),
    .A(\desk_clock.clk_gen_inst.refclk_div[2] ),
    .B(_0330_));
 sg13g2_nor2_1 _0966_ (.A(_0310_),
    .B(_0331_),
    .Y(_0013_));
 sg13g2_nand2_1 _0967_ (.Y(_0332_),
    .A(\desk_clock.clk_gen_inst.refclk_div[2] ),
    .B(_0330_));
 sg13g2_xor2_1 _0968_ (.B(_0332_),
    .A(\desk_clock.clk_gen_inst.refclk_div[3] ),
    .X(_0333_));
 sg13g2_nor2_1 _0969_ (.A(_0310_),
    .B(_0333_),
    .Y(_0014_));
 sg13g2_nor2_1 _0970_ (.A(_0308_),
    .B(_0312_),
    .Y(_0334_));
 sg13g2_xnor2_1 _0971_ (.Y(_0335_),
    .A(\desk_clock.clk_gen_inst.refclk_div[4] ),
    .B(_0334_));
 sg13g2_nor2_1 _0972_ (.A(net24),
    .B(_0335_),
    .Y(_0015_));
 sg13g2_nor3_2 _0973_ (.A(_0311_),
    .B(_0308_),
    .C(_0312_),
    .Y(_0336_));
 sg13g2_xnor2_1 _0974_ (.Y(_0337_),
    .A(\desk_clock.clk_gen_inst.refclk_div[5] ),
    .B(_0336_));
 sg13g2_nor2_1 _0975_ (.A(net24),
    .B(_0337_),
    .Y(_0016_));
 sg13g2_nand2_1 _0976_ (.Y(_0338_),
    .A(\desk_clock.clk_gen_inst.refclk_div[5] ),
    .B(_0336_));
 sg13g2_xor2_1 _0977_ (.B(_0338_),
    .A(\desk_clock.clk_gen_inst.refclk_div[6] ),
    .X(_0339_));
 sg13g2_nor2_1 _0978_ (.A(net24),
    .B(_0339_),
    .Y(_0017_));
 sg13g2_buf_1 _0979_ (.A(_0138_),
    .X(_0340_));
 sg13g2_nand3_1 _0980_ (.B(\desk_clock.clk_gen_inst.refclk_div[6] ),
    .C(_0336_),
    .A(\desk_clock.clk_gen_inst.refclk_div[5] ),
    .Y(_0341_));
 sg13g2_xor2_1 _0981_ (.B(_0341_),
    .A(\desk_clock.clk_gen_inst.refclk_div[7] ),
    .X(_0342_));
 sg13g2_nor2_1 _0982_ (.A(net29),
    .B(_0342_),
    .Y(_0018_));
 sg13g2_nand4_1 _0983_ (.B(\desk_clock.clk_gen_inst.refclk_div[6] ),
    .C(\desk_clock.clk_gen_inst.refclk_div[7] ),
    .A(\desk_clock.clk_gen_inst.refclk_div[5] ),
    .Y(_0343_),
    .D(_0336_));
 sg13g2_xor2_1 _0984_ (.B(_0343_),
    .A(\desk_clock.clk_gen_inst.refclk_div[8] ),
    .X(_0344_));
 sg13g2_nor2_1 _0985_ (.A(net29),
    .B(_0344_),
    .Y(_0019_));
 sg13g2_xnor2_1 _0986_ (.Y(_0345_),
    .A(\desk_clock.clk_gen_inst.refclk_div[9] ),
    .B(_0314_));
 sg13g2_nor2_1 _0987_ (.A(_0340_),
    .B(_0345_),
    .Y(_0020_));
 sg13g2_and2_1 _0988_ (.A(net33),
    .B(\desk_clock.clk_gen_inst.refclk_div[14] ),
    .X(_0021_));
 sg13g2_and2_1 _0989_ (.A(net33),
    .B(\desk_clock.clk_gen_inst.refclk_div[3] ),
    .X(_0022_));
 sg13g2_and2_1 _0990_ (.A(net33),
    .B(\desk_clock.clk_gen_inst.refclk_div[11] ),
    .X(_0023_));
 sg13g2_and2_1 _0991_ (.A(_0168_),
    .B(\desk_clock.clk_gen_inst.i_refclk ),
    .X(_0024_));
 sg13g2_nor2_1 _0992_ (.A(_0340_),
    .B(_0322_),
    .Y(_0025_));
 sg13g2_inv_1 _0993_ (.Y(_0346_),
    .A(\desk_clock.display_control_inst.o_write_config ));
 sg13g2_o21ai_1 _0994_ (.B1(net33),
    .Y(_0044_),
    .A1(_0346_),
    .A2(_0215_));
 sg13g2_buf_1 _0995_ (.A(_0227_),
    .X(\desk_clock.display_inst.disp_driver.o_serial_load ));
 sg13g2_and2_1 _0996_ (.A(net15),
    .B(net19),
    .X(_0347_));
 sg13g2_nand2_1 _0997_ (.Y(_0348_),
    .A(\desk_clock.display_inst.disp_driver.i_data[0] ),
    .B(_0347_));
 sg13g2_nand3_1 _0998_ (.B(_0234_),
    .C(net18),
    .A(\desk_clock.display_inst.disp_driver.data_reg[0] ),
    .Y(_0349_));
 sg13g2_a21oi_1 _0999_ (.A1(_0348_),
    .A2(_0349_),
    .Y(_0045_),
    .B1(net29));
 sg13g2_buf_1 _1000_ (.A(_0138_),
    .X(_0350_));
 sg13g2_nor2_1 _1001_ (.A(\desk_clock.display_inst.disp_driver.i_addr[2] ),
    .B(_0247_),
    .Y(_0351_));
 sg13g2_buf_1 _1002_ (.A(_0236_),
    .X(_0352_));
 sg13g2_nor2b_1 _1003_ (.A(net16),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[9] ),
    .Y(_0353_));
 sg13g2_a221oi_1 _1004_ (.B2(\desk_clock.display_inst.disp_driver.data_reg[10] ),
    .C1(_0353_),
    .B1(net18),
    .A1(net15),
    .Y(_0354_),
    .A2(net19));
 sg13g2_nor3_1 _1005_ (.A(net28),
    .B(_0351_),
    .C(_0354_),
    .Y(_0046_));
 sg13g2_nor2_1 _1006_ (.A(\desk_clock.display_inst.disp_driver.i_addr[3] ),
    .B(_0247_),
    .Y(_0355_));
 sg13g2_nor2b_1 _1007_ (.A(net16),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[10] ),
    .Y(_0356_));
 sg13g2_a221oi_1 _1008_ (.B2(\desk_clock.display_inst.disp_driver.data_reg[11] ),
    .C1(_0356_),
    .B1(net17),
    .A1(net15),
    .Y(_0357_),
    .A2(net19));
 sg13g2_nor3_1 _1009_ (.A(net28),
    .B(_0355_),
    .C(_0357_),
    .Y(_0047_));
 sg13g2_nand2_1 _1010_ (.Y(_0358_),
    .A(\desk_clock.display_inst.disp_driver.i_data[1] ),
    .B(_0347_));
 sg13g2_mux2_1 _1011_ (.A0(\desk_clock.display_inst.disp_driver.data_reg[0] ),
    .A1(\desk_clock.display_inst.disp_driver.data_reg[1] ),
    .S(_0236_),
    .X(_0359_));
 sg13g2_nand2_1 _1012_ (.Y(_0360_),
    .A(net12),
    .B(_0359_));
 sg13g2_a21oi_1 _1013_ (.A1(_0358_),
    .A2(_0360_),
    .Y(_0052_),
    .B1(net29));
 sg13g2_nor2_1 _1014_ (.A(\desk_clock.display_inst.disp_driver.i_data[2] ),
    .B(net12),
    .Y(_0361_));
 sg13g2_nor2b_1 _1015_ (.A(net16),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[1] ),
    .Y(_0362_));
 sg13g2_a221oi_1 _1016_ (.B2(\desk_clock.display_inst.disp_driver.data_reg[2] ),
    .C1(_0362_),
    .B1(net17),
    .A1(net15),
    .Y(_0363_),
    .A2(net19));
 sg13g2_nor3_1 _1017_ (.A(net31),
    .B(_0361_),
    .C(_0363_),
    .Y(_0053_));
 sg13g2_nor2_1 _1018_ (.A(\desk_clock.display_inst.disp_driver.i_data[3] ),
    .B(net12),
    .Y(_0364_));
 sg13g2_nor2b_1 _1019_ (.A(net16),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[2] ),
    .Y(_0365_));
 sg13g2_a221oi_1 _1020_ (.B2(\desk_clock.display_inst.disp_driver.data_reg[3] ),
    .C1(_0365_),
    .B1(net17),
    .A1(net15),
    .Y(_0366_),
    .A2(net19));
 sg13g2_nor3_1 _1021_ (.A(net31),
    .B(_0364_),
    .C(_0366_),
    .Y(_0054_));
 sg13g2_nand2b_1 _1022_ (.Y(_0367_),
    .B(net16),
    .A_N(\desk_clock.display_inst.disp_driver.data_reg[4] ));
 sg13g2_o21ai_1 _1023_ (.B1(_0367_),
    .Y(_0368_),
    .A1(\desk_clock.display_inst.disp_driver.data_reg[3] ),
    .A2(net18));
 sg13g2_o21ai_1 _1024_ (.B1(net36),
    .Y(_0369_),
    .A1(\desk_clock.display_inst.disp_driver.i_data[4] ),
    .A2(_0234_));
 sg13g2_a21oi_1 _1025_ (.A1(net12),
    .A2(_0368_),
    .Y(_0055_),
    .B1(_0369_));
 sg13g2_nand2b_1 _1026_ (.Y(_0370_),
    .B(net16),
    .A_N(\desk_clock.display_inst.disp_driver.data_reg[5] ));
 sg13g2_o21ai_1 _1027_ (.B1(_0370_),
    .Y(_0371_),
    .A1(\desk_clock.display_inst.disp_driver.data_reg[4] ),
    .A2(net18));
 sg13g2_a21oi_1 _1028_ (.A1(net12),
    .A2(_0371_),
    .Y(_0056_),
    .B1(_0369_));
 sg13g2_nand2b_1 _1029_ (.Y(_0372_),
    .B(net16),
    .A_N(\desk_clock.display_inst.disp_driver.data_reg[6] ));
 sg13g2_o21ai_1 _1030_ (.B1(_0372_),
    .Y(_0373_),
    .A1(\desk_clock.display_inst.disp_driver.data_reg[5] ),
    .A2(_0237_));
 sg13g2_a21oi_1 _1031_ (.A1(net12),
    .A2(_0373_),
    .Y(_0057_),
    .B1(_0369_));
 sg13g2_nor2_1 _1032_ (.A(\desk_clock.display_inst.disp_driver.i_data[7] ),
    .B(net12),
    .Y(_0374_));
 sg13g2_nor2b_1 _1033_ (.A(net16),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[6] ),
    .Y(_0375_));
 sg13g2_a221oi_1 _1034_ (.B2(\desk_clock.display_inst.disp_driver.data_reg[7] ),
    .C1(_0375_),
    .B1(_0238_),
    .A1(net15),
    .Y(_0376_),
    .A2(net19));
 sg13g2_nor3_1 _1035_ (.A(net31),
    .B(_0374_),
    .C(_0376_),
    .Y(_0058_));
 sg13g2_nor2_1 _1036_ (.A(\desk_clock.display_inst.disp_driver.i_addr[0] ),
    .B(_0234_),
    .Y(_0377_));
 sg13g2_nor2b_1 _1037_ (.A(_0352_),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[7] ),
    .Y(_0378_));
 sg13g2_a221oi_1 _1038_ (.B2(\desk_clock.display_inst.disp_driver.data_reg[8] ),
    .C1(_0378_),
    .B1(net17),
    .A1(net15),
    .Y(_0379_),
    .A2(net19));
 sg13g2_nor3_1 _1039_ (.A(net31),
    .B(_0377_),
    .C(_0379_),
    .Y(_0059_));
 sg13g2_nor2_1 _1040_ (.A(\desk_clock.display_inst.disp_driver.i_addr[1] ),
    .B(_0234_),
    .Y(_0380_));
 sg13g2_nor2b_1 _1041_ (.A(_0352_),
    .B_N(\desk_clock.display_inst.disp_driver.data_reg[8] ),
    .Y(_0381_));
 sg13g2_a221oi_1 _1042_ (.B2(\desk_clock.display_inst.disp_driver.data_reg[9] ),
    .C1(_0381_),
    .B1(net17),
    .A1(net15),
    .Y(_0382_),
    .A2(_0233_));
 sg13g2_nor3_1 _1043_ (.A(net31),
    .B(_0380_),
    .C(_0382_),
    .Y(_0060_));
 sg13g2_a21oi_2 _1044_ (.B1(_0263_),
    .Y(_0383_),
    .A2(_0135_),
    .A1(_0214_));
 sg13g2_a21o_1 _1045_ (.A2(_0135_),
    .A1(_0214_),
    .B1(_0263_),
    .X(_0384_));
 sg13g2_buf_2 _1046_ (.A(_0384_),
    .X(_0385_));
 sg13g2_nand2_1 _1047_ (.Y(_0386_),
    .A(_0287_),
    .B(net11));
 sg13g2_or3_1 _1048_ (.A(_0130_),
    .B(_0131_),
    .C(_0265_),
    .X(_0387_));
 sg13g2_and3_1 _1049_ (.X(_0388_),
    .A(_0385_),
    .B(_0386_),
    .C(_0387_));
 sg13g2_a21oi_1 _1050_ (.A1(\desk_clock.display_inst.disp_driver.i_addr[0] ),
    .A2(_0383_),
    .Y(_0389_),
    .B1(_0388_));
 sg13g2_nor2_1 _1051_ (.A(net29),
    .B(_0389_),
    .Y(_0066_));
 sg13g2_nor2_1 _1052_ (.A(\desk_clock.display_inst.disp_driver.i_addr[1] ),
    .B(_0385_),
    .Y(_0390_));
 sg13g2_nand2_1 _1053_ (.Y(_0391_),
    .A(net35),
    .B(net37));
 sg13g2_nand2b_1 _1054_ (.Y(_0392_),
    .B(net34),
    .A_N(net35));
 sg13g2_o21ai_1 _1055_ (.B1(_0392_),
    .Y(_0393_),
    .A1(net34),
    .A2(_0391_));
 sg13g2_a221oi_1 _1056_ (.B2(_0231_),
    .C1(_0383_),
    .B1(_0393_),
    .A1(net40),
    .Y(_0394_),
    .A2(net11));
 sg13g2_nor3_1 _1057_ (.A(net31),
    .B(_0390_),
    .C(_0394_),
    .Y(_0067_));
 sg13g2_nor2_1 _1058_ (.A(\desk_clock.display_inst.disp_driver.i_addr[2] ),
    .B(_0385_),
    .Y(_0395_));
 sg13g2_buf_1 _1059_ (.A(_0126_),
    .X(_0396_));
 sg13g2_nor2_1 _1060_ (.A(_0130_),
    .B(net34),
    .Y(_0397_));
 sg13g2_a221oi_1 _1061_ (.B2(net35),
    .C1(_0383_),
    .B1(_0397_),
    .A1(net27),
    .Y(_0398_),
    .A2(_0260_));
 sg13g2_nor3_1 _1062_ (.A(net31),
    .B(_0395_),
    .C(_0398_),
    .Y(_0068_));
 sg13g2_a21oi_1 _1063_ (.A1(_0125_),
    .A2(_0260_),
    .Y(_0399_),
    .B1(_0383_));
 sg13g2_a21oi_1 _1064_ (.A1(\desk_clock.display_inst.disp_driver.i_addr[3] ),
    .A2(_0383_),
    .Y(_0400_),
    .B1(_0399_));
 sg13g2_nor2_1 _1065_ (.A(net29),
    .B(_0400_),
    .Y(_0069_));
 sg13g2_nor2_1 _1066_ (.A(net27),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[3] ),
    .Y(_0401_));
 sg13g2_nor2b_1 _1067_ (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[3] ),
    .B_N(net27),
    .Y(_0402_));
 sg13g2_nor2_2 _1068_ (.A(net40),
    .B(net39),
    .Y(_0403_));
 sg13g2_a22oi_1 _1069_ (.Y(_0404_),
    .B1(_0402_),
    .B2(_0403_),
    .A2(_0401_),
    .A1(_0297_));
 sg13g2_xor2_1 _1070_ (.B(net39),
    .A(\desk_clock.display_inst.state[1] ),
    .X(_0405_));
 sg13g2_nand2_1 _1071_ (.Y(_0406_),
    .A(_0396_),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[3] ));
 sg13g2_nand2b_1 _1072_ (.Y(_0407_),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[3] ),
    .A_N(_0396_));
 sg13g2_nand3_1 _1073_ (.B(_0406_),
    .C(_0407_),
    .A(_0405_),
    .Y(_0408_));
 sg13g2_nand2_1 _1074_ (.Y(_0409_),
    .A(_0404_),
    .B(_0408_));
 sg13g2_nand2_1 _1075_ (.Y(_0410_),
    .A(_0123_),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[5] ));
 sg13g2_o21ai_1 _1076_ (.B1(net40),
    .Y(_0411_),
    .A1(_0123_),
    .A2(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[5] ));
 sg13g2_a21o_1 _1077_ (.A2(_0411_),
    .A1(_0410_),
    .B1(_0302_),
    .X(_0412_));
 sg13g2_buf_1 _1078_ (.A(_0412_),
    .X(_0413_));
 sg13g2_nand2b_1 _1079_ (.Y(_0414_),
    .B(net27),
    .A_N(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[5] ));
 sg13g2_and3_1 _1080_ (.X(_0415_),
    .A(net40),
    .B(net39),
    .C(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[5] ));
 sg13g2_a21oi_2 _1081_ (.B1(_0415_),
    .Y(_0416_),
    .A2(_0414_),
    .A1(_0403_));
 sg13g2_and2_1 _1082_ (.A(_0413_),
    .B(_0416_),
    .X(_0417_));
 sg13g2_nor2_1 _1083_ (.A(net38),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[1] ),
    .Y(_0418_));
 sg13g2_nor2b_1 _1084_ (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[1] ),
    .B_N(\desk_clock.display_inst.state[2] ),
    .Y(_0419_));
 sg13g2_a22oi_1 _1085_ (.Y(_0420_),
    .B1(_0419_),
    .B2(_0403_),
    .A2(_0418_),
    .A1(_0297_));
 sg13g2_nand2_1 _1086_ (.Y(_0421_),
    .A(\desk_clock.display_inst.state[2] ),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[1] ));
 sg13g2_nand2b_1 _1087_ (.Y(_0422_),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[1] ),
    .A_N(\desk_clock.display_inst.state[2] ));
 sg13g2_nand3_1 _1088_ (.B(_0421_),
    .C(_0422_),
    .A(_0405_),
    .Y(_0423_));
 sg13g2_buf_1 _1089_ (.A(_0423_),
    .X(_0424_));
 sg13g2_a22oi_1 _1090_ (.Y(_0425_),
    .B1(_0420_),
    .B2(_0424_),
    .A2(_0416_),
    .A1(_0413_));
 sg13g2_inv_1 _1091_ (.Y(_0426_),
    .A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[4] ));
 sg13g2_mux2_1 _1092_ (.A0(_0403_),
    .A1(_0297_),
    .S(_0302_),
    .X(_0427_));
 sg13g2_nor2_1 _1093_ (.A(net38),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[2] ),
    .Y(_0428_));
 sg13g2_nor2b_1 _1094_ (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[2] ),
    .B_N(net38),
    .Y(_0429_));
 sg13g2_a22oi_1 _1095_ (.Y(_0430_),
    .B1(_0429_),
    .B2(_0403_),
    .A2(_0428_),
    .A1(_0297_));
 sg13g2_nand2_1 _1096_ (.Y(_0431_),
    .A(net38),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[2] ));
 sg13g2_nand2b_1 _1097_ (.Y(_0432_),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[2] ),
    .A_N(net38));
 sg13g2_nand3_1 _1098_ (.B(_0431_),
    .C(_0432_),
    .A(_0405_),
    .Y(_0433_));
 sg13g2_buf_1 _1099_ (.A(_0433_),
    .X(_0434_));
 sg13g2_nand2_1 _1100_ (.Y(_0435_),
    .A(net38),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[4] ));
 sg13g2_nand2b_1 _1101_ (.Y(_0436_),
    .B(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[4] ),
    .A_N(net38));
 sg13g2_and3_1 _1102_ (.X(_0437_),
    .A(_0405_),
    .B(_0435_),
    .C(_0436_));
 sg13g2_buf_1 _1103_ (.A(_0437_),
    .X(_0438_));
 sg13g2_a221oi_1 _1104_ (.B2(_0434_),
    .C1(_0438_),
    .B1(_0430_),
    .A1(_0426_),
    .Y(_0439_),
    .A2(_0427_));
 sg13g2_buf_1 _1105_ (.A(_0439_),
    .X(_0440_));
 sg13g2_mux2_1 _1106_ (.A0(_0417_),
    .A1(_0425_),
    .S(_0440_),
    .X(_0441_));
 sg13g2_nand3_1 _1107_ (.B(net14),
    .C(_0441_),
    .A(net30),
    .Y(_0442_));
 sg13g2_mux2_1 _1108_ (.A0(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[0] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[0] ),
    .S(net40),
    .X(_0443_));
 sg13g2_nor2_1 _1109_ (.A(_0302_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_nor3_1 _1110_ (.A(net27),
    .B(_0304_),
    .C(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[0] ),
    .Y(_0445_));
 sg13g2_o21ai_1 _1111_ (.B1(_0287_),
    .Y(_0446_),
    .A1(_0444_),
    .A2(_0445_));
 sg13g2_and2_1 _1112_ (.A(_0430_),
    .B(_0434_),
    .X(_0447_));
 sg13g2_and2_1 _1113_ (.A(_0420_),
    .B(_0424_),
    .X(_0448_));
 sg13g2_buf_1 _1114_ (.A(_0448_),
    .X(_0449_));
 sg13g2_buf_1 _1115_ (.A(_0449_),
    .X(_0450_));
 sg13g2_nand3_1 _1116_ (.B(_0417_),
    .C(net8),
    .A(_0447_),
    .Y(_0451_));
 sg13g2_a21oi_1 _1117_ (.A1(_0426_),
    .A2(_0427_),
    .Y(_0452_),
    .B1(_0438_));
 sg13g2_nand2_2 _1118_ (.Y(_0453_),
    .A(_0413_),
    .B(_0416_));
 sg13g2_a22oi_1 _1119_ (.Y(_0454_),
    .B1(_0420_),
    .B2(_0424_),
    .A2(_0434_),
    .A1(_0430_));
 sg13g2_or3_1 _1120_ (.A(_0452_),
    .B(_0453_),
    .C(_0454_),
    .X(_0455_));
 sg13g2_nand3_1 _1121_ (.B(_0404_),
    .C(_0408_),
    .A(net30),
    .Y(_0456_));
 sg13g2_a21oi_1 _1122_ (.A1(_0440_),
    .A2(_0453_),
    .Y(_0457_),
    .B1(_0456_));
 sg13g2_nand3_1 _1123_ (.B(_0455_),
    .C(_0457_),
    .A(_0451_),
    .Y(_0458_));
 sg13g2_nand4_1 _1124_ (.B(_0442_),
    .C(_0446_),
    .A(net11),
    .Y(_0459_),
    .D(_0458_));
 sg13g2_nor2b_1 _1125_ (.A(_0397_),
    .B_N(_0129_),
    .Y(_0460_));
 sg13g2_nor2_1 _1126_ (.A(_0231_),
    .B(_0129_),
    .Y(_0461_));
 sg13g2_nor4_1 _1127_ (.A(_0228_),
    .B(_0130_),
    .C(_0229_),
    .D(_0131_),
    .Y(_0462_));
 sg13g2_nor3_1 _1128_ (.A(_0121_),
    .B(_0461_),
    .C(_0462_),
    .Y(_0463_));
 sg13g2_o21ai_1 _1129_ (.B1(_0463_),
    .Y(_0464_),
    .A1(_0391_),
    .A2(_0460_));
 sg13g2_and2_1 _1130_ (.A(_0385_),
    .B(_0464_),
    .X(_0465_));
 sg13g2_o21ai_1 _1131_ (.B1(net32),
    .Y(_0466_),
    .A1(\desk_clock.display_inst.disp_driver.i_data[0] ),
    .A2(_0385_));
 sg13g2_a21oi_1 _1132_ (.A1(_0459_),
    .A2(_0465_),
    .Y(_0070_),
    .B1(_0466_));
 sg13g2_nand2_2 _1133_ (.Y(_0467_),
    .A(_0430_),
    .B(_0434_));
 sg13g2_a21oi_1 _1134_ (.A1(net14),
    .A2(_0467_),
    .Y(_0468_),
    .B1(_0453_));
 sg13g2_o21ai_1 _1135_ (.B1(net13),
    .Y(_0469_),
    .A1(net14),
    .A2(_0467_));
 sg13g2_or2_1 _1136_ (.X(_0470_),
    .B(_0469_),
    .A(_0468_));
 sg13g2_a22oi_1 _1137_ (.Y(_0471_),
    .B1(_0413_),
    .B2(_0416_),
    .A2(_0408_),
    .A1(_0404_));
 sg13g2_buf_1 _1138_ (.A(_0471_),
    .X(_0472_));
 sg13g2_nor2_1 _1139_ (.A(net13),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_nor2_1 _1140_ (.A(_0287_),
    .B(_0473_),
    .Y(_0474_));
 sg13g2_nor3_1 _1141_ (.A(net30),
    .B(_0467_),
    .C(net8),
    .Y(_0475_));
 sg13g2_a21o_1 _1142_ (.A2(_0427_),
    .A1(_0426_),
    .B1(_0438_),
    .X(_0476_));
 sg13g2_buf_1 _1143_ (.A(_0476_),
    .X(_0477_));
 sg13g2_and4_1 _1144_ (.A(_0404_),
    .B(_0408_),
    .C(_0413_),
    .D(_0416_),
    .X(_0478_));
 sg13g2_a21o_1 _1145_ (.A2(_0478_),
    .A1(_0477_),
    .B1(_0472_),
    .X(_0479_));
 sg13g2_xnor2_1 _1146_ (.Y(_0480_),
    .A(_0440_),
    .B(net8));
 sg13g2_nor4_1 _1147_ (.A(net30),
    .B(_0472_),
    .C(_0478_),
    .D(_0480_),
    .Y(_0481_));
 sg13g2_a221oi_1 _1148_ (.B2(_0479_),
    .C1(_0481_),
    .B1(_0475_),
    .A1(_0470_),
    .Y(_0482_),
    .A2(_0474_));
 sg13g2_nand2b_1 _1149_ (.Y(_0483_),
    .B(net34),
    .A_N(net37));
 sg13g2_a21o_1 _1150_ (.A2(_0135_),
    .A1(_0214_),
    .B1(_0266_),
    .X(_0484_));
 sg13g2_o21ai_1 _1151_ (.B1(_0484_),
    .Y(_0485_),
    .A1(_0135_),
    .A2(_0483_));
 sg13g2_nand2_1 _1152_ (.Y(_0486_),
    .A(_0477_),
    .B(_0472_));
 sg13g2_nand3_1 _1153_ (.B(net8),
    .C(_0478_),
    .A(_0440_),
    .Y(_0487_));
 sg13g2_o21ai_1 _1154_ (.B1(_0487_),
    .Y(_0488_),
    .A1(net8),
    .A2(_0486_));
 sg13g2_nor2_1 _1155_ (.A(_0485_),
    .B(_0488_),
    .Y(_0489_));
 sg13g2_inv_1 _1156_ (.Y(_0490_),
    .A(\desk_clock.display_inst.disp_driver.i_data[1] ));
 sg13g2_a21oi_1 _1157_ (.A1(_0490_),
    .A2(_0383_),
    .Y(_0491_),
    .B1(_0138_));
 sg13g2_o21ai_1 _1158_ (.B1(_0491_),
    .Y(_0492_),
    .A1(net11),
    .A2(_0485_));
 sg13g2_a21oi_1 _1159_ (.A1(_0482_),
    .A2(_0489_),
    .Y(_0071_),
    .B1(_0492_));
 sg13g2_a21oi_1 _1160_ (.A1(_0409_),
    .A2(_0477_),
    .Y(_0493_),
    .B1(_0417_));
 sg13g2_nand2b_1 _1161_ (.Y(_0494_),
    .B(net30),
    .A_N(_0493_));
 sg13g2_a221oi_1 _1162_ (.B2(_0449_),
    .C1(_0477_),
    .B1(_0453_),
    .A1(_0430_),
    .Y(_0495_),
    .A2(_0434_));
 sg13g2_nand2_1 _1163_ (.Y(_0496_),
    .A(_0410_),
    .B(_0411_));
 sg13g2_a21o_1 _1164_ (.A2(_0414_),
    .A1(_0403_),
    .B1(_0415_),
    .X(_0497_));
 sg13g2_a221oi_1 _1165_ (.B2(_0424_),
    .C1(_0497_),
    .B1(_0420_),
    .A1(net27),
    .Y(_0498_),
    .A2(_0496_));
 sg13g2_nor3_1 _1166_ (.A(_0467_),
    .B(net13),
    .C(_0498_),
    .Y(_0499_));
 sg13g2_or4_1 _1167_ (.A(net30),
    .B(net14),
    .C(_0495_),
    .D(_0499_),
    .X(_0500_));
 sg13g2_and3_1 _1168_ (.X(_0501_),
    .A(_0447_),
    .B(_0450_),
    .C(_0472_));
 sg13g2_a21oi_1 _1169_ (.A1(_0453_),
    .A2(net8),
    .Y(_0502_),
    .B1(_0447_));
 sg13g2_nor2_1 _1170_ (.A(net30),
    .B(net13),
    .Y(_0503_));
 sg13g2_o21ai_1 _1171_ (.B1(_0503_),
    .Y(_0504_),
    .A1(_0501_),
    .A2(_0502_));
 sg13g2_nand3_1 _1172_ (.B(_0500_),
    .C(_0504_),
    .A(_0494_),
    .Y(_0505_));
 sg13g2_and2_1 _1173_ (.A(_0467_),
    .B(_0498_),
    .X(_0506_));
 sg13g2_and3_1 _1174_ (.X(_0507_),
    .A(_0447_),
    .B(_0453_),
    .C(_0449_));
 sg13g2_nand2_1 _1175_ (.Y(_0508_),
    .A(net14),
    .B(net13));
 sg13g2_or4_1 _1176_ (.A(net30),
    .B(_0506_),
    .C(_0507_),
    .D(_0508_),
    .X(_0509_));
 sg13g2_nand4_1 _1177_ (.B(net11),
    .C(_0385_),
    .A(net36),
    .Y(_0510_),
    .D(_0509_));
 sg13g2_nand2b_1 _1178_ (.Y(_0511_),
    .B(net37),
    .A_N(_0228_));
 sg13g2_a21oi_1 _1179_ (.A1(_0483_),
    .A2(_0511_),
    .Y(_0512_),
    .B1(_0130_));
 sg13g2_o21ai_1 _1180_ (.B1(\desk_clock.display_inst.display_settings.write_config ),
    .Y(_0513_),
    .A1(_0460_),
    .A2(_0512_));
 sg13g2_nor2_1 _1181_ (.A(_0383_),
    .B(_0513_),
    .Y(_0514_));
 sg13g2_and2_1 _1182_ (.A(net36),
    .B(\desk_clock.display_inst.disp_driver.i_data[2] ),
    .X(_0515_));
 sg13g2_a22oi_1 _1183_ (.Y(_0516_),
    .B1(_0515_),
    .B2(_0383_),
    .A2(_0514_),
    .A1(net36));
 sg13g2_o21ai_1 _1184_ (.B1(_0516_),
    .Y(_0072_),
    .A1(_0505_),
    .A2(_0510_));
 sg13g2_or3_1 _1185_ (.A(net14),
    .B(net13),
    .C(_0449_),
    .X(_0517_));
 sg13g2_nand3_1 _1186_ (.B(net13),
    .C(net8),
    .A(net14),
    .Y(_0518_));
 sg13g2_a21oi_1 _1187_ (.A1(_0517_),
    .A2(_0518_),
    .Y(_0519_),
    .B1(_0453_));
 sg13g2_xnor2_1 _1188_ (.Y(_0520_),
    .A(net14),
    .B(net8));
 sg13g2_nand2_1 _1189_ (.Y(_0521_),
    .A(net13),
    .B(_0453_));
 sg13g2_o21ai_1 _1190_ (.B1(_0467_),
    .Y(_0522_),
    .A1(_0520_),
    .A2(_0521_));
 sg13g2_nand3_1 _1191_ (.B(_0450_),
    .C(_0472_),
    .A(_0477_),
    .Y(_0523_));
 sg13g2_a221oi_1 _1192_ (.B2(_0424_),
    .C1(_0438_),
    .B1(_0420_),
    .A1(_0426_),
    .Y(_0524_),
    .A2(_0427_));
 sg13g2_a21oi_1 _1193_ (.A1(_0524_),
    .A2(_0478_),
    .Y(_0525_),
    .B1(_0467_));
 sg13g2_a21oi_1 _1194_ (.A1(_0523_),
    .A2(_0525_),
    .Y(_0526_),
    .B1(_0386_));
 sg13g2_o21ai_1 _1195_ (.B1(_0526_),
    .Y(_0527_),
    .A1(_0519_),
    .A2(_0522_));
 sg13g2_o21ai_1 _1196_ (.B1(net32),
    .Y(_0528_),
    .A1(\desk_clock.display_inst.disp_driver.i_data[3] ),
    .A2(_0385_));
 sg13g2_a21oi_1 _1197_ (.A1(_0484_),
    .A2(_0527_),
    .Y(_0073_),
    .B1(_0528_));
 sg13g2_nor2_1 _1198_ (.A(net40),
    .B(_0287_),
    .Y(_0529_));
 sg13g2_nor2_1 _1199_ (.A(_0304_),
    .B(\desk_clock.clk_seconds[0] ),
    .Y(_0530_));
 sg13g2_a221oi_1 _1200_ (.B2(_0218_),
    .C1(net27),
    .B1(_0530_),
    .A1(_0003_),
    .Y(_0531_),
    .A2(_0529_));
 sg13g2_nand2_1 _1201_ (.Y(_0532_),
    .A(_0304_),
    .B(_0218_));
 sg13g2_nand2_1 _1202_ (.Y(_0533_),
    .A(net27),
    .B(_0294_));
 sg13g2_a21oi_1 _1203_ (.A1(_0003_),
    .A2(_0532_),
    .Y(_0534_),
    .B1(_0533_));
 sg13g2_o21ai_1 _1204_ (.B1(net11),
    .Y(_0535_),
    .A1(_0531_),
    .A2(_0534_));
 sg13g2_o21ai_1 _1205_ (.B1(net32),
    .Y(_0536_),
    .A1(\desk_clock.display_inst.disp_driver.i_data[7] ),
    .A2(_0385_));
 sg13g2_a21oi_1 _1206_ (.A1(_0484_),
    .A2(_0535_),
    .Y(_0075_),
    .B1(_0536_));
 sg13g2_buf_1 _1207_ (.A(_0284_),
    .X(_0537_));
 sg13g2_mux2_1 _1208_ (.A0(\desk_clock.clk_hours[0] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[0] ),
    .S(net9),
    .X(_0538_));
 sg13g2_and2_1 _1209_ (.A(_0168_),
    .B(_0538_),
    .X(_0080_));
 sg13g2_buf_1 _1210_ (.A(_0167_),
    .X(_0539_));
 sg13g2_mux2_1 _1211_ (.A0(\desk_clock.clk_hours[1] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[1] ),
    .S(_0537_),
    .X(_0540_));
 sg13g2_and2_1 _1212_ (.A(net26),
    .B(_0540_),
    .X(_0081_));
 sg13g2_mux2_1 _1213_ (.A0(\desk_clock.clk_hours[2] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[2] ),
    .S(_0537_),
    .X(_0541_));
 sg13g2_and2_1 _1214_ (.A(net26),
    .B(_0541_),
    .X(_0082_));
 sg13g2_mux2_1 _1215_ (.A0(\desk_clock.clk_hours[3] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[3] ),
    .S(net9),
    .X(_0542_));
 sg13g2_and2_1 _1216_ (.A(_0539_),
    .B(_0542_),
    .X(_0083_));
 sg13g2_nor2_1 _1217_ (.A(_0175_),
    .B(_0285_),
    .Y(_0543_));
 sg13g2_a21oi_1 _1218_ (.A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[4] ),
    .A2(_0285_),
    .Y(_0544_),
    .B1(_0543_));
 sg13g2_nor2_1 _1219_ (.A(net29),
    .B(_0544_),
    .Y(_0084_));
 sg13g2_mux2_1 _1220_ (.A0(_0146_),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[0] ),
    .S(net9),
    .X(_0545_));
 sg13g2_and2_1 _1221_ (.A(net26),
    .B(_0545_),
    .X(_0085_));
 sg13g2_mux2_1 _1222_ (.A0(\desk_clock.clk_minutes[1] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[1] ),
    .S(net9),
    .X(_0546_));
 sg13g2_and2_1 _1223_ (.A(net26),
    .B(_0546_),
    .X(_0086_));
 sg13g2_mux2_1 _1224_ (.A0(\desk_clock.clk_minutes[2] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[2] ),
    .S(net9),
    .X(_0547_));
 sg13g2_and2_1 _1225_ (.A(net26),
    .B(_0547_),
    .X(_0087_));
 sg13g2_mux2_1 _1226_ (.A0(\desk_clock.clk_minutes[3] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[3] ),
    .S(net9),
    .X(_0548_));
 sg13g2_and2_1 _1227_ (.A(net26),
    .B(_0548_),
    .X(_0088_));
 sg13g2_mux2_1 _1228_ (.A0(\desk_clock.clk_minutes[4] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[4] ),
    .S(net9),
    .X(_0549_));
 sg13g2_and2_1 _1229_ (.A(net26),
    .B(_0549_),
    .X(_0089_));
 sg13g2_nor2_1 _1230_ (.A(_0182_),
    .B(net10),
    .Y(_0550_));
 sg13g2_a21oi_1 _1231_ (.A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[5] ),
    .A2(net10),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_nor2_1 _1232_ (.A(net29),
    .B(_0551_),
    .Y(_0090_));
 sg13g2_mux2_1 _1233_ (.A0(\desk_clock.clk_seconds[0] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[0] ),
    .S(net9),
    .X(_0552_));
 sg13g2_and2_1 _1234_ (.A(net26),
    .B(_0552_),
    .X(_0091_));
 sg13g2_mux2_1 _1235_ (.A0(\desk_clock.clk_seconds[1] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[1] ),
    .S(_0284_),
    .X(_0553_));
 sg13g2_and2_1 _1236_ (.A(_0539_),
    .B(_0553_),
    .X(_0092_));
 sg13g2_mux2_1 _1237_ (.A0(\desk_clock.clk_seconds[2] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[2] ),
    .S(_0284_),
    .X(_0554_));
 sg13g2_and2_1 _1238_ (.A(net32),
    .B(_0554_),
    .X(_0093_));
 sg13g2_mux2_1 _1239_ (.A0(\desk_clock.clk_seconds[3] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[3] ),
    .S(_0284_),
    .X(_0555_));
 sg13g2_and2_1 _1240_ (.A(net32),
    .B(_0555_),
    .X(_0094_));
 sg13g2_mux2_1 _1241_ (.A0(\desk_clock.clk_seconds[4] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[4] ),
    .S(_0284_),
    .X(_0556_));
 sg13g2_and2_1 _1242_ (.A(_0248_),
    .B(_0556_),
    .X(_0095_));
 sg13g2_mux2_1 _1243_ (.A0(\desk_clock.clk_seconds[5] ),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[5] ),
    .S(_0284_),
    .X(_0557_));
 sg13g2_and2_1 _1244_ (.A(_0248_),
    .B(_0557_),
    .X(_0096_));
 sg13g2_nor2b_1 _1245_ (.A(\desk_clock.clk_gen_inst.stb_gen_debounce_clk.sig_hold ),
    .B_N(\desk_clock.clk_gen_inst.refclk_div[3] ),
    .Y(_0558_));
 sg13g2_buf_1 _1246_ (.A(_0558_),
    .X(_0559_));
 sg13g2_buf_1 _1247_ (.A(_0559_),
    .X(_0560_));
 sg13g2_nand2_1 _1248_ (.Y(_0561_),
    .A(\desk_clock.input_debounce.fast_set_reg[1] ),
    .B(net23));
 sg13g2_buf_1 _1249_ (.A(net25),
    .X(_0562_));
 sg13g2_nand2b_1 _1250_ (.Y(_0563_),
    .B(\desk_clock.input_debounce.fast_set_reg[0] ),
    .A_N(_0562_));
 sg13g2_buf_1 _1251_ (.A(_0258_),
    .X(_0564_));
 sg13g2_a21oi_1 _1252_ (.A1(_0561_),
    .A2(_0563_),
    .Y(_0101_),
    .B1(net21));
 sg13g2_nand2_1 _1253_ (.Y(_0565_),
    .A(\desk_clock.input_debounce.fast_set_reg[2] ),
    .B(net23));
 sg13g2_nand2b_1 _1254_ (.Y(_0566_),
    .B(\desk_clock.input_debounce.fast_set_reg[1] ),
    .A_N(_0562_));
 sg13g2_a21oi_1 _1255_ (.A1(_0565_),
    .A2(_0566_),
    .Y(_0102_),
    .B1(net21));
 sg13g2_nand2_1 _1256_ (.Y(_0567_),
    .A(\desk_clock.input_debounce.fast_set_reg[3] ),
    .B(net23));
 sg13g2_buf_1 _1257_ (.A(net25),
    .X(_0568_));
 sg13g2_nand2b_1 _1258_ (.Y(_0569_),
    .B(\desk_clock.input_debounce.fast_set_reg[2] ),
    .A_N(net20));
 sg13g2_a21oi_1 _1259_ (.A1(_0567_),
    .A2(_0569_),
    .Y(_0103_),
    .B1(net21));
 sg13g2_nand2_1 _1260_ (.Y(_0570_),
    .A(\desk_clock.input_debounce.fast_set_reg[4] ),
    .B(net23));
 sg13g2_nand2b_1 _1261_ (.Y(_0571_),
    .B(\desk_clock.input_debounce.fast_set_reg[3] ),
    .A_N(_0568_));
 sg13g2_a21oi_1 _1262_ (.A1(_0570_),
    .A2(_0571_),
    .Y(_0104_),
    .B1(net21));
 sg13g2_nand2_1 _1263_ (.Y(_0572_),
    .A(\desk_clock.input_debounce.fast_set_reg[5] ),
    .B(_0560_));
 sg13g2_nand2b_1 _1264_ (.Y(_0573_),
    .B(\desk_clock.input_debounce.fast_set_reg[4] ),
    .A_N(_0568_));
 sg13g2_a21oi_1 _1265_ (.A1(_0572_),
    .A2(_0573_),
    .Y(_0105_),
    .B1(_0564_));
 sg13g2_nand2_1 _1266_ (.Y(_0574_),
    .A(net2),
    .B(_0560_));
 sg13g2_nand2b_1 _1267_ (.Y(_0575_),
    .B(\desk_clock.input_debounce.fast_set_reg[5] ),
    .A_N(net20));
 sg13g2_a21oi_1 _1268_ (.A1(_0574_),
    .A2(_0575_),
    .Y(_0106_),
    .B1(_0564_));
 sg13g2_nand2_1 _1269_ (.Y(_0576_),
    .A(\desk_clock.input_debounce.set_hours_reg[1] ),
    .B(net23));
 sg13g2_nand2b_1 _1270_ (.Y(_0577_),
    .B(\desk_clock.input_debounce.set_hours_reg[0] ),
    .A_N(net20));
 sg13g2_a21oi_1 _1271_ (.A1(_0576_),
    .A2(_0577_),
    .Y(_0107_),
    .B1(net21));
 sg13g2_nand2_1 _1272_ (.Y(_0578_),
    .A(\desk_clock.input_debounce.set_hours_reg[2] ),
    .B(net23));
 sg13g2_nand2b_1 _1273_ (.Y(_0579_),
    .B(\desk_clock.input_debounce.set_hours_reg[1] ),
    .A_N(net20));
 sg13g2_a21oi_1 _1274_ (.A1(_0578_),
    .A2(_0579_),
    .Y(_0108_),
    .B1(net21));
 sg13g2_nand2_1 _1275_ (.Y(_0580_),
    .A(\desk_clock.input_debounce.set_hours_reg[3] ),
    .B(net23));
 sg13g2_nand2b_1 _1276_ (.Y(_0581_),
    .B(\desk_clock.input_debounce.set_hours_reg[2] ),
    .A_N(net20));
 sg13g2_a21oi_1 _1277_ (.A1(_0580_),
    .A2(_0581_),
    .Y(_0109_),
    .B1(net21));
 sg13g2_nand2_1 _1278_ (.Y(_0582_),
    .A(\desk_clock.input_debounce.set_hours_reg[4] ),
    .B(net23));
 sg13g2_nand2b_1 _1279_ (.Y(_0583_),
    .B(\desk_clock.input_debounce.set_hours_reg[3] ),
    .A_N(net20));
 sg13g2_a21oi_1 _1280_ (.A1(_0582_),
    .A2(_0583_),
    .Y(_0110_),
    .B1(net21));
 sg13g2_nand2_1 _1281_ (.Y(_0584_),
    .A(\desk_clock.input_debounce.set_hours_reg[5] ),
    .B(net22));
 sg13g2_nand2b_1 _1282_ (.Y(_0585_),
    .B(\desk_clock.input_debounce.set_hours_reg[4] ),
    .A_N(net20));
 sg13g2_a21oi_1 _1283_ (.A1(_0584_),
    .A2(_0585_),
    .Y(_0111_),
    .B1(net28));
 sg13g2_nand2_1 _1284_ (.Y(_0586_),
    .A(net3),
    .B(net22));
 sg13g2_nand2b_1 _1285_ (.Y(_0587_),
    .B(\desk_clock.input_debounce.set_hours_reg[5] ),
    .A_N(net20));
 sg13g2_a21oi_1 _1286_ (.A1(_0586_),
    .A2(_0587_),
    .Y(_0112_),
    .B1(net28));
 sg13g2_nand2_1 _1287_ (.Y(_0588_),
    .A(\desk_clock.input_debounce.set_minutes_reg[1] ),
    .B(net22));
 sg13g2_nand2b_1 _1288_ (.Y(_0589_),
    .B(\desk_clock.input_debounce.set_minutes_reg[0] ),
    .A_N(net25));
 sg13g2_a21oi_1 _1289_ (.A1(_0588_),
    .A2(_0589_),
    .Y(_0113_),
    .B1(net28));
 sg13g2_nand2_1 _1290_ (.Y(_0590_),
    .A(\desk_clock.input_debounce.set_minutes_reg[2] ),
    .B(net22));
 sg13g2_nand2b_1 _1291_ (.Y(_0591_),
    .B(\desk_clock.input_debounce.set_minutes_reg[1] ),
    .A_N(net25));
 sg13g2_a21oi_1 _1292_ (.A1(_0590_),
    .A2(_0591_),
    .Y(_0114_),
    .B1(net28));
 sg13g2_nand2_1 _1293_ (.Y(_0592_),
    .A(\desk_clock.input_debounce.set_minutes_reg[3] ),
    .B(net22));
 sg13g2_nand2b_1 _1294_ (.Y(_0593_),
    .B(\desk_clock.input_debounce.set_minutes_reg[2] ),
    .A_N(net25));
 sg13g2_a21oi_1 _1295_ (.A1(_0592_),
    .A2(_0593_),
    .Y(_0115_),
    .B1(net28));
 sg13g2_nand2_1 _1296_ (.Y(_0594_),
    .A(\desk_clock.input_debounce.set_minutes_reg[4] ),
    .B(net22));
 sg13g2_nand2b_1 _1297_ (.Y(_0595_),
    .B(\desk_clock.input_debounce.set_minutes_reg[3] ),
    .A_N(net25));
 sg13g2_a21oi_1 _1298_ (.A1(_0594_),
    .A2(_0595_),
    .Y(_0116_),
    .B1(net28));
 sg13g2_nand2_1 _1299_ (.Y(_0596_),
    .A(\desk_clock.input_debounce.set_minutes_reg[5] ),
    .B(net22));
 sg13g2_nand2b_1 _1300_ (.Y(_0597_),
    .B(\desk_clock.input_debounce.set_minutes_reg[4] ),
    .A_N(net25));
 sg13g2_a21oi_1 _1301_ (.A1(_0596_),
    .A2(_0597_),
    .Y(_0117_),
    .B1(_0350_));
 sg13g2_nand2_1 _1302_ (.Y(_0598_),
    .A(net4),
    .B(net22));
 sg13g2_nand2b_1 _1303_ (.Y(_0599_),
    .B(\desk_clock.input_debounce.set_minutes_reg[5] ),
    .A_N(net25));
 sg13g2_a21oi_1 _1304_ (.A1(_0598_),
    .A2(_0599_),
    .Y(_0118_),
    .B1(_0350_));
 sg13g2_and2_1 _1305_ (.A(net32),
    .B(net1),
    .X(_0119_));
 sg13g2_and2_1 _1306_ (.A(net32),
    .B(\desk_clock.refclk_sync_inst.refclk_sync_reg[0] ),
    .X(_0120_));
 sg13g2_nor2_1 _1307_ (.A(clknet_5_14__leaf_clk),
    .B(\desk_clock.display_inst.disp_driver.o_serial_load ),
    .Y(\desk_clock.display_inst.disp_driver.o_serial_clk ));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _1310__60 (.L_HI(net60));
 sg13g2_buf_1 _1310_ (.A(net60),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1311_ (.A(net61),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1312_ (.A(net41),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1313_ (.A(net62),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1314_ (.A(net42),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1315_ (.A(net43),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1316_ (.A(net44),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1317_ (.A(net45),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1318_ (.A(\desk_clock.display_inst.disp_driver.o_serial_load ),
    .X(net5));
 sg13g2_buf_1 _1319_ (.A(\desk_clock.display_inst.disp_driver.data_reg[15] ),
    .X(net6));
 sg13g2_buf_1 _1320_ (.A(net46),
    .X(uio_out[2]));
 sg13g2_buf_1 _1321_ (.A(\desk_clock.display_inst.disp_driver.o_serial_clk ),
    .X(net7));
 sg13g2_buf_1 _1322_ (.A(net47),
    .X(uio_out[4]));
 sg13g2_buf_1 _1323_ (.A(net48),
    .X(uio_out[5]));
 sg13g2_buf_1 _1324_ (.A(net49),
    .X(uio_out[6]));
 sg13g2_buf_1 _1325_ (.A(net50),
    .X(uio_out[7]));
 sg13g2_buf_1 _1326_ (.A(net51),
    .X(uo_out[0]));
 sg13g2_buf_1 _1327_ (.A(net52),
    .X(uo_out[1]));
 sg13g2_buf_1 _1328_ (.A(net53),
    .X(uo_out[2]));
 sg13g2_buf_1 _1329_ (.A(net54),
    .X(uo_out[3]));
 sg13g2_buf_1 _1330_ (.A(net55),
    .X(uo_out[4]));
 sg13g2_buf_1 _1331_ (.A(net56),
    .X(uo_out[5]));
 sg13g2_buf_1 _1332_ (.A(net57),
    .X(uo_out[6]));
 sg13g2_buf_1 _1333_ (.A(net58),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[0]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net63),
    .D(_0006_),
    .Q_N(_0005_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[0] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[10]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net64),
    .D(_0007_),
    .Q_N(_0709_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[10] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[11]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net65),
    .D(_0008_),
    .Q_N(_0708_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[11] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[12]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net66),
    .D(_0009_),
    .Q_N(_0707_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[12] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[13]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net67),
    .D(_0010_),
    .Q_N(_0706_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[13] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[14]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net68),
    .D(_0011_),
    .Q_N(_0705_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[14] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[1]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net69),
    .D(_0012_),
    .Q_N(_0704_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[1] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[2]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net70),
    .D(_0013_),
    .Q_N(_0703_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[2] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[3]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net71),
    .D(_0014_),
    .Q_N(_0702_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[3] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[4]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net72),
    .D(_0015_),
    .Q_N(_0701_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[4] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[5]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net73),
    .D(_0016_),
    .Q_N(_0700_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[5] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[6]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net74),
    .D(_0017_),
    .Q_N(_0699_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[6] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[7]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net75),
    .D(_0018_),
    .Q_N(_0698_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[7] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[8]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net76),
    .D(_0019_),
    .Q_N(_0697_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[8] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.refclk_div[9]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net77),
    .D(_0020_),
    .Q_N(_0696_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[9] ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.stb_gen_1hz.sig_hold$_SDFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net78),
    .D(_0021_),
    .Q_N(_0695_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_1hz.sig_hold ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.stb_gen_debounce_clk.sig_hold$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net79),
    .D(_0022_),
    .Q_N(_0694_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_debounce_clk.sig_hold ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.stb_gen_fast_clk.sig_hold$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net80),
    .D(_0023_),
    .Q_N(_0693_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_fast_clk.sig_hold ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.stb_gen_refclk.sig_hold$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net81),
    .D(_0024_),
    .Q_N(_0692_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_refclk.sig_hold ));
 sg13g2_dfrbp_1 \desk_clock.clk_gen_inst.stb_gen_slow_clk.sig_hold$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net82),
    .D(_0025_),
    .Q_N(_0691_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_slow_clk.sig_hold ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_hours[0]$_SDFFE_PP0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net83),
    .D(_0026_),
    .Q_N(_0690_),
    .Q(\desk_clock.clk_hours[0] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_hours[1]$_SDFFE_PP0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net84),
    .D(_0027_),
    .Q_N(_0689_),
    .Q(\desk_clock.clk_hours[1] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_hours[2]$_SDFFE_PP0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net85),
    .D(_0028_),
    .Q_N(_0688_),
    .Q(\desk_clock.clk_hours[2] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_hours[3]$_SDFFE_PP0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net86),
    .D(_0029_),
    .Q_N(_0687_),
    .Q(\desk_clock.clk_hours[3] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_hours[4]$_SDFFE_PP0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net87),
    .D(_0030_),
    .Q_N(_0686_),
    .Q(\desk_clock.clk_hours[4] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_minutes[0]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net88),
    .D(_0031_),
    .Q_N(_0685_),
    .Q(\desk_clock.clk_minutes[0] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_minutes[1]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net89),
    .D(_0032_),
    .Q_N(_0684_),
    .Q(\desk_clock.clk_minutes[1] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_minutes[2]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net90),
    .D(_0033_),
    .Q_N(_0683_),
    .Q(\desk_clock.clk_minutes[2] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_minutes[3]$_SDFFE_PP0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net91),
    .D(_0034_),
    .Q_N(_0682_),
    .Q(\desk_clock.clk_minutes[3] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_minutes[4]$_SDFFE_PP0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net92),
    .D(_0035_),
    .Q_N(_0681_),
    .Q(\desk_clock.clk_minutes[4] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_minutes[5]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net93),
    .D(_0036_),
    .Q_N(_0680_),
    .Q(\desk_clock.clk_minutes[5] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_seconds[0]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net94),
    .D(_0037_),
    .Q_N(_0679_),
    .Q(\desk_clock.clk_seconds[0] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_seconds[1]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net95),
    .D(_0038_),
    .Q_N(_0678_),
    .Q(\desk_clock.clk_seconds[1] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_seconds[2]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net96),
    .D(_0039_),
    .Q_N(_0677_),
    .Q(\desk_clock.clk_seconds[2] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_seconds[3]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net97),
    .D(_0040_),
    .Q_N(_0676_),
    .Q(\desk_clock.clk_seconds[3] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_seconds[4]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net98),
    .D(_0041_),
    .Q_N(_0675_),
    .Q(\desk_clock.clk_seconds[4] ));
 sg13g2_dfrbp_1 \desk_clock.clock_reg_inst.o_seconds[5]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net99),
    .D(_0042_),
    .Q_N(_0674_),
    .Q(\desk_clock.clk_seconds[5] ));
 sg13g2_dfrbp_1 \desk_clock.display_control_inst.display_update$_SDFF_PP1_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net100),
    .D(_0043_),
    .Q_N(_0673_),
    .Q(\desk_clock.display_control_inst.display_update ));
 sg13g2_dfrbp_1 \desk_clock.display_control_inst.startup$_SDFFE_PN1P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net101),
    .D(_0044_),
    .Q_N(_0000_),
    .Q(\desk_clock.display_control_inst.o_write_config ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net102),
    .D(_0045_),
    .Q_N(_0672_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[0] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[10]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net103),
    .D(_0046_),
    .Q_N(_0671_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[10] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[11]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net104),
    .D(_0047_),
    .Q_N(_0670_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[11] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[12]$_SDFFE_PP0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net105),
    .D(_0048_),
    .Q_N(_0669_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[12] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[13]$_SDFFE_PP0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net106),
    .D(_0049_),
    .Q_N(_0668_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[13] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[14]$_SDFFE_PP0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net107),
    .D(_0050_),
    .Q_N(_0667_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[14] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[15]$_SDFFE_PP0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net108),
    .D(_0051_),
    .Q_N(_0666_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[15] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net109),
    .D(_0052_),
    .Q_N(_0665_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[1] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net110),
    .D(_0053_),
    .Q_N(_0664_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[2] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net111),
    .D(_0054_),
    .Q_N(_0663_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[3] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net112),
    .D(_0055_),
    .Q_N(_0662_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[4] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net113),
    .D(_0056_),
    .Q_N(_0661_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[5] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[6]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net114),
    .D(_0057_),
    .Q_N(_0660_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[6] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[7]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net115),
    .D(_0058_),
    .Q_N(_0659_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[7] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[8]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net116),
    .D(_0059_),
    .Q_N(_0658_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[8] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.data_reg[9]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net117),
    .D(_0060_),
    .Q_N(_0657_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[9] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.transfer_state[0]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net118),
    .D(_0061_),
    .Q_N(_0001_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[0] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.transfer_state[1]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net119),
    .D(_0062_),
    .Q_N(_0656_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[1] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.transfer_state[2]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net120),
    .D(_0063_),
    .Q_N(_0655_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[2] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.transfer_state[3]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net121),
    .D(_0064_),
    .Q_N(_0654_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[3] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.disp_driver.transfer_state[4]$_SDFFE_PP0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net122),
    .D(_0065_),
    .Q_N(_0653_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[4] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_addr[0]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net123),
    .D(_0066_),
    .Q_N(_0652_),
    .Q(\desk_clock.display_inst.disp_driver.i_addr[0] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_addr[1]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net124),
    .D(_0067_),
    .Q_N(_0651_),
    .Q(\desk_clock.display_inst.disp_driver.i_addr[1] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_addr[2]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net125),
    .D(_0068_),
    .Q_N(_0650_),
    .Q(\desk_clock.display_inst.disp_driver.i_addr[2] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_addr[3]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net126),
    .D(_0069_),
    .Q_N(_0649_),
    .Q(\desk_clock.display_inst.disp_driver.i_addr[3] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_data[0]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net127),
    .D(_0070_),
    .Q_N(_0648_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[0] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_data[1]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net128),
    .D(_0071_),
    .Q_N(_0647_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[1] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_data[2]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net129),
    .D(_0072_),
    .Q_N(_0646_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[2] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_data[3]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net130),
    .D(_0073_),
    .Q_N(_0645_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[3] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_data[5]$_SDFFE_PP0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net131),
    .D(_0074_),
    .Q_N(_0644_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[4] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.o_data[7]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net132),
    .D(_0075_),
    .Q_N(_0643_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[7] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.transfer_state[0]$_SDFFE_PP0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net133),
    .D(_0076_),
    .Q_N(_0004_),
    .Q(\desk_clock.display_inst.display_settings.transfer_state[0] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.transfer_state[1]$_SDFFE_PP0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net134),
    .D(_0077_),
    .Q_N(_0642_),
    .Q(\desk_clock.display_inst.display_settings.transfer_state[1] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.transfer_state[2]$_SDFFE_PP0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net135),
    .D(_0078_),
    .Q_N(_0641_),
    .Q(\desk_clock.display_inst.display_settings.transfer_state[2] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.transfer_state[3]$_SDFFE_PP0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net136),
    .D(net59),
    .Q_N(_0640_),
    .Q(\desk_clock.display_inst.display_settings.transfer_state[3] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.display_settings.write_config$_DFFE_PP_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net137),
    .D(_0079_),
    .Q_N(_0639_),
    .Q(\desk_clock.display_inst.display_settings.write_config ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.hours_int[0]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net138),
    .D(_0080_),
    .Q_N(_0638_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[0] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.hours_int[1]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net139),
    .D(_0081_),
    .Q_N(_0637_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[1] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.hours_int[2]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net140),
    .D(_0082_),
    .Q_N(_0636_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[2] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.hours_int[3]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net141),
    .D(_0083_),
    .Q_N(_0635_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[3] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.hours_int[4]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net142),
    .D(_0084_),
    .Q_N(_0634_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[4] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.minutes_int[0]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net143),
    .D(_0085_),
    .Q_N(_0633_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[0] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.minutes_int[1]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net144),
    .D(_0086_),
    .Q_N(_0632_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[1] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.minutes_int[2]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net145),
    .D(_0087_),
    .Q_N(_0631_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[2] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.minutes_int[3]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net146),
    .D(_0088_),
    .Q_N(_0630_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[3] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.minutes_int[4]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net147),
    .D(_0089_),
    .Q_N(_0629_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[4] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.minutes_int[5]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net148),
    .D(_0090_),
    .Q_N(_0628_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[5] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.seconds_int[0]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net149),
    .D(_0091_),
    .Q_N(_0627_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[0] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.seconds_int[1]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net150),
    .D(_0092_),
    .Q_N(_0626_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[1] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.seconds_int[2]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net151),
    .D(_0093_),
    .Q_N(_0625_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[2] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.seconds_int[3]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net152),
    .D(_0094_),
    .Q_N(_0624_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[3] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.seconds_int[4]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net153),
    .D(_0095_),
    .Q_N(_0623_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[4] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.seconds_int[5]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net154),
    .D(_0096_),
    .Q_N(_0622_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[5] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.state[0]$_SDFFE_PP0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net155),
    .D(_0097_),
    .Q_N(_0002_),
    .Q(\desk_clock.display_inst.state[0] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.state[1]$_SDFFE_PP0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net156),
    .D(_0098_),
    .Q_N(_0003_),
    .Q(\desk_clock.display_inst.state[1] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.state[2]$_SDFFE_PP0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net157),
    .D(_0099_),
    .Q_N(_0621_),
    .Q(\desk_clock.display_inst.state[2] ));
 sg13g2_dfrbp_1 \desk_clock.display_inst.state[3]$_SDFFE_PP0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net158),
    .D(_0100_),
    .Q_N(_0620_),
    .Q(\desk_clock.display_inst.state[3] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.fast_set_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net159),
    .D(_0101_),
    .Q_N(_0619_),
    .Q(\desk_clock.input_debounce.fast_set_reg[0] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.fast_set_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net160),
    .D(_0102_),
    .Q_N(_0618_),
    .Q(\desk_clock.input_debounce.fast_set_reg[1] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.fast_set_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net161),
    .D(_0103_),
    .Q_N(_0617_),
    .Q(\desk_clock.input_debounce.fast_set_reg[2] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.fast_set_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net162),
    .D(_0104_),
    .Q_N(_0616_),
    .Q(\desk_clock.input_debounce.fast_set_reg[3] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.fast_set_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net163),
    .D(_0105_),
    .Q_N(_0615_),
    .Q(\desk_clock.input_debounce.fast_set_reg[4] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.fast_set_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net164),
    .D(_0106_),
    .Q_N(_0614_),
    .Q(\desk_clock.input_debounce.fast_set_reg[5] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_hours_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net165),
    .D(_0107_),
    .Q_N(_0613_),
    .Q(\desk_clock.input_debounce.set_hours_reg[0] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_hours_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net166),
    .D(_0108_),
    .Q_N(_0612_),
    .Q(\desk_clock.input_debounce.set_hours_reg[1] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_hours_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net167),
    .D(_0109_),
    .Q_N(_0611_),
    .Q(\desk_clock.input_debounce.set_hours_reg[2] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_hours_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net168),
    .D(_0110_),
    .Q_N(_0610_),
    .Q(\desk_clock.input_debounce.set_hours_reg[3] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_hours_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net169),
    .D(_0111_),
    .Q_N(_0609_),
    .Q(\desk_clock.input_debounce.set_hours_reg[4] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_hours_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net170),
    .D(_0112_),
    .Q_N(_0608_),
    .Q(\desk_clock.input_debounce.set_hours_reg[5] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_minutes_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net171),
    .D(_0113_),
    .Q_N(_0607_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[0] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_minutes_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net172),
    .D(_0114_),
    .Q_N(_0606_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[1] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_minutes_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net173),
    .D(_0115_),
    .Q_N(_0605_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[2] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_minutes_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net174),
    .D(_0116_),
    .Q_N(_0604_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[3] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_minutes_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net175),
    .D(_0117_),
    .Q_N(_0603_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[4] ));
 sg13g2_dfrbp_1 \desk_clock.input_debounce.set_minutes_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net176),
    .D(_0118_),
    .Q_N(_0602_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[5] ));
 sg13g2_dfrbp_1 \desk_clock.refclk_sync_inst.refclk_sync_reg[0]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net177),
    .D(_0119_),
    .Q_N(_0601_),
    .Q(\desk_clock.refclk_sync_inst.refclk_sync_reg[0] ));
 sg13g2_dfrbp_1 \desk_clock.refclk_sync_inst.refclk_sync_reg[1]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net178),
    .D(_0120_),
    .Q_N(_0600_),
    .Q(\desk_clock.clk_gen_inst.i_refclk ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[0]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[1]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[3]));
 sg13g2_buf_2 fanout8 (.A(_0450_),
    .X(net8));
 sg13g2_buf_4 fanout9 (.X(net9),
    .A(_0537_));
 sg13g2_buf_2 fanout10 (.A(_0285_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_0260_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0247_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0452_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0409_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(\desk_clock.display_inst.disp_driver.o_serial_load ),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0352_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0238_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0237_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0233_),
    .X(net19));
 sg13g2_buf_1 fanout20 (.A(_0568_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0564_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0562_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0560_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0310_),
    .X(net24));
 sg13g2_buf_1 fanout25 (.A(_0559_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0539_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0396_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0350_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0340_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0294_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0258_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0248_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0168_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0229_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0228_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0167_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0131_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0126_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0123_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0122_),
    .X(net40));
 sg13g2_tielo _1312__41 (.L_LO(net41));
 sg13g2_tielo _1314__42 (.L_LO(net42));
 sg13g2_tielo _1315__43 (.L_LO(net43));
 sg13g2_tielo _1316__44 (.L_LO(net44));
 sg13g2_tielo _1317__45 (.L_LO(net45));
 sg13g2_tielo _1320__46 (.L_LO(net46));
 sg13g2_tielo _1322__47 (.L_LO(net47));
 sg13g2_tielo _1323__48 (.L_LO(net48));
 sg13g2_tielo _1324__49 (.L_LO(net49));
 sg13g2_tielo _1325__50 (.L_LO(net50));
 sg13g2_tielo _1326__51 (.L_LO(net51));
 sg13g2_tielo _1327__52 (.L_LO(net52));
 sg13g2_tielo _1328__53 (.L_LO(net53));
 sg13g2_tielo _1329__54 (.L_LO(net54));
 sg13g2_tielo _1330__55 (.L_LO(net55));
 sg13g2_tielo _1331__56 (.L_LO(net56));
 sg13g2_tielo _1332__57 (.L_LO(net57));
 sg13g2_tielo _1333__58 (.L_LO(net58));
 sg13g2_tielo \desk_clock.display_inst.display_settings.transfer_state[3]$_SDFFE_PP0P__59  (.L_LO(net59));
 sg13g2_tiehi _1311__61 (.L_HI(net61));
 sg13g2_tiehi _1313__62 (.L_HI(net62));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[0]$_SDFFE_PN0P__63  (.L_HI(net63));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[10]$_SDFFE_PN0P__64  (.L_HI(net64));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[11]$_SDFFE_PN0P__65  (.L_HI(net65));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[12]$_SDFFE_PN0P__66  (.L_HI(net66));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[13]$_SDFFE_PN0P__67  (.L_HI(net67));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[14]$_SDFFE_PN0P__68  (.L_HI(net68));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[1]$_SDFFE_PN0P__69  (.L_HI(net69));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[2]$_SDFFE_PN0P__70  (.L_HI(net70));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[3]$_SDFFE_PN0P__71  (.L_HI(net71));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[4]$_SDFFE_PN0P__72  (.L_HI(net72));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[5]$_SDFFE_PN0P__73  (.L_HI(net73));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[6]$_SDFFE_PN0P__74  (.L_HI(net74));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[7]$_SDFFE_PN0P__75  (.L_HI(net75));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[8]$_SDFFE_PN0P__76  (.L_HI(net76));
 sg13g2_tiehi \desk_clock.clk_gen_inst.refclk_div[9]$_SDFFE_PN0P__77  (.L_HI(net77));
 sg13g2_tiehi \desk_clock.clk_gen_inst.stb_gen_1hz.sig_hold$_SDFF_PN0__78  (.L_HI(net78));
 sg13g2_tiehi \desk_clock.clk_gen_inst.stb_gen_debounce_clk.sig_hold$_SDFF_PN0__79  (.L_HI(net79));
 sg13g2_tiehi \desk_clock.clk_gen_inst.stb_gen_fast_clk.sig_hold$_SDFF_PN0__80  (.L_HI(net80));
 sg13g2_tiehi \desk_clock.clk_gen_inst.stb_gen_refclk.sig_hold$_SDFF_PN0__81  (.L_HI(net81));
 sg13g2_tiehi \desk_clock.clk_gen_inst.stb_gen_slow_clk.sig_hold$_SDFF_PN0__82  (.L_HI(net82));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_hours[0]$_SDFFE_PP0P__83  (.L_HI(net83));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_hours[1]$_SDFFE_PP0P__84  (.L_HI(net84));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_hours[2]$_SDFFE_PP0P__85  (.L_HI(net85));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_hours[3]$_SDFFE_PP0P__86  (.L_HI(net86));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_hours[4]$_SDFFE_PP0P__87  (.L_HI(net87));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_minutes[0]$_SDFFE_PP0P__88  (.L_HI(net88));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_minutes[1]$_SDFFE_PP0P__89  (.L_HI(net89));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_minutes[2]$_SDFFE_PP0P__90  (.L_HI(net90));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_minutes[3]$_SDFFE_PP0P__91  (.L_HI(net91));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_minutes[4]$_SDFFE_PP0P__92  (.L_HI(net92));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_minutes[5]$_SDFFE_PP0P__93  (.L_HI(net93));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_seconds[0]$_SDFFE_PP0P__94  (.L_HI(net94));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_seconds[1]$_SDFFE_PP0P__95  (.L_HI(net95));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_seconds[2]$_SDFFE_PP0P__96  (.L_HI(net96));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_seconds[3]$_SDFFE_PP0P__97  (.L_HI(net97));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_seconds[4]$_SDFFE_PP0P__98  (.L_HI(net98));
 sg13g2_tiehi \desk_clock.clock_reg_inst.o_seconds[5]$_SDFFE_PP0P__99  (.L_HI(net99));
 sg13g2_tiehi \desk_clock.display_control_inst.display_update$_SDFF_PP1__100  (.L_HI(net100));
 sg13g2_tiehi \desk_clock.display_control_inst.startup$_SDFFE_PN1P__101  (.L_HI(net101));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[0]$_SDFFE_PN0P__102  (.L_HI(net102));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[10]$_SDFFE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[11]$_SDFFE_PN0P__104  (.L_HI(net104));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[12]$_SDFFE_PP0P__105  (.L_HI(net105));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[13]$_SDFFE_PP0P__106  (.L_HI(net106));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[14]$_SDFFE_PP0P__107  (.L_HI(net107));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[15]$_SDFFE_PP0P__108  (.L_HI(net108));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[1]$_SDFFE_PN0P__109  (.L_HI(net109));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[2]$_SDFFE_PN0P__110  (.L_HI(net110));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[3]$_SDFFE_PN0P__111  (.L_HI(net111));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[4]$_SDFFE_PN0P__112  (.L_HI(net112));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[5]$_SDFFE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[6]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[7]$_SDFFE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[8]$_SDFFE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.data_reg[9]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.transfer_state[0]$_SDFFE_PP0P__118  (.L_HI(net118));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.transfer_state[1]$_SDFFE_PP0P__119  (.L_HI(net119));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.transfer_state[2]$_SDFFE_PP0P__120  (.L_HI(net120));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.transfer_state[3]$_SDFFE_PP0P__121  (.L_HI(net121));
 sg13g2_tiehi \desk_clock.display_inst.disp_driver.transfer_state[4]$_SDFFE_PP0P__122  (.L_HI(net122));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_addr[0]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_addr[1]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_addr[2]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_addr[3]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_data[0]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_data[1]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_data[2]$_SDFFE_PN0P__129  (.L_HI(net129));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_data[3]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_data[5]$_SDFFE_PP0P__131  (.L_HI(net131));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.o_data[7]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.transfer_state[0]$_SDFFE_PP0P__133  (.L_HI(net133));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.transfer_state[1]$_SDFFE_PP0P__134  (.L_HI(net134));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.transfer_state[2]$_SDFFE_PP0P__135  (.L_HI(net135));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.transfer_state[3]$_SDFFE_PP0P__136  (.L_HI(net136));
 sg13g2_tiehi \desk_clock.display_inst.display_settings.write_config$_DFFE_PP__137  (.L_HI(net137));
 sg13g2_tiehi \desk_clock.display_inst.hours_int[0]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \desk_clock.display_inst.hours_int[1]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \desk_clock.display_inst.hours_int[2]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \desk_clock.display_inst.hours_int[3]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \desk_clock.display_inst.hours_int[4]$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \desk_clock.display_inst.minutes_int[0]$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \desk_clock.display_inst.minutes_int[1]$_SDFFE_PN0P__144  (.L_HI(net144));
 sg13g2_tiehi \desk_clock.display_inst.minutes_int[2]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \desk_clock.display_inst.minutes_int[3]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \desk_clock.display_inst.minutes_int[4]$_SDFFE_PN0P__147  (.L_HI(net147));
 sg13g2_tiehi \desk_clock.display_inst.minutes_int[5]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \desk_clock.display_inst.seconds_int[0]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \desk_clock.display_inst.seconds_int[1]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \desk_clock.display_inst.seconds_int[2]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \desk_clock.display_inst.seconds_int[3]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \desk_clock.display_inst.seconds_int[4]$_SDFFE_PN0P__153  (.L_HI(net153));
 sg13g2_tiehi \desk_clock.display_inst.seconds_int[5]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \desk_clock.display_inst.state[0]$_SDFFE_PP0P__155  (.L_HI(net155));
 sg13g2_tiehi \desk_clock.display_inst.state[1]$_SDFFE_PP0P__156  (.L_HI(net156));
 sg13g2_tiehi \desk_clock.display_inst.state[2]$_SDFFE_PP0P__157  (.L_HI(net157));
 sg13g2_tiehi \desk_clock.display_inst.state[3]$_SDFFE_PP0P__158  (.L_HI(net158));
 sg13g2_tiehi \desk_clock.input_debounce.fast_set_reg[0]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \desk_clock.input_debounce.fast_set_reg[1]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \desk_clock.input_debounce.fast_set_reg[2]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \desk_clock.input_debounce.fast_set_reg[3]$_SDFFE_PN0P__162  (.L_HI(net162));
 sg13g2_tiehi \desk_clock.input_debounce.fast_set_reg[4]$_SDFFE_PN0P__163  (.L_HI(net163));
 sg13g2_tiehi \desk_clock.input_debounce.fast_set_reg[5]$_SDFFE_PN0P__164  (.L_HI(net164));
 sg13g2_tiehi \desk_clock.input_debounce.set_hours_reg[0]$_SDFFE_PN0P__165  (.L_HI(net165));
 sg13g2_tiehi \desk_clock.input_debounce.set_hours_reg[1]$_SDFFE_PN0P__166  (.L_HI(net166));
 sg13g2_tiehi \desk_clock.input_debounce.set_hours_reg[2]$_SDFFE_PN0P__167  (.L_HI(net167));
 sg13g2_tiehi \desk_clock.input_debounce.set_hours_reg[3]$_SDFFE_PN0P__168  (.L_HI(net168));
 sg13g2_tiehi \desk_clock.input_debounce.set_hours_reg[4]$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \desk_clock.input_debounce.set_hours_reg[5]$_SDFFE_PN0P__170  (.L_HI(net170));
 sg13g2_tiehi \desk_clock.input_debounce.set_minutes_reg[0]$_SDFFE_PN0P__171  (.L_HI(net171));
 sg13g2_tiehi \desk_clock.input_debounce.set_minutes_reg[1]$_SDFFE_PN0P__172  (.L_HI(net172));
 sg13g2_tiehi \desk_clock.input_debounce.set_minutes_reg[2]$_SDFFE_PN0P__173  (.L_HI(net173));
 sg13g2_tiehi \desk_clock.input_debounce.set_minutes_reg[3]$_SDFFE_PN0P__174  (.L_HI(net174));
 sg13g2_tiehi \desk_clock.input_debounce.set_minutes_reg[4]$_SDFFE_PN0P__175  (.L_HI(net175));
 sg13g2_tiehi \desk_clock.input_debounce.set_minutes_reg[5]$_SDFFE_PN0P__176  (.L_HI(net176));
 sg13g2_tiehi \desk_clock.refclk_sync_inst.refclk_sync_reg[0]$_SDFF_PN0__177  (.L_HI(net177));
 sg13g2_tiehi \desk_clock.refclk_sync_inst.refclk_sync_reg[1]$_SDFF_PN0__178  (.L_HI(net178));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_31__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_4 FILLER_10_203 ();
 sg13g2_decap_4 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_decap_8 FILLER_10_227 ();
 sg13g2_decap_8 FILLER_10_234 ();
 sg13g2_decap_4 FILLER_10_241 ();
 sg13g2_decap_4 FILLER_10_250 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_decap_8 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_321 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_8 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_10_412 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_decap_4 FILLER_10_426 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_163 ();
 sg13g2_fill_2 FILLER_11_170 ();
 sg13g2_fill_1 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_decap_8 FILLER_11_191 ();
 sg13g2_fill_2 FILLER_11_198 ();
 sg13g2_fill_1 FILLER_11_200 ();
 sg13g2_decap_4 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_4 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_11_409 ();
 sg13g2_decap_8 FILLER_11_416 ();
 sg13g2_decap_8 FILLER_11_423 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_4 FILLER_12_126 ();
 sg13g2_fill_2 FILLER_12_130 ();
 sg13g2_fill_2 FILLER_12_158 ();
 sg13g2_fill_1 FILLER_12_160 ();
 sg13g2_fill_1 FILLER_12_202 ();
 sg13g2_fill_2 FILLER_12_223 ();
 sg13g2_decap_8 FILLER_12_229 ();
 sg13g2_decap_4 FILLER_12_236 ();
 sg13g2_decap_4 FILLER_12_252 ();
 sg13g2_fill_2 FILLER_12_256 ();
 sg13g2_fill_2 FILLER_12_275 ();
 sg13g2_fill_1 FILLER_12_277 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_decap_8 FILLER_12_332 ();
 sg13g2_decap_8 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_12_409 ();
 sg13g2_decap_8 FILLER_12_416 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_121 ();
 sg13g2_decap_8 FILLER_13_128 ();
 sg13g2_decap_4 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_139 ();
 sg13g2_decap_8 FILLER_13_144 ();
 sg13g2_decap_4 FILLER_13_151 ();
 sg13g2_decap_4 FILLER_13_164 ();
 sg13g2_fill_2 FILLER_13_168 ();
 sg13g2_decap_4 FILLER_13_180 ();
 sg13g2_fill_2 FILLER_13_184 ();
 sg13g2_decap_4 FILLER_13_191 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_213 ();
 sg13g2_fill_1 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_4 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_fill_2 FILLER_13_306 ();
 sg13g2_fill_1 FILLER_13_312 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_fill_2 FILLER_13_327 ();
 sg13g2_fill_2 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_4 FILLER_13_424 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_4 FILLER_14_105 ();
 sg13g2_fill_1 FILLER_14_109 ();
 sg13g2_fill_2 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_138 ();
 sg13g2_decap_4 FILLER_14_180 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_fill_2 FILLER_14_211 ();
 sg13g2_fill_1 FILLER_14_213 ();
 sg13g2_decap_4 FILLER_14_219 ();
 sg13g2_fill_1 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_fill_2 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_274 ();
 sg13g2_fill_2 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_317 ();
 sg13g2_fill_2 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_fill_2 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_121 ();
 sg13g2_decap_4 FILLER_15_125 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_decap_8 FILLER_15_162 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_decap_8 FILLER_15_180 ();
 sg13g2_decap_4 FILLER_15_187 ();
 sg13g2_decap_4 FILLER_15_195 ();
 sg13g2_fill_2 FILLER_15_199 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_228 ();
 sg13g2_fill_1 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_fill_1 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_fill_2 FILLER_15_326 ();
 sg13g2_fill_1 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_366 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_decap_8 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_4 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_79 ();
 sg13g2_fill_2 FILLER_16_86 ();
 sg13g2_decap_4 FILLER_16_92 ();
 sg13g2_fill_2 FILLER_16_96 ();
 sg13g2_decap_4 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_113 ();
 sg13g2_decap_8 FILLER_16_120 ();
 sg13g2_decap_4 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_131 ();
 sg13g2_fill_2 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_fill_1 FILLER_16_159 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_fill_2 FILLER_16_187 ();
 sg13g2_decap_8 FILLER_16_229 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_decap_4 FILLER_16_245 ();
 sg13g2_decap_4 FILLER_16_253 ();
 sg13g2_decap_4 FILLER_16_267 ();
 sg13g2_decap_4 FILLER_16_278 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_decap_4 FILLER_16_293 ();
 sg13g2_fill_2 FILLER_16_312 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_decap_4 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_16_409 ();
 sg13g2_decap_8 FILLER_16_416 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_118 ();
 sg13g2_decap_4 FILLER_17_127 ();
 sg13g2_decap_8 FILLER_17_135 ();
 sg13g2_fill_2 FILLER_17_142 ();
 sg13g2_fill_1 FILLER_17_144 ();
 sg13g2_decap_8 FILLER_17_180 ();
 sg13g2_decap_8 FILLER_17_187 ();
 sg13g2_fill_2 FILLER_17_194 ();
 sg13g2_fill_1 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_fill_2 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_270 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_decap_4 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_295 ();
 sg13g2_fill_1 FILLER_17_302 ();
 sg13g2_fill_2 FILLER_17_311 ();
 sg13g2_fill_1 FILLER_17_313 ();
 sg13g2_decap_4 FILLER_17_321 ();
 sg13g2_fill_2 FILLER_17_325 ();
 sg13g2_fill_2 FILLER_17_332 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_decap_4 FILLER_17_361 ();
 sg13g2_fill_2 FILLER_17_365 ();
 sg13g2_decap_4 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_decap_8 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_17_415 ();
 sg13g2_decap_8 FILLER_17_422 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_fill_2 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_37 ();
 sg13g2_fill_2 FILLER_18_51 ();
 sg13g2_fill_1 FILLER_18_53 ();
 sg13g2_fill_2 FILLER_18_76 ();
 sg13g2_fill_1 FILLER_18_86 ();
 sg13g2_fill_1 FILLER_18_92 ();
 sg13g2_fill_2 FILLER_18_98 ();
 sg13g2_fill_2 FILLER_18_106 ();
 sg13g2_fill_2 FILLER_18_112 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_fill_2 FILLER_18_164 ();
 sg13g2_decap_4 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_189 ();
 sg13g2_fill_1 FILLER_18_195 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_4 FILLER_18_224 ();
 sg13g2_decap_4 FILLER_18_232 ();
 sg13g2_decap_4 FILLER_18_240 ();
 sg13g2_decap_4 FILLER_18_248 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_decap_4 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_4 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_decap_4 FILLER_18_376 ();
 sg13g2_fill_1 FILLER_18_392 ();
 sg13g2_fill_2 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_59 ();
 sg13g2_fill_2 FILLER_19_87 ();
 sg13g2_fill_2 FILLER_19_94 ();
 sg13g2_decap_4 FILLER_19_103 ();
 sg13g2_fill_2 FILLER_19_121 ();
 sg13g2_decap_4 FILLER_19_132 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_180 ();
 sg13g2_fill_1 FILLER_19_193 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_decap_4 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_243 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_4 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_283 ();
 sg13g2_decap_8 FILLER_19_290 ();
 sg13g2_fill_1 FILLER_19_297 ();
 sg13g2_fill_1 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_4 FILLER_19_375 ();
 sg13g2_fill_1 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_2 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_421 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_fill_1 FILLER_20_47 ();
 sg13g2_fill_2 FILLER_20_61 ();
 sg13g2_fill_2 FILLER_20_67 ();
 sg13g2_fill_1 FILLER_20_69 ();
 sg13g2_fill_2 FILLER_20_79 ();
 sg13g2_decap_4 FILLER_20_86 ();
 sg13g2_decap_4 FILLER_20_100 ();
 sg13g2_fill_2 FILLER_20_104 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_fill_2 FILLER_20_151 ();
 sg13g2_fill_1 FILLER_20_153 ();
 sg13g2_fill_2 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_fill_2 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_181 ();
 sg13g2_decap_8 FILLER_20_212 ();
 sg13g2_decap_8 FILLER_20_219 ();
 sg13g2_fill_2 FILLER_20_226 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_fill_1 FILLER_20_251 ();
 sg13g2_fill_1 FILLER_20_283 ();
 sg13g2_decap_4 FILLER_20_289 ();
 sg13g2_fill_1 FILLER_20_293 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_4 FILLER_20_312 ();
 sg13g2_decap_4 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_330 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_fill_2 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_386 ();
 sg13g2_fill_2 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_42 ();
 sg13g2_fill_2 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_66 ();
 sg13g2_decap_4 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_85 ();
 sg13g2_decap_8 FILLER_21_92 ();
 sg13g2_decap_4 FILLER_21_99 ();
 sg13g2_fill_2 FILLER_21_103 ();
 sg13g2_decap_8 FILLER_21_110 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_157 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_240 ();
 sg13g2_decap_4 FILLER_21_247 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_274 ();
 sg13g2_fill_1 FILLER_21_276 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_fill_1 FILLER_21_402 ();
 sg13g2_decap_4 FILLER_21_407 ();
 sg13g2_fill_2 FILLER_21_411 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_decap_4 FILLER_21_424 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_39 ();
 sg13g2_decap_4 FILLER_22_49 ();
 sg13g2_decap_4 FILLER_22_57 ();
 sg13g2_fill_1 FILLER_22_61 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_1 FILLER_22_76 ();
 sg13g2_decap_8 FILLER_22_103 ();
 sg13g2_decap_8 FILLER_22_110 ();
 sg13g2_decap_8 FILLER_22_125 ();
 sg13g2_decap_8 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_fill_2 FILLER_22_165 ();
 sg13g2_decap_4 FILLER_22_171 ();
 sg13g2_fill_2 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_186 ();
 sg13g2_fill_2 FILLER_22_190 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_decap_4 FILLER_22_247 ();
 sg13g2_fill_2 FILLER_22_251 ();
 sg13g2_decap_8 FILLER_22_292 ();
 sg13g2_decap_4 FILLER_22_299 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_4 FILLER_22_327 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_fill_1 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_16 ();
 sg13g2_decap_8 FILLER_23_23 ();
 sg13g2_decap_4 FILLER_23_30 ();
 sg13g2_fill_2 FILLER_23_34 ();
 sg13g2_fill_2 FILLER_23_65 ();
 sg13g2_decap_4 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_90 ();
 sg13g2_fill_2 FILLER_23_97 ();
 sg13g2_decap_4 FILLER_23_140 ();
 sg13g2_decap_4 FILLER_23_157 ();
 sg13g2_decap_4 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_169 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_decap_8 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_218 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_decap_4 FILLER_23_260 ();
 sg13g2_fill_1 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_269 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_fill_2 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_4 FILLER_23_392 ();
 sg13g2_fill_2 FILLER_23_396 ();
 sg13g2_fill_2 FILLER_23_409 ();
 sg13g2_decap_8 FILLER_23_415 ();
 sg13g2_decap_8 FILLER_23_422 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_31 ();
 sg13g2_decap_4 FILLER_24_38 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_55 ();
 sg13g2_decap_8 FILLER_24_79 ();
 sg13g2_fill_1 FILLER_24_86 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_131 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_decap_4 FILLER_24_190 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_4 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_4 FILLER_24_314 ();
 sg13g2_decap_8 FILLER_24_344 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_394 ();
 sg13g2_fill_1 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_decap_4 FILLER_25_31 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_59 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_fill_1 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_141 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_185 ();
 sg13g2_decap_8 FILLER_25_192 ();
 sg13g2_decap_8 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_216 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_4 FILLER_25_232 ();
 sg13g2_fill_1 FILLER_25_236 ();
 sg13g2_decap_4 FILLER_25_291 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_fill_2 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_13 ();
 sg13g2_decap_8 FILLER_26_20 ();
 sg13g2_decap_8 FILLER_26_27 ();
 sg13g2_fill_1 FILLER_26_34 ();
 sg13g2_fill_1 FILLER_26_40 ();
 sg13g2_decap_4 FILLER_26_80 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_fill_1 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_110 ();
 sg13g2_fill_1 FILLER_26_118 ();
 sg13g2_decap_4 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_137 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_decap_4 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_decap_8 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_decap_8 FILLER_26_222 ();
 sg13g2_decap_4 FILLER_26_229 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_fill_2 FILLER_26_241 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_fill_2 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_fill_2 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_fill_2 FILLER_26_376 ();
 sg13g2_decap_4 FILLER_26_386 ();
 sg13g2_fill_2 FILLER_26_390 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_20 ();
 sg13g2_decap_8 FILLER_27_27 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_decap_4 FILLER_27_42 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_108 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_fill_2 FILLER_27_135 ();
 sg13g2_fill_2 FILLER_27_142 ();
 sg13g2_decap_8 FILLER_27_148 ();
 sg13g2_decap_8 FILLER_27_155 ();
 sg13g2_fill_2 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_decap_8 FILLER_27_181 ();
 sg13g2_decap_8 FILLER_27_188 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_4 FILLER_27_275 ();
 sg13g2_decap_8 FILLER_27_293 ();
 sg13g2_decap_8 FILLER_27_304 ();
 sg13g2_decap_4 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_315 ();
 sg13g2_decap_4 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_371 ();
 sg13g2_fill_1 FILLER_27_403 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_4 FILLER_28_74 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_decap_4 FILLER_28_91 ();
 sg13g2_fill_2 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_decap_8 FILLER_28_110 ();
 sg13g2_decap_8 FILLER_28_117 ();
 sg13g2_decap_8 FILLER_28_124 ();
 sg13g2_fill_2 FILLER_28_131 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_fill_2 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_201 ();
 sg13g2_decap_4 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_decap_4 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_264 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_347 ();
 sg13g2_fill_1 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_fill_2 FILLER_28_374 ();
 sg13g2_decap_4 FILLER_28_384 ();
 sg13g2_fill_1 FILLER_28_392 ();
 sg13g2_fill_2 FILLER_28_408 ();
 sg13g2_fill_1 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_415 ();
 sg13g2_decap_8 FILLER_28_422 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_4 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_37 ();
 sg13g2_fill_2 FILLER_29_44 ();
 sg13g2_fill_1 FILLER_29_46 ();
 sg13g2_decap_8 FILLER_29_57 ();
 sg13g2_fill_2 FILLER_29_64 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_4 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_decap_8 FILLER_29_124 ();
 sg13g2_fill_2 FILLER_29_131 ();
 sg13g2_decap_8 FILLER_29_143 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_decap_4 FILLER_29_156 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_1 FILLER_29_165 ();
 sg13g2_decap_8 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_187 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_decap_4 FILLER_29_220 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_279 ();
 sg13g2_fill_1 FILLER_29_281 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_decap_8 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_344 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_52 ();
 sg13g2_fill_1 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_83 ();
 sg13g2_decap_8 FILLER_30_90 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_99 ();
 sg13g2_decap_4 FILLER_30_108 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_117 ();
 sg13g2_decap_4 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_128 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_216 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_decap_4 FILLER_30_245 ();
 sg13g2_decap_4 FILLER_30_253 ();
 sg13g2_fill_1 FILLER_30_257 ();
 sg13g2_decap_4 FILLER_30_298 ();
 sg13g2_fill_1 FILLER_30_302 ();
 sg13g2_decap_8 FILLER_30_307 ();
 sg13g2_decap_8 FILLER_30_314 ();
 sg13g2_decap_4 FILLER_30_321 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_fill_2 FILLER_30_359 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_fill_1 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_30_376 ();
 sg13g2_fill_1 FILLER_30_378 ();
 sg13g2_decap_4 FILLER_30_387 ();
 sg13g2_fill_1 FILLER_30_391 ();
 sg13g2_fill_2 FILLER_30_400 ();
 sg13g2_decap_4 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_410 ();
 sg13g2_decap_8 FILLER_30_415 ();
 sg13g2_decap_8 FILLER_30_422 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_59 ();
 sg13g2_decap_4 FILLER_31_66 ();
 sg13g2_fill_2 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_76 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_90 ();
 sg13g2_decap_4 FILLER_31_95 ();
 sg13g2_fill_1 FILLER_31_99 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_132 ();
 sg13g2_decap_4 FILLER_31_142 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_fill_1 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_fill_2 FILLER_31_194 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_decap_8 FILLER_31_243 ();
 sg13g2_decap_8 FILLER_31_250 ();
 sg13g2_decap_4 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_291 ();
 sg13g2_decap_4 FILLER_31_324 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_decap_4 FILLER_31_333 ();
 sg13g2_fill_2 FILLER_31_353 ();
 sg13g2_decap_4 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_32 ();
 sg13g2_decap_4 FILLER_32_37 ();
 sg13g2_fill_2 FILLER_32_45 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_fill_1 FILLER_32_99 ();
 sg13g2_decap_4 FILLER_32_117 ();
 sg13g2_fill_1 FILLER_32_121 ();
 sg13g2_fill_2 FILLER_32_127 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_2 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_202 ();
 sg13g2_decap_4 FILLER_32_216 ();
 sg13g2_decap_8 FILLER_32_225 ();
 sg13g2_decap_8 FILLER_32_232 ();
 sg13g2_decap_8 FILLER_32_239 ();
 sg13g2_decap_8 FILLER_32_246 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_fill_1 FILLER_32_264 ();
 sg13g2_fill_2 FILLER_32_275 ();
 sg13g2_decap_4 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_decap_4 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_373 ();
 sg13g2_decap_4 FILLER_32_379 ();
 sg13g2_fill_1 FILLER_32_383 ();
 sg13g2_decap_4 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_32_423 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_60 ();
 sg13g2_fill_1 FILLER_33_62 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_79 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_153 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_decap_4 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_decap_4 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_decap_4 FILLER_33_221 ();
 sg13g2_fill_2 FILLER_33_225 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_fill_1 FILLER_33_291 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_339 ();
 sg13g2_decap_8 FILLER_33_345 ();
 sg13g2_decap_4 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_1 FILLER_33_409 ();
 sg13g2_decap_8 FILLER_33_414 ();
 sg13g2_decap_8 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_fill_2 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_41 ();
 sg13g2_decap_4 FILLER_34_60 ();
 sg13g2_fill_1 FILLER_34_64 ();
 sg13g2_decap_4 FILLER_34_74 ();
 sg13g2_decap_8 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_99 ();
 sg13g2_decap_8 FILLER_34_131 ();
 sg13g2_decap_4 FILLER_34_138 ();
 sg13g2_decap_4 FILLER_34_146 ();
 sg13g2_decap_8 FILLER_34_165 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_fill_2 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_decap_4 FILLER_34_214 ();
 sg13g2_decap_4 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_fill_2 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_decap_8 FILLER_34_306 ();
 sg13g2_decap_8 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_326 ();
 sg13g2_fill_2 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_fill_1 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_45 ();
 sg13g2_fill_1 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_71 ();
 sg13g2_decap_4 FILLER_35_78 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_fill_2 FILLER_35_108 ();
 sg13g2_decap_4 FILLER_35_114 ();
 sg13g2_decap_4 FILLER_35_121 ();
 sg13g2_decap_4 FILLER_35_161 ();
 sg13g2_fill_1 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_201 ();
 sg13g2_fill_1 FILLER_35_203 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_fill_2 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_decap_4 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_fill_2 FILLER_35_427 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_20 ();
 sg13g2_decap_8 FILLER_36_27 ();
 sg13g2_decap_4 FILLER_36_34 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_44 ();
 sg13g2_decap_4 FILLER_36_53 ();
 sg13g2_fill_2 FILLER_36_61 ();
 sg13g2_fill_1 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_68 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_fill_2 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_127 ();
 sg13g2_decap_8 FILLER_36_138 ();
 sg13g2_fill_1 FILLER_36_145 ();
 sg13g2_decap_8 FILLER_36_155 ();
 sg13g2_decap_8 FILLER_36_162 ();
 sg13g2_decap_4 FILLER_36_169 ();
 sg13g2_fill_2 FILLER_36_173 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_decap_4 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_211 ();
 sg13g2_decap_4 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_decap_4 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_decap_4 FILLER_36_253 ();
 sg13g2_decap_4 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_decap_8 FILLER_36_279 ();
 sg13g2_decap_8 FILLER_36_286 ();
 sg13g2_fill_2 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_decap_8 FILLER_36_306 ();
 sg13g2_fill_2 FILLER_36_313 ();
 sg13g2_decap_4 FILLER_36_320 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_342 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_350 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_fill_1 FILLER_36_401 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_40 ();
 sg13g2_decap_4 FILLER_37_47 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_fill_2 FILLER_37_92 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_100 ();
 sg13g2_fill_1 FILLER_37_127 ();
 sg13g2_fill_2 FILLER_37_154 ();
 sg13g2_fill_1 FILLER_37_156 ();
 sg13g2_fill_2 FILLER_37_161 ();
 sg13g2_fill_2 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_230 ();
 sg13g2_decap_4 FILLER_37_237 ();
 sg13g2_fill_2 FILLER_37_241 ();
 sg13g2_fill_2 FILLER_37_269 ();
 sg13g2_fill_2 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_fill_2 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_342 ();
 sg13g2_decap_4 FILLER_37_347 ();
 sg13g2_fill_2 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_358 ();
 sg13g2_fill_1 FILLER_37_360 ();
 sg13g2_fill_2 FILLER_37_365 ();
 sg13g2_fill_1 FILLER_37_397 ();
 sg13g2_fill_1 FILLER_37_403 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_79 ();
 sg13g2_fill_1 FILLER_38_81 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_decap_4 FILLER_38_276 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_decap_4 FILLER_38_291 ();
 sg13g2_fill_2 FILLER_38_312 ();
 sg13g2_decap_8 FILLER_38_321 ();
 sg13g2_fill_2 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_fill_1 FILLER_38_376 ();
 sg13g2_fill_2 FILLER_38_390 ();
 sg13g2_decap_4 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_405 ();
 sg13g2_fill_1 FILLER_38_409 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_421 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
